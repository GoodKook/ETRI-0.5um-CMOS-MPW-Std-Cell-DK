VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 843.000 BY 834.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 819.300 840.450 821.700 ;
        RECT 8.700 815.400 10.500 819.300 ;
        RECT 16.200 812.400 18.000 819.300 ;
        RECT 34.500 809.400 36.300 819.300 ;
        RECT 49.800 815.400 51.600 819.300 ;
        RECT 57.000 812.400 58.800 819.300 ;
        RECT 64.500 815.400 66.300 819.300 ;
        RECT 85.500 812.400 87.300 819.300 ;
        RECT 97.800 815.400 99.600 819.300 ;
        RECT 103.800 815.400 105.600 819.300 ;
        RECT 110.700 812.400 112.500 819.300 ;
        RECT 133.800 814.200 135.600 819.300 ;
        RECT 154.500 812.400 156.300 819.300 ;
        RECT 169.500 812.400 171.300 819.300 ;
        RECT 189.300 812.400 191.100 819.300 ;
        RECT 214.500 809.400 216.300 819.300 ;
        RECT 225.000 812.400 226.800 819.300 ;
        RECT 232.500 815.400 234.300 819.300 ;
        RECT 245.700 809.400 247.500 819.300 ;
        RECT 269.400 814.200 271.200 819.300 ;
        RECT 287.400 815.400 289.200 819.300 ;
        RECT 310.800 814.200 312.600 819.300 ;
        RECT 328.800 814.200 330.600 819.300 ;
        RECT 344.700 815.400 346.500 819.300 ;
        RECT 352.200 812.400 354.000 819.300 ;
        RECT 359.700 809.400 361.500 819.300 ;
        RECT 391.500 809.400 393.300 819.300 ;
        RECT 404.700 815.400 406.500 819.300 ;
        RECT 412.200 812.400 414.000 819.300 ;
        RECT 433.500 809.400 435.300 819.300 ;
        RECT 443.700 815.400 445.500 819.300 ;
        RECT 451.200 812.400 453.000 819.300 ;
        RECT 462.000 812.400 463.800 819.300 ;
        RECT 469.500 815.400 471.300 819.300 ;
        RECT 479.400 815.400 481.200 819.300 ;
        RECT 499.800 814.200 501.600 819.300 ;
        RECT 515.400 814.200 517.200 819.300 ;
        RECT 533.700 809.400 535.500 819.300 ;
        RECT 552.000 812.400 553.800 819.300 ;
        RECT 559.500 815.400 561.300 819.300 ;
        RECT 575.400 814.200 577.200 819.300 ;
        RECT 604.500 809.400 606.300 819.300 ;
        RECT 615.000 812.400 616.800 819.300 ;
        RECT 622.500 815.400 624.300 819.300 ;
        RECT 635.700 812.400 637.500 819.300 ;
        RECT 658.500 812.400 660.300 819.300 ;
        RECT 679.500 812.400 681.300 819.300 ;
        RECT 687.000 812.400 688.800 819.300 ;
        RECT 694.500 815.400 696.300 819.300 ;
        RECT 709.800 815.400 711.600 819.300 ;
        RECT 715.800 815.400 717.600 819.300 ;
        RECT 722.700 812.400 724.500 819.300 ;
        RECT 740.400 814.200 742.200 819.300 ;
        RECT 761.400 814.200 763.200 819.300 ;
        RECT 779.700 809.400 781.500 819.300 ;
        RECT 808.500 809.400 810.300 819.300 ;
        RECT 816.000 812.400 817.800 819.300 ;
        RECT 823.500 815.400 825.300 819.300 ;
        RECT 13.800 743.700 15.600 748.800 ;
        RECT 23.400 743.700 25.200 747.600 ;
        RECT 38.400 743.700 40.200 748.800 ;
        RECT 59.700 743.700 61.500 747.600 ;
        RECT 67.200 743.700 69.000 750.600 ;
        RECT 74.700 743.700 76.500 753.600 ;
        RECT 95.700 743.700 97.500 753.600 ;
        RECT 113.700 743.700 115.500 750.600 ;
        RECT 128.700 743.700 130.500 750.600 ;
        RECT 147.000 743.700 148.800 750.600 ;
        RECT 155.400 743.700 157.200 750.600 ;
        RECT 173.700 743.700 175.500 747.600 ;
        RECT 181.200 743.700 183.000 750.600 ;
        RECT 188.700 743.700 190.500 753.600 ;
        RECT 217.800 743.700 219.600 748.800 ;
        RECT 235.800 743.700 237.600 748.800 ;
        RECT 259.500 743.700 261.300 753.600 ;
        RECT 272.700 743.700 274.500 747.600 ;
        RECT 280.200 743.700 282.000 750.600 ;
        RECT 291.000 743.700 292.800 750.600 ;
        RECT 298.500 743.700 300.300 747.600 ;
        RECT 319.500 743.700 321.300 753.600 ;
        RECT 337.500 743.700 339.300 753.600 ;
        RECT 358.500 743.700 360.300 753.600 ;
        RECT 370.800 743.700 372.600 747.600 ;
        RECT 383.700 743.700 385.500 747.600 ;
        RECT 391.200 743.700 393.000 750.600 ;
        RECT 409.500 743.700 411.300 753.600 ;
        RECT 416.400 743.700 418.200 747.600 ;
        RECT 436.800 743.700 438.600 750.600 ;
        RECT 445.200 743.700 447.000 750.600 ;
        RECT 452.700 743.700 454.500 750.600 ;
        RECT 470.400 743.700 472.200 748.800 ;
        RECT 496.500 743.700 498.300 753.600 ;
        RECT 506.700 743.700 508.500 747.600 ;
        RECT 514.200 743.700 516.000 750.600 ;
        RECT 524.700 743.700 526.500 753.600 ;
        RECT 553.500 743.700 555.300 750.600 ;
        RECT 568.800 743.700 570.600 748.800 ;
        RECT 578.400 743.700 580.200 747.600 ;
        RECT 591.000 743.700 592.800 750.600 ;
        RECT 599.400 743.700 601.200 750.600 ;
        RECT 616.800 743.700 618.600 747.600 ;
        RECT 634.500 743.700 636.300 750.600 ;
        RECT 649.500 743.700 651.300 750.600 ;
        RECT 659.400 743.700 661.200 747.600 ;
        RECT 665.400 743.700 667.200 747.600 ;
        RECT 674.700 743.700 676.500 750.600 ;
        RECT 700.800 743.700 702.600 748.800 ;
        RECT 713.400 743.700 715.200 748.800 ;
        RECT 732.000 743.700 733.800 750.600 ;
        RECT 739.500 743.700 741.300 747.600 ;
        RECT 755.400 743.700 757.200 748.800 ;
        RECT 784.500 743.700 786.300 753.600 ;
        RECT 795.000 743.700 796.800 750.600 ;
        RECT 802.500 743.700 804.300 747.600 ;
        RECT 818.400 743.700 820.200 748.800 ;
        RECT 831.450 743.700 840.450 819.300 ;
        RECT 0.600 741.300 840.450 743.700 ;
        RECT 19.500 731.400 21.300 741.300 ;
        RECT 30.000 734.400 31.800 741.300 ;
        RECT 37.500 737.400 39.300 741.300 ;
        RECT 61.500 731.400 63.300 741.300 ;
        RECT 82.500 731.400 84.300 741.300 ;
        RECT 93.000 734.400 94.800 741.300 ;
        RECT 100.500 737.400 102.300 741.300 ;
        RECT 118.800 736.200 120.600 741.300 ;
        RECT 135.300 734.400 137.100 741.300 ;
        RECT 154.500 734.400 156.300 741.300 ;
        RECT 175.800 736.200 177.600 741.300 ;
        RECT 188.400 736.200 190.200 741.300 ;
        RECT 214.500 731.400 216.300 741.300 ;
        RECT 221.700 731.400 223.500 741.300 ;
        RECT 240.000 734.400 241.800 741.300 ;
        RECT 247.500 737.400 249.300 741.300 ;
        RECT 263.400 736.200 265.200 741.300 ;
        RECT 284.700 737.400 286.500 741.300 ;
        RECT 292.200 734.400 294.000 741.300 ;
        RECT 302.700 731.400 304.500 741.300 ;
        RECT 330.300 734.400 332.100 741.300 ;
        RECT 344.700 734.400 346.500 741.300 ;
        RECT 373.500 731.400 375.300 741.300 ;
        RECT 394.500 731.400 396.300 741.300 ;
        RECT 407.400 736.200 409.200 741.300 ;
        RECT 430.500 734.400 432.300 741.300 ;
        RECT 444.300 734.400 446.100 741.300 ;
        RECT 463.800 734.400 465.600 741.300 ;
        RECT 472.200 734.400 474.000 741.300 ;
        RECT 486.900 734.400 488.700 741.300 ;
        RECT 507.300 734.400 509.100 741.300 ;
        RECT 522.900 734.400 524.700 741.300 ;
        RECT 544.800 734.400 546.600 741.300 ;
        RECT 553.200 734.400 555.000 741.300 ;
        RECT 567.900 734.400 569.700 741.300 ;
        RECT 584.700 734.400 586.500 741.300 ;
        RECT 602.700 737.400 604.500 741.300 ;
        RECT 610.200 734.400 612.000 741.300 ;
        RECT 624.900 734.400 626.700 741.300 ;
        RECT 643.800 737.400 645.600 741.300 ;
        RECT 649.800 737.400 651.600 741.300 ;
        RECT 659.700 734.400 661.500 741.300 ;
        RECT 678.000 734.400 679.800 741.300 ;
        RECT 685.500 737.400 687.300 741.300 ;
        RECT 695.400 737.400 697.200 741.300 ;
        RECT 715.800 737.400 717.600 741.300 ;
        RECT 722.400 737.400 724.200 741.300 ;
        RECT 748.500 731.400 750.300 741.300 ;
        RECT 758.700 731.400 760.500 741.300 ;
        RECT 779.700 731.400 781.500 741.300 ;
        RECT 805.500 734.400 807.300 741.300 ;
        RECT 823.500 731.400 825.300 741.300 ;
        RECT 16.500 665.700 18.300 672.600 ;
        RECT 23.700 665.700 25.500 675.600 ;
        RECT 42.000 665.700 43.800 672.600 ;
        RECT 49.500 665.700 51.300 669.600 ;
        RECT 65.400 665.700 67.200 670.800 ;
        RECT 86.700 665.700 88.500 669.600 ;
        RECT 94.200 665.700 96.000 672.600 ;
        RECT 104.400 665.700 106.200 669.600 ;
        RECT 123.300 665.700 125.100 672.600 ;
        RECT 134.700 665.700 136.500 672.600 ;
        RECT 163.500 665.700 165.300 675.600 ;
        RECT 184.500 665.700 186.300 675.600 ;
        RECT 192.000 665.700 193.800 672.600 ;
        RECT 199.500 665.700 201.300 669.600 ;
        RECT 215.700 665.700 217.500 669.600 ;
        RECT 223.200 665.700 225.000 672.600 ;
        RECT 241.500 665.700 243.300 675.600 ;
        RECT 251.400 665.700 253.200 669.600 ;
        RECT 264.000 665.700 265.800 672.600 ;
        RECT 272.400 665.700 274.200 672.600 ;
        RECT 287.400 665.700 289.200 669.600 ;
        RECT 293.400 665.700 295.200 669.600 ;
        RECT 302.700 665.700 304.500 675.600 ;
        RECT 328.500 665.700 330.300 672.600 ;
        RECT 346.500 665.700 348.300 672.600 ;
        RECT 356.700 665.700 358.500 669.600 ;
        RECT 364.200 665.700 366.000 672.600 ;
        RECT 385.500 665.700 387.300 675.600 ;
        RECT 398.400 665.700 400.200 670.800 ;
        RECT 419.400 665.700 421.200 670.800 ;
        RECT 448.500 665.700 450.300 675.600 ;
        RECT 463.500 665.700 465.300 672.600 ;
        RECT 473.700 665.700 475.500 672.600 ;
        RECT 485.400 665.700 487.200 672.600 ;
        RECT 502.500 665.700 504.300 672.600 ;
        RECT 518.400 665.700 520.200 670.800 ;
        RECT 541.800 665.700 543.600 672.600 ;
        RECT 550.200 665.700 552.000 672.600 ;
        RECT 560.700 665.700 562.500 672.600 ;
        RECT 580.800 665.700 582.600 669.600 ;
        RECT 593.400 665.700 595.200 670.800 ;
        RECT 616.800 665.700 618.600 669.600 ;
        RECT 626.400 665.700 628.200 670.800 ;
        RECT 652.500 665.700 654.300 675.600 ;
        RECT 659.700 665.700 661.500 675.600 ;
        RECT 680.700 665.700 682.500 675.600 ;
        RECT 701.700 665.700 703.500 675.600 ;
        RECT 719.700 665.700 721.500 675.600 ;
        RECT 741.000 665.700 742.800 672.600 ;
        RECT 749.400 665.700 751.200 672.600 ;
        RECT 763.800 665.700 765.600 669.600 ;
        RECT 769.800 665.700 771.600 669.600 ;
        RECT 782.400 665.700 784.200 670.800 ;
        RECT 808.500 665.700 810.300 672.600 ;
        RECT 816.000 665.700 817.800 672.600 ;
        RECT 823.500 665.700 825.300 669.600 ;
        RECT 831.450 665.700 840.450 741.300 ;
        RECT 0.600 663.300 840.450 665.700 ;
        RECT 16.500 656.400 18.300 663.300 ;
        RECT 37.500 653.400 39.300 663.300 ;
        RECT 47.700 653.400 49.500 663.300 ;
        RECT 65.400 659.400 67.200 663.300 ;
        RECT 81.000 656.400 82.800 663.300 ;
        RECT 88.500 659.400 90.300 663.300 ;
        RECT 106.800 659.400 108.600 663.300 ;
        RECT 124.800 658.200 126.600 663.300 ;
        RECT 139.800 659.400 141.600 663.300 ;
        RECT 145.800 659.400 147.600 663.300 ;
        RECT 160.500 656.400 162.300 663.300 ;
        RECT 175.500 656.400 177.300 663.300 ;
        RECT 190.500 656.400 192.300 663.300 ;
        RECT 211.800 658.200 213.600 663.300 ;
        RECT 232.800 658.200 234.600 663.300 ;
        RECT 250.800 658.200 252.600 663.300 ;
        RECT 271.500 656.400 273.300 663.300 ;
        RECT 289.800 658.200 291.600 663.300 ;
        RECT 302.400 659.400 304.200 663.300 ;
        RECT 314.700 653.400 316.500 663.300 ;
        RECT 340.800 659.400 342.600 663.300 ;
        RECT 347.700 656.400 349.500 663.300 ;
        RECT 367.800 656.400 369.600 663.300 ;
        RECT 382.500 656.400 384.300 663.300 ;
        RECT 397.800 659.400 399.600 663.300 ;
        RECT 407.700 653.400 409.500 663.300 ;
        RECT 439.500 653.400 441.300 663.300 ;
        RECT 446.700 656.400 448.500 663.300 ;
        RECT 469.800 656.400 471.600 663.300 ;
        RECT 478.200 656.400 480.000 663.300 ;
        RECT 493.800 659.400 495.600 663.300 ;
        RECT 500.400 659.400 502.200 663.300 ;
        RECT 523.800 657.900 525.600 663.300 ;
        RECT 536.400 659.400 538.200 663.300 ;
        RECT 542.400 659.400 544.200 663.300 ;
        RECT 552.000 656.400 553.800 663.300 ;
        RECT 559.500 659.400 561.300 663.300 ;
        RECT 572.700 653.400 574.500 663.300 ;
        RECT 590.700 656.400 592.500 663.300 ;
        RECT 611.400 658.200 613.200 663.300 ;
        RECT 626.400 659.400 628.200 663.300 ;
        RECT 641.700 656.400 643.500 663.300 ;
        RECT 664.800 659.400 666.600 663.300 ;
        RECT 677.400 658.200 679.200 663.300 ;
        RECT 695.400 658.200 697.200 663.300 ;
        RECT 718.800 659.400 720.600 663.300 ;
        RECT 728.700 653.400 730.500 663.300 ;
        RECT 760.500 653.400 762.300 663.300 ;
        RECT 775.500 656.400 777.300 663.300 ;
        RECT 784.800 659.400 786.600 663.300 ;
        RECT 790.800 659.400 792.600 663.300 ;
        RECT 805.500 656.400 807.300 663.300 ;
        RECT 815.700 653.400 817.500 663.300 ;
        RECT 13.500 587.700 15.300 594.600 ;
        RECT 34.500 587.700 36.300 597.600 ;
        RECT 49.800 587.700 51.600 591.600 ;
        RECT 70.500 587.700 72.300 597.600 ;
        RECT 88.800 587.700 90.600 592.800 ;
        RECT 101.700 587.700 103.500 597.600 ;
        RECT 122.700 587.700 124.500 594.600 ;
        RECT 140.400 587.700 142.200 592.800 ;
        RECT 156.000 587.700 157.800 594.600 ;
        RECT 164.400 587.700 166.200 594.600 ;
        RECT 180.000 587.700 181.800 594.600 ;
        RECT 188.400 587.700 190.200 594.600 ;
        RECT 200.400 587.700 202.200 594.600 ;
        RECT 215.700 587.700 217.500 597.600 ;
        RECT 241.800 587.700 243.600 591.600 ;
        RECT 248.700 587.700 250.500 597.600 ;
        RECT 269.700 587.700 271.500 594.600 ;
        RECT 295.800 587.700 297.600 592.800 ;
        RECT 315.300 587.700 317.100 594.600 ;
        RECT 326.700 587.700 328.500 594.600 ;
        RECT 352.500 587.700 354.300 597.600 ;
        RECT 362.700 587.700 364.500 594.600 ;
        RECT 380.400 587.700 382.200 592.800 ;
        RECT 405.300 587.700 407.100 594.600 ;
        RECT 419.400 587.700 421.200 592.800 ;
        RECT 434.700 587.700 436.500 594.600 ;
        RECT 452.400 587.700 454.200 592.800 ;
        RECT 477.300 587.700 479.100 594.600 ;
        RECT 499.500 587.700 501.300 594.600 ;
        RECT 509.400 587.700 511.200 591.600 ;
        RECT 515.400 587.700 517.200 591.600 ;
        RECT 527.400 587.700 529.200 592.800 ;
        RECT 553.500 587.700 555.300 594.600 ;
        RECT 563.700 587.700 565.500 597.600 ;
        RECT 586.800 587.700 588.600 594.600 ;
        RECT 601.500 587.700 603.300 594.600 ;
        RECT 619.500 587.700 621.300 594.600 ;
        RECT 629.700 587.700 631.500 597.600 ;
        RECT 648.000 587.700 649.800 594.600 ;
        RECT 655.500 587.700 657.300 591.600 ;
        RECT 669.000 587.700 670.800 594.600 ;
        RECT 676.500 587.700 678.300 591.600 ;
        RECT 689.700 587.700 691.500 597.600 ;
        RECT 713.700 587.700 715.500 591.600 ;
        RECT 721.200 587.700 723.000 594.600 ;
        RECT 733.800 587.700 735.600 591.600 ;
        RECT 751.800 587.700 753.600 592.800 ;
        RECT 766.800 587.700 768.600 591.600 ;
        RECT 773.400 587.700 775.200 591.600 ;
        RECT 788.700 587.700 790.500 597.600 ;
        RECT 817.500 587.700 819.300 597.600 ;
        RECT 831.450 587.700 840.450 663.300 ;
        RECT 0.600 585.300 840.450 587.700 ;
        RECT 8.700 581.400 10.500 585.300 ;
        RECT 16.200 578.400 18.000 585.300 ;
        RECT 34.500 575.400 36.300 585.300 ;
        RECT 44.700 581.400 46.500 585.300 ;
        RECT 52.200 578.400 54.000 585.300 ;
        RECT 67.500 578.400 69.300 585.300 ;
        RECT 80.700 581.400 82.500 585.300 ;
        RECT 88.200 578.400 90.000 585.300 ;
        RECT 109.500 575.400 111.300 585.300 ;
        RECT 123.300 578.400 125.100 585.300 ;
        RECT 142.500 578.400 144.300 585.300 ;
        RECT 157.500 578.400 159.300 585.300 ;
        RECT 174.900 578.400 176.700 585.300 ;
        RECT 196.500 578.400 198.300 585.300 ;
        RECT 209.400 580.200 211.200 585.300 ;
        RECT 227.700 578.400 229.500 585.300 ;
        RECT 253.800 580.200 255.600 585.300 ;
        RECT 263.400 578.400 265.200 585.300 ;
        RECT 275.400 578.400 277.200 585.300 ;
        RECT 292.800 578.400 294.600 585.300 ;
        RECT 306.900 578.400 308.700 585.300 ;
        RECT 331.800 580.200 333.600 585.300 ;
        RECT 352.500 578.400 354.300 585.300 ;
        RECT 367.800 580.200 369.600 585.300 ;
        RECT 387.300 578.400 389.100 585.300 ;
        RECT 406.800 580.200 408.600 585.300 ;
        RECT 424.500 578.400 426.300 585.300 ;
        RECT 442.800 580.200 444.600 585.300 ;
        RECT 460.800 578.400 462.600 585.300 ;
        RECT 478.500 578.400 480.300 585.300 ;
        RECT 491.400 580.200 493.200 585.300 ;
        RECT 514.800 578.400 516.600 585.300 ;
        RECT 529.800 580.200 531.600 585.300 ;
        RECT 550.800 580.200 552.600 585.300 ;
        RECT 566.400 580.200 568.200 585.300 ;
        RECT 592.800 580.200 594.600 585.300 ;
        RECT 602.400 584.400 603.600 585.300 ;
        RECT 602.400 581.400 604.200 584.400 ;
        RECT 608.400 581.400 610.200 585.300 ;
        RECT 623.400 580.200 625.200 585.300 ;
        RECT 638.700 578.400 640.500 585.300 ;
        RECT 659.400 580.200 661.200 585.300 ;
        RECT 680.700 578.400 682.500 585.300 ;
        RECT 692.700 578.400 694.500 585.300 ;
        RECT 712.800 581.400 714.600 585.300 ;
        RECT 718.800 581.400 720.600 585.300 ;
        RECT 729.900 578.400 731.700 585.300 ;
        RECT 751.800 581.400 753.600 585.300 ;
        RECT 761.400 581.400 763.200 585.300 ;
        RECT 776.400 581.400 778.200 585.300 ;
        RECT 782.400 581.400 784.200 585.300 ;
        RECT 791.400 581.400 793.200 585.300 ;
        RECT 797.400 581.400 799.200 585.300 ;
        RECT 809.400 581.400 811.200 585.300 ;
        RECT 815.400 581.400 817.200 585.300 ;
        RECT 11.700 509.700 13.500 513.600 ;
        RECT 19.200 509.700 21.000 516.600 ;
        RECT 29.700 509.700 31.500 519.600 ;
        RECT 52.800 509.700 54.600 513.600 ;
        RECT 70.800 509.700 72.600 514.800 ;
        RECT 83.400 509.700 85.200 514.800 ;
        RECT 109.800 509.700 111.600 514.800 ;
        RECT 122.400 509.700 124.200 514.800 ;
        RECT 148.500 509.700 150.300 516.600 ;
        RECT 161.700 509.700 163.500 513.600 ;
        RECT 169.200 509.700 171.000 516.600 ;
        RECT 187.800 509.700 189.600 514.800 ;
        RECT 200.700 509.700 202.500 516.600 ;
        RECT 221.400 509.700 223.200 514.800 ;
        RECT 241.500 509.700 243.300 516.600 ;
        RECT 254.400 509.700 256.200 514.800 ;
        RECT 277.800 509.700 279.600 514.800 ;
        RECT 295.500 509.700 297.300 516.600 ;
        RECT 302.700 509.700 304.500 516.600 ;
        RECT 320.700 509.700 322.500 516.600 ;
        RECT 346.800 509.700 348.600 514.800 ;
        RECT 367.500 509.700 369.300 516.600 ;
        RECT 380.400 509.700 382.200 514.800 ;
        RECT 396.150 509.700 397.950 513.600 ;
        RECT 405.450 509.700 407.250 513.600 ;
        RECT 412.350 509.700 414.150 513.600 ;
        RECT 421.350 509.700 423.150 513.600 ;
        RECT 434.700 509.700 436.500 516.600 ;
        RECT 457.800 509.700 459.600 514.800 ;
        RECT 468.150 509.700 469.950 513.600 ;
        RECT 477.450 509.700 479.250 513.600 ;
        RECT 484.350 509.700 486.150 513.600 ;
        RECT 493.350 509.700 495.150 513.600 ;
        RECT 504.150 509.700 505.950 513.600 ;
        RECT 513.450 509.700 515.250 513.600 ;
        RECT 520.350 509.700 522.150 513.600 ;
        RECT 529.350 509.700 531.150 513.600 ;
        RECT 550.500 509.700 552.300 516.600 ;
        RECT 561.900 509.700 563.700 516.600 ;
        RECT 575.700 509.700 577.500 519.600 ;
        RECT 593.700 509.700 595.500 516.600 ;
        RECT 608.700 509.700 610.500 516.600 ;
        RECT 629.400 509.700 631.200 514.800 ;
        RECT 651.900 509.700 653.700 516.600 ;
        RECT 676.500 509.700 678.300 516.600 ;
        RECT 683.400 510.600 685.200 513.600 ;
        RECT 683.400 509.700 684.600 510.600 ;
        RECT 689.400 509.700 691.200 513.600 ;
        RECT 707.700 509.700 709.500 513.600 ;
        RECT 715.200 509.700 717.000 516.600 ;
        RECT 724.800 509.700 726.600 513.600 ;
        RECT 730.800 509.700 732.600 513.600 ;
        RECT 740.400 509.700 742.200 514.800 ;
        RECT 759.000 509.700 760.800 516.600 ;
        RECT 766.500 509.700 768.300 513.600 ;
        RECT 776.700 509.700 778.500 516.600 ;
        RECT 805.500 509.700 807.300 519.600 ;
        RECT 818.700 509.700 820.500 516.600 ;
        RECT 831.450 509.700 840.450 585.300 ;
        RECT 0.600 507.300 840.450 509.700 ;
        RECT 8.400 502.200 10.200 507.300 ;
        RECT 31.800 503.400 33.600 507.300 ;
        RECT 38.700 497.400 40.500 507.300 ;
        RECT 64.800 503.400 66.600 507.300 ;
        RECT 74.700 503.400 76.500 507.300 ;
        RECT 82.200 500.400 84.000 507.300 ;
        RECT 103.500 497.400 105.300 507.300 ;
        RECT 116.700 503.400 118.500 507.300 ;
        RECT 124.200 500.400 126.000 507.300 ;
        RECT 131.400 503.400 133.200 507.300 ;
        RECT 146.400 503.400 148.200 507.300 ;
        RECT 163.800 503.400 165.600 507.300 ;
        RECT 169.800 503.400 171.600 507.300 ;
        RECT 179.700 500.400 181.500 507.300 ;
        RECT 208.500 497.400 210.300 507.300 ;
        RECT 218.700 500.400 220.500 507.300 ;
        RECT 240.300 500.400 242.100 507.300 ;
        RECT 254.400 503.400 256.200 507.300 ;
        RECT 271.800 503.400 273.600 507.300 ;
        RECT 289.500 497.400 291.300 507.300 ;
        RECT 299.700 500.400 301.500 507.300 ;
        RECT 317.400 502.200 319.200 507.300 ;
        RECT 332.700 500.400 334.500 507.300 ;
        RECT 347.850 503.400 349.650 507.300 ;
        RECT 356.850 503.400 358.650 507.300 ;
        RECT 363.750 503.400 365.550 507.300 ;
        RECT 373.050 503.400 374.850 507.300 ;
        RECT 389.400 502.200 391.200 507.300 ;
        RECT 412.500 500.400 414.300 507.300 ;
        RECT 427.500 500.400 429.300 507.300 ;
        RECT 437.700 500.400 439.500 507.300 ;
        RECT 460.500 500.400 462.300 507.300 ;
        RECT 475.800 502.200 477.600 507.300 ;
        RECT 496.800 502.200 498.600 507.300 ;
        RECT 512.400 502.200 514.200 507.300 ;
        RECT 527.400 503.400 529.200 507.300 ;
        RECT 533.400 503.400 535.200 507.300 ;
        RECT 543.000 500.400 544.800 507.300 ;
        RECT 550.500 503.400 552.300 507.300 ;
        RECT 560.400 503.400 562.200 507.300 ;
        RECT 566.400 503.400 568.200 507.300 ;
        RECT 578.400 503.400 580.200 507.300 ;
        RECT 601.500 500.400 603.300 507.300 ;
        RECT 616.800 503.400 618.600 507.300 ;
        RECT 623.700 497.400 625.500 507.300 ;
        RECT 649.800 503.400 651.600 507.300 ;
        RECT 659.400 502.200 661.200 507.300 ;
        RECT 677.400 502.200 679.200 507.300 ;
        RECT 703.500 497.400 705.300 507.300 ;
        RECT 716.400 502.200 718.200 507.300 ;
        RECT 739.800 503.400 741.600 507.300 ;
        RECT 749.700 500.400 751.500 507.300 ;
        RECT 770.400 502.200 772.200 507.300 ;
        RECT 793.500 500.400 795.300 507.300 ;
        RECT 811.500 497.400 813.300 507.300 ;
        RECT 821.400 503.400 823.200 507.300 ;
        RECT 16.500 431.700 18.300 441.600 ;
        RECT 24.000 431.700 25.800 438.600 ;
        RECT 31.500 431.700 33.300 435.600 ;
        RECT 52.800 431.700 54.600 436.800 ;
        RECT 73.500 431.700 75.300 441.600 ;
        RECT 94.500 431.700 96.300 441.600 ;
        RECT 112.800 431.700 114.600 436.800 ;
        RECT 128.400 431.700 130.200 436.800 ;
        RECT 151.800 431.700 153.600 435.600 ;
        RECT 166.800 431.700 168.600 436.800 ;
        RECT 176.400 431.700 178.200 435.600 ;
        RECT 182.400 431.700 184.200 435.600 ;
        RECT 194.700 431.700 196.500 438.600 ;
        RECT 212.700 431.700 214.500 438.600 ;
        RECT 231.000 431.700 232.800 438.600 ;
        RECT 239.400 431.700 241.200 438.600 ;
        RECT 256.800 431.700 258.600 435.600 ;
        RECT 267.900 431.700 269.700 438.600 ;
        RECT 287.700 431.700 289.500 435.600 ;
        RECT 295.200 431.700 297.000 438.600 ;
        RECT 305.700 431.700 307.500 441.600 ;
        RECT 326.400 431.700 328.200 436.800 ;
        RECT 341.850 431.700 343.650 435.600 ;
        RECT 350.850 431.700 352.650 435.600 ;
        RECT 357.750 431.700 359.550 435.600 ;
        RECT 367.050 431.700 368.850 435.600 ;
        RECT 380.700 431.700 382.500 438.600 ;
        RECT 393.150 431.700 394.950 435.600 ;
        RECT 402.450 431.700 404.250 435.600 ;
        RECT 409.350 431.700 411.150 435.600 ;
        RECT 418.350 431.700 420.150 435.600 ;
        RECT 434.700 431.700 436.500 438.600 ;
        RECT 447.150 431.700 448.950 435.600 ;
        RECT 456.450 431.700 458.250 435.600 ;
        RECT 463.350 431.700 465.150 435.600 ;
        RECT 472.350 431.700 474.150 435.600 ;
        RECT 493.500 431.700 495.300 438.600 ;
        RECT 506.400 431.700 508.200 436.800 ;
        RECT 521.400 431.700 523.200 438.600 ;
        RECT 534.150 431.700 535.950 435.600 ;
        RECT 543.450 431.700 545.250 435.600 ;
        RECT 550.350 431.700 552.150 435.600 ;
        RECT 559.350 431.700 561.150 435.600 ;
        RECT 575.400 431.700 577.200 436.800 ;
        RECT 593.400 431.700 595.200 438.600 ;
        RECT 599.400 431.700 601.200 438.600 ;
        RECT 605.400 431.700 607.200 438.600 ;
        RECT 611.400 431.700 613.200 438.600 ;
        RECT 617.400 431.700 619.200 438.600 ;
        RECT 637.800 431.700 639.600 436.800 ;
        RECT 655.800 431.700 657.600 435.600 ;
        RECT 662.700 431.700 664.500 438.600 ;
        RECT 680.700 431.700 682.500 438.600 ;
        RECT 695.400 432.600 697.200 435.600 ;
        RECT 695.400 431.700 696.600 432.600 ;
        RECT 701.400 431.700 703.200 435.600 ;
        RECT 716.400 431.700 718.200 435.600 ;
        RECT 731.400 431.700 733.200 435.600 ;
        RECT 737.400 431.700 739.200 435.600 ;
        RECT 748.800 431.700 750.600 435.600 ;
        RECT 754.800 431.700 756.600 435.600 ;
        RECT 762.000 431.700 763.800 438.600 ;
        RECT 769.500 431.700 771.300 435.600 ;
        RECT 782.400 431.700 784.200 435.600 ;
        RECT 797.700 431.700 799.500 441.600 ;
        RECT 821.700 431.700 823.500 438.600 ;
        RECT 831.450 431.700 840.450 507.300 ;
        RECT 0.600 429.300 840.450 431.700 ;
        RECT 13.800 425.400 15.600 429.300 ;
        RECT 23.700 425.400 25.500 429.300 ;
        RECT 31.200 422.400 33.000 429.300 ;
        RECT 49.500 419.400 51.300 429.300 ;
        RECT 64.800 422.400 66.600 429.300 ;
        RECT 73.200 422.400 75.000 429.300 ;
        RECT 80.700 422.400 82.500 429.300 ;
        RECT 106.500 419.400 108.300 429.300 ;
        RECT 116.700 425.400 118.500 429.300 ;
        RECT 124.200 422.400 126.000 429.300 ;
        RECT 139.800 425.400 141.600 429.300 ;
        RECT 154.800 424.200 156.600 429.300 ;
        RECT 166.800 425.400 168.600 429.300 ;
        RECT 172.800 425.400 174.600 429.300 ;
        RECT 179.700 422.400 181.500 429.300 ;
        RECT 205.800 424.200 207.600 429.300 ;
        RECT 218.400 425.400 220.200 429.300 ;
        RECT 224.400 425.400 226.200 429.300 ;
        RECT 233.400 425.400 235.200 429.300 ;
        RECT 248.400 424.200 250.200 429.300 ;
        RECT 274.800 424.200 276.600 429.300 ;
        RECT 287.400 425.400 289.200 429.300 ;
        RECT 293.400 425.400 295.200 429.300 ;
        RECT 305.400 424.200 307.200 429.300 ;
        RECT 323.700 422.400 325.500 429.300 ;
        RECT 339.150 425.400 340.950 429.300 ;
        RECT 348.450 425.400 350.250 429.300 ;
        RECT 355.350 425.400 357.150 429.300 ;
        RECT 364.350 425.400 366.150 429.300 ;
        RECT 376.800 422.400 378.600 429.300 ;
        RECT 382.800 422.400 384.600 429.300 ;
        RECT 388.800 422.400 390.600 429.300 ;
        RECT 394.800 422.400 396.600 429.300 ;
        RECT 400.800 422.400 402.600 429.300 ;
        RECT 407.700 422.400 409.500 429.300 ;
        RECT 433.800 424.200 435.600 429.300 ;
        RECT 451.500 422.400 453.300 429.300 ;
        RECT 466.500 422.400 468.300 429.300 ;
        RECT 487.800 424.200 489.600 429.300 ;
        RECT 498.150 425.400 499.950 429.300 ;
        RECT 507.450 425.400 509.250 429.300 ;
        RECT 514.350 425.400 516.150 429.300 ;
        RECT 523.350 425.400 525.150 429.300 ;
        RECT 541.800 425.400 543.600 429.300 ;
        RECT 548.400 425.400 550.200 429.300 ;
        RECT 554.400 425.400 556.200 429.300 ;
        RECT 571.800 425.400 573.600 429.300 ;
        RECT 581.400 425.400 583.200 429.300 ;
        RECT 587.400 425.400 589.200 429.300 ;
        RECT 597.150 425.400 598.950 429.300 ;
        RECT 606.450 425.400 608.250 429.300 ;
        RECT 613.350 425.400 615.150 429.300 ;
        RECT 622.350 425.400 624.150 429.300 ;
        RECT 643.800 423.900 645.600 429.300 ;
        RECT 661.800 425.400 663.600 429.300 ;
        RECT 668.850 425.400 670.650 429.300 ;
        RECT 677.850 425.400 679.650 429.300 ;
        RECT 684.750 425.400 686.550 429.300 ;
        RECT 694.050 425.400 695.850 429.300 ;
        RECT 715.800 424.200 717.600 429.300 ;
        RECT 733.800 425.400 735.600 429.300 ;
        RECT 748.800 422.400 750.600 429.300 ;
        RECT 757.200 422.400 759.000 429.300 ;
        RECT 765.150 425.400 766.950 429.300 ;
        RECT 774.450 425.400 776.250 429.300 ;
        RECT 781.350 425.400 783.150 429.300 ;
        RECT 790.350 425.400 792.150 429.300 ;
        RECT 803.400 425.400 805.200 429.300 ;
        RECT 818.700 422.400 820.500 429.300 ;
        RECT 11.700 353.700 13.500 357.600 ;
        RECT 19.200 353.700 21.000 360.600 ;
        RECT 40.500 353.700 42.300 363.600 ;
        RECT 49.800 353.700 51.600 357.600 ;
        RECT 55.800 353.700 57.600 357.600 ;
        RECT 67.800 353.700 69.600 357.600 ;
        RECT 80.700 353.700 82.500 357.600 ;
        RECT 88.200 353.700 90.000 360.600 ;
        RECT 109.500 353.700 111.300 363.600 ;
        RECT 119.400 353.700 121.200 357.600 ;
        RECT 142.500 353.700 144.300 363.600 ;
        RECT 155.700 353.700 157.500 360.600 ;
        RECT 181.500 353.700 183.300 363.600 ;
        RECT 199.800 353.700 201.600 358.800 ;
        RECT 223.800 353.700 225.600 359.100 ;
        RECT 241.800 353.700 243.600 358.800 ;
        RECT 253.800 353.700 255.600 360.600 ;
        RECT 259.800 353.700 261.600 360.600 ;
        RECT 265.800 353.700 267.600 360.600 ;
        RECT 271.800 353.700 273.600 360.600 ;
        RECT 277.800 353.700 279.600 360.600 ;
        RECT 286.800 353.700 288.600 357.600 ;
        RECT 292.800 353.700 294.600 357.600 ;
        RECT 299.850 353.700 301.650 357.600 ;
        RECT 308.850 353.700 310.650 357.600 ;
        RECT 315.750 353.700 317.550 357.600 ;
        RECT 325.050 353.700 326.850 357.600 ;
        RECT 341.700 353.700 343.500 357.600 ;
        RECT 349.200 353.700 351.000 360.600 ;
        RECT 356.400 353.700 358.200 360.600 ;
        RECT 362.400 353.700 364.200 360.600 ;
        RECT 368.400 353.700 370.200 360.600 ;
        RECT 374.400 353.700 376.200 360.600 ;
        RECT 380.400 353.700 382.200 360.600 ;
        RECT 390.150 353.700 391.950 357.600 ;
        RECT 399.450 353.700 401.250 357.600 ;
        RECT 406.350 353.700 408.150 357.600 ;
        RECT 415.350 353.700 417.150 357.600 ;
        RECT 428.700 353.700 430.500 357.600 ;
        RECT 436.200 353.700 438.000 360.600 ;
        RECT 446.400 353.700 448.200 357.600 ;
        RECT 452.400 353.700 454.200 357.600 ;
        RECT 462.000 353.700 463.800 360.600 ;
        RECT 469.500 353.700 471.300 357.600 ;
        RECT 480.150 353.700 481.950 357.600 ;
        RECT 489.450 353.700 491.250 357.600 ;
        RECT 496.350 353.700 498.150 357.600 ;
        RECT 505.350 353.700 507.150 357.600 ;
        RECT 516.150 353.700 517.950 357.600 ;
        RECT 525.450 353.700 527.250 357.600 ;
        RECT 532.350 353.700 534.150 357.600 ;
        RECT 541.350 353.700 543.150 357.600 ;
        RECT 551.400 353.700 553.200 357.600 ;
        RECT 557.400 353.700 559.200 357.600 ;
        RECT 574.800 353.700 576.600 357.600 ;
        RECT 581.850 353.700 583.650 357.600 ;
        RECT 590.850 353.700 592.650 357.600 ;
        RECT 597.750 353.700 599.550 357.600 ;
        RECT 607.050 353.700 608.850 357.600 ;
        RECT 625.800 353.700 627.600 358.800 ;
        RECT 635.400 353.700 637.200 357.600 ;
        RECT 647.400 353.700 649.200 357.600 ;
        RECT 653.400 353.700 655.200 357.600 ;
        RECT 665.400 353.700 667.200 357.600 ;
        RECT 671.400 353.700 673.200 357.600 ;
        RECT 683.400 353.700 685.200 359.100 ;
        RECT 704.700 353.700 706.500 357.600 ;
        RECT 712.200 353.700 714.000 360.600 ;
        RECT 722.400 354.600 724.200 357.600 ;
        RECT 722.400 353.700 723.600 354.600 ;
        RECT 728.400 353.700 730.200 357.600 ;
        RECT 741.150 353.700 742.950 357.600 ;
        RECT 750.450 353.700 752.250 357.600 ;
        RECT 757.350 353.700 759.150 357.600 ;
        RECT 766.350 353.700 768.150 357.600 ;
        RECT 781.800 353.700 783.600 357.600 ;
        RECT 787.800 353.700 789.600 357.600 ;
        RECT 802.800 353.700 804.600 357.600 ;
        RECT 812.400 353.700 814.200 358.800 ;
        RECT 831.450 353.700 840.450 429.300 ;
        RECT 0.600 351.300 840.450 353.700 ;
        RECT 13.500 344.400 15.300 351.300 ;
        RECT 28.800 347.400 30.600 351.300 ;
        RECT 41.700 347.400 43.500 351.300 ;
        RECT 49.200 344.400 51.000 351.300 ;
        RECT 56.700 341.400 58.500 351.300 ;
        RECT 74.700 344.400 76.500 351.300 ;
        RECT 92.400 350.400 93.600 351.300 ;
        RECT 92.400 347.400 94.200 350.400 ;
        RECT 98.400 347.400 100.200 351.300 ;
        RECT 124.500 341.400 126.300 351.300 ;
        RECT 142.500 344.400 144.300 351.300 ;
        RECT 152.400 346.200 154.200 351.300 ;
        RECT 175.500 344.400 177.300 351.300 ;
        RECT 196.800 345.900 198.600 351.300 ;
        RECT 207.150 347.400 208.950 351.300 ;
        RECT 216.450 347.400 218.250 351.300 ;
        RECT 223.350 347.400 225.150 351.300 ;
        RECT 232.350 347.400 234.150 351.300 ;
        RECT 242.400 347.400 244.200 351.300 ;
        RECT 259.800 347.400 261.600 351.300 ;
        RECT 265.800 347.400 267.600 351.300 ;
        RECT 280.800 347.400 282.600 351.300 ;
        RECT 287.850 347.400 289.650 351.300 ;
        RECT 296.850 347.400 298.650 351.300 ;
        RECT 303.750 347.400 305.550 351.300 ;
        RECT 313.050 347.400 314.850 351.300 ;
        RECT 334.800 346.200 336.600 351.300 ;
        RECT 352.500 344.400 354.300 351.300 ;
        RECT 362.700 344.400 364.500 351.300 ;
        RECT 377.850 347.400 379.650 351.300 ;
        RECT 386.850 347.400 388.650 351.300 ;
        RECT 393.750 347.400 395.550 351.300 ;
        RECT 403.050 347.400 404.850 351.300 ;
        RECT 414.150 347.400 415.950 351.300 ;
        RECT 423.450 347.400 425.250 351.300 ;
        RECT 430.350 347.400 432.150 351.300 ;
        RECT 439.350 347.400 441.150 351.300 ;
        RECT 452.700 347.400 454.500 351.300 ;
        RECT 460.200 344.400 462.000 351.300 ;
        RECT 470.400 347.400 472.200 351.300 ;
        RECT 476.400 347.400 478.200 351.300 ;
        RECT 490.800 347.400 492.600 351.300 ;
        RECT 496.800 347.400 498.600 351.300 ;
        RECT 514.500 344.400 516.300 351.300 ;
        RECT 532.800 346.200 534.600 351.300 ;
        RECT 547.800 347.400 549.600 351.300 ;
        RECT 555.150 347.400 556.950 351.300 ;
        RECT 564.450 347.400 566.250 351.300 ;
        RECT 571.350 347.400 573.150 351.300 ;
        RECT 580.350 347.400 582.150 351.300 ;
        RECT 593.400 347.400 595.200 351.300 ;
        RECT 599.400 347.400 601.200 351.300 ;
        RECT 619.500 344.400 621.300 351.300 ;
        RECT 637.500 344.400 639.300 351.300 ;
        RECT 650.700 344.400 652.500 351.300 ;
        RECT 670.800 346.200 672.600 351.300 ;
        RECT 681.150 347.400 682.950 351.300 ;
        RECT 690.450 347.400 692.250 351.300 ;
        RECT 697.350 347.400 699.150 351.300 ;
        RECT 706.350 347.400 708.150 351.300 ;
        RECT 716.400 347.400 718.200 351.300 ;
        RECT 736.800 344.400 738.600 351.300 ;
        RECT 745.200 344.400 747.000 351.300 ;
        RECT 753.150 347.400 754.950 351.300 ;
        RECT 762.450 347.400 764.250 351.300 ;
        RECT 769.350 347.400 771.150 351.300 ;
        RECT 778.350 347.400 780.150 351.300 ;
        RECT 788.400 347.400 790.200 351.300 ;
        RECT 794.400 347.400 796.200 351.300 ;
        RECT 806.400 347.400 808.200 351.300 ;
        RECT 812.400 347.400 814.200 351.300 ;
        RECT 6.150 275.700 7.950 279.600 ;
        RECT 15.450 275.700 17.250 279.600 ;
        RECT 22.350 275.700 24.150 279.600 ;
        RECT 31.350 275.700 33.150 279.600 ;
        RECT 41.700 275.700 43.500 282.600 ;
        RECT 56.850 275.700 58.650 279.600 ;
        RECT 65.850 275.700 67.650 279.600 ;
        RECT 72.750 275.700 74.550 279.600 ;
        RECT 82.050 275.700 83.850 279.600 ;
        RECT 98.400 275.700 100.200 280.800 ;
        RECT 121.800 275.700 123.600 280.800 ;
        RECT 136.800 275.700 138.600 279.600 ;
        RECT 143.850 275.700 145.650 279.600 ;
        RECT 152.850 275.700 154.650 279.600 ;
        RECT 159.750 275.700 161.550 279.600 ;
        RECT 169.050 275.700 170.850 279.600 ;
        RECT 180.150 275.700 181.950 279.600 ;
        RECT 189.450 275.700 191.250 279.600 ;
        RECT 196.350 275.700 198.150 279.600 ;
        RECT 205.350 275.700 207.150 279.600 ;
        RECT 216.150 275.700 217.950 279.600 ;
        RECT 225.450 275.700 227.250 279.600 ;
        RECT 232.350 275.700 234.150 279.600 ;
        RECT 241.350 275.700 243.150 279.600 ;
        RECT 251.400 275.700 253.200 279.600 ;
        RECT 268.800 275.700 270.600 279.600 ;
        RECT 274.800 275.700 276.600 279.600 ;
        RECT 283.800 275.700 285.600 279.600 ;
        RECT 289.800 275.700 291.600 279.600 ;
        RECT 301.800 275.700 303.600 279.600 ;
        RECT 307.800 275.700 309.600 279.600 ;
        RECT 322.800 275.700 324.600 279.600 ;
        RECT 329.850 275.700 331.650 279.600 ;
        RECT 338.850 275.700 340.650 279.600 ;
        RECT 345.750 275.700 347.550 279.600 ;
        RECT 355.050 275.700 356.850 279.600 ;
        RECT 371.400 275.700 373.200 280.800 ;
        RECT 392.400 275.700 394.200 280.800 ;
        RECT 418.800 275.700 420.600 280.800 ;
        RECT 428.700 275.700 430.500 282.600 ;
        RECT 446.400 275.700 448.200 280.800 ;
        RECT 461.850 275.700 463.650 279.600 ;
        RECT 470.850 275.700 472.650 279.600 ;
        RECT 477.750 275.700 479.550 279.600 ;
        RECT 487.050 275.700 488.850 279.600 ;
        RECT 497.700 275.700 499.500 282.600 ;
        RECT 517.800 275.700 519.600 279.600 ;
        RECT 523.800 275.700 525.600 279.600 ;
        RECT 531.000 275.700 532.800 282.600 ;
        RECT 538.500 275.700 540.300 279.600 ;
        RECT 551.700 275.700 553.500 282.600 ;
        RECT 571.800 275.700 573.600 280.800 ;
        RECT 584.700 275.700 586.500 282.600 ;
        RECT 599.400 275.700 601.200 279.600 ;
        RECT 605.400 275.700 607.200 279.600 ;
        RECT 617.400 275.700 619.200 279.600 ;
        RECT 623.400 275.700 625.200 279.600 ;
        RECT 633.000 275.700 634.800 282.600 ;
        RECT 640.500 275.700 642.300 279.600 ;
        RECT 661.800 275.700 663.600 280.800 ;
        RECT 678.300 275.700 680.100 282.600 ;
        RECT 694.800 275.700 696.600 279.600 ;
        RECT 700.800 275.700 702.600 279.600 ;
        RECT 707.400 275.700 709.200 279.600 ;
        RECT 713.400 275.700 715.200 279.600 ;
        RECT 725.400 275.700 727.200 280.800 ;
        RECT 751.800 275.700 753.600 280.800 ;
        RECT 764.400 275.700 766.200 279.600 ;
        RECT 770.400 275.700 772.200 279.600 ;
        RECT 782.400 275.700 784.200 279.600 ;
        RECT 802.500 275.700 804.300 282.600 ;
        RECT 815.400 275.700 817.200 280.800 ;
        RECT 831.450 275.700 840.450 351.300 ;
        RECT 0.600 273.300 840.450 275.700 ;
        RECT 6.150 269.400 7.950 273.300 ;
        RECT 15.450 269.400 17.250 273.300 ;
        RECT 22.350 269.400 24.150 273.300 ;
        RECT 31.350 269.400 33.150 273.300 ;
        RECT 52.800 268.200 54.600 273.300 ;
        RECT 65.400 269.400 67.200 273.300 ;
        RECT 80.400 269.400 82.200 273.300 ;
        RECT 93.150 269.400 94.950 273.300 ;
        RECT 102.450 269.400 104.250 273.300 ;
        RECT 109.350 269.400 111.150 273.300 ;
        RECT 118.350 269.400 120.150 273.300 ;
        RECT 131.400 269.400 133.200 273.300 ;
        RECT 144.150 269.400 145.950 273.300 ;
        RECT 153.450 269.400 155.250 273.300 ;
        RECT 160.350 269.400 162.150 273.300 ;
        RECT 169.350 269.400 171.150 273.300 ;
        RECT 182.400 268.200 184.200 273.300 ;
        RECT 205.800 269.400 207.600 273.300 ;
        RECT 215.400 269.400 217.200 273.300 ;
        RECT 221.400 269.400 223.200 273.300 ;
        RECT 238.800 269.400 240.600 273.300 ;
        RECT 248.400 269.400 250.200 273.300 ;
        RECT 254.400 269.400 256.200 273.300 ;
        RECT 263.400 269.400 265.200 273.300 ;
        RECT 269.400 269.400 271.200 273.300 ;
        RECT 281.400 269.400 283.200 273.300 ;
        RECT 293.400 269.400 295.200 273.300 ;
        RECT 299.400 269.400 301.200 273.300 ;
        RECT 314.400 268.200 316.200 273.300 ;
        RECT 329.400 269.400 331.200 273.300 ;
        RECT 344.700 266.400 346.500 273.300 ;
        RECT 359.850 269.400 361.650 273.300 ;
        RECT 368.850 269.400 370.650 273.300 ;
        RECT 375.750 269.400 377.550 273.300 ;
        RECT 385.050 269.400 386.850 273.300 ;
        RECT 406.800 268.200 408.600 273.300 ;
        RECT 424.800 268.200 426.600 273.300 ;
        RECT 437.400 269.400 439.200 273.300 ;
        RECT 460.800 268.200 462.600 273.300 ;
        RECT 470.400 269.400 472.200 273.300 ;
        RECT 476.400 269.400 478.200 273.300 ;
        RECT 496.800 268.200 498.600 273.300 ;
        RECT 514.800 269.400 516.600 273.300 ;
        RECT 521.850 269.400 523.650 273.300 ;
        RECT 530.850 269.400 532.650 273.300 ;
        RECT 537.750 269.400 539.550 273.300 ;
        RECT 547.050 269.400 548.850 273.300 ;
        RECT 557.400 269.400 559.200 273.300 ;
        RECT 563.400 269.400 565.200 273.300 ;
        RECT 576.000 266.400 577.800 273.300 ;
        RECT 583.500 269.400 585.300 273.300 ;
        RECT 601.800 269.400 603.600 273.300 ;
        RECT 616.800 268.200 618.600 273.300 ;
        RECT 626.400 269.400 628.200 273.300 ;
        RECT 641.400 269.400 643.200 273.300 ;
        RECT 653.400 269.400 655.200 273.300 ;
        RECT 659.400 269.400 661.200 273.300 ;
        RECT 672.900 266.400 674.700 273.300 ;
        RECT 686.700 266.400 688.500 273.300 ;
        RECT 705.000 266.400 706.800 273.300 ;
        RECT 712.500 269.400 714.300 273.300 ;
        RECT 725.700 266.400 727.500 273.300 ;
        RECT 743.700 266.400 745.500 273.300 ;
        RECT 763.800 269.400 765.600 273.300 ;
        RECT 769.800 269.400 771.600 273.300 ;
        RECT 782.700 269.400 784.500 273.300 ;
        RECT 790.200 266.400 792.000 273.300 ;
        RECT 797.850 269.400 799.650 273.300 ;
        RECT 806.850 269.400 808.650 273.300 ;
        RECT 813.750 269.400 815.550 273.300 ;
        RECT 823.050 269.400 824.850 273.300 ;
        RECT 19.800 197.700 21.600 203.100 ;
        RECT 34.800 197.700 36.600 201.600 ;
        RECT 40.800 197.700 42.600 201.600 ;
        RECT 58.500 197.700 60.300 204.600 ;
        RECT 67.800 197.700 69.600 201.600 ;
        RECT 73.800 197.700 75.600 201.600 ;
        RECT 82.800 197.700 84.600 201.600 ;
        RECT 88.800 197.700 90.600 201.600 ;
        RECT 101.700 197.700 103.500 201.600 ;
        RECT 109.200 197.700 111.000 204.600 ;
        RECT 124.500 197.700 126.300 204.600 ;
        RECT 136.800 197.700 138.600 201.600 ;
        RECT 142.800 197.700 144.600 201.600 ;
        RECT 149.400 197.700 151.200 201.600 ;
        RECT 155.400 197.700 157.200 201.600 ;
        RECT 167.400 197.700 169.200 201.600 ;
        RECT 173.400 197.700 175.200 201.600 ;
        RECT 185.400 197.700 187.200 202.800 ;
        RECT 211.500 197.700 213.300 204.600 ;
        RECT 221.700 197.700 223.500 201.600 ;
        RECT 229.200 197.700 231.000 204.600 ;
        RECT 240.900 197.700 242.700 204.600 ;
        RECT 257.700 197.700 259.500 207.600 ;
        RECT 279.000 197.700 280.800 204.600 ;
        RECT 286.500 197.700 288.300 201.600 ;
        RECT 300.900 197.700 302.700 204.600 ;
        RECT 315.150 197.700 316.950 201.600 ;
        RECT 324.450 197.700 326.250 201.600 ;
        RECT 331.350 197.700 333.150 201.600 ;
        RECT 340.350 197.700 342.150 201.600 ;
        RECT 361.500 197.700 363.300 204.600 ;
        RECT 371.400 197.700 373.200 202.800 ;
        RECT 397.800 197.700 399.600 202.800 ;
        RECT 415.800 197.700 417.600 204.600 ;
        RECT 425.700 197.700 427.500 204.600 ;
        RECT 438.150 197.700 439.950 201.600 ;
        RECT 447.450 197.700 449.250 201.600 ;
        RECT 454.350 197.700 456.150 201.600 ;
        RECT 463.350 197.700 465.150 201.600 ;
        RECT 481.800 197.700 483.600 201.600 ;
        RECT 488.700 197.700 490.500 204.600 ;
        RECT 506.400 197.700 508.200 201.600 ;
        RECT 512.400 197.700 514.200 201.600 ;
        RECT 529.800 197.700 531.600 202.800 ;
        RECT 547.800 197.700 549.600 201.600 ;
        RECT 557.400 197.700 559.200 201.600 ;
        RECT 563.400 197.700 565.200 201.600 ;
        RECT 575.400 197.700 577.200 201.600 ;
        RECT 590.400 197.700 592.200 204.600 ;
        RECT 596.400 197.700 598.200 204.600 ;
        RECT 602.400 197.700 604.200 204.600 ;
        RECT 608.400 197.700 610.200 204.600 ;
        RECT 614.400 197.700 616.200 204.600 ;
        RECT 624.150 197.700 625.950 201.600 ;
        RECT 633.450 197.700 635.250 201.600 ;
        RECT 640.350 197.700 642.150 201.600 ;
        RECT 649.350 197.700 651.150 201.600 ;
        RECT 662.400 197.700 664.200 202.800 ;
        RECT 682.800 197.700 684.600 201.600 ;
        RECT 688.800 197.700 690.600 201.600 ;
        RECT 697.800 197.700 699.600 201.600 ;
        RECT 703.800 197.700 705.600 201.600 ;
        RECT 710.400 198.600 712.200 201.600 ;
        RECT 710.400 197.700 711.600 198.600 ;
        RECT 716.400 197.700 718.200 201.600 ;
        RECT 736.500 197.700 738.300 204.600 ;
        RECT 743.850 197.700 745.650 201.600 ;
        RECT 752.850 197.700 754.650 201.600 ;
        RECT 759.750 197.700 761.550 201.600 ;
        RECT 769.050 197.700 770.850 201.600 ;
        RECT 779.700 197.700 781.500 204.600 ;
        RECT 797.400 197.700 799.200 201.600 ;
        RECT 812.400 197.700 814.200 201.600 ;
        RECT 831.450 197.700 840.450 273.300 ;
        RECT 0.600 195.300 840.450 197.700 ;
        RECT 10.800 191.400 12.600 195.300 ;
        RECT 17.850 191.400 19.650 195.300 ;
        RECT 26.850 191.400 28.650 195.300 ;
        RECT 33.750 191.400 35.550 195.300 ;
        RECT 43.050 191.400 44.850 195.300 ;
        RECT 59.400 190.200 61.200 195.300 ;
        RECT 77.700 188.400 79.500 195.300 ;
        RECT 98.400 190.200 100.200 195.300 ;
        RECT 113.850 191.400 115.650 195.300 ;
        RECT 122.850 191.400 124.650 195.300 ;
        RECT 129.750 191.400 131.550 195.300 ;
        RECT 139.050 191.400 140.850 195.300 ;
        RECT 154.500 188.400 156.300 195.300 ;
        RECT 169.800 191.400 171.600 195.300 ;
        RECT 176.850 191.400 178.650 195.300 ;
        RECT 185.850 191.400 187.650 195.300 ;
        RECT 192.750 191.400 194.550 195.300 ;
        RECT 202.050 191.400 203.850 195.300 ;
        RECT 215.400 190.200 217.200 195.300 ;
        RECT 235.800 188.400 237.600 195.300 ;
        RECT 241.800 188.400 243.600 195.300 ;
        RECT 247.800 188.400 249.600 195.300 ;
        RECT 253.800 188.400 255.600 195.300 ;
        RECT 259.800 188.400 261.600 195.300 ;
        RECT 272.400 190.200 274.200 195.300 ;
        RECT 297.300 188.400 299.100 195.300 ;
        RECT 311.400 191.400 313.200 195.300 ;
        RECT 317.400 191.400 319.200 195.300 ;
        RECT 329.400 190.200 331.200 195.300 ;
        RECT 347.400 191.400 349.200 195.300 ;
        RECT 359.850 191.400 361.650 195.300 ;
        RECT 368.850 191.400 370.650 195.300 ;
        RECT 375.750 191.400 377.550 195.300 ;
        RECT 385.050 191.400 386.850 195.300 ;
        RECT 397.800 191.400 399.600 195.300 ;
        RECT 403.800 191.400 405.600 195.300 ;
        RECT 416.700 191.400 418.500 195.300 ;
        RECT 424.200 188.400 426.000 195.300 ;
        RECT 433.800 188.400 435.600 195.300 ;
        RECT 439.800 188.400 441.600 195.300 ;
        RECT 445.800 188.400 447.600 195.300 ;
        RECT 451.800 188.400 453.600 195.300 ;
        RECT 457.800 188.400 459.600 195.300 ;
        RECT 467.400 188.400 469.200 195.300 ;
        RECT 473.400 188.400 475.200 195.300 ;
        RECT 479.400 188.400 481.200 195.300 ;
        RECT 485.400 188.400 487.200 195.300 ;
        RECT 491.400 188.400 493.200 195.300 ;
        RECT 511.500 188.400 513.300 195.300 ;
        RECT 529.800 190.200 531.600 195.300 ;
        RECT 539.850 191.400 541.650 195.300 ;
        RECT 548.850 191.400 550.650 195.300 ;
        RECT 555.750 191.400 557.550 195.300 ;
        RECT 565.050 191.400 566.850 195.300 ;
        RECT 586.800 190.200 588.600 195.300 ;
        RECT 606.300 188.400 608.100 195.300 ;
        RECT 620.400 190.200 622.200 195.300 ;
        RECT 638.700 188.400 640.500 195.300 ;
        RECT 650.400 191.400 652.200 195.300 ;
        RECT 665.400 191.400 667.200 195.300 ;
        RECT 685.800 190.200 687.600 195.300 ;
        RECT 698.400 191.400 700.200 195.300 ;
        RECT 704.400 191.400 706.200 195.300 ;
        RECT 716.400 191.400 718.200 195.300 ;
        RECT 722.400 191.400 724.200 195.300 ;
        RECT 734.400 191.400 736.200 195.300 ;
        RECT 751.800 191.400 753.600 195.300 ;
        RECT 764.400 190.200 766.200 195.300 ;
        RECT 787.500 188.400 789.300 195.300 ;
        RECT 795.150 191.400 796.950 195.300 ;
        RECT 804.450 191.400 806.250 195.300 ;
        RECT 811.350 191.400 813.150 195.300 ;
        RECT 820.350 191.400 822.150 195.300 ;
        RECT 6.150 119.700 7.950 123.600 ;
        RECT 15.450 119.700 17.250 123.600 ;
        RECT 22.350 119.700 24.150 123.600 ;
        RECT 31.350 119.700 33.150 123.600 ;
        RECT 43.800 119.700 45.600 123.600 ;
        RECT 49.800 119.700 51.600 123.600 ;
        RECT 56.400 119.700 58.200 123.600 ;
        RECT 71.400 119.700 73.200 124.800 ;
        RECT 91.800 119.700 93.600 123.600 ;
        RECT 97.800 119.700 99.600 123.600 ;
        RECT 110.400 119.700 112.200 124.800 ;
        RECT 133.500 119.700 135.300 126.600 ;
        RECT 142.800 119.700 144.600 123.600 ;
        RECT 148.800 119.700 150.600 123.600 ;
        RECT 163.500 119.700 165.300 126.600 ;
        RECT 178.800 119.700 180.600 123.600 ;
        RECT 191.400 119.700 193.200 124.800 ;
        RECT 217.800 119.700 219.600 124.800 ;
        RECT 235.800 119.700 237.600 123.600 ;
        RECT 242.700 119.700 244.500 126.600 ;
        RECT 257.700 119.700 259.500 126.600 ;
        RECT 275.700 119.700 277.500 126.600 ;
        RECT 293.400 120.600 295.200 123.600 ;
        RECT 293.400 119.700 294.600 120.600 ;
        RECT 299.400 119.700 301.200 123.600 ;
        RECT 317.700 119.700 319.500 123.600 ;
        RECT 325.200 119.700 327.000 126.600 ;
        RECT 332.700 119.700 334.500 126.600 ;
        RECT 350.700 119.700 352.500 126.600 ;
        RECT 371.400 119.700 373.200 124.800 ;
        RECT 394.500 119.700 396.300 126.600 ;
        RECT 402.150 119.700 403.950 123.600 ;
        RECT 411.450 119.700 413.250 123.600 ;
        RECT 418.350 119.700 420.150 123.600 ;
        RECT 427.350 119.700 429.150 123.600 ;
        RECT 441.000 119.700 442.800 126.600 ;
        RECT 449.400 119.700 451.200 126.600 ;
        RECT 467.700 119.700 469.500 126.600 ;
        RECT 487.800 119.700 489.600 124.800 ;
        RECT 497.850 119.700 499.650 123.600 ;
        RECT 506.850 119.700 508.650 123.600 ;
        RECT 513.750 119.700 515.550 123.600 ;
        RECT 523.050 119.700 524.850 123.600 ;
        RECT 533.400 119.700 535.200 123.600 ;
        RECT 539.400 119.700 541.200 123.600 ;
        RECT 548.850 119.700 550.650 123.600 ;
        RECT 557.850 119.700 559.650 123.600 ;
        RECT 564.750 119.700 566.550 123.600 ;
        RECT 574.050 119.700 575.850 123.600 ;
        RECT 587.700 119.700 589.500 123.600 ;
        RECT 595.200 119.700 597.000 126.600 ;
        RECT 610.800 119.700 612.600 123.600 ;
        RECT 616.800 120.600 618.600 123.600 ;
        RECT 617.400 119.700 618.600 120.600 ;
        RECT 626.400 119.700 628.200 123.600 ;
        RECT 641.700 119.700 643.500 126.600 ;
        RECT 656.850 119.700 658.650 123.600 ;
        RECT 665.850 119.700 667.650 123.600 ;
        RECT 672.750 119.700 674.550 123.600 ;
        RECT 682.050 119.700 683.850 123.600 ;
        RECT 692.700 119.700 694.500 126.600 ;
        RECT 718.800 119.700 720.600 124.800 ;
        RECT 736.800 119.700 738.600 124.800 ;
        RECT 750.000 119.700 751.800 126.600 ;
        RECT 757.500 119.700 759.300 123.600 ;
        RECT 775.800 119.700 777.600 124.800 ;
        RECT 785.400 119.700 787.200 123.600 ;
        RECT 791.400 119.700 793.200 123.600 ;
        RECT 803.400 119.700 805.200 123.600 ;
        RECT 815.700 119.700 817.500 126.600 ;
        RECT 831.450 119.700 840.450 195.300 ;
        RECT 0.600 117.300 840.450 119.700 ;
        RECT 10.800 113.400 12.600 117.300 ;
        RECT 16.800 113.400 18.600 117.300 ;
        RECT 26.400 113.400 28.200 117.300 ;
        RECT 32.400 113.400 34.200 117.300 ;
        RECT 44.700 113.400 46.500 117.300 ;
        RECT 52.200 110.400 54.000 117.300 ;
        RECT 62.400 116.400 63.600 117.300 ;
        RECT 62.400 113.400 64.200 116.400 ;
        RECT 68.400 113.400 70.200 117.300 ;
        RECT 80.700 110.400 82.500 117.300 ;
        RECT 95.700 110.400 97.500 117.300 ;
        RECT 110.700 110.400 112.500 117.300 ;
        RECT 136.800 112.200 138.600 117.300 ;
        RECT 149.400 113.400 151.200 117.300 ;
        RECT 172.500 110.400 174.300 117.300 ;
        RECT 179.850 113.400 181.650 117.300 ;
        RECT 188.850 113.400 190.650 117.300 ;
        RECT 195.750 113.400 197.550 117.300 ;
        RECT 205.050 113.400 206.850 117.300 ;
        RECT 219.900 110.400 221.700 117.300 ;
        RECT 236.400 112.200 238.200 117.300 ;
        RECT 251.700 110.400 253.500 117.300 ;
        RECT 271.500 110.400 273.300 117.300 ;
        RECT 291.300 110.400 293.100 117.300 ;
        RECT 302.400 113.400 304.200 117.300 ;
        RECT 308.400 113.400 310.200 117.300 ;
        RECT 323.400 112.200 325.200 117.300 ;
        RECT 346.500 110.400 348.300 117.300 ;
        RECT 362.400 112.200 364.200 117.300 ;
        RECT 378.150 113.400 379.950 117.300 ;
        RECT 387.450 113.400 389.250 117.300 ;
        RECT 394.350 113.400 396.150 117.300 ;
        RECT 403.350 113.400 405.150 117.300 ;
        RECT 413.700 110.400 415.500 117.300 ;
        RECT 429.150 113.400 430.950 117.300 ;
        RECT 438.450 113.400 440.250 117.300 ;
        RECT 445.350 113.400 447.150 117.300 ;
        RECT 454.350 113.400 456.150 117.300 ;
        RECT 469.800 113.400 471.600 117.300 ;
        RECT 475.800 113.400 477.600 117.300 ;
        RECT 490.800 112.200 492.600 117.300 ;
        RECT 500.700 107.400 502.500 117.300 ;
        RECT 518.850 113.400 520.650 117.300 ;
        RECT 527.850 113.400 529.650 117.300 ;
        RECT 534.750 113.400 536.550 117.300 ;
        RECT 544.050 113.400 545.850 117.300 ;
        RECT 557.700 110.400 559.500 117.300 ;
        RECT 576.000 110.400 577.800 117.300 ;
        RECT 584.400 110.400 586.200 117.300 ;
        RECT 599.400 112.200 601.200 117.300 ;
        RECT 617.700 110.400 619.500 117.300 ;
        RECT 638.400 112.200 640.200 117.300 ;
        RECT 656.700 110.400 658.500 117.300 ;
        RECT 668.850 113.400 670.650 117.300 ;
        RECT 677.850 113.400 679.650 117.300 ;
        RECT 684.750 113.400 686.550 117.300 ;
        RECT 694.050 113.400 695.850 117.300 ;
        RECT 705.000 110.400 706.800 117.300 ;
        RECT 713.400 110.400 715.200 117.300 ;
        RECT 731.700 113.400 733.500 117.300 ;
        RECT 739.200 110.400 741.000 117.300 ;
        RECT 746.400 116.400 747.600 117.300 ;
        RECT 746.400 113.400 748.200 116.400 ;
        RECT 752.400 113.400 754.200 117.300 ;
        RECT 764.850 113.400 766.650 117.300 ;
        RECT 773.850 113.400 775.650 117.300 ;
        RECT 780.750 113.400 782.550 117.300 ;
        RECT 790.050 113.400 791.850 117.300 ;
        RECT 806.400 112.200 808.200 117.300 ;
        RECT 6.150 41.700 7.950 45.600 ;
        RECT 15.450 41.700 17.250 45.600 ;
        RECT 22.350 41.700 24.150 45.600 ;
        RECT 31.350 41.700 33.150 45.600 ;
        RECT 41.850 41.700 43.650 45.600 ;
        RECT 50.850 41.700 52.650 45.600 ;
        RECT 57.750 41.700 59.550 45.600 ;
        RECT 67.050 41.700 68.850 45.600 ;
        RECT 83.400 41.700 85.200 46.800 ;
        RECT 99.150 41.700 100.950 45.600 ;
        RECT 108.450 41.700 110.250 45.600 ;
        RECT 115.350 41.700 117.150 45.600 ;
        RECT 124.350 41.700 126.150 45.600 ;
        RECT 137.700 41.700 139.500 48.600 ;
        RECT 155.400 41.700 157.200 46.800 ;
        RECT 171.150 41.700 172.950 45.600 ;
        RECT 180.450 41.700 182.250 45.600 ;
        RECT 187.350 41.700 189.150 45.600 ;
        RECT 196.350 41.700 198.150 45.600 ;
        RECT 209.700 41.700 211.500 48.600 ;
        RECT 225.150 41.700 226.950 45.600 ;
        RECT 234.450 41.700 236.250 45.600 ;
        RECT 241.350 41.700 243.150 45.600 ;
        RECT 250.350 41.700 252.150 45.600 ;
        RECT 260.700 41.700 262.500 48.600 ;
        RECT 283.800 41.700 285.600 46.800 ;
        RECT 296.700 41.700 298.500 48.600 ;
        RECT 312.000 41.700 313.800 48.600 ;
        RECT 320.400 41.700 322.200 48.600 ;
        RECT 343.800 41.700 345.600 46.800 ;
        RECT 358.800 41.700 360.600 45.600 ;
        RECT 366.150 41.700 367.950 45.600 ;
        RECT 375.450 41.700 377.250 45.600 ;
        RECT 382.350 41.700 384.150 45.600 ;
        RECT 391.350 41.700 393.150 45.600 ;
        RECT 406.800 41.700 408.600 48.600 ;
        RECT 415.200 41.700 417.000 48.600 ;
        RECT 430.500 41.700 432.300 48.600 ;
        RECT 443.400 41.700 445.200 45.600 ;
        RECT 449.400 41.700 451.200 45.600 ;
        RECT 461.400 41.700 463.200 45.600 ;
        RECT 479.400 41.700 481.200 46.800 ;
        RECT 505.800 41.700 507.600 46.800 ;
        RECT 523.800 41.700 525.600 45.600 ;
        RECT 531.150 41.700 532.950 45.600 ;
        RECT 540.450 41.700 542.250 45.600 ;
        RECT 547.350 41.700 549.150 45.600 ;
        RECT 556.350 41.700 558.150 45.600 ;
        RECT 569.400 41.700 571.200 45.600 ;
        RECT 582.150 41.700 583.950 45.600 ;
        RECT 591.450 41.700 593.250 45.600 ;
        RECT 598.350 41.700 600.150 45.600 ;
        RECT 607.350 41.700 609.150 45.600 ;
        RECT 628.800 41.700 630.600 46.800 ;
        RECT 640.800 41.700 642.600 48.600 ;
        RECT 646.800 41.700 648.600 48.600 ;
        RECT 652.800 41.700 654.600 48.600 ;
        RECT 665.700 41.700 667.500 48.600 ;
        RECT 688.500 41.700 690.300 48.600 ;
        RECT 698.400 41.700 700.200 45.600 ;
        RECT 721.800 41.700 723.600 46.800 ;
        RECT 731.700 41.700 733.500 48.600 ;
        RECT 752.400 41.700 754.200 46.800 ;
        RECT 778.800 41.700 780.600 46.800 ;
        RECT 788.400 41.700 790.200 45.600 ;
        RECT 803.400 41.700 805.200 45.600 ;
        RECT 818.700 41.700 820.500 48.600 ;
        RECT 831.450 41.700 840.450 117.300 ;
        RECT 0.600 39.300 840.450 41.700 ;
        RECT 10.800 35.400 12.600 39.300 ;
        RECT 22.800 35.400 24.600 39.300 ;
        RECT 28.800 35.400 30.600 39.300 ;
        RECT 43.800 35.400 45.600 39.300 ;
        RECT 52.800 35.400 54.600 39.300 ;
        RECT 58.800 35.400 60.600 39.300 ;
        RECT 71.400 34.200 73.200 39.300 ;
        RECT 89.400 35.400 91.200 39.300 ;
        RECT 109.800 35.400 111.600 39.300 ;
        RECT 119.400 34.200 121.200 39.300 ;
        RECT 134.400 35.400 136.200 39.300 ;
        RECT 146.700 29.400 148.500 39.300 ;
        RECT 175.500 32.400 177.300 39.300 ;
        RECT 182.700 32.400 184.500 39.300 ;
        RECT 203.400 34.200 205.200 39.300 ;
        RECT 219.150 35.400 220.950 39.300 ;
        RECT 228.450 35.400 230.250 39.300 ;
        RECT 235.350 35.400 237.150 39.300 ;
        RECT 244.350 35.400 246.150 39.300 ;
        RECT 255.150 35.400 256.950 39.300 ;
        RECT 264.450 35.400 266.250 39.300 ;
        RECT 271.350 35.400 273.150 39.300 ;
        RECT 280.350 35.400 282.150 39.300 ;
        RECT 295.800 32.400 297.600 39.300 ;
        RECT 304.200 32.400 306.000 39.300 ;
        RECT 316.800 35.400 318.600 39.300 ;
        RECT 322.800 35.400 324.600 39.300 ;
        RECT 329.850 35.400 331.650 39.300 ;
        RECT 338.850 35.400 340.650 39.300 ;
        RECT 345.750 35.400 347.550 39.300 ;
        RECT 355.050 35.400 356.850 39.300 ;
        RECT 368.700 35.400 370.500 39.300 ;
        RECT 376.200 32.400 378.000 39.300 ;
        RECT 384.150 35.400 385.950 39.300 ;
        RECT 393.450 35.400 395.250 39.300 ;
        RECT 400.350 35.400 402.150 39.300 ;
        RECT 409.350 35.400 411.150 39.300 ;
        RECT 427.500 32.400 429.300 39.300 ;
        RECT 448.800 34.200 450.600 39.300 ;
        RECT 463.500 32.400 465.300 39.300 ;
        RECT 484.800 34.200 486.600 39.300 ;
        RECT 500.700 32.400 502.500 39.300 ;
        RECT 515.700 32.400 517.500 39.300 ;
        RECT 532.800 35.400 534.600 39.300 ;
        RECT 539.400 35.400 541.200 39.300 ;
        RECT 545.400 35.400 547.200 39.300 ;
        RECT 565.800 34.200 567.600 39.300 ;
        RECT 575.700 32.400 577.500 39.300 ;
        RECT 590.850 35.400 592.650 39.300 ;
        RECT 599.850 35.400 601.650 39.300 ;
        RECT 606.750 35.400 608.550 39.300 ;
        RECT 616.050 35.400 617.850 39.300 ;
        RECT 629.700 32.400 631.500 39.300 ;
        RECT 655.500 32.400 657.300 39.300 ;
        RECT 662.850 35.400 664.650 39.300 ;
        RECT 671.850 35.400 673.650 39.300 ;
        RECT 678.750 35.400 680.550 39.300 ;
        RECT 688.050 35.400 689.850 39.300 ;
        RECT 706.800 34.200 708.600 39.300 ;
        RECT 721.800 35.400 723.600 39.300 ;
        RECT 727.800 35.400 729.600 39.300 ;
        RECT 745.500 29.400 747.300 39.300 ;
        RECT 752.850 35.400 754.650 39.300 ;
        RECT 761.850 35.400 763.650 39.300 ;
        RECT 768.750 35.400 770.550 39.300 ;
        RECT 778.050 35.400 779.850 39.300 ;
        RECT 791.700 32.400 793.500 39.300 ;
        RECT 806.700 32.400 808.500 39.300 ;
        RECT 831.450 0.300 840.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 782.700 -0.450 821.700 ;
        RECT 13.800 782.700 15.600 793.800 ;
        RECT 28.800 782.700 30.600 789.000 ;
        RECT 34.800 782.700 36.600 789.600 ;
        RECT 49.800 782.700 51.600 789.600 ;
        RECT 59.400 782.700 61.200 793.800 ;
        RECT 79.800 782.700 81.600 789.600 ;
        RECT 85.800 782.700 87.600 789.600 ;
        RECT 103.800 782.700 105.600 795.600 ;
        RECT 110.400 782.700 112.200 789.600 ;
        RECT 116.400 782.700 118.200 789.600 ;
        RECT 128.400 782.700 130.200 789.600 ;
        RECT 135.900 782.700 137.700 795.600 ;
        RECT 148.800 782.700 150.600 789.600 ;
        RECT 154.800 782.700 156.600 789.600 ;
        RECT 169.500 782.700 171.300 795.600 ;
        RECT 187.200 782.700 189.000 795.600 ;
        RECT 193.800 782.700 195.600 789.600 ;
        RECT 208.800 782.700 210.600 789.000 ;
        RECT 214.800 782.700 216.600 789.600 ;
        RECT 227.400 782.700 229.200 793.800 ;
        RECT 245.400 782.700 247.200 789.600 ;
        RECT 251.400 782.700 253.200 789.000 ;
        RECT 267.300 782.700 269.100 795.600 ;
        RECT 274.800 782.700 276.600 789.600 ;
        RECT 287.400 782.700 289.200 789.600 ;
        RECT 305.400 782.700 307.200 789.600 ;
        RECT 312.900 782.700 314.700 795.600 ;
        RECT 323.400 782.700 325.200 789.600 ;
        RECT 330.900 782.700 332.700 795.600 ;
        RECT 349.800 782.700 351.600 793.800 ;
        RECT 359.400 782.700 361.200 789.600 ;
        RECT 365.400 782.700 367.200 789.000 ;
        RECT 385.800 782.700 387.600 789.000 ;
        RECT 391.800 782.700 393.600 789.600 ;
        RECT 409.800 782.700 411.600 793.800 ;
        RECT 427.800 782.700 429.600 789.000 ;
        RECT 433.800 782.700 435.600 789.600 ;
        RECT 448.800 782.700 450.600 793.800 ;
        RECT 464.400 782.700 466.200 793.800 ;
        RECT 479.400 782.700 481.200 789.600 ;
        RECT 494.400 782.700 496.200 789.600 ;
        RECT 501.900 782.700 503.700 795.600 ;
        RECT 513.300 782.700 515.100 795.600 ;
        RECT 520.800 782.700 522.600 789.600 ;
        RECT 533.400 782.700 535.200 789.600 ;
        RECT 539.400 782.700 541.200 789.000 ;
        RECT 554.400 782.700 556.200 793.800 ;
        RECT 573.300 782.700 575.100 795.600 ;
        RECT 580.800 782.700 582.600 789.600 ;
        RECT 598.800 782.700 600.600 789.000 ;
        RECT 604.800 782.700 606.600 789.600 ;
        RECT 617.400 782.700 619.200 793.800 ;
        RECT 635.400 782.700 637.200 789.600 ;
        RECT 641.400 782.700 643.200 789.600 ;
        RECT 658.500 782.700 660.300 795.600 ;
        RECT 673.800 782.700 675.600 789.600 ;
        RECT 679.800 782.700 681.600 789.600 ;
        RECT 689.400 782.700 691.200 793.800 ;
        RECT 715.800 782.700 717.600 795.600 ;
        RECT 722.400 782.700 724.200 789.600 ;
        RECT 728.400 782.700 730.200 789.600 ;
        RECT 738.300 782.700 740.100 795.600 ;
        RECT 745.800 782.700 747.600 789.600 ;
        RECT 759.300 782.700 761.100 795.600 ;
        RECT 766.800 782.700 768.600 789.600 ;
        RECT 779.400 782.700 781.200 789.600 ;
        RECT 785.400 782.700 787.200 789.000 ;
        RECT 802.800 782.700 804.600 789.000 ;
        RECT 808.800 782.700 810.600 789.600 ;
        RECT 818.400 782.700 820.200 793.800 ;
        RECT -9.450 780.300 830.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT 8.400 773.400 10.200 780.300 ;
        RECT 15.900 767.400 17.700 780.300 ;
        RECT 23.400 773.400 25.200 780.300 ;
        RECT 36.300 767.400 38.100 780.300 ;
        RECT 43.800 773.400 45.600 780.300 ;
        RECT 64.800 769.200 66.600 780.300 ;
        RECT 74.400 773.400 76.200 780.300 ;
        RECT 80.400 774.000 82.200 780.300 ;
        RECT 95.400 773.400 97.200 780.300 ;
        RECT 101.400 774.000 103.200 780.300 ;
        RECT 113.400 773.400 115.200 780.300 ;
        RECT 119.400 773.400 121.200 780.300 ;
        RECT 128.400 773.400 130.200 780.300 ;
        RECT 134.400 773.400 136.200 780.300 ;
        RECT 149.400 769.500 151.200 780.300 ;
        RECT 178.800 769.200 180.600 780.300 ;
        RECT 188.400 773.400 190.200 780.300 ;
        RECT 194.400 774.000 196.200 780.300 ;
        RECT 212.400 773.400 214.200 780.300 ;
        RECT 219.900 767.400 221.700 780.300 ;
        RECT 230.400 773.400 232.200 780.300 ;
        RECT 237.900 767.400 239.700 780.300 ;
        RECT 253.800 774.000 255.600 780.300 ;
        RECT 259.800 773.400 261.600 780.300 ;
        RECT 277.800 769.200 279.600 780.300 ;
        RECT 293.400 769.200 295.200 780.300 ;
        RECT 313.800 774.000 315.600 780.300 ;
        RECT 319.800 773.400 321.600 780.300 ;
        RECT 331.800 774.000 333.600 780.300 ;
        RECT 337.800 773.400 339.600 780.300 ;
        RECT 352.800 774.000 354.600 780.300 ;
        RECT 358.800 773.400 360.600 780.300 ;
        RECT 370.800 773.400 372.600 780.300 ;
        RECT 388.800 769.200 390.600 780.300 ;
        RECT 403.800 774.000 405.600 780.300 ;
        RECT 409.800 773.400 411.600 780.300 ;
        RECT 416.400 773.400 418.200 780.300 ;
        RECT 442.800 769.500 444.600 780.300 ;
        RECT 452.400 773.400 454.200 780.300 ;
        RECT 458.400 773.400 460.200 780.300 ;
        RECT 468.300 767.400 470.100 780.300 ;
        RECT 475.800 773.400 477.600 780.300 ;
        RECT 490.800 774.000 492.600 780.300 ;
        RECT 496.800 773.400 498.600 780.300 ;
        RECT 511.800 769.200 513.600 780.300 ;
        RECT 524.400 773.400 526.200 780.300 ;
        RECT 530.400 774.000 532.200 780.300 ;
        RECT 547.800 773.400 549.600 780.300 ;
        RECT 553.800 773.400 555.600 780.300 ;
        RECT 563.400 773.400 565.200 780.300 ;
        RECT 570.900 767.400 572.700 780.300 ;
        RECT 578.400 773.400 580.200 780.300 ;
        RECT 593.400 769.500 595.200 780.300 ;
        RECT 616.800 773.400 618.600 780.300 ;
        RECT 628.800 773.400 630.600 780.300 ;
        RECT 634.800 773.400 636.600 780.300 ;
        RECT 643.800 773.400 645.600 780.300 ;
        RECT 649.800 773.400 651.600 780.300 ;
        RECT 659.400 767.400 661.200 780.300 ;
        RECT 674.400 773.400 676.200 780.300 ;
        RECT 680.400 773.400 682.200 780.300 ;
        RECT 695.400 773.400 697.200 780.300 ;
        RECT 702.900 767.400 704.700 780.300 ;
        RECT 711.300 767.400 713.100 780.300 ;
        RECT 718.800 773.400 720.600 780.300 ;
        RECT 734.400 769.200 736.200 780.300 ;
        RECT 753.300 767.400 755.100 780.300 ;
        RECT 760.800 773.400 762.600 780.300 ;
        RECT 778.800 774.000 780.600 780.300 ;
        RECT 784.800 773.400 786.600 780.300 ;
        RECT 797.400 769.200 799.200 780.300 ;
        RECT 816.300 767.400 818.100 780.300 ;
        RECT 823.800 773.400 825.600 780.300 ;
        RECT 13.800 704.700 15.600 711.000 ;
        RECT 19.800 704.700 21.600 711.600 ;
        RECT 32.400 704.700 34.200 715.800 ;
        RECT 55.800 704.700 57.600 711.000 ;
        RECT 61.800 704.700 63.600 711.600 ;
        RECT 76.800 704.700 78.600 711.000 ;
        RECT 82.800 704.700 84.600 711.600 ;
        RECT 95.400 704.700 97.200 715.800 ;
        RECT 113.400 704.700 115.200 711.600 ;
        RECT 120.900 704.700 122.700 717.600 ;
        RECT 133.200 704.700 135.000 717.600 ;
        RECT 139.800 704.700 141.600 711.600 ;
        RECT 154.500 704.700 156.300 717.600 ;
        RECT 170.400 704.700 172.200 711.600 ;
        RECT 177.900 704.700 179.700 717.600 ;
        RECT 186.300 704.700 188.100 717.600 ;
        RECT 193.800 704.700 195.600 711.600 ;
        RECT 208.800 704.700 210.600 711.000 ;
        RECT 214.800 704.700 216.600 711.600 ;
        RECT 221.400 704.700 223.200 711.600 ;
        RECT 227.400 704.700 229.200 711.000 ;
        RECT 242.400 704.700 244.200 715.800 ;
        RECT 261.300 704.700 263.100 717.600 ;
        RECT 268.800 704.700 270.600 711.600 ;
        RECT 289.800 704.700 291.600 715.800 ;
        RECT 302.400 704.700 304.200 711.600 ;
        RECT 308.400 704.700 310.200 711.000 ;
        RECT 328.200 704.700 330.000 717.600 ;
        RECT 334.800 704.700 336.600 711.600 ;
        RECT 344.400 704.700 346.200 711.600 ;
        RECT 350.400 704.700 352.200 711.600 ;
        RECT 367.800 704.700 369.600 711.000 ;
        RECT 373.800 704.700 375.600 711.600 ;
        RECT 388.800 704.700 390.600 711.000 ;
        RECT 394.800 704.700 396.600 711.600 ;
        RECT 405.300 704.700 407.100 717.600 ;
        RECT 412.800 704.700 414.600 711.600 ;
        RECT 424.800 704.700 426.600 711.600 ;
        RECT 430.800 704.700 432.600 711.600 ;
        RECT 442.200 704.700 444.000 717.600 ;
        RECT 448.800 704.700 450.600 711.600 ;
        RECT 469.800 704.700 471.600 715.500 ;
        RECT 482.400 704.700 484.200 711.600 ;
        RECT 489.000 704.700 490.800 717.600 ;
        RECT 505.200 704.700 507.000 717.600 ;
        RECT 511.800 704.700 513.600 711.600 ;
        RECT 518.400 704.700 520.200 711.600 ;
        RECT 525.000 704.700 526.800 717.600 ;
        RECT 550.800 704.700 552.600 715.500 ;
        RECT 563.400 704.700 565.200 711.600 ;
        RECT 570.000 704.700 571.800 717.600 ;
        RECT 584.400 704.700 586.200 711.600 ;
        RECT 590.400 704.700 592.200 711.600 ;
        RECT 607.800 704.700 609.600 715.800 ;
        RECT 620.400 704.700 622.200 711.600 ;
        RECT 627.000 704.700 628.800 717.600 ;
        RECT 649.800 704.700 651.600 717.600 ;
        RECT 659.400 704.700 661.200 711.600 ;
        RECT 665.400 704.700 667.200 711.600 ;
        RECT 680.400 704.700 682.200 715.800 ;
        RECT 695.400 704.700 697.200 711.600 ;
        RECT 715.800 704.700 717.600 711.600 ;
        RECT 722.400 704.700 724.200 711.600 ;
        RECT 742.800 704.700 744.600 711.000 ;
        RECT 748.800 704.700 750.600 711.600 ;
        RECT 758.400 704.700 760.200 711.600 ;
        RECT 764.400 704.700 766.200 711.000 ;
        RECT 779.400 704.700 781.200 711.600 ;
        RECT 785.400 704.700 787.200 711.000 ;
        RECT 799.800 704.700 801.600 711.600 ;
        RECT 805.800 704.700 807.600 711.600 ;
        RECT 817.800 704.700 819.600 711.000 ;
        RECT 823.800 704.700 825.600 711.600 ;
        RECT -9.450 702.300 830.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT 10.800 695.400 12.600 702.300 ;
        RECT 16.800 695.400 18.600 702.300 ;
        RECT 23.400 695.400 25.200 702.300 ;
        RECT 29.400 696.000 31.200 702.300 ;
        RECT 44.400 691.200 46.200 702.300 ;
        RECT 63.300 689.400 65.100 702.300 ;
        RECT 70.800 695.400 72.600 702.300 ;
        RECT 91.800 691.200 93.600 702.300 ;
        RECT 104.400 695.400 106.200 702.300 ;
        RECT 121.200 689.400 123.000 702.300 ;
        RECT 127.800 695.400 129.600 702.300 ;
        RECT 134.400 695.400 136.200 702.300 ;
        RECT 140.400 695.400 142.200 702.300 ;
        RECT 157.800 696.000 159.600 702.300 ;
        RECT 163.800 695.400 165.600 702.300 ;
        RECT 178.800 696.000 180.600 702.300 ;
        RECT 184.800 695.400 186.600 702.300 ;
        RECT 194.400 691.200 196.200 702.300 ;
        RECT 220.800 691.200 222.600 702.300 ;
        RECT 235.800 696.000 237.600 702.300 ;
        RECT 241.800 695.400 243.600 702.300 ;
        RECT 251.400 695.400 253.200 702.300 ;
        RECT 266.400 691.500 268.200 702.300 ;
        RECT 287.400 689.400 289.200 702.300 ;
        RECT 302.400 695.400 304.200 702.300 ;
        RECT 308.400 696.000 310.200 702.300 ;
        RECT 322.800 695.400 324.600 702.300 ;
        RECT 328.800 695.400 330.600 702.300 ;
        RECT 340.800 695.400 342.600 702.300 ;
        RECT 346.800 695.400 348.600 702.300 ;
        RECT 361.800 691.200 363.600 702.300 ;
        RECT 379.800 696.000 381.600 702.300 ;
        RECT 385.800 695.400 387.600 702.300 ;
        RECT 396.300 689.400 398.100 702.300 ;
        RECT 403.800 695.400 405.600 702.300 ;
        RECT 417.300 689.400 419.100 702.300 ;
        RECT 424.800 695.400 426.600 702.300 ;
        RECT 442.800 696.000 444.600 702.300 ;
        RECT 448.800 695.400 450.600 702.300 ;
        RECT 457.800 695.400 459.600 702.300 ;
        RECT 463.800 695.400 465.600 702.300 ;
        RECT 473.700 689.400 475.500 702.300 ;
        RECT 485.400 689.400 487.200 702.300 ;
        RECT 502.500 689.400 504.300 702.300 ;
        RECT 516.300 689.400 518.100 702.300 ;
        RECT 523.800 695.400 525.600 702.300 ;
        RECT 547.800 691.500 549.600 702.300 ;
        RECT 560.400 695.400 562.200 702.300 ;
        RECT 566.400 695.400 568.200 702.300 ;
        RECT 580.800 695.400 582.600 702.300 ;
        RECT 591.300 689.400 593.100 702.300 ;
        RECT 598.800 695.400 600.600 702.300 ;
        RECT 616.800 695.400 618.600 702.300 ;
        RECT 624.300 689.400 626.100 702.300 ;
        RECT 631.800 695.400 633.600 702.300 ;
        RECT 646.800 696.000 648.600 702.300 ;
        RECT 652.800 695.400 654.600 702.300 ;
        RECT 659.400 695.400 661.200 702.300 ;
        RECT 665.400 696.000 667.200 702.300 ;
        RECT 680.400 695.400 682.200 702.300 ;
        RECT 686.400 696.000 688.200 702.300 ;
        RECT 701.400 695.400 703.200 702.300 ;
        RECT 707.400 696.000 709.200 702.300 ;
        RECT 719.400 695.400 721.200 702.300 ;
        RECT 725.400 696.000 727.200 702.300 ;
        RECT 743.400 691.500 745.200 702.300 ;
        RECT 769.800 689.400 771.600 702.300 ;
        RECT 780.300 689.400 782.100 702.300 ;
        RECT 787.800 695.400 789.600 702.300 ;
        RECT 802.800 695.400 804.600 702.300 ;
        RECT 808.800 695.400 810.600 702.300 ;
        RECT 818.400 691.200 820.200 702.300 ;
        RECT 10.800 626.700 12.600 633.600 ;
        RECT 16.800 626.700 18.600 633.600 ;
        RECT 31.800 626.700 33.600 633.000 ;
        RECT 37.800 626.700 39.600 633.600 ;
        RECT 47.400 626.700 49.200 633.600 ;
        RECT 53.400 626.700 55.200 633.000 ;
        RECT 65.400 626.700 67.200 633.600 ;
        RECT 83.400 626.700 85.200 637.800 ;
        RECT 106.800 626.700 108.600 633.600 ;
        RECT 119.400 626.700 121.200 633.600 ;
        RECT 126.900 626.700 128.700 639.600 ;
        RECT 145.800 626.700 147.600 639.600 ;
        RECT 154.800 626.700 156.600 633.600 ;
        RECT 160.800 626.700 162.600 633.600 ;
        RECT 169.800 626.700 171.600 633.600 ;
        RECT 175.800 626.700 177.600 633.600 ;
        RECT 190.500 626.700 192.300 639.600 ;
        RECT 206.400 626.700 208.200 633.600 ;
        RECT 213.900 626.700 215.700 639.600 ;
        RECT 227.400 626.700 229.200 633.600 ;
        RECT 234.900 626.700 236.700 639.600 ;
        RECT 245.400 626.700 247.200 633.600 ;
        RECT 252.900 626.700 254.700 639.600 ;
        RECT 265.800 626.700 267.600 633.600 ;
        RECT 271.800 626.700 273.600 633.600 ;
        RECT 284.400 626.700 286.200 633.600 ;
        RECT 291.900 626.700 293.700 639.600 ;
        RECT 302.400 626.700 304.200 633.600 ;
        RECT 314.400 626.700 316.200 633.600 ;
        RECT 320.400 626.700 322.200 633.000 ;
        RECT 340.800 626.700 342.600 633.600 ;
        RECT 347.400 626.700 349.200 633.600 ;
        RECT 353.400 626.700 355.200 633.600 ;
        RECT 367.800 626.700 369.600 639.600 ;
        RECT 376.800 626.700 378.600 633.600 ;
        RECT 382.800 626.700 384.600 633.600 ;
        RECT 397.800 626.700 399.600 633.600 ;
        RECT 407.400 626.700 409.200 633.600 ;
        RECT 413.400 626.700 415.200 633.000 ;
        RECT 433.800 626.700 435.600 633.000 ;
        RECT 439.800 626.700 441.600 633.600 ;
        RECT 446.400 626.700 448.200 633.600 ;
        RECT 452.400 626.700 454.200 633.600 ;
        RECT 475.800 626.700 477.600 637.500 ;
        RECT 493.800 626.700 495.600 633.600 ;
        RECT 500.400 626.700 502.200 633.600 ;
        RECT 516.300 626.700 518.100 639.600 ;
        RECT 526.800 626.700 528.600 639.600 ;
        RECT 536.400 626.700 538.200 639.600 ;
        RECT 554.400 626.700 556.200 637.800 ;
        RECT 572.400 626.700 574.200 633.600 ;
        RECT 578.400 626.700 580.200 633.000 ;
        RECT 590.400 626.700 592.200 633.600 ;
        RECT 596.400 626.700 598.200 633.600 ;
        RECT 609.300 626.700 611.100 639.600 ;
        RECT 616.800 626.700 618.600 633.600 ;
        RECT 626.400 626.700 628.200 633.600 ;
        RECT 641.400 626.700 643.200 633.600 ;
        RECT 647.400 626.700 649.200 633.600 ;
        RECT 664.800 626.700 666.600 633.600 ;
        RECT 675.300 626.700 677.100 639.600 ;
        RECT 682.800 626.700 684.600 633.600 ;
        RECT 693.300 626.700 695.100 639.600 ;
        RECT 700.800 626.700 702.600 633.600 ;
        RECT 718.800 626.700 720.600 633.600 ;
        RECT 728.400 626.700 730.200 633.600 ;
        RECT 734.400 626.700 736.200 633.000 ;
        RECT 754.800 626.700 756.600 633.000 ;
        RECT 760.800 626.700 762.600 633.600 ;
        RECT 769.800 626.700 771.600 633.600 ;
        RECT 775.800 626.700 777.600 633.600 ;
        RECT 790.800 626.700 792.600 639.600 ;
        RECT 799.800 626.700 801.600 633.600 ;
        RECT 805.800 626.700 807.600 633.600 ;
        RECT 815.400 626.700 817.200 633.600 ;
        RECT 821.400 626.700 823.200 633.000 ;
        RECT -9.450 624.300 830.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT 7.800 617.400 9.600 624.300 ;
        RECT 13.800 617.400 15.600 624.300 ;
        RECT 28.800 618.000 30.600 624.300 ;
        RECT 34.800 617.400 36.600 624.300 ;
        RECT 49.800 617.400 51.600 624.300 ;
        RECT 64.800 618.000 66.600 624.300 ;
        RECT 70.800 617.400 72.600 624.300 ;
        RECT 83.400 617.400 85.200 624.300 ;
        RECT 90.900 611.400 92.700 624.300 ;
        RECT 101.400 617.400 103.200 624.300 ;
        RECT 107.400 618.000 109.200 624.300 ;
        RECT 122.400 617.400 124.200 624.300 ;
        RECT 128.400 617.400 130.200 624.300 ;
        RECT 138.300 611.400 140.100 624.300 ;
        RECT 145.800 617.400 147.600 624.300 ;
        RECT 158.400 613.500 160.200 624.300 ;
        RECT 182.400 613.500 184.200 624.300 ;
        RECT 200.400 611.400 202.200 624.300 ;
        RECT 215.400 617.400 217.200 624.300 ;
        RECT 221.400 618.000 223.200 624.300 ;
        RECT 241.800 617.400 243.600 624.300 ;
        RECT 248.400 617.400 250.200 624.300 ;
        RECT 254.400 618.000 256.200 624.300 ;
        RECT 269.400 617.400 271.200 624.300 ;
        RECT 275.400 617.400 277.200 624.300 ;
        RECT 290.400 617.400 292.200 624.300 ;
        RECT 297.900 611.400 299.700 624.300 ;
        RECT 313.200 611.400 315.000 624.300 ;
        RECT 319.800 617.400 321.600 624.300 ;
        RECT 326.400 617.400 328.200 624.300 ;
        RECT 332.400 617.400 334.200 624.300 ;
        RECT 346.800 618.000 348.600 624.300 ;
        RECT 352.800 617.400 354.600 624.300 ;
        RECT 362.400 617.400 364.200 624.300 ;
        RECT 368.400 617.400 370.200 624.300 ;
        RECT 378.300 611.400 380.100 624.300 ;
        RECT 385.800 617.400 387.600 624.300 ;
        RECT 403.200 611.400 405.000 624.300 ;
        RECT 409.800 617.400 411.600 624.300 ;
        RECT 417.300 611.400 419.100 624.300 ;
        RECT 424.800 617.400 426.600 624.300 ;
        RECT 434.400 617.400 436.200 624.300 ;
        RECT 440.400 617.400 442.200 624.300 ;
        RECT 450.300 611.400 452.100 624.300 ;
        RECT 457.800 617.400 459.600 624.300 ;
        RECT 475.200 611.400 477.000 624.300 ;
        RECT 481.800 617.400 483.600 624.300 ;
        RECT 493.800 617.400 495.600 624.300 ;
        RECT 499.800 617.400 501.600 624.300 ;
        RECT 509.400 611.400 511.200 624.300 ;
        RECT 525.300 611.400 527.100 624.300 ;
        RECT 532.800 617.400 534.600 624.300 ;
        RECT 547.800 617.400 549.600 624.300 ;
        RECT 553.800 617.400 555.600 624.300 ;
        RECT 563.400 617.400 565.200 624.300 ;
        RECT 569.400 618.000 571.200 624.300 ;
        RECT 586.800 611.400 588.600 624.300 ;
        RECT 595.800 617.400 597.600 624.300 ;
        RECT 601.800 617.400 603.600 624.300 ;
        RECT 613.800 617.400 615.600 624.300 ;
        RECT 619.800 617.400 621.600 624.300 ;
        RECT 629.400 617.400 631.200 624.300 ;
        RECT 635.400 618.000 637.200 624.300 ;
        RECT 650.400 613.200 652.200 624.300 ;
        RECT 671.400 613.200 673.200 624.300 ;
        RECT 689.400 617.400 691.200 624.300 ;
        RECT 695.400 618.000 697.200 624.300 ;
        RECT 718.800 613.200 720.600 624.300 ;
        RECT 733.800 617.400 735.600 624.300 ;
        RECT 746.400 617.400 748.200 624.300 ;
        RECT 753.900 611.400 755.700 624.300 ;
        RECT 766.800 617.400 768.600 624.300 ;
        RECT 773.400 617.400 775.200 624.300 ;
        RECT 788.400 617.400 790.200 624.300 ;
        RECT 794.400 618.000 796.200 624.300 ;
        RECT 811.800 618.000 813.600 624.300 ;
        RECT 817.800 617.400 819.600 624.300 ;
        RECT 13.800 548.700 15.600 559.800 ;
        RECT 28.800 548.700 30.600 555.000 ;
        RECT 34.800 548.700 36.600 555.600 ;
        RECT 49.800 548.700 51.600 559.800 ;
        RECT 61.800 548.700 63.600 555.600 ;
        RECT 67.800 548.700 69.600 555.600 ;
        RECT 85.800 548.700 87.600 559.800 ;
        RECT 103.800 548.700 105.600 555.000 ;
        RECT 109.800 548.700 111.600 555.600 ;
        RECT 121.200 548.700 123.000 561.600 ;
        RECT 127.800 548.700 129.600 555.600 ;
        RECT 136.800 548.700 138.600 555.600 ;
        RECT 142.800 548.700 144.600 555.600 ;
        RECT 157.500 548.700 159.300 561.600 ;
        RECT 170.400 548.700 172.200 555.600 ;
        RECT 177.000 548.700 178.800 561.600 ;
        RECT 190.800 548.700 192.600 555.600 ;
        RECT 196.800 548.700 198.600 555.600 ;
        RECT 207.300 548.700 209.100 561.600 ;
        RECT 214.800 548.700 216.600 555.600 ;
        RECT 227.400 548.700 229.200 555.600 ;
        RECT 233.400 548.700 235.200 555.600 ;
        RECT 248.400 548.700 250.200 555.600 ;
        RECT 255.900 548.700 257.700 561.600 ;
        RECT 263.400 548.700 265.200 561.600 ;
        RECT 275.400 548.700 277.200 561.600 ;
        RECT 292.800 548.700 294.600 561.600 ;
        RECT 302.400 548.700 304.200 555.600 ;
        RECT 309.000 548.700 310.800 561.600 ;
        RECT 326.400 548.700 328.200 555.600 ;
        RECT 333.900 548.700 335.700 561.600 ;
        RECT 346.800 548.700 348.600 555.600 ;
        RECT 352.800 548.700 354.600 555.600 ;
        RECT 362.400 548.700 364.200 555.600 ;
        RECT 369.900 548.700 371.700 561.600 ;
        RECT 385.200 548.700 387.000 561.600 ;
        RECT 391.800 548.700 393.600 555.600 ;
        RECT 401.400 548.700 403.200 555.600 ;
        RECT 408.900 548.700 410.700 561.600 ;
        RECT 418.800 548.700 420.600 555.600 ;
        RECT 424.800 548.700 426.600 555.600 ;
        RECT 437.400 548.700 439.200 555.600 ;
        RECT 444.900 548.700 446.700 561.600 ;
        RECT 460.800 548.700 462.600 561.600 ;
        RECT 472.800 548.700 474.600 555.600 ;
        RECT 478.800 548.700 480.600 555.600 ;
        RECT 489.300 548.700 491.100 561.600 ;
        RECT 496.800 548.700 498.600 555.600 ;
        RECT 514.800 548.700 516.600 561.600 ;
        RECT 524.400 548.700 526.200 555.600 ;
        RECT 531.900 548.700 533.700 561.600 ;
        RECT 545.400 548.700 547.200 555.600 ;
        RECT 552.900 548.700 554.700 561.600 ;
        RECT 564.300 548.700 566.100 561.600 ;
        RECT 571.800 548.700 573.600 555.600 ;
        RECT 587.400 548.700 589.200 555.600 ;
        RECT 594.900 548.700 596.700 561.600 ;
        RECT 606.900 548.700 608.700 561.600 ;
        RECT 621.300 548.700 623.100 561.600 ;
        RECT 628.800 548.700 630.600 555.600 ;
        RECT 638.400 548.700 640.200 555.600 ;
        RECT 644.400 548.700 646.200 555.600 ;
        RECT 657.300 548.700 659.100 561.600 ;
        RECT 664.800 548.700 666.600 555.600 ;
        RECT 680.700 548.700 682.500 561.600 ;
        RECT 692.400 548.700 694.200 555.600 ;
        RECT 698.400 548.700 700.200 555.600 ;
        RECT 718.800 548.700 720.600 561.600 ;
        RECT 725.400 548.700 727.200 555.600 ;
        RECT 732.000 548.700 733.800 561.600 ;
        RECT 751.800 548.700 753.600 555.600 ;
        RECT 761.400 548.700 763.200 555.600 ;
        RECT 776.400 548.700 778.200 561.600 ;
        RECT 791.400 548.700 793.200 561.600 ;
        RECT 809.400 548.700 811.200 561.600 ;
        RECT -9.450 546.300 830.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT 16.800 535.200 18.600 546.300 ;
        RECT 29.400 539.400 31.200 546.300 ;
        RECT 35.400 540.000 37.200 546.300 ;
        RECT 52.800 539.400 54.600 546.300 ;
        RECT 65.400 539.400 67.200 546.300 ;
        RECT 72.900 533.400 74.700 546.300 ;
        RECT 81.300 533.400 83.100 546.300 ;
        RECT 88.800 539.400 90.600 546.300 ;
        RECT 104.400 539.400 106.200 546.300 ;
        RECT 111.900 533.400 113.700 546.300 ;
        RECT 120.300 533.400 122.100 546.300 ;
        RECT 127.800 539.400 129.600 546.300 ;
        RECT 142.800 539.400 144.600 546.300 ;
        RECT 148.800 539.400 150.600 546.300 ;
        RECT 166.800 535.200 168.600 546.300 ;
        RECT 182.400 539.400 184.200 546.300 ;
        RECT 189.900 533.400 191.700 546.300 ;
        RECT 200.400 539.400 202.200 546.300 ;
        RECT 206.400 539.400 208.200 546.300 ;
        RECT 219.300 533.400 221.100 546.300 ;
        RECT 226.800 539.400 228.600 546.300 ;
        RECT 241.500 533.400 243.300 546.300 ;
        RECT 252.300 533.400 254.100 546.300 ;
        RECT 259.800 539.400 261.600 546.300 ;
        RECT 272.400 539.400 274.200 546.300 ;
        RECT 279.900 533.400 281.700 546.300 ;
        RECT 289.800 539.400 291.600 546.300 ;
        RECT 295.800 539.400 297.600 546.300 ;
        RECT 302.400 539.400 304.200 546.300 ;
        RECT 308.400 539.400 310.200 546.300 ;
        RECT 320.400 539.400 322.200 546.300 ;
        RECT 326.400 539.400 328.200 546.300 ;
        RECT 341.400 539.400 343.200 546.300 ;
        RECT 348.900 533.400 350.700 546.300 ;
        RECT 361.800 539.400 363.600 546.300 ;
        RECT 367.800 539.400 369.600 546.300 ;
        RECT 378.300 533.400 380.100 546.300 ;
        RECT 385.800 539.400 387.600 546.300 ;
        RECT 396.150 539.400 397.950 546.300 ;
        RECT 406.350 539.400 408.150 546.300 ;
        RECT 412.950 539.400 414.750 546.300 ;
        RECT 421.650 542.400 423.450 546.300 ;
        RECT 434.400 539.400 436.200 546.300 ;
        RECT 440.400 539.400 442.200 546.300 ;
        RECT 452.400 539.400 454.200 546.300 ;
        RECT 459.900 533.400 461.700 546.300 ;
        RECT 468.150 539.400 469.950 546.300 ;
        RECT 478.350 539.400 480.150 546.300 ;
        RECT 484.950 539.400 486.750 546.300 ;
        RECT 493.650 542.400 495.450 546.300 ;
        RECT 504.150 539.400 505.950 546.300 ;
        RECT 514.350 539.400 516.150 546.300 ;
        RECT 520.950 539.400 522.750 546.300 ;
        RECT 529.650 542.400 531.450 546.300 ;
        RECT 544.800 539.400 546.600 546.300 ;
        RECT 550.800 539.400 552.600 546.300 ;
        RECT 557.400 539.400 559.200 546.300 ;
        RECT 564.000 533.400 565.800 546.300 ;
        RECT 575.400 539.400 577.200 546.300 ;
        RECT 581.400 540.000 583.200 546.300 ;
        RECT 593.400 539.400 595.200 546.300 ;
        RECT 599.400 539.400 601.200 546.300 ;
        RECT 608.400 539.400 610.200 546.300 ;
        RECT 614.400 539.400 616.200 546.300 ;
        RECT 627.300 533.400 629.100 546.300 ;
        RECT 634.800 539.400 636.600 546.300 ;
        RECT 647.400 539.400 649.200 546.300 ;
        RECT 654.000 533.400 655.800 546.300 ;
        RECT 670.800 539.400 672.600 546.300 ;
        RECT 676.800 539.400 678.600 546.300 ;
        RECT 687.900 533.400 689.700 546.300 ;
        RECT 712.800 535.200 714.600 546.300 ;
        RECT 730.800 533.400 732.600 546.300 ;
        RECT 738.300 533.400 740.100 546.300 ;
        RECT 745.800 539.400 747.600 546.300 ;
        RECT 761.400 535.200 763.200 546.300 ;
        RECT 776.400 539.400 778.200 546.300 ;
        RECT 782.400 539.400 784.200 546.300 ;
        RECT 799.800 540.000 801.600 546.300 ;
        RECT 805.800 539.400 807.600 546.300 ;
        RECT 818.700 533.400 820.500 546.300 ;
        RECT 6.300 470.700 8.100 483.600 ;
        RECT 13.800 470.700 15.600 477.600 ;
        RECT 31.800 470.700 33.600 477.600 ;
        RECT 38.400 470.700 40.200 477.600 ;
        RECT 44.400 470.700 46.200 477.000 ;
        RECT 64.800 470.700 66.600 477.600 ;
        RECT 79.800 470.700 81.600 481.800 ;
        RECT 97.800 470.700 99.600 477.000 ;
        RECT 103.800 470.700 105.600 477.600 ;
        RECT 121.800 470.700 123.600 481.800 ;
        RECT 131.400 470.700 133.200 477.600 ;
        RECT 146.400 470.700 148.200 477.600 ;
        RECT 169.800 470.700 171.600 483.600 ;
        RECT 179.400 470.700 181.200 477.600 ;
        RECT 185.400 470.700 187.200 477.600 ;
        RECT 202.800 470.700 204.600 477.000 ;
        RECT 208.800 470.700 210.600 477.600 ;
        RECT 218.400 470.700 220.200 477.600 ;
        RECT 224.400 470.700 226.200 477.600 ;
        RECT 238.200 470.700 240.000 483.600 ;
        RECT 244.800 470.700 246.600 477.600 ;
        RECT 254.400 470.700 256.200 477.600 ;
        RECT 271.800 470.700 273.600 477.600 ;
        RECT 283.800 470.700 285.600 477.000 ;
        RECT 289.800 470.700 291.600 477.600 ;
        RECT 299.400 470.700 301.200 477.600 ;
        RECT 305.400 470.700 307.200 477.600 ;
        RECT 315.300 470.700 317.100 483.600 ;
        RECT 322.800 470.700 324.600 477.600 ;
        RECT 332.400 470.700 334.200 477.600 ;
        RECT 338.400 470.700 340.200 477.600 ;
        RECT 347.550 470.700 349.350 474.600 ;
        RECT 356.250 470.700 358.050 477.600 ;
        RECT 362.850 470.700 364.650 477.600 ;
        RECT 373.050 470.700 374.850 477.600 ;
        RECT 387.300 470.700 389.100 483.600 ;
        RECT 394.800 470.700 396.600 477.600 ;
        RECT 406.800 470.700 408.600 477.600 ;
        RECT 412.800 470.700 414.600 477.600 ;
        RECT 421.800 470.700 423.600 477.600 ;
        RECT 427.800 470.700 429.600 477.600 ;
        RECT 437.400 470.700 439.200 477.600 ;
        RECT 443.400 470.700 445.200 477.600 ;
        RECT 454.800 470.700 456.600 477.600 ;
        RECT 460.800 470.700 462.600 477.600 ;
        RECT 470.400 470.700 472.200 477.600 ;
        RECT 477.900 470.700 479.700 483.600 ;
        RECT 491.400 470.700 493.200 477.600 ;
        RECT 498.900 470.700 500.700 483.600 ;
        RECT 510.300 470.700 512.100 483.600 ;
        RECT 517.800 470.700 519.600 477.600 ;
        RECT 527.400 470.700 529.200 483.600 ;
        RECT 545.400 470.700 547.200 481.800 ;
        RECT 560.400 470.700 562.200 483.600 ;
        RECT 578.400 470.700 580.200 477.600 ;
        RECT 595.800 470.700 597.600 477.600 ;
        RECT 601.800 470.700 603.600 477.600 ;
        RECT 616.800 470.700 618.600 477.600 ;
        RECT 623.400 470.700 625.200 477.600 ;
        RECT 629.400 470.700 631.200 477.000 ;
        RECT 649.800 470.700 651.600 477.600 ;
        RECT 657.300 470.700 659.100 483.600 ;
        RECT 664.800 470.700 666.600 477.600 ;
        RECT 675.300 470.700 677.100 483.600 ;
        RECT 682.800 470.700 684.600 477.600 ;
        RECT 697.800 470.700 699.600 477.000 ;
        RECT 703.800 470.700 705.600 477.600 ;
        RECT 714.300 470.700 716.100 483.600 ;
        RECT 721.800 470.700 723.600 477.600 ;
        RECT 739.800 470.700 741.600 477.600 ;
        RECT 749.400 470.700 751.200 477.600 ;
        RECT 755.400 470.700 757.200 477.600 ;
        RECT 768.300 470.700 770.100 483.600 ;
        RECT 775.800 470.700 777.600 477.600 ;
        RECT 787.800 470.700 789.600 477.600 ;
        RECT 793.800 470.700 795.600 477.600 ;
        RECT 805.800 470.700 807.600 477.000 ;
        RECT 811.800 470.700 813.600 477.600 ;
        RECT 821.400 470.700 823.200 477.600 ;
        RECT -9.450 468.300 830.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT 10.800 462.000 12.600 468.300 ;
        RECT 16.800 461.400 18.600 468.300 ;
        RECT 26.400 457.200 28.200 468.300 ;
        RECT 47.400 461.400 49.200 468.300 ;
        RECT 54.900 455.400 56.700 468.300 ;
        RECT 67.800 462.000 69.600 468.300 ;
        RECT 73.800 461.400 75.600 468.300 ;
        RECT 88.800 462.000 90.600 468.300 ;
        RECT 94.800 461.400 96.600 468.300 ;
        RECT 107.400 461.400 109.200 468.300 ;
        RECT 114.900 455.400 116.700 468.300 ;
        RECT 126.300 455.400 128.100 468.300 ;
        RECT 133.800 461.400 135.600 468.300 ;
        RECT 151.800 461.400 153.600 468.300 ;
        RECT 161.400 461.400 163.200 468.300 ;
        RECT 168.900 455.400 170.700 468.300 ;
        RECT 176.400 455.400 178.200 468.300 ;
        RECT 194.400 461.400 196.200 468.300 ;
        RECT 200.400 461.400 202.200 468.300 ;
        RECT 212.400 461.400 214.200 468.300 ;
        RECT 218.400 461.400 220.200 468.300 ;
        RECT 233.400 457.500 235.200 468.300 ;
        RECT 256.800 461.400 258.600 468.300 ;
        RECT 263.400 461.400 265.200 468.300 ;
        RECT 270.000 455.400 271.800 468.300 ;
        RECT 292.800 457.200 294.600 468.300 ;
        RECT 305.400 461.400 307.200 468.300 ;
        RECT 311.400 462.000 313.200 468.300 ;
        RECT 324.300 455.400 326.100 468.300 ;
        RECT 331.800 461.400 333.600 468.300 ;
        RECT 341.550 464.400 343.350 468.300 ;
        RECT 350.250 461.400 352.050 468.300 ;
        RECT 356.850 461.400 358.650 468.300 ;
        RECT 367.050 461.400 368.850 468.300 ;
        RECT 380.700 455.400 382.500 468.300 ;
        RECT 393.150 461.400 394.950 468.300 ;
        RECT 403.350 461.400 405.150 468.300 ;
        RECT 409.950 461.400 411.750 468.300 ;
        RECT 418.650 464.400 420.450 468.300 ;
        RECT 434.700 455.400 436.500 468.300 ;
        RECT 447.150 461.400 448.950 468.300 ;
        RECT 457.350 461.400 459.150 468.300 ;
        RECT 463.950 461.400 465.750 468.300 ;
        RECT 472.650 464.400 474.450 468.300 ;
        RECT 487.800 461.400 489.600 468.300 ;
        RECT 493.800 461.400 495.600 468.300 ;
        RECT 504.300 455.400 506.100 468.300 ;
        RECT 511.800 461.400 513.600 468.300 ;
        RECT 521.400 455.400 523.200 468.300 ;
        RECT 534.150 461.400 535.950 468.300 ;
        RECT 544.350 461.400 546.150 468.300 ;
        RECT 550.950 461.400 552.750 468.300 ;
        RECT 559.650 464.400 561.450 468.300 ;
        RECT 573.300 455.400 575.100 468.300 ;
        RECT 580.800 461.400 582.600 468.300 ;
        RECT 593.400 455.400 595.200 468.300 ;
        RECT 599.400 455.400 601.200 468.300 ;
        RECT 605.400 455.400 607.200 468.300 ;
        RECT 611.400 455.400 613.200 468.300 ;
        RECT 617.400 455.400 619.200 468.300 ;
        RECT 632.400 461.400 634.200 468.300 ;
        RECT 639.900 455.400 641.700 468.300 ;
        RECT 655.800 461.400 657.600 468.300 ;
        RECT 662.400 461.400 664.200 468.300 ;
        RECT 668.400 461.400 670.200 468.300 ;
        RECT 680.400 461.400 682.200 468.300 ;
        RECT 686.400 461.400 688.200 468.300 ;
        RECT 699.900 455.400 701.700 468.300 ;
        RECT 716.400 461.400 718.200 468.300 ;
        RECT 731.400 455.400 733.200 468.300 ;
        RECT 754.800 455.400 756.600 468.300 ;
        RECT 764.400 457.200 766.200 468.300 ;
        RECT 782.400 461.400 784.200 468.300 ;
        RECT 797.400 461.400 799.200 468.300 ;
        RECT 803.400 462.000 805.200 468.300 ;
        RECT 821.700 455.400 823.500 468.300 ;
        RECT 13.800 392.700 15.600 399.600 ;
        RECT 28.800 392.700 30.600 403.800 ;
        RECT 43.800 392.700 45.600 399.000 ;
        RECT 49.800 392.700 51.600 399.600 ;
        RECT 70.800 392.700 72.600 403.500 ;
        RECT 80.400 392.700 82.200 399.600 ;
        RECT 86.400 392.700 88.200 399.600 ;
        RECT 100.800 392.700 102.600 399.000 ;
        RECT 106.800 392.700 108.600 399.600 ;
        RECT 121.800 392.700 123.600 403.800 ;
        RECT 139.800 392.700 141.600 399.600 ;
        RECT 149.400 392.700 151.200 399.600 ;
        RECT 156.900 392.700 158.700 405.600 ;
        RECT 172.800 392.700 174.600 405.600 ;
        RECT 179.400 392.700 181.200 399.600 ;
        RECT 185.400 392.700 187.200 399.600 ;
        RECT 200.400 392.700 202.200 399.600 ;
        RECT 207.900 392.700 209.700 405.600 ;
        RECT 218.400 392.700 220.200 405.600 ;
        RECT 233.400 392.700 235.200 399.600 ;
        RECT 246.300 392.700 248.100 405.600 ;
        RECT 253.800 392.700 255.600 399.600 ;
        RECT 269.400 392.700 271.200 399.600 ;
        RECT 276.900 392.700 278.700 405.600 ;
        RECT 287.400 392.700 289.200 405.600 ;
        RECT 303.300 392.700 305.100 405.600 ;
        RECT 310.800 392.700 312.600 399.600 ;
        RECT 323.400 392.700 325.200 399.600 ;
        RECT 329.400 392.700 331.200 399.600 ;
        RECT 339.150 392.700 340.950 399.600 ;
        RECT 349.350 392.700 351.150 399.600 ;
        RECT 355.950 392.700 357.750 399.600 ;
        RECT 364.650 392.700 366.450 396.600 ;
        RECT 376.800 392.700 378.600 405.600 ;
        RECT 382.800 392.700 384.600 405.600 ;
        RECT 388.800 392.700 390.600 405.600 ;
        RECT 394.800 392.700 396.600 405.600 ;
        RECT 400.800 392.700 402.600 405.600 ;
        RECT 407.400 392.700 409.200 399.600 ;
        RECT 413.400 392.700 415.200 399.600 ;
        RECT 428.400 392.700 430.200 399.600 ;
        RECT 435.900 392.700 437.700 405.600 ;
        RECT 445.800 392.700 447.600 399.600 ;
        RECT 451.800 392.700 453.600 399.600 ;
        RECT 466.500 392.700 468.300 405.600 ;
        RECT 482.400 392.700 484.200 399.600 ;
        RECT 489.900 392.700 491.700 405.600 ;
        RECT 498.150 392.700 499.950 399.600 ;
        RECT 508.350 392.700 510.150 399.600 ;
        RECT 514.950 392.700 516.750 399.600 ;
        RECT 523.650 392.700 525.450 396.600 ;
        RECT 541.800 392.700 543.600 399.600 ;
        RECT 548.400 392.700 550.200 405.600 ;
        RECT 571.800 392.700 573.600 399.600 ;
        RECT 581.400 392.700 583.200 405.600 ;
        RECT 597.150 392.700 598.950 399.600 ;
        RECT 607.350 392.700 609.150 399.600 ;
        RECT 613.950 392.700 615.750 399.600 ;
        RECT 622.650 392.700 624.450 396.600 ;
        RECT 636.300 392.700 638.100 405.600 ;
        RECT 646.800 392.700 648.600 405.600 ;
        RECT 661.800 392.700 663.600 399.600 ;
        RECT 668.550 392.700 670.350 396.600 ;
        RECT 677.250 392.700 679.050 399.600 ;
        RECT 683.850 392.700 685.650 399.600 ;
        RECT 694.050 392.700 695.850 399.600 ;
        RECT 710.400 392.700 712.200 399.600 ;
        RECT 717.900 392.700 719.700 405.600 ;
        RECT 733.800 392.700 735.600 399.600 ;
        RECT 754.800 392.700 756.600 403.500 ;
        RECT 765.150 392.700 766.950 399.600 ;
        RECT 775.350 392.700 777.150 399.600 ;
        RECT 781.950 392.700 783.750 399.600 ;
        RECT 790.650 392.700 792.450 396.600 ;
        RECT 803.400 392.700 805.200 399.600 ;
        RECT 818.400 392.700 820.200 399.600 ;
        RECT 824.400 392.700 826.200 399.600 ;
        RECT -9.450 390.300 830.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT 16.800 379.200 18.600 390.300 ;
        RECT 34.800 384.000 36.600 390.300 ;
        RECT 40.800 383.400 42.600 390.300 ;
        RECT 55.800 377.400 57.600 390.300 ;
        RECT 67.800 383.400 69.600 390.300 ;
        RECT 85.800 379.200 87.600 390.300 ;
        RECT 103.800 384.000 105.600 390.300 ;
        RECT 109.800 383.400 111.600 390.300 ;
        RECT 119.400 383.400 121.200 390.300 ;
        RECT 136.800 384.000 138.600 390.300 ;
        RECT 142.800 383.400 144.600 390.300 ;
        RECT 155.700 377.400 157.500 390.300 ;
        RECT 175.800 384.000 177.600 390.300 ;
        RECT 181.800 383.400 183.600 390.300 ;
        RECT 194.400 383.400 196.200 390.300 ;
        RECT 201.900 377.400 203.700 390.300 ;
        RECT 216.300 377.400 218.100 390.300 ;
        RECT 226.800 377.400 228.600 390.300 ;
        RECT 236.400 383.400 238.200 390.300 ;
        RECT 243.900 377.400 245.700 390.300 ;
        RECT 253.800 377.400 255.600 390.300 ;
        RECT 259.800 377.400 261.600 390.300 ;
        RECT 265.800 377.400 267.600 390.300 ;
        RECT 271.800 377.400 273.600 390.300 ;
        RECT 277.800 377.400 279.600 390.300 ;
        RECT 292.800 377.400 294.600 390.300 ;
        RECT 299.550 386.400 301.350 390.300 ;
        RECT 308.250 383.400 310.050 390.300 ;
        RECT 314.850 383.400 316.650 390.300 ;
        RECT 325.050 383.400 326.850 390.300 ;
        RECT 346.800 379.200 348.600 390.300 ;
        RECT 356.400 377.400 358.200 390.300 ;
        RECT 362.400 377.400 364.200 390.300 ;
        RECT 368.400 377.400 370.200 390.300 ;
        RECT 374.400 377.400 376.200 390.300 ;
        RECT 380.400 377.400 382.200 390.300 ;
        RECT 390.150 383.400 391.950 390.300 ;
        RECT 400.350 383.400 402.150 390.300 ;
        RECT 406.950 383.400 408.750 390.300 ;
        RECT 415.650 386.400 417.450 390.300 ;
        RECT 433.800 379.200 435.600 390.300 ;
        RECT 446.400 377.400 448.200 390.300 ;
        RECT 464.400 379.200 466.200 390.300 ;
        RECT 480.150 383.400 481.950 390.300 ;
        RECT 490.350 383.400 492.150 390.300 ;
        RECT 496.950 383.400 498.750 390.300 ;
        RECT 505.650 386.400 507.450 390.300 ;
        RECT 516.150 383.400 517.950 390.300 ;
        RECT 526.350 383.400 528.150 390.300 ;
        RECT 532.950 383.400 534.750 390.300 ;
        RECT 541.650 386.400 543.450 390.300 ;
        RECT 551.400 377.400 553.200 390.300 ;
        RECT 574.800 383.400 576.600 390.300 ;
        RECT 581.550 386.400 583.350 390.300 ;
        RECT 590.250 383.400 592.050 390.300 ;
        RECT 596.850 383.400 598.650 390.300 ;
        RECT 607.050 383.400 608.850 390.300 ;
        RECT 620.400 383.400 622.200 390.300 ;
        RECT 627.900 377.400 629.700 390.300 ;
        RECT 635.400 383.400 637.200 390.300 ;
        RECT 647.400 377.400 649.200 390.300 ;
        RECT 665.400 377.400 667.200 390.300 ;
        RECT 680.400 377.400 682.200 390.300 ;
        RECT 690.900 377.400 692.700 390.300 ;
        RECT 709.800 379.200 711.600 390.300 ;
        RECT 726.900 377.400 728.700 390.300 ;
        RECT 741.150 383.400 742.950 390.300 ;
        RECT 751.350 383.400 753.150 390.300 ;
        RECT 757.950 383.400 759.750 390.300 ;
        RECT 766.650 386.400 768.450 390.300 ;
        RECT 787.800 377.400 789.600 390.300 ;
        RECT 802.800 383.400 804.600 390.300 ;
        RECT 810.300 377.400 812.100 390.300 ;
        RECT 817.800 383.400 819.600 390.300 ;
        RECT 7.800 314.700 9.600 321.600 ;
        RECT 13.800 314.700 15.600 321.600 ;
        RECT 28.800 314.700 30.600 321.600 ;
        RECT 46.800 314.700 48.600 325.800 ;
        RECT 56.400 314.700 58.200 321.600 ;
        RECT 62.400 314.700 64.200 321.000 ;
        RECT 74.400 314.700 76.200 321.600 ;
        RECT 80.400 314.700 82.200 321.600 ;
        RECT 96.900 314.700 98.700 327.600 ;
        RECT 118.800 314.700 120.600 321.000 ;
        RECT 124.800 314.700 126.600 321.600 ;
        RECT 136.800 314.700 138.600 321.600 ;
        RECT 142.800 314.700 144.600 321.600 ;
        RECT 150.300 314.700 152.100 327.600 ;
        RECT 157.800 314.700 159.600 321.600 ;
        RECT 175.500 314.700 177.300 327.600 ;
        RECT 189.300 314.700 191.100 327.600 ;
        RECT 199.800 314.700 201.600 327.600 ;
        RECT 207.150 314.700 208.950 321.600 ;
        RECT 217.350 314.700 219.150 321.600 ;
        RECT 223.950 314.700 225.750 321.600 ;
        RECT 232.650 314.700 234.450 318.600 ;
        RECT 242.400 314.700 244.200 321.600 ;
        RECT 265.800 314.700 267.600 327.600 ;
        RECT 280.800 314.700 282.600 321.600 ;
        RECT 287.550 314.700 289.350 318.600 ;
        RECT 296.250 314.700 298.050 321.600 ;
        RECT 302.850 314.700 304.650 321.600 ;
        RECT 313.050 314.700 314.850 321.600 ;
        RECT 329.400 314.700 331.200 321.600 ;
        RECT 336.900 314.700 338.700 327.600 ;
        RECT 352.500 314.700 354.300 327.600 ;
        RECT 362.400 314.700 364.200 321.600 ;
        RECT 368.400 314.700 370.200 321.600 ;
        RECT 377.550 314.700 379.350 318.600 ;
        RECT 386.250 314.700 388.050 321.600 ;
        RECT 392.850 314.700 394.650 321.600 ;
        RECT 403.050 314.700 404.850 321.600 ;
        RECT 414.150 314.700 415.950 321.600 ;
        RECT 424.350 314.700 426.150 321.600 ;
        RECT 430.950 314.700 432.750 321.600 ;
        RECT 439.650 314.700 441.450 318.600 ;
        RECT 457.800 314.700 459.600 325.800 ;
        RECT 470.400 314.700 472.200 327.600 ;
        RECT 496.800 314.700 498.600 327.600 ;
        RECT 508.800 314.700 510.600 321.600 ;
        RECT 514.800 314.700 516.600 321.600 ;
        RECT 527.400 314.700 529.200 321.600 ;
        RECT 534.900 314.700 536.700 327.600 ;
        RECT 547.800 314.700 549.600 321.600 ;
        RECT 555.150 314.700 556.950 321.600 ;
        RECT 565.350 314.700 567.150 321.600 ;
        RECT 571.950 314.700 573.750 321.600 ;
        RECT 580.650 314.700 582.450 318.600 ;
        RECT 593.400 314.700 595.200 327.600 ;
        RECT 613.800 314.700 615.600 321.600 ;
        RECT 619.800 314.700 621.600 321.600 ;
        RECT 631.800 314.700 633.600 321.600 ;
        RECT 637.800 314.700 639.600 321.600 ;
        RECT 650.700 314.700 652.500 327.600 ;
        RECT 665.400 314.700 667.200 321.600 ;
        RECT 672.900 314.700 674.700 327.600 ;
        RECT 681.150 314.700 682.950 321.600 ;
        RECT 691.350 314.700 693.150 321.600 ;
        RECT 697.950 314.700 699.750 321.600 ;
        RECT 706.650 314.700 708.450 318.600 ;
        RECT 716.400 314.700 718.200 321.600 ;
        RECT 742.800 314.700 744.600 325.500 ;
        RECT 753.150 314.700 754.950 321.600 ;
        RECT 763.350 314.700 765.150 321.600 ;
        RECT 769.950 314.700 771.750 321.600 ;
        RECT 778.650 314.700 780.450 318.600 ;
        RECT 788.400 314.700 790.200 327.600 ;
        RECT 806.400 314.700 808.200 327.600 ;
        RECT -9.450 312.300 830.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT 6.150 305.400 7.950 312.300 ;
        RECT 16.350 305.400 18.150 312.300 ;
        RECT 22.950 305.400 24.750 312.300 ;
        RECT 31.650 308.400 33.450 312.300 ;
        RECT 41.400 305.400 43.200 312.300 ;
        RECT 47.400 305.400 49.200 312.300 ;
        RECT 56.550 308.400 58.350 312.300 ;
        RECT 65.250 305.400 67.050 312.300 ;
        RECT 71.850 305.400 73.650 312.300 ;
        RECT 82.050 305.400 83.850 312.300 ;
        RECT 96.300 299.400 98.100 312.300 ;
        RECT 103.800 305.400 105.600 312.300 ;
        RECT 116.400 305.400 118.200 312.300 ;
        RECT 123.900 299.400 125.700 312.300 ;
        RECT 136.800 305.400 138.600 312.300 ;
        RECT 143.550 308.400 145.350 312.300 ;
        RECT 152.250 305.400 154.050 312.300 ;
        RECT 158.850 305.400 160.650 312.300 ;
        RECT 169.050 305.400 170.850 312.300 ;
        RECT 180.150 305.400 181.950 312.300 ;
        RECT 190.350 305.400 192.150 312.300 ;
        RECT 196.950 305.400 198.750 312.300 ;
        RECT 205.650 308.400 207.450 312.300 ;
        RECT 216.150 305.400 217.950 312.300 ;
        RECT 226.350 305.400 228.150 312.300 ;
        RECT 232.950 305.400 234.750 312.300 ;
        RECT 241.650 308.400 243.450 312.300 ;
        RECT 251.400 305.400 253.200 312.300 ;
        RECT 274.800 299.400 276.600 312.300 ;
        RECT 289.800 299.400 291.600 312.300 ;
        RECT 307.800 299.400 309.600 312.300 ;
        RECT 322.800 305.400 324.600 312.300 ;
        RECT 329.550 308.400 331.350 312.300 ;
        RECT 338.250 305.400 340.050 312.300 ;
        RECT 344.850 305.400 346.650 312.300 ;
        RECT 355.050 305.400 356.850 312.300 ;
        RECT 369.300 299.400 371.100 312.300 ;
        RECT 376.800 305.400 378.600 312.300 ;
        RECT 390.300 299.400 392.100 312.300 ;
        RECT 397.800 305.400 399.600 312.300 ;
        RECT 413.400 305.400 415.200 312.300 ;
        RECT 420.900 299.400 422.700 312.300 ;
        RECT 428.400 305.400 430.200 312.300 ;
        RECT 434.400 305.400 436.200 312.300 ;
        RECT 444.300 299.400 446.100 312.300 ;
        RECT 451.800 305.400 453.600 312.300 ;
        RECT 461.550 308.400 463.350 312.300 ;
        RECT 470.250 305.400 472.050 312.300 ;
        RECT 476.850 305.400 478.650 312.300 ;
        RECT 487.050 305.400 488.850 312.300 ;
        RECT 497.400 305.400 499.200 312.300 ;
        RECT 503.400 305.400 505.200 312.300 ;
        RECT 523.800 299.400 525.600 312.300 ;
        RECT 533.400 301.200 535.200 312.300 ;
        RECT 551.700 299.400 553.500 312.300 ;
        RECT 566.400 305.400 568.200 312.300 ;
        RECT 573.900 299.400 575.700 312.300 ;
        RECT 584.400 305.400 586.200 312.300 ;
        RECT 590.400 305.400 592.200 312.300 ;
        RECT 599.400 299.400 601.200 312.300 ;
        RECT 617.400 299.400 619.200 312.300 ;
        RECT 635.400 301.200 637.200 312.300 ;
        RECT 656.400 305.400 658.200 312.300 ;
        RECT 663.900 299.400 665.700 312.300 ;
        RECT 676.200 299.400 678.000 312.300 ;
        RECT 682.800 305.400 684.600 312.300 ;
        RECT 700.800 299.400 702.600 312.300 ;
        RECT 707.400 299.400 709.200 312.300 ;
        RECT 723.300 299.400 725.100 312.300 ;
        RECT 730.800 305.400 732.600 312.300 ;
        RECT 746.400 305.400 748.200 312.300 ;
        RECT 753.900 299.400 755.700 312.300 ;
        RECT 764.400 299.400 766.200 312.300 ;
        RECT 782.400 305.400 784.200 312.300 ;
        RECT 796.800 305.400 798.600 312.300 ;
        RECT 802.800 305.400 804.600 312.300 ;
        RECT 813.300 299.400 815.100 312.300 ;
        RECT 820.800 305.400 822.600 312.300 ;
        RECT 6.150 236.700 7.950 243.600 ;
        RECT 16.350 236.700 18.150 243.600 ;
        RECT 22.950 236.700 24.750 243.600 ;
        RECT 31.650 236.700 33.450 240.600 ;
        RECT 47.400 236.700 49.200 243.600 ;
        RECT 54.900 236.700 56.700 249.600 ;
        RECT 65.400 236.700 67.200 243.600 ;
        RECT 80.400 236.700 82.200 243.600 ;
        RECT 93.150 236.700 94.950 243.600 ;
        RECT 103.350 236.700 105.150 243.600 ;
        RECT 109.950 236.700 111.750 243.600 ;
        RECT 118.650 236.700 120.450 240.600 ;
        RECT 131.400 236.700 133.200 243.600 ;
        RECT 144.150 236.700 145.950 243.600 ;
        RECT 154.350 236.700 156.150 243.600 ;
        RECT 160.950 236.700 162.750 243.600 ;
        RECT 169.650 236.700 171.450 240.600 ;
        RECT 180.300 236.700 182.100 249.600 ;
        RECT 187.800 236.700 189.600 243.600 ;
        RECT 205.800 236.700 207.600 243.600 ;
        RECT 215.400 236.700 217.200 249.600 ;
        RECT 238.800 236.700 240.600 243.600 ;
        RECT 248.400 236.700 250.200 249.600 ;
        RECT 263.400 236.700 265.200 249.600 ;
        RECT 281.400 236.700 283.200 243.600 ;
        RECT 293.400 236.700 295.200 249.600 ;
        RECT 312.300 236.700 314.100 249.600 ;
        RECT 319.800 236.700 321.600 243.600 ;
        RECT 329.400 236.700 331.200 243.600 ;
        RECT 344.400 236.700 346.200 243.600 ;
        RECT 350.400 236.700 352.200 243.600 ;
        RECT 359.550 236.700 361.350 240.600 ;
        RECT 368.250 236.700 370.050 243.600 ;
        RECT 374.850 236.700 376.650 243.600 ;
        RECT 385.050 236.700 386.850 243.600 ;
        RECT 401.400 236.700 403.200 243.600 ;
        RECT 408.900 236.700 410.700 249.600 ;
        RECT 419.400 236.700 421.200 243.600 ;
        RECT 426.900 236.700 428.700 249.600 ;
        RECT 437.400 236.700 439.200 243.600 ;
        RECT 455.400 236.700 457.200 243.600 ;
        RECT 462.900 236.700 464.700 249.600 ;
        RECT 470.400 236.700 472.200 249.600 ;
        RECT 491.400 236.700 493.200 243.600 ;
        RECT 498.900 236.700 500.700 249.600 ;
        RECT 514.800 236.700 516.600 243.600 ;
        RECT 521.550 236.700 523.350 240.600 ;
        RECT 530.250 236.700 532.050 243.600 ;
        RECT 536.850 236.700 538.650 243.600 ;
        RECT 547.050 236.700 548.850 243.600 ;
        RECT 557.400 236.700 559.200 249.600 ;
        RECT 578.400 236.700 580.200 247.800 ;
        RECT 601.800 236.700 603.600 243.600 ;
        RECT 611.400 236.700 613.200 243.600 ;
        RECT 618.900 236.700 620.700 249.600 ;
        RECT 626.400 236.700 628.200 243.600 ;
        RECT 641.400 236.700 643.200 243.600 ;
        RECT 653.400 236.700 655.200 249.600 ;
        RECT 668.400 236.700 670.200 243.600 ;
        RECT 675.000 236.700 676.800 249.600 ;
        RECT 686.400 236.700 688.200 243.600 ;
        RECT 692.400 236.700 694.200 243.600 ;
        RECT 707.400 236.700 709.200 247.800 ;
        RECT 725.400 236.700 727.200 243.600 ;
        RECT 731.400 236.700 733.200 243.600 ;
        RECT 743.400 236.700 745.200 243.600 ;
        RECT 749.400 236.700 751.200 243.600 ;
        RECT 769.800 236.700 771.600 249.600 ;
        RECT 787.800 236.700 789.600 247.800 ;
        RECT 797.550 236.700 799.350 240.600 ;
        RECT 806.250 236.700 808.050 243.600 ;
        RECT 812.850 236.700 814.650 243.600 ;
        RECT 823.050 236.700 824.850 243.600 ;
        RECT -9.450 234.300 830.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT 12.300 221.400 14.100 234.300 ;
        RECT 22.800 221.400 24.600 234.300 ;
        RECT 40.800 221.400 42.600 234.300 ;
        RECT 52.800 227.400 54.600 234.300 ;
        RECT 58.800 227.400 60.600 234.300 ;
        RECT 73.800 221.400 75.600 234.300 ;
        RECT 88.800 221.400 90.600 234.300 ;
        RECT 106.800 223.200 108.600 234.300 ;
        RECT 124.500 221.400 126.300 234.300 ;
        RECT 142.800 221.400 144.600 234.300 ;
        RECT 149.400 221.400 151.200 234.300 ;
        RECT 167.400 221.400 169.200 234.300 ;
        RECT 183.300 221.400 185.100 234.300 ;
        RECT 190.800 227.400 192.600 234.300 ;
        RECT 205.800 227.400 207.600 234.300 ;
        RECT 211.800 227.400 213.600 234.300 ;
        RECT 226.800 223.200 228.600 234.300 ;
        RECT 236.400 227.400 238.200 234.300 ;
        RECT 243.000 221.400 244.800 234.300 ;
        RECT 257.400 227.400 259.200 234.300 ;
        RECT 263.400 228.000 265.200 234.300 ;
        RECT 281.400 223.200 283.200 234.300 ;
        RECT 296.400 227.400 298.200 234.300 ;
        RECT 303.000 221.400 304.800 234.300 ;
        RECT 315.150 227.400 316.950 234.300 ;
        RECT 325.350 227.400 327.150 234.300 ;
        RECT 331.950 227.400 333.750 234.300 ;
        RECT 340.650 230.400 342.450 234.300 ;
        RECT 355.800 227.400 357.600 234.300 ;
        RECT 361.800 227.400 363.600 234.300 ;
        RECT 369.300 221.400 371.100 234.300 ;
        RECT 376.800 227.400 378.600 234.300 ;
        RECT 392.400 227.400 394.200 234.300 ;
        RECT 399.900 221.400 401.700 234.300 ;
        RECT 415.800 221.400 417.600 234.300 ;
        RECT 425.700 221.400 427.500 234.300 ;
        RECT 438.150 227.400 439.950 234.300 ;
        RECT 448.350 227.400 450.150 234.300 ;
        RECT 454.950 227.400 456.750 234.300 ;
        RECT 463.650 230.400 465.450 234.300 ;
        RECT 481.800 227.400 483.600 234.300 ;
        RECT 488.400 227.400 490.200 234.300 ;
        RECT 494.400 227.400 496.200 234.300 ;
        RECT 506.400 221.400 508.200 234.300 ;
        RECT 524.400 227.400 526.200 234.300 ;
        RECT 531.900 221.400 533.700 234.300 ;
        RECT 547.800 227.400 549.600 234.300 ;
        RECT 557.400 221.400 559.200 234.300 ;
        RECT 575.400 227.400 577.200 234.300 ;
        RECT 590.400 221.400 592.200 234.300 ;
        RECT 596.400 221.400 598.200 234.300 ;
        RECT 602.400 221.400 604.200 234.300 ;
        RECT 608.400 221.400 610.200 234.300 ;
        RECT 614.400 221.400 616.200 234.300 ;
        RECT 624.150 227.400 625.950 234.300 ;
        RECT 634.350 227.400 636.150 234.300 ;
        RECT 640.950 227.400 642.750 234.300 ;
        RECT 649.650 230.400 651.450 234.300 ;
        RECT 660.300 221.400 662.100 234.300 ;
        RECT 667.800 227.400 669.600 234.300 ;
        RECT 688.800 221.400 690.600 234.300 ;
        RECT 703.800 221.400 705.600 234.300 ;
        RECT 714.900 221.400 716.700 234.300 ;
        RECT 730.800 227.400 732.600 234.300 ;
        RECT 736.800 227.400 738.600 234.300 ;
        RECT 743.550 230.400 745.350 234.300 ;
        RECT 752.250 227.400 754.050 234.300 ;
        RECT 758.850 227.400 760.650 234.300 ;
        RECT 769.050 227.400 770.850 234.300 ;
        RECT 779.400 227.400 781.200 234.300 ;
        RECT 785.400 227.400 787.200 234.300 ;
        RECT 797.400 227.400 799.200 234.300 ;
        RECT 812.400 227.400 814.200 234.300 ;
        RECT 10.800 158.700 12.600 165.600 ;
        RECT 17.550 158.700 19.350 162.600 ;
        RECT 26.250 158.700 28.050 165.600 ;
        RECT 32.850 158.700 34.650 165.600 ;
        RECT 43.050 158.700 44.850 165.600 ;
        RECT 57.300 158.700 59.100 171.600 ;
        RECT 64.800 158.700 66.600 165.600 ;
        RECT 77.400 158.700 79.200 165.600 ;
        RECT 83.400 158.700 85.200 165.600 ;
        RECT 96.300 158.700 98.100 171.600 ;
        RECT 103.800 158.700 105.600 165.600 ;
        RECT 113.550 158.700 115.350 162.600 ;
        RECT 122.250 158.700 124.050 165.600 ;
        RECT 128.850 158.700 130.650 165.600 ;
        RECT 139.050 158.700 140.850 165.600 ;
        RECT 154.500 158.700 156.300 171.600 ;
        RECT 169.800 158.700 171.600 165.600 ;
        RECT 176.550 158.700 178.350 162.600 ;
        RECT 185.250 158.700 187.050 165.600 ;
        RECT 191.850 158.700 193.650 165.600 ;
        RECT 202.050 158.700 203.850 165.600 ;
        RECT 213.300 158.700 215.100 171.600 ;
        RECT 220.800 158.700 222.600 165.600 ;
        RECT 235.800 158.700 237.600 171.600 ;
        RECT 241.800 158.700 243.600 171.600 ;
        RECT 247.800 158.700 249.600 171.600 ;
        RECT 253.800 158.700 255.600 171.600 ;
        RECT 259.800 158.700 261.600 171.600 ;
        RECT 270.300 158.700 272.100 171.600 ;
        RECT 277.800 158.700 279.600 165.600 ;
        RECT 295.200 158.700 297.000 171.600 ;
        RECT 301.800 158.700 303.600 165.600 ;
        RECT 311.400 158.700 313.200 171.600 ;
        RECT 327.300 158.700 329.100 171.600 ;
        RECT 334.800 158.700 336.600 165.600 ;
        RECT 347.400 158.700 349.200 165.600 ;
        RECT 359.550 158.700 361.350 162.600 ;
        RECT 368.250 158.700 370.050 165.600 ;
        RECT 374.850 158.700 376.650 165.600 ;
        RECT 385.050 158.700 386.850 165.600 ;
        RECT 403.800 158.700 405.600 171.600 ;
        RECT 421.800 158.700 423.600 169.800 ;
        RECT 433.800 158.700 435.600 171.600 ;
        RECT 439.800 158.700 441.600 171.600 ;
        RECT 445.800 158.700 447.600 171.600 ;
        RECT 451.800 158.700 453.600 171.600 ;
        RECT 457.800 158.700 459.600 171.600 ;
        RECT 467.400 158.700 469.200 171.600 ;
        RECT 473.400 158.700 475.200 171.600 ;
        RECT 479.400 158.700 481.200 171.600 ;
        RECT 485.400 158.700 487.200 171.600 ;
        RECT 491.400 158.700 493.200 171.600 ;
        RECT 505.800 158.700 507.600 165.600 ;
        RECT 511.800 158.700 513.600 165.600 ;
        RECT 524.400 158.700 526.200 165.600 ;
        RECT 531.900 158.700 533.700 171.600 ;
        RECT 539.550 158.700 541.350 162.600 ;
        RECT 548.250 158.700 550.050 165.600 ;
        RECT 554.850 158.700 556.650 165.600 ;
        RECT 565.050 158.700 566.850 165.600 ;
        RECT 581.400 158.700 583.200 165.600 ;
        RECT 588.900 158.700 590.700 171.600 ;
        RECT 604.200 158.700 606.000 171.600 ;
        RECT 610.800 158.700 612.600 165.600 ;
        RECT 618.300 158.700 620.100 171.600 ;
        RECT 625.800 158.700 627.600 165.600 ;
        RECT 638.700 158.700 640.500 171.600 ;
        RECT 650.400 158.700 652.200 165.600 ;
        RECT 665.400 158.700 667.200 165.600 ;
        RECT 680.400 158.700 682.200 165.600 ;
        RECT 687.900 158.700 689.700 171.600 ;
        RECT 698.400 158.700 700.200 171.600 ;
        RECT 716.400 158.700 718.200 171.600 ;
        RECT 734.400 158.700 736.200 165.600 ;
        RECT 751.800 158.700 753.600 165.600 ;
        RECT 762.300 158.700 764.100 171.600 ;
        RECT 769.800 158.700 771.600 165.600 ;
        RECT 781.800 158.700 783.600 165.600 ;
        RECT 787.800 158.700 789.600 165.600 ;
        RECT 795.150 158.700 796.950 165.600 ;
        RECT 805.350 158.700 807.150 165.600 ;
        RECT 811.950 158.700 813.750 165.600 ;
        RECT 820.650 158.700 822.450 162.600 ;
        RECT -9.450 156.300 830.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT 6.150 149.400 7.950 156.300 ;
        RECT 16.350 149.400 18.150 156.300 ;
        RECT 22.950 149.400 24.750 156.300 ;
        RECT 31.650 152.400 33.450 156.300 ;
        RECT 49.800 143.400 51.600 156.300 ;
        RECT 56.400 149.400 58.200 156.300 ;
        RECT 69.300 143.400 71.100 156.300 ;
        RECT 76.800 149.400 78.600 156.300 ;
        RECT 97.800 143.400 99.600 156.300 ;
        RECT 108.300 143.400 110.100 156.300 ;
        RECT 115.800 149.400 117.600 156.300 ;
        RECT 127.800 149.400 129.600 156.300 ;
        RECT 133.800 149.400 135.600 156.300 ;
        RECT 148.800 143.400 150.600 156.300 ;
        RECT 157.800 149.400 159.600 156.300 ;
        RECT 163.800 149.400 165.600 156.300 ;
        RECT 178.800 149.400 180.600 156.300 ;
        RECT 189.300 143.400 191.100 156.300 ;
        RECT 196.800 149.400 198.600 156.300 ;
        RECT 212.400 149.400 214.200 156.300 ;
        RECT 219.900 143.400 221.700 156.300 ;
        RECT 235.800 149.400 237.600 156.300 ;
        RECT 242.400 149.400 244.200 156.300 ;
        RECT 248.400 149.400 250.200 156.300 ;
        RECT 257.400 149.400 259.200 156.300 ;
        RECT 263.400 149.400 265.200 156.300 ;
        RECT 275.400 149.400 277.200 156.300 ;
        RECT 281.400 149.400 283.200 156.300 ;
        RECT 297.900 143.400 299.700 156.300 ;
        RECT 322.800 145.200 324.600 156.300 ;
        RECT 332.400 149.400 334.200 156.300 ;
        RECT 338.400 149.400 340.200 156.300 ;
        RECT 350.400 149.400 352.200 156.300 ;
        RECT 356.400 149.400 358.200 156.300 ;
        RECT 369.300 143.400 371.100 156.300 ;
        RECT 376.800 149.400 378.600 156.300 ;
        RECT 388.800 149.400 390.600 156.300 ;
        RECT 394.800 149.400 396.600 156.300 ;
        RECT 402.150 149.400 403.950 156.300 ;
        RECT 412.350 149.400 414.150 156.300 ;
        RECT 418.950 149.400 420.750 156.300 ;
        RECT 427.650 152.400 429.450 156.300 ;
        RECT 443.400 145.500 445.200 156.300 ;
        RECT 467.700 143.400 469.500 156.300 ;
        RECT 482.400 149.400 484.200 156.300 ;
        RECT 489.900 143.400 491.700 156.300 ;
        RECT 497.550 152.400 499.350 156.300 ;
        RECT 506.250 149.400 508.050 156.300 ;
        RECT 512.850 149.400 514.650 156.300 ;
        RECT 523.050 149.400 524.850 156.300 ;
        RECT 533.400 143.400 535.200 156.300 ;
        RECT 548.550 152.400 550.350 156.300 ;
        RECT 557.250 149.400 559.050 156.300 ;
        RECT 563.850 149.400 565.650 156.300 ;
        RECT 574.050 149.400 575.850 156.300 ;
        RECT 592.800 145.200 594.600 156.300 ;
        RECT 612.300 143.400 614.100 156.300 ;
        RECT 626.400 149.400 628.200 156.300 ;
        RECT 641.400 149.400 643.200 156.300 ;
        RECT 647.400 149.400 649.200 156.300 ;
        RECT 656.550 152.400 658.350 156.300 ;
        RECT 665.250 149.400 667.050 156.300 ;
        RECT 671.850 149.400 673.650 156.300 ;
        RECT 682.050 149.400 683.850 156.300 ;
        RECT 692.400 149.400 694.200 156.300 ;
        RECT 698.400 149.400 700.200 156.300 ;
        RECT 713.400 149.400 715.200 156.300 ;
        RECT 720.900 143.400 722.700 156.300 ;
        RECT 731.400 149.400 733.200 156.300 ;
        RECT 738.900 143.400 740.700 156.300 ;
        RECT 752.400 145.200 754.200 156.300 ;
        RECT 770.400 149.400 772.200 156.300 ;
        RECT 777.900 143.400 779.700 156.300 ;
        RECT 785.400 143.400 787.200 156.300 ;
        RECT 803.400 149.400 805.200 156.300 ;
        RECT 815.400 149.400 817.200 156.300 ;
        RECT 821.400 149.400 823.200 156.300 ;
        RECT 16.800 80.700 18.600 93.600 ;
        RECT 26.400 80.700 28.200 93.600 ;
        RECT 49.800 80.700 51.600 91.800 ;
        RECT 66.900 80.700 68.700 93.600 ;
        RECT 80.400 80.700 82.200 87.600 ;
        RECT 86.400 80.700 88.200 87.600 ;
        RECT 95.400 80.700 97.200 87.600 ;
        RECT 101.400 80.700 103.200 87.600 ;
        RECT 110.400 80.700 112.200 87.600 ;
        RECT 116.400 80.700 118.200 87.600 ;
        RECT 131.400 80.700 133.200 87.600 ;
        RECT 138.900 80.700 140.700 93.600 ;
        RECT 149.400 80.700 151.200 87.600 ;
        RECT 166.800 80.700 168.600 87.600 ;
        RECT 172.800 80.700 174.600 87.600 ;
        RECT 179.550 80.700 181.350 84.600 ;
        RECT 188.250 80.700 190.050 87.600 ;
        RECT 194.850 80.700 196.650 87.600 ;
        RECT 205.050 80.700 206.850 87.600 ;
        RECT 215.400 80.700 217.200 87.600 ;
        RECT 222.000 80.700 223.800 93.600 ;
        RECT 234.300 80.700 236.100 93.600 ;
        RECT 241.800 80.700 243.600 87.600 ;
        RECT 251.400 80.700 253.200 87.600 ;
        RECT 257.400 80.700 259.200 87.600 ;
        RECT 271.500 80.700 273.300 93.600 ;
        RECT 289.200 80.700 291.000 93.600 ;
        RECT 295.800 80.700 297.600 87.600 ;
        RECT 302.400 80.700 304.200 93.600 ;
        RECT 321.300 80.700 323.100 93.600 ;
        RECT 328.800 80.700 330.600 87.600 ;
        RECT 346.500 80.700 348.300 93.600 ;
        RECT 360.300 80.700 362.100 93.600 ;
        RECT 367.800 80.700 369.600 87.600 ;
        RECT 378.150 80.700 379.950 87.600 ;
        RECT 388.350 80.700 390.150 87.600 ;
        RECT 394.950 80.700 396.750 87.600 ;
        RECT 403.650 80.700 405.450 84.600 ;
        RECT 413.400 80.700 415.200 87.600 ;
        RECT 419.400 80.700 421.200 87.600 ;
        RECT 429.150 80.700 430.950 87.600 ;
        RECT 439.350 80.700 441.150 87.600 ;
        RECT 445.950 80.700 447.750 87.600 ;
        RECT 454.650 80.700 456.450 84.600 ;
        RECT 475.800 80.700 477.600 93.600 ;
        RECT 485.400 80.700 487.200 87.600 ;
        RECT 492.900 80.700 494.700 93.600 ;
        RECT 500.400 80.700 502.200 87.600 ;
        RECT 506.400 80.700 508.200 87.000 ;
        RECT 518.550 80.700 520.350 84.600 ;
        RECT 527.250 80.700 529.050 87.600 ;
        RECT 533.850 80.700 535.650 87.600 ;
        RECT 544.050 80.700 545.850 87.600 ;
        RECT 557.400 80.700 559.200 87.600 ;
        RECT 563.400 80.700 565.200 87.600 ;
        RECT 578.400 80.700 580.200 91.500 ;
        RECT 597.300 80.700 599.100 93.600 ;
        RECT 604.800 80.700 606.600 87.600 ;
        RECT 617.400 80.700 619.200 87.600 ;
        RECT 623.400 80.700 625.200 87.600 ;
        RECT 636.300 80.700 638.100 93.600 ;
        RECT 643.800 80.700 645.600 87.600 ;
        RECT 656.700 80.700 658.500 93.600 ;
        RECT 668.550 80.700 670.350 84.600 ;
        RECT 677.250 80.700 679.050 87.600 ;
        RECT 683.850 80.700 685.650 87.600 ;
        RECT 694.050 80.700 695.850 87.600 ;
        RECT 707.400 80.700 709.200 91.500 ;
        RECT 736.800 80.700 738.600 91.800 ;
        RECT 750.900 80.700 752.700 93.600 ;
        RECT 764.550 80.700 766.350 84.600 ;
        RECT 773.250 80.700 775.050 87.600 ;
        RECT 779.850 80.700 781.650 87.600 ;
        RECT 790.050 80.700 791.850 87.600 ;
        RECT 804.300 80.700 806.100 93.600 ;
        RECT 811.800 80.700 813.600 87.600 ;
        RECT -9.450 78.300 830.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT 6.150 71.400 7.950 78.300 ;
        RECT 16.350 71.400 18.150 78.300 ;
        RECT 22.950 71.400 24.750 78.300 ;
        RECT 31.650 74.400 33.450 78.300 ;
        RECT 41.550 74.400 43.350 78.300 ;
        RECT 50.250 71.400 52.050 78.300 ;
        RECT 56.850 71.400 58.650 78.300 ;
        RECT 67.050 71.400 68.850 78.300 ;
        RECT 81.300 65.400 83.100 78.300 ;
        RECT 88.800 71.400 90.600 78.300 ;
        RECT 99.150 71.400 100.950 78.300 ;
        RECT 109.350 71.400 111.150 78.300 ;
        RECT 115.950 71.400 117.750 78.300 ;
        RECT 124.650 74.400 126.450 78.300 ;
        RECT 137.400 71.400 139.200 78.300 ;
        RECT 143.400 71.400 145.200 78.300 ;
        RECT 153.300 65.400 155.100 78.300 ;
        RECT 160.800 71.400 162.600 78.300 ;
        RECT 171.150 71.400 172.950 78.300 ;
        RECT 181.350 71.400 183.150 78.300 ;
        RECT 187.950 71.400 189.750 78.300 ;
        RECT 196.650 74.400 198.450 78.300 ;
        RECT 209.400 71.400 211.200 78.300 ;
        RECT 215.400 71.400 217.200 78.300 ;
        RECT 225.150 71.400 226.950 78.300 ;
        RECT 235.350 71.400 237.150 78.300 ;
        RECT 241.950 71.400 243.750 78.300 ;
        RECT 250.650 74.400 252.450 78.300 ;
        RECT 260.400 71.400 262.200 78.300 ;
        RECT 266.400 71.400 268.200 78.300 ;
        RECT 278.400 71.400 280.200 78.300 ;
        RECT 285.900 65.400 287.700 78.300 ;
        RECT 296.400 71.400 298.200 78.300 ;
        RECT 302.400 71.400 304.200 78.300 ;
        RECT 314.400 67.500 316.200 78.300 ;
        RECT 338.400 71.400 340.200 78.300 ;
        RECT 345.900 65.400 347.700 78.300 ;
        RECT 358.800 71.400 360.600 78.300 ;
        RECT 366.150 71.400 367.950 78.300 ;
        RECT 376.350 71.400 378.150 78.300 ;
        RECT 382.950 71.400 384.750 78.300 ;
        RECT 391.650 74.400 393.450 78.300 ;
        RECT 412.800 67.500 414.600 78.300 ;
        RECT 430.500 65.400 432.300 78.300 ;
        RECT 443.400 65.400 445.200 78.300 ;
        RECT 461.400 71.400 463.200 78.300 ;
        RECT 477.300 65.400 479.100 78.300 ;
        RECT 484.800 71.400 486.600 78.300 ;
        RECT 500.400 71.400 502.200 78.300 ;
        RECT 507.900 65.400 509.700 78.300 ;
        RECT 523.800 71.400 525.600 78.300 ;
        RECT 531.150 71.400 532.950 78.300 ;
        RECT 541.350 71.400 543.150 78.300 ;
        RECT 547.950 71.400 549.750 78.300 ;
        RECT 556.650 74.400 558.450 78.300 ;
        RECT 569.400 71.400 571.200 78.300 ;
        RECT 582.150 71.400 583.950 78.300 ;
        RECT 592.350 71.400 594.150 78.300 ;
        RECT 598.950 71.400 600.750 78.300 ;
        RECT 607.650 74.400 609.450 78.300 ;
        RECT 623.400 71.400 625.200 78.300 ;
        RECT 630.900 65.400 632.700 78.300 ;
        RECT 640.800 65.400 642.600 78.300 ;
        RECT 646.800 65.400 648.600 78.300 ;
        RECT 652.800 65.400 654.600 78.300 ;
        RECT 665.700 65.400 667.500 78.300 ;
        RECT 682.800 71.400 684.600 78.300 ;
        RECT 688.800 71.400 690.600 78.300 ;
        RECT 698.400 71.400 700.200 78.300 ;
        RECT 716.400 71.400 718.200 78.300 ;
        RECT 723.900 65.400 725.700 78.300 ;
        RECT 731.400 71.400 733.200 78.300 ;
        RECT 737.400 71.400 739.200 78.300 ;
        RECT 750.300 65.400 752.100 78.300 ;
        RECT 757.800 71.400 759.600 78.300 ;
        RECT 773.400 71.400 775.200 78.300 ;
        RECT 780.900 65.400 782.700 78.300 ;
        RECT 788.400 71.400 790.200 78.300 ;
        RECT 803.400 71.400 805.200 78.300 ;
        RECT 818.700 65.400 820.500 78.300 ;
        RECT 10.800 2.700 12.600 9.600 ;
        RECT 28.800 2.700 30.600 15.600 ;
        RECT 43.800 2.700 45.600 9.600 ;
        RECT 58.800 2.700 60.600 15.600 ;
        RECT 69.300 2.700 71.100 15.600 ;
        RECT 76.800 2.700 78.600 9.600 ;
        RECT 89.400 2.700 91.200 9.600 ;
        RECT 109.800 2.700 111.600 9.600 ;
        RECT 117.300 2.700 119.100 15.600 ;
        RECT 124.800 2.700 126.600 9.600 ;
        RECT 134.400 2.700 136.200 9.600 ;
        RECT 146.400 2.700 148.200 9.600 ;
        RECT 152.400 2.700 154.200 9.000 ;
        RECT 169.800 2.700 171.600 9.600 ;
        RECT 175.800 2.700 177.600 9.600 ;
        RECT 182.400 2.700 184.200 9.600 ;
        RECT 188.400 2.700 190.200 9.600 ;
        RECT 201.300 2.700 203.100 15.600 ;
        RECT 208.800 2.700 210.600 9.600 ;
        RECT 219.150 2.700 220.950 9.600 ;
        RECT 229.350 2.700 231.150 9.600 ;
        RECT 235.950 2.700 237.750 9.600 ;
        RECT 244.650 2.700 246.450 6.600 ;
        RECT 255.150 2.700 256.950 9.600 ;
        RECT 265.350 2.700 267.150 9.600 ;
        RECT 271.950 2.700 273.750 9.600 ;
        RECT 280.650 2.700 282.450 6.600 ;
        RECT 301.800 2.700 303.600 13.500 ;
        RECT 322.800 2.700 324.600 15.600 ;
        RECT 329.550 2.700 331.350 6.600 ;
        RECT 338.250 2.700 340.050 9.600 ;
        RECT 344.850 2.700 346.650 9.600 ;
        RECT 355.050 2.700 356.850 9.600 ;
        RECT 373.800 2.700 375.600 13.800 ;
        RECT 384.150 2.700 385.950 9.600 ;
        RECT 394.350 2.700 396.150 9.600 ;
        RECT 400.950 2.700 402.750 9.600 ;
        RECT 409.650 2.700 411.450 6.600 ;
        RECT 427.500 2.700 429.300 15.600 ;
        RECT 443.400 2.700 445.200 9.600 ;
        RECT 450.900 2.700 452.700 15.600 ;
        RECT 463.500 2.700 465.300 15.600 ;
        RECT 479.400 2.700 481.200 9.600 ;
        RECT 486.900 2.700 488.700 15.600 ;
        RECT 500.700 2.700 502.500 15.600 ;
        RECT 515.700 2.700 517.500 15.600 ;
        RECT 532.800 2.700 534.600 9.600 ;
        RECT 539.400 2.700 541.200 15.600 ;
        RECT 560.400 2.700 562.200 9.600 ;
        RECT 567.900 2.700 569.700 15.600 ;
        RECT 575.400 2.700 577.200 9.600 ;
        RECT 581.400 2.700 583.200 9.600 ;
        RECT 590.550 2.700 592.350 6.600 ;
        RECT 599.250 2.700 601.050 9.600 ;
        RECT 605.850 2.700 607.650 9.600 ;
        RECT 616.050 2.700 617.850 9.600 ;
        RECT 629.400 2.700 631.200 9.600 ;
        RECT 635.400 2.700 637.200 9.600 ;
        RECT 649.800 2.700 651.600 9.600 ;
        RECT 655.800 2.700 657.600 9.600 ;
        RECT 662.550 2.700 664.350 6.600 ;
        RECT 671.250 2.700 673.050 9.600 ;
        RECT 677.850 2.700 679.650 9.600 ;
        RECT 688.050 2.700 689.850 9.600 ;
        RECT 701.400 2.700 703.200 9.600 ;
        RECT 708.900 2.700 710.700 15.600 ;
        RECT 727.800 2.700 729.600 15.600 ;
        RECT 739.800 2.700 741.600 9.000 ;
        RECT 745.800 2.700 747.600 9.600 ;
        RECT 752.550 2.700 754.350 6.600 ;
        RECT 761.250 2.700 763.050 9.600 ;
        RECT 767.850 2.700 769.650 9.600 ;
        RECT 778.050 2.700 779.850 9.600 ;
        RECT 791.700 2.700 793.500 15.600 ;
        RECT 806.400 2.700 808.200 9.600 ;
        RECT 812.400 2.700 814.200 9.600 ;
        RECT -9.450 0.300 830.400 2.700 ;
    END
  END vdd
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 352.950 642.450 355.050 643.050 ;
        RECT 361.950 642.450 364.050 643.050 ;
        RECT 352.950 641.550 364.050 642.450 ;
        RECT 352.950 640.950 355.050 641.550 ;
        RECT 361.950 640.950 364.050 641.550 ;
        RECT 376.950 640.950 379.050 643.050 ;
        RECT 367.950 607.950 370.050 610.050 ;
        RECT 595.950 607.950 598.050 610.050 ;
        RECT 586.950 604.950 589.050 607.050 ;
      LAYER metal2 ;
        RECT 377.400 827.400 381.450 828.450 ;
        RECT 377.400 789.450 378.450 827.400 ;
        RECT 377.400 788.400 381.450 789.450 ;
        RECT 380.400 745.050 381.450 788.400 ;
        RECT 355.950 742.950 358.050 745.050 ;
        RECT 379.950 742.950 382.050 745.050 ;
        RECT 356.400 703.050 357.450 742.950 ;
        RECT 355.950 700.950 358.050 703.050 ;
        RECT 382.950 700.950 385.050 703.050 ;
        RECT 383.400 693.450 384.450 700.950 ;
        RECT 380.400 692.400 384.450 693.450 ;
        RECT 380.400 684.450 381.450 692.400 ;
        RECT 377.400 683.400 381.450 684.450 ;
        RECT 377.400 646.050 378.450 683.400 ;
        RECT 361.950 640.950 364.050 646.050 ;
        RECT 376.950 640.950 379.050 646.050 ;
        RECT 362.400 616.050 363.450 640.950 ;
        RECT 586.950 631.950 589.050 634.050 ;
        RECT 503.100 628.950 505.200 631.050 ;
        RECT 503.400 625.050 504.450 628.950 ;
        RECT 430.950 622.950 433.050 625.050 ;
        RECT 502.950 622.950 505.050 625.050 ;
        RECT 431.400 616.050 432.450 622.950 ;
        RECT 361.950 613.950 364.050 616.050 ;
        RECT 367.950 613.950 370.050 616.050 ;
        RECT 430.950 613.950 433.050 616.050 ;
        RECT 368.400 610.050 369.450 613.950 ;
        RECT 587.400 610.050 588.450 631.950 ;
        RECT 367.950 607.950 370.050 610.050 ;
        RECT 586.950 604.950 589.050 610.050 ;
        RECT 592.950 607.950 598.050 610.050 ;
      LAYER metal3 ;
        RECT 355.950 744.600 358.050 745.050 ;
        RECT 379.950 744.600 382.050 745.050 ;
        RECT 355.950 743.400 382.050 744.600 ;
        RECT 355.950 742.950 358.050 743.400 ;
        RECT 379.950 742.950 382.050 743.400 ;
        RECT 355.950 702.600 358.050 703.050 ;
        RECT 382.950 702.600 385.050 703.050 ;
        RECT 355.950 701.400 385.050 702.600 ;
        RECT 355.950 700.950 358.050 701.400 ;
        RECT 382.950 700.950 385.050 701.400 ;
        RECT 361.950 645.600 364.050 646.050 ;
        RECT 376.950 645.600 379.050 646.050 ;
        RECT 361.950 644.400 379.050 645.600 ;
        RECT 361.950 643.950 364.050 644.400 ;
        RECT 376.950 643.950 379.050 644.400 ;
        RECT 586.950 633.600 589.050 634.050 ;
        RECT 578.400 632.400 589.050 633.600 ;
        RECT 503.100 630.600 505.200 631.050 ;
        RECT 578.400 630.600 579.600 632.400 ;
        RECT 586.950 631.950 589.050 632.400 ;
        RECT 503.100 629.400 579.600 630.600 ;
        RECT 503.100 628.950 505.200 629.400 ;
        RECT 430.950 624.600 433.050 625.050 ;
        RECT 502.950 624.600 505.050 625.050 ;
        RECT 430.950 623.400 505.050 624.600 ;
        RECT 430.950 622.950 433.050 623.400 ;
        RECT 502.950 622.950 505.050 623.400 ;
        RECT 361.950 615.600 364.050 616.050 ;
        RECT 367.950 615.600 370.050 616.050 ;
        RECT 430.950 615.600 433.050 616.050 ;
        RECT 361.950 614.400 433.050 615.600 ;
        RECT 361.950 613.950 364.050 614.400 ;
        RECT 367.950 613.950 370.050 614.400 ;
        RECT 430.950 613.950 433.050 614.400 ;
        RECT 586.950 609.600 589.050 610.050 ;
        RECT 592.950 609.600 595.050 610.050 ;
        RECT 586.950 608.400 595.050 609.600 ;
        RECT 586.950 607.950 589.050 608.400 ;
        RECT 592.950 607.950 595.050 608.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 475.950 645.450 478.050 646.200 ;
        RECT 484.950 645.450 487.050 646.050 ;
        RECT 475.950 644.550 487.050 645.450 ;
        RECT 475.950 643.950 478.050 644.550 ;
        RECT 484.950 643.950 487.050 644.550 ;
        RECT 265.950 637.950 268.050 643.050 ;
        RECT 313.950 604.950 316.050 607.050 ;
        RECT 565.950 604.950 568.050 607.050 ;
        RECT 262.950 565.950 265.050 568.200 ;
        RECT 307.950 565.950 310.050 568.050 ;
        RECT 385.950 565.950 388.050 568.050 ;
        RECT 232.950 562.950 235.050 565.050 ;
        RECT 418.950 562.950 421.050 565.050 ;
        RECT 544.950 529.950 547.050 532.050 ;
        RECT 613.950 529.950 616.050 532.050 ;
      LAYER metal2 ;
        RECT 467.400 804.450 468.450 828.450 ;
        RECT 464.400 803.400 468.450 804.450 ;
        RECT 464.400 784.050 465.450 803.400 ;
        RECT 463.950 781.950 466.050 784.050 ;
        RECT 481.950 781.800 484.050 783.900 ;
        RECT 482.400 732.450 483.450 781.800 ;
        RECT 479.400 731.400 483.450 732.450 ;
        RECT 479.400 682.050 480.450 731.400 ;
        RECT 478.950 679.950 481.050 682.050 ;
        RECT 484.950 679.800 487.050 681.900 ;
        RECT 475.950 646.050 478.050 646.200 ;
        RECT 485.400 646.050 486.450 679.800 ;
        RECT 475.950 645.600 480.000 646.050 ;
        RECT 475.950 644.100 480.450 645.600 ;
        RECT 477.000 643.950 480.450 644.100 ;
        RECT 484.950 643.950 487.050 646.050 ;
        RECT 265.950 637.950 268.050 640.050 ;
        RECT 266.400 625.050 267.450 637.950 ;
        RECT 265.950 622.950 268.050 625.050 ;
        RECT 307.950 622.950 310.050 625.050 ;
        RECT 313.950 622.950 316.050 625.050 ;
        RECT 266.400 580.050 267.450 622.950 ;
        RECT 232.950 577.950 235.050 580.050 ;
        RECT 265.950 577.950 268.050 580.050 ;
        RECT 233.400 571.050 234.450 577.950 ;
        RECT 232.950 568.950 235.050 571.050 ;
        RECT 233.400 565.050 234.450 568.950 ;
        RECT 262.950 566.100 265.050 571.050 ;
        RECT 308.400 568.050 309.450 622.950 ;
        RECT 314.400 619.050 315.450 622.950 ;
        RECT 479.400 619.050 480.450 643.950 ;
        RECT 313.950 616.950 316.050 619.050 ;
        RECT 478.950 616.950 481.050 619.050 ;
        RECT 541.950 616.950 544.050 619.050 ;
        RECT 314.400 607.050 315.450 616.950 ;
        RECT 313.950 604.950 316.050 607.050 ;
        RECT 542.400 604.050 543.450 616.950 ;
        RECT 541.950 601.950 544.050 604.050 ;
        RECT 565.950 601.950 568.050 607.050 ;
        RECT 542.400 570.450 543.450 601.950 ;
        RECT 542.400 569.400 546.450 570.450 ;
        RECT 307.950 565.950 310.050 568.050 ;
        RECT 385.950 565.950 388.050 568.050 ;
        RECT 232.950 562.950 235.050 565.050 ;
        RECT 308.400 559.050 309.450 565.950 ;
        RECT 307.950 556.950 310.050 559.050 ;
        RECT 346.800 556.950 348.900 559.050 ;
        RECT 347.400 541.050 348.450 556.950 ;
        RECT 386.400 553.050 387.450 565.950 ;
        RECT 418.950 562.950 421.050 565.050 ;
        RECT 419.400 553.050 420.450 562.950 ;
        RECT 385.950 550.950 388.050 553.050 ;
        RECT 418.950 550.950 421.050 553.050 ;
        RECT 386.400 541.050 387.450 550.950 ;
        RECT 346.950 538.950 349.050 541.050 ;
        RECT 385.950 538.950 388.050 541.050 ;
        RECT 545.400 532.050 546.450 569.400 ;
        RECT 544.950 529.950 547.050 532.050 ;
        RECT 610.950 529.950 616.050 532.050 ;
      LAYER metal3 ;
        RECT 463.950 783.600 466.050 784.050 ;
        RECT 481.950 783.600 484.050 783.900 ;
        RECT 463.950 782.400 484.050 783.600 ;
        RECT 463.950 781.950 466.050 782.400 ;
        RECT 481.950 781.800 484.050 782.400 ;
        RECT 478.950 681.600 481.050 682.050 ;
        RECT 484.950 681.600 487.050 681.900 ;
        RECT 478.950 680.400 487.050 681.600 ;
        RECT 478.950 679.950 481.050 680.400 ;
        RECT 484.950 679.800 487.050 680.400 ;
        RECT 265.950 624.600 268.050 625.050 ;
        RECT 307.950 624.600 310.050 625.050 ;
        RECT 313.950 624.600 316.050 625.050 ;
        RECT 265.950 623.400 316.050 624.600 ;
        RECT 265.950 622.950 268.050 623.400 ;
        RECT 307.950 622.950 310.050 623.400 ;
        RECT 313.950 622.950 316.050 623.400 ;
        RECT 313.950 618.600 316.050 619.050 ;
        RECT 478.950 618.600 481.050 619.050 ;
        RECT 541.950 618.600 544.050 619.050 ;
        RECT 313.950 617.400 544.050 618.600 ;
        RECT 313.950 616.950 316.050 617.400 ;
        RECT 478.950 616.950 481.050 617.400 ;
        RECT 541.950 616.950 544.050 617.400 ;
        RECT 541.950 603.600 544.050 604.050 ;
        RECT 565.950 603.600 568.050 604.050 ;
        RECT 541.950 602.400 568.050 603.600 ;
        RECT 541.950 601.950 544.050 602.400 ;
        RECT 565.950 601.950 568.050 602.400 ;
        RECT 232.950 579.600 235.050 580.050 ;
        RECT 265.950 579.600 268.050 580.050 ;
        RECT 232.950 578.400 268.050 579.600 ;
        RECT 232.950 577.950 235.050 578.400 ;
        RECT 265.950 577.950 268.050 578.400 ;
        RECT 232.950 570.600 235.050 571.050 ;
        RECT 262.950 570.600 265.050 571.050 ;
        RECT 232.950 569.400 265.050 570.600 ;
        RECT 232.950 568.950 235.050 569.400 ;
        RECT 262.950 568.950 265.050 569.400 ;
        RECT 307.950 558.600 310.050 559.050 ;
        RECT 346.800 558.600 348.900 559.050 ;
        RECT 307.950 557.400 348.900 558.600 ;
        RECT 307.950 556.950 310.050 557.400 ;
        RECT 346.800 556.950 348.900 557.400 ;
        RECT 385.950 552.600 388.050 553.050 ;
        RECT 418.950 552.600 421.050 553.050 ;
        RECT 385.950 551.400 421.050 552.600 ;
        RECT 385.950 550.950 388.050 551.400 ;
        RECT 418.950 550.950 421.050 551.400 ;
        RECT 346.950 540.600 349.050 541.050 ;
        RECT 385.950 540.600 388.050 541.050 ;
        RECT 346.950 539.400 388.050 540.600 ;
        RECT 346.950 538.950 349.050 539.400 ;
        RECT 385.950 538.950 388.050 539.400 ;
        RECT 544.950 531.600 547.050 532.050 ;
        RECT 610.950 531.600 613.050 532.050 ;
        RECT 544.950 530.400 613.050 531.600 ;
        RECT 544.950 529.950 547.050 530.400 ;
        RECT 610.950 529.950 613.050 530.400 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 469.950 643.950 472.050 646.050 ;
        RECT 274.950 607.950 277.050 610.050 ;
        RECT 403.950 604.950 406.050 610.050 ;
        RECT 493.950 607.950 496.050 610.050 ;
        RECT 547.950 607.950 550.050 610.050 ;
        RECT 475.950 604.950 478.050 607.050 ;
        RECT 175.950 565.800 178.050 568.050 ;
        RECT 274.950 565.950 277.050 568.050 ;
        RECT 472.950 562.950 475.050 565.050 ;
        RECT 562.950 526.950 565.050 529.050 ;
        RECT 223.950 484.950 226.050 487.050 ;
      LAYER metal2 ;
        RECT 482.400 787.200 483.450 828.450 ;
        RECT 460.950 784.950 463.050 787.050 ;
        RECT 481.950 785.100 484.050 787.200 ;
        RECT 461.400 736.050 462.450 784.950 ;
        RECT 454.950 733.950 457.050 736.050 ;
        RECT 460.950 733.950 463.050 736.050 ;
        RECT 455.400 715.050 456.450 733.950 ;
        RECT 439.950 712.950 442.050 715.050 ;
        RECT 454.950 712.950 457.050 715.050 ;
        RECT 440.400 664.050 441.450 712.950 ;
        RECT 427.950 661.950 430.050 664.050 ;
        RECT 439.950 661.950 442.050 664.050 ;
        RECT 428.400 643.050 429.450 661.950 ;
        RECT 427.950 640.950 430.050 643.050 ;
        RECT 469.950 640.950 472.050 646.050 ;
        RECT 428.400 637.050 429.450 640.950 ;
        RECT 475.950 640.800 478.050 642.900 ;
        RECT 403.950 634.950 406.050 637.050 ;
        RECT 427.950 634.950 430.050 637.050 ;
        RECT 404.400 610.050 405.450 634.950 ;
        RECT 274.950 607.950 277.050 610.050 ;
        RECT 403.950 607.950 406.050 610.050 ;
        RECT 275.400 571.050 276.450 607.950 ;
        RECT 404.400 580.050 405.450 607.950 ;
        RECT 476.400 607.050 477.450 640.800 ;
        RECT 475.950 604.950 478.050 607.050 ;
        RECT 493.950 604.950 496.050 610.050 ;
        RECT 547.950 607.950 550.050 610.050 ;
        RECT 494.400 595.050 495.450 604.950 ;
        RECT 493.950 592.950 496.050 595.050 ;
        RECT 373.950 577.950 376.050 580.050 ;
        RECT 403.950 577.950 406.050 580.050 ;
        RECT 175.950 565.800 178.050 567.900 ;
        RECT 274.950 565.950 277.050 571.050 ;
        RECT 286.950 568.950 289.050 571.050 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 176.400 550.050 177.450 565.800 ;
        RECT 175.950 547.950 178.050 550.050 ;
        RECT 190.800 547.950 192.900 550.050 ;
        RECT 191.400 526.200 192.450 547.950 ;
        RECT 190.950 524.100 193.050 526.200 ;
        RECT 287.400 523.050 288.450 568.950 ;
        RECT 311.400 553.050 312.450 568.950 ;
        RECT 374.400 553.050 375.450 577.950 ;
        RECT 494.400 577.050 495.450 592.950 ;
        RECT 548.400 592.050 549.450 607.950 ;
        RECT 547.950 589.950 550.050 592.050 ;
        RECT 472.950 574.950 475.050 577.050 ;
        RECT 493.950 574.950 496.050 577.050 ;
        RECT 473.400 565.050 474.450 574.950 ;
        RECT 472.950 562.950 475.050 565.050 ;
        RECT 310.950 550.950 313.050 553.050 ;
        RECT 373.950 550.950 376.050 553.050 ;
        RECT 548.400 544.050 549.450 589.950 ;
        RECT 547.950 541.950 550.050 544.050 ;
        RECT 562.950 541.950 565.050 544.050 ;
        RECT 563.400 529.050 564.450 541.950 ;
        RECT 562.950 526.950 565.050 529.050 ;
        RECT 205.950 520.950 208.050 523.050 ;
        RECT 226.950 520.950 229.050 523.050 ;
        RECT 286.950 520.950 289.050 523.050 ;
        RECT 206.400 517.050 207.450 520.950 ;
        RECT 227.400 517.050 228.450 520.950 ;
        RECT 205.950 514.950 208.050 517.050 ;
        RECT 226.950 514.950 229.050 517.050 ;
        RECT 227.400 498.450 228.450 514.950 ;
        RECT 224.400 497.400 228.450 498.450 ;
        RECT 224.400 487.050 225.450 497.400 ;
        RECT 223.950 484.950 226.050 487.050 ;
      LAYER metal3 ;
        RECT 460.950 786.600 463.050 787.050 ;
        RECT 481.950 786.600 484.050 787.200 ;
        RECT 460.950 785.400 484.050 786.600 ;
        RECT 460.950 784.950 463.050 785.400 ;
        RECT 481.950 785.100 484.050 785.400 ;
        RECT 454.950 735.600 457.050 736.050 ;
        RECT 460.950 735.600 463.050 736.050 ;
        RECT 454.950 734.400 463.050 735.600 ;
        RECT 454.950 733.950 457.050 734.400 ;
        RECT 460.950 733.950 463.050 734.400 ;
        RECT 439.950 714.600 442.050 715.050 ;
        RECT 454.950 714.600 457.050 715.050 ;
        RECT 439.950 713.400 457.050 714.600 ;
        RECT 439.950 712.950 442.050 713.400 ;
        RECT 454.950 712.950 457.050 713.400 ;
        RECT 427.950 663.600 430.050 664.050 ;
        RECT 439.950 663.600 442.050 664.050 ;
        RECT 427.950 662.400 442.050 663.600 ;
        RECT 427.950 661.950 430.050 662.400 ;
        RECT 439.950 661.950 442.050 662.400 ;
        RECT 427.950 642.600 430.050 643.050 ;
        RECT 469.950 642.600 472.050 643.050 ;
        RECT 475.950 642.600 478.050 642.900 ;
        RECT 427.950 641.400 478.050 642.600 ;
        RECT 427.950 640.950 430.050 641.400 ;
        RECT 469.950 640.950 472.050 641.400 ;
        RECT 475.950 640.800 478.050 641.400 ;
        RECT 403.950 636.600 406.050 637.050 ;
        RECT 427.950 636.600 430.050 637.050 ;
        RECT 403.950 635.400 430.050 636.600 ;
        RECT 403.950 634.950 406.050 635.400 ;
        RECT 427.950 634.950 430.050 635.400 ;
        RECT 475.950 606.600 478.050 607.050 ;
        RECT 493.950 606.600 496.050 607.050 ;
        RECT 475.950 605.400 496.050 606.600 ;
        RECT 475.950 604.950 478.050 605.400 ;
        RECT 493.950 604.950 496.050 605.400 ;
        RECT 493.950 594.600 496.050 595.050 ;
        RECT 493.950 593.400 534.600 594.600 ;
        RECT 493.950 592.950 496.050 593.400 ;
        RECT 533.400 591.600 534.600 593.400 ;
        RECT 547.950 591.600 550.050 592.050 ;
        RECT 533.400 590.400 550.050 591.600 ;
        RECT 547.950 589.950 550.050 590.400 ;
        RECT 373.950 579.600 376.050 580.050 ;
        RECT 403.950 579.600 406.050 580.050 ;
        RECT 373.950 578.400 406.050 579.600 ;
        RECT 373.950 577.950 376.050 578.400 ;
        RECT 403.950 577.950 406.050 578.400 ;
        RECT 472.950 576.600 475.050 577.050 ;
        RECT 493.950 576.600 496.050 577.050 ;
        RECT 472.950 575.400 496.050 576.600 ;
        RECT 472.950 574.950 475.050 575.400 ;
        RECT 493.950 574.950 496.050 575.400 ;
        RECT 274.950 570.600 277.050 571.050 ;
        RECT 286.950 570.600 289.050 571.050 ;
        RECT 310.950 570.600 313.050 571.050 ;
        RECT 274.950 569.400 313.050 570.600 ;
        RECT 274.950 568.950 277.050 569.400 ;
        RECT 286.950 568.950 289.050 569.400 ;
        RECT 310.950 568.950 313.050 569.400 ;
        RECT 310.950 552.600 313.050 553.050 ;
        RECT 373.950 552.600 376.050 553.050 ;
        RECT 310.950 551.400 376.050 552.600 ;
        RECT 310.950 550.950 313.050 551.400 ;
        RECT 373.950 550.950 376.050 551.400 ;
        RECT 175.950 549.600 178.050 550.050 ;
        RECT 190.800 549.600 192.900 550.050 ;
        RECT 175.950 548.400 192.900 549.600 ;
        RECT 175.950 547.950 178.050 548.400 ;
        RECT 190.800 547.950 192.900 548.400 ;
        RECT 547.950 543.600 550.050 544.050 ;
        RECT 562.950 543.600 565.050 544.050 ;
        RECT 547.950 542.400 565.050 543.600 ;
        RECT 547.950 541.950 550.050 542.400 ;
        RECT 562.950 541.950 565.050 542.400 ;
        RECT 190.950 522.600 193.050 526.200 ;
        RECT 205.950 522.600 208.050 523.050 ;
        RECT 190.950 522.000 208.050 522.600 ;
        RECT 191.400 521.400 208.050 522.000 ;
        RECT 205.950 520.950 208.050 521.400 ;
        RECT 226.950 522.600 229.050 523.050 ;
        RECT 286.950 522.600 289.050 523.050 ;
        RECT 226.950 521.400 289.050 522.600 ;
        RECT 226.950 520.950 229.050 521.400 ;
        RECT 286.950 520.950 289.050 521.400 ;
        RECT 205.950 516.600 208.050 517.050 ;
        RECT 226.950 516.600 229.050 517.050 ;
        RECT 205.950 515.400 229.050 516.600 ;
        RECT 205.950 514.950 208.050 515.400 ;
        RECT 226.950 514.950 229.050 515.400 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 640.950 798.450 643.050 799.050 ;
        RECT 645.000 798.450 649.050 799.050 ;
        RECT 640.950 797.550 649.050 798.450 ;
        RECT 640.950 796.950 643.050 797.550 ;
        RECT 645.000 796.950 649.050 797.550 ;
        RECT 133.950 763.950 136.050 766.050 ;
        RECT 337.950 685.950 343.050 688.050 ;
        RECT 547.950 682.950 550.050 685.050 ;
        RECT 154.950 640.800 157.050 643.050 ;
        RECT 595.950 640.950 598.050 643.050 ;
        RECT 205.950 531.450 208.050 532.050 ;
        RECT 210.000 531.450 214.050 532.050 ;
        RECT 205.950 530.550 214.050 531.450 ;
        RECT 205.950 529.950 208.050 530.550 ;
        RECT 210.000 529.950 214.050 530.550 ;
        RECT 199.950 451.950 202.050 454.050 ;
      LAYER metal2 ;
        RECT 638.400 823.050 639.450 828.450 ;
        RECT 637.950 820.950 640.050 823.050 ;
        RECT 646.950 820.950 649.050 823.050 ;
        RECT 647.400 799.050 648.450 820.950 ;
        RECT 640.950 796.950 643.050 799.050 ;
        RECT 646.950 796.950 649.050 799.050 ;
        RECT 641.400 781.050 642.450 796.950 ;
        RECT 631.950 778.950 634.050 781.050 ;
        RECT 640.950 778.950 643.050 781.050 ;
        RECT 133.950 763.950 136.050 766.050 ;
        RECT 134.400 754.050 135.450 763.950 ;
        RECT 632.400 754.050 633.450 778.950 ;
        RECT 133.950 751.950 136.050 754.050 ;
        RECT 604.950 751.950 607.050 754.050 ;
        RECT 631.950 751.950 634.050 754.050 ;
        RECT 148.950 748.950 151.050 751.050 ;
        RECT 149.400 712.050 150.450 748.950 ;
        RECT 605.400 736.050 606.450 751.950 ;
        RECT 592.950 733.950 595.050 736.050 ;
        RECT 604.950 733.950 607.050 736.050 ;
        RECT 593.400 712.050 594.450 733.950 ;
        RECT 148.950 709.950 151.050 712.050 ;
        RECT 172.950 709.950 175.050 712.050 ;
        RECT 559.950 709.950 562.050 712.050 ;
        RECT 592.950 709.950 595.050 712.050 ;
        RECT 173.400 673.050 174.450 709.950 ;
        RECT 560.400 705.450 561.450 709.950 ;
        RECT 557.400 704.400 561.450 705.450 ;
        RECT 337.950 685.950 340.050 688.050 ;
        RECT 338.400 673.050 339.450 685.950 ;
        RECT 547.950 679.950 550.050 685.050 ;
        RECT 557.400 682.050 558.450 704.400 ;
        RECT 556.950 679.950 559.050 682.050 ;
        RECT 157.950 670.950 160.050 673.050 ;
        RECT 172.950 670.950 175.050 673.050 ;
        RECT 208.950 670.950 211.050 673.050 ;
        RECT 337.950 670.950 340.050 673.050 ;
        RECT 457.950 670.950 460.050 673.050 ;
        RECT 502.950 670.950 505.050 673.050 ;
        RECT 158.400 643.050 159.450 670.950 ;
        RECT 156.000 642.900 159.450 643.050 ;
        RECT 154.950 641.250 159.450 642.900 ;
        RECT 154.950 640.950 159.000 641.250 ;
        RECT 154.950 640.800 157.050 640.950 ;
        RECT 209.400 588.450 210.450 670.950 ;
        RECT 338.400 655.050 339.450 670.950 ;
        RECT 458.400 655.050 459.450 670.950 ;
        RECT 503.400 664.050 504.450 670.950 ;
        RECT 557.400 664.050 558.450 679.950 ;
        RECT 502.950 661.950 505.050 664.050 ;
        RECT 556.950 661.950 559.050 664.050 ;
        RECT 595.950 661.950 598.050 664.050 ;
        RECT 337.950 652.950 340.050 655.050 ;
        RECT 457.950 652.950 460.050 655.050 ;
        RECT 596.400 643.050 597.450 661.950 ;
        RECT 595.950 640.950 598.050 643.050 ;
        RECT 206.400 587.400 210.450 588.450 ;
        RECT 206.400 580.050 207.450 587.400 ;
        RECT 205.950 577.950 208.050 580.050 ;
        RECT 199.950 574.950 202.050 577.050 ;
        RECT 200.400 564.450 201.450 574.950 ;
        RECT 200.400 563.400 204.450 564.450 ;
        RECT 203.400 532.050 204.450 563.400 ;
        RECT 203.400 530.400 208.050 532.050 ;
        RECT 204.000 529.950 208.050 530.400 ;
        RECT 211.950 529.950 214.050 532.050 ;
        RECT 212.400 487.050 213.450 529.950 ;
        RECT 199.950 484.950 202.050 487.050 ;
        RECT 211.950 484.950 214.050 487.050 ;
        RECT 200.400 454.050 201.450 484.950 ;
        RECT 199.950 451.950 202.050 454.050 ;
      LAYER metal3 ;
        RECT 637.950 822.600 640.050 823.050 ;
        RECT 646.950 822.600 649.050 823.050 ;
        RECT 637.950 821.400 649.050 822.600 ;
        RECT 637.950 820.950 640.050 821.400 ;
        RECT 646.950 820.950 649.050 821.400 ;
        RECT 631.950 780.600 634.050 781.050 ;
        RECT 640.950 780.600 643.050 781.050 ;
        RECT 631.950 779.400 643.050 780.600 ;
        RECT 631.950 778.950 634.050 779.400 ;
        RECT 640.950 778.950 643.050 779.400 ;
        RECT 133.950 753.600 136.050 754.050 ;
        RECT 604.950 753.600 607.050 754.050 ;
        RECT 631.950 753.600 634.050 754.050 ;
        RECT 133.950 752.400 144.600 753.600 ;
        RECT 133.950 751.950 136.050 752.400 ;
        RECT 143.400 750.600 144.600 752.400 ;
        RECT 604.950 752.400 634.050 753.600 ;
        RECT 604.950 751.950 607.050 752.400 ;
        RECT 631.950 751.950 634.050 752.400 ;
        RECT 148.950 750.600 151.050 751.050 ;
        RECT 143.400 749.400 151.050 750.600 ;
        RECT 148.950 748.950 151.050 749.400 ;
        RECT 592.950 735.600 595.050 736.050 ;
        RECT 604.950 735.600 607.050 736.050 ;
        RECT 592.950 734.400 607.050 735.600 ;
        RECT 592.950 733.950 595.050 734.400 ;
        RECT 604.950 733.950 607.050 734.400 ;
        RECT 148.950 711.600 151.050 712.050 ;
        RECT 172.950 711.600 175.050 712.050 ;
        RECT 148.950 710.400 175.050 711.600 ;
        RECT 148.950 709.950 151.050 710.400 ;
        RECT 172.950 709.950 175.050 710.400 ;
        RECT 559.950 711.600 562.050 712.050 ;
        RECT 592.950 711.600 595.050 712.050 ;
        RECT 559.950 710.400 595.050 711.600 ;
        RECT 559.950 709.950 562.050 710.400 ;
        RECT 592.950 709.950 595.050 710.400 ;
        RECT 547.950 681.600 550.050 682.050 ;
        RECT 556.950 681.600 559.050 682.050 ;
        RECT 547.950 680.400 559.050 681.600 ;
        RECT 547.950 679.950 550.050 680.400 ;
        RECT 556.950 679.950 559.050 680.400 ;
        RECT 157.950 672.600 160.050 673.050 ;
        RECT 172.950 672.600 175.050 673.050 ;
        RECT 208.950 672.600 211.050 673.050 ;
        RECT 337.950 672.600 340.050 673.050 ;
        RECT 157.950 671.400 340.050 672.600 ;
        RECT 157.950 670.950 160.050 671.400 ;
        RECT 172.950 670.950 175.050 671.400 ;
        RECT 208.950 670.950 211.050 671.400 ;
        RECT 337.950 670.950 340.050 671.400 ;
        RECT 457.950 672.600 460.050 673.050 ;
        RECT 502.950 672.600 505.050 673.050 ;
        RECT 457.950 671.400 505.050 672.600 ;
        RECT 457.950 670.950 460.050 671.400 ;
        RECT 502.950 670.950 505.050 671.400 ;
        RECT 502.950 663.600 505.050 664.050 ;
        RECT 556.950 663.600 559.050 664.050 ;
        RECT 595.950 663.600 598.050 664.050 ;
        RECT 502.950 662.400 598.050 663.600 ;
        RECT 502.950 661.950 505.050 662.400 ;
        RECT 556.950 661.950 559.050 662.400 ;
        RECT 595.950 661.950 598.050 662.400 ;
        RECT 337.950 654.600 340.050 655.050 ;
        RECT 457.950 654.600 460.050 655.050 ;
        RECT 337.950 653.400 460.050 654.600 ;
        RECT 337.950 652.950 340.050 653.400 ;
        RECT 457.950 652.950 460.050 653.400 ;
        RECT 204.000 579.600 208.050 580.050 ;
        RECT 203.400 577.950 208.050 579.600 ;
        RECT 203.400 577.050 204.600 577.950 ;
        RECT 199.950 575.400 204.600 577.050 ;
        RECT 199.950 574.950 204.000 575.400 ;
        RECT 199.950 486.600 202.050 487.050 ;
        RECT 211.950 486.600 214.050 487.050 ;
        RECT 199.950 485.400 214.050 486.600 ;
        RECT 199.950 484.950 202.050 485.400 ;
        RECT 211.950 484.950 214.050 485.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal1 ;
        RECT 661.950 802.950 664.050 808.050 ;
        RECT 157.950 724.950 160.050 727.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 193.950 646.950 196.050 649.050 ;
      LAYER metal2 ;
        RECT 656.400 814.050 657.450 828.450 ;
        RECT 655.950 811.950 658.050 814.050 ;
        RECT 661.950 811.950 664.050 814.050 ;
        RECT 662.400 808.050 663.450 811.950 ;
        RECT 661.950 805.950 664.050 808.050 ;
        RECT 662.400 748.050 663.450 805.950 ;
        RECT 457.950 745.050 460.050 748.050 ;
        RECT 661.950 745.950 664.050 748.050 ;
        RECT 442.950 742.950 445.050 745.050 ;
        RECT 454.950 744.000 460.050 745.050 ;
        RECT 454.950 743.400 459.450 744.000 ;
        RECT 454.950 742.950 459.000 743.400 ;
        RECT 166.950 730.950 169.050 733.050 ;
        RECT 167.400 727.050 168.450 730.950 ;
        RECT 205.950 730.800 208.050 732.900 ;
        RECT 157.950 724.950 163.050 727.050 ;
        RECT 166.950 724.950 169.050 727.050 ;
        RECT 206.400 658.050 207.450 730.800 ;
        RECT 443.400 730.050 444.450 742.950 ;
        RECT 442.950 727.950 445.050 730.050 ;
        RECT 436.950 724.950 439.050 727.050 ;
        RECT 437.400 703.050 438.450 724.950 ;
        RECT 436.950 700.950 439.050 703.050 ;
        RECT 469.950 700.950 472.050 703.050 ;
        RECT 470.400 682.050 471.450 700.950 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 193.950 655.950 196.050 658.050 ;
        RECT 205.950 655.950 208.050 658.050 ;
        RECT 194.400 649.050 195.450 655.950 ;
        RECT 193.950 646.950 196.050 649.050 ;
      LAYER metal3 ;
        RECT 655.950 813.600 658.050 814.050 ;
        RECT 661.950 813.600 664.050 814.050 ;
        RECT 655.950 812.400 664.050 813.600 ;
        RECT 655.950 811.950 658.050 812.400 ;
        RECT 661.950 811.950 664.050 812.400 ;
        RECT 457.950 747.600 460.050 748.050 ;
        RECT 661.950 747.600 664.050 748.050 ;
        RECT 457.950 746.400 664.050 747.600 ;
        RECT 457.950 745.950 460.050 746.400 ;
        RECT 661.950 745.950 664.050 746.400 ;
        RECT 442.950 744.600 445.050 745.050 ;
        RECT 454.950 744.600 457.050 745.050 ;
        RECT 442.950 743.400 457.050 744.600 ;
        RECT 442.950 742.950 445.050 743.400 ;
        RECT 454.950 742.950 457.050 743.400 ;
        RECT 166.950 732.600 169.050 733.050 ;
        RECT 205.950 732.600 208.050 732.900 ;
        RECT 166.950 731.400 444.600 732.600 ;
        RECT 166.950 730.950 169.050 731.400 ;
        RECT 205.950 730.800 208.050 731.400 ;
        RECT 443.400 730.050 444.600 731.400 ;
        RECT 442.950 729.600 445.050 730.050 ;
        RECT 437.400 729.000 445.050 729.600 ;
        RECT 436.950 728.400 445.050 729.000 ;
        RECT 160.950 726.600 163.050 727.050 ;
        RECT 166.950 726.600 169.050 727.050 ;
        RECT 160.950 725.400 169.050 726.600 ;
        RECT 160.950 724.950 163.050 725.400 ;
        RECT 166.950 724.950 169.050 725.400 ;
        RECT 436.950 724.950 439.050 728.400 ;
        RECT 442.950 727.950 445.050 728.400 ;
        RECT 436.950 702.600 439.050 703.050 ;
        RECT 469.950 702.600 472.050 703.050 ;
        RECT 436.950 701.400 472.050 702.600 ;
        RECT 436.950 700.950 439.050 701.400 ;
        RECT 469.950 700.950 472.050 701.400 ;
        RECT 193.950 657.600 196.050 658.050 ;
        RECT 205.950 657.600 208.050 658.050 ;
        RECT 193.950 656.400 208.050 657.600 ;
        RECT 193.950 655.950 196.050 656.400 ;
        RECT 205.950 655.950 208.050 656.400 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal1 ;
        RECT 172.950 802.950 175.050 805.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 244.950 523.950 247.050 526.050 ;
      LAYER metal2 ;
        RECT 662.400 820.050 663.450 828.450 ;
        RECT 661.950 817.950 664.050 820.050 ;
        RECT 670.950 817.950 673.050 820.050 ;
        RECT 171.000 804.450 175.050 805.050 ;
        RECT 170.400 802.950 175.050 804.450 ;
        RECT 170.400 754.050 171.450 802.950 ;
        RECT 154.950 751.950 157.050 754.050 ;
        RECT 169.950 751.950 172.050 754.050 ;
        RECT 155.400 652.050 156.450 751.950 ;
        RECT 671.400 697.050 672.450 817.950 ;
        RECT 505.950 694.950 508.050 697.050 ;
        RECT 670.950 694.950 673.050 697.050 ;
        RECT 506.400 682.050 507.450 694.950 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 506.400 670.050 507.450 679.950 ;
        RECT 361.950 667.950 364.050 670.050 ;
        RECT 505.950 667.950 508.050 670.050 ;
        RECT 362.400 661.050 363.450 667.950 ;
        RECT 283.950 658.950 286.050 661.050 ;
        RECT 361.950 658.950 364.050 661.050 ;
        RECT 284.400 652.050 285.450 658.950 ;
        RECT 154.950 649.950 157.050 652.050 ;
        RECT 283.950 649.950 286.050 652.050 ;
        RECT 155.400 646.200 156.450 649.950 ;
        RECT 155.100 644.100 157.200 646.200 ;
        RECT 151.950 640.800 154.050 642.900 ;
        RECT 152.400 589.050 153.450 640.800 ;
        RECT 151.950 586.950 154.050 589.050 ;
        RECT 160.950 586.950 163.050 589.050 ;
        RECT 244.950 586.950 247.050 589.050 ;
        RECT 161.400 571.050 162.450 586.950 ;
        RECT 160.950 568.950 163.050 571.050 ;
        RECT 245.400 526.050 246.450 586.950 ;
        RECT 244.950 523.950 247.050 526.050 ;
      LAYER metal3 ;
        RECT 661.950 819.600 664.050 820.050 ;
        RECT 670.950 819.600 673.050 820.050 ;
        RECT 661.950 818.400 673.050 819.600 ;
        RECT 661.950 817.950 664.050 818.400 ;
        RECT 670.950 817.950 673.050 818.400 ;
        RECT 154.950 753.600 157.050 754.050 ;
        RECT 169.950 753.600 172.050 754.050 ;
        RECT 154.950 752.400 172.050 753.600 ;
        RECT 154.950 751.950 157.050 752.400 ;
        RECT 169.950 751.950 172.050 752.400 ;
        RECT 505.950 696.600 508.050 697.050 ;
        RECT 670.950 696.600 673.050 697.050 ;
        RECT 505.950 695.400 673.050 696.600 ;
        RECT 505.950 694.950 508.050 695.400 ;
        RECT 670.950 694.950 673.050 695.400 ;
        RECT 361.950 669.600 364.050 670.050 ;
        RECT 505.950 669.600 508.050 670.050 ;
        RECT 361.950 668.400 508.050 669.600 ;
        RECT 361.950 667.950 364.050 668.400 ;
        RECT 505.950 667.950 508.050 668.400 ;
        RECT 283.950 660.600 286.050 661.050 ;
        RECT 361.950 660.600 364.050 661.050 ;
        RECT 283.950 659.400 364.050 660.600 ;
        RECT 283.950 658.950 286.050 659.400 ;
        RECT 361.950 658.950 364.050 659.400 ;
        RECT 154.950 651.600 157.050 652.050 ;
        RECT 283.950 651.600 286.050 652.050 ;
        RECT 154.950 650.400 286.050 651.600 ;
        RECT 154.950 649.950 157.050 650.400 ;
        RECT 283.950 649.950 286.050 650.400 ;
        RECT 155.100 645.000 157.200 646.200 ;
        RECT 154.950 644.100 157.200 645.000 ;
        RECT 154.950 643.050 157.050 644.100 ;
        RECT 153.000 642.900 157.050 643.050 ;
        RECT 151.950 642.000 157.050 642.900 ;
        RECT 151.950 641.400 156.600 642.000 ;
        RECT 151.950 640.950 156.000 641.400 ;
        RECT 151.950 640.800 154.050 640.950 ;
        RECT 151.950 588.600 154.050 589.050 ;
        RECT 160.950 588.600 163.050 589.050 ;
        RECT 244.950 588.600 247.050 589.050 ;
        RECT 151.950 587.400 247.050 588.600 ;
        RECT 151.950 586.950 154.050 587.400 ;
        RECT 160.950 586.950 163.050 587.400 ;
        RECT 244.950 586.950 247.050 587.400 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal1 ;
        RECT 13.950 292.950 16.050 295.050 ;
      LAYER metal2 ;
        RECT 13.950 292.950 19.050 295.050 ;
      LAYER metal3 ;
        RECT 16.950 294.600 19.050 295.050 ;
        RECT -3.600 293.400 19.050 294.600 ;
        RECT 16.950 292.950 19.050 293.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal1 ;
        RECT 820.950 52.950 823.050 55.050 ;
      LAYER metal2 ;
        RECT 820.950 58.950 823.050 61.050 ;
        RECT 821.400 55.050 822.450 58.950 ;
        RECT 820.950 52.950 823.050 55.050 ;
      LAYER metal3 ;
        RECT 820.950 60.600 823.050 61.050 ;
        RECT 820.950 59.400 837.600 60.600 ;
        RECT 820.950 58.950 823.050 59.400 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal1 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 436.950 484.950 439.050 487.200 ;
      LAYER metal2 ;
        RECT 7.950 532.950 10.050 535.050 ;
        RECT 8.400 511.050 9.450 532.950 ;
        RECT 7.950 508.950 10.050 511.050 ;
        RECT 88.950 508.950 91.050 511.050 ;
        RECT 89.400 475.050 90.450 508.950 ;
        RECT 406.950 499.950 409.050 502.050 ;
        RECT 436.950 499.950 439.050 502.050 ;
        RECT 407.400 487.050 408.450 499.950 ;
        RECT 437.400 487.200 438.450 499.950 ;
        RECT 406.950 484.950 409.050 487.050 ;
        RECT 436.950 485.100 439.050 487.200 ;
        RECT 407.400 475.050 408.450 484.950 ;
        RECT 88.950 472.950 91.050 475.050 ;
        RECT 406.950 472.950 409.050 475.050 ;
      LAYER metal3 ;
        RECT 7.950 534.600 10.050 535.050 ;
        RECT -3.600 533.400 10.050 534.600 ;
        RECT 7.950 532.950 10.050 533.400 ;
        RECT 7.950 510.600 10.050 511.050 ;
        RECT 88.950 510.600 91.050 511.050 ;
        RECT 7.950 509.400 91.050 510.600 ;
        RECT 7.950 508.950 10.050 509.400 ;
        RECT 88.950 508.950 91.050 509.400 ;
        RECT 406.950 501.600 409.050 502.050 ;
        RECT 436.950 501.600 439.050 502.050 ;
        RECT 406.950 500.400 439.050 501.600 ;
        RECT 406.950 499.950 409.050 500.400 ;
        RECT 436.950 499.950 439.050 500.400 ;
        RECT 88.950 474.600 91.050 475.050 ;
        RECT 406.950 474.600 409.050 475.050 ;
        RECT 88.950 473.400 409.050 474.600 ;
        RECT 88.950 472.950 91.050 473.400 ;
        RECT 406.950 472.950 409.050 473.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal1 ;
        RECT 361.950 529.950 364.050 535.050 ;
        RECT 433.950 529.950 436.050 532.050 ;
      LAYER metal2 ;
        RECT 1.950 541.950 4.050 544.050 ;
        RECT 361.950 541.950 364.050 544.050 ;
        RECT 433.950 541.950 436.050 544.050 ;
        RECT 2.400 529.050 3.450 541.950 ;
        RECT 362.400 535.050 363.450 541.950 ;
        RECT 361.950 532.950 364.050 535.050 ;
        RECT 434.400 532.050 435.450 541.950 ;
        RECT 433.950 529.950 436.050 532.050 ;
        RECT 1.950 526.950 4.050 529.050 ;
      LAYER metal3 ;
        RECT 1.950 543.600 4.050 544.050 ;
        RECT 361.950 543.600 364.050 544.050 ;
        RECT 433.950 543.600 436.050 544.050 ;
        RECT 1.950 542.400 436.050 543.600 ;
        RECT 1.950 541.950 4.050 542.400 ;
        RECT 361.950 541.950 364.050 542.400 ;
        RECT 433.950 541.950 436.050 542.400 ;
        RECT 1.950 528.600 4.050 529.050 ;
        RECT -3.600 527.400 4.050 528.600 ;
        RECT 1.950 526.950 4.050 527.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 304.950 484.950 307.050 487.050 ;
        RECT 331.950 484.950 334.050 487.050 ;
        RECT 305.550 483.000 306.450 484.950 ;
        RECT 304.950 478.950 307.050 483.000 ;
      LAYER metal2 ;
        RECT 1.950 487.950 4.050 490.050 ;
        RECT 2.400 478.050 3.450 487.950 ;
        RECT 304.950 478.950 307.050 484.050 ;
        RECT 331.950 481.950 334.050 487.050 ;
        RECT 1.950 475.950 4.050 478.050 ;
        RECT 76.950 475.950 79.050 478.050 ;
        RECT 77.400 469.050 78.450 475.950 ;
        RECT 305.400 472.050 306.450 478.950 ;
        RECT 304.950 469.950 307.050 472.050 ;
        RECT 76.950 466.950 79.050 469.050 ;
      LAYER metal3 ;
        RECT 1.950 489.600 4.050 490.050 ;
        RECT -3.600 488.400 4.050 489.600 ;
        RECT 1.950 487.950 4.050 488.400 ;
        RECT 304.950 483.600 307.050 484.050 ;
        RECT 331.950 483.600 334.050 484.050 ;
        RECT 304.950 482.400 334.050 483.600 ;
        RECT 304.950 481.950 307.050 482.400 ;
        RECT 331.950 481.950 334.050 482.400 ;
        RECT 1.950 477.600 4.050 478.050 ;
        RECT 76.950 477.600 79.050 478.050 ;
        RECT 1.950 476.400 79.050 477.600 ;
        RECT 1.950 475.950 4.050 476.400 ;
        RECT 76.950 475.950 79.050 476.400 ;
        RECT 304.950 471.600 307.050 472.050 ;
        RECT 221.400 470.400 307.050 471.600 ;
        RECT 76.950 468.600 79.050 469.050 ;
        RECT 221.400 468.600 222.600 470.400 ;
        RECT 304.950 469.950 307.050 470.400 ;
        RECT 76.950 467.400 222.600 468.600 ;
        RECT 76.950 466.950 79.050 467.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal1 ;
        RECT 328.950 406.950 334.050 409.050 ;
        RECT 406.950 406.950 409.050 409.050 ;
      LAYER metal2 ;
        RECT 4.950 409.950 7.050 412.050 ;
        RECT 5.400 403.050 6.450 409.950 ;
        RECT 328.950 406.950 334.050 409.050 ;
        RECT 403.950 406.950 409.050 409.050 ;
        RECT 329.400 403.050 330.450 406.950 ;
        RECT 4.950 400.950 7.050 403.050 ;
        RECT 328.950 400.950 331.050 403.050 ;
      LAYER metal3 ;
        RECT 4.950 411.600 7.050 412.050 ;
        RECT -3.600 410.400 7.050 411.600 ;
        RECT 4.950 409.950 7.050 410.400 ;
        RECT 328.950 408.600 331.050 409.050 ;
        RECT 403.950 408.600 406.050 409.050 ;
        RECT 328.950 407.400 406.050 408.600 ;
        RECT 328.950 406.950 331.050 407.400 ;
        RECT 403.950 406.950 406.050 407.400 ;
        RECT 4.950 402.600 7.050 403.050 ;
        RECT 328.950 402.600 331.050 403.050 ;
        RECT 4.950 401.400 331.050 402.600 ;
        RECT 4.950 400.950 7.050 401.400 ;
        RECT 328.950 400.950 331.050 401.400 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal1 ;
        RECT 682.950 571.950 688.050 574.050 ;
      LAYER metal2 ;
        RECT 685.950 571.950 688.050 574.050 ;
        RECT 686.400 556.050 687.450 571.950 ;
        RECT 829.950 565.950 832.050 568.050 ;
        RECT 830.400 556.050 831.450 565.950 ;
        RECT 685.950 553.950 688.050 556.050 ;
        RECT 829.950 553.950 832.050 556.050 ;
      LAYER metal3 ;
        RECT 829.950 567.600 832.050 568.050 ;
        RECT 829.950 566.400 837.600 567.600 ;
        RECT 829.950 565.950 832.050 566.400 ;
        RECT 685.950 555.600 688.050 556.050 ;
        RECT 829.950 555.600 832.050 556.050 ;
        RECT 685.950 554.400 832.050 555.600 ;
        RECT 685.950 553.950 688.050 554.400 ;
        RECT 829.950 553.950 832.050 554.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal1 ;
        RECT 820.950 520.950 826.050 523.050 ;
      LAYER metal2 ;
        RECT 823.950 526.950 826.050 529.050 ;
        RECT 824.400 523.050 825.450 526.950 ;
        RECT 823.950 520.950 826.050 523.050 ;
      LAYER metal3 ;
        RECT 823.950 528.600 826.050 529.050 ;
        RECT 823.950 527.400 837.600 528.600 ;
        RECT 823.950 526.950 826.050 527.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal1 ;
        RECT 793.950 27.450 796.050 28.050 ;
        RECT 798.000 27.450 802.050 28.050 ;
        RECT 793.950 26.550 802.050 27.450 ;
        RECT 793.950 25.950 796.050 26.550 ;
        RECT 798.000 25.950 802.050 26.550 ;
      LAYER metal2 ;
        RECT 829.950 454.950 832.050 457.050 ;
        RECT 830.400 49.050 831.450 454.950 ;
        RECT 799.950 46.950 802.050 49.050 ;
        RECT 829.950 46.950 832.050 49.050 ;
        RECT 800.400 28.050 801.450 46.950 ;
        RECT 799.950 25.950 802.050 28.050 ;
      LAYER metal3 ;
        RECT 829.950 456.600 832.050 457.050 ;
        RECT 829.950 455.400 837.600 456.600 ;
        RECT 829.950 454.950 832.050 455.400 ;
        RECT 799.950 48.600 802.050 49.050 ;
        RECT 829.950 48.600 832.050 49.050 ;
        RECT 799.950 47.400 832.050 48.600 ;
        RECT 799.950 46.950 802.050 47.400 ;
        RECT 829.950 46.950 832.050 47.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal1 ;
        RECT 823.950 442.950 829.050 445.050 ;
      LAYER metal2 ;
        RECT 826.950 448.950 829.050 451.050 ;
        RECT 827.400 445.050 828.450 448.950 ;
        RECT 826.950 442.950 829.050 445.050 ;
      LAYER metal3 ;
        RECT 826.950 450.600 829.050 451.050 ;
        RECT 826.950 449.400 837.600 450.600 ;
        RECT 826.950 448.950 829.050 449.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal1 ;
        RECT 532.950 25.950 535.050 28.050 ;
      LAYER metal2 ;
        RECT 532.950 25.950 535.050 28.050 ;
        RECT 533.400 -2.550 534.450 25.950 ;
        RECT 530.400 -3.600 534.450 -2.550 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal1 ;
        RECT 691.950 54.450 696.000 55.050 ;
        RECT 697.950 54.450 700.050 55.050 ;
        RECT 691.950 53.550 700.050 54.450 ;
        RECT 691.950 52.950 696.000 53.550 ;
        RECT 697.950 52.950 700.050 53.550 ;
      LAYER metal2 ;
        RECT 691.950 52.950 694.050 55.050 ;
        RECT 692.400 7.050 693.450 52.950 ;
        RECT 691.950 4.950 694.050 7.050 ;
        RECT 700.950 4.950 703.050 7.050 ;
        RECT 701.400 -3.600 702.450 4.950 ;
      LAYER metal3 ;
        RECT 691.950 6.600 694.050 7.050 ;
        RECT 700.950 6.600 703.050 7.050 ;
        RECT 691.950 5.400 703.050 6.600 ;
        RECT 691.950 4.950 694.050 5.400 ;
        RECT 700.950 4.950 703.050 5.400 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal1 ;
        RECT 811.950 205.800 814.050 211.050 ;
      LAYER metal2 ;
        RECT 811.950 205.800 814.050 207.900 ;
        RECT 812.400 187.050 813.450 205.800 ;
        RECT 811.950 184.950 814.050 187.050 ;
        RECT 823.950 184.950 826.050 187.050 ;
        RECT 824.400 7.050 825.450 184.950 ;
        RECT 808.950 4.950 811.050 7.050 ;
        RECT 823.950 4.950 826.050 7.050 ;
        RECT 809.400 -3.600 810.450 4.950 ;
      LAYER metal3 ;
        RECT 811.950 186.600 814.050 187.050 ;
        RECT 823.950 186.600 826.050 187.050 ;
        RECT 811.950 185.400 826.050 186.600 ;
        RECT 811.950 184.950 814.050 185.400 ;
        RECT 823.950 184.950 826.050 185.400 ;
        RECT 808.950 6.600 811.050 7.050 ;
        RECT 823.950 6.600 826.050 7.050 ;
        RECT 808.950 5.400 826.050 6.600 ;
        RECT 808.950 4.950 811.050 5.400 ;
        RECT 823.950 4.950 826.050 5.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal1 ;
        RECT 625.950 127.950 628.050 133.050 ;
      LAYER metal2 ;
        RECT 625.950 127.950 628.050 130.050 ;
        RECT 626.400 70.050 627.450 127.950 ;
        RECT 625.950 67.950 628.050 70.050 ;
        RECT 637.950 67.950 640.050 70.050 ;
        RECT 638.400 4.050 639.450 67.950 ;
        RECT 637.950 1.950 640.050 4.050 ;
        RECT 814.950 1.950 817.050 4.050 ;
        RECT 815.400 -3.600 816.450 1.950 ;
      LAYER metal3 ;
        RECT 625.950 69.600 628.050 70.050 ;
        RECT 637.950 69.600 640.050 70.050 ;
        RECT 625.950 68.400 640.050 69.600 ;
        RECT 625.950 67.950 628.050 68.400 ;
        RECT 637.950 67.950 640.050 68.400 ;
        RECT 637.950 3.600 640.050 4.050 ;
        RECT 814.950 3.600 817.050 4.050 ;
        RECT 637.950 2.400 817.050 3.600 ;
        RECT 637.950 1.950 640.050 2.400 ;
        RECT 814.950 1.950 817.050 2.400 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal1 ;
        RECT 424.950 25.950 427.050 28.050 ;
      LAYER metal2 ;
        RECT 424.950 25.950 427.050 28.050 ;
        RECT 425.400 -3.600 426.450 25.950 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal1 ;
        RECT 460.950 25.950 463.050 28.050 ;
      LAYER metal2 ;
        RECT 460.950 25.950 463.050 28.050 ;
        RECT 461.400 -3.600 462.450 25.950 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal1 ;
        RECT 502.950 25.950 505.050 28.050 ;
      LAYER metal2 ;
        RECT 502.950 25.950 505.050 28.050 ;
        RECT 503.400 -2.550 504.450 25.950 ;
        RECT 500.400 -3.600 504.450 -2.550 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal1 ;
        RECT 517.950 25.950 520.050 28.050 ;
      LAYER metal2 ;
        RECT 517.950 25.950 520.050 28.050 ;
        RECT 518.400 -2.550 519.450 25.950 ;
        RECT 515.400 -3.600 519.450 -2.550 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 274.950 369.450 277.050 370.050 ;
        RECT 280.950 369.450 283.050 373.050 ;
        RECT 274.950 369.000 283.050 369.450 ;
        RECT 274.950 368.550 282.450 369.000 ;
        RECT 274.950 367.950 277.050 368.550 ;
        RECT 358.950 367.950 361.050 370.050 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 469.950 178.950 472.050 181.050 ;
      LAYER metal2 ;
        RECT 665.400 827.400 669.450 828.450 ;
        RECT 665.400 790.050 666.450 827.400 ;
        RECT 637.950 787.950 640.050 790.050 ;
        RECT 664.950 787.950 667.050 790.050 ;
        RECT 638.400 655.050 639.450 787.950 ;
        RECT 511.950 652.950 514.050 655.050 ;
        RECT 637.950 652.950 640.050 655.050 ;
        RECT 512.400 577.200 513.450 652.950 ;
        RECT 502.950 574.950 505.050 577.050 ;
        RECT 511.950 575.100 514.050 577.200 ;
        RECT 503.400 547.050 504.450 574.950 ;
        RECT 484.950 544.950 487.050 547.050 ;
        RECT 502.950 544.950 505.050 547.050 ;
        RECT 485.400 475.050 486.450 544.950 ;
        RECT 484.950 472.950 487.050 475.050 ;
        RECT 514.950 472.950 517.050 475.050 ;
        RECT 515.400 442.050 516.450 472.950 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 596.400 442.050 597.450 445.950 ;
        RECT 514.950 439.950 517.050 442.050 ;
        RECT 595.950 439.950 598.050 442.050 ;
        RECT 515.400 418.050 516.450 439.950 ;
        RECT 397.950 412.950 400.050 418.050 ;
        RECT 514.950 415.950 517.050 418.050 ;
        RECT 398.400 388.050 399.450 412.950 ;
        RECT 358.950 385.950 361.050 388.050 ;
        RECT 397.950 385.950 400.050 388.050 ;
        RECT 274.950 367.950 277.050 370.050 ;
        RECT 280.950 367.950 283.050 373.050 ;
        RECT 359.400 370.050 360.450 385.950 ;
        RECT 355.950 367.950 361.050 370.050 ;
        RECT 275.400 340.050 276.450 367.950 ;
        RECT 262.950 337.950 265.050 340.050 ;
        RECT 274.950 337.950 277.050 340.050 ;
        RECT 263.400 298.050 264.450 337.950 ;
        RECT 262.950 295.950 265.050 298.050 ;
        RECT 271.950 295.950 274.050 298.050 ;
        RECT 272.400 270.450 273.450 295.950 ;
        RECT 272.400 269.400 276.450 270.450 ;
        RECT 275.400 232.050 276.450 269.400 ;
        RECT 265.950 229.950 268.050 232.050 ;
        RECT 274.950 229.950 277.050 232.050 ;
        RECT 266.400 199.050 267.450 229.950 ;
        RECT 592.950 211.950 595.050 214.050 ;
        RECT 593.400 208.050 594.450 211.950 ;
        RECT 502.950 205.950 505.050 208.050 ;
        RECT 592.950 205.950 595.050 208.050 ;
        RECT 256.950 196.950 259.050 199.050 ;
        RECT 265.950 196.950 268.050 199.050 ;
        RECT 257.400 181.050 258.450 196.950 ;
        RECT 256.950 178.950 259.050 181.050 ;
        RECT 454.950 178.950 457.050 181.050 ;
        RECT 469.950 178.950 472.050 181.050 ;
        RECT 257.400 175.050 258.450 178.950 ;
        RECT 455.400 175.050 456.450 178.950 ;
        RECT 470.400 175.050 471.450 178.950 ;
        RECT 503.400 175.050 504.450 205.950 ;
        RECT 256.950 172.950 259.050 175.050 ;
        RECT 454.950 172.950 457.050 175.050 ;
        RECT 469.950 172.950 472.050 175.050 ;
        RECT 502.950 172.950 505.050 175.050 ;
      LAYER metal3 ;
        RECT 637.950 789.600 640.050 790.050 ;
        RECT 664.950 789.600 667.050 790.050 ;
        RECT 637.950 788.400 667.050 789.600 ;
        RECT 637.950 787.950 640.050 788.400 ;
        RECT 664.950 787.950 667.050 788.400 ;
        RECT 511.950 654.600 514.050 655.050 ;
        RECT 637.950 654.600 640.050 655.050 ;
        RECT 511.950 653.400 640.050 654.600 ;
        RECT 511.950 652.950 514.050 653.400 ;
        RECT 637.950 652.950 640.050 653.400 ;
        RECT 502.950 576.600 505.050 577.050 ;
        RECT 511.950 576.600 514.050 577.200 ;
        RECT 502.950 575.400 514.050 576.600 ;
        RECT 502.950 574.950 505.050 575.400 ;
        RECT 511.950 575.100 514.050 575.400 ;
        RECT 484.950 546.600 487.050 547.050 ;
        RECT 502.950 546.600 505.050 547.050 ;
        RECT 484.950 545.400 505.050 546.600 ;
        RECT 484.950 544.950 487.050 545.400 ;
        RECT 502.950 544.950 505.050 545.400 ;
        RECT 484.950 474.600 487.050 475.050 ;
        RECT 514.950 474.600 517.050 475.050 ;
        RECT 484.950 473.400 517.050 474.600 ;
        RECT 484.950 472.950 487.050 473.400 ;
        RECT 514.950 472.950 517.050 473.400 ;
        RECT 514.950 441.600 517.050 442.050 ;
        RECT 595.950 441.600 598.050 442.050 ;
        RECT 514.950 440.400 598.050 441.600 ;
        RECT 514.950 439.950 517.050 440.400 ;
        RECT 595.950 439.950 598.050 440.400 ;
        RECT 397.950 417.600 400.050 418.050 ;
        RECT 514.950 417.600 517.050 418.050 ;
        RECT 397.950 416.400 517.050 417.600 ;
        RECT 397.950 415.950 400.050 416.400 ;
        RECT 514.950 415.950 517.050 416.400 ;
        RECT 358.950 387.600 361.050 388.050 ;
        RECT 397.950 387.600 400.050 388.050 ;
        RECT 358.950 386.400 400.050 387.600 ;
        RECT 358.950 385.950 361.050 386.400 ;
        RECT 397.950 385.950 400.050 386.400 ;
        RECT 280.950 369.600 283.050 370.050 ;
        RECT 355.950 369.600 358.050 370.050 ;
        RECT 280.950 368.400 358.050 369.600 ;
        RECT 280.950 367.950 283.050 368.400 ;
        RECT 355.950 367.950 358.050 368.400 ;
        RECT 262.950 339.600 265.050 340.050 ;
        RECT 274.950 339.600 277.050 340.050 ;
        RECT 262.950 338.400 277.050 339.600 ;
        RECT 262.950 337.950 265.050 338.400 ;
        RECT 274.950 337.950 277.050 338.400 ;
        RECT 262.950 297.600 265.050 298.050 ;
        RECT 271.950 297.600 274.050 298.050 ;
        RECT 262.950 296.400 274.050 297.600 ;
        RECT 262.950 295.950 265.050 296.400 ;
        RECT 271.950 295.950 274.050 296.400 ;
        RECT 265.950 231.600 268.050 232.050 ;
        RECT 274.950 231.600 277.050 232.050 ;
        RECT 265.950 230.400 277.050 231.600 ;
        RECT 265.950 229.950 268.050 230.400 ;
        RECT 274.950 229.950 277.050 230.400 ;
        RECT 502.950 207.600 505.050 208.050 ;
        RECT 592.950 207.600 595.050 208.050 ;
        RECT 502.950 206.400 595.050 207.600 ;
        RECT 502.950 205.950 505.050 206.400 ;
        RECT 592.950 205.950 595.050 206.400 ;
        RECT 256.950 198.600 259.050 199.050 ;
        RECT 265.950 198.600 268.050 199.050 ;
        RECT 256.950 197.400 268.050 198.600 ;
        RECT 256.950 196.950 259.050 197.400 ;
        RECT 265.950 196.950 268.050 197.400 ;
        RECT 256.950 174.600 259.050 175.050 ;
        RECT 454.950 174.600 457.050 175.050 ;
        RECT 469.950 174.600 472.050 175.050 ;
        RECT 502.950 174.600 505.050 175.050 ;
        RECT 256.950 173.400 505.050 174.600 ;
        RECT 256.950 172.950 259.050 173.400 ;
        RECT 454.950 172.950 457.050 173.400 ;
        RECT 469.950 172.950 472.050 173.400 ;
        RECT 502.950 172.950 505.050 173.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 12.000 814.050 13.800 818.400 ;
        RECT 8.400 812.400 13.800 814.050 ;
        RECT 8.400 809.100 9.300 812.400 ;
        RECT 29.100 810.000 30.900 818.400 ;
        RECT 46.800 815.400 48.600 818.400 ;
        RECT 26.700 808.350 30.900 810.000 ;
        RECT 4.950 805.950 10.050 808.050 ;
        RECT 13.950 805.950 16.050 808.050 ;
        RECT 8.400 795.600 9.300 804.900 ;
        RECT 14.100 804.150 15.900 804.900 ;
        RECT 11.100 803.100 12.900 803.850 ;
        RECT 17.100 803.100 18.900 803.850 ;
        RECT 10.950 799.950 13.050 802.050 ;
        RECT 16.950 799.950 19.050 802.050 ;
        RECT 26.700 800.100 27.600 808.350 ;
        RECT 29.100 806.100 30.900 806.850 ;
        RECT 28.950 802.950 31.050 805.050 ;
        RECT 47.400 803.100 48.600 815.400 ;
        RECT 61.200 814.050 63.000 818.400 ;
        RECT 61.200 812.400 66.600 814.050 ;
        RECT 65.700 809.100 66.600 812.400 ;
        RECT 81.000 811.200 82.800 818.400 ;
        RECT 100.800 815.400 102.600 818.400 ;
        RECT 101.400 812.100 102.600 815.400 ;
        RECT 115.200 811.200 117.000 818.400 ;
        RECT 127.800 812.400 129.600 818.400 ;
        RECT 81.000 810.300 84.600 811.200 ;
        RECT 49.950 805.950 52.050 808.050 ;
        RECT 58.950 805.950 61.050 808.050 ;
        RECT 64.950 807.450 67.050 808.050 ;
        RECT 76.950 807.450 79.050 808.050 ;
        RECT 64.950 806.550 79.050 807.450 ;
        RECT 64.950 805.950 67.050 806.550 ;
        RECT 76.950 805.950 79.050 806.550 ;
        RECT 83.400 806.100 84.600 810.300 ;
        RECT 94.950 810.450 99.000 811.050 ;
        RECT 100.950 810.450 103.050 811.050 ;
        RECT 94.950 809.550 103.050 810.450 ;
        RECT 94.950 808.950 99.000 809.550 ;
        RECT 100.950 808.950 103.050 809.550 ;
        RECT 113.400 810.300 117.000 811.200 ;
        RECT 128.400 810.300 129.600 812.400 ;
        RECT 130.800 813.300 132.600 818.400 ;
        RECT 136.800 813.300 138.600 818.400 ;
        RECT 130.800 811.950 138.600 813.300 ;
        RECT 150.000 811.200 151.800 818.400 ;
        RECT 166.500 812.400 168.300 818.400 ;
        RECT 172.800 815.400 174.600 818.400 ;
        RECT 150.000 810.300 153.600 811.200 ;
        RECT 100.950 806.100 102.300 807.900 ;
        RECT 113.400 806.100 114.600 810.300 ;
        RECT 128.400 809.250 132.150 810.300 ;
        RECT 130.950 809.100 132.150 809.250 ;
        RECT 50.100 804.150 51.900 804.900 ;
        RECT 59.100 804.150 60.900 804.900 ;
        RECT 56.100 803.100 57.900 803.850 ;
        RECT 62.100 803.100 63.900 803.850 ;
        RECT 31.950 799.950 34.050 802.050 ;
        RECT 46.950 799.950 49.050 802.050 ;
        RECT 52.950 799.950 58.050 802.050 ;
        RECT 61.950 799.950 64.050 802.050 ;
        RECT 25.950 796.950 28.050 799.050 ;
        RECT 32.100 798.150 33.900 798.900 ;
        RECT 35.100 797.100 36.900 797.850 ;
        RECT 7.800 783.600 9.600 795.600 ;
        RECT 10.800 794.700 18.600 795.600 ;
        RECT 10.800 783.600 12.600 794.700 ;
        RECT 16.800 783.600 18.600 794.700 ;
        RECT 26.700 790.800 27.600 795.900 ;
        RECT 34.950 793.950 37.050 796.050 ;
        RECT 26.700 789.900 33.300 790.800 ;
        RECT 26.700 789.600 27.600 789.900 ;
        RECT 25.800 783.600 27.600 789.600 ;
        RECT 31.800 789.600 33.300 789.900 ;
        RECT 47.400 789.600 48.600 798.900 ;
        RECT 65.700 795.600 66.600 804.900 ;
        RECT 70.950 804.450 73.050 805.050 ;
        RECT 82.950 804.450 85.050 805.050 ;
        RECT 70.950 803.550 85.050 804.450 ;
        RECT 70.950 802.950 73.050 803.550 ;
        RECT 82.950 802.950 85.050 803.550 ;
        RECT 88.950 804.450 91.050 805.050 ;
        RECT 97.950 804.450 100.050 805.050 ;
        RECT 88.950 803.550 100.050 804.450 ;
        RECT 88.950 802.950 91.050 803.550 ;
        RECT 97.950 802.950 100.050 803.550 ;
        RECT 101.100 801.900 102.300 806.100 ;
        RECT 130.950 805.950 133.050 808.050 ;
        RECT 136.950 805.950 139.050 808.050 ;
        RECT 152.400 806.100 153.600 810.300 ;
        RECT 166.800 809.100 168.000 812.400 ;
        RECT 172.800 811.500 174.000 815.400 ;
        RECT 186.300 814.200 188.100 818.400 ;
        RECT 168.900 810.600 174.000 811.500 ;
        RECT 186.150 812.400 188.100 814.200 ;
        RECT 168.900 809.700 170.850 810.600 ;
        RECT 169.950 809.100 170.850 809.700 ;
        RECT 186.150 809.100 187.050 812.400 ;
        RECT 188.100 810.600 189.900 811.500 ;
        RECT 193.800 810.600 195.600 818.400 ;
        RECT 188.100 809.700 195.600 810.600 ;
        RECT 209.100 810.000 210.900 818.400 ;
        RECT 229.200 814.050 231.000 818.400 ;
        RECT 229.200 812.400 234.600 814.050 ;
        RECT 166.950 805.950 169.050 808.050 ;
        RECT 112.950 802.950 115.050 805.050 ;
        RECT 128.100 803.100 129.900 803.850 ;
        RECT 131.850 803.100 133.050 804.900 ;
        RECT 137.100 804.150 138.900 804.900 ;
        RECT 134.100 803.100 135.900 803.850 ;
        RECT 80.100 800.100 81.900 800.850 ;
        RECT 79.950 796.950 82.050 799.050 ;
        RECT 31.800 783.600 33.600 789.600 ;
        RECT 46.800 783.600 48.600 789.600 ;
        RECT 56.400 794.700 64.200 795.600 ;
        RECT 56.400 783.600 58.200 794.700 ;
        RECT 62.400 783.600 64.200 794.700 ;
        RECT 65.400 783.600 67.200 795.600 ;
        RECT 83.400 789.600 84.600 801.900 ;
        RECT 98.100 801.150 99.900 801.900 ;
        RECT 86.100 800.100 87.900 800.850 ;
        RECT 85.950 796.950 88.050 799.050 ;
        RECT 100.950 796.650 102.300 801.900 ;
        RECT 103.950 799.950 106.050 802.050 ;
        RECT 110.100 800.100 111.900 800.850 ;
        RECT 104.100 798.150 105.900 798.900 ;
        RECT 109.950 796.950 112.050 799.050 ;
        RECT 82.800 783.600 84.600 789.600 ;
        RECT 99.600 795.600 102.300 796.650 ;
        RECT 99.600 783.600 101.400 795.600 ;
        RECT 113.400 789.600 114.600 801.900 ;
        RECT 121.950 801.450 126.000 802.050 ;
        RECT 127.950 801.450 130.050 802.050 ;
        RECT 116.100 800.100 117.900 800.850 ;
        RECT 121.950 800.550 130.050 801.450 ;
        RECT 121.950 799.950 126.000 800.550 ;
        RECT 127.950 799.950 130.050 800.550 ;
        RECT 115.950 796.950 118.050 799.050 ;
        RECT 131.850 798.900 132.900 803.100 ;
        RECT 151.950 802.950 154.050 805.050 ;
        RECT 170.100 804.900 170.850 809.100 ;
        RECT 184.950 805.950 187.050 808.050 ;
        RECT 133.950 799.950 136.050 802.050 ;
        RECT 149.100 800.100 150.900 800.850 ;
        RECT 131.850 795.600 133.050 798.900 ;
        RECT 148.950 796.950 151.050 799.050 ;
        RECT 113.400 783.600 115.200 789.600 ;
        RECT 131.700 783.600 133.500 795.600 ;
        RECT 152.400 789.600 153.600 801.900 ;
        RECT 155.100 800.100 156.900 800.850 ;
        RECT 154.950 796.950 157.050 799.050 ;
        RECT 166.800 795.600 168.000 804.900 ;
        RECT 169.950 798.300 170.850 804.900 ;
        RECT 173.100 801.150 174.900 801.900 ;
        RECT 168.900 797.400 170.850 798.300 ;
        RECT 168.900 796.500 174.600 797.400 ;
        RECT 151.800 783.600 153.600 789.600 ;
        RECT 166.500 783.600 168.300 795.600 ;
        RECT 173.400 789.600 174.600 796.500 ;
        RECT 184.950 795.600 186.000 804.900 ;
        RECT 188.100 803.100 189.900 803.850 ;
        RECT 187.950 799.950 190.050 802.050 ;
        RECT 172.800 783.600 174.600 789.600 ;
        RECT 184.200 783.600 186.000 795.600 ;
        RECT 191.550 789.600 192.600 809.700 ;
        RECT 206.700 808.350 210.900 810.000 ;
        RECT 233.700 809.100 234.600 812.400 ;
        RECT 251.100 810.000 252.900 818.400 ;
        RECT 266.400 813.300 268.200 818.400 ;
        RECT 272.400 813.300 274.200 818.400 ;
        RECT 266.400 811.950 274.200 813.300 ;
        RECT 275.400 812.400 277.200 818.400 ;
        RECT 290.400 815.400 292.200 818.400 ;
        RECT 275.400 810.300 276.600 812.400 ;
        RECT 251.100 808.350 255.300 810.000 ;
        RECT 272.850 809.250 276.600 810.300 ;
        RECT 272.850 809.100 274.050 809.250 ;
        RECT 193.950 802.950 196.050 805.050 ;
        RECT 194.100 801.150 195.900 801.900 ;
        RECT 206.700 800.100 207.600 808.350 ;
        RECT 209.100 806.100 210.900 806.850 ;
        RECT 226.950 805.950 229.050 808.050 ;
        RECT 232.950 807.450 235.050 808.050 ;
        RECT 241.950 807.450 244.050 808.050 ;
        RECT 232.950 806.550 244.050 807.450 ;
        RECT 232.950 805.950 235.050 806.550 ;
        RECT 241.950 805.950 244.050 806.550 ;
        RECT 251.100 806.100 252.900 806.850 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 227.100 804.150 228.900 804.900 ;
        RECT 224.100 803.100 225.900 803.850 ;
        RECT 230.100 803.100 231.900 803.850 ;
        RECT 211.950 799.950 214.050 802.050 ;
        RECT 223.950 799.950 226.050 802.050 ;
        RECT 229.950 799.950 232.050 802.050 ;
        RECT 193.950 798.450 196.050 798.900 ;
        RECT 205.950 798.450 208.050 799.050 ;
        RECT 193.950 797.550 208.050 798.450 ;
        RECT 212.100 798.150 213.900 798.900 ;
        RECT 193.950 796.800 196.050 797.550 ;
        RECT 205.950 796.950 208.050 797.550 ;
        RECT 215.100 797.100 216.900 797.850 ;
        RECT 206.700 790.800 207.600 795.900 ;
        RECT 214.950 793.950 217.050 796.050 ;
        RECT 233.700 795.600 234.600 804.900 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 247.950 799.950 250.050 802.050 ;
        RECT 254.400 800.100 255.300 808.350 ;
        RECT 265.950 805.950 268.050 808.050 ;
        RECT 271.950 807.450 274.050 808.050 ;
        RECT 280.950 807.450 283.050 808.050 ;
        RECT 271.950 806.550 283.050 807.450 ;
        RECT 271.950 805.950 274.050 806.550 ;
        RECT 280.950 805.950 283.050 806.550 ;
        RECT 286.950 805.950 289.050 808.050 ;
        RECT 266.100 804.150 267.900 804.900 ;
        RECT 269.100 803.100 270.900 803.850 ;
        RECT 271.950 803.100 273.150 804.900 ;
        RECT 287.100 804.150 288.900 804.900 ;
        RECT 275.100 803.100 276.900 803.850 ;
        RECT 290.400 803.100 291.600 815.400 ;
        RECT 304.800 812.400 306.600 818.400 ;
        RECT 305.400 810.300 306.600 812.400 ;
        RECT 307.800 813.300 309.600 818.400 ;
        RECT 313.800 813.300 315.600 818.400 ;
        RECT 307.800 811.950 315.600 813.300 ;
        RECT 322.800 812.400 324.600 818.400 ;
        RECT 323.400 810.300 324.600 812.400 ;
        RECT 325.800 813.300 327.600 818.400 ;
        RECT 331.800 813.300 333.600 818.400 ;
        RECT 348.000 814.050 349.800 818.400 ;
        RECT 325.800 811.950 333.600 813.300 ;
        RECT 344.400 812.400 349.800 814.050 ;
        RECT 305.400 809.250 309.150 810.300 ;
        RECT 323.400 809.250 327.150 810.300 ;
        RECT 307.950 809.100 309.150 809.250 ;
        RECT 325.950 809.100 327.150 809.250 ;
        RECT 344.400 809.100 345.300 812.400 ;
        RECT 365.100 810.000 366.900 818.400 ;
        RECT 386.100 810.000 387.900 818.400 ;
        RECT 408.000 814.050 409.800 818.400 ;
        RECT 365.100 808.350 369.300 810.000 ;
        RECT 307.950 805.950 310.050 808.050 ;
        RECT 313.950 805.950 316.050 808.050 ;
        RECT 322.950 805.950 328.050 808.050 ;
        RECT 331.950 805.950 334.050 808.050 ;
        RECT 340.950 805.950 346.050 808.050 ;
        RECT 349.950 805.950 352.050 808.050 ;
        RECT 365.100 806.100 366.900 806.850 ;
        RECT 305.100 803.100 306.900 803.850 ;
        RECT 308.850 803.100 310.050 804.900 ;
        RECT 314.100 804.150 315.900 804.900 ;
        RECT 311.100 803.100 312.900 803.850 ;
        RECT 323.100 803.100 324.900 803.850 ;
        RECT 326.850 803.100 328.050 804.900 ;
        RECT 332.100 804.150 333.900 804.900 ;
        RECT 329.100 803.100 330.900 803.850 ;
        RECT 259.950 801.450 262.050 802.050 ;
        RECT 268.950 801.450 271.050 802.050 ;
        RECT 259.950 800.550 271.050 801.450 ;
        RECT 259.950 799.950 262.050 800.550 ;
        RECT 268.950 799.950 271.050 800.550 ;
        RECT 248.100 798.150 249.900 798.900 ;
        RECT 253.950 798.450 256.050 799.050 ;
        RECT 262.950 798.450 265.050 799.050 ;
        RECT 272.100 798.900 273.150 803.100 ;
        RECT 274.950 799.950 277.050 802.050 ;
        RECT 289.950 799.950 295.050 802.050 ;
        RECT 304.950 799.950 307.050 802.050 ;
        RECT 308.850 798.900 309.900 803.100 ;
        RECT 310.950 799.950 313.050 802.050 ;
        RECT 322.950 799.800 325.050 802.050 ;
        RECT 326.850 798.900 327.900 803.100 ;
        RECT 328.950 799.950 331.050 802.050 ;
        RECT 245.100 797.100 246.900 797.850 ;
        RECT 253.950 797.550 265.050 798.450 ;
        RECT 253.950 796.950 256.050 797.550 ;
        RECT 262.950 796.950 265.050 797.550 ;
        RECT 224.400 794.700 232.200 795.600 ;
        RECT 206.700 789.900 213.300 790.800 ;
        RECT 206.700 789.600 207.600 789.900 ;
        RECT 190.800 783.600 192.600 789.600 ;
        RECT 205.800 783.600 207.600 789.600 ;
        RECT 211.800 789.600 213.300 789.900 ;
        RECT 211.800 783.600 213.600 789.600 ;
        RECT 224.400 783.600 226.200 794.700 ;
        RECT 230.400 783.600 232.200 794.700 ;
        RECT 233.400 783.600 235.200 795.600 ;
        RECT 244.950 793.950 247.050 796.050 ;
        RECT 254.400 790.800 255.300 795.900 ;
        RECT 271.950 795.600 273.150 798.900 ;
        RECT 248.700 789.900 255.300 790.800 ;
        RECT 248.700 789.600 250.200 789.900 ;
        RECT 248.400 783.600 250.200 789.600 ;
        RECT 254.400 789.600 255.300 789.900 ;
        RECT 254.400 783.600 256.200 789.600 ;
        RECT 271.500 783.600 273.300 795.600 ;
        RECT 290.400 789.600 291.600 798.900 ;
        RECT 308.850 795.600 310.050 798.900 ;
        RECT 326.850 795.600 328.050 798.900 ;
        RECT 344.400 795.600 345.300 804.900 ;
        RECT 350.100 804.150 351.900 804.900 ;
        RECT 347.100 803.100 348.900 803.850 ;
        RECT 353.100 803.100 354.900 803.850 ;
        RECT 364.950 802.950 367.050 805.200 ;
        RECT 346.950 799.950 349.050 802.050 ;
        RECT 352.950 799.950 355.050 802.050 ;
        RECT 361.950 799.950 364.050 802.050 ;
        RECT 368.400 800.100 369.300 808.350 ;
        RECT 383.700 808.350 387.900 810.000 ;
        RECT 404.400 812.400 409.800 814.050 ;
        RECT 404.400 809.100 405.300 812.400 ;
        RECT 428.100 810.000 429.900 818.400 ;
        RECT 447.000 814.050 448.800 818.400 ;
        RECT 425.700 808.350 429.900 810.000 ;
        RECT 443.400 812.400 448.800 814.050 ;
        RECT 466.200 814.050 468.000 818.400 ;
        RECT 482.400 815.400 484.200 818.400 ;
        RECT 466.200 812.400 471.600 814.050 ;
        RECT 443.400 809.100 444.300 812.400 ;
        RECT 470.700 809.100 471.600 812.400 ;
        RECT 383.700 800.100 384.600 808.350 ;
        RECT 397.950 807.450 402.000 808.050 ;
        RECT 403.950 807.450 406.050 808.050 ;
        RECT 386.100 806.100 387.900 806.850 ;
        RECT 397.950 806.550 406.050 807.450 ;
        RECT 397.950 805.950 402.000 806.550 ;
        RECT 403.950 805.950 406.050 806.550 ;
        RECT 409.950 805.950 412.050 808.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 388.950 799.950 391.050 802.050 ;
        RECT 362.100 798.150 363.900 798.900 ;
        RECT 359.100 797.100 360.900 797.850 ;
        RECT 367.950 796.950 372.900 799.050 ;
        RECT 373.950 798.450 376.050 799.050 ;
        RECT 382.950 798.450 385.050 799.050 ;
        RECT 373.950 797.550 385.050 798.450 ;
        RECT 389.100 798.150 390.900 798.900 ;
        RECT 373.950 796.950 376.050 797.550 ;
        RECT 382.950 796.950 385.050 797.550 ;
        RECT 392.100 797.100 393.900 797.850 ;
        RECT 290.400 783.600 292.200 789.600 ;
        RECT 308.700 783.600 310.500 795.600 ;
        RECT 326.700 783.600 328.500 795.600 ;
        RECT 343.800 783.600 345.600 795.600 ;
        RECT 346.800 794.700 354.600 795.600 ;
        RECT 346.800 783.600 348.600 794.700 ;
        RECT 352.800 783.600 354.600 794.700 ;
        RECT 358.950 793.950 361.050 796.050 ;
        RECT 368.400 790.800 369.300 795.900 ;
        RECT 362.700 789.900 369.300 790.800 ;
        RECT 362.700 789.600 364.200 789.900 ;
        RECT 362.400 783.600 364.200 789.600 ;
        RECT 368.400 789.600 369.300 789.900 ;
        RECT 383.700 790.800 384.600 795.900 ;
        RECT 391.950 793.950 394.050 796.050 ;
        RECT 404.400 795.600 405.300 804.900 ;
        RECT 410.100 804.150 411.900 804.900 ;
        RECT 407.100 803.100 408.900 803.850 ;
        RECT 413.100 803.100 414.900 803.850 ;
        RECT 406.950 799.950 409.050 802.050 ;
        RECT 412.950 799.950 415.050 802.050 ;
        RECT 425.700 800.100 426.600 808.350 ;
        RECT 433.950 807.450 436.050 808.050 ;
        RECT 442.950 807.450 445.050 808.050 ;
        RECT 428.100 806.100 429.900 806.850 ;
        RECT 433.950 806.550 445.050 807.450 ;
        RECT 433.950 805.950 436.050 806.550 ;
        RECT 442.950 805.950 445.050 806.550 ;
        RECT 448.950 805.950 451.050 808.050 ;
        RECT 454.950 807.450 457.050 808.050 ;
        RECT 463.950 807.450 466.050 808.050 ;
        RECT 454.950 806.550 466.050 807.450 ;
        RECT 454.950 805.950 457.050 806.550 ;
        RECT 463.950 805.950 466.050 806.550 ;
        RECT 469.950 805.950 475.050 808.050 ;
        RECT 478.950 805.950 481.050 808.050 ;
        RECT 427.950 802.950 430.050 805.050 ;
        RECT 430.950 799.950 433.050 802.050 ;
        RECT 418.950 798.450 423.000 799.050 ;
        RECT 424.950 798.450 427.050 799.050 ;
        RECT 418.950 797.550 427.050 798.450 ;
        RECT 431.100 798.150 432.900 798.900 ;
        RECT 418.950 796.950 423.000 797.550 ;
        RECT 424.950 796.950 427.050 797.550 ;
        RECT 434.100 797.100 435.900 797.850 ;
        RECT 383.700 789.900 390.300 790.800 ;
        RECT 383.700 789.600 384.600 789.900 ;
        RECT 368.400 783.600 370.200 789.600 ;
        RECT 382.800 783.600 384.600 789.600 ;
        RECT 388.800 789.600 390.300 789.900 ;
        RECT 388.800 783.600 390.600 789.600 ;
        RECT 403.800 783.600 405.600 795.600 ;
        RECT 406.800 794.700 414.600 795.600 ;
        RECT 406.800 783.600 408.600 794.700 ;
        RECT 412.800 783.600 414.600 794.700 ;
        RECT 425.700 790.800 426.600 795.900 ;
        RECT 433.950 793.950 436.050 796.050 ;
        RECT 443.400 795.600 444.300 804.900 ;
        RECT 449.100 804.150 450.900 804.900 ;
        RECT 464.100 804.150 465.900 804.900 ;
        RECT 446.100 803.100 447.900 803.850 ;
        RECT 452.100 803.100 453.900 803.850 ;
        RECT 461.100 803.100 462.900 803.850 ;
        RECT 467.100 803.100 468.900 803.850 ;
        RECT 445.950 799.950 448.050 802.050 ;
        RECT 451.950 799.950 454.050 802.050 ;
        RECT 460.950 799.950 463.050 802.050 ;
        RECT 466.950 799.950 469.050 802.050 ;
        RECT 470.700 795.600 471.600 804.900 ;
        RECT 479.100 804.150 480.900 804.900 ;
        RECT 482.400 803.100 483.600 815.400 ;
        RECT 493.800 812.400 495.600 818.400 ;
        RECT 494.400 810.300 495.600 812.400 ;
        RECT 496.800 813.300 498.600 818.400 ;
        RECT 502.800 813.300 504.600 818.400 ;
        RECT 496.800 811.950 504.600 813.300 ;
        RECT 512.400 813.300 514.200 818.400 ;
        RECT 518.400 813.300 520.200 818.400 ;
        RECT 512.400 811.950 520.200 813.300 ;
        RECT 521.400 812.400 523.200 818.400 ;
        RECT 521.400 810.300 522.600 812.400 ;
        RECT 494.400 809.250 498.150 810.300 ;
        RECT 496.950 809.100 498.150 809.250 ;
        RECT 518.850 809.250 522.600 810.300 ;
        RECT 539.100 810.000 540.900 818.400 ;
        RECT 556.200 814.050 558.000 818.400 ;
        RECT 556.200 812.400 561.600 814.050 ;
        RECT 518.850 809.100 520.050 809.250 ;
        RECT 539.100 808.350 543.300 810.000 ;
        RECT 560.700 809.100 561.600 812.400 ;
        RECT 572.400 813.300 574.200 818.400 ;
        RECT 578.400 813.300 580.200 818.400 ;
        RECT 572.400 811.950 580.200 813.300 ;
        RECT 581.400 812.400 583.200 818.400 ;
        RECT 581.400 810.300 582.600 812.400 ;
        RECT 578.850 809.250 582.600 810.300 ;
        RECT 599.100 810.000 600.900 818.400 ;
        RECT 619.200 814.050 621.000 818.400 ;
        RECT 619.200 812.400 624.600 814.050 ;
        RECT 578.850 809.100 580.050 809.250 ;
        RECT 484.950 807.450 487.050 808.050 ;
        RECT 496.950 807.450 499.050 808.050 ;
        RECT 484.950 806.550 499.050 807.450 ;
        RECT 484.950 805.950 487.050 806.550 ;
        RECT 496.950 805.950 499.050 806.550 ;
        RECT 502.950 805.950 505.050 808.050 ;
        RECT 511.950 805.950 514.050 808.050 ;
        RECT 517.950 805.950 520.050 808.050 ;
        RECT 539.100 806.100 540.900 806.850 ;
        RECT 494.100 803.100 495.900 803.850 ;
        RECT 497.850 803.100 499.050 804.900 ;
        RECT 503.100 804.150 504.900 804.900 ;
        RECT 512.100 804.150 513.900 804.900 ;
        RECT 500.100 803.100 501.900 803.850 ;
        RECT 515.100 803.100 516.900 803.850 ;
        RECT 517.950 803.100 519.150 804.900 ;
        RECT 521.100 803.100 522.900 803.850 ;
        RECT 475.950 801.450 480.000 802.050 ;
        RECT 481.950 801.450 484.050 802.050 ;
        RECT 475.950 800.550 484.050 801.450 ;
        RECT 475.950 799.950 480.000 800.550 ;
        RECT 481.950 799.950 484.050 800.550 ;
        RECT 493.950 799.950 496.050 802.050 ;
        RECT 497.850 798.900 498.900 803.100 ;
        RECT 499.950 799.950 502.050 802.050 ;
        RECT 514.950 799.950 517.050 802.050 ;
        RECT 518.100 798.900 519.150 803.100 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 520.950 799.950 523.050 802.050 ;
        RECT 535.950 799.950 538.050 802.050 ;
        RECT 542.400 800.100 543.300 808.350 ;
        RECT 596.700 808.350 600.900 810.000 ;
        RECT 623.700 809.100 624.600 812.400 ;
        RECT 640.200 811.200 642.000 818.400 ;
        RECT 655.500 812.400 657.300 818.400 ;
        RECT 661.800 815.400 663.600 818.400 ;
        RECT 638.400 810.300 642.000 811.200 ;
        RECT 553.950 805.950 556.050 808.050 ;
        RECT 559.950 807.450 562.050 808.050 ;
        RECT 564.000 807.450 568.050 808.050 ;
        RECT 559.950 806.550 568.050 807.450 ;
        RECT 559.950 805.950 562.050 806.550 ;
        RECT 564.000 805.950 568.050 806.550 ;
        RECT 571.950 805.950 574.050 808.050 ;
        RECT 577.950 807.450 580.050 808.050 ;
        RECT 592.950 807.450 595.050 808.050 ;
        RECT 577.950 806.550 595.050 807.450 ;
        RECT 577.950 805.950 580.050 806.550 ;
        RECT 592.950 805.950 595.050 806.550 ;
        RECT 554.100 804.150 555.900 804.900 ;
        RECT 551.100 803.100 552.900 803.850 ;
        RECT 557.100 803.100 558.900 803.850 ;
        RECT 550.950 799.950 553.050 802.050 ;
        RECT 556.950 799.950 559.050 802.050 ;
        RECT 425.700 789.900 432.300 790.800 ;
        RECT 425.700 789.600 426.600 789.900 ;
        RECT 424.800 783.600 426.600 789.600 ;
        RECT 430.800 789.600 432.300 789.900 ;
        RECT 430.800 783.600 432.600 789.600 ;
        RECT 442.800 783.600 444.600 795.600 ;
        RECT 445.800 794.700 453.600 795.600 ;
        RECT 445.800 783.600 447.600 794.700 ;
        RECT 451.800 783.600 453.600 794.700 ;
        RECT 461.400 794.700 469.200 795.600 ;
        RECT 461.400 783.600 463.200 794.700 ;
        RECT 467.400 783.600 469.200 794.700 ;
        RECT 470.400 783.600 472.200 795.600 ;
        RECT 482.400 789.600 483.600 798.900 ;
        RECT 497.850 795.600 499.050 798.900 ;
        RECT 517.950 795.600 519.150 798.900 ;
        RECT 536.100 798.150 537.900 798.900 ;
        RECT 533.100 797.100 534.900 797.850 ;
        RECT 541.950 796.950 547.050 799.050 ;
        RECT 482.400 783.600 484.200 789.600 ;
        RECT 497.700 783.600 499.500 795.600 ;
        RECT 517.500 783.600 519.300 795.600 ;
        RECT 532.950 793.950 535.050 796.050 ;
        RECT 542.400 790.800 543.300 795.900 ;
        RECT 560.700 795.600 561.600 804.900 ;
        RECT 572.100 804.150 573.900 804.900 ;
        RECT 575.100 803.100 576.900 803.850 ;
        RECT 577.950 803.100 579.150 804.900 ;
        RECT 581.100 803.100 582.900 803.850 ;
        RECT 574.950 799.950 577.050 802.050 ;
        RECT 578.100 798.900 579.150 803.100 ;
        RECT 580.950 799.950 583.050 802.050 ;
        RECT 596.700 800.100 597.600 808.350 ;
        RECT 599.100 806.100 600.900 806.850 ;
        RECT 616.950 805.950 619.050 808.050 ;
        RECT 622.950 805.950 625.050 808.050 ;
        RECT 638.400 806.100 639.600 810.300 ;
        RECT 655.800 809.100 657.000 812.400 ;
        RECT 661.800 811.500 663.000 815.400 ;
        RECT 657.900 810.600 663.000 811.500 ;
        RECT 675.000 811.200 676.800 818.400 ;
        RECT 691.200 814.050 693.000 818.400 ;
        RECT 712.800 815.400 714.600 818.400 ;
        RECT 691.200 812.400 696.600 814.050 ;
        RECT 657.900 809.700 659.850 810.600 ;
        RECT 675.000 810.300 678.600 811.200 ;
        RECT 658.950 809.100 659.850 809.700 ;
        RECT 643.950 807.450 646.050 808.050 ;
        RECT 655.950 807.450 658.050 808.050 ;
        RECT 643.950 806.550 658.050 807.450 ;
        RECT 643.950 805.950 646.050 806.550 ;
        RECT 655.950 805.950 658.050 806.550 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 617.100 804.150 618.900 804.900 ;
        RECT 614.100 803.100 615.900 803.850 ;
        RECT 620.100 803.100 621.900 803.850 ;
        RECT 601.950 799.950 604.050 802.050 ;
        RECT 613.950 799.950 616.050 802.050 ;
        RECT 619.950 799.950 622.050 802.050 ;
        RECT 577.950 795.600 579.150 798.900 ;
        RECT 586.950 798.450 589.050 799.050 ;
        RECT 595.950 798.450 598.050 799.050 ;
        RECT 586.950 797.550 598.050 798.450 ;
        RECT 602.100 798.150 603.900 798.900 ;
        RECT 586.950 796.950 589.050 797.550 ;
        RECT 595.950 796.950 598.050 797.550 ;
        RECT 605.100 797.100 606.900 797.850 ;
        RECT 536.700 789.900 543.300 790.800 ;
        RECT 536.700 789.600 538.200 789.900 ;
        RECT 536.400 783.600 538.200 789.600 ;
        RECT 542.400 789.600 543.300 789.900 ;
        RECT 551.400 794.700 559.200 795.600 ;
        RECT 542.400 783.600 544.200 789.600 ;
        RECT 551.400 783.600 553.200 794.700 ;
        RECT 557.400 783.600 559.200 794.700 ;
        RECT 560.400 783.600 562.200 795.600 ;
        RECT 577.500 783.600 579.300 795.600 ;
        RECT 596.700 790.800 597.600 795.900 ;
        RECT 604.950 793.950 607.050 796.050 ;
        RECT 623.700 795.600 624.600 804.900 ;
        RECT 628.950 804.450 631.050 805.050 ;
        RECT 637.950 804.450 640.050 805.050 ;
        RECT 659.100 804.900 659.850 809.100 ;
        RECT 677.400 806.100 678.600 810.300 ;
        RECT 695.700 809.100 696.600 812.400 ;
        RECT 713.400 812.100 714.600 815.400 ;
        RECT 727.200 811.200 729.000 818.400 ;
        RECT 737.400 813.300 739.200 818.400 ;
        RECT 743.400 813.300 745.200 818.400 ;
        RECT 737.400 811.950 745.200 813.300 ;
        RECT 746.400 812.400 748.200 818.400 ;
        RECT 758.400 813.300 760.200 818.400 ;
        RECT 764.400 813.300 766.200 818.400 ;
        RECT 712.950 810.450 715.050 811.050 ;
        RECT 721.950 810.450 724.050 811.050 ;
        RECT 712.950 809.550 724.050 810.450 ;
        RECT 712.950 808.950 715.050 809.550 ;
        RECT 721.950 808.950 724.050 809.550 ;
        RECT 725.400 810.300 729.000 811.200 ;
        RECT 746.400 810.300 747.600 812.400 ;
        RECT 758.400 811.950 766.200 813.300 ;
        RECT 767.400 812.400 769.200 818.400 ;
        RECT 767.400 810.300 768.600 812.400 ;
        RECT 688.950 805.950 691.050 808.050 ;
        RECT 694.950 807.450 697.050 808.050 ;
        RECT 703.950 807.450 706.050 808.050 ;
        RECT 694.950 806.550 706.050 807.450 ;
        RECT 694.950 805.950 697.050 806.550 ;
        RECT 703.950 805.950 706.050 806.550 ;
        RECT 712.950 806.100 714.300 807.900 ;
        RECT 725.400 806.100 726.600 810.300 ;
        RECT 743.850 809.250 747.600 810.300 ;
        RECT 764.850 809.250 768.600 810.300 ;
        RECT 785.100 810.000 786.900 818.400 ;
        RECT 803.100 810.000 804.900 818.400 ;
        RECT 820.200 814.050 822.000 818.400 ;
        RECT 820.200 812.400 825.600 814.050 ;
        RECT 743.850 809.100 745.050 809.250 ;
        RECT 764.850 809.100 766.050 809.250 ;
        RECT 785.100 808.350 789.300 810.000 ;
        RECT 628.950 803.550 640.050 804.450 ;
        RECT 628.950 802.950 631.050 803.550 ;
        RECT 637.950 802.950 640.050 803.550 ;
        RECT 635.100 800.100 636.900 800.850 ;
        RECT 634.950 796.950 637.050 799.050 ;
        RECT 614.400 794.700 622.200 795.600 ;
        RECT 596.700 789.900 603.300 790.800 ;
        RECT 596.700 789.600 597.600 789.900 ;
        RECT 595.800 783.600 597.600 789.600 ;
        RECT 601.800 789.600 603.300 789.900 ;
        RECT 601.800 783.600 603.600 789.600 ;
        RECT 614.400 783.600 616.200 794.700 ;
        RECT 620.400 783.600 622.200 794.700 ;
        RECT 623.400 783.600 625.200 795.600 ;
        RECT 638.400 789.600 639.600 801.900 ;
        RECT 641.100 800.100 642.900 800.850 ;
        RECT 655.800 795.600 657.000 804.900 ;
        RECT 658.950 798.300 659.850 804.900 ;
        RECT 676.950 802.950 682.050 805.050 ;
        RECT 689.100 804.150 690.900 804.900 ;
        RECT 686.100 803.100 687.900 803.850 ;
        RECT 692.100 803.100 693.900 803.850 ;
        RECT 662.100 801.150 663.900 801.900 ;
        RECT 674.100 800.100 675.900 800.850 ;
        RECT 657.900 797.400 659.850 798.300 ;
        RECT 657.900 796.500 663.600 797.400 ;
        RECT 673.950 796.950 676.050 799.050 ;
        RECT 638.400 783.600 640.200 789.600 ;
        RECT 655.500 783.600 657.300 795.600 ;
        RECT 662.400 789.600 663.600 796.500 ;
        RECT 677.400 789.600 678.600 801.900 ;
        RECT 680.100 800.100 681.900 800.850 ;
        RECT 685.950 799.950 688.050 802.050 ;
        RECT 691.950 799.950 694.050 802.050 ;
        RECT 679.950 796.800 682.050 799.050 ;
        RECT 695.700 795.600 696.600 804.900 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 713.100 801.900 714.300 806.100 ;
        RECT 736.950 805.950 739.050 808.050 ;
        RECT 742.950 807.450 745.050 808.050 ;
        RECT 747.000 807.450 751.050 808.050 ;
        RECT 742.950 806.550 751.050 807.450 ;
        RECT 742.950 805.950 745.050 806.550 ;
        RECT 747.000 805.950 751.050 806.550 ;
        RECT 757.950 805.950 760.050 808.050 ;
        RECT 763.950 807.450 766.050 808.050 ;
        RECT 778.950 807.450 781.050 808.050 ;
        RECT 763.950 806.550 781.050 807.450 ;
        RECT 763.950 805.950 766.050 806.550 ;
        RECT 778.950 805.950 781.050 806.550 ;
        RECT 785.100 806.100 786.900 806.850 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 737.100 804.150 738.900 804.900 ;
        RECT 740.100 803.100 741.900 803.850 ;
        RECT 742.950 803.100 744.150 804.900 ;
        RECT 758.100 804.150 759.900 804.900 ;
        RECT 746.100 803.100 747.900 803.850 ;
        RECT 761.100 803.100 762.900 803.850 ;
        RECT 763.950 803.100 765.150 804.900 ;
        RECT 767.100 803.100 768.900 803.850 ;
        RECT 710.100 801.150 711.900 801.900 ;
        RECT 712.950 796.650 714.300 801.900 ;
        RECT 715.950 799.950 718.050 802.050 ;
        RECT 722.100 800.100 723.900 800.850 ;
        RECT 716.100 798.150 717.900 798.900 ;
        RECT 721.950 796.950 724.050 799.050 ;
        RECT 711.600 795.600 714.300 796.650 ;
        RECT 661.800 783.600 663.600 789.600 ;
        RECT 676.800 783.600 678.600 789.600 ;
        RECT 686.400 794.700 694.200 795.600 ;
        RECT 686.400 783.600 688.200 794.700 ;
        RECT 692.400 783.600 694.200 794.700 ;
        RECT 695.400 783.600 697.200 795.600 ;
        RECT 711.600 783.600 713.400 795.600 ;
        RECT 725.400 789.600 726.600 801.900 ;
        RECT 728.100 800.100 729.900 800.850 ;
        RECT 739.950 799.950 742.050 802.050 ;
        RECT 727.950 796.950 730.050 799.050 ;
        RECT 743.100 798.900 744.150 803.100 ;
        RECT 745.950 799.950 748.050 802.050 ;
        RECT 760.950 799.950 763.050 802.050 ;
        RECT 764.100 798.900 765.150 803.100 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 766.950 799.950 769.050 802.050 ;
        RECT 781.950 799.950 784.050 802.050 ;
        RECT 788.400 800.100 789.300 808.350 ;
        RECT 800.700 808.350 804.900 810.000 ;
        RECT 824.700 809.100 825.600 812.400 ;
        RECT 800.700 800.100 801.600 808.350 ;
        RECT 803.100 806.100 804.900 806.850 ;
        RECT 817.950 805.950 820.050 808.050 ;
        RECT 823.950 805.950 826.050 808.050 ;
        RECT 802.950 802.950 805.050 805.200 ;
        RECT 818.100 804.150 819.900 804.900 ;
        RECT 815.100 803.100 816.900 803.850 ;
        RECT 821.100 803.100 822.900 803.850 ;
        RECT 805.950 799.950 808.050 802.050 ;
        RECT 814.950 799.950 817.050 802.050 ;
        RECT 820.950 799.950 823.050 802.050 ;
        RECT 742.950 795.600 744.150 798.900 ;
        RECT 763.950 795.600 765.150 798.900 ;
        RECT 782.100 798.150 783.900 798.900 ;
        RECT 787.950 798.450 790.050 799.050 ;
        RECT 792.000 798.450 796.050 799.050 ;
        RECT 779.100 797.100 780.900 797.850 ;
        RECT 787.950 797.550 796.050 798.450 ;
        RECT 787.950 796.950 790.050 797.550 ;
        RECT 792.000 796.950 796.050 797.550 ;
        RECT 799.950 796.950 802.050 799.050 ;
        RECT 806.100 798.150 807.900 798.900 ;
        RECT 809.100 797.100 810.900 797.850 ;
        RECT 725.400 783.600 727.200 789.600 ;
        RECT 742.500 783.600 744.300 795.600 ;
        RECT 763.500 783.600 765.300 795.600 ;
        RECT 778.950 793.950 781.050 796.050 ;
        RECT 788.400 790.800 789.300 795.900 ;
        RECT 782.700 789.900 789.300 790.800 ;
        RECT 782.700 789.600 784.200 789.900 ;
        RECT 782.400 783.600 784.200 789.600 ;
        RECT 788.400 789.600 789.300 789.900 ;
        RECT 800.700 790.800 801.600 795.900 ;
        RECT 808.950 793.950 811.050 796.050 ;
        RECT 824.700 795.600 825.600 804.900 ;
        RECT 815.400 794.700 823.200 795.600 ;
        RECT 800.700 789.900 807.300 790.800 ;
        RECT 800.700 789.600 801.600 789.900 ;
        RECT 788.400 783.600 790.200 789.600 ;
        RECT 799.800 783.600 801.600 789.600 ;
        RECT 805.800 789.600 807.300 789.900 ;
        RECT 805.800 783.600 807.600 789.600 ;
        RECT 815.400 783.600 817.200 794.700 ;
        RECT 821.400 783.600 823.200 794.700 ;
        RECT 824.400 783.600 826.200 795.600 ;
        RECT 11.700 767.400 13.500 779.400 ;
        RECT 26.400 773.400 28.200 779.400 ;
        RECT 11.850 764.100 13.050 767.400 ;
        RECT 26.400 764.100 27.600 773.400 ;
        RECT 40.500 767.400 42.300 779.400 ;
        RECT 58.800 767.400 60.600 779.400 ;
        RECT 61.800 768.300 63.600 779.400 ;
        RECT 67.800 768.300 69.600 779.400 ;
        RECT 77.400 773.400 79.200 779.400 ;
        RECT 77.700 773.100 79.200 773.400 ;
        RECT 83.400 773.400 85.200 779.400 ;
        RECT 98.400 773.400 100.200 779.400 ;
        RECT 83.400 773.100 84.300 773.400 ;
        RECT 77.700 772.200 84.300 773.100 ;
        RECT 98.700 773.100 100.200 773.400 ;
        RECT 104.400 773.400 106.200 779.400 ;
        RECT 116.400 773.400 118.200 779.400 ;
        RECT 131.400 773.400 133.200 779.400 ;
        RECT 104.400 773.100 105.300 773.400 ;
        RECT 98.700 772.200 105.300 773.100 ;
        RECT 61.800 767.400 69.600 768.300 ;
        RECT 40.950 764.100 42.150 767.400 ;
        RECT 7.950 760.950 10.050 763.050 ;
        RECT 11.850 759.900 12.900 764.100 ;
        RECT 13.950 760.950 16.050 763.050 ;
        RECT 25.950 760.950 31.050 763.050 ;
        RECT 37.950 760.950 40.050 763.050 ;
        RECT 41.100 759.900 42.150 764.100 ;
        RECT 43.950 760.950 46.050 763.050 ;
        RECT 8.100 759.150 9.900 759.900 ;
        RECT 11.850 758.100 13.050 759.900 ;
        RECT 14.100 759.150 15.900 759.900 ;
        RECT 17.100 758.100 18.900 758.850 ;
        RECT 23.100 758.100 24.900 758.850 ;
        RECT 10.950 754.950 13.050 757.050 ;
        RECT 16.950 754.950 19.050 757.050 ;
        RECT 10.950 753.750 12.150 753.900 ;
        RECT 8.400 752.700 12.150 753.750 ;
        RECT 8.400 750.600 9.600 752.700 ;
        RECT 22.950 751.950 25.050 757.050 ;
        RECT 7.800 744.600 9.600 750.600 ;
        RECT 10.800 749.700 18.600 751.050 ;
        RECT 10.800 744.600 12.600 749.700 ;
        RECT 16.800 744.600 18.600 749.700 ;
        RECT 26.400 747.600 27.600 759.900 ;
        RECT 38.100 759.150 39.900 759.900 ;
        RECT 35.100 758.100 36.900 758.850 ;
        RECT 40.950 758.100 42.150 759.900 ;
        RECT 44.100 759.150 45.900 759.900 ;
        RECT 59.400 758.100 60.300 767.400 ;
        RECT 73.950 766.950 76.050 769.050 ;
        RECT 83.400 767.100 84.300 772.200 ;
        RECT 94.950 766.950 97.050 769.050 ;
        RECT 104.400 767.100 105.300 772.200 ;
        RECT 74.100 765.150 75.900 765.900 ;
        RECT 77.100 764.100 78.900 764.850 ;
        RECT 82.950 763.950 85.050 766.050 ;
        RECT 95.100 765.150 96.900 765.900 ;
        RECT 98.100 764.100 99.900 764.850 ;
        RECT 103.950 763.950 106.050 766.050 ;
        RECT 112.950 763.950 115.050 766.050 ;
        RECT 61.950 760.950 64.050 763.050 ;
        RECT 67.950 760.950 70.050 763.050 ;
        RECT 76.950 760.950 79.050 763.050 ;
        RECT 62.100 759.150 63.900 759.900 ;
        RECT 68.100 759.150 69.900 759.900 ;
        RECT 65.100 758.100 66.900 758.850 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 34.950 754.950 37.050 757.050 ;
        RECT 40.950 754.950 45.900 757.050 ;
        RECT 58.950 756.450 61.050 757.050 ;
        RECT 47.550 756.000 61.050 756.450 ;
        RECT 46.950 755.550 61.050 756.000 ;
        RECT 41.850 753.750 43.050 753.900 ;
        RECT 41.850 752.700 45.600 753.750 ;
        RECT 35.400 749.700 43.200 751.050 ;
        RECT 26.400 744.600 28.200 747.600 ;
        RECT 35.400 744.600 37.200 749.700 ;
        RECT 41.400 744.600 43.200 749.700 ;
        RECT 44.400 750.600 45.600 752.700 ;
        RECT 46.950 751.950 49.050 755.550 ;
        RECT 58.950 754.950 61.050 755.550 ;
        RECT 64.950 754.950 67.050 757.050 ;
        RECT 80.100 756.150 81.900 756.900 ;
        RECT 83.400 754.650 84.300 762.900 ;
        RECT 97.950 760.950 100.050 763.200 ;
        RECT 100.950 757.950 103.050 760.200 ;
        RECT 101.100 756.150 102.900 756.900 ;
        RECT 104.400 754.650 105.300 762.900 ;
        RECT 113.100 762.150 114.900 762.900 ;
        RECT 116.400 761.100 117.600 773.400 ;
        RECT 118.950 763.950 121.050 766.050 ;
        RECT 127.950 763.950 130.050 766.050 ;
        RECT 119.100 762.150 120.900 762.900 ;
        RECT 128.100 762.150 129.900 762.900 ;
        RECT 131.400 761.100 132.600 773.400 ;
        RECT 146.400 768.600 148.200 779.400 ;
        RECT 152.400 778.500 160.200 779.400 ;
        RECT 152.400 768.600 154.200 778.500 ;
        RECT 146.400 767.700 154.200 768.600 ;
        RECT 155.400 766.500 157.200 777.600 ;
        RECT 158.400 767.400 160.200 778.500 ;
        RECT 172.800 767.400 174.600 779.400 ;
        RECT 175.800 768.300 177.600 779.400 ;
        RECT 181.800 768.300 183.600 779.400 ;
        RECT 191.400 773.400 193.200 779.400 ;
        RECT 191.700 773.100 193.200 773.400 ;
        RECT 197.400 773.400 199.200 779.400 ;
        RECT 197.400 773.100 198.300 773.400 ;
        RECT 191.700 772.200 198.300 773.100 ;
        RECT 175.800 767.400 183.600 768.300 ;
        RECT 153.150 765.600 157.200 766.500 ;
        RECT 153.150 764.100 154.050 765.600 ;
        RECT 134.100 762.150 135.900 762.900 ;
        RECT 148.950 760.800 151.050 763.050 ;
        RECT 106.950 759.450 109.050 760.050 ;
        RECT 115.950 759.450 118.050 760.050 ;
        RECT 106.950 758.550 118.050 759.450 ;
        RECT 106.950 757.950 109.050 758.550 ;
        RECT 115.950 757.950 118.050 758.550 ;
        RECT 130.950 757.950 133.050 760.050 ;
        RECT 153.150 759.900 153.900 764.100 ;
        RECT 154.950 762.450 157.050 763.050 ;
        RECT 166.950 762.450 169.050 763.050 ;
        RECT 154.950 761.550 169.050 762.450 ;
        RECT 154.950 760.950 157.050 761.550 ;
        RECT 166.950 760.950 169.050 761.550 ;
        RECT 149.250 759.150 151.050 759.900 ;
        RECT 146.250 758.100 148.050 758.850 ;
        RECT 153.150 758.100 154.050 759.900 ;
        RECT 154.950 759.150 156.750 759.900 ;
        RECT 158.100 758.100 159.900 758.850 ;
        RECT 173.400 758.100 174.300 767.400 ;
        RECT 187.950 766.950 190.050 769.050 ;
        RECT 197.400 767.100 198.300 772.200 ;
        RECT 215.700 767.400 217.500 779.400 ;
        RECT 233.700 767.400 235.500 779.400 ;
        RECT 250.800 773.400 252.600 779.400 ;
        RECT 251.700 773.100 252.600 773.400 ;
        RECT 256.800 773.400 258.600 779.400 ;
        RECT 256.800 773.100 258.300 773.400 ;
        RECT 251.700 772.200 258.300 773.100 ;
        RECT 188.100 765.150 189.900 765.900 ;
        RECT 196.950 765.450 199.050 766.050 ;
        RECT 205.950 765.450 208.050 766.050 ;
        RECT 191.100 764.100 192.900 764.850 ;
        RECT 196.950 764.550 208.050 765.450 ;
        RECT 196.950 763.950 199.050 764.550 ;
        RECT 205.950 763.950 208.050 764.550 ;
        RECT 215.850 764.100 217.050 767.400 ;
        RECT 233.850 764.100 235.050 767.400 ;
        RECT 251.700 767.100 252.600 772.200 ;
        RECT 259.950 766.950 262.050 769.050 ;
        RECT 271.800 767.400 273.600 779.400 ;
        RECT 274.800 768.300 276.600 779.400 ;
        RECT 280.800 768.300 282.600 779.400 ;
        RECT 274.800 767.400 282.600 768.300 ;
        RECT 290.400 768.300 292.200 779.400 ;
        RECT 296.400 768.300 298.200 779.400 ;
        RECT 290.400 767.400 298.200 768.300 ;
        RECT 299.400 767.400 301.200 779.400 ;
        RECT 310.800 773.400 312.600 779.400 ;
        RECT 311.700 773.100 312.600 773.400 ;
        RECT 316.800 773.400 318.600 779.400 ;
        RECT 328.800 773.400 330.600 779.400 ;
        RECT 316.800 773.100 318.300 773.400 ;
        RECT 311.700 772.200 318.300 773.100 ;
        RECT 329.700 773.100 330.600 773.400 ;
        RECT 334.800 773.400 336.600 779.400 ;
        RECT 349.800 773.400 351.600 779.400 ;
        RECT 334.800 773.100 336.300 773.400 ;
        RECT 329.700 772.200 336.300 773.100 ;
        RECT 350.700 773.100 351.600 773.400 ;
        RECT 355.800 773.400 357.600 779.400 ;
        RECT 367.800 773.400 369.600 779.400 ;
        RECT 355.800 773.100 357.300 773.400 ;
        RECT 350.700 772.200 357.300 773.100 ;
        RECT 241.950 765.450 244.050 766.050 ;
        RECT 250.950 765.450 253.050 766.050 ;
        RECT 241.950 764.550 253.050 765.450 ;
        RECT 260.100 765.150 261.900 765.900 ;
        RECT 175.950 760.950 178.050 763.050 ;
        RECT 181.950 760.950 184.050 763.050 ;
        RECT 190.950 760.950 193.050 763.050 ;
        RECT 176.100 759.150 177.900 759.900 ;
        RECT 182.100 759.150 183.900 759.900 ;
        RECT 179.100 758.100 180.900 758.850 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 59.400 750.600 60.300 753.900 ;
        RECT 80.100 753.000 84.300 754.650 ;
        RECT 101.100 753.000 105.300 754.650 ;
        RECT 44.400 744.600 46.200 750.600 ;
        RECT 59.400 748.950 64.800 750.600 ;
        RECT 63.000 744.600 64.800 748.950 ;
        RECT 80.100 744.600 81.900 753.000 ;
        RECT 101.100 744.600 102.900 753.000 ;
        RECT 116.400 752.700 117.600 756.900 ;
        RECT 131.400 752.700 132.600 756.900 ;
        RECT 145.950 754.950 148.050 757.050 ;
        RECT 151.950 754.950 154.050 757.050 ;
        RECT 157.950 756.450 160.050 757.050 ;
        RECT 162.000 756.450 166.050 757.050 ;
        RECT 157.950 755.550 166.050 756.450 ;
        RECT 157.950 754.950 160.050 755.550 ;
        RECT 162.000 754.950 166.050 755.550 ;
        RECT 172.950 754.950 175.050 757.050 ;
        RECT 178.950 754.950 181.050 757.050 ;
        RECT 194.100 756.150 195.900 756.900 ;
        RECT 197.400 754.650 198.300 762.900 ;
        RECT 211.950 760.950 214.050 763.050 ;
        RECT 215.850 759.900 216.900 764.100 ;
        RECT 217.950 760.950 220.050 763.050 ;
        RECT 229.950 760.950 232.050 763.200 ;
        RECT 233.850 759.900 234.900 764.100 ;
        RECT 241.950 763.950 244.050 764.550 ;
        RECT 250.950 763.950 253.050 764.550 ;
        RECT 257.100 764.100 258.900 764.850 ;
        RECT 235.950 760.950 238.050 763.050 ;
        RECT 212.100 759.150 213.900 759.900 ;
        RECT 215.850 758.100 217.050 759.900 ;
        RECT 218.100 759.150 219.900 759.900 ;
        RECT 230.100 759.150 231.900 759.900 ;
        RECT 221.100 758.100 222.900 758.850 ;
        RECT 233.850 758.100 235.050 759.900 ;
        RECT 236.100 759.150 237.900 759.900 ;
        RECT 239.100 758.100 240.900 758.850 ;
        RECT 199.950 756.450 202.050 757.050 ;
        RECT 214.950 756.450 217.050 757.050 ;
        RECT 199.950 755.550 217.050 756.450 ;
        RECT 199.950 754.950 202.050 755.550 ;
        RECT 214.950 754.950 217.050 755.550 ;
        RECT 220.950 754.950 223.050 757.050 ;
        RECT 229.950 754.950 235.050 757.050 ;
        RECT 238.950 754.950 241.050 757.050 ;
        RECT 116.400 751.800 120.000 752.700 ;
        RECT 131.400 751.800 135.000 752.700 ;
        RECT 118.200 744.600 120.000 751.800 ;
        RECT 133.200 744.600 135.000 751.800 ;
        RECT 151.950 750.600 153.000 753.900 ;
        RECT 151.200 744.600 153.000 750.600 ;
        RECT 173.400 750.600 174.300 753.900 ;
        RECT 194.100 753.000 198.300 754.650 ;
        RECT 251.700 754.650 252.600 762.900 ;
        RECT 256.950 760.950 259.050 763.050 ;
        RECT 253.950 757.950 256.050 760.050 ;
        RECT 272.400 758.100 273.300 767.400 ;
        RECT 274.950 760.950 277.050 763.050 ;
        RECT 280.950 760.950 283.050 763.050 ;
        RECT 289.950 760.950 292.050 763.050 ;
        RECT 295.950 760.950 298.050 763.050 ;
        RECT 275.100 759.150 276.900 759.900 ;
        RECT 281.100 759.150 282.900 759.900 ;
        RECT 290.100 759.150 291.900 759.900 ;
        RECT 296.100 759.150 297.900 759.900 ;
        RECT 278.100 758.100 279.900 758.850 ;
        RECT 293.100 758.100 294.900 758.850 ;
        RECT 299.700 758.100 300.600 767.400 ;
        RECT 311.700 767.100 312.600 772.200 ;
        RECT 319.950 766.950 322.050 769.050 ;
        RECT 329.700 767.100 330.600 772.200 ;
        RECT 337.950 766.950 340.050 769.050 ;
        RECT 350.700 767.100 351.600 772.200 ;
        RECT 358.950 766.950 361.050 769.050 ;
        RECT 304.950 765.450 309.000 766.050 ;
        RECT 310.950 765.450 313.050 766.050 ;
        RECT 304.950 764.550 313.050 765.450 ;
        RECT 320.100 765.150 321.900 765.900 ;
        RECT 304.950 763.950 309.000 764.550 ;
        RECT 310.950 763.950 313.050 764.550 ;
        RECT 317.100 764.100 318.900 764.850 ;
        RECT 325.950 763.950 331.050 766.050 ;
        RECT 338.100 765.150 339.900 765.900 ;
        RECT 343.950 765.450 348.000 766.050 ;
        RECT 349.950 765.450 352.050 766.050 ;
        RECT 335.100 764.100 336.900 764.850 ;
        RECT 343.950 764.550 352.050 765.450 ;
        RECT 359.100 765.150 360.900 765.900 ;
        RECT 343.950 763.950 348.000 764.550 ;
        RECT 349.950 763.950 352.050 764.550 ;
        RECT 356.100 764.100 357.900 764.850 ;
        RECT 368.400 764.100 369.600 773.400 ;
        RECT 382.800 767.400 384.600 779.400 ;
        RECT 385.800 768.300 387.600 779.400 ;
        RECT 391.800 768.300 393.600 779.400 ;
        RECT 400.800 773.400 402.600 779.400 ;
        RECT 385.800 767.400 393.600 768.300 ;
        RECT 401.700 773.100 402.600 773.400 ;
        RECT 406.800 773.400 408.600 779.400 ;
        RECT 419.400 773.400 421.200 779.400 ;
        RECT 433.800 778.500 441.600 779.400 ;
        RECT 406.800 773.100 408.300 773.400 ;
        RECT 401.700 772.200 408.300 773.100 ;
        RECT 254.100 756.150 255.900 756.900 ;
        RECT 265.950 756.450 270.000 757.050 ;
        RECT 271.950 756.450 274.050 757.050 ;
        RECT 265.950 755.550 274.050 756.450 ;
        RECT 265.950 754.950 270.000 755.550 ;
        RECT 271.950 754.950 274.050 755.550 ;
        RECT 277.950 754.950 280.050 757.050 ;
        RECT 292.950 754.950 295.050 757.050 ;
        RECT 298.950 754.950 304.050 757.050 ;
        RECT 311.700 754.650 312.600 762.900 ;
        RECT 316.950 760.950 319.050 763.200 ;
        RECT 313.950 757.950 316.050 760.050 ;
        RECT 314.100 756.150 315.900 756.900 ;
        RECT 329.700 754.650 330.600 762.900 ;
        RECT 334.950 760.950 337.050 763.200 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 332.100 756.150 333.900 756.900 ;
        RECT 337.950 756.450 340.050 757.050 ;
        RECT 346.950 756.450 349.050 757.050 ;
        RECT 337.950 755.550 349.050 756.450 ;
        RECT 337.950 754.950 340.050 755.550 ;
        RECT 346.950 754.950 349.050 755.550 ;
        RECT 350.700 754.650 351.600 762.900 ;
        RECT 355.950 760.950 358.050 763.050 ;
        RECT 364.950 760.950 370.050 763.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 353.100 756.150 354.900 756.900 ;
        RECT 214.950 753.750 216.150 753.900 ;
        RECT 232.950 753.750 234.150 753.900 ;
        RECT 173.400 748.950 178.800 750.600 ;
        RECT 177.000 744.600 178.800 748.950 ;
        RECT 194.100 744.600 195.900 753.000 ;
        RECT 212.400 752.700 216.150 753.750 ;
        RECT 230.400 752.700 234.150 753.750 ;
        RECT 251.700 753.000 255.900 754.650 ;
        RECT 212.400 750.600 213.600 752.700 ;
        RECT 211.800 744.600 213.600 750.600 ;
        RECT 214.800 749.700 222.600 751.050 ;
        RECT 230.400 750.600 231.600 752.700 ;
        RECT 214.800 744.600 216.600 749.700 ;
        RECT 220.800 744.600 222.600 749.700 ;
        RECT 229.800 744.600 231.600 750.600 ;
        RECT 232.800 749.700 240.600 751.050 ;
        RECT 232.800 744.600 234.600 749.700 ;
        RECT 238.800 744.600 240.600 749.700 ;
        RECT 254.100 744.600 255.900 753.000 ;
        RECT 272.400 750.600 273.300 753.900 ;
        RECT 299.700 750.600 300.600 753.900 ;
        RECT 311.700 753.000 315.900 754.650 ;
        RECT 329.700 753.000 333.900 754.650 ;
        RECT 350.700 753.000 354.900 754.650 ;
        RECT 272.400 748.950 277.800 750.600 ;
        RECT 276.000 744.600 277.800 748.950 ;
        RECT 295.200 748.950 300.600 750.600 ;
        RECT 295.200 744.600 297.000 748.950 ;
        RECT 314.100 744.600 315.900 753.000 ;
        RECT 332.100 744.600 333.900 753.000 ;
        RECT 353.100 744.600 354.900 753.000 ;
        RECT 368.400 747.600 369.600 759.900 ;
        RECT 371.100 758.100 372.900 758.850 ;
        RECT 383.400 758.100 384.300 767.400 ;
        RECT 401.700 767.100 402.600 772.200 ;
        RECT 409.950 766.950 412.050 769.050 ;
        RECT 397.950 763.950 403.050 766.050 ;
        RECT 410.100 765.150 411.900 765.900 ;
        RECT 407.100 764.100 408.900 764.850 ;
        RECT 419.400 764.100 420.600 773.400 ;
        RECT 433.800 767.400 435.600 778.500 ;
        RECT 436.800 766.500 438.600 777.600 ;
        RECT 439.800 768.600 441.600 778.500 ;
        RECT 445.800 768.600 447.600 779.400 ;
        RECT 439.800 767.700 447.600 768.600 ;
        RECT 455.400 773.400 457.200 779.400 ;
        RECT 436.800 765.600 440.850 766.500 ;
        RECT 439.950 764.100 440.850 765.600 ;
        RECT 385.950 760.950 388.050 763.200 ;
        RECT 391.950 760.950 394.050 763.050 ;
        RECT 386.100 759.150 387.900 759.900 ;
        RECT 392.100 759.150 393.900 759.900 ;
        RECT 389.100 758.100 390.900 758.850 ;
        RECT 370.950 754.950 373.050 757.200 ;
        RECT 382.950 756.450 385.050 757.050 ;
        RECT 377.550 755.550 385.050 756.450 ;
        RECT 370.950 750.450 373.050 751.050 ;
        RECT 377.550 750.450 378.450 755.550 ;
        RECT 382.950 754.950 385.050 755.550 ;
        RECT 388.950 754.950 391.050 757.050 ;
        RECT 401.700 754.650 402.600 762.900 ;
        RECT 406.950 760.950 409.050 763.050 ;
        RECT 409.950 762.450 412.050 763.050 ;
        RECT 418.950 762.450 421.050 763.050 ;
        RECT 409.950 761.550 421.050 762.450 ;
        RECT 409.950 760.950 412.050 761.550 ;
        RECT 418.950 760.950 421.050 761.550 ;
        RECT 436.950 760.950 439.050 763.050 ;
        RECT 403.950 757.950 406.050 760.050 ;
        RECT 440.100 759.900 440.850 764.100 ;
        RECT 448.950 763.950 454.050 766.050 ;
        RECT 442.950 760.950 445.050 763.050 ;
        RECT 452.100 762.150 453.900 762.900 ;
        RECT 455.400 761.100 456.600 773.400 ;
        RECT 472.500 767.400 474.300 779.400 ;
        RECT 487.800 773.400 489.600 779.400 ;
        RECT 488.700 773.100 489.600 773.400 ;
        RECT 493.800 773.400 495.600 779.400 ;
        RECT 493.800 773.100 495.300 773.400 ;
        RECT 488.700 772.200 495.300 773.100 ;
        RECT 457.950 763.950 460.050 766.050 ;
        RECT 472.950 764.100 474.150 767.400 ;
        RECT 488.700 767.100 489.600 772.200 ;
        RECT 496.950 766.950 499.050 769.050 ;
        RECT 505.800 767.400 507.600 779.400 ;
        RECT 508.800 768.300 510.600 779.400 ;
        RECT 514.800 768.300 516.600 779.400 ;
        RECT 527.400 773.400 529.200 779.400 ;
        RECT 527.700 773.100 529.200 773.400 ;
        RECT 533.400 773.400 535.200 779.400 ;
        RECT 550.800 773.400 552.600 779.400 ;
        RECT 533.400 773.100 534.300 773.400 ;
        RECT 527.700 772.200 534.300 773.100 ;
        RECT 508.800 767.400 516.600 768.300 ;
        RECT 458.100 762.150 459.900 762.900 ;
        RECT 469.950 760.950 472.050 763.050 ;
        RECT 454.950 759.900 459.450 760.050 ;
        RECT 473.100 759.900 474.150 764.100 ;
        RECT 484.950 763.950 490.050 766.050 ;
        RECT 497.100 765.150 498.900 765.900 ;
        RECT 494.100 764.100 495.900 764.850 ;
        RECT 475.950 760.950 478.050 763.050 ;
        RECT 416.100 758.100 417.900 758.850 ;
        RECT 404.100 756.150 405.900 756.900 ;
        RECT 415.950 754.950 418.050 757.050 ;
        RECT 370.950 749.550 378.450 750.450 ;
        RECT 383.400 750.600 384.300 753.900 ;
        RECT 401.700 753.000 405.900 754.650 ;
        RECT 370.950 748.950 373.050 749.550 ;
        RECT 383.400 748.950 388.800 750.600 ;
        RECT 367.800 744.600 369.600 747.600 ;
        RECT 387.000 744.600 388.800 748.950 ;
        RECT 404.100 744.600 405.900 753.000 ;
        RECT 419.400 747.600 420.600 759.900 ;
        RECT 437.250 759.150 439.050 759.900 ;
        RECT 434.100 758.100 435.900 758.850 ;
        RECT 439.950 758.100 440.850 759.900 ;
        RECT 442.950 759.150 444.750 759.900 ;
        RECT 445.950 758.100 447.750 758.850 ;
        RECT 454.950 757.950 460.050 759.900 ;
        RECT 470.100 759.150 471.900 759.900 ;
        RECT 467.100 758.100 468.900 758.850 ;
        RECT 472.950 758.100 474.150 759.900 ;
        RECT 476.100 759.150 477.900 759.900 ;
        RECT 457.950 757.800 460.050 757.950 ;
        RECT 433.950 754.950 436.050 757.050 ;
        RECT 439.950 754.950 442.050 757.050 ;
        RECT 445.950 754.950 448.050 757.050 ;
        RECT 441.000 750.600 442.050 753.900 ;
        RECT 455.400 752.700 456.600 756.900 ;
        RECT 466.950 754.950 469.050 757.050 ;
        RECT 472.950 756.450 475.050 757.050 ;
        RECT 484.950 756.450 487.050 757.050 ;
        RECT 472.950 755.550 487.050 756.450 ;
        RECT 472.950 754.950 475.050 755.550 ;
        RECT 484.950 754.950 487.050 755.550 ;
        RECT 488.700 754.650 489.600 762.900 ;
        RECT 493.950 760.950 496.050 763.050 ;
        RECT 490.950 757.950 493.050 760.050 ;
        RECT 506.400 758.100 507.300 767.400 ;
        RECT 523.950 766.950 526.050 769.050 ;
        RECT 533.400 767.100 534.300 772.200 ;
        RECT 524.100 765.150 525.900 765.900 ;
        RECT 532.950 765.450 535.050 766.050 ;
        RECT 537.000 765.450 541.050 766.050 ;
        RECT 527.100 764.100 528.900 764.850 ;
        RECT 532.950 764.550 541.050 765.450 ;
        RECT 532.950 763.950 535.050 764.550 ;
        RECT 537.000 763.950 541.050 764.550 ;
        RECT 547.950 763.950 550.050 766.050 ;
        RECT 508.950 760.950 511.050 763.050 ;
        RECT 514.950 760.950 517.050 763.050 ;
        RECT 526.950 760.950 529.050 763.050 ;
        RECT 509.100 759.150 510.900 759.900 ;
        RECT 515.100 759.150 516.900 759.900 ;
        RECT 512.100 758.100 513.900 758.850 ;
        RECT 529.950 757.950 532.050 760.050 ;
        RECT 491.100 756.150 492.900 756.900 ;
        RECT 499.950 756.450 504.000 757.050 ;
        RECT 505.950 756.450 508.050 757.050 ;
        RECT 499.950 755.550 508.050 756.450 ;
        RECT 499.950 754.950 504.000 755.550 ;
        RECT 505.950 754.950 508.050 755.550 ;
        RECT 511.950 754.950 514.050 757.050 ;
        RECT 530.100 756.150 531.900 756.900 ;
        RECT 533.400 754.650 534.300 762.900 ;
        RECT 548.100 762.150 549.900 762.900 ;
        RECT 551.400 761.100 552.600 773.400 ;
        RECT 566.700 767.400 568.500 779.400 ;
        RECT 581.400 773.400 583.200 779.400 ;
        RECT 553.950 763.950 556.050 766.050 ;
        RECT 566.850 764.100 568.050 767.400 ;
        RECT 581.400 764.100 582.600 773.400 ;
        RECT 590.400 768.600 592.200 779.400 ;
        RECT 596.400 778.500 604.200 779.400 ;
        RECT 596.400 768.600 598.200 778.500 ;
        RECT 590.400 767.700 598.200 768.600 ;
        RECT 599.400 766.500 601.200 777.600 ;
        RECT 602.400 767.400 604.200 778.500 ;
        RECT 613.800 773.400 615.600 779.400 ;
        RECT 631.800 773.400 633.600 779.400 ;
        RECT 646.800 773.400 648.600 779.400 ;
        RECT 597.150 765.600 601.200 766.500 ;
        RECT 597.150 764.100 598.050 765.600 ;
        RECT 614.400 764.100 615.600 773.400 ;
        RECT 554.100 762.150 555.900 762.900 ;
        RECT 562.950 760.950 565.050 763.050 ;
        RECT 550.950 759.450 553.050 760.050 ;
        RECT 566.850 759.900 567.900 764.100 ;
        RECT 568.950 760.950 571.050 763.050 ;
        RECT 580.950 762.450 583.050 763.050 ;
        RECT 585.000 762.450 589.050 763.050 ;
        RECT 580.950 761.550 589.050 762.450 ;
        RECT 580.950 760.950 583.050 761.550 ;
        RECT 585.000 760.950 589.050 761.550 ;
        RECT 592.950 760.950 595.050 763.050 ;
        RECT 597.150 759.900 597.900 764.100 ;
        RECT 628.950 763.800 631.050 766.050 ;
        RECT 598.950 760.950 601.050 763.050 ;
        RECT 604.950 762.450 607.050 763.050 ;
        RECT 613.950 762.450 616.050 763.050 ;
        RECT 604.950 761.550 616.050 762.450 ;
        RECT 629.100 762.150 630.900 762.900 ;
        RECT 604.950 760.950 607.050 761.550 ;
        RECT 613.950 760.950 616.050 761.550 ;
        RECT 632.400 761.100 633.600 773.400 ;
        RECT 634.950 763.950 637.050 766.050 ;
        RECT 643.950 763.950 646.050 766.050 ;
        RECT 635.100 762.150 636.900 762.900 ;
        RECT 644.100 762.150 645.900 762.900 ;
        RECT 647.400 761.100 648.600 773.400 ;
        RECT 663.600 767.400 665.400 779.400 ;
        RECT 662.700 766.350 665.400 767.400 ;
        RECT 677.400 773.400 679.200 779.400 ;
        RECT 649.950 763.950 652.050 766.050 ;
        RECT 659.100 764.100 660.900 764.850 ;
        RECT 650.100 762.150 651.900 762.900 ;
        RECT 658.950 760.950 661.050 763.050 ;
        RECT 662.700 761.100 664.050 766.350 ;
        RECT 673.950 763.950 676.050 766.050 ;
        RECT 674.100 762.150 675.900 762.900 ;
        RECT 665.100 761.100 666.900 761.850 ;
        RECT 677.400 761.100 678.600 773.400 ;
        RECT 698.700 767.400 700.500 779.400 ;
        RECT 715.500 767.400 717.300 779.400 ;
        RECT 731.400 768.300 733.200 779.400 ;
        RECT 737.400 768.300 739.200 779.400 ;
        RECT 731.400 767.400 739.200 768.300 ;
        RECT 740.400 767.400 742.200 779.400 ;
        RECT 757.500 767.400 759.300 779.400 ;
        RECT 775.800 773.400 777.600 779.400 ;
        RECT 776.700 773.100 777.600 773.400 ;
        RECT 781.800 773.400 783.600 779.400 ;
        RECT 781.800 773.100 783.300 773.400 ;
        RECT 776.700 772.200 783.300 773.100 ;
        RECT 679.950 763.950 682.050 766.050 ;
        RECT 698.850 764.100 700.050 767.400 ;
        RECT 715.950 764.100 717.150 767.400 ;
        RECT 680.100 762.150 681.900 762.900 ;
        RECT 550.950 759.000 558.450 759.450 ;
        RECT 563.100 759.150 564.900 759.900 ;
        RECT 550.950 758.550 559.050 759.000 ;
        RECT 550.950 757.950 553.050 758.550 ;
        RECT 473.850 753.750 475.050 753.900 ;
        RECT 473.850 752.700 477.600 753.750 ;
        RECT 488.700 753.000 492.900 754.650 ;
        RECT 455.400 751.800 459.000 752.700 ;
        RECT 419.400 744.600 421.200 747.600 ;
        RECT 441.000 744.600 442.800 750.600 ;
        RECT 457.200 744.600 459.000 751.800 ;
        RECT 467.400 749.700 475.200 751.050 ;
        RECT 467.400 744.600 469.200 749.700 ;
        RECT 473.400 744.600 475.200 749.700 ;
        RECT 476.400 750.600 477.600 752.700 ;
        RECT 476.400 744.600 478.200 750.600 ;
        RECT 491.100 744.600 492.900 753.000 ;
        RECT 506.400 750.600 507.300 753.900 ;
        RECT 530.100 753.000 534.300 754.650 ;
        RECT 506.400 748.950 511.800 750.600 ;
        RECT 510.000 744.600 511.800 748.950 ;
        RECT 530.100 744.600 531.900 753.000 ;
        RECT 551.400 752.700 552.600 756.900 ;
        RECT 556.950 754.950 559.050 758.550 ;
        RECT 566.850 758.100 568.050 759.900 ;
        RECT 569.100 759.150 570.900 759.900 ;
        RECT 572.100 758.100 573.900 758.850 ;
        RECT 578.100 758.100 579.900 758.850 ;
        RECT 565.950 754.950 568.050 757.050 ;
        RECT 571.950 754.950 574.050 757.050 ;
        RECT 577.950 754.950 580.050 757.050 ;
        RECT 565.950 753.750 567.150 753.900 ;
        RECT 549.000 751.800 552.600 752.700 ;
        RECT 563.400 752.700 567.150 753.750 ;
        RECT 549.000 744.600 550.800 751.800 ;
        RECT 563.400 750.600 564.600 752.700 ;
        RECT 562.800 744.600 564.600 750.600 ;
        RECT 565.800 749.700 573.600 751.050 ;
        RECT 565.800 744.600 567.600 749.700 ;
        RECT 571.800 744.600 573.600 749.700 ;
        RECT 581.400 747.600 582.600 759.900 ;
        RECT 593.250 759.150 595.050 759.900 ;
        RECT 590.250 758.100 592.050 758.850 ;
        RECT 597.150 758.100 598.050 759.900 ;
        RECT 598.950 759.150 600.750 759.900 ;
        RECT 602.100 758.100 603.900 758.850 ;
        RECT 589.950 754.950 592.050 757.050 ;
        RECT 595.950 754.950 598.050 757.050 ;
        RECT 601.950 756.450 604.050 757.050 ;
        RECT 610.950 756.450 613.050 757.050 ;
        RECT 601.950 755.550 613.050 756.450 ;
        RECT 601.950 754.950 604.050 755.550 ;
        RECT 610.950 754.950 613.050 755.550 ;
        RECT 595.950 750.600 597.000 753.900 ;
        RECT 581.400 744.600 583.200 747.600 ;
        RECT 595.200 744.600 597.000 750.600 ;
        RECT 614.400 747.600 615.600 759.900 ;
        RECT 631.950 759.450 634.050 760.050 ;
        RECT 640.950 759.450 643.050 760.050 ;
        RECT 617.100 758.100 618.900 758.850 ;
        RECT 631.950 758.550 643.050 759.450 ;
        RECT 631.950 757.950 634.050 758.550 ;
        RECT 640.950 757.950 643.050 758.550 ;
        RECT 646.950 759.450 649.050 760.050 ;
        RECT 651.000 759.450 655.050 760.050 ;
        RECT 646.950 758.550 655.050 759.450 ;
        RECT 646.950 757.950 649.050 758.550 ;
        RECT 651.000 757.950 655.050 758.550 ;
        RECT 616.950 754.950 619.050 757.050 ;
        RECT 662.700 756.900 663.900 761.100 ;
        RECT 694.950 760.950 697.050 763.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 676.950 759.450 679.050 760.050 ;
        RECT 681.000 759.450 685.050 760.050 ;
        RECT 698.850 759.900 699.900 764.100 ;
        RECT 700.950 760.950 703.050 763.050 ;
        RECT 712.950 760.950 715.050 763.050 ;
        RECT 716.100 759.900 717.150 764.100 ;
        RECT 718.950 760.950 721.050 763.050 ;
        RECT 730.950 760.950 733.050 763.050 ;
        RECT 736.950 760.950 739.050 763.050 ;
        RECT 676.950 758.550 685.050 759.450 ;
        RECT 695.100 759.150 696.900 759.900 ;
        RECT 676.950 757.950 679.050 758.550 ;
        RECT 681.000 757.950 685.050 758.550 ;
        RECT 698.850 758.100 700.050 759.900 ;
        RECT 701.100 759.150 702.900 759.900 ;
        RECT 713.100 759.150 714.900 759.900 ;
        RECT 704.100 758.100 705.900 758.850 ;
        RECT 710.100 758.100 711.900 758.850 ;
        RECT 715.950 758.100 717.150 759.900 ;
        RECT 719.100 759.150 720.900 759.900 ;
        RECT 731.100 759.150 732.900 759.900 ;
        RECT 737.100 759.150 738.900 759.900 ;
        RECT 734.100 758.100 735.900 758.850 ;
        RECT 740.700 758.100 741.600 767.400 ;
        RECT 757.950 764.100 759.150 767.400 ;
        RECT 776.700 767.100 777.600 772.200 ;
        RECT 784.950 766.800 787.050 769.050 ;
        RECT 794.400 768.300 796.200 779.400 ;
        RECT 800.400 768.300 802.200 779.400 ;
        RECT 794.400 767.400 802.200 768.300 ;
        RECT 803.400 767.400 805.200 779.400 ;
        RECT 820.500 767.400 822.300 779.400 ;
        RECT 754.950 760.950 757.050 763.050 ;
        RECT 758.100 759.900 759.150 764.100 ;
        RECT 775.950 763.950 778.050 766.050 ;
        RECT 785.100 765.150 786.900 765.900 ;
        RECT 782.100 764.100 783.900 764.850 ;
        RECT 760.950 760.950 763.050 763.050 ;
        RECT 755.100 759.150 756.900 759.900 ;
        RECT 752.100 758.100 753.900 758.850 ;
        RECT 757.950 758.100 759.150 759.900 ;
        RECT 761.100 759.150 762.900 759.900 ;
        RECT 632.400 752.700 633.600 756.900 ;
        RECT 647.400 752.700 648.600 756.900 ;
        RECT 662.700 755.100 664.050 756.900 ;
        RECT 613.800 744.600 615.600 747.600 ;
        RECT 630.000 751.800 633.600 752.700 ;
        RECT 645.000 751.800 648.600 752.700 ;
        RECT 661.950 753.450 664.050 754.050 ;
        RECT 673.950 753.450 676.050 754.050 ;
        RECT 661.950 752.550 676.050 753.450 ;
        RECT 661.950 751.950 664.050 752.550 ;
        RECT 673.950 751.950 676.050 752.550 ;
        RECT 677.400 752.700 678.600 756.900 ;
        RECT 697.950 754.950 700.050 757.050 ;
        RECT 703.950 754.950 706.050 757.050 ;
        RECT 709.950 754.950 712.050 757.050 ;
        RECT 715.950 756.450 718.050 757.050 ;
        RECT 727.950 756.450 730.050 757.050 ;
        RECT 715.950 755.550 730.050 756.450 ;
        RECT 715.950 754.950 718.050 755.550 ;
        RECT 727.950 754.950 730.050 755.550 ;
        RECT 733.950 754.950 736.050 757.050 ;
        RECT 739.950 754.950 745.050 757.050 ;
        RECT 751.950 754.950 754.050 757.050 ;
        RECT 757.950 754.950 760.050 757.050 ;
        RECT 776.700 754.650 777.600 762.900 ;
        RECT 781.950 760.950 784.050 763.050 ;
        RECT 793.950 760.950 796.050 763.050 ;
        RECT 799.950 760.950 802.050 763.050 ;
        RECT 778.950 757.800 781.050 760.050 ;
        RECT 794.100 759.150 795.900 759.900 ;
        RECT 800.100 759.150 801.900 759.900 ;
        RECT 797.100 758.100 798.900 758.850 ;
        RECT 803.700 758.100 804.600 767.400 ;
        RECT 820.950 764.100 822.150 767.400 ;
        RECT 817.950 760.950 820.050 763.050 ;
        RECT 821.100 759.900 822.150 764.100 ;
        RECT 823.950 760.950 826.050 763.050 ;
        RECT 818.100 759.150 819.900 759.900 ;
        RECT 815.100 758.100 816.900 758.850 ;
        RECT 820.950 758.100 822.150 759.900 ;
        RECT 824.100 759.150 825.900 759.900 ;
        RECT 779.100 756.150 780.900 756.900 ;
        RECT 796.950 754.950 799.050 757.050 ;
        RECT 802.950 754.950 807.900 757.050 ;
        RECT 808.950 756.450 813.000 757.050 ;
        RECT 814.950 756.450 817.050 757.050 ;
        RECT 808.950 755.550 817.050 756.450 ;
        RECT 808.950 754.950 813.000 755.550 ;
        RECT 814.950 754.950 817.050 755.550 ;
        RECT 820.950 754.950 823.050 757.050 ;
        RECT 697.950 753.750 699.150 753.900 ;
        RECT 695.400 752.700 699.150 753.750 ;
        RECT 716.850 753.750 718.050 753.900 ;
        RECT 716.850 752.700 720.600 753.750 ;
        RECT 677.400 751.800 681.000 752.700 ;
        RECT 630.000 744.600 631.800 751.800 ;
        RECT 645.000 744.600 646.800 751.800 ;
        RECT 662.400 747.600 663.600 750.900 ;
        RECT 662.400 744.600 664.200 747.600 ;
        RECT 679.200 744.600 681.000 751.800 ;
        RECT 695.400 750.600 696.600 752.700 ;
        RECT 694.800 744.600 696.600 750.600 ;
        RECT 697.800 749.700 705.600 751.050 ;
        RECT 697.800 744.600 699.600 749.700 ;
        RECT 703.800 744.600 705.600 749.700 ;
        RECT 710.400 749.700 718.200 751.050 ;
        RECT 710.400 744.600 712.200 749.700 ;
        RECT 716.400 744.600 718.200 749.700 ;
        RECT 719.400 750.600 720.600 752.700 ;
        RECT 740.700 750.600 741.600 753.900 ;
        RECT 758.850 753.750 760.050 753.900 ;
        RECT 758.850 752.700 762.600 753.750 ;
        RECT 776.700 753.000 780.900 754.650 ;
        RECT 719.400 744.600 721.200 750.600 ;
        RECT 736.200 748.950 741.600 750.600 ;
        RECT 752.400 749.700 760.200 751.050 ;
        RECT 736.200 744.600 738.000 748.950 ;
        RECT 752.400 744.600 754.200 749.700 ;
        RECT 758.400 744.600 760.200 749.700 ;
        RECT 761.400 750.600 762.600 752.700 ;
        RECT 761.400 744.600 763.200 750.600 ;
        RECT 779.100 744.600 780.900 753.000 ;
        RECT 803.700 750.600 804.600 753.900 ;
        RECT 821.850 753.750 823.050 753.900 ;
        RECT 821.850 752.700 825.600 753.750 ;
        RECT 799.200 748.950 804.600 750.600 ;
        RECT 815.400 749.700 823.200 751.050 ;
        RECT 799.200 744.600 801.000 748.950 ;
        RECT 815.400 744.600 817.200 749.700 ;
        RECT 821.400 744.600 823.200 749.700 ;
        RECT 824.400 750.600 825.600 752.700 ;
        RECT 824.400 744.600 826.200 750.600 ;
        RECT 14.100 732.000 15.900 740.400 ;
        RECT 34.200 736.050 36.000 740.400 ;
        RECT 34.200 734.400 39.600 736.050 ;
        RECT 11.700 730.350 15.900 732.000 ;
        RECT 38.700 731.100 39.600 734.400 ;
        RECT 56.100 732.000 57.900 740.400 ;
        RECT 77.100 732.000 78.900 740.400 ;
        RECT 97.200 736.050 99.000 740.400 ;
        RECT 97.200 734.400 102.600 736.050 ;
        RECT 112.800 734.400 114.600 740.400 ;
        RECT 53.700 730.350 57.900 732.000 ;
        RECT 74.700 730.350 78.900 732.000 ;
        RECT 11.700 722.100 12.600 730.350 ;
        RECT 19.950 729.450 22.050 730.200 ;
        RECT 31.950 729.450 34.050 730.050 ;
        RECT 14.100 728.100 15.900 728.850 ;
        RECT 19.950 728.550 34.050 729.450 ;
        RECT 19.950 728.100 22.050 728.550 ;
        RECT 31.950 727.950 34.050 728.550 ;
        RECT 37.950 729.450 40.050 730.050 ;
        RECT 46.950 729.450 49.050 730.050 ;
        RECT 37.950 728.550 49.050 729.450 ;
        RECT 37.950 727.950 40.050 728.550 ;
        RECT 46.950 727.950 49.050 728.550 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 32.100 726.150 33.900 726.900 ;
        RECT 29.100 725.100 30.900 725.850 ;
        RECT 35.100 725.100 36.900 725.850 ;
        RECT 16.950 721.950 19.050 724.050 ;
        RECT 25.950 721.950 31.050 724.050 ;
        RECT 34.950 721.950 37.050 724.050 ;
        RECT 10.950 718.950 13.050 721.050 ;
        RECT 17.100 720.150 18.900 720.900 ;
        RECT 20.100 719.100 21.900 719.850 ;
        RECT 11.700 712.800 12.600 717.900 ;
        RECT 19.950 715.950 22.050 718.050 ;
        RECT 38.700 717.600 39.600 726.900 ;
        RECT 53.700 722.100 54.600 730.350 ;
        RECT 56.100 728.100 57.900 728.850 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 58.950 721.950 61.050 724.050 ;
        RECT 74.700 722.100 75.600 730.350 ;
        RECT 82.950 729.450 85.050 730.050 ;
        RECT 94.950 729.450 97.050 733.050 ;
        RECT 101.700 731.100 102.600 734.400 ;
        RECT 113.400 732.300 114.600 734.400 ;
        RECT 115.800 735.300 117.600 740.400 ;
        RECT 121.800 735.300 123.600 740.400 ;
        RECT 132.300 736.200 134.100 740.400 ;
        RECT 115.800 733.950 123.600 735.300 ;
        RECT 132.150 734.400 134.100 736.200 ;
        RECT 113.400 731.250 117.150 732.300 ;
        RECT 115.950 731.100 117.150 731.250 ;
        RECT 132.150 731.100 133.050 734.400 ;
        RECT 134.100 732.600 135.900 733.500 ;
        RECT 139.800 732.600 141.600 740.400 ;
        RECT 151.500 734.400 153.300 740.400 ;
        RECT 157.800 737.400 159.600 740.400 ;
        RECT 134.100 731.700 141.600 732.600 ;
        RECT 142.950 732.450 147.000 733.050 ;
        RECT 77.100 728.100 78.900 728.850 ;
        RECT 82.950 728.550 97.050 729.450 ;
        RECT 82.950 727.950 85.050 728.550 ;
        RECT 94.950 727.950 97.050 728.550 ;
        RECT 100.950 729.450 103.050 730.050 ;
        RECT 109.950 729.450 112.050 730.050 ;
        RECT 100.950 728.550 112.050 729.450 ;
        RECT 100.950 727.950 103.050 728.550 ;
        RECT 109.950 727.950 112.050 728.550 ;
        RECT 115.950 727.950 118.050 730.050 ;
        RECT 121.950 727.950 124.050 730.050 ;
        RECT 127.950 727.950 133.050 730.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 95.100 726.150 96.900 726.900 ;
        RECT 92.100 725.100 93.900 725.850 ;
        RECT 98.100 725.100 99.900 725.850 ;
        RECT 79.950 721.950 82.050 724.050 ;
        RECT 85.950 723.450 90.000 724.050 ;
        RECT 91.950 723.450 94.050 724.050 ;
        RECT 85.950 722.550 94.050 723.450 ;
        RECT 85.950 721.950 90.000 722.550 ;
        RECT 91.950 721.950 94.050 722.550 ;
        RECT 97.950 721.950 100.050 724.050 ;
        RECT 52.950 718.950 55.050 721.050 ;
        RECT 59.100 720.150 60.900 720.900 ;
        RECT 67.950 720.450 72.000 721.050 ;
        RECT 73.950 720.450 76.050 721.050 ;
        RECT 62.100 719.100 63.900 719.850 ;
        RECT 67.950 719.550 76.050 720.450 ;
        RECT 80.100 720.150 81.900 720.900 ;
        RECT 67.950 718.950 72.000 719.550 ;
        RECT 73.950 718.950 76.050 719.550 ;
        RECT 83.100 719.100 84.900 719.850 ;
        RECT 29.400 716.700 37.200 717.600 ;
        RECT 11.700 711.900 18.300 712.800 ;
        RECT 11.700 711.600 12.600 711.900 ;
        RECT 10.800 705.600 12.600 711.600 ;
        RECT 16.800 711.600 18.300 711.900 ;
        RECT 16.800 705.600 18.600 711.600 ;
        RECT 29.400 705.600 31.200 716.700 ;
        RECT 35.400 705.600 37.200 716.700 ;
        RECT 38.400 705.600 40.200 717.600 ;
        RECT 53.700 712.800 54.600 717.900 ;
        RECT 61.950 715.950 64.050 718.050 ;
        RECT 74.700 712.800 75.600 717.900 ;
        RECT 82.950 715.950 85.050 718.050 ;
        RECT 101.700 717.600 102.600 726.900 ;
        RECT 113.100 725.100 114.900 725.850 ;
        RECT 116.850 725.100 118.050 726.900 ;
        RECT 122.100 726.150 123.900 726.900 ;
        RECT 119.100 725.100 120.900 725.850 ;
        RECT 112.950 721.950 115.050 724.050 ;
        RECT 116.850 720.900 117.900 725.100 ;
        RECT 118.950 721.950 121.050 724.050 ;
        RECT 116.850 717.600 118.050 720.900 ;
        RECT 130.950 717.600 132.000 726.900 ;
        RECT 134.100 725.100 135.900 725.850 ;
        RECT 133.950 721.950 136.050 724.050 ;
        RECT 92.400 716.700 100.200 717.600 ;
        RECT 53.700 711.900 60.300 712.800 ;
        RECT 53.700 711.600 54.600 711.900 ;
        RECT 52.800 705.600 54.600 711.600 ;
        RECT 58.800 711.600 60.300 711.900 ;
        RECT 74.700 711.900 81.300 712.800 ;
        RECT 74.700 711.600 75.600 711.900 ;
        RECT 58.800 705.600 60.600 711.600 ;
        RECT 73.800 705.600 75.600 711.600 ;
        RECT 79.800 711.600 81.300 711.900 ;
        RECT 79.800 705.600 81.600 711.600 ;
        RECT 92.400 705.600 94.200 716.700 ;
        RECT 98.400 705.600 100.200 716.700 ;
        RECT 101.400 705.600 103.200 717.600 ;
        RECT 116.700 705.600 118.500 717.600 ;
        RECT 130.200 705.600 132.000 717.600 ;
        RECT 137.550 711.600 138.600 731.700 ;
        RECT 142.950 730.950 147.450 732.450 ;
        RECT 151.800 731.100 153.000 734.400 ;
        RECT 157.800 733.500 159.000 737.400 ;
        RECT 169.800 734.400 171.600 740.400 ;
        RECT 153.900 732.600 159.000 733.500 ;
        RECT 153.900 731.700 155.850 732.600 ;
        RECT 154.950 731.100 155.850 731.700 ;
        RECT 170.400 732.300 171.600 734.400 ;
        RECT 172.800 735.300 174.600 740.400 ;
        RECT 178.800 735.300 180.600 740.400 ;
        RECT 172.800 733.950 180.600 735.300 ;
        RECT 185.400 735.300 187.200 740.400 ;
        RECT 191.400 735.300 193.200 740.400 ;
        RECT 185.400 733.950 193.200 735.300 ;
        RECT 194.400 734.400 196.200 740.400 ;
        RECT 194.400 732.300 195.600 734.400 ;
        RECT 170.400 731.250 174.150 732.300 ;
        RECT 172.950 731.100 174.150 731.250 ;
        RECT 191.850 731.250 195.600 732.300 ;
        RECT 209.100 732.000 210.900 740.400 ;
        RECT 191.850 731.100 193.050 731.250 ;
        RECT 139.950 724.950 142.050 727.050 ;
        RECT 146.550 723.900 147.450 730.950 ;
        RECT 151.950 727.950 154.050 730.050 ;
        RECT 155.100 726.900 155.850 731.100 ;
        RECT 206.700 730.350 210.900 732.000 ;
        RECT 227.100 732.000 228.900 740.400 ;
        RECT 244.200 736.050 246.000 740.400 ;
        RECT 244.200 734.400 249.600 736.050 ;
        RECT 227.100 730.350 231.300 732.000 ;
        RECT 248.700 731.100 249.600 734.400 ;
        RECT 260.400 735.300 262.200 740.400 ;
        RECT 266.400 735.300 268.200 740.400 ;
        RECT 260.400 733.950 268.200 735.300 ;
        RECT 269.400 734.400 271.200 740.400 ;
        RECT 288.000 736.050 289.800 740.400 ;
        RECT 284.400 734.400 289.800 736.050 ;
        RECT 269.400 732.300 270.600 734.400 ;
        RECT 266.850 731.250 270.600 732.300 ;
        RECT 266.850 731.100 268.050 731.250 ;
        RECT 284.400 731.100 285.300 734.400 ;
        RECT 308.100 732.000 309.900 740.400 ;
        RECT 327.300 736.200 329.100 740.400 ;
        RECT 327.150 734.400 329.100 736.200 ;
        RECT 308.100 730.350 312.300 732.000 ;
        RECT 327.150 731.100 328.050 734.400 ;
        RECT 329.100 732.600 330.900 733.500 ;
        RECT 334.800 732.600 336.600 740.400 ;
        RECT 349.200 733.200 351.000 740.400 ;
        RECT 329.100 731.700 336.600 732.600 ;
        RECT 347.400 732.300 351.000 733.200 ;
        RECT 163.950 729.450 166.050 730.050 ;
        RECT 172.950 729.450 175.050 730.050 ;
        RECT 163.950 728.550 175.050 729.450 ;
        RECT 163.950 727.950 166.050 728.550 ;
        RECT 172.950 727.950 175.050 728.550 ;
        RECT 178.950 729.450 181.050 730.050 ;
        RECT 184.950 729.450 187.050 730.050 ;
        RECT 178.950 728.550 187.050 729.450 ;
        RECT 178.950 727.950 181.050 728.550 ;
        RECT 184.950 727.950 187.050 728.550 ;
        RECT 190.950 727.950 193.050 730.050 ;
        RECT 140.100 723.150 141.900 723.900 ;
        RECT 145.950 721.800 148.050 723.900 ;
        RECT 151.800 717.600 153.000 726.900 ;
        RECT 154.950 720.300 155.850 726.900 ;
        RECT 170.100 725.100 171.900 725.850 ;
        RECT 173.850 725.100 175.050 726.900 ;
        RECT 179.100 726.150 180.900 726.900 ;
        RECT 185.100 726.150 186.900 726.900 ;
        RECT 176.100 725.100 177.900 725.850 ;
        RECT 188.100 725.100 189.900 725.850 ;
        RECT 190.950 725.100 192.150 726.900 ;
        RECT 194.100 725.100 195.900 725.850 ;
        RECT 158.100 723.150 159.900 723.900 ;
        RECT 169.950 721.950 172.050 724.050 ;
        RECT 153.900 719.400 155.850 720.300 ;
        RECT 173.850 720.900 174.900 725.100 ;
        RECT 175.950 721.950 178.050 724.050 ;
        RECT 187.950 721.950 190.050 724.050 ;
        RECT 191.100 720.900 192.150 725.100 ;
        RECT 193.950 721.950 196.050 724.050 ;
        RECT 206.700 722.100 207.600 730.350 ;
        RECT 209.100 728.100 210.900 728.850 ;
        RECT 227.100 728.100 228.900 728.850 ;
        RECT 208.950 724.950 211.050 727.200 ;
        RECT 226.950 724.950 229.050 727.050 ;
        RECT 211.950 721.950 214.050 724.050 ;
        RECT 223.950 721.950 226.050 724.050 ;
        RECT 230.400 722.100 231.300 730.350 ;
        RECT 241.950 727.950 244.050 730.050 ;
        RECT 247.950 727.950 253.050 730.050 ;
        RECT 259.950 727.950 262.050 730.050 ;
        RECT 265.950 729.450 268.050 730.050 ;
        RECT 277.800 729.450 279.900 730.050 ;
        RECT 265.950 728.550 279.900 729.450 ;
        RECT 265.950 727.950 268.050 728.550 ;
        RECT 277.800 727.950 279.900 728.550 ;
        RECT 280.950 727.950 286.050 730.050 ;
        RECT 289.950 727.950 292.050 730.050 ;
        RECT 308.100 728.100 309.900 728.850 ;
        RECT 242.100 726.150 243.900 726.900 ;
        RECT 239.100 725.100 240.900 725.850 ;
        RECT 245.100 725.100 246.900 725.850 ;
        RECT 238.950 721.950 241.050 724.050 ;
        RECT 244.950 721.950 247.050 724.050 ;
        RECT 153.900 718.500 159.600 719.400 ;
        RECT 136.800 705.600 138.600 711.600 ;
        RECT 151.500 705.600 153.300 717.600 ;
        RECT 158.400 711.600 159.600 718.500 ;
        RECT 173.850 717.600 175.050 720.900 ;
        RECT 190.950 717.600 192.150 720.900 ;
        RECT 202.950 718.950 208.050 721.050 ;
        RECT 212.100 720.150 213.900 720.900 ;
        RECT 224.100 720.150 225.900 720.900 ;
        RECT 215.100 719.100 216.900 719.850 ;
        RECT 221.100 719.100 222.900 719.850 ;
        RECT 229.950 718.950 232.050 721.050 ;
        RECT 157.800 705.600 159.600 711.600 ;
        RECT 173.700 705.600 175.500 717.600 ;
        RECT 190.500 705.600 192.300 717.600 ;
        RECT 206.700 712.800 207.600 717.900 ;
        RECT 214.950 717.450 217.050 718.050 ;
        RECT 220.950 717.450 223.050 718.050 ;
        RECT 214.950 716.550 223.050 717.450 ;
        RECT 214.950 715.950 217.050 716.550 ;
        RECT 220.950 715.950 223.050 716.550 ;
        RECT 230.400 712.800 231.300 717.900 ;
        RECT 248.700 717.600 249.600 726.900 ;
        RECT 260.100 726.150 261.900 726.900 ;
        RECT 263.100 725.100 264.900 725.850 ;
        RECT 265.950 725.100 267.150 726.900 ;
        RECT 269.100 725.100 270.900 725.850 ;
        RECT 262.950 721.950 265.050 724.050 ;
        RECT 266.100 720.900 267.150 725.100 ;
        RECT 268.950 721.950 271.050 724.050 ;
        RECT 265.950 717.600 267.150 720.900 ;
        RECT 284.400 717.600 285.300 726.900 ;
        RECT 290.100 726.150 291.900 726.900 ;
        RECT 287.100 725.100 288.900 725.850 ;
        RECT 293.100 725.100 294.900 725.850 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 286.950 721.950 289.050 724.050 ;
        RECT 292.950 721.950 295.050 724.050 ;
        RECT 304.950 721.950 307.050 724.050 ;
        RECT 311.400 722.100 312.300 730.350 ;
        RECT 313.950 729.450 316.050 730.050 ;
        RECT 325.950 729.450 328.050 730.050 ;
        RECT 313.950 728.550 328.050 729.450 ;
        RECT 313.950 727.950 316.050 728.550 ;
        RECT 325.950 727.950 328.050 728.550 ;
        RECT 305.100 720.150 306.900 720.900 ;
        RECT 310.950 720.450 313.050 721.050 ;
        RECT 315.000 720.450 319.050 721.050 ;
        RECT 302.100 719.100 303.900 719.850 ;
        RECT 310.950 719.550 319.050 720.450 ;
        RECT 310.950 718.950 313.050 719.550 ;
        RECT 315.000 718.950 319.050 719.550 ;
        RECT 206.700 711.900 213.300 712.800 ;
        RECT 206.700 711.600 207.600 711.900 ;
        RECT 205.800 705.600 207.600 711.600 ;
        RECT 211.800 711.600 213.300 711.900 ;
        RECT 224.700 711.900 231.300 712.800 ;
        RECT 224.700 711.600 226.200 711.900 ;
        RECT 211.800 705.600 213.600 711.600 ;
        RECT 224.400 705.600 226.200 711.600 ;
        RECT 230.400 711.600 231.300 711.900 ;
        RECT 239.400 716.700 247.200 717.600 ;
        RECT 230.400 705.600 232.200 711.600 ;
        RECT 239.400 705.600 241.200 716.700 ;
        RECT 245.400 705.600 247.200 716.700 ;
        RECT 248.400 705.600 250.200 717.600 ;
        RECT 265.500 705.600 267.300 717.600 ;
        RECT 271.950 708.450 274.050 709.050 ;
        RECT 277.950 708.450 280.050 709.050 ;
        RECT 271.950 707.550 280.050 708.450 ;
        RECT 271.950 706.950 274.050 707.550 ;
        RECT 277.950 706.950 280.050 707.550 ;
        RECT 283.800 705.600 285.600 717.600 ;
        RECT 286.800 716.700 294.600 717.600 ;
        RECT 286.800 705.600 288.600 716.700 ;
        RECT 292.800 705.600 294.600 716.700 ;
        RECT 301.950 715.950 304.050 718.050 ;
        RECT 311.400 712.800 312.300 717.900 ;
        RECT 325.950 717.600 327.000 726.900 ;
        RECT 329.100 725.100 330.900 725.850 ;
        RECT 328.950 721.950 331.050 724.050 ;
        RECT 305.700 711.900 312.300 712.800 ;
        RECT 305.700 711.600 307.200 711.900 ;
        RECT 305.400 705.600 307.200 711.600 ;
        RECT 311.400 711.600 312.300 711.900 ;
        RECT 311.400 705.600 313.200 711.600 ;
        RECT 325.200 705.600 327.000 717.600 ;
        RECT 332.550 711.600 333.600 731.700 ;
        RECT 347.400 728.100 348.600 732.300 ;
        RECT 368.100 732.000 369.900 740.400 ;
        RECT 389.100 732.000 390.900 740.400 ;
        RECT 404.400 735.300 406.200 740.400 ;
        RECT 410.400 735.300 412.200 740.400 ;
        RECT 404.400 733.950 412.200 735.300 ;
        RECT 413.400 734.400 415.200 740.400 ;
        RECT 413.400 732.300 414.600 734.400 ;
        RECT 426.000 733.200 427.800 740.400 ;
        RECT 441.300 736.200 443.100 740.400 ;
        RECT 441.150 734.400 443.100 736.200 ;
        RECT 426.000 732.300 429.600 733.200 ;
        RECT 365.700 730.350 369.900 732.000 ;
        RECT 386.700 730.350 390.900 732.000 ;
        RECT 410.850 731.250 414.600 732.300 ;
        RECT 410.850 731.100 412.050 731.250 ;
        RECT 334.950 724.950 337.050 727.050 ;
        RECT 343.950 724.950 349.050 727.050 ;
        RECT 335.100 723.150 336.900 723.900 ;
        RECT 344.100 722.100 345.900 722.850 ;
        RECT 343.950 718.950 346.050 721.050 ;
        RECT 331.800 705.600 333.600 711.600 ;
        RECT 347.400 711.600 348.600 723.900 ;
        RECT 350.100 722.100 351.900 722.850 ;
        RECT 365.700 722.100 366.600 730.350 ;
        RECT 368.100 728.100 369.900 728.850 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 721.950 373.050 724.050 ;
        RECT 386.700 722.100 387.600 730.350 ;
        RECT 394.950 729.450 397.050 730.050 ;
        RECT 403.950 729.450 406.050 730.050 ;
        RECT 389.100 728.100 390.900 728.850 ;
        RECT 394.950 728.550 406.050 729.450 ;
        RECT 394.950 727.950 397.050 728.550 ;
        RECT 403.950 727.950 406.050 728.550 ;
        RECT 409.950 729.450 412.050 730.050 ;
        RECT 418.950 729.450 421.050 730.050 ;
        RECT 409.950 728.550 421.050 729.450 ;
        RECT 409.950 727.950 412.050 728.550 ;
        RECT 418.950 727.950 421.050 728.550 ;
        RECT 428.400 728.100 429.600 732.300 ;
        RECT 433.950 729.450 436.050 733.050 ;
        RECT 441.150 731.100 442.050 734.400 ;
        RECT 443.100 732.600 444.900 733.500 ;
        RECT 448.800 732.600 450.600 740.400 ;
        RECT 443.100 731.700 450.600 732.600 ;
        RECT 468.000 734.400 469.800 740.400 ;
        RECT 439.950 729.450 442.050 730.050 ;
        RECT 433.950 729.000 442.050 729.450 ;
        RECT 434.550 728.550 442.050 729.000 ;
        RECT 439.950 727.950 442.050 728.550 ;
        RECT 388.950 724.950 391.050 727.200 ;
        RECT 404.100 726.150 405.900 726.900 ;
        RECT 407.100 725.100 408.900 725.850 ;
        RECT 409.950 725.100 411.150 726.900 ;
        RECT 413.100 725.100 414.900 725.850 ;
        RECT 391.950 721.950 394.050 724.050 ;
        RECT 406.950 721.950 409.050 724.050 ;
        RECT 349.950 718.950 352.050 721.050 ;
        RECT 358.950 720.450 363.000 721.050 ;
        RECT 364.950 720.450 367.050 721.050 ;
        RECT 358.950 719.550 367.050 720.450 ;
        RECT 371.100 720.150 372.900 720.900 ;
        RECT 379.950 720.450 384.000 721.050 ;
        RECT 385.950 720.450 388.050 721.050 ;
        RECT 410.100 720.900 411.150 725.100 ;
        RECT 424.950 724.950 430.050 727.050 ;
        RECT 412.950 721.950 415.050 724.050 ;
        RECT 425.100 722.100 426.900 722.850 ;
        RECT 358.950 718.950 363.000 719.550 ;
        RECT 364.950 718.950 367.050 719.550 ;
        RECT 374.100 719.100 375.900 719.850 ;
        RECT 379.950 719.550 388.050 720.450 ;
        RECT 392.100 720.150 393.900 720.900 ;
        RECT 379.950 718.950 384.000 719.550 ;
        RECT 385.950 718.950 388.050 719.550 ;
        RECT 395.100 719.100 396.900 719.850 ;
        RECT 365.700 712.800 366.600 717.900 ;
        RECT 373.950 715.950 376.050 718.050 ;
        RECT 386.700 712.800 387.600 717.900 ;
        RECT 394.950 715.950 397.050 718.050 ;
        RECT 409.950 717.600 411.150 720.900 ;
        RECT 424.950 718.950 427.050 721.050 ;
        RECT 365.700 711.900 372.300 712.800 ;
        RECT 365.700 711.600 366.600 711.900 ;
        RECT 347.400 705.600 349.200 711.600 ;
        RECT 364.800 705.600 366.600 711.600 ;
        RECT 370.800 711.600 372.300 711.900 ;
        RECT 386.700 711.900 393.300 712.800 ;
        RECT 386.700 711.600 387.600 711.900 ;
        RECT 370.800 705.600 372.600 711.600 ;
        RECT 385.800 705.600 387.600 711.600 ;
        RECT 391.800 711.600 393.300 711.900 ;
        RECT 391.800 705.600 393.600 711.600 ;
        RECT 409.500 705.600 411.300 717.600 ;
        RECT 428.400 711.600 429.600 723.900 ;
        RECT 431.100 722.100 432.900 722.850 ;
        RECT 430.950 718.950 433.050 721.050 ;
        RECT 439.950 717.600 441.000 726.900 ;
        RECT 443.100 725.100 444.900 725.850 ;
        RECT 442.950 721.950 445.050 724.050 ;
        RECT 427.800 705.600 429.600 711.600 ;
        RECT 439.200 705.600 441.000 717.600 ;
        RECT 446.550 711.600 447.600 731.700 ;
        RECT 468.000 731.100 469.050 734.400 ;
        RECT 482.400 732.600 484.200 740.400 ;
        RECT 489.900 736.200 491.700 740.400 ;
        RECT 504.300 736.200 506.100 740.400 ;
        RECT 489.900 734.400 491.850 736.200 ;
        RECT 488.100 732.600 489.900 733.500 ;
        RECT 482.400 731.700 489.900 732.600 ;
        RECT 460.950 727.950 463.050 730.050 ;
        RECT 466.950 727.950 469.050 730.050 ;
        RECT 472.950 727.950 478.050 730.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 461.100 726.150 462.900 726.900 ;
        RECT 464.250 725.100 466.050 725.850 ;
        RECT 466.950 725.100 467.850 726.900 ;
        RECT 472.950 726.150 474.750 726.900 ;
        RECT 469.950 725.100 471.750 725.850 ;
        RECT 449.100 723.150 450.900 723.900 ;
        RECT 463.950 721.950 466.050 724.050 ;
        RECT 467.100 720.900 467.850 725.100 ;
        RECT 481.950 724.950 484.050 727.050 ;
        RECT 469.950 721.950 472.050 724.050 ;
        RECT 482.100 723.150 483.900 723.900 ;
        RECT 466.950 719.400 467.850 720.900 ;
        RECT 463.800 718.500 467.850 719.400 ;
        RECT 445.800 705.600 447.600 711.600 ;
        RECT 460.800 706.500 462.600 717.600 ;
        RECT 463.800 707.400 465.600 718.500 ;
        RECT 466.800 716.400 474.600 717.300 ;
        RECT 466.800 706.500 468.600 716.400 ;
        RECT 460.800 705.600 468.600 706.500 ;
        RECT 472.800 705.600 474.600 716.400 ;
        RECT 485.400 711.600 486.450 731.700 ;
        RECT 490.950 731.100 491.850 734.400 ;
        RECT 504.150 734.400 506.100 736.200 ;
        RECT 504.150 731.100 505.050 734.400 ;
        RECT 506.100 732.600 507.900 733.500 ;
        RECT 511.800 732.600 513.600 740.400 ;
        RECT 506.100 731.700 513.600 732.600 ;
        RECT 518.400 732.600 520.200 740.400 ;
        RECT 525.900 736.200 527.700 740.400 ;
        RECT 525.900 734.400 527.850 736.200 ;
        RECT 524.100 732.600 525.900 733.500 ;
        RECT 518.400 731.700 525.900 732.600 ;
        RECT 487.950 727.950 493.050 730.050 ;
        RECT 502.950 727.950 505.050 730.050 ;
        RECT 488.100 725.100 489.900 725.850 ;
        RECT 487.950 721.950 490.050 724.050 ;
        RECT 492.000 717.600 493.050 726.900 ;
        RECT 502.950 717.600 504.000 726.900 ;
        RECT 506.100 725.100 507.900 725.850 ;
        RECT 505.950 721.950 508.050 724.050 ;
        RECT 485.400 705.600 487.200 711.600 ;
        RECT 492.000 705.600 493.800 717.600 ;
        RECT 502.200 705.600 504.000 717.600 ;
        RECT 509.550 711.600 510.600 731.700 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 517.950 724.950 520.050 727.050 ;
        RECT 512.100 723.150 513.900 723.900 ;
        RECT 518.100 723.150 519.900 723.900 ;
        RECT 508.800 705.600 510.600 711.600 ;
        RECT 521.400 711.600 522.450 731.700 ;
        RECT 526.950 731.100 527.850 734.400 ;
        RECT 549.000 734.400 550.800 740.400 ;
        RECT 549.000 731.100 550.050 734.400 ;
        RECT 563.400 732.600 565.200 740.400 ;
        RECT 570.900 736.200 572.700 740.400 ;
        RECT 570.900 734.400 572.850 736.200 ;
        RECT 569.100 732.600 570.900 733.500 ;
        RECT 563.400 731.700 570.900 732.600 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 541.950 727.950 544.050 730.050 ;
        RECT 547.950 727.950 550.050 730.050 ;
        RECT 553.950 727.950 556.050 730.050 ;
        RECT 524.100 725.100 525.900 725.850 ;
        RECT 523.950 721.950 526.050 724.050 ;
        RECT 528.000 717.600 529.050 726.900 ;
        RECT 542.100 726.150 543.900 726.900 ;
        RECT 545.250 725.100 547.050 725.850 ;
        RECT 547.950 725.100 548.850 726.900 ;
        RECT 553.950 726.150 555.750 726.900 ;
        RECT 550.950 725.100 552.750 725.850 ;
        RECT 544.950 721.950 547.050 724.050 ;
        RECT 548.100 720.900 548.850 725.100 ;
        RECT 562.950 724.950 565.050 727.050 ;
        RECT 550.950 721.950 553.050 724.050 ;
        RECT 563.100 723.150 564.900 723.900 ;
        RECT 547.950 719.400 548.850 720.900 ;
        RECT 544.800 718.500 548.850 719.400 ;
        RECT 521.400 705.600 523.200 711.600 ;
        RECT 528.000 705.600 529.800 717.600 ;
        RECT 541.800 706.500 543.600 717.600 ;
        RECT 544.800 707.400 546.600 718.500 ;
        RECT 547.800 716.400 555.600 717.300 ;
        RECT 547.800 706.500 549.600 716.400 ;
        RECT 541.800 705.600 549.600 706.500 ;
        RECT 553.800 705.600 555.600 716.400 ;
        RECT 566.400 711.600 567.450 731.700 ;
        RECT 571.950 731.100 572.850 734.400 ;
        RECT 589.200 733.200 591.000 740.400 ;
        RECT 606.000 736.050 607.800 740.400 ;
        RECT 587.400 732.300 591.000 733.200 ;
        RECT 602.400 734.400 607.800 736.050 ;
        RECT 568.950 727.950 574.050 730.050 ;
        RECT 587.400 728.100 588.600 732.300 ;
        RECT 602.400 731.100 603.300 734.400 ;
        RECT 620.400 732.600 622.200 740.400 ;
        RECT 627.900 736.200 629.700 740.400 ;
        RECT 646.800 737.400 648.600 740.400 ;
        RECT 627.900 734.400 629.850 736.200 ;
        RECT 626.100 732.600 627.900 733.500 ;
        RECT 620.400 731.700 627.900 732.600 ;
        RECT 569.100 725.100 570.900 725.850 ;
        RECT 568.950 721.950 571.050 724.050 ;
        RECT 573.000 717.600 574.050 726.900 ;
        RECT 586.950 726.450 589.050 727.050 ;
        RECT 595.950 726.450 598.050 730.050 ;
        RECT 601.950 727.950 604.050 730.050 ;
        RECT 607.950 727.950 610.050 730.050 ;
        RECT 586.950 726.000 598.050 726.450 ;
        RECT 586.950 725.550 597.450 726.000 ;
        RECT 586.950 724.950 589.050 725.550 ;
        RECT 584.100 722.100 585.900 722.850 ;
        RECT 583.950 718.950 586.050 721.050 ;
        RECT 566.400 705.600 568.200 711.600 ;
        RECT 573.000 705.600 574.800 717.600 ;
        RECT 587.400 711.600 588.600 723.900 ;
        RECT 590.100 722.100 591.900 722.850 ;
        RECT 589.950 718.950 592.050 721.050 ;
        RECT 602.400 717.600 603.300 726.900 ;
        RECT 608.100 726.150 609.900 726.900 ;
        RECT 605.100 725.100 606.900 725.850 ;
        RECT 611.100 725.100 612.900 725.850 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 604.950 721.950 607.050 724.050 ;
        RECT 610.950 721.950 613.050 724.050 ;
        RECT 620.100 723.150 621.900 723.900 ;
        RECT 587.400 705.600 589.200 711.600 ;
        RECT 601.800 705.600 603.600 717.600 ;
        RECT 604.800 716.700 612.600 717.600 ;
        RECT 604.800 705.600 606.600 716.700 ;
        RECT 610.800 705.600 612.600 716.700 ;
        RECT 623.400 711.600 624.450 731.700 ;
        RECT 628.950 731.100 629.850 734.400 ;
        RECT 647.400 734.100 648.600 737.400 ;
        RECT 664.200 733.200 666.000 740.400 ;
        RECT 682.200 736.050 684.000 740.400 ;
        RECT 698.400 737.400 700.200 740.400 ;
        RECT 712.800 737.400 714.600 740.400 ;
        RECT 682.200 734.400 687.600 736.050 ;
        RECT 646.950 732.450 649.050 733.050 ;
        RECT 658.950 732.450 661.050 733.050 ;
        RECT 646.950 731.550 661.050 732.450 ;
        RECT 646.950 730.950 649.050 731.550 ;
        RECT 658.950 730.950 661.050 731.550 ;
        RECT 662.400 732.300 666.000 733.200 ;
        RECT 634.950 730.050 637.050 730.200 ;
        RECT 628.950 729.450 631.050 730.050 ;
        RECT 633.000 729.450 637.050 730.050 ;
        RECT 628.950 728.550 637.050 729.450 ;
        RECT 628.950 727.950 631.050 728.550 ;
        RECT 633.000 728.100 637.050 728.550 ;
        RECT 646.950 728.100 648.300 729.900 ;
        RECT 662.400 728.100 663.600 732.300 ;
        RECT 686.700 731.100 687.600 734.400 ;
        RECT 679.950 729.450 682.050 730.050 ;
        RECT 671.550 728.550 682.050 729.450 ;
        RECT 633.000 727.950 636.000 728.100 ;
        RECT 626.100 725.100 627.900 725.850 ;
        RECT 625.950 721.950 628.050 724.050 ;
        RECT 630.000 717.600 631.050 726.900 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 647.100 723.900 648.300 728.100 ;
        RECT 661.950 726.450 664.050 727.050 ;
        RECT 671.550 726.450 672.450 728.550 ;
        RECT 679.950 727.950 682.050 728.550 ;
        RECT 685.950 727.950 688.050 730.050 ;
        RECT 694.950 727.950 697.050 730.050 ;
        RECT 661.950 725.550 672.450 726.450 ;
        RECT 680.100 726.150 681.900 726.900 ;
        RECT 661.950 724.950 664.050 725.550 ;
        RECT 677.100 725.100 678.900 725.850 ;
        RECT 683.100 725.100 684.900 725.850 ;
        RECT 644.100 723.150 645.900 723.900 ;
        RECT 646.950 718.650 648.300 723.900 ;
        RECT 649.950 721.950 652.050 724.050 ;
        RECT 659.100 722.100 660.900 722.850 ;
        RECT 650.100 720.150 651.900 720.900 ;
        RECT 658.950 718.950 661.050 721.050 ;
        RECT 645.600 717.600 648.300 718.650 ;
        RECT 623.400 705.600 625.200 711.600 ;
        RECT 630.000 705.600 631.800 717.600 ;
        RECT 645.600 705.600 647.400 717.600 ;
        RECT 662.400 711.600 663.600 723.900 ;
        RECT 665.100 722.100 666.900 722.850 ;
        RECT 676.950 721.950 679.050 724.050 ;
        RECT 682.950 721.950 685.050 724.050 ;
        RECT 664.950 718.950 667.050 721.050 ;
        RECT 686.700 717.600 687.600 726.900 ;
        RECT 695.100 726.150 696.900 726.900 ;
        RECT 698.400 725.100 699.600 737.400 ;
        RECT 713.400 725.100 714.600 737.400 ;
        RECT 725.400 737.400 727.200 740.400 ;
        RECT 715.950 727.950 718.050 730.050 ;
        RECT 721.950 727.950 724.050 730.050 ;
        RECT 716.100 726.150 717.900 726.900 ;
        RECT 722.100 726.150 723.900 726.900 ;
        RECT 725.400 725.100 726.600 737.400 ;
        RECT 743.100 732.000 744.900 740.400 ;
        RECT 740.700 730.350 744.900 732.000 ;
        RECT 764.100 732.000 765.900 740.400 ;
        RECT 785.100 732.000 786.900 740.400 ;
        RECT 801.000 733.200 802.800 740.400 ;
        RECT 801.000 732.300 804.600 733.200 ;
        RECT 764.100 730.350 768.300 732.000 ;
        RECT 785.100 730.350 789.300 732.000 ;
        RECT 697.950 723.450 700.050 724.050 ;
        RECT 706.950 723.450 709.050 724.050 ;
        RECT 697.950 722.550 709.050 723.450 ;
        RECT 697.950 721.950 700.050 722.550 ;
        RECT 706.950 721.950 709.050 722.550 ;
        RECT 712.950 721.950 715.050 724.050 ;
        RECT 724.950 721.950 727.050 724.050 ;
        RECT 740.700 722.100 741.600 730.350 ;
        RECT 743.100 728.100 744.900 728.850 ;
        RECT 764.100 728.100 765.900 728.850 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 763.950 724.950 766.050 727.050 ;
        RECT 745.950 721.950 748.050 724.050 ;
        RECT 760.950 721.950 763.050 724.050 ;
        RECT 767.400 722.100 768.300 730.350 ;
        RECT 785.100 728.100 786.900 728.850 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 781.950 721.950 784.050 724.050 ;
        RECT 788.400 722.100 789.300 730.350 ;
        RECT 803.400 728.100 804.600 732.300 ;
        RECT 818.100 732.000 819.900 740.400 ;
        RECT 815.700 730.350 819.900 732.000 ;
        RECT 793.950 726.450 796.050 727.050 ;
        RECT 802.950 726.450 805.050 727.050 ;
        RECT 793.950 725.550 805.050 726.450 ;
        RECT 793.950 724.950 796.050 725.550 ;
        RECT 802.950 724.950 805.050 725.550 ;
        RECT 800.100 722.100 801.900 722.850 ;
        RECT 677.400 716.700 685.200 717.600 ;
        RECT 662.400 705.600 664.200 711.600 ;
        RECT 677.400 705.600 679.200 716.700 ;
        RECT 683.400 705.600 685.200 716.700 ;
        RECT 686.400 705.600 688.200 717.600 ;
        RECT 698.400 711.600 699.600 720.900 ;
        RECT 713.400 711.600 714.600 720.900 ;
        RECT 698.400 705.600 700.200 711.600 ;
        RECT 712.800 705.600 714.600 711.600 ;
        RECT 725.400 711.600 726.600 720.900 ;
        RECT 739.950 718.950 742.050 721.050 ;
        RECT 746.100 720.150 747.900 720.900 ;
        RECT 761.100 720.150 762.900 720.900 ;
        RECT 749.100 719.100 750.900 719.850 ;
        RECT 758.100 719.100 759.900 719.850 ;
        RECT 766.950 718.950 769.050 721.050 ;
        RECT 782.100 720.150 783.900 720.900 ;
        RECT 779.100 719.100 780.900 719.850 ;
        RECT 787.950 718.950 793.050 721.050 ;
        RECT 799.950 718.950 802.050 721.050 ;
        RECT 740.700 712.800 741.600 717.900 ;
        RECT 748.950 715.950 751.050 718.050 ;
        RECT 757.950 715.950 760.050 718.050 ;
        RECT 767.400 712.800 768.300 717.900 ;
        RECT 778.950 715.950 781.050 718.050 ;
        RECT 788.400 712.800 789.300 717.900 ;
        RECT 740.700 711.900 747.300 712.800 ;
        RECT 740.700 711.600 741.600 711.900 ;
        RECT 725.400 705.600 727.200 711.600 ;
        RECT 739.800 705.600 741.600 711.600 ;
        RECT 745.800 711.600 747.300 711.900 ;
        RECT 761.700 711.900 768.300 712.800 ;
        RECT 761.700 711.600 763.200 711.900 ;
        RECT 745.800 705.600 747.600 711.600 ;
        RECT 761.400 705.600 763.200 711.600 ;
        RECT 767.400 711.600 768.300 711.900 ;
        RECT 782.700 711.900 789.300 712.800 ;
        RECT 782.700 711.600 784.200 711.900 ;
        RECT 767.400 705.600 769.200 711.600 ;
        RECT 782.400 705.600 784.200 711.600 ;
        RECT 788.400 711.600 789.300 711.900 ;
        RECT 803.400 711.600 804.600 723.900 ;
        RECT 806.100 722.100 807.900 722.850 ;
        RECT 815.700 722.100 816.600 730.350 ;
        RECT 818.100 728.100 819.900 728.850 ;
        RECT 817.950 724.950 820.050 727.050 ;
        RECT 820.950 721.800 823.050 724.050 ;
        RECT 805.950 718.950 808.050 721.050 ;
        RECT 811.950 718.950 817.050 721.050 ;
        RECT 821.100 720.150 822.900 720.900 ;
        RECT 824.100 719.100 825.900 719.850 ;
        RECT 815.700 712.800 816.600 717.900 ;
        RECT 823.950 715.950 826.050 718.050 ;
        RECT 815.700 711.900 822.300 712.800 ;
        RECT 815.700 711.600 816.600 711.900 ;
        RECT 788.400 705.600 790.200 711.600 ;
        RECT 802.800 705.600 804.600 711.600 ;
        RECT 814.800 705.600 816.600 711.600 ;
        RECT 820.800 711.600 822.300 711.900 ;
        RECT 820.800 705.600 822.600 711.600 ;
        RECT 13.800 695.400 15.600 701.400 ;
        RECT 26.400 695.400 28.200 701.400 ;
        RECT 10.950 685.950 13.050 688.050 ;
        RECT 11.100 684.150 12.900 684.900 ;
        RECT 14.400 683.100 15.600 695.400 ;
        RECT 26.700 695.100 28.200 695.400 ;
        RECT 32.400 695.400 34.200 701.400 ;
        RECT 32.400 695.100 33.300 695.400 ;
        RECT 26.700 694.200 33.300 695.100 ;
        RECT 22.950 688.950 25.050 691.050 ;
        RECT 32.400 689.100 33.300 694.200 ;
        RECT 41.400 690.300 43.200 701.400 ;
        RECT 47.400 690.300 49.200 701.400 ;
        RECT 41.400 689.400 49.200 690.300 ;
        RECT 50.400 689.400 52.200 701.400 ;
        RECT 67.500 689.400 69.300 701.400 ;
        RECT 85.800 689.400 87.600 701.400 ;
        RECT 88.800 690.300 90.600 701.400 ;
        RECT 94.800 690.300 96.600 701.400 ;
        RECT 88.800 689.400 96.600 690.300 ;
        RECT 107.400 695.400 109.200 701.400 ;
        RECT 16.950 685.950 19.050 688.050 ;
        RECT 23.100 687.150 24.900 687.900 ;
        RECT 26.100 686.100 27.900 686.850 ;
        RECT 31.950 685.950 34.050 688.050 ;
        RECT 17.100 684.150 18.900 684.900 ;
        RECT 25.950 682.950 28.050 685.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 28.950 679.800 31.050 682.050 ;
        RECT 14.400 674.700 15.600 678.900 ;
        RECT 29.100 678.150 30.900 678.900 ;
        RECT 32.400 676.650 33.300 684.900 ;
        RECT 37.950 682.950 43.050 685.050 ;
        RECT 46.950 682.950 49.050 685.050 ;
        RECT 41.100 681.150 42.900 681.900 ;
        RECT 47.100 681.150 48.900 681.900 ;
        RECT 44.100 680.100 45.900 680.850 ;
        RECT 50.700 680.100 51.600 689.400 ;
        RECT 67.950 686.100 69.150 689.400 ;
        RECT 64.950 682.950 67.050 685.050 ;
        RECT 68.100 681.900 69.150 686.100 ;
        RECT 70.950 682.950 73.050 685.050 ;
        RECT 65.100 681.150 66.900 681.900 ;
        RECT 62.100 680.100 63.900 680.850 ;
        RECT 67.950 680.100 69.150 681.900 ;
        RECT 71.100 681.150 72.900 681.900 ;
        RECT 86.400 680.100 87.300 689.400 ;
        RECT 88.950 682.950 91.050 685.050 ;
        RECT 94.950 682.950 97.050 685.050 ;
        RECT 100.950 684.450 103.050 688.050 ;
        RECT 107.400 686.100 108.600 695.400 ;
        RECT 118.200 689.400 120.000 701.400 ;
        RECT 124.800 695.400 126.600 701.400 ;
        RECT 106.950 684.450 109.050 685.050 ;
        RECT 100.950 684.000 109.050 684.450 ;
        RECT 101.550 683.550 109.050 684.000 ;
        RECT 106.950 682.950 109.050 683.550 ;
        RECT 89.100 681.150 90.900 681.900 ;
        RECT 95.100 681.150 96.900 681.900 ;
        RECT 92.100 680.100 93.900 680.850 ;
        RECT 104.100 680.100 105.900 680.850 ;
        RECT 34.950 678.450 37.050 679.050 ;
        RECT 43.950 678.450 46.050 679.050 ;
        RECT 34.950 677.550 46.050 678.450 ;
        RECT 34.950 676.950 37.050 677.550 ;
        RECT 43.950 676.950 46.050 677.550 ;
        RECT 49.950 676.950 54.900 679.050 ;
        RECT 55.950 678.450 60.000 679.050 ;
        RECT 61.950 678.450 64.050 679.050 ;
        RECT 55.950 677.550 64.050 678.450 ;
        RECT 55.950 676.950 60.000 677.550 ;
        RECT 61.950 676.950 64.050 677.550 ;
        RECT 67.950 678.450 70.050 679.050 ;
        RECT 76.800 678.450 78.900 679.050 ;
        RECT 67.950 677.550 78.900 678.450 ;
        RECT 67.950 676.950 70.050 677.550 ;
        RECT 76.800 676.950 78.900 677.550 ;
        RECT 79.950 678.450 84.000 679.050 ;
        RECT 85.950 678.450 88.050 679.050 ;
        RECT 79.950 677.550 88.050 678.450 ;
        RECT 79.950 676.950 84.000 677.550 ;
        RECT 85.950 676.950 88.050 677.550 ;
        RECT 91.950 676.950 94.050 679.050 ;
        RECT 103.950 676.950 106.050 679.050 ;
        RECT 12.000 673.800 15.600 674.700 ;
        RECT 29.100 675.000 33.300 676.650 ;
        RECT 12.000 666.600 13.800 673.800 ;
        RECT 29.100 666.600 30.900 675.000 ;
        RECT 50.700 672.600 51.600 675.900 ;
        RECT 68.850 675.750 70.050 675.900 ;
        RECT 68.850 674.700 72.600 675.750 ;
        RECT 46.200 670.950 51.600 672.600 ;
        RECT 62.400 671.700 70.200 673.050 ;
        RECT 46.200 666.600 48.000 670.950 ;
        RECT 62.400 666.600 64.200 671.700 ;
        RECT 68.400 666.600 70.200 671.700 ;
        RECT 71.400 672.600 72.600 674.700 ;
        RECT 86.400 672.600 87.300 675.900 ;
        RECT 71.400 666.600 73.200 672.600 ;
        RECT 86.400 670.950 91.800 672.600 ;
        RECT 90.000 666.600 91.800 670.950 ;
        RECT 107.400 669.600 108.600 681.900 ;
        RECT 118.950 680.100 120.000 689.400 ;
        RECT 121.950 682.950 124.050 685.050 ;
        RECT 122.100 681.150 123.900 681.900 ;
        RECT 118.950 676.950 121.050 679.050 ;
        RECT 120.150 672.600 121.050 675.900 ;
        RECT 125.550 675.300 126.600 695.400 ;
        RECT 137.400 695.400 139.200 701.400 ;
        RECT 154.800 695.400 156.600 701.400 ;
        RECT 133.950 685.950 136.050 688.050 ;
        RECT 134.100 684.150 135.900 684.900 ;
        RECT 128.100 683.100 129.900 683.850 ;
        RECT 137.400 683.100 138.600 695.400 ;
        RECT 155.700 695.100 156.600 695.400 ;
        RECT 160.800 695.400 162.600 701.400 ;
        RECT 175.800 695.400 177.600 701.400 ;
        RECT 160.800 695.100 162.300 695.400 ;
        RECT 155.700 694.200 162.300 695.100 ;
        RECT 176.700 695.100 177.600 695.400 ;
        RECT 181.800 695.400 183.600 701.400 ;
        RECT 181.800 695.100 183.300 695.400 ;
        RECT 176.700 694.200 183.300 695.100 ;
        RECT 155.700 689.100 156.600 694.200 ;
        RECT 163.950 688.950 166.050 691.050 ;
        RECT 176.700 689.100 177.600 694.200 ;
        RECT 184.950 688.950 187.050 691.050 ;
        RECT 191.400 690.300 193.200 701.400 ;
        RECT 197.400 690.300 199.200 701.400 ;
        RECT 191.400 689.400 199.200 690.300 ;
        RECT 200.400 689.400 202.200 701.400 ;
        RECT 214.800 689.400 216.600 701.400 ;
        RECT 217.800 690.300 219.600 701.400 ;
        RECT 223.800 690.300 225.600 701.400 ;
        RECT 232.800 695.400 234.600 701.400 ;
        RECT 217.800 689.400 225.600 690.300 ;
        RECT 233.700 695.100 234.600 695.400 ;
        RECT 238.800 695.400 240.600 701.400 ;
        RECT 254.400 695.400 256.200 701.400 ;
        RECT 238.800 695.100 240.300 695.400 ;
        RECT 233.700 694.200 240.300 695.100 ;
        RECT 139.950 685.950 142.050 688.050 ;
        RECT 151.950 685.950 157.050 688.050 ;
        RECT 164.100 687.150 165.900 687.900 ;
        RECT 169.950 687.450 174.000 688.050 ;
        RECT 175.950 687.450 178.050 688.050 ;
        RECT 161.100 686.100 162.900 686.850 ;
        RECT 169.950 686.550 178.050 687.450 ;
        RECT 185.100 687.150 186.900 687.900 ;
        RECT 169.950 685.950 174.000 686.550 ;
        RECT 175.950 685.950 178.050 686.550 ;
        RECT 182.100 686.100 183.900 686.850 ;
        RECT 140.100 684.150 141.900 684.900 ;
        RECT 127.950 679.950 130.050 682.050 ;
        RECT 136.950 679.950 139.050 682.050 ;
        RECT 122.100 674.400 129.600 675.300 ;
        RECT 122.100 673.500 123.900 674.400 ;
        RECT 120.150 670.800 122.100 672.600 ;
        RECT 107.400 666.600 109.200 669.600 ;
        RECT 120.300 666.600 122.100 670.800 ;
        RECT 127.800 666.600 129.600 674.400 ;
        RECT 137.400 674.700 138.600 678.900 ;
        RECT 155.700 676.650 156.600 684.900 ;
        RECT 160.950 682.950 163.050 685.200 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 158.100 678.150 159.900 678.900 ;
        RECT 176.700 676.650 177.600 684.900 ;
        RECT 181.950 682.950 184.050 685.050 ;
        RECT 190.950 682.950 193.050 685.050 ;
        RECT 196.950 682.950 199.050 685.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 191.100 681.150 192.900 681.900 ;
        RECT 197.100 681.150 198.900 681.900 ;
        RECT 194.100 680.100 195.900 680.850 ;
        RECT 200.700 680.100 201.600 689.400 ;
        RECT 215.400 680.100 216.300 689.400 ;
        RECT 233.700 689.100 234.600 694.200 ;
        RECT 241.950 688.950 244.050 691.050 ;
        RECT 230.550 687.900 235.050 688.050 ;
        RECT 229.950 685.950 235.050 687.900 ;
        RECT 242.100 687.150 243.900 687.900 ;
        RECT 239.100 686.100 240.900 686.850 ;
        RECT 254.400 686.100 255.600 695.400 ;
        RECT 263.400 690.600 265.200 701.400 ;
        RECT 269.400 700.500 277.200 701.400 ;
        RECT 269.400 690.600 271.200 700.500 ;
        RECT 263.400 689.700 271.200 690.600 ;
        RECT 272.400 688.500 274.200 699.600 ;
        RECT 275.400 689.400 277.200 700.500 ;
        RECT 291.600 689.400 293.400 701.400 ;
        RECT 305.400 695.400 307.200 701.400 ;
        RECT 305.700 695.100 307.200 695.400 ;
        RECT 311.400 695.400 313.200 701.400 ;
        RECT 325.800 695.400 327.600 701.400 ;
        RECT 343.800 695.400 345.600 701.400 ;
        RECT 311.400 695.100 312.300 695.400 ;
        RECT 305.700 694.200 312.300 695.100 ;
        RECT 270.150 687.600 274.200 688.500 ;
        RECT 290.700 688.350 293.400 689.400 ;
        RECT 301.950 688.950 304.050 691.050 ;
        RECT 311.400 689.100 312.300 694.200 ;
        RECT 270.150 686.100 271.050 687.600 ;
        RECT 287.100 686.100 288.900 686.850 ;
        RECT 229.950 685.800 232.050 685.950 ;
        RECT 217.950 682.950 220.050 685.050 ;
        RECT 223.950 682.950 226.050 685.050 ;
        RECT 218.100 681.150 219.900 681.900 ;
        RECT 224.100 681.150 225.900 681.900 ;
        RECT 221.100 680.100 222.900 680.850 ;
        RECT 179.100 678.150 180.900 678.900 ;
        RECT 193.950 676.950 196.050 679.050 ;
        RECT 199.950 676.950 205.050 679.050 ;
        RECT 214.950 676.950 217.050 679.050 ;
        RECT 220.950 676.950 223.050 679.050 ;
        RECT 233.700 676.650 234.600 684.900 ;
        RECT 238.950 682.950 241.050 685.050 ;
        RECT 253.950 682.950 259.050 685.050 ;
        RECT 265.950 682.950 268.050 685.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 270.150 681.900 270.900 686.100 ;
        RECT 271.950 682.950 274.050 685.050 ;
        RECT 286.950 682.950 289.050 685.050 ;
        RECT 290.700 683.100 292.050 688.350 ;
        RECT 302.100 687.150 303.900 687.900 ;
        RECT 305.100 686.100 306.900 686.850 ;
        RECT 310.950 685.950 313.050 688.050 ;
        RECT 322.950 685.950 325.050 688.050 ;
        RECT 293.100 683.100 294.900 683.850 ;
        RECT 251.100 680.100 252.900 680.850 ;
        RECT 236.100 678.150 237.900 678.900 ;
        RECT 250.950 676.950 253.050 679.050 ;
        RECT 155.700 675.000 159.900 676.650 ;
        RECT 176.700 675.000 180.900 676.650 ;
        RECT 137.400 673.800 141.000 674.700 ;
        RECT 139.200 666.600 141.000 673.800 ;
        RECT 142.950 669.450 145.050 670.050 ;
        RECT 151.950 669.450 154.050 670.050 ;
        RECT 142.950 668.550 154.050 669.450 ;
        RECT 142.950 667.950 145.050 668.550 ;
        RECT 151.950 667.950 154.050 668.550 ;
        RECT 158.100 666.600 159.900 675.000 ;
        RECT 179.100 666.600 180.900 675.000 ;
        RECT 200.700 672.600 201.600 675.900 ;
        RECT 196.200 670.950 201.600 672.600 ;
        RECT 215.400 672.600 216.300 675.900 ;
        RECT 233.700 675.000 237.900 676.650 ;
        RECT 215.400 670.950 220.800 672.600 ;
        RECT 196.200 666.600 198.000 670.950 ;
        RECT 219.000 666.600 220.800 670.950 ;
        RECT 236.100 666.600 237.900 675.000 ;
        RECT 254.400 669.600 255.600 681.900 ;
        RECT 266.250 681.150 268.050 681.900 ;
        RECT 263.250 680.100 265.050 680.850 ;
        RECT 270.150 680.100 271.050 681.900 ;
        RECT 271.950 681.150 273.750 681.900 ;
        RECT 275.100 680.100 276.900 680.850 ;
        RECT 262.950 676.950 265.050 679.050 ;
        RECT 268.950 676.950 271.050 679.050 ;
        RECT 274.950 676.950 277.050 679.050 ;
        RECT 290.700 678.900 291.900 683.100 ;
        RECT 304.950 682.950 307.050 685.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 290.700 677.100 292.050 678.900 ;
        RECT 308.100 678.150 309.900 678.900 ;
        RECT 311.400 676.650 312.300 684.900 ;
        RECT 323.100 684.150 324.900 684.900 ;
        RECT 326.400 683.100 327.600 695.400 ;
        RECT 328.950 685.950 331.050 688.050 ;
        RECT 329.100 684.150 330.900 684.900 ;
        RECT 341.100 684.150 342.900 684.900 ;
        RECT 344.400 683.100 345.600 695.400 ;
        RECT 346.950 685.950 349.050 691.050 ;
        RECT 355.800 689.400 357.600 701.400 ;
        RECT 358.800 690.300 360.600 701.400 ;
        RECT 364.800 690.300 366.600 701.400 ;
        RECT 376.800 695.400 378.600 701.400 ;
        RECT 358.800 689.400 366.600 690.300 ;
        RECT 377.700 695.100 378.600 695.400 ;
        RECT 382.800 695.400 384.600 701.400 ;
        RECT 382.800 695.100 384.300 695.400 ;
        RECT 377.700 694.200 384.300 695.100 ;
        RECT 347.100 684.150 348.900 684.900 ;
        RECT 325.950 681.450 328.050 682.050 ;
        RECT 334.950 681.450 337.050 682.200 ;
        RECT 325.950 680.550 337.050 681.450 ;
        RECT 325.950 679.950 328.050 680.550 ;
        RECT 334.950 680.100 337.050 680.550 ;
        RECT 343.950 679.950 349.050 682.050 ;
        RECT 356.400 680.100 357.300 689.400 ;
        RECT 377.700 689.100 378.600 694.200 ;
        RECT 385.950 688.950 388.050 691.050 ;
        RECT 400.500 689.400 402.300 701.400 ;
        RECT 406.950 693.450 409.050 694.050 ;
        RECT 412.950 693.450 415.050 694.050 ;
        RECT 406.950 692.550 415.050 693.450 ;
        RECT 406.950 691.950 409.050 692.550 ;
        RECT 412.950 691.950 415.050 692.550 ;
        RECT 421.500 689.400 423.300 701.400 ;
        RECT 439.800 695.400 441.600 701.400 ;
        RECT 440.700 695.100 441.600 695.400 ;
        RECT 445.800 695.400 447.600 701.400 ;
        RECT 460.800 695.400 462.600 701.400 ;
        RECT 445.800 695.100 447.300 695.400 ;
        RECT 440.700 694.200 447.300 695.100 ;
        RECT 424.950 690.450 427.050 691.050 ;
        RECT 424.950 689.550 432.450 690.450 ;
        RECT 376.950 685.950 379.050 688.050 ;
        RECT 386.100 687.150 387.900 687.900 ;
        RECT 383.100 686.100 384.900 686.850 ;
        RECT 400.950 686.100 402.150 689.400 ;
        RECT 421.950 686.100 423.150 689.400 ;
        RECT 424.950 688.950 427.050 689.550 ;
        RECT 358.950 682.950 361.050 685.050 ;
        RECT 364.950 682.950 367.050 685.050 ;
        RECT 359.100 681.150 360.900 681.900 ;
        RECT 365.100 681.150 366.900 681.900 ;
        RECT 362.100 680.100 363.900 680.850 ;
        RECT 268.950 672.600 270.000 675.900 ;
        RECT 280.950 675.450 283.050 676.050 ;
        RECT 289.950 675.450 292.050 676.050 ;
        RECT 280.950 674.550 292.050 675.450 ;
        RECT 280.950 673.950 283.050 674.550 ;
        RECT 289.950 673.950 292.050 674.550 ;
        RECT 308.100 675.000 312.300 676.650 ;
        RECT 254.400 666.600 256.200 669.600 ;
        RECT 268.200 666.600 270.000 672.600 ;
        RECT 290.400 669.600 291.600 672.900 ;
        RECT 290.400 666.600 292.200 669.600 ;
        RECT 308.100 666.600 309.900 675.000 ;
        RECT 326.400 674.700 327.600 678.900 ;
        RECT 344.400 674.700 345.600 678.900 ;
        RECT 352.950 676.950 358.050 679.050 ;
        RECT 361.950 676.950 364.050 679.050 ;
        RECT 377.700 676.650 378.600 684.900 ;
        RECT 382.950 682.950 385.050 685.200 ;
        RECT 397.950 682.950 400.050 685.050 ;
        RECT 379.950 679.950 382.050 682.050 ;
        RECT 401.100 681.900 402.150 686.100 ;
        RECT 403.950 682.950 406.050 685.050 ;
        RECT 418.950 682.950 421.050 685.050 ;
        RECT 422.100 681.900 423.150 686.100 ;
        RECT 424.950 682.950 427.050 685.050 ;
        RECT 398.100 681.150 399.900 681.900 ;
        RECT 395.100 680.100 396.900 680.850 ;
        RECT 400.950 680.100 402.150 681.900 ;
        RECT 404.100 681.150 405.900 681.900 ;
        RECT 419.100 681.150 420.900 681.900 ;
        RECT 416.100 680.100 417.900 680.850 ;
        RECT 421.950 680.100 423.150 681.900 ;
        RECT 425.100 681.150 426.900 681.900 ;
        RECT 431.550 681.450 432.450 689.550 ;
        RECT 440.700 689.100 441.600 694.200 ;
        RECT 448.950 688.950 454.050 691.050 ;
        RECT 436.950 685.950 442.050 688.050 ;
        RECT 449.100 687.150 450.900 687.900 ;
        RECT 446.100 686.100 447.900 686.850 ;
        RECT 457.950 685.950 460.050 688.050 ;
        RECT 436.950 681.450 439.050 682.050 ;
        RECT 431.550 680.550 439.050 681.450 ;
        RECT 436.950 679.950 439.050 680.550 ;
        RECT 380.100 678.150 381.900 678.900 ;
        RECT 394.950 676.950 397.050 679.050 ;
        RECT 400.950 678.450 403.050 679.050 ;
        RECT 409.950 678.450 412.050 679.050 ;
        RECT 400.950 677.550 412.050 678.450 ;
        RECT 400.950 676.950 403.050 677.550 ;
        RECT 409.950 676.950 412.050 677.550 ;
        RECT 415.950 676.950 418.050 679.050 ;
        RECT 421.950 678.450 424.050 679.050 ;
        RECT 430.950 678.450 433.050 679.050 ;
        RECT 421.950 677.550 433.050 678.450 ;
        RECT 421.950 676.950 424.050 677.550 ;
        RECT 430.950 676.950 433.050 677.550 ;
        RECT 440.700 676.650 441.600 684.900 ;
        RECT 445.950 682.950 448.050 685.200 ;
        RECT 458.100 684.150 459.900 684.900 ;
        RECT 461.400 683.100 462.600 695.400 ;
        RECT 470.400 695.400 472.200 701.400 ;
        RECT 470.400 688.500 471.600 695.400 ;
        RECT 476.700 689.400 478.500 701.400 ;
        RECT 488.400 689.400 490.200 701.400 ;
        RECT 499.500 689.400 501.300 701.400 ;
        RECT 505.800 695.400 507.600 701.400 ;
        RECT 463.950 685.950 466.050 688.050 ;
        RECT 470.400 687.600 476.100 688.500 ;
        RECT 474.150 686.700 476.100 687.600 ;
        RECT 464.100 684.150 465.900 684.900 ;
        RECT 470.100 683.100 471.900 683.850 ;
        RECT 442.950 679.950 445.050 682.050 ;
        RECT 460.950 681.450 463.050 682.050 ;
        RECT 455.550 681.000 463.050 681.450 ;
        RECT 454.950 680.550 463.050 681.000 ;
        RECT 443.100 678.150 444.900 678.900 ;
        RECT 454.950 676.950 457.050 680.550 ;
        RECT 460.950 679.950 463.050 680.550 ;
        RECT 474.150 680.100 475.050 686.700 ;
        RECT 477.000 680.100 478.200 689.400 ;
        RECT 484.950 682.950 487.050 685.200 ;
        RECT 485.100 681.150 486.900 681.900 ;
        RECT 488.400 680.100 489.600 689.400 ;
        RECT 499.800 680.100 501.000 689.400 ;
        RECT 506.400 688.500 507.600 695.400 ;
        RECT 520.500 689.400 522.300 701.400 ;
        RECT 538.800 700.500 546.600 701.400 ;
        RECT 538.800 689.400 540.600 700.500 ;
        RECT 501.900 687.600 507.600 688.500 ;
        RECT 501.900 686.700 503.850 687.600 ;
        RECT 502.950 680.100 503.850 686.700 ;
        RECT 520.950 686.100 522.150 689.400 ;
        RECT 541.800 688.500 543.600 699.600 ;
        RECT 544.800 690.600 546.600 700.500 ;
        RECT 550.800 690.600 552.600 701.400 ;
        RECT 544.800 689.700 552.600 690.600 ;
        RECT 563.400 695.400 565.200 701.400 ;
        RECT 577.800 695.400 579.600 701.400 ;
        RECT 541.800 687.600 545.850 688.500 ;
        RECT 544.950 686.100 545.850 687.600 ;
        RECT 506.100 683.100 507.900 683.850 ;
        RECT 517.950 682.950 520.050 685.050 ;
        RECT 521.100 681.900 522.150 686.100 ;
        RECT 523.950 682.950 526.050 685.050 ;
        RECT 541.950 682.950 544.050 685.200 ;
        RECT 518.100 681.150 519.900 681.900 ;
        RECT 515.100 680.100 516.900 680.850 ;
        RECT 520.950 680.100 522.150 681.900 ;
        RECT 524.100 681.150 525.900 681.900 ;
        RECT 324.000 673.800 327.600 674.700 ;
        RECT 342.000 673.800 345.600 674.700 ;
        RECT 324.000 666.600 325.800 673.800 ;
        RECT 342.000 666.600 343.800 673.800 ;
        RECT 356.400 672.600 357.300 675.900 ;
        RECT 377.700 675.000 381.900 676.650 ;
        RECT 356.400 670.950 361.800 672.600 ;
        RECT 360.000 666.600 361.800 670.950 ;
        RECT 380.100 666.600 381.900 675.000 ;
        RECT 401.850 675.750 403.050 675.900 ;
        RECT 422.850 675.750 424.050 675.900 ;
        RECT 401.850 674.700 405.600 675.750 ;
        RECT 422.850 674.700 426.600 675.750 ;
        RECT 440.700 675.000 444.900 676.650 ;
        RECT 395.400 671.700 403.200 673.050 ;
        RECT 395.400 666.600 397.200 671.700 ;
        RECT 401.400 666.600 403.200 671.700 ;
        RECT 404.400 672.600 405.600 674.700 ;
        RECT 404.400 666.600 406.200 672.600 ;
        RECT 416.400 671.700 424.200 673.050 ;
        RECT 416.400 666.600 418.200 671.700 ;
        RECT 422.400 666.600 424.200 671.700 ;
        RECT 425.400 672.600 426.600 674.700 ;
        RECT 425.400 666.600 427.200 672.600 ;
        RECT 443.100 666.600 444.900 675.000 ;
        RECT 461.400 674.700 462.600 678.900 ;
        RECT 459.000 673.800 462.600 674.700 ;
        RECT 474.150 675.900 474.900 680.100 ;
        RECT 475.950 678.450 478.050 679.050 ;
        RECT 480.000 678.450 484.050 679.050 ;
        RECT 475.950 677.550 484.050 678.450 ;
        RECT 475.950 676.950 478.050 677.550 ;
        RECT 480.000 676.950 484.050 677.550 ;
        RECT 487.950 676.950 490.050 679.050 ;
        RECT 496.950 676.950 502.050 679.050 ;
        RECT 503.100 675.900 503.850 680.100 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 545.100 681.900 545.850 686.100 ;
        RECT 559.950 685.950 562.050 688.050 ;
        RECT 560.100 684.150 561.900 684.900 ;
        RECT 563.400 683.100 564.600 695.400 ;
        RECT 565.950 685.950 568.050 688.050 ;
        RECT 578.400 686.100 579.600 695.400 ;
        RECT 595.500 689.400 597.300 701.400 ;
        RECT 613.800 695.400 615.600 701.400 ;
        RECT 595.950 686.100 597.150 689.400 ;
        RECT 614.400 686.100 615.600 695.400 ;
        RECT 628.500 689.400 630.300 701.400 ;
        RECT 643.800 695.400 645.600 701.400 ;
        RECT 644.700 695.100 645.600 695.400 ;
        RECT 649.800 695.400 651.600 701.400 ;
        RECT 662.400 695.400 664.200 701.400 ;
        RECT 649.800 695.100 651.300 695.400 ;
        RECT 644.700 694.200 651.300 695.100 ;
        RECT 662.700 695.100 664.200 695.400 ;
        RECT 668.400 695.400 670.200 701.400 ;
        RECT 683.400 695.400 685.200 701.400 ;
        RECT 668.400 695.100 669.300 695.400 ;
        RECT 662.700 694.200 669.300 695.100 ;
        RECT 683.700 695.100 685.200 695.400 ;
        RECT 689.400 695.400 691.200 701.400 ;
        RECT 704.400 695.400 706.200 701.400 ;
        RECT 689.400 695.100 690.300 695.400 ;
        RECT 683.700 694.200 690.300 695.100 ;
        RECT 704.700 695.100 706.200 695.400 ;
        RECT 710.400 695.400 712.200 701.400 ;
        RECT 722.400 695.400 724.200 701.400 ;
        RECT 710.400 695.100 711.300 695.400 ;
        RECT 704.700 694.200 711.300 695.100 ;
        RECT 722.700 695.100 724.200 695.400 ;
        RECT 728.400 695.400 730.200 701.400 ;
        RECT 728.400 695.100 729.300 695.400 ;
        RECT 722.700 694.200 729.300 695.100 ;
        RECT 628.950 686.100 630.150 689.400 ;
        RECT 644.700 689.100 645.600 694.200 ;
        RECT 652.950 688.950 655.050 691.050 ;
        RECT 658.950 688.950 661.050 691.050 ;
        RECT 668.400 689.100 669.300 694.200 ;
        RECT 679.950 688.950 682.050 691.050 ;
        RECT 689.400 689.100 690.300 694.200 ;
        RECT 700.950 688.950 703.050 691.050 ;
        RECT 710.400 689.100 711.300 694.200 ;
        RECT 718.950 688.950 721.050 691.050 ;
        RECT 728.400 689.100 729.300 694.200 ;
        RECT 740.400 690.600 742.200 701.400 ;
        RECT 746.400 700.500 754.200 701.400 ;
        RECT 746.400 690.600 748.200 700.500 ;
        RECT 740.400 689.700 748.200 690.600 ;
        RECT 749.400 688.500 751.200 699.600 ;
        RECT 752.400 689.400 754.200 700.500 ;
        RECT 765.600 689.400 767.400 701.400 ;
        RECT 784.500 689.400 786.300 701.400 ;
        RECT 805.800 695.400 807.600 701.400 ;
        RECT 566.100 684.150 567.900 684.900 ;
        RECT 577.950 684.450 580.050 685.050 ;
        RECT 586.950 684.450 589.050 685.050 ;
        RECT 577.950 683.550 589.050 684.450 ;
        RECT 577.950 682.950 580.050 683.550 ;
        RECT 586.950 682.950 589.050 683.550 ;
        RECT 592.950 682.950 595.050 685.050 ;
        RECT 542.250 681.150 544.050 681.900 ;
        RECT 539.100 680.100 540.900 680.850 ;
        RECT 544.950 680.100 545.850 681.900 ;
        RECT 547.950 681.150 549.750 681.900 ;
        RECT 562.950 681.450 565.050 682.050 ;
        RECT 571.950 681.450 574.050 682.050 ;
        RECT 596.100 681.900 597.150 686.100 ;
        RECT 598.950 682.950 601.050 685.050 ;
        RECT 604.950 684.450 607.050 685.050 ;
        RECT 610.950 684.450 616.050 685.050 ;
        RECT 604.950 683.550 616.050 684.450 ;
        RECT 604.950 682.950 607.050 683.550 ;
        RECT 610.950 682.950 616.050 683.550 ;
        RECT 625.950 682.950 628.050 685.050 ;
        RECT 629.100 681.900 630.150 686.100 ;
        RECT 643.950 685.950 646.050 688.050 ;
        RECT 653.100 687.150 654.900 687.900 ;
        RECT 659.100 687.150 660.900 687.900 ;
        RECT 650.100 686.100 651.900 686.850 ;
        RECT 662.100 686.100 663.900 686.850 ;
        RECT 667.950 685.950 673.050 688.050 ;
        RECT 680.100 687.150 681.900 687.900 ;
        RECT 683.100 686.100 684.900 686.850 ;
        RECT 688.950 685.950 694.050 688.050 ;
        RECT 701.100 687.150 702.900 687.900 ;
        RECT 704.100 686.100 705.900 686.850 ;
        RECT 709.950 685.950 715.050 688.050 ;
        RECT 719.100 687.150 720.900 687.900 ;
        RECT 727.950 687.450 730.050 688.050 ;
        RECT 736.950 687.450 739.050 688.050 ;
        RECT 722.100 686.100 723.900 686.850 ;
        RECT 727.950 686.550 739.050 687.450 ;
        RECT 727.950 685.950 730.050 686.550 ;
        RECT 736.950 685.950 739.050 686.550 ;
        RECT 747.150 687.600 751.200 688.500 ;
        RECT 765.600 688.350 768.300 689.400 ;
        RECT 747.150 686.100 748.050 687.600 ;
        RECT 631.950 682.950 634.050 685.200 ;
        RECT 550.950 680.100 552.750 680.850 ;
        RECT 562.950 680.550 574.050 681.450 ;
        RECT 562.950 679.950 565.050 680.550 ;
        RECT 571.950 679.950 574.050 680.550 ;
        RECT 511.950 676.950 517.050 679.050 ;
        RECT 520.950 678.450 523.050 679.050 ;
        RECT 529.950 678.450 532.050 679.050 ;
        RECT 520.950 677.550 532.050 678.450 ;
        RECT 520.950 676.950 523.050 677.550 ;
        RECT 529.950 676.950 532.050 677.550 ;
        RECT 533.550 676.050 534.450 679.950 ;
        RECT 538.950 676.950 541.050 679.050 ;
        RECT 544.950 676.950 547.050 679.050 ;
        RECT 550.950 676.950 553.050 679.050 ;
        RECT 474.150 675.300 475.050 675.900 ;
        RECT 474.150 674.400 476.100 675.300 ;
        RECT 459.000 666.600 460.800 673.800 ;
        RECT 471.000 673.500 476.100 674.400 ;
        RECT 471.000 669.600 472.200 673.500 ;
        RECT 477.000 672.600 478.200 675.900 ;
        RECT 488.400 672.600 489.600 675.900 ;
        RECT 499.800 672.600 501.000 675.900 ;
        RECT 502.950 675.300 503.850 675.900 ;
        RECT 501.900 674.400 503.850 675.300 ;
        RECT 521.850 675.750 523.050 675.900 ;
        RECT 521.850 674.700 525.600 675.750 ;
        RECT 501.900 673.500 507.000 674.400 ;
        RECT 470.400 666.600 472.200 669.600 ;
        RECT 476.700 666.600 478.500 672.600 ;
        RECT 488.400 666.600 490.200 672.600 ;
        RECT 499.500 666.600 501.300 672.600 ;
        RECT 505.800 669.600 507.000 673.500 ;
        RECT 515.400 671.700 523.200 673.050 ;
        RECT 505.800 666.600 507.600 669.600 ;
        RECT 515.400 666.600 517.200 671.700 ;
        RECT 521.400 666.600 523.200 671.700 ;
        RECT 524.400 672.600 525.600 674.700 ;
        RECT 532.950 673.950 535.050 676.050 ;
        RECT 546.000 672.600 547.050 675.900 ;
        RECT 563.400 674.700 564.600 678.900 ;
        RECT 568.950 675.450 571.050 676.200 ;
        RECT 574.950 675.450 577.050 676.050 ;
        RECT 563.400 673.800 567.000 674.700 ;
        RECT 568.950 674.550 577.050 675.450 ;
        RECT 568.950 674.100 571.050 674.550 ;
        RECT 574.950 673.950 577.050 674.550 ;
        RECT 524.400 666.600 526.200 672.600 ;
        RECT 546.000 666.600 547.800 672.600 ;
        RECT 565.200 666.600 567.000 673.800 ;
        RECT 578.400 669.600 579.600 681.900 ;
        RECT 593.100 681.150 594.900 681.900 ;
        RECT 581.100 680.100 582.900 680.850 ;
        RECT 590.100 680.100 591.900 680.850 ;
        RECT 595.950 680.100 597.150 681.900 ;
        RECT 599.100 681.150 600.900 681.900 ;
        RECT 580.950 676.950 583.050 679.050 ;
        RECT 589.950 676.950 592.050 679.050 ;
        RECT 595.950 678.450 598.050 679.050 ;
        RECT 610.950 678.450 613.050 679.050 ;
        RECT 595.950 677.550 613.050 678.450 ;
        RECT 595.950 676.950 598.050 677.550 ;
        RECT 610.950 676.950 613.050 677.550 ;
        RECT 596.850 675.750 598.050 675.900 ;
        RECT 596.850 674.700 600.600 675.750 ;
        RECT 577.800 666.600 579.600 669.600 ;
        RECT 590.400 671.700 598.200 673.050 ;
        RECT 590.400 666.600 592.200 671.700 ;
        RECT 596.400 666.600 598.200 671.700 ;
        RECT 599.400 672.600 600.600 674.700 ;
        RECT 599.400 666.600 601.200 672.600 ;
        RECT 614.400 669.600 615.600 681.900 ;
        RECT 626.100 681.150 627.900 681.900 ;
        RECT 617.100 680.100 618.900 680.850 ;
        RECT 623.100 680.100 624.900 680.850 ;
        RECT 628.950 680.100 630.150 681.900 ;
        RECT 632.100 681.150 633.900 681.900 ;
        RECT 616.950 676.950 619.050 679.050 ;
        RECT 622.950 676.950 625.050 679.050 ;
        RECT 628.950 676.950 634.050 679.050 ;
        RECT 644.700 676.650 645.600 684.900 ;
        RECT 649.950 682.950 652.050 685.050 ;
        RECT 661.950 682.950 664.050 685.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 664.950 679.950 667.050 682.050 ;
        RECT 647.100 678.150 648.900 678.900 ;
        RECT 665.100 678.150 666.900 678.900 ;
        RECT 668.400 676.650 669.300 684.900 ;
        RECT 682.950 682.950 685.050 685.200 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 686.100 678.150 687.900 678.900 ;
        RECT 689.400 676.650 690.300 684.900 ;
        RECT 703.950 682.950 706.050 685.200 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 707.100 678.150 708.900 678.900 ;
        RECT 710.400 676.650 711.300 684.900 ;
        RECT 721.950 682.950 724.050 685.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 725.100 678.150 726.900 678.900 ;
        RECT 728.400 676.650 729.300 684.900 ;
        RECT 742.950 682.950 745.050 685.050 ;
        RECT 747.150 681.900 747.900 686.100 ;
        RECT 748.950 682.950 751.050 685.050 ;
        RECT 764.100 683.100 765.900 683.850 ;
        RECT 766.950 683.100 768.300 688.350 ;
        RECT 770.100 686.100 771.900 686.850 ;
        RECT 784.950 686.100 786.150 689.400 ;
        RECT 743.250 681.150 745.050 681.900 ;
        RECT 740.250 680.100 742.050 680.850 ;
        RECT 747.150 680.100 748.050 681.900 ;
        RECT 748.950 681.150 750.750 681.900 ;
        RECT 752.100 680.100 753.900 680.850 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 739.950 676.950 742.050 679.050 ;
        RECT 745.950 676.950 748.050 679.050 ;
        RECT 751.950 676.950 754.050 679.050 ;
        RECT 767.100 678.900 768.300 683.100 ;
        RECT 769.950 682.950 772.050 685.050 ;
        RECT 781.950 682.950 784.050 685.050 ;
        RECT 785.100 681.900 786.150 686.100 ;
        RECT 802.950 685.950 805.050 688.050 ;
        RECT 787.950 682.950 790.050 685.050 ;
        RECT 803.100 684.150 804.900 684.900 ;
        RECT 806.400 683.100 807.600 695.400 ;
        RECT 815.400 690.300 817.200 701.400 ;
        RECT 821.400 690.300 823.200 701.400 ;
        RECT 815.400 689.400 823.200 690.300 ;
        RECT 824.400 689.400 826.200 701.400 ;
        RECT 808.950 685.950 811.050 688.050 ;
        RECT 809.100 684.150 810.900 684.900 ;
        RECT 814.950 682.950 817.050 685.050 ;
        RECT 820.950 682.950 823.050 685.050 ;
        RECT 782.100 681.150 783.900 681.900 ;
        RECT 779.100 680.100 780.900 680.850 ;
        RECT 784.950 680.100 786.150 681.900 ;
        RECT 788.100 681.150 789.900 681.900 ;
        RECT 793.950 681.450 796.050 682.050 ;
        RECT 805.950 681.450 808.050 682.050 ;
        RECT 793.950 680.550 808.050 681.450 ;
        RECT 815.100 681.150 816.900 681.900 ;
        RECT 821.100 681.150 822.900 681.900 ;
        RECT 793.950 679.950 796.050 680.550 ;
        RECT 805.950 679.950 808.050 680.550 ;
        RECT 818.100 680.100 819.900 680.850 ;
        RECT 824.700 680.100 825.600 689.400 ;
        RECT 766.950 677.100 768.300 678.900 ;
        RECT 778.950 676.950 781.050 679.050 ;
        RECT 784.950 676.950 787.050 679.050 ;
        RECT 629.850 675.750 631.050 675.900 ;
        RECT 629.850 674.700 633.600 675.750 ;
        RECT 644.700 675.000 648.900 676.650 ;
        RECT 613.800 666.600 615.600 669.600 ;
        RECT 623.400 671.700 631.200 673.050 ;
        RECT 623.400 666.600 625.200 671.700 ;
        RECT 629.400 666.600 631.200 671.700 ;
        RECT 632.400 672.600 633.600 674.700 ;
        RECT 632.400 666.600 634.200 672.600 ;
        RECT 647.100 666.600 648.900 675.000 ;
        RECT 665.100 675.000 669.300 676.650 ;
        RECT 686.100 675.000 690.300 676.650 ;
        RECT 707.100 675.000 711.300 676.650 ;
        RECT 725.100 675.000 729.300 676.650 ;
        RECT 665.100 666.600 666.900 675.000 ;
        RECT 686.100 666.600 687.900 675.000 ;
        RECT 707.100 666.600 708.900 675.000 ;
        RECT 725.100 666.600 726.900 675.000 ;
        RECT 745.950 672.600 747.000 675.900 ;
        RECT 766.950 675.450 769.050 676.050 ;
        RECT 758.550 674.550 769.050 675.450 ;
        RECT 785.850 675.750 787.050 675.900 ;
        RECT 785.850 674.700 789.600 675.750 ;
        RECT 806.400 674.700 807.600 678.900 ;
        RECT 817.950 676.950 820.050 679.050 ;
        RECT 823.950 676.950 826.050 679.050 ;
        RECT 758.550 673.050 759.450 674.550 ;
        RECT 766.950 673.950 769.050 674.550 ;
        RECT 745.200 666.600 747.000 672.600 ;
        RECT 754.950 671.550 759.450 673.050 ;
        RECT 754.950 670.950 759.000 671.550 ;
        RECT 767.400 669.600 768.600 672.900 ;
        RECT 766.800 666.600 768.600 669.600 ;
        RECT 779.400 671.700 787.200 673.050 ;
        RECT 779.400 666.600 781.200 671.700 ;
        RECT 785.400 666.600 787.200 671.700 ;
        RECT 788.400 672.600 789.600 674.700 ;
        RECT 804.000 673.800 807.600 674.700 ;
        RECT 788.400 666.600 790.200 672.600 ;
        RECT 804.000 666.600 805.800 673.800 ;
        RECT 824.700 672.600 825.600 675.900 ;
        RECT 820.200 670.950 825.600 672.600 ;
        RECT 820.200 666.600 822.000 670.950 ;
        RECT 12.000 655.200 13.800 662.400 ;
        RECT 12.000 654.300 15.600 655.200 ;
        RECT 14.400 650.100 15.600 654.300 ;
        RECT 32.100 654.000 33.900 662.400 ;
        RECT 29.700 652.350 33.900 654.000 ;
        RECT 53.100 654.000 54.900 662.400 ;
        RECT 68.400 659.400 70.200 662.400 ;
        RECT 53.100 652.350 57.300 654.000 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 11.100 644.100 12.900 644.850 ;
        RECT 7.950 640.950 13.050 643.050 ;
        RECT 14.400 633.600 15.600 645.900 ;
        RECT 17.100 644.100 18.900 644.850 ;
        RECT 29.700 644.100 30.600 652.350 ;
        RECT 32.100 650.100 33.900 650.850 ;
        RECT 53.100 650.100 54.900 650.850 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 52.950 646.950 55.050 649.200 ;
        RECT 34.950 643.950 37.050 646.050 ;
        RECT 49.950 643.950 52.050 646.050 ;
        RECT 56.400 644.100 57.300 652.350 ;
        RECT 64.950 649.950 67.050 652.050 ;
        RECT 65.100 648.150 66.900 648.900 ;
        RECT 68.400 647.100 69.600 659.400 ;
        RECT 85.200 658.050 87.000 662.400 ;
        RECT 103.800 659.400 105.600 662.400 ;
        RECT 85.200 656.400 90.600 658.050 ;
        RECT 89.700 653.100 90.600 656.400 ;
        RECT 70.950 651.450 73.050 652.050 ;
        RECT 82.950 651.450 85.050 652.050 ;
        RECT 70.950 650.550 85.050 651.450 ;
        RECT 70.950 649.950 73.050 650.550 ;
        RECT 82.950 649.950 85.050 650.550 ;
        RECT 88.950 651.450 91.050 652.050 ;
        RECT 93.000 651.450 97.050 652.050 ;
        RECT 88.950 650.550 97.050 651.450 ;
        RECT 88.950 649.950 91.050 650.550 ;
        RECT 93.000 649.950 97.050 650.550 ;
        RECT 83.100 648.150 84.900 648.900 ;
        RECT 80.100 647.100 81.900 647.850 ;
        RECT 86.100 647.100 87.900 647.850 ;
        RECT 67.950 643.950 73.050 646.050 ;
        RECT 76.950 643.950 82.050 646.050 ;
        RECT 85.950 643.950 88.050 646.050 ;
        RECT 16.950 640.950 19.050 643.050 ;
        RECT 22.950 642.450 27.000 643.050 ;
        RECT 28.950 642.450 31.050 643.050 ;
        RECT 22.950 641.550 31.050 642.450 ;
        RECT 35.100 642.150 36.900 642.900 ;
        RECT 50.100 642.150 51.900 642.900 ;
        RECT 22.950 640.950 27.000 641.550 ;
        RECT 28.950 640.950 31.050 641.550 ;
        RECT 38.100 641.100 39.900 641.850 ;
        RECT 47.100 641.100 48.900 641.850 ;
        RECT 55.950 640.950 58.050 643.050 ;
        RECT 29.700 634.800 30.600 639.900 ;
        RECT 37.950 637.950 40.050 640.050 ;
        RECT 46.950 637.950 52.050 640.050 ;
        RECT 56.400 634.800 57.300 639.900 ;
        RECT 29.700 633.900 36.300 634.800 ;
        RECT 29.700 633.600 30.600 633.900 ;
        RECT 13.800 627.600 15.600 633.600 ;
        RECT 28.800 627.600 30.600 633.600 ;
        RECT 34.800 633.600 36.300 633.900 ;
        RECT 50.700 633.900 57.300 634.800 ;
        RECT 50.700 633.600 52.200 633.900 ;
        RECT 34.800 627.600 36.600 633.600 ;
        RECT 50.400 627.600 52.200 633.600 ;
        RECT 56.400 633.600 57.300 633.900 ;
        RECT 68.400 633.600 69.600 642.900 ;
        RECT 89.700 639.600 90.600 648.900 ;
        RECT 104.400 647.100 105.600 659.400 ;
        RECT 118.800 656.400 120.600 662.400 ;
        RECT 119.400 654.300 120.600 656.400 ;
        RECT 121.800 657.300 123.600 662.400 ;
        RECT 127.800 657.300 129.600 662.400 ;
        RECT 142.800 659.400 144.600 662.400 ;
        RECT 121.800 655.950 129.600 657.300 ;
        RECT 143.400 656.100 144.600 659.400 ;
        RECT 156.000 655.200 157.800 662.400 ;
        RECT 171.000 655.200 172.800 662.400 ;
        RECT 187.500 656.400 189.300 662.400 ;
        RECT 193.800 659.400 195.600 662.400 ;
        RECT 136.950 654.450 141.000 655.050 ;
        RECT 142.950 654.450 145.050 655.050 ;
        RECT 119.400 653.250 123.150 654.300 ;
        RECT 121.950 653.100 123.150 653.250 ;
        RECT 136.950 653.550 145.050 654.450 ;
        RECT 156.000 654.300 159.600 655.200 ;
        RECT 171.000 654.300 174.600 655.200 ;
        RECT 136.950 652.950 141.000 653.550 ;
        RECT 142.950 652.950 145.050 653.550 ;
        RECT 106.950 649.950 109.050 652.050 ;
        RECT 121.950 649.950 124.050 652.050 ;
        RECT 127.950 649.800 130.050 652.050 ;
        RECT 142.950 650.100 144.300 651.900 ;
        RECT 158.400 650.100 159.600 654.300 ;
        RECT 173.400 650.100 174.600 654.300 ;
        RECT 187.800 653.100 189.000 656.400 ;
        RECT 193.800 655.500 195.000 659.400 ;
        RECT 205.800 656.400 207.600 662.400 ;
        RECT 189.900 654.600 195.000 655.500 ;
        RECT 189.900 653.700 191.850 654.600 ;
        RECT 190.950 653.100 191.850 653.700 ;
        RECT 206.400 654.300 207.600 656.400 ;
        RECT 208.800 657.300 210.600 662.400 ;
        RECT 214.800 657.300 216.600 662.400 ;
        RECT 208.800 655.950 216.600 657.300 ;
        RECT 226.800 656.400 228.600 662.400 ;
        RECT 227.400 654.300 228.600 656.400 ;
        RECT 229.800 657.300 231.600 662.400 ;
        RECT 235.800 657.300 237.600 662.400 ;
        RECT 229.800 655.950 237.600 657.300 ;
        RECT 244.800 656.400 246.600 662.400 ;
        RECT 245.400 654.300 246.600 656.400 ;
        RECT 247.800 657.300 249.600 662.400 ;
        RECT 253.800 657.300 255.600 662.400 ;
        RECT 247.800 655.950 255.600 657.300 ;
        RECT 267.000 655.200 268.800 662.400 ;
        RECT 283.800 656.400 285.600 662.400 ;
        RECT 267.000 654.300 270.600 655.200 ;
        RECT 206.400 653.250 210.150 654.300 ;
        RECT 227.400 653.250 231.150 654.300 ;
        RECT 245.400 653.250 249.150 654.300 ;
        RECT 208.950 653.100 210.150 653.250 ;
        RECT 229.950 653.100 231.150 653.250 ;
        RECT 247.950 653.100 249.150 653.250 ;
        RECT 107.100 648.150 108.900 648.900 ;
        RECT 119.100 647.100 120.900 647.850 ;
        RECT 122.850 647.100 124.050 648.900 ;
        RECT 128.100 648.150 129.900 648.900 ;
        RECT 125.100 647.100 126.900 647.850 ;
        RECT 100.950 643.950 106.050 646.050 ;
        RECT 118.950 643.950 121.050 646.050 ;
        RECT 122.850 642.900 123.900 647.100 ;
        RECT 139.950 646.950 142.050 649.050 ;
        RECT 124.950 643.950 127.050 646.050 ;
        RECT 143.100 645.900 144.300 650.100 ;
        RECT 184.950 649.950 190.050 652.050 ;
        RECT 151.950 648.450 156.000 649.050 ;
        RECT 157.950 648.450 160.050 649.050 ;
        RECT 151.950 647.550 160.050 648.450 ;
        RECT 151.950 646.950 156.000 647.550 ;
        RECT 157.950 646.950 160.050 647.550 ;
        RECT 172.950 648.450 175.050 649.050 ;
        RECT 181.950 648.450 184.050 649.050 ;
        RECT 191.100 648.900 191.850 653.100 ;
        RECT 204.000 651.900 207.000 652.050 ;
        RECT 202.950 651.450 207.000 651.900 ;
        RECT 208.950 651.450 211.050 652.050 ;
        RECT 202.950 650.550 211.050 651.450 ;
        RECT 202.950 649.950 207.000 650.550 ;
        RECT 208.950 649.950 211.050 650.550 ;
        RECT 214.950 649.950 217.050 652.050 ;
        RECT 229.950 649.950 232.050 652.050 ;
        RECT 235.950 649.950 238.050 652.050 ;
        RECT 247.950 649.950 250.050 652.050 ;
        RECT 253.950 649.950 259.050 652.050 ;
        RECT 269.400 650.100 270.600 654.300 ;
        RECT 284.400 654.300 285.600 656.400 ;
        RECT 286.800 657.300 288.600 662.400 ;
        RECT 292.800 657.300 294.600 662.400 ;
        RECT 286.800 655.950 294.600 657.300 ;
        RECT 305.400 659.400 307.200 662.400 ;
        RECT 284.400 653.250 288.150 654.300 ;
        RECT 286.950 653.100 288.150 653.250 ;
        RECT 286.950 649.950 289.050 652.050 ;
        RECT 292.950 649.950 295.050 652.050 ;
        RECT 301.950 649.950 304.050 652.050 ;
        RECT 202.950 649.800 205.050 649.950 ;
        RECT 172.950 647.550 184.050 648.450 ;
        RECT 172.950 646.950 175.050 647.550 ;
        RECT 181.950 646.950 184.050 647.550 ;
        RECT 140.100 645.150 141.900 645.900 ;
        RECT 80.400 638.700 88.200 639.600 ;
        RECT 56.400 627.600 58.200 633.600 ;
        RECT 68.400 627.600 70.200 633.600 ;
        RECT 80.400 627.600 82.200 638.700 ;
        RECT 86.400 627.600 88.200 638.700 ;
        RECT 89.400 627.600 91.200 639.600 ;
        RECT 104.400 633.600 105.600 642.900 ;
        RECT 122.850 639.600 124.050 642.900 ;
        RECT 142.950 640.650 144.300 645.900 ;
        RECT 145.950 643.800 148.050 646.050 ;
        RECT 155.100 644.100 156.900 644.850 ;
        RECT 146.100 642.150 147.900 642.900 ;
        RECT 141.600 639.600 144.300 640.650 ;
        RECT 103.800 627.600 105.600 633.600 ;
        RECT 122.700 627.600 124.500 639.600 ;
        RECT 141.600 627.600 143.400 639.600 ;
        RECT 158.400 633.600 159.600 645.900 ;
        RECT 161.100 644.100 162.900 644.850 ;
        RECT 170.100 644.100 171.900 644.850 ;
        RECT 160.950 640.950 163.050 643.050 ;
        RECT 169.950 640.950 172.050 643.050 ;
        RECT 173.400 633.600 174.600 645.900 ;
        RECT 176.100 644.100 177.900 644.850 ;
        RECT 175.950 640.950 178.050 643.050 ;
        RECT 187.800 639.600 189.000 648.900 ;
        RECT 190.950 642.300 191.850 648.900 ;
        RECT 206.100 647.100 207.900 647.850 ;
        RECT 209.850 647.100 211.050 648.900 ;
        RECT 215.100 648.150 216.900 648.900 ;
        RECT 212.100 647.100 213.900 647.850 ;
        RECT 227.100 647.100 228.900 647.850 ;
        RECT 230.850 647.100 232.050 648.900 ;
        RECT 236.100 648.150 237.900 648.900 ;
        RECT 233.100 647.100 234.900 647.850 ;
        RECT 245.100 647.100 246.900 647.850 ;
        RECT 248.850 647.100 250.050 648.900 ;
        RECT 254.100 648.150 255.900 648.900 ;
        RECT 268.950 648.450 271.050 649.050 ;
        RECT 277.950 648.450 280.050 649.050 ;
        RECT 251.100 647.100 252.900 647.850 ;
        RECT 268.950 647.550 280.050 648.450 ;
        RECT 194.100 645.150 195.900 645.900 ;
        RECT 205.950 643.950 208.050 646.050 ;
        RECT 189.900 641.400 191.850 642.300 ;
        RECT 209.850 642.900 210.900 647.100 ;
        RECT 211.950 643.950 214.050 646.050 ;
        RECT 226.950 643.950 229.050 646.050 ;
        RECT 230.850 642.900 231.900 647.100 ;
        RECT 232.950 643.950 235.050 646.050 ;
        RECT 241.950 643.950 247.050 646.050 ;
        RECT 189.900 640.500 195.600 641.400 ;
        RECT 157.800 627.600 159.600 633.600 ;
        RECT 172.800 627.600 174.600 633.600 ;
        RECT 187.500 627.600 189.300 639.600 ;
        RECT 194.400 633.600 195.600 640.500 ;
        RECT 209.850 639.600 211.050 642.900 ;
        RECT 230.850 639.600 232.050 642.900 ;
        RECT 244.950 640.950 247.050 643.950 ;
        RECT 248.850 642.900 249.900 647.100 ;
        RECT 268.950 646.950 271.050 647.550 ;
        RECT 277.950 646.950 280.050 647.550 ;
        RECT 284.100 647.100 285.900 647.850 ;
        RECT 287.850 647.100 289.050 648.900 ;
        RECT 293.100 648.150 294.900 648.900 ;
        RECT 302.100 648.150 303.900 648.900 ;
        RECT 290.100 647.100 291.900 647.850 ;
        RECT 305.400 647.100 306.600 659.400 ;
        RECT 320.100 654.000 321.900 662.400 ;
        RECT 337.800 659.400 339.600 662.400 ;
        RECT 320.100 652.350 324.300 654.000 ;
        RECT 320.100 650.100 321.900 650.850 ;
        RECT 250.950 643.950 253.050 646.050 ;
        RECT 266.100 644.100 267.900 644.850 ;
        RECT 248.850 639.600 250.050 642.900 ;
        RECT 193.800 627.600 195.600 633.600 ;
        RECT 209.700 627.600 211.500 639.600 ;
        RECT 230.700 627.600 232.500 639.600 ;
        RECT 248.700 627.600 250.500 639.600 ;
        RECT 269.400 633.600 270.600 645.900 ;
        RECT 272.100 644.100 273.900 644.850 ;
        RECT 283.950 643.950 286.050 646.050 ;
        RECT 271.950 642.450 274.050 643.050 ;
        RECT 276.000 642.900 279.000 643.050 ;
        RECT 287.850 642.900 288.900 647.100 ;
        RECT 319.950 646.950 322.050 649.200 ;
        RECT 289.950 643.950 292.050 646.050 ;
        RECT 304.950 643.950 307.050 646.050 ;
        RECT 316.950 643.950 319.050 646.050 ;
        RECT 323.400 644.100 324.300 652.350 ;
        RECT 328.950 645.450 331.050 649.050 ;
        RECT 338.400 647.100 339.600 659.400 ;
        RECT 352.200 655.200 354.000 662.400 ;
        RECT 364.800 656.400 366.600 662.400 ;
        RECT 350.400 654.300 354.000 655.200 ;
        RECT 340.950 649.950 343.050 652.200 ;
        RECT 350.400 650.100 351.600 654.300 ;
        RECT 365.400 653.100 366.600 656.400 ;
        RECT 378.000 655.200 379.800 662.400 ;
        RECT 394.800 659.400 396.600 662.400 ;
        RECT 378.000 654.300 381.600 655.200 ;
        RECT 364.950 649.950 367.050 652.050 ;
        RECT 380.400 650.100 381.600 654.300 ;
        RECT 341.100 648.150 342.900 648.900 ;
        RECT 349.950 646.950 355.050 649.050 ;
        RECT 337.950 645.450 340.050 646.050 ;
        RECT 328.950 645.000 340.050 645.450 ;
        RECT 329.550 644.550 340.050 645.000 ;
        RECT 337.950 643.950 340.050 644.550 ;
        RECT 347.100 644.100 348.900 644.850 ;
        RECT 276.000 642.450 280.050 642.900 ;
        RECT 271.950 641.550 280.050 642.450 ;
        RECT 271.950 640.950 274.050 641.550 ;
        RECT 276.000 640.950 280.050 641.550 ;
        RECT 277.950 640.800 280.050 640.950 ;
        RECT 287.850 639.600 289.050 642.900 ;
        RECT 268.800 627.600 270.600 633.600 ;
        RECT 287.700 627.600 289.500 639.600 ;
        RECT 305.400 633.600 306.600 642.900 ;
        RECT 317.100 642.150 318.900 642.900 ;
        RECT 322.950 642.450 325.050 643.050 ;
        RECT 331.950 642.450 334.050 643.050 ;
        RECT 314.100 641.100 315.900 641.850 ;
        RECT 322.950 641.550 334.050 642.450 ;
        RECT 322.950 640.950 325.050 641.550 ;
        RECT 331.950 640.950 334.050 641.550 ;
        RECT 313.950 637.950 316.050 640.050 ;
        RECT 323.400 634.800 324.300 639.900 ;
        RECT 317.700 633.900 324.300 634.800 ;
        RECT 317.700 633.600 319.200 633.900 ;
        RECT 305.400 627.600 307.200 633.600 ;
        RECT 317.400 627.600 319.200 633.600 ;
        RECT 323.400 633.600 324.300 633.900 ;
        RECT 338.400 633.600 339.600 642.900 ;
        RECT 346.950 637.950 349.050 643.050 ;
        RECT 323.400 627.600 325.200 633.600 ;
        RECT 337.800 627.600 339.600 633.600 ;
        RECT 350.400 633.600 351.600 645.900 ;
        RECT 353.100 644.100 354.900 644.850 ;
        RECT 365.400 639.600 366.600 648.900 ;
        RECT 379.950 648.450 382.050 649.050 ;
        RECT 388.950 648.450 391.050 649.050 ;
        RECT 368.100 647.100 369.900 647.850 ;
        RECT 379.950 647.550 391.050 648.450 ;
        RECT 379.950 646.950 382.050 647.550 ;
        RECT 388.950 646.950 391.050 647.550 ;
        RECT 395.400 647.100 396.600 659.400 ;
        RECT 413.100 654.000 414.900 662.400 ;
        RECT 434.100 654.000 435.900 662.400 ;
        RECT 451.200 655.200 453.000 662.400 ;
        RECT 413.100 652.350 417.300 654.000 ;
        RECT 397.950 651.450 400.050 652.050 ;
        RECT 406.950 651.450 409.050 652.050 ;
        RECT 397.950 650.550 409.050 651.450 ;
        RECT 397.950 649.950 400.050 650.550 ;
        RECT 406.950 649.950 409.050 650.550 ;
        RECT 413.100 650.100 414.900 650.850 ;
        RECT 398.100 648.150 399.900 648.900 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 367.950 643.950 370.050 646.050 ;
        RECT 377.100 644.100 378.900 644.850 ;
        RECT 350.400 627.600 352.200 633.600 ;
        RECT 364.800 627.600 366.600 639.600 ;
        RECT 380.400 633.600 381.600 645.900 ;
        RECT 394.950 645.450 397.050 646.050 ;
        RECT 403.950 645.450 406.050 646.050 ;
        RECT 383.100 644.100 384.900 644.850 ;
        RECT 394.950 644.550 406.050 645.450 ;
        RECT 394.950 643.950 397.050 644.550 ;
        RECT 403.950 643.950 406.050 644.550 ;
        RECT 409.950 643.950 412.050 646.050 ;
        RECT 416.400 644.100 417.300 652.350 ;
        RECT 431.700 652.350 435.900 654.000 ;
        RECT 449.400 654.300 453.000 655.200 ;
        RECT 474.000 656.400 475.800 662.400 ;
        RECT 490.800 659.400 492.600 662.400 ;
        RECT 431.700 644.100 432.600 652.350 ;
        RECT 434.100 650.100 435.900 650.850 ;
        RECT 449.400 650.100 450.600 654.300 ;
        RECT 474.000 653.100 475.050 656.400 ;
        RECT 466.950 649.950 469.050 652.050 ;
        RECT 472.950 649.950 475.050 652.050 ;
        RECT 478.950 649.950 481.050 652.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 448.950 648.450 451.050 649.050 ;
        RECT 460.950 648.450 463.050 649.050 ;
        RECT 448.950 647.550 463.050 648.450 ;
        RECT 467.100 648.150 468.900 648.900 ;
        RECT 448.950 646.950 451.050 647.550 ;
        RECT 460.950 646.950 463.050 647.550 ;
        RECT 470.250 647.100 472.050 647.850 ;
        RECT 472.950 647.100 473.850 648.900 ;
        RECT 478.950 648.150 480.750 648.900 ;
        RECT 475.950 647.100 477.750 647.850 ;
        RECT 491.400 647.100 492.600 659.400 ;
        RECT 503.400 659.400 505.200 662.400 ;
        RECT 514.800 661.500 522.600 662.400 ;
        RECT 493.950 649.950 496.050 652.050 ;
        RECT 499.950 649.950 502.050 652.050 ;
        RECT 494.100 648.150 495.900 648.900 ;
        RECT 500.100 648.150 501.900 648.900 ;
        RECT 503.400 647.100 504.600 659.400 ;
        RECT 514.800 656.400 516.600 661.500 ;
        RECT 517.800 656.400 519.600 660.600 ;
        RECT 520.800 657.000 522.600 661.500 ;
        RECT 526.800 657.000 528.600 662.400 ;
        RECT 514.950 649.950 517.050 655.050 ;
        RECT 518.400 654.900 519.300 656.400 ;
        RECT 520.800 656.100 528.600 657.000 ;
        RECT 539.400 659.400 541.200 662.400 ;
        RECT 539.400 656.100 540.600 659.400 ;
        RECT 556.200 658.050 558.000 662.400 ;
        RECT 556.200 656.400 561.600 658.050 ;
        RECT 518.400 653.700 522.600 654.900 ;
        RECT 538.950 654.450 541.050 655.050 ;
        RECT 547.950 654.450 550.050 655.050 ;
        RECT 521.400 653.100 522.600 653.700 ;
        RECT 526.950 653.100 528.750 653.850 ;
        RECT 538.950 653.550 550.050 654.450 ;
        RECT 538.950 652.950 541.050 653.550 ;
        RECT 547.950 652.950 550.050 653.550 ;
        RECT 560.700 653.100 561.600 656.400 ;
        RECT 578.100 654.000 579.900 662.400 ;
        RECT 595.200 655.200 597.000 662.400 ;
        RECT 608.400 657.300 610.200 662.400 ;
        RECT 614.400 657.300 616.200 662.400 ;
        RECT 608.400 655.950 616.200 657.300 ;
        RECT 617.400 656.400 619.200 662.400 ;
        RECT 629.400 659.400 631.200 662.400 ;
        RECT 593.400 654.300 597.000 655.200 ;
        RECT 617.400 654.300 618.600 656.400 ;
        RECT 578.100 652.350 582.300 654.000 ;
        RECT 520.950 649.950 523.050 652.050 ;
        RECT 526.950 649.950 529.050 652.050 ;
        RECT 539.700 650.100 541.050 651.900 ;
        RECT 436.950 643.950 439.050 646.050 ;
        RECT 446.100 644.100 447.900 644.850 ;
        RECT 382.950 640.950 385.050 643.050 ;
        RECT 395.400 633.600 396.600 642.900 ;
        RECT 410.100 642.150 411.900 642.900 ;
        RECT 415.950 642.450 418.050 643.050 ;
        RECT 424.950 642.450 427.050 643.050 ;
        RECT 407.100 641.100 408.900 641.850 ;
        RECT 415.950 641.550 427.050 642.450 ;
        RECT 415.950 640.950 418.050 641.550 ;
        RECT 424.950 640.950 427.050 641.550 ;
        RECT 430.950 640.950 433.050 643.050 ;
        RECT 437.100 642.150 438.900 642.900 ;
        RECT 440.100 641.100 441.900 641.850 ;
        RECT 445.950 640.950 448.050 643.050 ;
        RECT 406.950 637.950 409.050 640.050 ;
        RECT 416.400 634.800 417.300 639.900 ;
        RECT 410.700 633.900 417.300 634.800 ;
        RECT 410.700 633.600 412.200 633.900 ;
        RECT 379.800 627.600 381.600 633.600 ;
        RECT 394.800 627.600 396.600 633.600 ;
        RECT 410.400 627.600 412.200 633.600 ;
        RECT 416.400 633.600 417.300 633.900 ;
        RECT 431.700 634.800 432.600 639.900 ;
        RECT 439.950 637.950 442.050 640.050 ;
        RECT 431.700 633.900 438.300 634.800 ;
        RECT 431.700 633.600 432.600 633.900 ;
        RECT 416.400 627.600 418.200 633.600 ;
        RECT 430.800 627.600 432.600 633.600 ;
        RECT 436.800 633.600 438.300 633.900 ;
        RECT 449.400 633.600 450.600 645.900 ;
        RECT 452.100 644.100 453.900 644.850 ;
        RECT 451.950 640.950 454.050 643.050 ;
        RECT 473.100 642.900 473.850 647.100 ;
        RECT 490.950 643.950 493.050 646.050 ;
        RECT 502.950 645.450 505.050 646.050 ;
        RECT 508.950 645.450 511.050 649.050 ;
        RECT 515.250 648.150 517.050 648.900 ;
        RECT 518.700 647.100 520.500 647.850 ;
        RECT 502.950 645.000 511.050 645.450 ;
        RECT 502.950 644.550 510.450 645.000 ;
        RECT 502.950 643.950 505.050 644.550 ;
        RECT 517.950 643.950 520.050 646.050 ;
        RECT 472.950 641.400 473.850 642.900 ;
        RECT 469.800 640.500 473.850 641.400 ;
        RECT 436.800 627.600 438.600 633.600 ;
        RECT 449.400 627.600 451.200 633.600 ;
        RECT 466.800 628.500 468.600 639.600 ;
        RECT 469.800 629.400 471.600 640.500 ;
        RECT 472.800 638.400 480.600 639.300 ;
        RECT 472.800 628.500 474.600 638.400 ;
        RECT 466.800 627.600 474.600 628.500 ;
        RECT 478.800 627.600 480.600 638.400 ;
        RECT 491.400 633.600 492.600 642.900 ;
        RECT 490.800 627.600 492.600 633.600 ;
        RECT 503.400 633.600 504.600 642.900 ;
        RECT 521.400 639.600 522.600 648.900 ;
        RECT 524.100 647.100 525.900 647.850 ;
        RECT 523.950 643.950 526.050 646.050 ;
        RECT 535.950 643.950 538.050 646.050 ;
        RECT 539.700 645.900 540.900 650.100 ;
        RECT 553.950 649.950 556.050 652.050 ;
        RECT 559.950 651.450 562.050 652.050 ;
        RECT 571.950 651.450 574.050 652.050 ;
        RECT 559.950 650.550 574.050 651.450 ;
        RECT 559.950 649.950 562.050 650.550 ;
        RECT 571.950 649.950 574.050 650.550 ;
        RECT 578.100 650.100 579.900 650.850 ;
        RECT 541.950 646.950 544.050 649.050 ;
        RECT 554.100 648.150 555.900 648.900 ;
        RECT 551.100 647.100 552.900 647.850 ;
        RECT 557.100 647.100 558.900 647.850 ;
        RECT 536.100 642.150 537.900 642.900 ;
        RECT 539.700 640.650 541.050 645.900 ;
        RECT 542.100 645.150 543.900 645.900 ;
        RECT 550.950 643.950 553.050 646.050 ;
        RECT 556.950 643.950 559.050 646.050 ;
        RECT 539.700 639.600 542.400 640.650 ;
        RECT 560.700 639.600 561.600 648.900 ;
        RECT 577.950 646.950 580.050 649.050 ;
        RECT 574.950 643.950 577.050 646.050 ;
        RECT 581.400 644.100 582.300 652.350 ;
        RECT 593.400 650.100 594.600 654.300 ;
        RECT 614.850 653.250 618.600 654.300 ;
        RECT 614.850 653.100 616.050 653.250 ;
        RECT 607.950 649.950 610.050 652.050 ;
        RECT 613.950 649.950 616.050 652.050 ;
        RECT 625.950 649.950 628.050 652.050 ;
        RECT 592.950 646.950 595.050 649.050 ;
        RECT 608.100 648.150 609.900 648.900 ;
        RECT 611.100 647.100 612.900 647.850 ;
        RECT 613.950 647.100 615.150 648.900 ;
        RECT 626.100 648.150 627.900 648.900 ;
        RECT 617.100 647.100 618.900 647.850 ;
        RECT 629.400 647.100 630.600 659.400 ;
        RECT 646.200 655.200 648.000 662.400 ;
        RECT 661.800 659.400 663.600 662.400 ;
        RECT 644.400 654.300 648.000 655.200 ;
        RECT 644.400 650.100 645.600 654.300 ;
        RECT 634.950 648.450 637.050 649.050 ;
        RECT 643.950 648.450 646.050 649.050 ;
        RECT 634.950 647.550 646.050 648.450 ;
        RECT 590.100 644.100 591.900 644.850 ;
        RECT 575.100 642.150 576.900 642.900 ;
        RECT 572.100 641.100 573.900 641.850 ;
        RECT 580.950 640.950 586.050 643.050 ;
        RECT 589.950 640.950 592.050 643.050 ;
        RECT 503.400 627.600 505.200 633.600 ;
        RECT 520.800 627.600 524.100 639.600 ;
        RECT 540.600 627.600 542.400 639.600 ;
        RECT 551.400 638.700 559.200 639.600 ;
        RECT 551.400 627.600 553.200 638.700 ;
        RECT 557.400 627.600 559.200 638.700 ;
        RECT 560.400 627.600 562.200 639.600 ;
        RECT 571.950 637.950 574.050 640.050 ;
        RECT 581.400 634.800 582.300 639.900 ;
        RECT 575.700 633.900 582.300 634.800 ;
        RECT 575.700 633.600 577.200 633.900 ;
        RECT 575.400 627.600 577.200 633.600 ;
        RECT 581.400 633.600 582.300 633.900 ;
        RECT 593.400 633.600 594.600 645.900 ;
        RECT 596.100 644.100 597.900 644.850 ;
        RECT 610.950 643.950 613.050 646.050 ;
        RECT 614.100 642.900 615.150 647.100 ;
        RECT 634.950 646.950 637.050 647.550 ;
        RECT 643.950 646.950 646.050 647.550 ;
        RECT 662.400 647.100 663.600 659.400 ;
        RECT 674.400 657.300 676.200 662.400 ;
        RECT 680.400 657.300 682.200 662.400 ;
        RECT 674.400 655.950 682.200 657.300 ;
        RECT 683.400 656.400 685.200 662.400 ;
        RECT 692.400 657.300 694.200 662.400 ;
        RECT 698.400 657.300 700.200 662.400 ;
        RECT 683.400 654.300 684.600 656.400 ;
        RECT 692.400 655.950 700.200 657.300 ;
        RECT 701.400 656.400 703.200 662.400 ;
        RECT 715.800 659.400 717.600 662.400 ;
        RECT 701.400 654.300 702.600 656.400 ;
        RECT 680.850 653.250 684.600 654.300 ;
        RECT 698.850 653.250 702.600 654.300 ;
        RECT 680.850 653.100 682.050 653.250 ;
        RECT 698.850 653.100 700.050 653.250 ;
        RECT 664.950 649.950 667.050 652.050 ;
        RECT 673.950 649.950 676.050 652.050 ;
        RECT 679.950 649.950 682.050 652.050 ;
        RECT 691.950 649.950 694.050 652.050 ;
        RECT 697.950 651.450 700.050 652.050 ;
        RECT 712.950 651.450 715.050 652.050 ;
        RECT 697.950 650.550 715.050 651.450 ;
        RECT 697.950 649.950 700.050 650.550 ;
        RECT 712.950 649.950 715.050 650.550 ;
        RECT 665.100 648.150 666.900 648.900 ;
        RECT 674.100 648.150 675.900 648.900 ;
        RECT 677.100 647.100 678.900 647.850 ;
        RECT 679.950 647.100 681.150 648.900 ;
        RECT 692.100 648.150 693.900 648.900 ;
        RECT 683.100 647.100 684.900 647.850 ;
        RECT 695.100 647.100 696.900 647.850 ;
        RECT 697.950 647.100 699.150 648.900 ;
        RECT 701.100 647.100 702.900 647.850 ;
        RECT 716.400 647.100 717.600 659.400 ;
        RECT 734.100 654.000 735.900 662.400 ;
        RECT 755.100 654.000 756.900 662.400 ;
        RECT 771.000 655.200 772.800 662.400 ;
        RECT 787.800 659.400 789.600 662.400 ;
        RECT 788.400 656.100 789.600 659.400 ;
        RECT 801.000 655.200 802.800 662.400 ;
        RECT 771.000 654.300 774.600 655.200 ;
        RECT 734.100 652.350 738.300 654.000 ;
        RECT 718.950 649.950 721.050 652.050 ;
        RECT 734.100 650.100 735.900 650.850 ;
        RECT 719.100 648.150 720.900 648.900 ;
        RECT 616.950 643.950 619.050 646.050 ;
        RECT 628.950 643.950 634.050 646.050 ;
        RECT 641.100 644.100 642.900 644.850 ;
        RECT 613.950 639.600 615.150 642.900 ;
        RECT 581.400 627.600 583.200 633.600 ;
        RECT 593.400 627.600 595.200 633.600 ;
        RECT 613.500 627.600 615.300 639.600 ;
        RECT 629.400 633.600 630.600 642.900 ;
        RECT 640.950 640.950 643.050 643.050 ;
        RECT 644.400 633.600 645.600 645.900 ;
        RECT 661.950 645.450 664.050 646.050 ;
        RECT 670.950 645.450 673.050 646.050 ;
        RECT 647.100 644.100 648.900 644.850 ;
        RECT 661.950 644.550 673.050 645.450 ;
        RECT 661.950 643.950 664.050 644.550 ;
        RECT 670.950 643.950 673.050 644.550 ;
        RECT 676.950 643.950 679.050 646.050 ;
        RECT 646.950 640.950 649.050 643.050 ;
        RECT 680.100 642.900 681.150 647.100 ;
        RECT 682.950 643.950 685.050 646.050 ;
        RECT 694.950 643.950 697.050 646.050 ;
        RECT 698.100 642.900 699.150 647.100 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 700.950 643.950 703.050 646.050 ;
        RECT 709.950 645.450 714.000 646.050 ;
        RECT 715.950 645.450 718.050 646.050 ;
        RECT 724.950 645.450 727.050 645.900 ;
        RECT 709.950 644.550 727.050 645.450 ;
        RECT 709.950 643.950 714.000 644.550 ;
        RECT 715.950 643.950 718.050 644.550 ;
        RECT 724.950 643.800 727.050 644.550 ;
        RECT 730.950 643.950 733.050 646.050 ;
        RECT 737.400 644.100 738.300 652.350 ;
        RECT 752.700 652.350 756.900 654.000 ;
        RECT 752.700 644.100 753.600 652.350 ;
        RECT 755.100 650.100 756.900 650.850 ;
        RECT 773.400 650.100 774.600 654.300 ;
        RECT 775.950 654.450 778.050 655.050 ;
        RECT 787.950 654.450 790.050 655.050 ;
        RECT 775.950 653.550 790.050 654.450 ;
        RECT 801.000 654.300 804.600 655.200 ;
        RECT 775.950 652.950 778.050 653.550 ;
        RECT 787.950 652.950 790.050 653.550 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 772.950 648.450 775.050 649.050 ;
        RECT 778.950 648.450 781.050 652.050 ;
        RECT 787.950 650.100 789.300 651.900 ;
        RECT 772.950 648.000 781.050 648.450 ;
        RECT 772.950 647.550 780.450 648.000 ;
        RECT 772.950 646.950 775.050 647.550 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 757.950 643.950 760.050 646.050 ;
        RECT 788.100 645.900 789.300 650.100 ;
        RECT 796.950 648.450 799.050 652.050 ;
        RECT 803.400 650.100 804.600 654.300 ;
        RECT 821.100 654.000 822.900 662.400 ;
        RECT 821.100 652.350 825.300 654.000 ;
        RECT 821.100 650.100 822.900 650.850 ;
        RECT 802.950 648.450 805.050 649.050 ;
        RECT 796.950 648.000 805.050 648.450 ;
        RECT 797.550 647.550 805.050 648.000 ;
        RECT 802.950 646.950 805.050 647.550 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 770.100 644.100 771.900 644.850 ;
        RECT 662.400 633.600 663.600 642.900 ;
        RECT 679.950 639.600 681.150 642.900 ;
        RECT 697.950 639.600 699.150 642.900 ;
        RECT 629.400 627.600 631.200 633.600 ;
        RECT 644.400 627.600 646.200 633.600 ;
        RECT 661.800 627.600 663.600 633.600 ;
        RECT 679.500 627.600 681.300 639.600 ;
        RECT 697.500 627.600 699.300 639.600 ;
        RECT 716.400 633.600 717.600 642.900 ;
        RECT 731.100 642.150 732.900 642.900 ;
        RECT 736.950 642.450 739.050 643.050 ;
        RECT 745.800 642.450 747.900 643.050 ;
        RECT 728.100 641.100 729.900 641.850 ;
        RECT 736.950 641.550 747.900 642.450 ;
        RECT 736.950 640.950 739.050 641.550 ;
        RECT 745.800 640.950 747.900 641.550 ;
        RECT 748.950 640.950 754.050 643.050 ;
        RECT 758.100 642.150 759.900 642.900 ;
        RECT 761.100 641.100 762.900 641.850 ;
        RECT 769.950 640.950 772.050 643.050 ;
        RECT 727.950 637.950 730.050 640.050 ;
        RECT 737.400 634.800 738.300 639.900 ;
        RECT 731.700 633.900 738.300 634.800 ;
        RECT 731.700 633.600 733.200 633.900 ;
        RECT 715.800 627.600 717.600 633.600 ;
        RECT 731.400 627.600 733.200 633.600 ;
        RECT 737.400 633.600 738.300 633.900 ;
        RECT 752.700 634.800 753.600 639.900 ;
        RECT 760.950 637.950 766.050 640.050 ;
        RECT 752.700 633.900 759.300 634.800 ;
        RECT 752.700 633.600 753.600 633.900 ;
        RECT 737.400 627.600 739.200 633.600 ;
        RECT 751.800 627.600 753.600 633.600 ;
        RECT 757.800 633.600 759.300 633.900 ;
        RECT 773.400 633.600 774.600 645.900 ;
        RECT 785.100 645.150 786.900 645.900 ;
        RECT 776.100 644.100 777.900 644.850 ;
        RECT 775.950 640.950 778.050 643.050 ;
        RECT 787.950 640.650 789.300 645.900 ;
        RECT 790.950 643.950 793.050 646.050 ;
        RECT 800.100 644.100 801.900 644.850 ;
        RECT 791.100 642.150 792.900 642.900 ;
        RECT 799.950 640.950 802.050 643.050 ;
        RECT 757.800 627.600 759.600 633.600 ;
        RECT 772.800 627.600 774.600 633.600 ;
        RECT 786.600 639.600 789.300 640.650 ;
        RECT 786.600 627.600 788.400 639.600 ;
        RECT 803.400 633.600 804.600 645.900 ;
        RECT 806.100 644.100 807.900 644.850 ;
        RECT 814.950 643.950 820.050 646.050 ;
        RECT 824.400 644.100 825.300 652.350 ;
        RECT 805.950 640.950 808.050 643.050 ;
        RECT 818.100 642.150 819.900 642.900 ;
        RECT 815.100 641.100 816.900 641.850 ;
        RECT 823.950 640.950 826.050 643.050 ;
        RECT 814.950 637.950 817.050 640.050 ;
        RECT 824.400 634.800 825.300 639.900 ;
        RECT 818.700 633.900 825.300 634.800 ;
        RECT 818.700 633.600 820.200 633.900 ;
        RECT 802.800 627.600 804.600 633.600 ;
        RECT 818.400 627.600 820.200 633.600 ;
        RECT 824.400 633.600 825.300 633.900 ;
        RECT 824.400 627.600 826.200 633.600 ;
        RECT 10.800 617.400 12.600 623.400 ;
        RECT 25.800 617.400 27.600 623.400 ;
        RECT 7.950 607.950 10.050 610.050 ;
        RECT 8.100 606.150 9.900 606.900 ;
        RECT 11.400 605.100 12.600 617.400 ;
        RECT 26.700 617.100 27.600 617.400 ;
        RECT 31.800 617.400 33.600 623.400 ;
        RECT 46.800 617.400 48.600 623.400 ;
        RECT 61.800 617.400 63.600 623.400 ;
        RECT 31.800 617.100 33.300 617.400 ;
        RECT 26.700 616.200 33.300 617.100 ;
        RECT 26.700 611.100 27.600 616.200 ;
        RECT 34.950 610.950 37.050 613.050 ;
        RECT 13.950 607.950 16.050 610.050 ;
        RECT 25.950 607.950 28.050 610.050 ;
        RECT 35.100 609.150 36.900 609.900 ;
        RECT 32.100 608.100 33.900 608.850 ;
        RECT 47.400 608.100 48.600 617.400 ;
        RECT 62.700 617.100 63.600 617.400 ;
        RECT 67.800 617.400 69.600 623.400 ;
        RECT 67.800 617.100 69.300 617.400 ;
        RECT 62.700 616.200 69.300 617.100 ;
        RECT 62.700 611.100 63.600 616.200 ;
        RECT 70.950 610.950 73.050 613.050 ;
        RECT 86.700 611.400 88.500 623.400 ;
        RECT 104.400 617.400 106.200 623.400 ;
        RECT 104.700 617.100 106.200 617.400 ;
        RECT 110.400 617.400 112.200 623.400 ;
        RECT 125.400 617.400 127.200 623.400 ;
        RECT 110.400 617.100 111.300 617.400 ;
        RECT 104.700 616.200 111.300 617.100 ;
        RECT 52.950 609.450 55.050 610.050 ;
        RECT 61.950 609.450 64.050 610.050 ;
        RECT 52.950 608.550 64.050 609.450 ;
        RECT 71.100 609.150 72.900 609.900 ;
        RECT 52.950 607.950 55.050 608.550 ;
        RECT 61.950 607.950 64.050 608.550 ;
        RECT 68.100 608.100 69.900 608.850 ;
        RECT 86.850 608.100 88.050 611.400 ;
        RECT 100.950 610.950 103.050 613.050 ;
        RECT 110.400 611.100 111.300 616.200 ;
        RECT 101.100 609.150 102.900 609.900 ;
        RECT 104.100 608.100 105.900 608.850 ;
        RECT 14.100 606.150 15.900 606.900 ;
        RECT 10.950 603.450 13.050 604.050 ;
        RECT 15.000 603.450 19.050 604.050 ;
        RECT 10.950 602.550 19.050 603.450 ;
        RECT 10.950 601.950 13.050 602.550 ;
        RECT 15.000 601.950 19.050 602.550 ;
        RECT 11.400 596.700 12.600 600.900 ;
        RECT 26.700 598.650 27.600 606.900 ;
        RECT 31.950 604.950 34.050 607.050 ;
        RECT 46.950 604.950 49.050 607.050 ;
        RECT 28.950 601.950 31.050 604.050 ;
        RECT 29.100 600.150 30.900 600.900 ;
        RECT 26.700 597.000 30.900 598.650 ;
        RECT 9.000 595.800 12.600 596.700 ;
        RECT 9.000 588.600 10.800 595.800 ;
        RECT 16.950 594.450 19.050 595.050 ;
        RECT 25.950 594.450 28.050 595.050 ;
        RECT 16.950 593.550 28.050 594.450 ;
        RECT 16.950 592.950 19.050 593.550 ;
        RECT 25.950 592.950 28.050 593.550 ;
        RECT 29.100 588.600 30.900 597.000 ;
        RECT 47.400 591.600 48.600 603.900 ;
        RECT 50.100 602.100 51.900 602.850 ;
        RECT 49.950 598.950 52.050 601.050 ;
        RECT 62.700 598.650 63.600 606.900 ;
        RECT 67.950 604.950 70.050 607.050 ;
        RECT 82.950 604.950 85.050 607.050 ;
        RECT 64.950 601.950 67.050 604.050 ;
        RECT 86.850 603.900 87.900 608.100 ;
        RECT 109.950 607.950 112.050 610.050 ;
        RECT 121.950 607.950 124.050 610.050 ;
        RECT 88.950 604.950 91.050 607.050 ;
        RECT 103.950 604.950 106.050 607.050 ;
        RECT 83.100 603.150 84.900 603.900 ;
        RECT 86.850 602.100 88.050 603.900 ;
        RECT 89.100 603.150 90.900 603.900 ;
        RECT 92.100 602.100 93.900 602.850 ;
        RECT 106.950 601.950 109.050 604.050 ;
        RECT 65.100 600.150 66.900 600.900 ;
        RECT 70.950 600.450 73.050 601.050 ;
        RECT 85.950 600.450 88.050 601.050 ;
        RECT 70.950 599.550 88.050 600.450 ;
        RECT 70.950 598.950 73.050 599.550 ;
        RECT 85.950 598.950 88.050 599.550 ;
        RECT 91.950 598.950 94.050 601.050 ;
        RECT 107.100 600.150 108.900 600.900 ;
        RECT 110.400 598.650 111.300 606.900 ;
        RECT 122.100 606.150 123.900 606.900 ;
        RECT 125.400 605.100 126.600 617.400 ;
        RECT 142.500 611.400 144.300 623.400 ;
        RECT 155.400 612.600 157.200 623.400 ;
        RECT 161.400 622.500 169.200 623.400 ;
        RECT 161.400 612.600 163.200 622.500 ;
        RECT 155.400 611.700 163.200 612.600 ;
        RECT 127.950 607.950 130.050 610.050 ;
        RECT 142.950 608.100 144.150 611.400 ;
        RECT 164.400 610.500 166.200 621.600 ;
        RECT 167.400 611.400 169.200 622.500 ;
        RECT 179.400 612.600 181.200 623.400 ;
        RECT 185.400 622.500 193.200 623.400 ;
        RECT 185.400 612.600 187.200 622.500 ;
        RECT 179.400 611.700 187.200 612.600 ;
        RECT 188.400 610.500 190.200 621.600 ;
        RECT 191.400 611.400 193.200 622.500 ;
        RECT 203.400 611.400 205.200 623.400 ;
        RECT 218.400 617.400 220.200 623.400 ;
        RECT 218.700 617.100 220.200 617.400 ;
        RECT 224.400 617.400 226.200 623.400 ;
        RECT 238.800 617.400 240.600 623.400 ;
        RECT 251.400 617.400 253.200 623.400 ;
        RECT 224.400 617.100 225.300 617.400 ;
        RECT 218.700 616.200 225.300 617.100 ;
        RECT 128.100 606.150 129.900 606.900 ;
        RECT 139.950 604.950 142.050 607.050 ;
        RECT 115.950 603.450 118.050 604.050 ;
        RECT 124.950 603.450 127.050 604.050 ;
        RECT 143.100 603.900 144.150 608.100 ;
        RECT 162.150 609.600 166.200 610.500 ;
        RECT 186.150 609.600 190.200 610.500 ;
        RECT 162.150 608.100 163.050 609.600 ;
        RECT 186.150 608.100 187.050 609.600 ;
        RECT 145.950 604.950 148.050 607.050 ;
        RECT 157.950 604.950 160.050 607.050 ;
        RECT 162.150 603.900 162.900 608.100 ;
        RECT 163.950 604.950 166.050 607.050 ;
        RECT 181.950 604.950 184.050 607.050 ;
        RECT 186.150 603.900 186.900 608.100 ;
        RECT 187.950 604.950 190.050 607.050 ;
        RECT 199.950 604.950 202.050 607.050 ;
        RECT 115.950 602.550 127.050 603.450 ;
        RECT 140.100 603.150 141.900 603.900 ;
        RECT 115.950 601.950 118.050 602.550 ;
        RECT 124.950 601.950 127.050 602.550 ;
        RECT 137.100 602.100 138.900 602.850 ;
        RECT 142.950 602.100 144.150 603.900 ;
        RECT 146.100 603.150 147.900 603.900 ;
        RECT 158.250 603.150 160.050 603.900 ;
        RECT 155.250 602.100 157.050 602.850 ;
        RECT 162.150 602.100 163.050 603.900 ;
        RECT 163.950 603.150 165.750 603.900 ;
        RECT 182.250 603.150 184.050 603.900 ;
        RECT 167.100 602.100 168.900 602.850 ;
        RECT 179.250 602.100 181.050 602.850 ;
        RECT 186.150 602.100 187.050 603.900 ;
        RECT 187.950 603.150 189.750 603.900 ;
        RECT 200.100 603.150 201.900 603.900 ;
        RECT 191.100 602.100 192.900 602.850 ;
        RECT 203.400 602.100 204.600 611.400 ;
        RECT 214.950 610.950 217.050 613.050 ;
        RECT 224.400 611.100 225.300 616.200 ;
        RECT 215.100 609.150 216.900 609.900 ;
        RECT 218.100 608.100 219.900 608.850 ;
        RECT 223.950 607.950 226.050 610.050 ;
        RECT 217.950 604.950 220.050 607.050 ;
        RECT 220.950 601.800 223.050 604.050 ;
        RECT 62.700 597.000 66.900 598.650 ;
        RECT 85.950 597.750 87.150 597.900 ;
        RECT 46.800 588.600 48.600 591.600 ;
        RECT 65.100 588.600 66.900 597.000 ;
        RECT 83.400 596.700 87.150 597.750 ;
        RECT 107.100 597.000 111.300 598.650 ;
        RECT 83.400 594.600 84.600 596.700 ;
        RECT 82.800 588.600 84.600 594.600 ;
        RECT 85.800 593.700 93.600 595.050 ;
        RECT 85.800 588.600 87.600 593.700 ;
        RECT 91.800 588.600 93.600 593.700 ;
        RECT 107.100 588.600 108.900 597.000 ;
        RECT 125.400 596.700 126.600 600.900 ;
        RECT 136.950 598.800 139.050 601.050 ;
        RECT 142.950 598.950 145.050 601.050 ;
        RECT 154.950 598.950 157.050 601.050 ;
        RECT 160.950 598.950 163.050 601.050 ;
        RECT 166.950 598.950 169.050 601.050 ;
        RECT 178.950 598.950 181.050 601.050 ;
        RECT 184.950 598.800 187.050 601.050 ;
        RECT 190.950 598.950 193.050 601.050 ;
        RECT 202.950 598.950 205.050 601.050 ;
        RECT 221.100 600.150 222.900 600.900 ;
        RECT 224.400 598.650 225.300 606.900 ;
        RECT 232.950 606.450 235.050 610.050 ;
        RECT 239.400 608.100 240.600 617.400 ;
        RECT 251.700 617.100 253.200 617.400 ;
        RECT 257.400 617.400 259.200 623.400 ;
        RECT 272.400 617.400 274.200 623.400 ;
        RECT 257.400 617.100 258.300 617.400 ;
        RECT 251.700 616.200 258.300 617.100 ;
        RECT 247.950 610.950 250.050 613.050 ;
        RECT 257.400 611.100 258.300 616.200 ;
        RECT 248.100 609.150 249.900 609.900 ;
        RECT 251.100 608.100 252.900 608.850 ;
        RECT 256.950 607.950 259.050 610.050 ;
        RECT 268.950 607.950 271.050 610.200 ;
        RECT 238.950 606.450 241.050 607.050 ;
        RECT 232.950 606.000 241.050 606.450 ;
        RECT 233.550 605.550 241.050 606.000 ;
        RECT 238.950 604.950 241.050 605.550 ;
        RECT 250.950 604.950 253.050 607.050 ;
        RECT 143.850 597.750 145.050 597.900 ;
        RECT 143.850 596.700 147.600 597.750 ;
        RECT 125.400 595.800 129.000 596.700 ;
        RECT 127.200 588.600 129.000 595.800 ;
        RECT 137.400 593.700 145.200 595.050 ;
        RECT 137.400 588.600 139.200 593.700 ;
        RECT 143.400 588.600 145.200 593.700 ;
        RECT 146.400 594.600 147.600 596.700 ;
        RECT 160.950 594.600 162.000 597.900 ;
        RECT 184.950 594.600 186.000 597.900 ;
        RECT 146.400 588.600 148.200 594.600 ;
        RECT 160.200 588.600 162.000 594.600 ;
        RECT 184.200 588.600 186.000 594.600 ;
        RECT 203.400 594.600 204.600 597.900 ;
        RECT 221.100 597.000 225.300 598.650 ;
        RECT 203.400 588.600 205.200 594.600 ;
        RECT 221.100 588.600 222.900 597.000 ;
        RECT 239.400 591.600 240.600 603.900 ;
        RECT 242.100 602.100 243.900 602.850 ;
        RECT 253.950 601.950 256.050 604.050 ;
        RECT 241.950 600.450 244.050 601.050 ;
        RECT 246.000 600.450 250.050 601.050 ;
        RECT 241.950 599.550 250.050 600.450 ;
        RECT 254.100 600.150 255.900 600.900 ;
        RECT 241.950 598.950 244.050 599.550 ;
        RECT 246.000 598.950 250.050 599.550 ;
        RECT 257.400 598.650 258.300 606.900 ;
        RECT 269.100 606.150 270.900 606.900 ;
        RECT 272.400 605.100 273.600 617.400 ;
        RECT 293.700 611.400 295.500 623.400 ;
        RECT 310.200 611.400 312.000 623.400 ;
        RECT 316.800 617.400 318.600 623.400 ;
        RECT 293.850 608.100 295.050 611.400 ;
        RECT 275.100 606.150 276.900 606.900 ;
        RECT 289.950 604.800 292.050 607.050 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 293.850 603.900 294.900 608.100 ;
        RECT 295.950 604.950 298.050 607.050 ;
        RECT 290.100 603.150 291.900 603.900 ;
        RECT 293.850 602.100 295.050 603.900 ;
        RECT 296.100 603.150 297.900 603.900 ;
        RECT 299.100 602.100 300.900 602.850 ;
        RECT 310.950 602.100 312.000 611.400 ;
        RECT 314.100 603.150 315.900 603.900 ;
        RECT 238.800 588.600 240.600 591.600 ;
        RECT 254.100 597.000 258.300 598.650 ;
        RECT 254.100 588.600 255.900 597.000 ;
        RECT 272.400 596.700 273.600 600.900 ;
        RECT 277.950 600.450 280.050 601.050 ;
        RECT 292.950 600.450 295.050 601.050 ;
        RECT 277.950 599.550 295.050 600.450 ;
        RECT 277.950 598.950 280.050 599.550 ;
        RECT 292.950 598.950 295.050 599.550 ;
        RECT 298.950 598.950 301.050 601.050 ;
        RECT 304.950 600.450 309.000 601.050 ;
        RECT 310.950 600.450 313.050 601.050 ;
        RECT 304.950 599.550 313.050 600.450 ;
        RECT 304.950 598.950 309.000 599.550 ;
        RECT 310.950 598.950 313.050 599.550 ;
        RECT 292.950 597.750 294.150 597.900 ;
        RECT 290.400 596.700 294.150 597.750 ;
        RECT 272.400 595.800 276.000 596.700 ;
        RECT 274.200 588.600 276.000 595.800 ;
        RECT 290.400 594.600 291.600 596.700 ;
        RECT 289.800 588.600 291.600 594.600 ;
        RECT 292.800 593.700 300.600 595.050 ;
        RECT 292.800 588.600 294.600 593.700 ;
        RECT 298.800 588.600 300.600 593.700 ;
        RECT 312.150 594.600 313.050 597.900 ;
        RECT 317.550 597.300 318.600 617.400 ;
        RECT 329.400 617.400 331.200 623.400 ;
        RECT 343.800 617.400 345.600 623.400 ;
        RECT 325.950 607.950 328.050 610.050 ;
        RECT 326.100 606.150 327.900 606.900 ;
        RECT 320.100 605.100 321.900 605.850 ;
        RECT 329.400 605.100 330.600 617.400 ;
        RECT 344.700 617.100 345.600 617.400 ;
        RECT 349.800 617.400 351.600 623.400 ;
        RECT 365.400 617.400 367.200 623.400 ;
        RECT 349.800 617.100 351.300 617.400 ;
        RECT 344.700 616.200 351.300 617.100 ;
        RECT 344.700 611.100 345.600 616.200 ;
        RECT 352.950 610.950 355.050 613.050 ;
        RECT 331.950 607.950 334.050 610.050 ;
        RECT 337.950 609.450 342.000 610.050 ;
        RECT 343.950 609.450 346.050 610.050 ;
        RECT 337.950 608.550 346.050 609.450 ;
        RECT 353.100 609.150 354.900 609.900 ;
        RECT 337.950 607.950 342.000 608.550 ;
        RECT 343.950 607.950 346.050 608.550 ;
        RECT 350.100 608.100 351.900 608.850 ;
        RECT 361.950 607.950 364.050 610.050 ;
        RECT 332.100 606.150 333.900 606.900 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 328.950 603.450 331.050 604.050 ;
        RECT 333.000 603.450 337.050 604.050 ;
        RECT 328.950 602.550 337.050 603.450 ;
        RECT 328.950 601.950 331.050 602.550 ;
        RECT 333.000 601.950 337.050 602.550 ;
        RECT 314.100 596.400 321.600 597.300 ;
        RECT 314.100 595.500 315.900 596.400 ;
        RECT 312.150 592.800 314.100 594.600 ;
        RECT 312.300 588.600 314.100 592.800 ;
        RECT 319.800 588.600 321.600 596.400 ;
        RECT 329.400 596.700 330.600 600.900 ;
        RECT 344.700 598.650 345.600 606.900 ;
        RECT 349.950 604.950 352.050 607.050 ;
        RECT 362.100 606.150 363.900 606.900 ;
        RECT 365.400 605.100 366.600 617.400 ;
        RECT 382.500 611.400 384.300 623.400 ;
        RECT 400.200 611.400 402.000 623.400 ;
        RECT 406.800 617.400 408.600 623.400 ;
        RECT 382.950 608.100 384.150 611.400 ;
        RECT 368.100 606.150 369.900 606.900 ;
        RECT 379.950 604.950 382.050 607.050 ;
        RECT 346.950 601.950 349.050 604.050 ;
        RECT 358.950 603.450 363.000 604.050 ;
        RECT 364.950 603.450 367.050 604.050 ;
        RECT 383.100 603.900 384.150 608.100 ;
        RECT 385.950 604.950 388.050 607.050 ;
        RECT 358.950 602.550 367.050 603.450 ;
        RECT 380.100 603.150 381.900 603.900 ;
        RECT 358.950 601.950 363.000 602.550 ;
        RECT 364.950 601.950 367.050 602.550 ;
        RECT 377.100 602.100 378.900 602.850 ;
        RECT 382.950 602.100 384.150 603.900 ;
        RECT 386.100 603.150 387.900 603.900 ;
        RECT 400.950 602.100 402.000 611.400 ;
        RECT 404.100 603.150 405.900 603.900 ;
        RECT 347.100 600.150 348.900 600.900 ;
        RECT 344.700 597.000 348.900 598.650 ;
        RECT 329.400 595.800 333.000 596.700 ;
        RECT 331.200 588.600 333.000 595.800 ;
        RECT 347.100 588.600 348.900 597.000 ;
        RECT 365.400 596.700 366.600 600.900 ;
        RECT 376.950 598.950 379.050 601.050 ;
        RECT 382.950 598.950 385.050 601.050 ;
        RECT 391.950 600.450 394.050 601.050 ;
        RECT 400.950 600.450 403.050 601.050 ;
        RECT 391.950 599.550 403.050 600.450 ;
        RECT 391.950 598.950 394.050 599.550 ;
        RECT 400.950 598.950 403.050 599.550 ;
        RECT 383.850 597.750 385.050 597.900 ;
        RECT 383.850 596.700 387.600 597.750 ;
        RECT 365.400 595.800 369.000 596.700 ;
        RECT 367.200 588.600 369.000 595.800 ;
        RECT 377.400 593.700 385.200 595.050 ;
        RECT 377.400 588.600 379.200 593.700 ;
        RECT 383.400 588.600 385.200 593.700 ;
        RECT 386.400 594.600 387.600 596.700 ;
        RECT 402.150 594.600 403.050 597.900 ;
        RECT 407.550 597.300 408.600 617.400 ;
        RECT 421.500 611.400 423.300 623.400 ;
        RECT 437.400 617.400 439.200 623.400 ;
        RECT 421.950 608.100 423.150 611.400 ;
        RECT 410.100 605.100 411.900 605.850 ;
        RECT 418.950 604.950 421.050 607.050 ;
        RECT 409.950 598.950 412.050 604.050 ;
        RECT 422.100 603.900 423.150 608.100 ;
        RECT 430.950 607.950 436.050 610.050 ;
        RECT 424.950 604.950 427.050 607.050 ;
        RECT 434.100 606.150 435.900 606.900 ;
        RECT 437.400 605.100 438.600 617.400 ;
        RECT 454.500 611.400 456.300 623.400 ;
        RECT 472.200 611.400 474.000 623.400 ;
        RECT 478.800 617.400 480.600 623.400 ;
        RECT 496.800 617.400 498.600 623.400 ;
        RECT 439.950 607.950 442.050 610.050 ;
        RECT 454.950 608.100 456.150 611.400 ;
        RECT 440.100 606.150 441.900 606.900 ;
        RECT 451.950 604.950 454.050 607.050 ;
        RECT 419.100 603.150 420.900 603.900 ;
        RECT 416.100 602.100 417.900 602.850 ;
        RECT 421.950 602.100 423.150 603.900 ;
        RECT 425.100 603.150 426.900 603.900 ;
        RECT 433.950 601.950 439.050 604.050 ;
        RECT 455.100 603.900 456.150 608.100 ;
        RECT 457.950 604.950 460.050 607.050 ;
        RECT 452.100 603.150 453.900 603.900 ;
        RECT 449.100 602.100 450.900 602.850 ;
        RECT 454.950 602.100 456.150 603.900 ;
        RECT 458.100 603.150 459.900 603.900 ;
        RECT 472.950 602.100 474.000 611.400 ;
        RECT 476.100 603.150 477.900 603.900 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 421.950 598.800 424.050 601.050 ;
        RECT 422.850 597.750 424.050 597.900 ;
        RECT 404.100 596.400 411.600 597.300 ;
        RECT 422.850 596.700 426.600 597.750 ;
        RECT 404.100 595.500 405.900 596.400 ;
        RECT 386.400 588.600 388.200 594.600 ;
        RECT 402.150 592.800 404.100 594.600 ;
        RECT 402.300 588.600 404.100 592.800 ;
        RECT 409.800 588.600 411.600 596.400 ;
        RECT 416.400 593.700 424.200 595.050 ;
        RECT 416.400 588.600 418.200 593.700 ;
        RECT 422.400 588.600 424.200 593.700 ;
        RECT 425.400 594.600 426.600 596.700 ;
        RECT 437.400 596.700 438.600 600.900 ;
        RECT 448.950 598.950 451.050 601.050 ;
        RECT 454.950 598.950 457.050 601.050 ;
        RECT 460.950 600.450 463.050 601.200 ;
        RECT 472.950 600.450 475.050 601.050 ;
        RECT 460.950 599.550 475.050 600.450 ;
        RECT 460.950 599.100 463.050 599.550 ;
        RECT 472.950 598.950 475.050 599.550 ;
        RECT 455.850 597.750 457.050 597.900 ;
        RECT 455.850 596.700 459.600 597.750 ;
        RECT 437.400 595.800 441.000 596.700 ;
        RECT 425.400 588.600 427.200 594.600 ;
        RECT 439.200 588.600 441.000 595.800 ;
        RECT 449.400 593.700 457.200 595.050 ;
        RECT 449.400 588.600 451.200 593.700 ;
        RECT 455.400 588.600 457.200 593.700 ;
        RECT 458.400 594.600 459.600 596.700 ;
        RECT 474.150 594.600 475.050 597.900 ;
        RECT 479.550 597.300 480.600 617.400 ;
        RECT 494.100 606.150 495.900 606.900 ;
        RECT 482.100 605.100 483.900 605.850 ;
        RECT 497.400 605.100 498.600 617.400 ;
        RECT 513.600 611.400 515.400 623.400 ;
        RECT 529.500 611.400 531.300 623.400 ;
        RECT 550.800 617.400 552.600 623.400 ;
        RECT 566.400 617.400 568.200 623.400 ;
        RECT 512.700 610.350 515.400 611.400 ;
        RECT 499.950 607.950 502.050 610.050 ;
        RECT 509.100 608.100 510.900 608.850 ;
        RECT 500.100 606.150 501.900 606.900 ;
        RECT 508.950 604.950 511.050 607.050 ;
        RECT 512.700 605.100 514.050 610.350 ;
        RECT 529.950 608.100 531.150 611.400 ;
        RECT 515.100 605.100 516.900 605.850 ;
        RECT 481.950 601.950 484.050 604.050 ;
        RECT 487.950 603.450 490.050 604.050 ;
        RECT 496.950 603.450 499.050 604.050 ;
        RECT 501.000 603.450 505.050 604.050 ;
        RECT 487.950 602.550 505.050 603.450 ;
        RECT 487.950 601.950 490.050 602.550 ;
        RECT 496.950 601.950 499.050 602.550 ;
        RECT 501.000 601.950 505.050 602.550 ;
        RECT 512.700 600.900 513.900 605.100 ;
        RECT 523.950 604.950 529.050 607.050 ;
        RECT 514.950 601.800 517.050 604.050 ;
        RECT 530.100 603.900 531.150 608.100 ;
        RECT 532.950 604.950 535.050 607.050 ;
        RECT 548.100 606.150 549.900 606.900 ;
        RECT 551.400 605.100 552.600 617.400 ;
        RECT 566.700 617.100 568.200 617.400 ;
        RECT 572.400 617.400 574.200 623.400 ;
        RECT 572.400 617.100 573.300 617.400 ;
        RECT 566.700 616.200 573.300 617.100 ;
        RECT 562.950 610.950 565.050 613.050 ;
        RECT 572.400 611.100 573.300 616.200 ;
        RECT 583.800 611.400 585.600 623.400 ;
        RECT 598.800 617.400 600.600 623.400 ;
        RECT 616.800 617.400 618.600 623.400 ;
        RECT 632.400 617.400 634.200 623.400 ;
        RECT 553.950 607.950 556.050 610.050 ;
        RECT 563.100 609.150 564.900 609.900 ;
        RECT 571.950 609.450 574.050 610.050 ;
        RECT 576.000 609.450 580.050 610.050 ;
        RECT 566.100 608.100 567.900 608.850 ;
        RECT 571.950 608.550 580.050 609.450 ;
        RECT 571.950 607.950 574.050 608.550 ;
        RECT 576.000 607.950 580.050 608.550 ;
        RECT 554.100 606.150 555.900 606.900 ;
        RECT 527.100 603.150 528.900 603.900 ;
        RECT 524.100 602.100 525.900 602.850 ;
        RECT 529.950 602.100 531.150 603.900 ;
        RECT 533.100 603.150 534.900 603.900 ;
        RECT 538.950 603.450 541.050 603.900 ;
        RECT 544.950 603.450 547.050 604.050 ;
        RECT 538.950 602.550 547.050 603.450 ;
        RECT 538.950 601.800 541.050 602.550 ;
        RECT 544.950 601.950 547.050 602.550 ;
        RECT 550.950 603.450 553.050 604.050 ;
        RECT 559.950 603.450 562.050 604.050 ;
        RECT 550.950 602.550 562.050 603.450 ;
        RECT 550.950 601.950 553.050 602.550 ;
        RECT 559.950 601.950 562.050 602.550 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 476.100 596.400 483.600 597.300 ;
        RECT 497.400 596.700 498.600 600.900 ;
        RECT 512.700 599.100 514.050 600.900 ;
        RECT 523.950 598.950 526.050 601.050 ;
        RECT 529.950 598.950 532.050 601.050 ;
        RECT 476.100 595.500 477.900 596.400 ;
        RECT 458.400 588.600 460.200 594.600 ;
        RECT 474.150 592.800 476.100 594.600 ;
        RECT 474.300 588.600 476.100 592.800 ;
        RECT 481.800 588.600 483.600 596.400 ;
        RECT 495.000 595.800 498.600 596.700 ;
        RECT 508.950 595.950 514.050 598.050 ;
        RECT 530.850 597.750 532.050 597.900 ;
        RECT 530.850 596.700 534.600 597.750 ;
        RECT 551.400 596.700 552.600 600.900 ;
        RECT 569.100 600.150 570.900 600.900 ;
        RECT 572.400 598.650 573.300 606.900 ;
        RECT 584.400 602.100 585.600 611.400 ;
        RECT 596.100 606.150 597.900 606.900 ;
        RECT 599.400 605.100 600.600 617.400 ;
        RECT 601.950 607.950 604.050 610.050 ;
        RECT 613.950 607.950 616.050 610.050 ;
        RECT 602.100 606.150 603.900 606.900 ;
        RECT 614.100 606.150 615.900 606.900 ;
        RECT 617.400 605.100 618.600 617.400 ;
        RECT 632.700 617.100 634.200 617.400 ;
        RECT 638.400 617.400 640.200 623.400 ;
        RECT 638.400 617.100 639.300 617.400 ;
        RECT 632.700 616.200 639.300 617.100 ;
        RECT 628.950 610.950 631.050 613.050 ;
        RECT 638.400 611.100 639.300 616.200 ;
        RECT 647.400 612.300 649.200 623.400 ;
        RECT 653.400 612.300 655.200 623.400 ;
        RECT 647.400 611.400 655.200 612.300 ;
        RECT 656.400 611.400 658.200 623.400 ;
        RECT 668.400 612.300 670.200 623.400 ;
        RECT 674.400 612.300 676.200 623.400 ;
        RECT 668.400 611.400 676.200 612.300 ;
        RECT 677.400 611.400 679.200 623.400 ;
        RECT 692.400 617.400 694.200 623.400 ;
        RECT 692.700 617.100 694.200 617.400 ;
        RECT 698.400 617.400 700.200 623.400 ;
        RECT 698.400 617.100 699.300 617.400 ;
        RECT 692.700 616.200 699.300 617.100 ;
        RECT 619.950 607.950 622.050 610.050 ;
        RECT 629.100 609.150 630.900 609.900 ;
        RECT 632.100 608.100 633.900 608.850 ;
        RECT 637.950 607.950 643.050 610.050 ;
        RECT 620.100 606.150 621.900 606.900 ;
        RECT 631.950 604.950 634.050 607.050 ;
        RECT 587.100 603.150 588.900 603.900 ;
        RECT 598.950 601.950 604.050 604.050 ;
        RECT 607.950 603.450 610.050 604.050 ;
        RECT 616.950 603.450 619.050 604.050 ;
        RECT 607.950 602.550 619.050 603.450 ;
        RECT 607.950 601.950 610.050 602.550 ;
        RECT 616.950 601.950 619.050 602.550 ;
        RECT 634.950 601.950 637.050 604.050 ;
        RECT 574.950 600.450 577.050 601.050 ;
        RECT 583.950 600.450 586.050 601.050 ;
        RECT 574.950 599.550 586.050 600.450 ;
        RECT 574.950 598.950 577.050 599.550 ;
        RECT 583.950 598.950 586.050 599.550 ;
        RECT 495.000 588.600 496.800 595.800 ;
        RECT 512.400 591.600 513.600 594.900 ;
        RECT 524.400 593.700 532.200 595.050 ;
        RECT 512.400 588.600 514.200 591.600 ;
        RECT 524.400 588.600 526.200 593.700 ;
        RECT 530.400 588.600 532.200 593.700 ;
        RECT 533.400 594.600 534.600 596.700 ;
        RECT 549.000 595.800 552.600 596.700 ;
        RECT 569.100 597.000 573.300 598.650 ;
        RECT 533.400 588.600 535.200 594.600 ;
        RECT 549.000 588.600 550.800 595.800 ;
        RECT 569.100 588.600 570.900 597.000 ;
        RECT 584.400 594.600 585.600 597.900 ;
        RECT 599.400 596.700 600.600 600.900 ;
        RECT 617.400 596.700 618.600 600.900 ;
        RECT 635.100 600.150 636.900 600.900 ;
        RECT 638.400 598.650 639.300 606.900 ;
        RECT 646.950 604.950 649.050 607.050 ;
        RECT 652.950 604.950 655.050 607.050 ;
        RECT 647.100 603.150 648.900 603.900 ;
        RECT 653.100 603.150 654.900 603.900 ;
        RECT 650.100 602.100 651.900 602.850 ;
        RECT 656.700 602.100 657.600 611.400 ;
        RECT 667.950 604.950 670.050 607.050 ;
        RECT 673.950 604.950 676.050 607.050 ;
        RECT 668.100 603.150 669.900 603.900 ;
        RECT 674.100 603.150 675.900 603.900 ;
        RECT 671.100 602.100 672.900 602.850 ;
        RECT 677.700 602.100 678.600 611.400 ;
        RECT 688.950 610.950 691.050 613.050 ;
        RECT 698.400 611.100 699.300 616.200 ;
        RECT 712.800 611.400 714.600 623.400 ;
        RECT 715.800 612.300 717.600 623.400 ;
        RECT 721.800 612.300 723.600 623.400 ;
        RECT 730.800 617.400 732.600 623.400 ;
        RECT 715.800 611.400 723.600 612.300 ;
        RECT 689.100 609.150 690.900 609.900 ;
        RECT 697.950 609.450 700.050 610.050 ;
        RECT 706.950 609.450 709.050 610.050 ;
        RECT 692.100 608.100 693.900 608.850 ;
        RECT 697.950 608.550 709.050 609.450 ;
        RECT 697.950 607.950 700.050 608.550 ;
        RECT 706.950 607.950 709.050 608.550 ;
        RECT 691.950 604.950 694.050 607.050 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 649.950 598.950 652.050 601.050 ;
        RECT 655.950 598.950 661.050 601.050 ;
        RECT 670.950 598.950 673.050 601.050 ;
        RECT 676.950 600.450 679.050 601.050 ;
        RECT 688.950 600.450 691.050 601.050 ;
        RECT 676.950 599.550 691.050 600.450 ;
        RECT 695.100 600.150 696.900 600.900 ;
        RECT 676.950 598.950 679.050 599.550 ;
        RECT 688.950 598.950 691.050 599.550 ;
        RECT 698.400 598.650 699.300 606.900 ;
        RECT 713.400 602.100 714.300 611.400 ;
        RECT 731.400 608.100 732.600 617.400 ;
        RECT 749.700 611.400 751.500 623.400 ;
        RECT 763.800 617.400 765.600 623.400 ;
        RECT 749.850 608.100 751.050 611.400 ;
        RECT 764.400 608.100 765.600 617.400 ;
        RECT 776.400 617.400 778.200 623.400 ;
        RECT 791.400 617.400 793.200 623.400 ;
        RECT 776.400 608.100 777.600 617.400 ;
        RECT 791.700 617.100 793.200 617.400 ;
        RECT 797.400 617.400 799.200 623.400 ;
        RECT 808.800 617.400 810.600 623.400 ;
        RECT 797.400 617.100 798.300 617.400 ;
        RECT 791.700 616.200 798.300 617.100 ;
        RECT 787.950 610.950 790.050 613.050 ;
        RECT 797.400 611.100 798.300 616.200 ;
        RECT 809.700 617.100 810.600 617.400 ;
        RECT 814.800 617.400 816.600 623.400 ;
        RECT 814.800 617.100 816.300 617.400 ;
        RECT 809.700 616.200 816.300 617.100 ;
        RECT 809.700 611.100 810.600 616.200 ;
        RECT 817.950 610.950 820.050 613.050 ;
        RECT 788.100 609.150 789.900 609.900 ;
        RECT 791.100 608.100 792.900 608.850 ;
        RECT 715.950 604.950 718.050 607.050 ;
        RECT 721.950 604.950 724.050 607.050 ;
        RECT 730.950 606.450 733.050 607.050 ;
        RECT 745.950 606.450 748.050 607.050 ;
        RECT 730.950 605.550 748.050 606.450 ;
        RECT 730.950 604.950 733.050 605.550 ;
        RECT 745.950 604.950 748.050 605.550 ;
        RECT 749.850 603.900 750.900 608.100 ;
        RECT 796.950 607.950 799.050 610.050 ;
        RECT 802.950 609.450 807.000 610.050 ;
        RECT 808.950 609.450 811.050 610.050 ;
        RECT 802.950 608.550 811.050 609.450 ;
        RECT 818.100 609.150 819.900 609.900 ;
        RECT 802.950 607.950 807.000 608.550 ;
        RECT 808.950 607.950 811.050 608.550 ;
        RECT 815.100 608.100 816.900 608.850 ;
        RECT 751.950 604.950 754.050 607.050 ;
        RECT 760.950 604.950 766.050 607.050 ;
        RECT 775.950 606.450 778.050 607.050 ;
        RECT 784.950 606.450 787.050 607.050 ;
        RECT 775.950 605.550 787.050 606.450 ;
        RECT 775.950 604.950 778.050 605.550 ;
        RECT 784.950 604.950 787.050 605.550 ;
        RECT 790.950 604.950 793.050 607.200 ;
        RECT 716.100 603.150 717.900 603.900 ;
        RECT 722.100 603.150 723.900 603.900 ;
        RECT 719.100 602.100 720.900 602.850 ;
        RECT 709.950 598.950 715.050 601.050 ;
        RECT 718.950 598.950 721.050 601.050 ;
        RECT 583.800 588.600 585.600 594.600 ;
        RECT 597.000 595.800 600.600 596.700 ;
        RECT 615.000 595.800 618.600 596.700 ;
        RECT 635.100 597.000 639.300 598.650 ;
        RECT 597.000 588.600 598.800 595.800 ;
        RECT 615.000 588.600 616.800 595.800 ;
        RECT 635.100 588.600 636.900 597.000 ;
        RECT 656.700 594.600 657.600 597.900 ;
        RECT 677.700 594.600 678.600 597.900 ;
        RECT 652.200 592.950 657.600 594.600 ;
        RECT 673.200 592.950 678.600 594.600 ;
        RECT 695.100 597.000 699.300 598.650 ;
        RECT 652.200 588.600 654.000 592.950 ;
        RECT 673.200 588.600 675.000 592.950 ;
        RECT 695.100 588.600 696.900 597.000 ;
        RECT 713.400 594.600 714.300 597.900 ;
        RECT 713.400 592.950 718.800 594.600 ;
        RECT 717.000 588.600 718.800 592.950 ;
        RECT 731.400 591.600 732.600 603.900 ;
        RECT 746.100 603.150 747.900 603.900 ;
        RECT 734.100 602.100 735.900 602.850 ;
        RECT 749.850 602.100 751.050 603.900 ;
        RECT 752.100 603.150 753.900 603.900 ;
        RECT 755.100 602.100 756.900 602.850 ;
        RECT 733.950 598.950 736.050 601.050 ;
        RECT 748.950 598.950 751.050 601.050 ;
        RECT 754.950 598.950 757.050 601.050 ;
        RECT 748.950 597.750 750.150 597.900 ;
        RECT 746.400 596.700 750.150 597.750 ;
        RECT 746.400 594.600 747.600 596.700 ;
        RECT 730.800 588.600 732.600 591.600 ;
        RECT 745.800 588.600 747.600 594.600 ;
        RECT 748.800 593.700 756.600 595.050 ;
        RECT 748.800 588.600 750.600 593.700 ;
        RECT 754.800 588.600 756.600 593.700 ;
        RECT 764.400 591.600 765.600 603.900 ;
        RECT 767.100 602.100 768.900 602.850 ;
        RECT 773.100 602.100 774.900 602.850 ;
        RECT 766.950 598.950 769.050 601.050 ;
        RECT 772.950 598.950 775.050 601.050 ;
        RECT 763.800 588.600 765.600 591.600 ;
        RECT 776.400 591.600 777.600 603.900 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 794.100 600.150 795.900 600.900 ;
        RECT 797.400 598.650 798.300 606.900 ;
        RECT 794.100 597.000 798.300 598.650 ;
        RECT 809.700 598.650 810.600 606.900 ;
        RECT 814.950 604.950 817.050 607.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 812.100 600.150 813.900 600.900 ;
        RECT 809.700 597.000 813.900 598.650 ;
        RECT 776.400 588.600 778.200 591.600 ;
        RECT 794.100 588.600 795.900 597.000 ;
        RECT 812.100 588.600 813.900 597.000 ;
        RECT 12.000 580.050 13.800 584.400 ;
        RECT 8.400 578.400 13.800 580.050 ;
        RECT 8.400 575.100 9.300 578.400 ;
        RECT 29.100 576.000 30.900 584.400 ;
        RECT 48.000 580.050 49.800 584.400 ;
        RECT 26.700 574.350 30.900 576.000 ;
        RECT 44.400 578.400 49.800 580.050 ;
        RECT 44.400 575.100 45.300 578.400 ;
        RECT 63.000 577.200 64.800 584.400 ;
        RECT 84.000 580.050 85.800 584.400 ;
        RECT 80.400 578.400 85.800 580.050 ;
        RECT 63.000 576.300 66.600 577.200 ;
        RECT 7.950 571.950 10.050 574.050 ;
        RECT 13.950 571.950 16.050 574.050 ;
        RECT 8.400 561.600 9.300 570.900 ;
        RECT 14.100 570.150 15.900 570.900 ;
        RECT 11.100 569.100 12.900 569.850 ;
        RECT 17.100 569.100 18.900 569.850 ;
        RECT 10.950 565.950 13.050 568.050 ;
        RECT 16.950 565.950 19.050 568.050 ;
        RECT 26.700 566.100 27.600 574.350 ;
        RECT 34.950 573.450 37.050 574.200 ;
        RECT 43.950 573.450 46.050 574.050 ;
        RECT 29.100 572.100 30.900 572.850 ;
        RECT 34.950 572.550 46.050 573.450 ;
        RECT 34.950 572.100 37.050 572.550 ;
        RECT 43.950 571.950 46.050 572.550 ;
        RECT 49.950 571.950 52.050 574.050 ;
        RECT 65.400 572.100 66.600 576.300 ;
        RECT 80.400 575.100 81.300 578.400 ;
        RECT 104.100 576.000 105.900 584.400 ;
        RECT 120.300 580.200 122.100 584.400 ;
        RECT 101.700 574.350 105.900 576.000 ;
        RECT 120.150 578.400 122.100 580.200 ;
        RECT 120.150 575.100 121.050 578.400 ;
        RECT 122.100 576.600 123.900 577.500 ;
        RECT 127.800 576.600 129.600 584.400 ;
        RECT 122.100 575.700 129.600 576.600 ;
        RECT 138.000 577.200 139.800 584.400 ;
        RECT 154.500 578.400 156.300 584.400 ;
        RECT 160.800 581.400 162.600 584.400 ;
        RECT 138.000 576.300 141.600 577.200 ;
        RECT 79.950 571.800 82.050 574.050 ;
        RECT 85.950 573.450 88.050 574.050 ;
        RECT 97.950 573.450 100.050 574.050 ;
        RECT 85.950 572.550 100.050 573.450 ;
        RECT 85.950 571.950 88.050 572.550 ;
        RECT 97.950 571.950 100.050 572.550 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 565.950 34.050 568.050 ;
        RECT 22.950 562.950 28.050 565.050 ;
        RECT 32.100 564.150 33.900 564.900 ;
        RECT 35.100 563.100 36.900 563.850 ;
        RECT 7.800 549.600 9.600 561.600 ;
        RECT 10.800 560.700 18.600 561.600 ;
        RECT 10.800 549.600 12.600 560.700 ;
        RECT 16.800 549.600 18.600 560.700 ;
        RECT 26.700 556.800 27.600 561.900 ;
        RECT 34.950 559.950 37.050 562.050 ;
        RECT 44.400 561.600 45.300 570.900 ;
        RECT 50.100 570.150 51.900 570.900 ;
        RECT 47.100 569.100 48.900 569.850 ;
        RECT 53.100 569.100 54.900 569.850 ;
        RECT 64.950 568.950 67.050 571.050 ;
        RECT 46.950 565.950 49.050 568.050 ;
        RECT 52.950 565.950 55.050 568.050 ;
        RECT 62.100 566.100 63.900 566.850 ;
        RECT 61.950 562.950 64.050 565.050 ;
        RECT 26.700 555.900 33.300 556.800 ;
        RECT 26.700 555.600 27.600 555.900 ;
        RECT 25.800 549.600 27.600 555.600 ;
        RECT 31.800 555.600 33.300 555.900 ;
        RECT 31.800 549.600 33.600 555.600 ;
        RECT 43.800 549.600 45.600 561.600 ;
        RECT 46.800 560.700 54.600 561.600 ;
        RECT 46.800 549.600 48.600 560.700 ;
        RECT 52.800 549.600 54.600 560.700 ;
        RECT 65.400 555.600 66.600 567.900 ;
        RECT 68.100 566.100 69.900 566.850 ;
        RECT 67.950 562.950 70.050 565.050 ;
        RECT 80.400 561.600 81.300 570.900 ;
        RECT 86.100 570.150 87.900 570.900 ;
        RECT 83.100 569.100 84.900 569.850 ;
        RECT 89.100 569.100 90.900 569.850 ;
        RECT 82.950 565.950 85.050 568.050 ;
        RECT 88.950 565.950 91.050 568.050 ;
        RECT 101.700 566.100 102.600 574.350 ;
        RECT 104.100 572.100 105.900 572.850 ;
        RECT 115.950 571.950 124.050 574.050 ;
        RECT 103.950 568.950 106.050 571.050 ;
        RECT 106.950 565.950 109.050 568.050 ;
        RECT 98.550 564.900 103.050 565.050 ;
        RECT 97.950 562.950 103.050 564.900 ;
        RECT 107.100 564.150 108.900 564.900 ;
        RECT 110.100 563.100 111.900 563.850 ;
        RECT 97.950 562.800 100.050 562.950 ;
        RECT 64.800 549.600 66.600 555.600 ;
        RECT 79.800 549.600 81.600 561.600 ;
        RECT 82.800 560.700 90.600 561.600 ;
        RECT 82.800 549.600 84.600 560.700 ;
        RECT 88.800 549.600 90.600 560.700 ;
        RECT 101.700 556.800 102.600 561.900 ;
        RECT 109.950 559.950 112.050 562.050 ;
        RECT 118.950 561.600 120.000 570.900 ;
        RECT 122.100 569.100 123.900 569.850 ;
        RECT 121.950 565.950 124.050 568.050 ;
        RECT 101.700 555.900 108.300 556.800 ;
        RECT 101.700 555.600 102.600 555.900 ;
        RECT 100.800 549.600 102.600 555.600 ;
        RECT 106.800 555.600 108.300 555.900 ;
        RECT 106.800 549.600 108.600 555.600 ;
        RECT 118.200 549.600 120.000 561.600 ;
        RECT 125.550 555.600 126.600 575.700 ;
        RECT 140.400 572.100 141.600 576.300 ;
        RECT 154.800 575.100 156.000 578.400 ;
        RECT 160.800 577.500 162.000 581.400 ;
        RECT 156.900 576.600 162.000 577.500 ;
        RECT 170.400 576.600 172.200 584.400 ;
        RECT 177.900 580.200 179.700 584.400 ;
        RECT 177.900 578.400 179.850 580.200 ;
        RECT 176.100 576.600 177.900 577.500 ;
        RECT 156.900 575.700 158.850 576.600 ;
        RECT 170.400 575.700 177.900 576.600 ;
        RECT 157.950 575.100 158.850 575.700 ;
        RECT 145.950 573.450 148.050 574.050 ;
        RECT 154.950 573.450 157.050 574.050 ;
        RECT 145.950 572.550 157.050 573.450 ;
        RECT 145.950 571.950 148.050 572.550 ;
        RECT 154.950 571.950 157.050 572.550 ;
        RECT 127.950 568.950 130.050 571.050 ;
        RECT 139.950 570.450 142.050 571.050 ;
        RECT 148.950 570.450 151.050 571.050 ;
        RECT 158.100 570.900 158.850 575.100 ;
        RECT 139.950 569.550 151.050 570.450 ;
        RECT 139.950 568.950 142.050 569.550 ;
        RECT 148.950 568.950 151.050 569.550 ;
        RECT 128.100 567.150 129.900 567.900 ;
        RECT 137.100 566.100 138.900 566.850 ;
        RECT 136.950 562.950 139.050 565.050 ;
        RECT 140.400 555.600 141.600 567.900 ;
        RECT 143.100 566.100 144.900 566.850 ;
        RECT 142.950 562.950 145.050 565.050 ;
        RECT 154.800 561.600 156.000 570.900 ;
        RECT 157.950 564.300 158.850 570.900 ;
        RECT 169.950 568.950 172.050 571.050 ;
        RECT 161.100 567.150 162.900 567.900 ;
        RECT 170.100 567.150 171.900 567.900 ;
        RECT 156.900 563.400 158.850 564.300 ;
        RECT 156.900 562.500 162.600 563.400 ;
        RECT 124.800 549.600 126.600 555.600 ;
        RECT 139.800 549.600 141.600 555.600 ;
        RECT 154.500 549.600 156.300 561.600 ;
        RECT 161.400 555.600 162.600 562.500 ;
        RECT 160.800 549.600 162.600 555.600 ;
        RECT 173.400 555.600 174.450 575.700 ;
        RECT 178.950 575.100 179.850 578.400 ;
        RECT 192.000 577.200 193.800 584.400 ;
        RECT 206.400 579.300 208.200 584.400 ;
        RECT 212.400 579.300 214.200 584.400 ;
        RECT 206.400 577.950 214.200 579.300 ;
        RECT 215.400 578.400 217.200 584.400 ;
        RECT 192.000 576.300 195.600 577.200 ;
        RECT 215.400 576.300 216.600 578.400 ;
        RECT 232.200 577.200 234.000 584.400 ;
        RECT 247.800 578.400 249.600 584.400 ;
        RECT 225.000 576.450 229.050 577.050 ;
        RECT 178.950 573.450 181.050 574.050 ;
        RECT 187.950 573.450 190.050 574.050 ;
        RECT 178.950 572.550 190.050 573.450 ;
        RECT 178.950 571.950 181.050 572.550 ;
        RECT 187.950 571.950 190.050 572.550 ;
        RECT 194.400 572.100 195.600 576.300 ;
        RECT 212.850 575.250 216.600 576.300 ;
        RECT 212.850 575.100 214.050 575.250 ;
        RECT 224.550 574.950 229.050 576.450 ;
        RECT 230.400 576.300 234.000 577.200 ;
        RECT 248.400 576.300 249.600 578.400 ;
        RECT 250.800 579.300 252.600 584.400 ;
        RECT 256.800 579.300 258.600 584.400 ;
        RECT 250.800 577.950 258.600 579.300 ;
        RECT 266.400 578.400 268.200 584.400 ;
        RECT 278.400 578.400 280.200 584.400 ;
        RECT 289.800 578.400 291.600 584.400 ;
        RECT 202.950 571.950 208.050 574.050 ;
        RECT 211.950 573.450 214.050 574.050 ;
        RECT 224.550 573.450 225.450 574.950 ;
        RECT 211.950 572.550 225.450 573.450 ;
        RECT 211.950 571.950 214.050 572.550 ;
        RECT 230.400 572.100 231.600 576.300 ;
        RECT 248.400 575.250 252.150 576.300 ;
        RECT 250.950 575.100 252.150 575.250 ;
        RECT 266.400 575.100 267.600 578.400 ;
        RECT 278.400 575.100 279.600 578.400 ;
        RECT 290.400 575.100 291.600 578.400 ;
        RECT 302.400 576.600 304.200 584.400 ;
        RECT 309.900 580.200 311.700 584.400 ;
        RECT 309.900 578.400 311.850 580.200 ;
        RECT 325.800 578.400 327.600 584.400 ;
        RECT 308.100 576.600 309.900 577.500 ;
        RECT 302.400 575.700 309.900 576.600 ;
        RECT 250.950 571.950 253.050 574.050 ;
        RECT 256.950 571.950 259.050 574.050 ;
        RECT 265.950 571.950 268.050 574.050 ;
        RECT 277.950 571.950 280.050 574.050 ;
        RECT 283.950 573.450 288.000 574.050 ;
        RECT 289.950 573.450 292.050 574.050 ;
        RECT 283.950 572.550 292.050 573.450 ;
        RECT 283.950 571.950 288.000 572.550 ;
        RECT 289.950 571.950 292.050 572.550 ;
        RECT 176.100 569.100 177.900 569.850 ;
        RECT 180.000 561.600 181.050 570.900 ;
        RECT 193.950 568.950 199.050 571.050 ;
        RECT 206.100 570.150 207.900 570.900 ;
        RECT 209.100 569.100 210.900 569.850 ;
        RECT 211.950 569.100 213.150 570.900 ;
        RECT 223.950 570.450 228.000 571.050 ;
        RECT 229.950 570.450 232.050 571.050 ;
        RECT 215.100 569.100 216.900 569.850 ;
        RECT 223.950 569.550 232.050 570.450 ;
        RECT 191.100 566.100 192.900 566.850 ;
        RECT 190.950 562.950 193.050 565.050 ;
        RECT 173.400 549.600 175.200 555.600 ;
        RECT 180.000 549.600 181.800 561.600 ;
        RECT 194.400 555.600 195.600 567.900 ;
        RECT 197.100 566.100 198.900 566.850 ;
        RECT 208.950 565.950 211.050 568.050 ;
        RECT 196.950 562.950 199.050 565.050 ;
        RECT 212.100 564.900 213.150 569.100 ;
        RECT 223.950 568.950 228.000 569.550 ;
        RECT 229.950 568.950 232.050 569.550 ;
        RECT 248.100 569.100 249.900 569.850 ;
        RECT 251.850 569.100 253.050 570.900 ;
        RECT 257.100 570.150 258.900 570.900 ;
        RECT 254.100 569.100 255.900 569.850 ;
        RECT 263.100 569.100 264.900 569.850 ;
        RECT 214.950 565.950 217.050 568.050 ;
        RECT 227.100 566.100 228.900 566.850 ;
        RECT 211.950 561.600 213.150 564.900 ;
        RECT 226.950 562.950 229.050 565.050 ;
        RECT 193.800 549.600 195.600 555.600 ;
        RECT 211.500 549.600 213.300 561.600 ;
        RECT 230.400 555.600 231.600 567.900 ;
        RECT 233.100 566.100 234.900 566.850 ;
        RECT 247.950 565.950 250.050 568.050 ;
        RECT 251.850 564.900 252.900 569.100 ;
        RECT 253.950 565.950 256.050 568.050 ;
        RECT 251.850 561.600 253.050 564.900 ;
        RECT 266.400 561.600 267.600 570.900 ;
        RECT 275.100 569.100 276.900 569.850 ;
        RECT 278.400 561.600 279.600 570.900 ;
        RECT 290.400 561.600 291.600 570.900 ;
        RECT 293.100 569.100 294.900 569.850 ;
        RECT 301.950 568.950 304.050 571.050 ;
        RECT 292.950 565.950 298.050 568.050 ;
        RECT 302.100 567.150 303.900 567.900 ;
        RECT 230.400 549.600 232.200 555.600 ;
        RECT 251.700 549.600 253.500 561.600 ;
        RECT 266.400 549.600 268.200 561.600 ;
        RECT 278.400 549.600 280.200 561.600 ;
        RECT 289.800 549.600 291.600 561.600 ;
        RECT 305.400 555.600 306.450 575.700 ;
        RECT 310.950 575.100 311.850 578.400 ;
        RECT 326.400 576.300 327.600 578.400 ;
        RECT 328.800 579.300 330.600 584.400 ;
        RECT 334.800 579.300 336.600 584.400 ;
        RECT 328.800 577.950 336.600 579.300 ;
        RECT 348.000 577.200 349.800 584.400 ;
        RECT 361.800 578.400 363.600 584.400 ;
        RECT 348.000 576.300 351.600 577.200 ;
        RECT 326.400 575.250 330.150 576.300 ;
        RECT 328.950 575.100 330.150 575.250 ;
        RECT 310.950 573.450 313.050 574.050 ;
        RECT 322.950 573.450 325.050 574.050 ;
        RECT 310.950 572.550 325.050 573.450 ;
        RECT 310.950 571.950 313.050 572.550 ;
        RECT 322.950 571.950 325.050 572.550 ;
        RECT 328.950 571.950 331.050 574.050 ;
        RECT 334.950 571.950 337.050 574.050 ;
        RECT 350.400 572.100 351.600 576.300 ;
        RECT 362.400 576.300 363.600 578.400 ;
        RECT 364.800 579.300 366.600 584.400 ;
        RECT 370.800 579.300 372.600 584.400 ;
        RECT 384.300 580.200 386.100 584.400 ;
        RECT 364.800 577.950 372.600 579.300 ;
        RECT 384.150 578.400 386.100 580.200 ;
        RECT 362.400 575.250 366.150 576.300 ;
        RECT 364.950 575.100 366.150 575.250 ;
        RECT 384.150 575.100 385.050 578.400 ;
        RECT 386.100 576.600 387.900 577.500 ;
        RECT 391.800 576.600 393.600 584.400 ;
        RECT 400.800 578.400 402.600 584.400 ;
        RECT 386.100 575.700 393.600 576.600 ;
        RECT 401.400 576.300 402.600 578.400 ;
        RECT 403.800 579.300 405.600 584.400 ;
        RECT 409.800 579.300 411.600 584.400 ;
        RECT 403.800 577.950 411.600 579.300 ;
        RECT 420.000 577.200 421.800 584.400 ;
        RECT 436.800 578.400 438.600 584.400 ;
        RECT 420.000 576.300 423.600 577.200 ;
        RECT 364.950 571.950 367.050 574.050 ;
        RECT 370.950 571.950 373.050 574.050 ;
        RECT 382.950 571.950 385.050 574.050 ;
        RECT 308.100 569.100 309.900 569.850 ;
        RECT 312.000 561.600 313.050 570.900 ;
        RECT 326.100 569.100 327.900 569.850 ;
        RECT 329.850 569.100 331.050 570.900 ;
        RECT 335.100 570.150 336.900 570.900 ;
        RECT 343.950 570.450 348.000 571.050 ;
        RECT 349.950 570.450 352.050 571.050 ;
        RECT 332.100 569.100 333.900 569.850 ;
        RECT 343.950 569.550 352.050 570.450 ;
        RECT 325.950 565.950 328.050 568.050 ;
        RECT 329.850 564.900 330.900 569.100 ;
        RECT 343.950 568.950 348.000 569.550 ;
        RECT 349.950 568.950 352.050 569.550 ;
        RECT 362.100 569.100 363.900 569.850 ;
        RECT 365.850 569.100 367.050 570.900 ;
        RECT 371.100 570.150 372.900 570.900 ;
        RECT 368.100 569.100 369.900 569.850 ;
        RECT 331.950 567.450 334.050 568.050 ;
        RECT 336.000 567.450 340.050 568.050 ;
        RECT 331.950 566.550 340.050 567.450 ;
        RECT 331.950 565.950 334.050 566.550 ;
        RECT 336.000 565.950 340.050 566.550 ;
        RECT 347.100 566.100 348.900 566.850 ;
        RECT 329.850 561.600 331.050 564.900 ;
        RECT 346.950 562.950 349.050 565.050 ;
        RECT 305.400 549.600 307.200 555.600 ;
        RECT 312.000 549.600 313.800 561.600 ;
        RECT 329.700 549.600 331.500 561.600 ;
        RECT 350.400 555.600 351.600 567.900 ;
        RECT 353.100 566.100 354.900 566.850 ;
        RECT 361.950 565.950 364.050 568.050 ;
        RECT 352.950 562.800 355.050 565.050 ;
        RECT 365.850 564.900 366.900 569.100 ;
        RECT 367.950 565.950 370.050 568.050 ;
        RECT 365.850 561.600 367.050 564.900 ;
        RECT 382.950 561.600 384.000 570.900 ;
        RECT 386.100 569.100 387.900 569.850 ;
        RECT 349.800 549.600 351.600 555.600 ;
        RECT 365.700 549.600 367.500 561.600 ;
        RECT 382.200 549.600 384.000 561.600 ;
        RECT 389.550 555.600 390.600 575.700 ;
        RECT 401.400 575.250 405.150 576.300 ;
        RECT 403.950 575.100 405.150 575.250 ;
        RECT 400.950 571.950 406.050 574.050 ;
        RECT 409.950 573.450 412.050 574.050 ;
        RECT 414.000 573.450 418.050 574.050 ;
        RECT 409.950 572.550 418.050 573.450 ;
        RECT 409.950 571.950 412.050 572.550 ;
        RECT 414.000 571.950 418.050 572.550 ;
        RECT 422.400 572.100 423.600 576.300 ;
        RECT 437.400 576.300 438.600 578.400 ;
        RECT 439.800 579.300 441.600 584.400 ;
        RECT 445.800 579.300 447.600 584.400 ;
        RECT 439.800 577.950 447.600 579.300 ;
        RECT 457.800 578.400 459.600 584.400 ;
        RECT 437.400 575.250 441.150 576.300 ;
        RECT 439.950 575.100 441.150 575.250 ;
        RECT 458.400 575.100 459.600 578.400 ;
        RECT 474.000 577.200 475.800 584.400 ;
        RECT 488.400 579.300 490.200 584.400 ;
        RECT 494.400 579.300 496.200 584.400 ;
        RECT 488.400 577.950 496.200 579.300 ;
        RECT 497.400 578.400 499.200 584.400 ;
        RECT 511.800 578.400 513.600 584.400 ;
        RECT 523.800 578.400 525.600 584.400 ;
        RECT 474.000 576.300 477.600 577.200 ;
        RECT 497.400 576.300 498.600 578.400 ;
        RECT 430.950 573.450 433.050 574.050 ;
        RECT 439.950 573.450 442.050 574.050 ;
        RECT 430.950 572.550 442.050 573.450 ;
        RECT 430.950 571.950 433.050 572.550 ;
        RECT 439.950 571.950 442.050 572.550 ;
        RECT 445.950 571.950 448.050 574.050 ;
        RECT 457.950 571.950 460.050 574.050 ;
        RECT 476.400 572.100 477.600 576.300 ;
        RECT 494.850 575.250 498.600 576.300 ;
        RECT 494.850 575.100 496.050 575.250 ;
        RECT 512.400 575.100 513.600 578.400 ;
        RECT 524.400 576.300 525.600 578.400 ;
        RECT 526.800 579.300 528.600 584.400 ;
        RECT 532.800 579.300 534.600 584.400 ;
        RECT 526.800 577.950 534.600 579.300 ;
        RECT 544.800 578.400 546.600 584.400 ;
        RECT 545.400 576.300 546.600 578.400 ;
        RECT 547.800 579.300 549.600 584.400 ;
        RECT 553.800 579.300 555.600 584.400 ;
        RECT 547.800 577.950 555.600 579.300 ;
        RECT 563.400 579.300 565.200 584.400 ;
        RECT 569.400 579.300 571.200 584.400 ;
        RECT 563.400 577.950 571.200 579.300 ;
        RECT 572.400 578.400 574.200 584.400 ;
        RECT 586.800 578.400 588.600 584.400 ;
        RECT 572.400 576.300 573.600 578.400 ;
        RECT 524.400 575.250 528.150 576.300 ;
        RECT 545.400 575.250 549.150 576.300 ;
        RECT 526.950 575.100 528.150 575.250 ;
        RECT 547.950 575.100 549.150 575.250 ;
        RECT 569.850 575.250 573.600 576.300 ;
        RECT 587.400 576.300 588.600 578.400 ;
        RECT 589.800 579.300 591.600 584.400 ;
        RECT 595.800 579.300 597.600 584.400 ;
        RECT 605.400 581.400 607.200 584.400 ;
        RECT 589.800 577.950 597.600 579.300 ;
        RECT 606.300 577.200 607.200 581.400 ;
        RECT 611.400 578.400 613.200 584.400 ;
        RECT 620.400 579.300 622.200 584.400 ;
        RECT 626.400 579.300 628.200 584.400 ;
        RECT 606.300 576.300 609.750 577.200 ;
        RECT 587.400 575.250 591.150 576.300 ;
        RECT 607.950 575.400 609.750 576.300 ;
        RECT 569.850 575.100 571.050 575.250 ;
        RECT 589.950 575.100 591.150 575.250 ;
        RECT 487.950 571.950 490.050 574.050 ;
        RECT 493.950 573.450 496.050 574.050 ;
        RECT 505.950 573.450 508.050 574.050 ;
        RECT 493.950 572.550 508.050 573.450 ;
        RECT 493.950 571.950 496.050 572.550 ;
        RECT 505.950 571.950 508.050 572.550 ;
        RECT 511.950 571.800 514.050 574.050 ;
        RECT 526.950 571.950 529.050 574.050 ;
        RECT 532.950 571.950 535.050 574.050 ;
        RECT 544.950 571.950 550.050 574.050 ;
        RECT 553.950 571.950 556.050 574.050 ;
        RECT 562.950 571.950 565.050 574.050 ;
        RECT 568.950 573.450 571.050 574.050 ;
        RECT 580.950 573.450 583.050 573.900 ;
        RECT 568.950 572.550 583.050 573.450 ;
        RECT 568.950 571.950 571.050 572.550 ;
        RECT 580.950 571.800 583.050 572.550 ;
        RECT 589.950 571.950 592.050 574.050 ;
        RECT 595.950 571.950 598.050 574.050 ;
        RECT 604.950 571.950 607.050 574.050 ;
        RECT 391.950 568.950 394.050 571.050 ;
        RECT 401.100 569.100 402.900 569.850 ;
        RECT 404.850 569.100 406.050 570.900 ;
        RECT 410.100 570.150 411.900 570.900 ;
        RECT 407.100 569.100 408.900 569.850 ;
        RECT 392.100 567.150 393.900 567.900 ;
        RECT 400.950 565.950 403.050 568.050 ;
        RECT 404.850 564.900 405.900 569.100 ;
        RECT 421.950 568.950 427.050 571.050 ;
        RECT 437.100 569.100 438.900 569.850 ;
        RECT 440.850 569.100 442.050 570.900 ;
        RECT 446.100 570.150 447.900 570.900 ;
        RECT 443.100 569.100 444.900 569.850 ;
        RECT 406.950 565.950 409.050 568.050 ;
        RECT 419.100 566.100 420.900 566.850 ;
        RECT 404.850 561.600 406.050 564.900 ;
        RECT 388.800 549.600 390.600 555.600 ;
        RECT 404.700 549.600 406.500 561.600 ;
        RECT 422.400 555.600 423.600 567.900 ;
        RECT 425.100 566.100 426.900 566.850 ;
        RECT 436.950 565.950 439.050 568.050 ;
        RECT 424.950 562.950 427.050 565.050 ;
        RECT 440.850 564.900 441.900 569.100 ;
        RECT 442.950 565.950 445.050 568.050 ;
        RECT 440.850 561.600 442.050 564.900 ;
        RECT 458.400 561.600 459.600 570.900 ;
        RECT 475.950 570.450 478.050 571.050 ;
        RECT 480.000 570.450 484.050 571.050 ;
        RECT 461.100 569.100 462.900 569.850 ;
        RECT 475.950 569.550 484.050 570.450 ;
        RECT 488.100 570.150 489.900 570.900 ;
        RECT 475.950 568.950 478.050 569.550 ;
        RECT 480.000 568.950 484.050 569.550 ;
        RECT 491.100 569.100 492.900 569.850 ;
        RECT 493.950 569.100 495.150 570.900 ;
        RECT 497.100 569.100 498.900 569.850 ;
        RECT 460.950 565.950 466.050 568.050 ;
        RECT 473.100 566.100 474.900 566.850 ;
        RECT 421.800 549.600 423.600 555.600 ;
        RECT 440.700 549.600 442.500 561.600 ;
        RECT 457.800 549.600 459.600 561.600 ;
        RECT 476.400 555.600 477.600 567.900 ;
        RECT 479.100 566.100 480.900 566.850 ;
        RECT 490.950 565.950 493.050 568.050 ;
        RECT 478.950 562.950 481.050 565.050 ;
        RECT 494.100 564.900 495.150 569.100 ;
        RECT 496.950 565.950 499.050 568.050 ;
        RECT 493.950 561.600 495.150 564.900 ;
        RECT 512.400 561.600 513.600 570.900 ;
        RECT 515.100 569.100 516.900 569.850 ;
        RECT 524.100 569.100 525.900 569.850 ;
        RECT 527.850 569.100 529.050 570.900 ;
        RECT 533.100 570.150 534.900 570.900 ;
        RECT 530.100 569.100 531.900 569.850 ;
        RECT 545.100 569.100 546.900 569.850 ;
        RECT 548.850 569.100 550.050 570.900 ;
        RECT 554.100 570.150 555.900 570.900 ;
        RECT 563.100 570.150 564.900 570.900 ;
        RECT 551.100 569.100 552.900 569.850 ;
        RECT 566.100 569.100 567.900 569.850 ;
        RECT 568.950 569.100 570.150 570.900 ;
        RECT 572.100 569.100 573.900 569.850 ;
        RECT 587.100 569.100 588.900 569.850 ;
        RECT 590.850 569.100 592.050 570.900 ;
        RECT 596.100 570.150 597.900 570.900 ;
        RECT 605.100 570.150 606.900 570.900 ;
        RECT 593.100 569.100 594.900 569.850 ;
        RECT 602.100 569.100 603.900 569.850 ;
        RECT 514.950 565.950 517.050 568.050 ;
        RECT 523.950 565.950 526.050 568.050 ;
        RECT 527.850 564.900 528.900 569.100 ;
        RECT 529.950 565.950 532.050 568.050 ;
        RECT 541.950 565.950 547.050 568.050 ;
        RECT 548.850 564.900 549.900 569.100 ;
        RECT 550.950 567.450 553.050 568.050 ;
        RECT 565.950 567.450 568.050 568.050 ;
        RECT 550.950 566.550 568.050 567.450 ;
        RECT 550.950 565.950 553.050 566.550 ;
        RECT 565.950 565.950 568.050 566.550 ;
        RECT 569.100 564.900 570.150 569.100 ;
        RECT 571.950 565.950 574.050 568.050 ;
        RECT 586.950 565.950 589.050 568.050 ;
        RECT 527.850 561.600 529.050 564.900 ;
        RECT 548.850 561.600 550.050 564.900 ;
        RECT 568.950 561.600 570.150 564.900 ;
        RECT 590.850 564.900 591.900 569.100 ;
        RECT 592.950 565.950 595.050 568.050 ;
        RECT 601.950 565.950 604.050 568.050 ;
        RECT 590.850 561.600 592.050 564.900 ;
        RECT 608.700 564.600 609.600 575.400 ;
        RECT 612.000 572.100 613.050 578.400 ;
        RECT 620.400 577.950 628.200 579.300 ;
        RECT 629.400 578.400 631.200 584.400 ;
        RECT 629.400 576.300 630.600 578.400 ;
        RECT 643.200 577.200 645.000 584.400 ;
        RECT 656.400 579.300 658.200 584.400 ;
        RECT 662.400 579.300 664.200 584.400 ;
        RECT 656.400 577.950 664.200 579.300 ;
        RECT 665.400 578.400 667.200 584.400 ;
        RECT 677.400 581.400 679.200 584.400 ;
        RECT 626.850 575.250 630.600 576.300 ;
        RECT 641.400 576.300 645.000 577.200 ;
        RECT 665.400 576.300 666.600 578.400 ;
        RECT 678.000 577.500 679.200 581.400 ;
        RECT 683.700 578.400 685.500 584.400 ;
        RECT 678.000 576.600 683.100 577.500 ;
        RECT 626.850 575.100 628.050 575.250 ;
        RECT 619.950 571.950 622.050 574.050 ;
        RECT 625.950 573.450 628.050 574.050 ;
        RECT 634.950 573.450 637.050 574.050 ;
        RECT 625.950 572.550 637.050 573.450 ;
        RECT 625.950 571.950 628.050 572.550 ;
        RECT 634.950 571.950 637.050 572.550 ;
        RECT 641.400 572.100 642.600 576.300 ;
        RECT 662.850 575.250 666.600 576.300 ;
        RECT 681.150 575.700 683.100 576.600 ;
        RECT 662.850 575.100 664.050 575.250 ;
        RECT 681.150 575.100 682.050 575.700 ;
        RECT 684.000 575.100 685.200 578.400 ;
        RECT 697.200 577.200 699.000 584.400 ;
        RECT 715.800 581.400 717.600 584.400 ;
        RECT 716.400 578.100 717.600 581.400 ;
        RECT 695.400 576.300 699.000 577.200 ;
        RECT 655.950 571.950 658.050 574.050 ;
        RECT 661.950 571.950 667.050 574.050 ;
        RECT 610.950 568.950 616.050 571.050 ;
        RECT 620.100 570.150 621.900 570.900 ;
        RECT 623.100 569.100 624.900 569.850 ;
        RECT 625.950 569.100 627.150 570.900 ;
        RECT 640.950 570.450 643.050 571.050 ;
        RECT 649.950 570.450 652.050 571.050 ;
        RECT 629.100 569.100 630.900 569.850 ;
        RECT 640.950 569.550 652.050 570.450 ;
        RECT 656.100 570.150 657.900 570.900 ;
        RECT 607.800 564.000 609.600 564.600 ;
        RECT 602.400 562.800 609.600 564.000 ;
        RECT 602.400 561.600 603.600 562.800 ;
        RECT 610.950 561.600 612.300 567.900 ;
        RECT 622.950 565.950 625.050 568.050 ;
        RECT 626.100 564.900 627.150 569.100 ;
        RECT 640.950 568.950 643.050 569.550 ;
        RECT 649.950 568.950 652.050 569.550 ;
        RECT 659.100 569.100 660.900 569.850 ;
        RECT 661.950 569.100 663.150 570.900 ;
        RECT 670.950 570.450 675.000 571.050 ;
        RECT 676.950 570.450 679.050 571.050 ;
        RECT 665.100 569.100 666.900 569.850 ;
        RECT 670.950 569.550 679.050 570.450 ;
        RECT 628.950 565.950 631.050 568.050 ;
        RECT 638.100 566.100 639.900 566.850 ;
        RECT 625.950 561.600 627.150 564.900 ;
        RECT 634.950 562.950 640.050 565.050 ;
        RECT 475.800 549.600 477.600 555.600 ;
        RECT 493.500 549.600 495.300 561.600 ;
        RECT 511.800 549.600 513.600 561.600 ;
        RECT 527.700 549.600 529.500 561.600 ;
        RECT 548.700 549.600 550.500 561.600 ;
        RECT 568.500 549.600 570.300 561.600 ;
        RECT 590.700 549.600 592.500 561.600 ;
        RECT 602.400 549.600 604.200 561.600 ;
        RECT 609.900 560.100 612.300 561.600 ;
        RECT 609.900 549.600 611.700 560.100 ;
        RECT 625.500 549.600 627.300 561.600 ;
        RECT 641.400 555.600 642.600 567.900 ;
        RECT 644.100 566.100 645.900 566.850 ;
        RECT 658.950 565.950 661.050 568.050 ;
        RECT 643.950 562.950 646.050 565.050 ;
        RECT 662.100 564.900 663.150 569.100 ;
        RECT 670.950 568.950 675.000 569.550 ;
        RECT 676.950 568.950 679.050 569.550 ;
        RECT 681.150 570.900 681.900 575.100 ;
        RECT 695.400 572.100 696.600 576.300 ;
        RECT 712.950 574.950 718.050 577.050 ;
        RECT 725.400 576.600 727.200 584.400 ;
        RECT 732.900 580.200 734.700 584.400 ;
        RECT 748.800 581.400 750.600 584.400 ;
        RECT 732.900 578.400 734.850 580.200 ;
        RECT 731.100 576.600 732.900 577.500 ;
        RECT 725.400 575.700 732.900 576.600 ;
        RECT 715.950 572.100 717.300 573.900 ;
        RECT 664.950 565.950 667.050 568.050 ;
        RECT 677.100 567.150 678.900 567.900 ;
        RECT 661.950 561.600 663.150 564.900 ;
        RECT 681.150 564.300 682.050 570.900 ;
        RECT 681.150 563.400 683.100 564.300 ;
        RECT 677.400 562.500 683.100 563.400 ;
        RECT 641.400 549.600 643.200 555.600 ;
        RECT 661.500 549.600 663.300 561.600 ;
        RECT 677.400 555.600 678.600 562.500 ;
        RECT 684.000 561.600 685.200 570.900 ;
        RECT 694.950 570.450 697.050 571.050 ;
        RECT 706.950 570.450 709.050 571.050 ;
        RECT 694.950 569.550 709.050 570.450 ;
        RECT 694.950 568.950 697.050 569.550 ;
        RECT 706.950 568.950 709.050 569.550 ;
        RECT 712.950 568.950 715.050 571.050 ;
        RECT 716.100 567.900 717.300 572.100 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 692.100 566.100 693.900 566.850 ;
        RECT 691.950 562.950 694.050 565.050 ;
        RECT 677.400 549.600 679.200 555.600 ;
        RECT 683.700 549.600 685.500 561.600 ;
        RECT 695.400 555.600 696.600 567.900 ;
        RECT 713.100 567.150 714.900 567.900 ;
        RECT 698.100 566.100 699.900 566.850 ;
        RECT 697.950 562.950 700.050 565.050 ;
        RECT 715.950 562.650 717.300 567.900 ;
        RECT 718.950 565.950 721.050 568.050 ;
        RECT 725.100 567.150 726.900 567.900 ;
        RECT 719.100 564.150 720.900 564.900 ;
        RECT 714.600 561.600 717.300 562.650 ;
        RECT 695.400 549.600 697.200 555.600 ;
        RECT 714.600 549.600 716.400 561.600 ;
        RECT 728.400 555.600 729.450 575.700 ;
        RECT 733.950 575.100 734.850 578.400 ;
        RECT 733.950 571.950 739.050 574.050 ;
        RECT 731.100 569.100 732.900 569.850 ;
        RECT 730.950 565.950 733.050 568.050 ;
        RECT 735.000 561.600 736.050 570.900 ;
        RECT 749.400 569.100 750.600 581.400 ;
        RECT 764.400 581.400 766.200 584.400 ;
        RECT 779.400 581.400 781.200 584.400 ;
        RECT 794.400 581.400 796.200 584.400 ;
        RECT 812.400 581.400 814.200 584.400 ;
        RECT 751.950 571.950 754.050 574.050 ;
        RECT 760.950 571.950 763.050 574.050 ;
        RECT 752.100 570.150 753.900 570.900 ;
        RECT 761.100 570.150 762.900 570.900 ;
        RECT 764.400 569.100 765.600 581.400 ;
        RECT 779.400 578.100 780.600 581.400 ;
        RECT 794.400 578.100 795.600 581.400 ;
        RECT 812.400 578.100 813.600 581.400 ;
        RECT 766.950 576.450 769.050 577.050 ;
        RECT 778.950 576.450 781.050 577.050 ;
        RECT 766.950 575.550 781.050 576.450 ;
        RECT 766.950 574.950 769.050 575.550 ;
        RECT 778.950 574.950 781.050 575.550 ;
        RECT 790.950 574.950 796.050 577.050 ;
        RECT 811.950 576.450 814.050 577.050 ;
        RECT 816.000 576.450 820.050 577.050 ;
        RECT 811.950 575.550 820.050 576.450 ;
        RECT 811.950 574.950 814.050 575.550 ;
        RECT 816.000 574.950 820.050 575.550 ;
        RECT 779.700 572.100 781.050 573.900 ;
        RECT 794.700 572.100 796.050 573.900 ;
        RECT 812.700 572.100 814.050 573.900 ;
        RECT 748.950 565.950 751.050 568.050 ;
        RECT 763.950 567.450 766.050 568.050 ;
        RECT 768.000 567.450 772.050 568.050 ;
        RECT 763.950 566.550 772.050 567.450 ;
        RECT 763.950 565.950 766.050 566.550 ;
        RECT 768.000 565.950 772.050 566.550 ;
        RECT 775.950 565.950 778.050 568.050 ;
        RECT 779.700 567.900 780.900 572.100 ;
        RECT 781.950 568.950 784.050 571.050 ;
        RECT 728.400 549.600 730.200 555.600 ;
        RECT 735.000 549.600 736.800 561.600 ;
        RECT 749.400 555.600 750.600 564.900 ;
        RECT 748.800 549.600 750.600 555.600 ;
        RECT 764.400 555.600 765.600 564.900 ;
        RECT 776.100 564.150 777.900 564.900 ;
        RECT 779.700 562.650 781.050 567.900 ;
        RECT 782.100 567.150 783.900 567.900 ;
        RECT 790.950 565.800 793.050 568.050 ;
        RECT 794.700 567.900 795.900 572.100 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 791.100 564.150 792.900 564.900 ;
        RECT 794.700 562.650 796.050 567.900 ;
        RECT 797.100 567.150 798.900 567.900 ;
        RECT 808.950 565.950 811.050 568.050 ;
        RECT 812.700 567.900 813.900 572.100 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 809.100 564.150 810.900 564.900 ;
        RECT 812.700 562.650 814.050 567.900 ;
        RECT 815.100 567.150 816.900 567.900 ;
        RECT 779.700 561.600 782.400 562.650 ;
        RECT 794.700 561.600 797.400 562.650 ;
        RECT 812.700 561.600 815.400 562.650 ;
        RECT 764.400 549.600 766.200 555.600 ;
        RECT 780.600 549.600 782.400 561.600 ;
        RECT 795.600 549.600 797.400 561.600 ;
        RECT 813.600 549.600 815.400 561.600 ;
        RECT 10.800 533.400 12.600 545.400 ;
        RECT 13.800 534.300 15.600 545.400 ;
        RECT 19.800 534.300 21.600 545.400 ;
        RECT 32.400 539.400 34.200 545.400 ;
        RECT 32.700 539.100 34.200 539.400 ;
        RECT 38.400 539.400 40.200 545.400 ;
        RECT 49.800 539.400 51.600 545.400 ;
        RECT 38.400 539.100 39.300 539.400 ;
        RECT 32.700 538.200 39.300 539.100 ;
        RECT 13.800 533.400 21.600 534.300 ;
        RECT 11.400 524.100 12.300 533.400 ;
        RECT 25.950 532.950 31.050 535.050 ;
        RECT 38.400 533.100 39.300 538.200 ;
        RECT 29.100 531.150 30.900 531.900 ;
        RECT 32.100 530.100 33.900 530.850 ;
        RECT 37.950 529.950 40.050 532.050 ;
        RECT 50.400 530.100 51.600 539.400 ;
        RECT 68.700 533.400 70.500 545.400 ;
        RECT 85.500 533.400 87.300 545.400 ;
        RECT 107.700 533.400 109.500 545.400 ;
        RECT 124.500 533.400 126.300 545.400 ;
        RECT 145.800 539.400 147.600 545.400 ;
        RECT 68.850 530.100 70.050 533.400 ;
        RECT 85.950 530.100 87.150 533.400 ;
        RECT 13.950 526.950 16.050 529.050 ;
        RECT 19.950 526.950 22.050 529.050 ;
        RECT 31.950 526.950 34.050 529.200 ;
        RECT 14.100 525.150 15.900 525.900 ;
        RECT 20.100 525.150 21.900 525.900 ;
        RECT 17.100 524.100 18.900 524.850 ;
        RECT 34.950 523.950 37.050 526.050 ;
        RECT 4.950 522.450 9.000 523.050 ;
        RECT 10.950 522.450 13.050 523.050 ;
        RECT 4.950 521.550 13.050 522.450 ;
        RECT 4.950 520.950 9.000 521.550 ;
        RECT 10.950 520.950 13.050 521.550 ;
        RECT 16.950 520.950 19.050 523.050 ;
        RECT 35.100 522.150 36.900 522.900 ;
        RECT 38.400 520.650 39.300 528.900 ;
        RECT 46.950 526.950 52.050 529.050 ;
        RECT 64.950 526.950 67.050 529.050 ;
        RECT 68.850 525.900 69.900 530.100 ;
        RECT 70.950 526.950 73.050 529.050 ;
        RECT 82.950 526.950 85.050 529.050 ;
        RECT 86.100 525.900 87.150 530.100 ;
        RECT 107.850 530.100 109.050 533.400 ;
        RECT 124.950 530.100 126.150 533.400 ;
        RECT 88.950 526.950 91.050 529.050 ;
        RECT 103.950 526.950 106.050 529.050 ;
        RECT 107.850 525.900 108.900 530.100 ;
        RECT 109.950 528.450 112.050 529.050 ;
        RECT 114.000 528.900 117.000 529.050 ;
        RECT 114.000 528.450 118.050 528.900 ;
        RECT 109.950 527.550 118.050 528.450 ;
        RECT 109.950 526.950 112.050 527.550 ;
        RECT 114.000 526.950 118.050 527.550 ;
        RECT 121.950 526.950 124.050 529.050 ;
        RECT 115.950 526.800 118.050 526.950 ;
        RECT 125.100 525.900 126.150 530.100 ;
        RECT 142.950 529.950 145.050 532.050 ;
        RECT 127.950 526.950 130.050 529.050 ;
        RECT 143.100 528.150 144.900 528.900 ;
        RECT 146.400 527.100 147.600 539.400 ;
        RECT 148.950 537.450 151.050 538.050 ;
        RECT 154.950 537.450 157.050 538.050 ;
        RECT 148.950 536.550 157.050 537.450 ;
        RECT 148.950 535.950 151.050 536.550 ;
        RECT 154.950 535.950 157.050 536.550 ;
        RECT 160.800 533.400 162.600 545.400 ;
        RECT 163.800 534.300 165.600 545.400 ;
        RECT 169.800 534.300 171.600 545.400 ;
        RECT 163.800 533.400 171.600 534.300 ;
        RECT 185.700 533.400 187.500 545.400 ;
        RECT 203.400 539.400 205.200 545.400 ;
        RECT 148.950 529.950 151.050 532.050 ;
        RECT 149.100 528.150 150.900 528.900 ;
        RECT 11.400 516.600 12.300 519.900 ;
        RECT 35.100 519.000 39.300 520.650 ;
        RECT 11.400 514.950 16.800 516.600 ;
        RECT 15.000 510.600 16.800 514.950 ;
        RECT 35.100 510.600 36.900 519.000 ;
        RECT 50.400 513.600 51.600 525.900 ;
        RECT 65.100 525.150 66.900 525.900 ;
        RECT 53.100 524.100 54.900 524.850 ;
        RECT 68.850 524.100 70.050 525.900 ;
        RECT 71.100 525.150 72.900 525.900 ;
        RECT 83.100 525.150 84.900 525.900 ;
        RECT 74.100 524.100 75.900 524.850 ;
        RECT 80.100 524.100 81.900 524.850 ;
        RECT 85.950 524.100 87.150 525.900 ;
        RECT 89.100 525.150 90.900 525.900 ;
        RECT 104.100 525.150 105.900 525.900 ;
        RECT 107.850 524.100 109.050 525.900 ;
        RECT 110.100 525.150 111.900 525.900 ;
        RECT 122.100 525.150 123.900 525.900 ;
        RECT 113.100 524.100 114.900 524.850 ;
        RECT 119.100 524.100 120.900 524.850 ;
        RECT 124.950 524.100 126.150 525.900 ;
        RECT 128.100 525.150 129.900 525.900 ;
        RECT 142.950 523.950 148.050 526.050 ;
        RECT 161.400 524.100 162.300 533.400 ;
        RECT 185.850 530.100 187.050 533.400 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 169.950 526.950 172.050 529.050 ;
        RECT 181.950 526.950 184.050 529.050 ;
        RECT 185.850 525.900 186.900 530.100 ;
        RECT 199.950 529.950 202.050 532.050 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 200.100 528.150 201.900 528.900 ;
        RECT 203.400 527.100 204.600 539.400 ;
        RECT 223.500 533.400 225.300 545.400 ;
        RECT 238.500 533.400 240.300 545.400 ;
        RECT 244.800 539.400 246.600 545.400 ;
        RECT 223.950 530.100 225.150 533.400 ;
        RECT 206.100 528.150 207.900 528.900 ;
        RECT 220.950 526.950 223.050 529.050 ;
        RECT 164.100 525.150 165.900 525.900 ;
        RECT 170.100 525.150 171.900 525.900 ;
        RECT 182.100 525.150 183.900 525.900 ;
        RECT 167.100 524.100 168.900 524.850 ;
        RECT 185.850 524.100 187.050 525.900 ;
        RECT 188.100 525.150 189.900 525.900 ;
        RECT 191.100 524.100 192.900 524.850 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 224.100 525.900 225.150 530.100 ;
        RECT 226.950 526.950 229.050 529.050 ;
        RECT 221.100 525.150 222.900 525.900 ;
        RECT 218.100 524.100 219.900 524.850 ;
        RECT 223.950 524.100 225.150 525.900 ;
        RECT 227.100 525.150 228.900 525.900 ;
        RECT 238.800 524.100 240.000 533.400 ;
        RECT 245.400 532.500 246.600 539.400 ;
        RECT 256.500 533.400 258.300 545.400 ;
        RECT 275.700 533.400 277.500 545.400 ;
        RECT 292.800 539.400 294.600 545.400 ;
        RECT 240.900 531.600 246.600 532.500 ;
        RECT 240.900 530.700 242.850 531.600 ;
        RECT 241.950 524.100 242.850 530.700 ;
        RECT 256.950 530.100 258.150 533.400 ;
        RECT 245.100 527.100 246.900 527.850 ;
        RECT 253.950 526.950 256.050 529.050 ;
        RECT 257.100 525.900 258.150 530.100 ;
        RECT 275.850 530.100 277.050 533.400 ;
        RECT 259.950 526.950 262.050 529.050 ;
        RECT 271.950 526.950 274.050 529.050 ;
        RECT 275.850 525.900 276.900 530.100 ;
        RECT 289.950 529.950 292.050 532.050 ;
        RECT 277.950 526.950 280.050 529.050 ;
        RECT 290.100 528.150 291.900 528.900 ;
        RECT 293.400 527.100 294.600 539.400 ;
        RECT 305.400 539.400 307.200 545.400 ;
        RECT 323.400 539.400 325.200 545.400 ;
        RECT 295.950 529.950 298.050 532.200 ;
        RECT 301.950 529.950 304.050 532.050 ;
        RECT 296.100 528.150 297.900 528.900 ;
        RECT 302.100 528.150 303.900 528.900 ;
        RECT 305.400 527.100 306.600 539.400 ;
        RECT 307.950 529.950 310.050 532.050 ;
        RECT 319.950 529.950 322.050 532.050 ;
        RECT 308.100 528.150 309.900 528.900 ;
        RECT 320.100 528.150 321.900 528.900 ;
        RECT 323.400 527.100 324.600 539.400 ;
        RECT 344.700 533.400 346.500 545.400 ;
        RECT 364.800 539.400 366.600 545.400 ;
        RECT 325.950 529.950 328.050 532.050 ;
        RECT 344.850 530.100 346.050 533.400 ;
        RECT 326.100 528.150 327.900 528.900 ;
        RECT 340.950 526.950 343.050 529.050 ;
        RECT 254.100 525.150 255.900 525.900 ;
        RECT 251.100 524.100 252.900 524.850 ;
        RECT 256.950 524.100 258.150 525.900 ;
        RECT 260.100 525.150 261.900 525.900 ;
        RECT 272.100 525.150 273.900 525.900 ;
        RECT 275.850 524.100 277.050 525.900 ;
        RECT 278.100 525.150 279.900 525.900 ;
        RECT 281.100 524.100 282.900 524.850 ;
        RECT 52.950 520.950 55.050 523.050 ;
        RECT 65.550 522.900 70.050 523.050 ;
        RECT 64.950 520.950 70.050 522.900 ;
        RECT 73.950 520.950 76.050 523.050 ;
        RECT 79.950 520.950 82.050 523.050 ;
        RECT 85.950 520.950 88.050 523.050 ;
        RECT 100.950 522.450 105.000 523.050 ;
        RECT 106.950 522.450 109.050 523.050 ;
        RECT 100.950 521.550 109.050 522.450 ;
        RECT 100.950 520.950 105.000 521.550 ;
        RECT 106.950 520.950 109.050 521.550 ;
        RECT 112.950 520.950 115.050 523.050 ;
        RECT 118.950 520.950 121.050 523.050 ;
        RECT 124.950 520.950 127.050 523.050 ;
        RECT 64.950 520.800 67.050 520.950 ;
        RECT 67.950 519.750 69.150 519.900 ;
        RECT 65.400 518.700 69.150 519.750 ;
        RECT 86.850 519.750 88.050 519.900 ;
        RECT 106.950 519.750 108.150 519.900 ;
        RECT 86.850 518.700 90.600 519.750 ;
        RECT 65.400 516.600 66.600 518.700 ;
        RECT 49.800 510.600 51.600 513.600 ;
        RECT 64.800 510.600 66.600 516.600 ;
        RECT 67.800 515.700 75.600 517.050 ;
        RECT 67.800 510.600 69.600 515.700 ;
        RECT 73.800 510.600 75.600 515.700 ;
        RECT 80.400 515.700 88.200 517.050 ;
        RECT 80.400 510.600 82.200 515.700 ;
        RECT 86.400 510.600 88.200 515.700 ;
        RECT 89.400 516.600 90.600 518.700 ;
        RECT 104.400 518.700 108.150 519.750 ;
        RECT 125.850 519.750 127.050 519.900 ;
        RECT 125.850 518.700 129.600 519.750 ;
        RECT 146.400 518.700 147.600 522.900 ;
        RECT 157.950 520.950 163.050 523.050 ;
        RECT 166.950 520.950 169.050 523.050 ;
        RECT 172.950 522.450 175.050 523.050 ;
        RECT 184.950 522.450 187.050 523.050 ;
        RECT 172.950 521.550 187.050 522.450 ;
        RECT 172.950 520.950 175.050 521.550 ;
        RECT 184.950 520.950 187.050 521.550 ;
        RECT 190.950 520.800 193.050 523.050 ;
        RECT 104.400 516.600 105.600 518.700 ;
        RECT 89.400 510.600 91.200 516.600 ;
        RECT 103.800 510.600 105.600 516.600 ;
        RECT 106.800 515.700 114.600 517.050 ;
        RECT 106.800 510.600 108.600 515.700 ;
        RECT 112.800 510.600 114.600 515.700 ;
        RECT 119.400 515.700 127.200 517.050 ;
        RECT 119.400 510.600 121.200 515.700 ;
        RECT 125.400 510.600 127.200 515.700 ;
        RECT 128.400 516.600 129.600 518.700 ;
        RECT 144.000 517.800 147.600 518.700 ;
        RECT 128.400 510.600 130.200 516.600 ;
        RECT 144.000 510.600 145.800 517.800 ;
        RECT 161.400 516.600 162.300 519.900 ;
        RECT 184.950 519.750 186.150 519.900 ;
        RECT 182.400 518.700 186.150 519.750 ;
        RECT 203.400 518.700 204.600 522.900 ;
        RECT 217.950 520.950 220.050 523.050 ;
        RECT 223.950 520.950 226.050 523.050 ;
        RECT 229.950 522.450 232.050 523.050 ;
        RECT 238.950 522.450 241.050 523.050 ;
        RECT 229.950 521.550 241.050 522.450 ;
        RECT 229.950 520.950 232.050 521.550 ;
        RECT 238.950 520.950 241.050 521.550 ;
        RECT 242.100 519.900 242.850 524.100 ;
        RECT 292.950 523.950 298.050 526.050 ;
        RECT 304.950 523.950 310.050 526.050 ;
        RECT 322.950 523.950 328.050 526.050 ;
        RECT 344.850 525.900 345.900 530.100 ;
        RECT 346.950 526.950 349.050 529.050 ;
        RECT 362.100 528.150 363.900 528.900 ;
        RECT 365.400 527.100 366.600 539.400 ;
        RECT 382.500 533.400 384.300 545.400 ;
        RECT 393.150 533.400 394.950 545.400 ;
        RECT 401.550 539.400 403.350 545.400 ;
        RECT 401.550 538.500 402.750 539.400 ;
        RECT 409.350 538.500 411.150 545.400 ;
        RECT 417.150 539.400 418.950 545.400 ;
        RECT 397.950 536.400 402.750 538.500 ;
        RECT 405.450 537.450 412.050 538.500 ;
        RECT 405.450 536.700 407.250 537.450 ;
        RECT 410.250 536.700 412.050 537.450 ;
        RECT 417.150 537.300 421.050 539.400 ;
        RECT 401.550 535.500 402.750 536.400 ;
        RECT 414.450 535.800 416.250 536.400 ;
        RECT 401.550 534.300 409.050 535.500 ;
        RECT 407.250 533.700 409.050 534.300 ;
        RECT 409.950 534.900 416.250 535.800 ;
        RECT 367.950 529.950 370.050 532.050 ;
        RECT 382.950 530.100 384.150 533.400 ;
        RECT 368.100 528.150 369.900 528.900 ;
        RECT 379.950 526.950 382.050 529.050 ;
        RECT 341.100 525.150 342.900 525.900 ;
        RECT 344.850 524.100 346.050 525.900 ;
        RECT 347.100 525.150 348.900 525.900 ;
        RECT 364.950 525.450 367.050 526.050 ;
        RECT 369.000 525.450 373.050 526.050 ;
        RECT 383.100 525.900 384.150 530.100 ;
        RECT 393.150 532.500 394.050 533.400 ;
        RECT 409.950 532.800 410.850 534.900 ;
        RECT 414.450 534.600 416.250 534.900 ;
        RECT 417.150 534.600 419.850 536.400 ;
        RECT 417.150 533.700 418.050 534.600 ;
        RECT 402.450 532.500 410.850 532.800 ;
        RECT 393.150 531.900 410.850 532.500 ;
        RECT 412.050 532.800 418.050 533.700 ;
        RECT 418.950 532.800 421.050 533.700 ;
        RECT 424.650 533.400 426.450 545.400 ;
        RECT 393.150 531.300 404.250 531.900 ;
        RECT 385.950 526.950 388.050 529.050 ;
        RECT 350.100 524.100 351.900 524.850 ;
        RECT 364.950 524.550 373.050 525.450 ;
        RECT 380.100 525.150 381.900 525.900 ;
        RECT 364.950 523.950 367.050 524.550 ;
        RECT 369.000 523.950 373.050 524.550 ;
        RECT 377.100 524.100 378.900 524.850 ;
        RECT 382.950 524.100 384.150 525.900 ;
        RECT 386.100 525.150 387.900 525.900 ;
        RECT 250.950 520.950 253.050 523.050 ;
        RECT 256.950 520.950 259.050 523.050 ;
        RECT 265.950 522.450 268.050 523.050 ;
        RECT 274.950 522.450 277.050 523.050 ;
        RECT 265.950 521.550 277.050 522.450 ;
        RECT 265.950 520.950 268.050 521.550 ;
        RECT 274.950 520.950 277.050 521.550 ;
        RECT 280.950 520.950 283.050 523.050 ;
        RECT 224.850 519.750 226.050 519.900 ;
        RECT 224.850 518.700 228.600 519.750 ;
        RECT 182.400 516.600 183.600 518.700 ;
        RECT 203.400 517.800 207.000 518.700 ;
        RECT 161.400 514.950 166.800 516.600 ;
        RECT 165.000 510.600 166.800 514.950 ;
        RECT 181.800 510.600 183.600 516.600 ;
        RECT 184.800 515.700 192.600 517.050 ;
        RECT 184.800 510.600 186.600 515.700 ;
        RECT 190.800 510.600 192.600 515.700 ;
        RECT 205.200 510.600 207.000 517.800 ;
        RECT 218.400 515.700 226.200 517.050 ;
        RECT 218.400 510.600 220.200 515.700 ;
        RECT 224.400 510.600 226.200 515.700 ;
        RECT 227.400 516.600 228.600 518.700 ;
        RECT 238.800 516.600 240.000 519.900 ;
        RECT 241.950 519.300 242.850 519.900 ;
        RECT 240.900 518.400 242.850 519.300 ;
        RECT 257.850 519.750 259.050 519.900 ;
        RECT 274.950 519.750 276.150 519.900 ;
        RECT 257.850 518.700 261.600 519.750 ;
        RECT 240.900 517.500 246.000 518.400 ;
        RECT 227.400 510.600 229.200 516.600 ;
        RECT 238.500 510.600 240.300 516.600 ;
        RECT 244.800 513.600 246.000 517.500 ;
        RECT 251.400 515.700 259.200 517.050 ;
        RECT 244.800 510.600 246.600 513.600 ;
        RECT 251.400 510.600 253.200 515.700 ;
        RECT 257.400 510.600 259.200 515.700 ;
        RECT 260.400 516.600 261.600 518.700 ;
        RECT 272.400 518.700 276.150 519.750 ;
        RECT 293.400 518.700 294.600 522.900 ;
        RECT 272.400 516.600 273.600 518.700 ;
        RECT 291.000 517.800 294.600 518.700 ;
        RECT 305.400 518.700 306.600 522.900 ;
        RECT 323.400 518.700 324.600 522.900 ;
        RECT 343.950 520.950 346.050 523.050 ;
        RECT 349.950 520.950 352.050 523.050 ;
        RECT 343.950 519.750 345.150 519.900 ;
        RECT 341.400 518.700 345.150 519.750 ;
        RECT 365.400 518.700 366.600 522.900 ;
        RECT 373.950 520.950 379.050 523.050 ;
        RECT 382.950 520.950 385.050 523.050 ;
        RECT 383.850 519.750 385.050 519.900 ;
        RECT 383.850 518.700 387.600 519.750 ;
        RECT 305.400 517.800 309.000 518.700 ;
        RECT 323.400 517.800 327.000 518.700 ;
        RECT 260.400 510.600 262.200 516.600 ;
        RECT 271.800 510.600 273.600 516.600 ;
        RECT 274.800 515.700 282.600 517.050 ;
        RECT 274.800 510.600 276.600 515.700 ;
        RECT 280.800 510.600 282.600 515.700 ;
        RECT 291.000 510.600 292.800 517.800 ;
        RECT 307.200 510.600 309.000 517.800 ;
        RECT 325.200 510.600 327.000 517.800 ;
        RECT 341.400 516.600 342.600 518.700 ;
        RECT 363.000 517.800 366.600 518.700 ;
        RECT 340.800 510.600 342.600 516.600 ;
        RECT 343.800 515.700 351.600 517.050 ;
        RECT 343.800 510.600 345.600 515.700 ;
        RECT 349.800 510.600 351.600 515.700 ;
        RECT 363.000 510.600 364.800 517.800 ;
        RECT 377.400 515.700 385.200 517.050 ;
        RECT 377.400 510.600 379.200 515.700 ;
        RECT 383.400 510.600 385.200 515.700 ;
        RECT 386.400 516.600 387.600 518.700 ;
        RECT 393.150 516.600 394.050 531.300 ;
        RECT 402.450 531.000 404.250 531.300 ;
        RECT 398.100 526.200 402.900 527.400 ;
        RECT 398.100 525.600 399.900 526.200 ;
        RECT 403.950 523.950 406.050 529.050 ;
        RECT 412.050 527.100 412.950 532.800 ;
        RECT 418.950 531.600 423.150 532.800 ;
        RECT 422.250 529.800 424.050 531.600 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 395.100 522.150 396.900 523.950 ;
        RECT 425.250 523.050 426.450 533.400 ;
        RECT 437.400 539.400 439.200 545.400 ;
        RECT 434.100 528.150 435.900 528.900 ;
        RECT 437.400 527.100 438.600 539.400 ;
        RECT 455.700 533.400 457.500 545.400 ;
        RECT 465.150 533.400 466.950 545.400 ;
        RECT 473.550 539.400 475.350 545.400 ;
        RECT 473.550 538.500 474.750 539.400 ;
        RECT 481.350 538.500 483.150 545.400 ;
        RECT 489.150 539.400 490.950 545.400 ;
        RECT 469.950 536.400 474.750 538.500 ;
        RECT 477.450 537.450 484.050 538.500 ;
        RECT 477.450 536.700 479.250 537.450 ;
        RECT 482.250 536.700 484.050 537.450 ;
        RECT 489.150 537.300 493.050 539.400 ;
        RECT 473.550 535.500 474.750 536.400 ;
        RECT 486.450 535.800 488.250 536.400 ;
        RECT 473.550 534.300 481.050 535.500 ;
        RECT 479.250 533.700 481.050 534.300 ;
        RECT 481.950 534.900 488.250 535.800 ;
        RECT 439.950 529.950 442.050 532.050 ;
        RECT 455.850 530.100 457.050 533.400 ;
        RECT 465.150 532.500 466.050 533.400 ;
        RECT 481.950 532.800 482.850 534.900 ;
        RECT 486.450 534.600 488.250 534.900 ;
        RECT 489.150 534.600 491.850 536.400 ;
        RECT 489.150 533.700 490.050 534.600 ;
        RECT 474.450 532.500 482.850 532.800 ;
        RECT 465.150 531.900 482.850 532.500 ;
        RECT 484.050 532.800 490.050 533.700 ;
        RECT 490.950 532.800 493.050 533.700 ;
        RECT 496.650 533.400 498.450 545.400 ;
        RECT 465.150 531.300 476.250 531.900 ;
        RECT 440.100 528.150 441.900 528.900 ;
        RECT 451.950 528.450 454.050 529.050 ;
        RECT 446.550 527.550 454.050 528.450 ;
        RECT 436.950 525.450 439.050 526.050 ;
        RECT 446.550 525.450 447.450 527.550 ;
        RECT 451.950 526.950 454.050 527.550 ;
        RECT 455.850 525.900 456.900 530.100 ;
        RECT 457.950 526.950 460.050 529.050 ;
        RECT 436.950 524.550 447.450 525.450 ;
        RECT 452.100 525.150 453.900 525.900 ;
        RECT 436.950 523.950 439.050 524.550 ;
        RECT 455.850 524.100 457.050 525.900 ;
        RECT 458.100 525.150 459.900 525.900 ;
        RECT 461.100 524.100 462.900 524.850 ;
        RECT 396.000 521.400 396.900 522.150 ;
        RECT 412.050 522.000 412.950 522.900 ;
        RECT 401.100 521.400 402.900 522.000 ;
        RECT 412.050 521.400 413.850 522.000 ;
        RECT 396.000 520.200 413.850 521.400 ;
        RECT 420.150 520.950 420.900 522.750 ;
        RECT 421.950 520.950 424.050 523.050 ;
        RECT 425.100 520.950 426.450 523.050 ;
        RECT 401.850 517.200 402.900 520.200 ;
        RECT 386.400 510.600 388.200 516.600 ;
        RECT 393.150 510.600 394.950 516.600 ;
        RECT 397.950 514.500 400.050 516.600 ;
        RECT 401.550 515.400 403.350 517.200 ;
        RECT 404.850 516.450 406.650 517.200 ;
        RECT 425.250 516.600 426.450 520.950 ;
        RECT 437.400 518.700 438.600 522.900 ;
        RECT 454.950 520.950 457.050 523.050 ;
        RECT 460.950 520.950 463.050 523.050 ;
        RECT 454.950 519.750 456.150 519.900 ;
        RECT 452.400 518.700 456.150 519.750 ;
        RECT 437.400 517.800 441.000 518.700 ;
        RECT 404.850 515.400 409.800 516.450 ;
        RECT 418.950 515.700 421.050 516.600 ;
        RECT 399.000 513.600 400.050 514.500 ;
        RECT 408.750 513.600 409.800 515.400 ;
        RECT 417.300 514.500 421.050 515.700 ;
        RECT 417.300 513.600 418.350 514.500 ;
        RECT 399.000 512.700 402.750 513.600 ;
        RECT 400.950 510.600 402.750 512.700 ;
        RECT 408.750 510.600 410.550 513.600 ;
        RECT 416.550 510.600 418.350 513.600 ;
        RECT 424.650 510.600 426.450 516.600 ;
        RECT 439.200 510.600 441.000 517.800 ;
        RECT 452.400 516.600 453.600 518.700 ;
        RECT 451.800 510.600 453.600 516.600 ;
        RECT 454.800 515.700 462.600 517.050 ;
        RECT 454.800 510.600 456.600 515.700 ;
        RECT 460.800 510.600 462.600 515.700 ;
        RECT 465.150 516.600 466.050 531.300 ;
        RECT 474.450 531.000 476.250 531.300 ;
        RECT 470.100 526.200 474.900 527.400 ;
        RECT 470.100 525.600 471.900 526.200 ;
        RECT 475.950 523.950 478.050 529.050 ;
        RECT 484.050 527.100 484.950 532.800 ;
        RECT 490.950 531.600 495.150 532.800 ;
        RECT 494.250 529.800 496.050 531.600 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 467.100 522.150 468.900 523.950 ;
        RECT 497.250 523.050 498.450 533.400 ;
        RECT 468.000 521.400 468.900 522.150 ;
        RECT 484.050 522.000 484.950 522.900 ;
        RECT 473.100 521.400 474.900 522.000 ;
        RECT 484.050 521.400 485.850 522.000 ;
        RECT 468.000 520.200 485.850 521.400 ;
        RECT 492.150 520.950 492.900 522.750 ;
        RECT 493.950 520.950 496.050 523.050 ;
        RECT 497.100 520.950 498.450 523.050 ;
        RECT 473.850 517.200 474.900 520.200 ;
        RECT 465.150 510.600 466.950 516.600 ;
        RECT 469.950 514.500 472.050 516.600 ;
        RECT 473.550 515.400 475.350 517.200 ;
        RECT 476.850 516.450 478.650 517.200 ;
        RECT 497.250 516.600 498.450 520.950 ;
        RECT 476.850 515.400 481.800 516.450 ;
        RECT 490.950 515.700 493.050 516.600 ;
        RECT 471.000 513.600 472.050 514.500 ;
        RECT 480.750 513.600 481.800 515.400 ;
        RECT 489.300 514.500 493.050 515.700 ;
        RECT 489.300 513.600 490.350 514.500 ;
        RECT 471.000 512.700 474.750 513.600 ;
        RECT 472.950 510.600 474.750 512.700 ;
        RECT 480.750 510.600 482.550 513.600 ;
        RECT 488.550 510.600 490.350 513.600 ;
        RECT 496.650 510.600 498.450 516.600 ;
        RECT 501.150 533.400 502.950 545.400 ;
        RECT 509.550 539.400 511.350 545.400 ;
        RECT 509.550 538.500 510.750 539.400 ;
        RECT 517.350 538.500 519.150 545.400 ;
        RECT 525.150 539.400 526.950 545.400 ;
        RECT 505.950 536.400 510.750 538.500 ;
        RECT 513.450 537.450 520.050 538.500 ;
        RECT 513.450 536.700 515.250 537.450 ;
        RECT 518.250 536.700 520.050 537.450 ;
        RECT 525.150 537.300 529.050 539.400 ;
        RECT 509.550 535.500 510.750 536.400 ;
        RECT 522.450 535.800 524.250 536.400 ;
        RECT 509.550 534.300 517.050 535.500 ;
        RECT 515.250 533.700 517.050 534.300 ;
        RECT 517.950 534.900 524.250 535.800 ;
        RECT 501.150 532.500 502.050 533.400 ;
        RECT 517.950 532.800 518.850 534.900 ;
        RECT 522.450 534.600 524.250 534.900 ;
        RECT 525.150 534.600 527.850 536.400 ;
        RECT 525.150 533.700 526.050 534.600 ;
        RECT 510.450 532.500 518.850 532.800 ;
        RECT 501.150 531.900 518.850 532.500 ;
        RECT 520.050 532.800 526.050 533.700 ;
        RECT 526.950 532.800 529.050 533.700 ;
        RECT 532.650 533.400 534.450 545.400 ;
        RECT 547.800 539.400 549.600 545.400 ;
        RECT 501.150 531.300 512.250 531.900 ;
        RECT 501.150 516.600 502.050 531.300 ;
        RECT 510.450 531.000 512.250 531.300 ;
        RECT 506.100 526.200 510.900 527.400 ;
        RECT 506.100 525.600 507.900 526.200 ;
        RECT 511.950 523.950 514.050 529.050 ;
        RECT 520.050 527.100 520.950 532.800 ;
        RECT 526.950 531.600 531.150 532.800 ;
        RECT 530.250 529.800 532.050 531.600 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 503.100 522.150 504.900 523.950 ;
        RECT 533.250 523.050 534.450 533.400 ;
        RECT 545.100 528.150 546.900 528.900 ;
        RECT 548.400 527.100 549.600 539.400 ;
        RECT 560.400 539.400 562.200 545.400 ;
        RECT 550.950 529.950 553.050 532.050 ;
        RECT 551.100 528.150 552.900 528.900 ;
        RECT 557.100 527.100 558.900 527.850 ;
        RECT 538.950 525.450 541.050 526.050 ;
        RECT 547.950 525.450 550.050 526.050 ;
        RECT 538.950 524.550 550.050 525.450 ;
        RECT 538.950 523.950 541.050 524.550 ;
        RECT 547.950 523.950 550.050 524.550 ;
        RECT 556.950 523.950 559.050 526.200 ;
        RECT 504.000 521.400 504.900 522.150 ;
        RECT 520.050 522.000 520.950 522.900 ;
        RECT 509.100 521.400 510.900 522.000 ;
        RECT 520.050 521.400 521.850 522.000 ;
        RECT 504.000 520.200 521.850 521.400 ;
        RECT 528.150 520.950 528.900 522.750 ;
        RECT 529.950 520.950 532.050 523.050 ;
        RECT 533.100 520.950 534.450 523.050 ;
        RECT 509.850 517.200 510.900 520.200 ;
        RECT 501.150 510.600 502.950 516.600 ;
        RECT 505.950 514.500 508.050 516.600 ;
        RECT 509.550 515.400 511.350 517.200 ;
        RECT 512.850 516.450 514.650 517.200 ;
        RECT 533.250 516.600 534.450 520.950 ;
        RECT 548.400 518.700 549.600 522.900 ;
        RECT 560.400 519.300 561.450 539.400 ;
        RECT 567.000 533.400 568.800 545.400 ;
        RECT 578.400 539.400 580.200 545.400 ;
        RECT 578.700 539.100 580.200 539.400 ;
        RECT 584.400 539.400 586.200 545.400 ;
        RECT 596.400 539.400 598.200 545.400 ;
        RECT 611.400 539.400 613.200 545.400 ;
        RECT 584.400 539.100 585.300 539.400 ;
        RECT 578.700 538.200 585.300 539.100 ;
        RECT 563.100 525.150 564.900 525.900 ;
        RECT 567.000 524.100 568.050 533.400 ;
        RECT 574.950 532.950 577.050 535.050 ;
        RECT 584.400 533.100 585.300 538.200 ;
        RECT 575.100 531.150 576.900 531.900 ;
        RECT 578.100 530.100 579.900 530.850 ;
        RECT 583.950 529.950 589.050 532.050 ;
        RECT 592.950 529.950 595.050 532.050 ;
        RECT 577.950 526.950 580.050 529.050 ;
        RECT 580.950 523.950 583.050 526.050 ;
        RECT 565.950 522.450 571.050 523.050 ;
        RECT 574.950 522.450 577.050 523.050 ;
        RECT 565.950 521.550 577.050 522.450 ;
        RECT 581.100 522.150 582.900 522.900 ;
        RECT 565.950 520.950 571.050 521.550 ;
        RECT 574.950 520.950 577.050 521.550 ;
        RECT 584.400 520.650 585.300 528.900 ;
        RECT 593.100 528.150 594.900 528.900 ;
        RECT 596.400 527.100 597.600 539.400 ;
        RECT 598.950 529.950 601.050 532.050 ;
        RECT 607.950 529.950 610.050 532.050 ;
        RECT 599.100 528.150 600.900 528.900 ;
        RECT 608.100 528.150 609.900 528.900 ;
        RECT 611.400 527.100 612.600 539.400 ;
        RECT 631.500 533.400 633.300 545.400 ;
        RECT 650.400 539.400 652.200 545.400 ;
        RECT 631.950 530.100 633.150 533.400 ;
        RECT 614.100 528.150 615.900 528.900 ;
        RECT 628.950 526.950 631.050 529.050 ;
        RECT 589.950 525.450 594.000 526.050 ;
        RECT 595.950 525.450 598.050 526.050 ;
        RECT 589.950 524.550 598.050 525.450 ;
        RECT 589.950 523.950 594.000 524.550 ;
        RECT 595.950 523.950 598.050 524.550 ;
        RECT 610.950 525.450 613.050 526.050 ;
        RECT 619.950 525.450 622.050 526.050 ;
        RECT 632.100 525.900 633.150 530.100 ;
        RECT 634.950 526.950 637.050 529.050 ;
        RECT 647.100 527.100 648.900 527.850 ;
        RECT 610.950 524.550 622.050 525.450 ;
        RECT 629.100 525.150 630.900 525.900 ;
        RECT 610.950 523.950 613.050 524.550 ;
        RECT 619.950 523.950 622.050 524.550 ;
        RECT 626.100 524.100 627.900 524.850 ;
        RECT 631.950 524.100 633.150 525.900 ;
        RECT 635.100 525.150 636.900 525.900 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 512.850 515.400 517.800 516.450 ;
        RECT 526.950 515.700 529.050 516.600 ;
        RECT 507.000 513.600 508.050 514.500 ;
        RECT 516.750 513.600 517.800 515.400 ;
        RECT 525.300 514.500 529.050 515.700 ;
        RECT 525.300 513.600 526.350 514.500 ;
        RECT 507.000 512.700 510.750 513.600 ;
        RECT 508.950 510.600 510.750 512.700 ;
        RECT 516.750 510.600 518.550 513.600 ;
        RECT 524.550 510.600 526.350 513.600 ;
        RECT 532.650 510.600 534.450 516.600 ;
        RECT 546.000 517.800 549.600 518.700 ;
        RECT 557.400 518.400 564.900 519.300 ;
        RECT 546.000 510.600 547.800 517.800 ;
        RECT 557.400 510.600 559.200 518.400 ;
        RECT 563.100 517.500 564.900 518.400 ;
        RECT 565.950 516.600 566.850 519.900 ;
        RECT 564.900 514.800 566.850 516.600 ;
        RECT 581.100 519.000 585.300 520.650 ;
        RECT 564.900 510.600 566.700 514.800 ;
        RECT 581.100 510.600 582.900 519.000 ;
        RECT 596.400 518.700 597.600 522.900 ;
        RECT 611.400 518.700 612.600 522.900 ;
        RECT 625.950 520.950 628.050 523.050 ;
        RECT 631.950 522.450 634.050 523.050 ;
        RECT 636.000 522.450 640.050 523.050 ;
        RECT 631.950 521.550 640.050 522.450 ;
        RECT 631.950 520.950 634.050 521.550 ;
        RECT 636.000 520.950 640.050 521.550 ;
        RECT 632.850 519.750 634.050 519.900 ;
        RECT 632.850 518.700 636.600 519.750 ;
        RECT 650.400 519.300 651.450 539.400 ;
        RECT 657.000 533.400 658.800 545.400 ;
        RECT 673.800 539.400 675.600 545.400 ;
        RECT 652.950 526.950 655.050 529.050 ;
        RECT 653.100 525.150 654.900 525.900 ;
        RECT 657.000 524.100 658.050 533.400 ;
        RECT 670.950 529.950 673.050 532.050 ;
        RECT 671.100 528.150 672.900 528.900 ;
        RECT 674.400 527.100 675.600 539.400 ;
        RECT 683.400 533.400 685.200 545.400 ;
        RECT 690.900 534.900 692.700 545.400 ;
        RECT 690.900 533.400 693.300 534.900 ;
        RECT 706.800 533.400 708.600 545.400 ;
        RECT 709.800 534.300 711.600 545.400 ;
        RECT 715.800 534.300 717.600 545.400 ;
        RECT 709.800 533.400 717.600 534.300 ;
        RECT 726.600 533.400 728.400 545.400 ;
        RECT 742.500 533.400 744.300 545.400 ;
        RECT 758.400 534.300 760.200 545.400 ;
        RECT 764.400 534.300 766.200 545.400 ;
        RECT 758.400 533.400 766.200 534.300 ;
        RECT 767.400 533.400 769.200 545.400 ;
        RECT 779.400 539.400 781.200 545.400 ;
        RECT 796.800 539.400 798.600 545.400 ;
        RECT 683.400 532.200 684.600 533.400 ;
        RECT 676.950 529.950 679.050 532.050 ;
        RECT 683.400 531.000 690.600 532.200 ;
        RECT 688.800 530.400 690.600 531.000 ;
        RECT 677.100 528.150 678.900 528.900 ;
        RECT 682.950 526.950 685.050 529.050 ;
        RECT 664.950 525.450 667.050 526.050 ;
        RECT 673.950 525.450 676.050 526.050 ;
        RECT 664.950 524.550 676.050 525.450 ;
        RECT 683.100 525.150 684.900 525.900 ;
        RECT 664.950 523.950 667.050 524.550 ;
        RECT 673.950 523.950 676.050 524.550 ;
        RECT 686.100 524.100 687.900 524.850 ;
        RECT 655.950 520.950 661.050 523.050 ;
        RECT 596.400 517.800 600.000 518.700 ;
        RECT 611.400 517.800 615.000 518.700 ;
        RECT 598.200 510.600 600.000 517.800 ;
        RECT 613.200 510.600 615.000 517.800 ;
        RECT 626.400 515.700 634.200 517.050 ;
        RECT 626.400 510.600 628.200 515.700 ;
        RECT 632.400 510.600 634.200 515.700 ;
        RECT 635.400 516.600 636.600 518.700 ;
        RECT 647.400 518.400 654.900 519.300 ;
        RECT 635.400 510.600 637.200 516.600 ;
        RECT 647.400 510.600 649.200 518.400 ;
        RECT 653.100 517.500 654.900 518.400 ;
        RECT 655.950 516.600 656.850 519.900 ;
        RECT 674.400 518.700 675.600 522.900 ;
        RECT 685.950 520.950 688.050 523.050 ;
        RECT 689.700 519.600 690.600 530.400 ;
        RECT 691.950 527.100 693.300 533.400 ;
        RECT 697.950 526.050 700.050 526.200 ;
        RECT 691.950 525.450 694.050 526.050 ;
        RECT 696.000 525.450 700.050 526.050 ;
        RECT 691.950 524.550 700.050 525.450 ;
        RECT 691.950 523.950 694.050 524.550 ;
        RECT 696.000 524.100 700.050 524.550 ;
        RECT 707.400 524.100 708.300 533.400 ;
        RECT 726.600 532.350 729.300 533.400 ;
        RECT 709.950 526.950 712.050 529.050 ;
        RECT 715.950 526.950 718.050 529.200 ;
        RECT 725.100 527.100 726.900 527.850 ;
        RECT 727.950 527.100 729.300 532.350 ;
        RECT 731.100 530.100 732.900 530.850 ;
        RECT 742.950 530.100 744.150 533.400 ;
        RECT 710.100 525.150 711.900 525.900 ;
        RECT 716.100 525.150 717.900 525.900 ;
        RECT 713.100 524.100 714.900 524.850 ;
        RECT 696.000 523.950 699.000 524.100 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 688.950 518.700 690.750 519.600 ;
        RECT 654.900 514.800 656.850 516.600 ;
        RECT 672.000 517.800 675.600 518.700 ;
        RECT 687.300 517.800 690.750 518.700 ;
        RECT 654.900 510.600 656.700 514.800 ;
        RECT 672.000 510.600 673.800 517.800 ;
        RECT 687.300 513.600 688.200 517.800 ;
        RECT 693.000 516.600 694.050 522.900 ;
        RECT 697.950 522.450 700.050 522.900 ;
        RECT 706.950 522.450 709.050 523.050 ;
        RECT 697.950 521.550 709.050 522.450 ;
        RECT 697.950 520.800 700.050 521.550 ;
        RECT 706.950 520.950 709.050 521.550 ;
        RECT 712.950 520.950 715.050 523.050 ;
        RECT 728.100 522.900 729.300 527.100 ;
        RECT 730.950 526.950 733.050 529.050 ;
        RECT 739.950 526.950 742.050 529.050 ;
        RECT 743.100 525.900 744.150 530.100 ;
        RECT 745.950 526.950 748.050 529.050 ;
        RECT 757.950 526.950 760.050 529.050 ;
        RECT 763.950 526.950 766.050 529.050 ;
        RECT 740.100 525.150 741.900 525.900 ;
        RECT 737.100 524.100 738.900 524.850 ;
        RECT 742.950 524.100 744.150 525.900 ;
        RECT 746.100 525.150 747.900 525.900 ;
        RECT 758.100 525.150 759.900 525.900 ;
        RECT 764.100 525.150 765.900 525.900 ;
        RECT 761.100 524.100 762.900 524.850 ;
        RECT 767.700 524.100 768.600 533.400 ;
        RECT 775.950 529.950 778.050 532.050 ;
        RECT 776.100 528.150 777.900 528.900 ;
        RECT 779.400 527.100 780.600 539.400 ;
        RECT 797.700 539.100 798.600 539.400 ;
        RECT 802.800 539.400 804.600 545.400 ;
        RECT 815.400 539.400 817.200 545.400 ;
        RECT 802.800 539.100 804.300 539.400 ;
        RECT 797.700 538.200 804.300 539.100 ;
        RECT 797.700 533.100 798.600 538.200 ;
        RECT 805.950 532.950 808.050 535.050 ;
        RECT 815.400 532.500 816.600 539.400 ;
        RECT 821.700 533.400 823.500 545.400 ;
        RECT 781.950 529.950 784.050 532.050 ;
        RECT 790.950 531.450 795.000 532.050 ;
        RECT 796.950 531.450 799.050 532.050 ;
        RECT 790.950 530.550 799.050 531.450 ;
        RECT 806.100 531.150 807.900 531.900 ;
        RECT 815.400 531.600 821.100 532.500 ;
        RECT 790.950 529.950 795.000 530.550 ;
        RECT 796.950 529.950 799.050 530.550 ;
        RECT 803.100 530.100 804.900 530.850 ;
        RECT 819.150 530.700 821.100 531.600 ;
        RECT 782.100 528.150 783.900 528.900 ;
        RECT 772.950 525.450 777.000 526.050 ;
        RECT 778.950 525.450 781.050 526.050 ;
        RECT 772.950 524.550 781.050 525.450 ;
        RECT 772.950 523.950 777.000 524.550 ;
        RECT 778.950 523.950 781.050 524.550 ;
        RECT 727.950 521.100 729.300 522.900 ;
        RECT 736.950 520.950 739.050 523.050 ;
        RECT 742.950 520.950 745.050 523.050 ;
        RECT 751.950 522.450 754.050 523.050 ;
        RECT 760.950 522.450 763.050 523.050 ;
        RECT 751.950 521.550 763.050 522.450 ;
        RECT 751.950 520.950 754.050 521.550 ;
        RECT 760.950 520.950 763.050 521.550 ;
        RECT 766.950 520.950 769.050 523.050 ;
        RECT 707.400 516.600 708.300 519.900 ;
        RECT 718.950 519.450 721.050 520.050 ;
        RECT 727.950 519.450 730.050 520.050 ;
        RECT 718.950 518.550 730.050 519.450 ;
        RECT 743.850 519.750 745.050 519.900 ;
        RECT 743.850 518.700 747.600 519.750 ;
        RECT 718.950 517.950 721.050 518.550 ;
        RECT 727.950 517.950 730.050 518.550 ;
        RECT 686.400 510.600 688.200 513.600 ;
        RECT 692.400 510.600 694.200 516.600 ;
        RECT 707.400 514.950 712.800 516.600 ;
        RECT 711.000 510.600 712.800 514.950 ;
        RECT 728.400 513.600 729.600 516.900 ;
        RECT 727.800 510.600 729.600 513.600 ;
        RECT 737.400 515.700 745.200 517.050 ;
        RECT 737.400 510.600 739.200 515.700 ;
        RECT 743.400 510.600 745.200 515.700 ;
        RECT 746.400 516.600 747.600 518.700 ;
        RECT 767.700 516.600 768.600 519.900 ;
        RECT 779.400 518.700 780.600 522.900 ;
        RECT 797.700 520.650 798.600 528.900 ;
        RECT 802.950 526.950 805.050 529.050 ;
        RECT 815.100 527.100 816.900 527.850 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 800.100 522.150 801.900 522.900 ;
        RECT 814.950 520.950 817.050 526.050 ;
        RECT 819.150 524.100 820.050 530.700 ;
        RECT 822.000 524.100 823.200 533.400 ;
        RECT 797.700 519.000 801.900 520.650 ;
        RECT 779.400 517.800 783.000 518.700 ;
        RECT 746.400 510.600 748.200 516.600 ;
        RECT 763.200 514.950 768.600 516.600 ;
        RECT 763.200 510.600 765.000 514.950 ;
        RECT 781.200 510.600 783.000 517.800 ;
        RECT 800.100 510.600 801.900 519.000 ;
        RECT 819.150 519.900 819.900 524.100 ;
        RECT 819.150 519.300 820.050 519.900 ;
        RECT 819.150 518.400 821.100 519.300 ;
        RECT 816.000 517.500 821.100 518.400 ;
        RECT 816.000 513.600 817.200 517.500 ;
        RECT 822.000 516.600 823.200 519.900 ;
        RECT 815.400 510.600 817.200 513.600 ;
        RECT 821.700 510.600 823.500 516.600 ;
        RECT 5.400 501.300 7.200 506.400 ;
        RECT 11.400 501.300 13.200 506.400 ;
        RECT 5.400 499.950 13.200 501.300 ;
        RECT 14.400 500.400 16.200 506.400 ;
        RECT 28.800 503.400 30.600 506.400 ;
        RECT 14.400 498.300 15.600 500.400 ;
        RECT 11.850 497.250 15.600 498.300 ;
        RECT 11.850 497.100 13.050 497.250 ;
        RECT 4.950 493.950 7.050 496.050 ;
        RECT 10.950 495.450 13.050 496.050 ;
        RECT 22.950 495.450 25.050 496.050 ;
        RECT 10.950 494.550 25.050 495.450 ;
        RECT 10.950 493.950 13.050 494.550 ;
        RECT 22.950 493.950 25.050 494.550 ;
        RECT 5.100 492.150 6.900 492.900 ;
        RECT 8.100 491.100 9.900 491.850 ;
        RECT 10.950 491.100 12.150 492.900 ;
        RECT 14.100 491.100 15.900 491.850 ;
        RECT 7.950 487.950 10.050 490.200 ;
        RECT 11.100 486.900 12.150 491.100 ;
        RECT 13.950 487.950 16.050 490.050 ;
        RECT 19.950 489.450 22.050 493.050 ;
        RECT 29.400 491.100 30.600 503.400 ;
        RECT 44.100 498.000 45.900 506.400 ;
        RECT 61.800 503.400 63.600 506.400 ;
        RECT 44.100 496.350 48.300 498.000 ;
        RECT 31.950 493.950 34.050 496.050 ;
        RECT 44.100 494.100 45.900 494.850 ;
        RECT 32.100 492.150 33.900 492.900 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 28.950 489.450 31.050 490.050 ;
        RECT 19.950 489.000 31.050 489.450 ;
        RECT 20.550 488.550 31.050 489.000 ;
        RECT 28.950 487.950 31.050 488.550 ;
        RECT 40.950 487.950 43.050 490.050 ;
        RECT 47.400 488.100 48.300 496.350 ;
        RECT 62.400 491.100 63.600 503.400 ;
        RECT 78.000 502.050 79.800 506.400 ;
        RECT 74.400 500.400 79.800 502.050 ;
        RECT 74.400 497.100 75.300 500.400 ;
        RECT 98.100 498.000 99.900 506.400 ;
        RECT 120.000 502.050 121.800 506.400 ;
        RECT 95.700 496.350 99.900 498.000 ;
        RECT 116.400 500.400 121.800 502.050 ;
        RECT 134.400 503.400 136.200 506.400 ;
        RECT 149.400 503.400 151.200 506.400 ;
        RECT 166.800 503.400 168.600 506.400 ;
        RECT 116.400 497.100 117.300 500.400 ;
        RECT 64.950 493.950 67.050 496.050 ;
        RECT 70.950 493.950 76.050 496.050 ;
        RECT 79.950 493.950 82.050 496.050 ;
        RECT 65.100 492.150 66.900 492.900 ;
        RECT 52.950 489.450 55.050 490.050 ;
        RECT 61.950 489.450 64.050 490.050 ;
        RECT 52.950 488.550 64.050 489.450 ;
        RECT 52.950 487.950 55.050 488.550 ;
        RECT 61.950 487.950 64.050 488.550 ;
        RECT 10.950 483.600 12.150 486.900 ;
        RECT 10.500 471.600 12.300 483.600 ;
        RECT 29.400 477.600 30.600 486.900 ;
        RECT 41.100 486.150 42.900 486.900 ;
        RECT 38.100 485.100 39.900 485.850 ;
        RECT 46.950 484.950 49.050 487.050 ;
        RECT 31.950 483.450 36.000 484.050 ;
        RECT 37.950 483.450 40.050 484.050 ;
        RECT 31.950 482.550 40.050 483.450 ;
        RECT 31.950 481.950 36.000 482.550 ;
        RECT 37.950 481.950 40.050 482.550 ;
        RECT 47.400 478.800 48.300 483.900 ;
        RECT 41.700 477.900 48.300 478.800 ;
        RECT 41.700 477.600 43.200 477.900 ;
        RECT 28.800 471.600 30.600 477.600 ;
        RECT 41.400 471.600 43.200 477.600 ;
        RECT 47.400 477.600 48.300 477.900 ;
        RECT 62.400 477.600 63.600 486.900 ;
        RECT 74.400 483.600 75.300 492.900 ;
        RECT 80.100 492.150 81.900 492.900 ;
        RECT 77.100 491.100 78.900 491.850 ;
        RECT 83.100 491.100 84.900 491.850 ;
        RECT 76.950 487.950 79.050 490.050 ;
        RECT 82.950 487.950 85.050 490.050 ;
        RECT 95.700 488.100 96.600 496.350 ;
        RECT 98.100 494.100 99.900 494.850 ;
        RECT 115.950 493.950 118.050 496.050 ;
        RECT 121.950 493.950 124.050 496.050 ;
        RECT 130.950 493.950 133.050 496.050 ;
        RECT 97.950 490.950 100.050 493.050 ;
        RECT 100.950 487.950 103.050 490.050 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 101.100 486.150 102.900 486.900 ;
        RECT 104.100 485.100 105.900 485.850 ;
        RECT 47.400 471.600 49.200 477.600 ;
        RECT 61.800 471.600 63.600 477.600 ;
        RECT 73.800 471.600 75.600 483.600 ;
        RECT 76.800 482.700 84.600 483.600 ;
        RECT 76.800 471.600 78.600 482.700 ;
        RECT 82.800 471.600 84.600 482.700 ;
        RECT 95.700 478.800 96.600 483.900 ;
        RECT 103.950 481.950 106.050 484.050 ;
        RECT 116.400 483.600 117.300 492.900 ;
        RECT 122.100 492.150 123.900 492.900 ;
        RECT 131.100 492.150 132.900 492.900 ;
        RECT 119.100 491.100 120.900 491.850 ;
        RECT 125.100 491.100 126.900 491.850 ;
        RECT 134.400 491.100 135.600 503.400 ;
        RECT 145.950 493.950 148.050 496.050 ;
        RECT 146.100 492.150 147.900 492.900 ;
        RECT 149.400 491.100 150.600 503.400 ;
        RECT 167.400 500.100 168.600 503.400 ;
        RECT 184.200 499.200 186.000 506.400 ;
        RECT 151.950 498.450 154.050 499.050 ;
        RECT 166.950 498.450 169.050 499.050 ;
        RECT 151.950 497.550 169.050 498.450 ;
        RECT 151.950 496.950 154.050 497.550 ;
        RECT 166.950 496.950 169.050 497.550 ;
        RECT 182.400 498.300 186.000 499.200 ;
        RECT 166.950 494.100 168.300 495.900 ;
        RECT 163.950 490.950 166.050 493.050 ;
        RECT 118.950 487.950 121.050 490.050 ;
        RECT 124.950 487.950 127.050 490.050 ;
        RECT 131.550 489.900 136.050 490.050 ;
        RECT 130.950 487.950 136.050 489.900 ;
        RECT 139.950 489.450 142.050 489.900 ;
        RECT 148.950 489.450 151.050 490.050 ;
        RECT 167.100 489.900 168.300 494.100 ;
        RECT 175.950 492.450 178.050 496.050 ;
        RECT 182.400 494.100 183.600 498.300 ;
        RECT 203.100 498.000 204.900 506.400 ;
        RECT 223.200 499.200 225.000 506.400 ;
        RECT 237.300 502.200 239.100 506.400 ;
        RECT 200.700 496.350 204.900 498.000 ;
        RECT 221.400 498.300 225.000 499.200 ;
        RECT 237.150 500.400 239.100 502.200 ;
        RECT 181.950 492.450 184.050 493.050 ;
        RECT 175.950 492.000 184.050 492.450 ;
        RECT 176.550 491.550 184.050 492.000 ;
        RECT 181.950 490.950 184.050 491.550 ;
        RECT 139.950 488.550 151.050 489.450 ;
        RECT 164.100 489.150 165.900 489.900 ;
        RECT 130.950 487.800 133.050 487.950 ;
        RECT 139.950 487.800 142.050 488.550 ;
        RECT 148.950 487.950 151.050 488.550 ;
        RECT 95.700 477.900 102.300 478.800 ;
        RECT 95.700 477.600 96.600 477.900 ;
        RECT 94.800 471.600 96.600 477.600 ;
        RECT 100.800 477.600 102.300 477.900 ;
        RECT 100.800 471.600 102.600 477.600 ;
        RECT 115.800 471.600 117.600 483.600 ;
        RECT 118.800 482.700 126.600 483.600 ;
        RECT 118.800 471.600 120.600 482.700 ;
        RECT 124.800 471.600 126.600 482.700 ;
        RECT 134.400 477.600 135.600 486.900 ;
        RECT 149.400 477.600 150.600 486.900 ;
        RECT 166.950 484.650 168.300 489.900 ;
        RECT 169.950 487.950 172.050 490.050 ;
        RECT 179.100 488.100 180.900 488.850 ;
        RECT 170.100 486.150 171.900 486.900 ;
        RECT 178.950 484.950 181.050 487.050 ;
        RECT 165.600 483.600 168.300 484.650 ;
        RECT 134.400 471.600 136.200 477.600 ;
        RECT 149.400 471.600 151.200 477.600 ;
        RECT 165.600 471.600 167.400 483.600 ;
        RECT 182.400 477.600 183.600 489.900 ;
        RECT 185.100 488.100 186.900 488.850 ;
        RECT 200.700 488.100 201.600 496.350 ;
        RECT 203.100 494.100 204.900 494.850 ;
        RECT 221.400 494.100 222.600 498.300 ;
        RECT 237.150 497.100 238.050 500.400 ;
        RECT 239.100 498.600 240.900 499.500 ;
        RECT 244.800 498.600 246.600 506.400 ;
        RECT 239.100 497.700 246.600 498.600 ;
        RECT 257.400 503.400 259.200 506.400 ;
        RECT 268.800 503.400 270.600 506.400 ;
        RECT 232.950 493.950 238.050 496.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 217.950 492.450 223.050 493.050 ;
        RECT 225.000 492.450 229.050 493.050 ;
        RECT 217.950 491.550 229.050 492.450 ;
        RECT 217.950 490.950 223.050 491.550 ;
        RECT 225.000 490.950 229.050 491.550 ;
        RECT 205.950 487.950 208.050 490.050 ;
        RECT 218.100 488.100 219.900 488.850 ;
        RECT 184.950 484.950 187.050 487.050 ;
        RECT 190.950 486.450 193.050 487.050 ;
        RECT 199.950 486.450 202.050 487.050 ;
        RECT 190.950 485.550 202.050 486.450 ;
        RECT 206.100 486.150 207.900 486.900 ;
        RECT 190.950 484.950 193.050 485.550 ;
        RECT 199.950 484.950 202.050 485.550 ;
        RECT 209.100 485.100 210.900 485.850 ;
        RECT 217.950 484.950 220.050 487.050 ;
        RECT 200.700 478.800 201.600 483.900 ;
        RECT 208.950 481.950 211.050 484.050 ;
        RECT 200.700 477.900 207.300 478.800 ;
        RECT 200.700 477.600 201.600 477.900 ;
        RECT 182.400 471.600 184.200 477.600 ;
        RECT 199.800 471.600 201.600 477.600 ;
        RECT 205.800 477.600 207.300 477.900 ;
        RECT 221.400 477.600 222.600 489.900 ;
        RECT 224.100 488.100 225.900 488.850 ;
        RECT 235.950 483.600 237.000 492.900 ;
        RECT 239.100 491.100 240.900 491.850 ;
        RECT 238.950 487.950 241.050 490.050 ;
        RECT 205.800 471.600 207.600 477.600 ;
        RECT 221.400 471.600 223.200 477.600 ;
        RECT 235.200 471.600 237.000 483.600 ;
        RECT 242.550 477.600 243.600 497.700 ;
        RECT 253.950 493.950 256.050 496.050 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 254.100 492.150 255.900 492.900 ;
        RECT 257.400 491.100 258.600 503.400 ;
        RECT 269.400 491.100 270.600 503.400 ;
        RECT 284.100 498.000 285.900 506.400 ;
        RECT 304.200 499.200 306.000 506.400 ;
        RECT 314.400 501.300 316.200 506.400 ;
        RECT 320.400 501.300 322.200 506.400 ;
        RECT 314.400 499.950 322.200 501.300 ;
        RECT 323.400 500.400 325.200 506.400 ;
        RECT 281.700 496.350 285.900 498.000 ;
        RECT 302.400 498.300 306.000 499.200 ;
        RECT 323.400 498.300 324.600 500.400 ;
        RECT 337.200 499.200 339.000 506.400 ;
        RECT 271.950 493.950 274.050 496.050 ;
        RECT 272.100 492.150 273.900 492.900 ;
        RECT 245.100 489.150 246.900 489.900 ;
        RECT 250.950 489.450 255.000 490.050 ;
        RECT 256.950 489.450 259.050 490.050 ;
        RECT 250.950 488.550 259.050 489.450 ;
        RECT 250.950 487.950 255.000 488.550 ;
        RECT 256.950 487.950 259.050 488.550 ;
        RECT 268.950 487.950 271.050 490.050 ;
        RECT 281.700 488.100 282.600 496.350 ;
        RECT 284.100 494.100 285.900 494.850 ;
        RECT 302.400 494.100 303.600 498.300 ;
        RECT 320.850 497.250 324.600 498.300 ;
        RECT 335.400 498.300 339.000 499.200 ;
        RECT 344.550 500.400 346.350 506.400 ;
        RECT 352.650 503.400 354.450 506.400 ;
        RECT 360.450 503.400 362.250 506.400 ;
        RECT 368.250 504.300 370.050 506.400 ;
        RECT 368.250 503.400 372.000 504.300 ;
        RECT 352.650 502.500 353.700 503.400 ;
        RECT 349.950 501.300 353.700 502.500 ;
        RECT 361.200 501.600 362.250 503.400 ;
        RECT 370.950 502.500 372.000 503.400 ;
        RECT 349.950 500.400 352.050 501.300 ;
        RECT 361.200 500.550 366.150 501.600 ;
        RECT 320.850 497.100 322.050 497.250 ;
        RECT 313.950 493.950 316.050 496.050 ;
        RECT 319.950 495.450 322.050 496.050 ;
        RECT 328.950 495.450 331.050 496.050 ;
        RECT 319.950 494.550 331.050 495.450 ;
        RECT 319.950 493.950 322.050 494.550 ;
        RECT 328.950 493.950 331.050 494.550 ;
        RECT 335.400 494.100 336.600 498.300 ;
        RECT 344.550 496.050 345.750 500.400 ;
        RECT 364.350 499.800 366.150 500.550 ;
        RECT 367.650 499.800 369.450 501.600 ;
        RECT 370.950 500.400 373.050 502.500 ;
        RECT 376.050 500.400 377.850 506.400 ;
        RECT 368.100 496.800 369.150 499.800 ;
        RECT 344.550 493.950 345.900 496.050 ;
        RECT 346.950 493.950 349.050 496.050 ;
        RECT 350.100 494.250 350.850 496.050 ;
        RECT 357.150 495.600 375.000 496.800 ;
        RECT 357.150 495.000 358.950 495.600 ;
        RECT 368.100 495.000 369.900 495.600 ;
        RECT 358.050 494.100 358.950 495.000 ;
        RECT 374.100 494.850 375.000 495.600 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 301.950 490.950 307.050 493.050 ;
        RECT 314.100 492.150 315.900 492.900 ;
        RECT 317.100 491.100 318.900 491.850 ;
        RECT 319.950 491.100 321.150 492.900 ;
        RECT 323.100 491.100 324.900 491.850 ;
        RECT 286.950 487.950 289.050 490.050 ;
        RECT 299.100 488.100 300.900 488.850 ;
        RECT 241.800 471.600 243.600 477.600 ;
        RECT 257.400 477.600 258.600 486.900 ;
        RECT 269.400 477.600 270.600 486.900 ;
        RECT 280.950 484.950 283.050 487.050 ;
        RECT 287.100 486.150 288.900 486.900 ;
        RECT 290.100 485.100 291.900 485.850 ;
        RECT 298.950 484.950 301.050 487.050 ;
        RECT 281.700 478.800 282.600 483.900 ;
        RECT 289.950 481.950 292.050 484.050 ;
        RECT 281.700 477.900 288.300 478.800 ;
        RECT 281.700 477.600 282.600 477.900 ;
        RECT 257.400 471.600 259.200 477.600 ;
        RECT 268.800 471.600 270.600 477.600 ;
        RECT 280.800 471.600 282.600 477.600 ;
        RECT 286.800 477.600 288.300 477.900 ;
        RECT 302.400 477.600 303.600 489.900 ;
        RECT 310.950 489.450 315.000 490.050 ;
        RECT 316.950 489.450 319.050 490.050 ;
        RECT 305.100 488.100 306.900 488.850 ;
        RECT 310.950 488.550 319.050 489.450 ;
        RECT 310.950 487.950 315.000 488.550 ;
        RECT 316.950 487.950 319.050 488.550 ;
        RECT 320.100 486.900 321.150 491.100 ;
        RECT 334.950 490.950 340.050 493.050 ;
        RECT 322.950 487.950 325.050 490.050 ;
        RECT 332.100 488.100 333.900 488.850 ;
        RECT 319.950 483.600 321.150 486.900 ;
        RECT 286.800 471.600 288.600 477.600 ;
        RECT 302.400 471.600 304.200 477.600 ;
        RECT 319.500 471.600 321.300 483.600 ;
        RECT 335.400 477.600 336.600 489.900 ;
        RECT 338.100 488.100 339.900 488.850 ;
        RECT 337.950 484.950 340.050 487.050 ;
        RECT 344.550 483.600 345.750 493.950 ;
        RECT 374.100 493.050 375.900 494.850 ;
        RECT 358.950 490.800 361.050 493.050 ;
        RECT 371.100 490.800 372.900 491.400 ;
        RECT 346.950 485.400 348.750 487.200 ;
        RECT 347.850 484.200 352.050 485.400 ;
        RECT 358.050 484.200 358.950 489.900 ;
        RECT 364.950 487.950 367.050 490.050 ;
        RECT 368.100 489.600 372.900 490.800 ;
        RECT 366.750 485.700 368.550 486.000 ;
        RECT 376.950 485.700 377.850 500.400 ;
        RECT 386.400 501.300 388.200 506.400 ;
        RECT 392.400 501.300 394.200 506.400 ;
        RECT 386.400 499.950 394.200 501.300 ;
        RECT 395.400 500.400 397.200 506.400 ;
        RECT 395.400 498.300 396.600 500.400 ;
        RECT 408.000 499.200 409.800 506.400 ;
        RECT 423.000 499.200 424.800 506.400 ;
        RECT 442.200 499.200 444.000 506.400 ;
        RECT 408.000 498.300 411.600 499.200 ;
        RECT 423.000 498.300 426.600 499.200 ;
        RECT 392.850 497.250 396.600 498.300 ;
        RECT 392.850 497.100 394.050 497.250 ;
        RECT 385.950 493.950 388.050 496.050 ;
        RECT 391.950 493.950 394.050 496.050 ;
        RECT 410.400 494.100 411.600 498.300 ;
        RECT 425.400 494.100 426.600 498.300 ;
        RECT 440.400 498.300 444.000 499.200 ;
        RECT 456.000 499.200 457.800 506.400 ;
        RECT 469.800 500.400 471.600 506.400 ;
        RECT 456.000 498.300 459.600 499.200 ;
        RECT 440.400 494.100 441.600 498.300 ;
        RECT 458.400 494.100 459.600 498.300 ;
        RECT 470.400 498.300 471.600 500.400 ;
        RECT 472.800 501.300 474.600 506.400 ;
        RECT 478.800 501.300 480.600 506.400 ;
        RECT 472.800 499.950 480.600 501.300 ;
        RECT 490.800 500.400 492.600 506.400 ;
        RECT 491.400 498.300 492.600 500.400 ;
        RECT 493.800 501.300 495.600 506.400 ;
        RECT 499.800 501.300 501.600 506.400 ;
        RECT 493.800 499.950 501.600 501.300 ;
        RECT 509.400 501.300 511.200 506.400 ;
        RECT 515.400 501.300 517.200 506.400 ;
        RECT 509.400 499.950 517.200 501.300 ;
        RECT 518.400 500.400 520.200 506.400 ;
        RECT 530.400 503.400 532.200 506.400 ;
        RECT 518.400 498.300 519.600 500.400 ;
        RECT 530.400 500.100 531.600 503.400 ;
        RECT 547.200 502.050 549.000 506.400 ;
        RECT 563.400 503.400 565.200 506.400 ;
        RECT 581.400 503.400 583.200 506.400 ;
        RECT 547.200 500.400 552.600 502.050 ;
        RECT 470.400 497.250 474.150 498.300 ;
        RECT 491.400 497.250 495.150 498.300 ;
        RECT 472.950 497.100 474.150 497.250 ;
        RECT 493.950 497.100 495.150 497.250 ;
        RECT 515.850 497.250 519.600 498.300 ;
        RECT 529.950 498.450 532.050 499.050 ;
        RECT 538.950 498.450 541.050 499.050 ;
        RECT 529.950 497.550 541.050 498.450 ;
        RECT 515.850 497.100 517.050 497.250 ;
        RECT 529.950 496.950 532.050 497.550 ;
        RECT 538.950 496.950 541.050 497.550 ;
        RECT 551.700 497.100 552.600 500.400 ;
        RECT 563.400 500.100 564.600 503.400 ;
        RECT 577.950 501.450 580.050 502.050 ;
        RECT 572.550 500.550 580.050 501.450 ;
        RECT 562.950 498.450 565.050 499.050 ;
        RECT 572.550 498.450 573.450 500.550 ;
        RECT 577.950 499.950 580.050 500.550 ;
        RECT 562.950 497.550 573.450 498.450 ;
        RECT 562.950 496.950 565.050 497.550 ;
        RECT 472.950 493.950 475.050 496.050 ;
        RECT 478.950 493.950 481.050 496.050 ;
        RECT 493.950 493.950 496.050 496.050 ;
        RECT 499.950 493.950 502.050 496.050 ;
        RECT 508.950 493.950 511.050 496.050 ;
        RECT 514.950 493.950 517.050 496.050 ;
        RECT 530.700 494.100 532.050 495.900 ;
        RECT 386.100 492.150 387.900 492.900 ;
        RECT 389.100 491.100 390.900 491.850 ;
        RECT 391.950 491.100 393.150 492.900 ;
        RECT 400.950 492.450 403.050 493.050 ;
        RECT 409.950 492.450 412.050 493.050 ;
        RECT 395.100 491.100 396.900 491.850 ;
        RECT 400.950 491.550 412.050 492.450 ;
        RECT 388.950 487.950 391.050 490.050 ;
        RECT 392.100 486.900 393.150 491.100 ;
        RECT 400.950 490.950 403.050 491.550 ;
        RECT 409.950 490.950 412.050 491.550 ;
        RECT 424.950 492.450 427.050 493.050 ;
        RECT 429.000 492.450 433.050 493.050 ;
        RECT 424.950 491.550 433.050 492.450 ;
        RECT 424.950 490.950 427.050 491.550 ;
        RECT 429.000 490.950 433.050 491.550 ;
        RECT 439.950 492.450 442.050 493.050 ;
        RECT 448.950 492.450 451.050 493.050 ;
        RECT 439.950 491.550 451.050 492.450 ;
        RECT 439.950 490.950 442.050 491.550 ;
        RECT 448.950 490.950 451.050 491.550 ;
        RECT 457.950 492.450 460.050 493.050 ;
        RECT 462.000 492.450 466.050 493.050 ;
        RECT 457.950 491.550 466.050 492.450 ;
        RECT 457.950 490.950 460.050 491.550 ;
        RECT 462.000 490.950 466.050 491.550 ;
        RECT 470.100 491.100 471.900 491.850 ;
        RECT 473.850 491.100 475.050 492.900 ;
        RECT 479.100 492.150 480.900 492.900 ;
        RECT 476.100 491.100 477.900 491.850 ;
        RECT 491.100 491.100 492.900 491.850 ;
        RECT 494.850 491.100 496.050 492.900 ;
        RECT 500.100 492.150 501.900 492.900 ;
        RECT 509.100 492.150 510.900 492.900 ;
        RECT 497.100 491.100 498.900 491.850 ;
        RECT 512.100 491.100 513.900 491.850 ;
        RECT 514.950 491.100 516.150 492.900 ;
        RECT 518.100 491.100 519.900 491.850 ;
        RECT 394.950 487.950 397.050 490.050 ;
        RECT 407.100 488.100 408.900 488.850 ;
        RECT 366.750 485.100 377.850 485.700 ;
        RECT 335.400 471.600 337.200 477.600 ;
        RECT 344.550 471.600 346.350 483.600 ;
        RECT 349.950 483.300 352.050 484.200 ;
        RECT 352.950 483.300 358.950 484.200 ;
        RECT 360.150 484.500 377.850 485.100 ;
        RECT 360.150 484.200 368.550 484.500 ;
        RECT 352.950 482.400 353.850 483.300 ;
        RECT 351.150 480.600 353.850 482.400 ;
        RECT 354.750 482.100 356.550 482.400 ;
        RECT 360.150 482.100 361.050 484.200 ;
        RECT 376.950 483.600 377.850 484.500 ;
        RECT 391.950 483.600 393.150 486.900 ;
        RECT 354.750 481.200 361.050 482.100 ;
        RECT 361.950 482.700 363.750 483.300 ;
        RECT 361.950 481.500 369.450 482.700 ;
        RECT 354.750 480.600 356.550 481.200 ;
        RECT 368.250 480.600 369.450 481.500 ;
        RECT 349.950 477.600 353.850 479.700 ;
        RECT 358.950 479.550 360.750 480.300 ;
        RECT 363.750 479.550 365.550 480.300 ;
        RECT 358.950 478.500 365.550 479.550 ;
        RECT 368.250 478.500 373.050 480.600 ;
        RECT 352.050 471.600 353.850 477.600 ;
        RECT 359.850 471.600 361.650 478.500 ;
        RECT 368.250 477.600 369.450 478.500 ;
        RECT 367.650 471.600 369.450 477.600 ;
        RECT 376.050 471.600 377.850 483.600 ;
        RECT 391.500 471.600 393.300 483.600 ;
        RECT 410.400 477.600 411.600 489.900 ;
        RECT 413.100 488.100 414.900 488.850 ;
        RECT 422.100 488.100 423.900 488.850 ;
        RECT 412.950 484.950 415.050 487.050 ;
        RECT 421.950 484.950 424.050 487.050 ;
        RECT 425.400 477.600 426.600 489.900 ;
        RECT 428.100 488.100 429.900 488.850 ;
        RECT 437.100 488.100 438.900 488.850 ;
        RECT 427.950 484.950 430.050 487.050 ;
        RECT 409.800 471.600 411.600 477.600 ;
        RECT 424.800 471.600 426.600 477.600 ;
        RECT 440.400 477.600 441.600 489.900 ;
        RECT 443.100 488.100 444.900 488.850 ;
        RECT 455.100 488.100 456.900 488.850 ;
        RECT 442.950 484.950 445.050 487.050 ;
        RECT 454.950 484.950 457.050 487.050 ;
        RECT 458.400 477.600 459.600 489.900 ;
        RECT 461.100 488.100 462.900 488.850 ;
        RECT 469.950 487.950 472.050 490.050 ;
        RECT 460.950 484.950 463.050 487.050 ;
        RECT 473.850 486.900 474.900 491.100 ;
        RECT 475.950 487.950 478.050 490.050 ;
        RECT 490.950 487.950 493.050 490.050 ;
        RECT 494.850 486.900 495.900 491.100 ;
        RECT 496.950 487.950 499.050 490.050 ;
        RECT 511.950 487.950 514.050 490.050 ;
        RECT 515.100 486.900 516.150 491.100 ;
        RECT 517.950 487.950 520.050 490.050 ;
        RECT 526.950 487.950 529.050 490.050 ;
        RECT 530.700 489.900 531.900 494.100 ;
        RECT 544.950 493.950 547.050 496.050 ;
        RECT 550.950 493.950 556.050 496.050 ;
        RECT 563.700 494.100 565.050 495.900 ;
        RECT 532.950 490.950 535.050 493.050 ;
        RECT 545.100 492.150 546.900 492.900 ;
        RECT 542.100 491.100 543.900 491.850 ;
        RECT 548.100 491.100 549.900 491.850 ;
        RECT 473.850 483.600 475.050 486.900 ;
        RECT 494.850 483.600 496.050 486.900 ;
        RECT 514.950 483.600 516.150 486.900 ;
        RECT 527.100 486.150 528.900 486.900 ;
        RECT 530.700 484.650 532.050 489.900 ;
        RECT 533.100 489.150 534.900 489.900 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 547.950 487.950 550.050 490.050 ;
        RECT 530.700 483.600 533.400 484.650 ;
        RECT 551.700 483.600 552.600 492.900 ;
        RECT 559.950 487.950 562.050 490.050 ;
        RECT 563.700 489.900 564.900 494.100 ;
        RECT 577.950 493.950 580.050 496.050 ;
        RECT 565.950 490.950 568.050 493.050 ;
        RECT 578.100 492.150 579.900 492.900 ;
        RECT 581.400 491.100 582.600 503.400 ;
        RECT 597.000 499.200 598.800 506.400 ;
        RECT 613.800 503.400 615.600 506.400 ;
        RECT 597.000 498.300 600.600 499.200 ;
        RECT 599.400 494.100 600.600 498.300 ;
        RECT 598.950 492.450 601.050 493.050 ;
        RECT 607.950 492.450 610.050 493.050 ;
        RECT 598.950 491.550 610.050 492.450 ;
        RECT 598.950 490.950 601.050 491.550 ;
        RECT 607.950 490.950 610.050 491.550 ;
        RECT 614.400 491.100 615.600 503.400 ;
        RECT 629.100 498.000 630.900 506.400 ;
        RECT 646.800 503.400 648.600 506.400 ;
        RECT 629.100 496.350 633.300 498.000 ;
        RECT 616.950 493.950 619.050 496.050 ;
        RECT 629.100 494.100 630.900 494.850 ;
        RECT 617.100 492.150 618.900 492.900 ;
        RECT 628.950 490.950 631.050 493.050 ;
        RECT 560.100 486.150 561.900 486.900 ;
        RECT 563.700 484.650 565.050 489.900 ;
        RECT 566.100 489.150 567.900 489.900 ;
        RECT 580.950 489.450 583.050 490.050 ;
        RECT 585.000 489.450 589.050 490.050 ;
        RECT 580.950 488.550 589.050 489.450 ;
        RECT 580.950 487.950 583.050 488.550 ;
        RECT 585.000 487.950 589.050 488.550 ;
        RECT 596.100 488.100 597.900 488.850 ;
        RECT 563.700 483.600 566.400 484.650 ;
        RECT 440.400 471.600 442.200 477.600 ;
        RECT 457.800 471.600 459.600 477.600 ;
        RECT 473.700 471.600 475.500 483.600 ;
        RECT 494.700 471.600 496.500 483.600 ;
        RECT 514.500 471.600 516.300 483.600 ;
        RECT 531.600 471.600 533.400 483.600 ;
        RECT 542.400 482.700 550.200 483.600 ;
        RECT 542.400 471.600 544.200 482.700 ;
        RECT 548.400 471.600 550.200 482.700 ;
        RECT 551.400 471.600 553.200 483.600 ;
        RECT 564.600 471.600 566.400 483.600 ;
        RECT 581.400 477.600 582.600 486.900 ;
        RECT 595.950 484.950 598.050 487.050 ;
        RECT 599.400 477.600 600.600 489.900 ;
        RECT 613.950 489.450 616.050 490.050 ;
        RECT 618.000 489.450 622.050 490.050 ;
        RECT 602.100 488.100 603.900 488.850 ;
        RECT 613.950 488.550 622.050 489.450 ;
        RECT 613.950 487.950 616.050 488.550 ;
        RECT 618.000 487.950 622.050 488.550 ;
        RECT 625.950 487.950 628.050 490.050 ;
        RECT 632.400 488.100 633.300 496.350 ;
        RECT 647.400 491.100 648.600 503.400 ;
        RECT 656.400 501.300 658.200 506.400 ;
        RECT 662.400 501.300 664.200 506.400 ;
        RECT 656.400 499.950 664.200 501.300 ;
        RECT 665.400 500.400 667.200 506.400 ;
        RECT 674.400 501.300 676.200 506.400 ;
        RECT 680.400 501.300 682.200 506.400 ;
        RECT 665.400 498.300 666.600 500.400 ;
        RECT 674.400 499.950 682.200 501.300 ;
        RECT 683.400 500.400 685.200 506.400 ;
        RECT 683.400 498.300 684.600 500.400 ;
        RECT 662.850 497.250 666.600 498.300 ;
        RECT 680.850 497.250 684.600 498.300 ;
        RECT 698.100 498.000 699.900 506.400 ;
        RECT 713.400 501.300 715.200 506.400 ;
        RECT 719.400 501.300 721.200 506.400 ;
        RECT 713.400 499.950 721.200 501.300 ;
        RECT 722.400 500.400 724.200 506.400 ;
        RECT 736.800 503.400 738.600 506.400 ;
        RECT 722.400 498.300 723.600 500.400 ;
        RECT 662.850 497.100 664.050 497.250 ;
        RECT 680.850 497.100 682.050 497.250 ;
        RECT 695.700 496.350 699.900 498.000 ;
        RECT 719.850 497.250 723.600 498.300 ;
        RECT 719.850 497.100 721.050 497.250 ;
        RECT 649.950 493.950 652.050 496.050 ;
        RECT 655.950 493.950 658.050 496.050 ;
        RECT 661.950 495.450 664.050 496.050 ;
        RECT 666.000 495.450 670.050 496.050 ;
        RECT 661.950 494.550 670.050 495.450 ;
        RECT 661.950 493.950 664.050 494.550 ;
        RECT 666.000 493.950 670.050 494.550 ;
        RECT 673.950 493.950 676.050 496.050 ;
        RECT 679.950 495.450 682.050 496.050 ;
        RECT 684.000 495.450 688.050 496.050 ;
        RECT 679.950 494.550 688.050 495.450 ;
        RECT 679.950 493.950 682.050 494.550 ;
        RECT 684.000 493.950 688.050 494.550 ;
        RECT 650.100 492.150 651.900 492.900 ;
        RECT 656.100 492.150 657.900 492.900 ;
        RECT 659.100 491.100 660.900 491.850 ;
        RECT 661.950 491.100 663.150 492.900 ;
        RECT 674.100 492.150 675.900 492.900 ;
        RECT 665.100 491.100 666.900 491.850 ;
        RECT 677.100 491.100 678.900 491.850 ;
        RECT 679.950 491.100 681.150 492.900 ;
        RECT 683.100 491.100 684.900 491.850 ;
        RECT 640.950 490.050 643.050 490.200 ;
        RECT 640.950 489.450 645.000 490.050 ;
        RECT 646.950 489.450 649.050 490.050 ;
        RECT 640.950 488.550 649.050 489.450 ;
        RECT 640.950 488.100 645.000 488.550 ;
        RECT 642.000 487.950 645.000 488.100 ;
        RECT 646.950 487.950 649.050 488.550 ;
        RECT 658.950 487.950 661.050 490.050 ;
        RECT 601.950 484.950 604.050 487.050 ;
        RECT 614.400 477.600 615.600 486.900 ;
        RECT 626.100 486.150 627.900 486.900 ;
        RECT 631.950 486.450 634.050 487.050 ;
        RECT 662.100 486.900 663.150 491.100 ;
        RECT 664.950 487.950 667.050 490.050 ;
        RECT 676.950 487.950 679.050 490.050 ;
        RECT 680.100 486.900 681.150 491.100 ;
        RECT 682.950 487.950 685.050 490.050 ;
        RECT 695.700 488.100 696.600 496.350 ;
        RECT 698.100 494.100 699.900 494.850 ;
        RECT 712.950 493.950 715.050 496.050 ;
        RECT 718.950 493.950 721.050 496.050 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 713.100 492.150 714.900 492.900 ;
        RECT 716.100 491.100 717.900 491.850 ;
        RECT 718.950 491.100 720.150 492.900 ;
        RECT 722.100 491.100 723.900 491.850 ;
        RECT 737.400 491.100 738.600 503.400 ;
        RECT 754.200 499.200 756.000 506.400 ;
        RECT 767.400 501.300 769.200 506.400 ;
        RECT 773.400 501.300 775.200 506.400 ;
        RECT 767.400 499.950 775.200 501.300 ;
        RECT 776.400 500.400 778.200 506.400 ;
        RECT 752.400 498.300 756.000 499.200 ;
        RECT 776.400 498.300 777.600 500.400 ;
        RECT 789.000 499.200 790.800 506.400 ;
        RECT 789.000 498.300 792.600 499.200 ;
        RECT 739.950 493.950 742.050 496.050 ;
        RECT 752.400 494.100 753.600 498.300 ;
        RECT 773.850 497.250 777.600 498.300 ;
        RECT 773.850 497.100 775.050 497.250 ;
        RECT 766.950 493.950 769.050 496.050 ;
        RECT 772.950 495.450 775.050 496.050 ;
        RECT 781.950 495.450 784.050 496.050 ;
        RECT 772.950 494.550 784.050 495.450 ;
        RECT 772.950 493.950 775.050 494.550 ;
        RECT 781.950 493.950 784.050 494.550 ;
        RECT 791.400 494.100 792.600 498.300 ;
        RECT 806.100 498.000 807.900 506.400 ;
        RECT 803.700 496.350 807.900 498.000 ;
        RECT 824.400 503.400 826.200 506.400 ;
        RECT 740.100 492.150 741.900 492.900 ;
        RECT 745.950 492.450 750.000 493.050 ;
        RECT 751.950 492.450 754.050 493.050 ;
        RECT 745.950 491.550 754.050 492.450 ;
        RECT 767.100 492.150 768.900 492.900 ;
        RECT 700.950 487.950 703.050 490.200 ;
        RECT 715.950 487.950 718.050 490.050 ;
        RECT 640.950 486.450 643.050 486.900 ;
        RECT 623.100 485.100 624.900 485.850 ;
        RECT 631.950 485.550 643.050 486.450 ;
        RECT 631.950 484.950 634.050 485.550 ;
        RECT 640.950 484.800 643.050 485.550 ;
        RECT 622.950 481.950 625.050 484.050 ;
        RECT 632.400 478.800 633.300 483.900 ;
        RECT 626.700 477.900 633.300 478.800 ;
        RECT 626.700 477.600 628.200 477.900 ;
        RECT 581.400 471.600 583.200 477.600 ;
        RECT 598.800 471.600 600.600 477.600 ;
        RECT 613.800 471.600 615.600 477.600 ;
        RECT 626.400 471.600 628.200 477.600 ;
        RECT 632.400 477.600 633.300 477.900 ;
        RECT 647.400 477.600 648.600 486.900 ;
        RECT 661.950 483.600 663.150 486.900 ;
        RECT 679.950 483.600 681.150 486.900 ;
        RECT 688.950 486.450 693.000 487.050 ;
        RECT 694.950 486.450 697.050 487.050 ;
        RECT 719.100 486.900 720.150 491.100 ;
        RECT 745.950 490.950 750.000 491.550 ;
        RECT 751.950 490.950 754.050 491.550 ;
        RECT 770.100 491.100 771.900 491.850 ;
        RECT 772.950 491.100 774.150 492.900 ;
        RECT 790.950 492.450 793.050 493.050 ;
        RECT 776.100 491.100 777.900 491.850 ;
        RECT 782.550 491.550 793.050 492.450 ;
        RECT 721.950 487.950 724.050 490.050 ;
        RECT 730.950 489.450 735.000 490.050 ;
        RECT 736.950 489.450 739.050 490.050 ;
        RECT 730.950 488.550 739.050 489.450 ;
        RECT 730.950 487.950 735.000 488.550 ;
        RECT 736.950 487.950 739.050 488.550 ;
        RECT 749.100 488.100 750.900 488.850 ;
        RECT 688.950 485.550 697.050 486.450 ;
        RECT 701.100 486.150 702.900 486.900 ;
        RECT 688.950 484.950 693.000 485.550 ;
        RECT 694.950 484.950 697.050 485.550 ;
        RECT 704.100 485.100 705.900 485.850 ;
        RECT 632.400 471.600 634.200 477.600 ;
        RECT 646.800 471.600 648.600 477.600 ;
        RECT 661.500 471.600 663.300 483.600 ;
        RECT 679.500 471.600 681.300 483.600 ;
        RECT 695.700 478.800 696.600 483.900 ;
        RECT 700.950 481.950 706.050 484.050 ;
        RECT 718.950 483.600 720.150 486.900 ;
        RECT 695.700 477.900 702.300 478.800 ;
        RECT 695.700 477.600 696.600 477.900 ;
        RECT 694.800 471.600 696.600 477.600 ;
        RECT 700.800 477.600 702.300 477.900 ;
        RECT 700.800 471.600 702.600 477.600 ;
        RECT 718.500 471.600 720.300 483.600 ;
        RECT 737.400 477.600 738.600 486.900 ;
        RECT 748.950 484.950 751.050 487.050 ;
        RECT 736.800 471.600 738.600 477.600 ;
        RECT 752.400 477.600 753.600 489.900 ;
        RECT 755.100 488.100 756.900 488.850 ;
        RECT 769.950 487.950 772.050 490.050 ;
        RECT 754.950 484.950 757.050 487.050 ;
        RECT 773.100 486.900 774.150 491.100 ;
        RECT 775.950 487.950 778.050 490.050 ;
        RECT 772.950 483.600 774.150 486.900 ;
        RECT 782.550 483.900 783.450 491.550 ;
        RECT 790.950 490.950 793.050 491.550 ;
        RECT 788.100 488.100 789.900 488.850 ;
        RECT 787.950 484.950 790.050 487.050 ;
        RECT 752.400 471.600 754.200 477.600 ;
        RECT 772.500 471.600 774.300 483.600 ;
        RECT 781.950 481.800 784.050 483.900 ;
        RECT 791.400 477.600 792.600 489.900 ;
        RECT 794.100 488.100 795.900 488.850 ;
        RECT 803.700 488.100 804.600 496.350 ;
        RECT 806.100 494.100 807.900 494.850 ;
        RECT 820.950 493.950 823.050 496.050 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 821.100 492.150 822.900 492.900 ;
        RECT 824.400 491.100 825.600 503.400 ;
        RECT 808.950 487.950 811.050 490.050 ;
        RECT 814.950 489.450 817.050 490.050 ;
        RECT 823.950 489.450 826.050 490.050 ;
        RECT 814.950 488.550 826.050 489.450 ;
        RECT 814.950 487.950 817.050 488.550 ;
        RECT 823.950 487.950 826.050 488.550 ;
        RECT 793.950 484.950 796.050 487.050 ;
        RECT 802.950 484.950 805.050 487.050 ;
        RECT 809.100 486.150 810.900 486.900 ;
        RECT 812.100 485.100 813.900 485.850 ;
        RECT 803.700 478.800 804.600 483.900 ;
        RECT 811.950 481.950 814.050 484.050 ;
        RECT 803.700 477.900 810.300 478.800 ;
        RECT 803.700 477.600 804.600 477.900 ;
        RECT 790.800 471.600 792.600 477.600 ;
        RECT 802.800 471.600 804.600 477.600 ;
        RECT 808.800 477.600 810.300 477.900 ;
        RECT 824.400 477.600 825.600 486.900 ;
        RECT 808.800 471.600 810.600 477.600 ;
        RECT 824.400 471.600 826.200 477.600 ;
        RECT 7.800 461.400 9.600 467.400 ;
        RECT 8.700 461.100 9.600 461.400 ;
        RECT 13.800 461.400 15.600 467.400 ;
        RECT 13.800 461.100 15.300 461.400 ;
        RECT 8.700 460.200 15.300 461.100 ;
        RECT 8.700 455.100 9.600 460.200 ;
        RECT 16.950 454.950 19.050 457.050 ;
        RECT 23.400 456.300 25.200 467.400 ;
        RECT 29.400 456.300 31.200 467.400 ;
        RECT 23.400 455.400 31.200 456.300 ;
        RECT 32.400 455.400 34.200 467.400 ;
        RECT 50.700 455.400 52.500 467.400 ;
        RECT 64.800 461.400 66.600 467.400 ;
        RECT 65.700 461.100 66.600 461.400 ;
        RECT 70.800 461.400 72.600 467.400 ;
        RECT 85.800 461.400 87.600 467.400 ;
        RECT 70.800 461.100 72.300 461.400 ;
        RECT 65.700 460.200 72.300 461.100 ;
        RECT 86.700 461.100 87.600 461.400 ;
        RECT 91.800 461.400 93.600 467.400 ;
        RECT 91.800 461.100 93.300 461.400 ;
        RECT 86.700 460.200 93.300 461.100 ;
        RECT 4.950 451.950 10.050 454.050 ;
        RECT 17.100 453.150 18.900 453.900 ;
        RECT 14.100 452.100 15.900 452.850 ;
        RECT 8.700 442.650 9.600 450.900 ;
        RECT 13.950 448.950 16.050 451.050 ;
        RECT 22.950 448.950 25.050 451.050 ;
        RECT 28.950 448.950 31.050 451.050 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 23.100 447.150 24.900 447.900 ;
        RECT 29.100 447.150 30.900 447.900 ;
        RECT 26.100 446.100 27.900 446.850 ;
        RECT 32.700 446.100 33.600 455.400 ;
        RECT 50.850 452.100 52.050 455.400 ;
        RECT 65.700 455.100 66.600 460.200 ;
        RECT 73.950 454.950 76.050 457.050 ;
        RECT 86.700 455.100 87.600 460.200 ;
        RECT 94.950 454.950 97.050 457.050 ;
        RECT 110.700 455.400 112.500 467.400 ;
        RECT 130.500 455.400 132.300 467.400 ;
        RECT 148.800 461.400 150.600 467.400 ;
        RECT 46.950 448.950 49.050 451.050 ;
        RECT 50.850 447.900 51.900 452.100 ;
        RECT 64.950 451.950 67.050 454.050 ;
        RECT 74.100 453.150 75.900 453.900 ;
        RECT 79.950 453.450 84.000 454.050 ;
        RECT 85.950 453.450 88.050 454.050 ;
        RECT 71.100 452.100 72.900 452.850 ;
        RECT 79.950 452.550 88.050 453.450 ;
        RECT 95.100 453.150 96.900 453.900 ;
        RECT 79.950 451.950 84.000 452.550 ;
        RECT 85.950 451.950 88.050 452.550 ;
        RECT 92.100 452.100 93.900 452.850 ;
        RECT 110.850 452.100 112.050 455.400 ;
        RECT 130.950 452.100 132.150 455.400 ;
        RECT 149.400 452.100 150.600 461.400 ;
        RECT 164.700 455.400 166.500 467.400 ;
        RECT 180.600 455.400 182.400 467.400 ;
        RECT 164.850 452.100 166.050 455.400 ;
        RECT 179.700 454.350 182.400 455.400 ;
        RECT 197.400 461.400 199.200 467.400 ;
        RECT 215.400 461.400 217.200 467.400 ;
        RECT 176.100 452.100 177.900 452.850 ;
        RECT 52.950 448.950 55.050 451.050 ;
        RECT 47.100 447.150 48.900 447.900 ;
        RECT 50.850 446.100 52.050 447.900 ;
        RECT 53.100 447.150 54.900 447.900 ;
        RECT 56.100 446.100 57.900 446.850 ;
        RECT 11.100 444.150 12.900 444.900 ;
        RECT 25.950 442.950 28.050 445.050 ;
        RECT 31.950 442.950 37.050 445.050 ;
        RECT 43.950 444.450 48.000 445.050 ;
        RECT 49.950 444.450 52.050 445.050 ;
        RECT 43.950 443.550 52.050 444.450 ;
        RECT 43.950 442.950 48.000 443.550 ;
        RECT 49.950 442.950 52.050 443.550 ;
        RECT 55.950 442.950 58.050 445.050 ;
        RECT 65.700 442.650 66.600 450.900 ;
        RECT 70.950 448.950 73.050 451.050 ;
        RECT 67.950 445.950 70.050 448.050 ;
        RECT 68.100 444.150 69.900 444.900 ;
        RECT 86.700 442.650 87.600 450.900 ;
        RECT 91.950 448.950 94.050 451.050 ;
        RECT 106.950 448.950 109.050 451.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 110.850 447.900 111.900 452.100 ;
        RECT 112.950 448.950 115.050 451.050 ;
        RECT 127.950 448.950 130.050 451.050 ;
        RECT 131.100 447.900 132.150 452.100 ;
        RECT 133.950 448.950 136.050 451.050 ;
        RECT 139.950 450.450 142.050 451.050 ;
        RECT 148.950 450.450 151.050 451.050 ;
        RECT 139.950 449.550 151.050 450.450 ;
        RECT 139.950 448.950 142.050 449.550 ;
        RECT 148.950 448.950 151.050 449.550 ;
        RECT 160.950 448.950 163.050 451.050 ;
        RECT 164.850 447.900 165.900 452.100 ;
        RECT 166.950 448.950 169.050 451.050 ;
        RECT 175.950 448.950 178.050 451.050 ;
        RECT 179.700 449.100 181.050 454.350 ;
        RECT 184.950 453.450 187.050 454.050 ;
        RECT 193.950 453.450 196.050 454.050 ;
        RECT 184.950 452.550 196.050 453.450 ;
        RECT 184.950 451.950 187.050 452.550 ;
        RECT 193.950 451.950 196.050 452.550 ;
        RECT 194.100 450.150 195.900 450.900 ;
        RECT 182.100 449.100 183.900 449.850 ;
        RECT 197.400 449.100 198.600 461.400 ;
        RECT 211.950 451.950 214.050 454.050 ;
        RECT 200.100 450.150 201.900 450.900 ;
        RECT 212.100 450.150 213.900 450.900 ;
        RECT 215.400 449.100 216.600 461.400 ;
        RECT 230.400 456.600 232.200 467.400 ;
        RECT 236.400 466.500 244.200 467.400 ;
        RECT 236.400 456.600 238.200 466.500 ;
        RECT 230.400 455.700 238.200 456.600 ;
        RECT 239.400 454.500 241.200 465.600 ;
        RECT 242.400 455.400 244.200 466.500 ;
        RECT 253.800 461.400 255.600 467.400 ;
        RECT 217.950 451.950 220.050 454.050 ;
        RECT 237.150 453.600 241.200 454.500 ;
        RECT 237.150 452.100 238.050 453.600 ;
        RECT 254.400 452.100 255.600 461.400 ;
        RECT 266.400 461.400 268.200 467.400 ;
        RECT 218.100 450.150 219.900 450.900 ;
        RECT 107.100 447.150 108.900 447.900 ;
        RECT 110.850 446.100 112.050 447.900 ;
        RECT 113.100 447.150 114.900 447.900 ;
        RECT 128.100 447.150 129.900 447.900 ;
        RECT 116.100 446.100 117.900 446.850 ;
        RECT 125.100 446.100 126.900 446.850 ;
        RECT 130.950 446.100 132.150 447.900 ;
        RECT 134.100 447.150 135.900 447.900 ;
        RECT 89.100 444.150 90.900 444.900 ;
        RECT 94.950 444.450 97.050 445.050 ;
        RECT 109.950 444.450 112.050 445.050 ;
        RECT 94.950 443.550 112.050 444.450 ;
        RECT 94.950 442.950 97.050 443.550 ;
        RECT 109.950 442.950 112.050 443.550 ;
        RECT 115.950 442.950 118.050 445.050 ;
        RECT 124.950 442.950 127.050 445.050 ;
        RECT 130.950 442.950 133.050 445.050 ;
        RECT 8.700 441.000 12.900 442.650 ;
        RECT 11.100 432.600 12.900 441.000 ;
        RECT 32.700 438.600 33.600 441.900 ;
        RECT 49.950 441.750 51.150 441.900 ;
        RECT 47.400 440.700 51.150 441.750 ;
        RECT 65.700 441.000 69.900 442.650 ;
        RECT 86.700 441.000 90.900 442.650 ;
        RECT 109.950 441.750 111.150 441.900 ;
        RECT 47.400 438.600 48.600 440.700 ;
        RECT 28.200 436.950 33.600 438.600 ;
        RECT 28.200 432.600 30.000 436.950 ;
        RECT 46.800 432.600 48.600 438.600 ;
        RECT 49.800 437.700 57.600 439.050 ;
        RECT 49.800 432.600 51.600 437.700 ;
        RECT 55.800 432.600 57.600 437.700 ;
        RECT 68.100 432.600 69.900 441.000 ;
        RECT 89.100 432.600 90.900 441.000 ;
        RECT 107.400 440.700 111.150 441.750 ;
        RECT 131.850 441.750 133.050 441.900 ;
        RECT 131.850 440.700 135.600 441.750 ;
        RECT 107.400 438.600 108.600 440.700 ;
        RECT 106.800 432.600 108.600 438.600 ;
        RECT 109.800 437.700 117.600 439.050 ;
        RECT 109.800 432.600 111.600 437.700 ;
        RECT 115.800 432.600 117.600 437.700 ;
        RECT 125.400 437.700 133.200 439.050 ;
        RECT 125.400 432.600 127.200 437.700 ;
        RECT 131.400 432.600 133.200 437.700 ;
        RECT 134.400 438.600 135.600 440.700 ;
        RECT 134.400 432.600 136.200 438.600 ;
        RECT 149.400 435.600 150.600 447.900 ;
        RECT 161.100 447.150 162.900 447.900 ;
        RECT 152.100 446.100 153.900 446.850 ;
        RECT 164.850 446.100 166.050 447.900 ;
        RECT 167.100 447.150 168.900 447.900 ;
        RECT 170.100 446.100 171.900 446.850 ;
        RECT 151.950 442.950 154.050 445.050 ;
        RECT 157.950 444.450 162.000 445.050 ;
        RECT 163.950 444.450 166.050 445.050 ;
        RECT 157.950 443.550 166.050 444.450 ;
        RECT 157.950 442.950 162.000 443.550 ;
        RECT 163.950 442.950 166.050 443.550 ;
        RECT 169.950 442.950 172.050 445.050 ;
        RECT 179.700 444.900 180.900 449.100 ;
        RECT 232.950 448.950 235.050 451.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 190.950 447.450 195.000 448.050 ;
        RECT 196.950 447.450 199.050 448.050 ;
        RECT 190.950 446.550 199.050 447.450 ;
        RECT 190.950 445.950 195.000 446.550 ;
        RECT 196.950 445.950 199.050 446.550 ;
        RECT 202.950 447.450 205.050 448.050 ;
        RECT 214.950 447.450 217.050 448.050 ;
        RECT 237.150 447.900 237.900 452.100 ;
        RECT 238.950 448.950 241.050 451.050 ;
        RECT 250.950 448.950 256.050 451.050 ;
        RECT 263.100 449.100 264.900 449.850 ;
        RECT 202.950 446.550 217.050 447.450 ;
        RECT 233.250 447.150 235.050 447.900 ;
        RECT 202.950 445.950 205.050 446.550 ;
        RECT 214.950 445.950 217.050 446.550 ;
        RECT 230.250 446.100 232.050 446.850 ;
        RECT 237.150 446.100 238.050 447.900 ;
        RECT 238.950 447.150 240.750 447.900 ;
        RECT 242.100 446.100 243.900 446.850 ;
        RECT 179.700 443.100 181.050 444.900 ;
        RECT 163.950 441.750 165.150 441.900 ;
        RECT 161.400 440.700 165.150 441.750 ;
        RECT 161.400 438.600 162.600 440.700 ;
        RECT 178.950 439.800 181.050 442.050 ;
        RECT 197.400 440.700 198.600 444.900 ;
        RECT 215.400 440.700 216.600 444.900 ;
        RECT 229.950 442.950 232.050 445.050 ;
        RECT 235.950 442.950 238.050 445.050 ;
        RECT 241.950 444.450 244.050 445.050 ;
        RECT 246.000 444.450 250.050 445.050 ;
        RECT 241.950 443.550 250.050 444.450 ;
        RECT 241.950 442.950 244.050 443.550 ;
        RECT 246.000 442.950 250.050 443.550 ;
        RECT 197.400 439.800 201.000 440.700 ;
        RECT 215.400 439.800 219.000 440.700 ;
        RECT 148.800 432.600 150.600 435.600 ;
        RECT 160.800 432.600 162.600 438.600 ;
        RECT 163.800 437.700 171.600 439.050 ;
        RECT 163.800 432.600 165.600 437.700 ;
        RECT 169.800 432.600 171.600 437.700 ;
        RECT 179.400 435.600 180.600 438.900 ;
        RECT 179.400 432.600 181.200 435.600 ;
        RECT 199.200 432.600 201.000 439.800 ;
        RECT 217.200 432.600 219.000 439.800 ;
        RECT 235.950 438.600 237.000 441.900 ;
        RECT 235.200 432.600 237.000 438.600 ;
        RECT 254.400 435.600 255.600 447.900 ;
        RECT 257.100 446.100 258.900 446.850 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 256.950 442.950 259.050 445.050 ;
        RECT 266.400 441.300 267.450 461.400 ;
        RECT 273.000 455.400 274.800 467.400 ;
        RECT 286.800 455.400 288.600 467.400 ;
        RECT 289.800 456.300 291.600 467.400 ;
        RECT 295.800 456.300 297.600 467.400 ;
        RECT 308.400 461.400 310.200 467.400 ;
        RECT 308.700 461.100 310.200 461.400 ;
        RECT 314.400 461.400 316.200 467.400 ;
        RECT 314.400 461.100 315.300 461.400 ;
        RECT 308.700 460.200 315.300 461.100 ;
        RECT 289.800 455.400 297.600 456.300 ;
        RECT 268.950 448.950 271.050 451.050 ;
        RECT 269.100 447.150 270.900 447.900 ;
        RECT 273.000 446.100 274.050 455.400 ;
        RECT 287.400 446.100 288.300 455.400 ;
        RECT 304.950 454.950 307.050 457.050 ;
        RECT 314.400 455.100 315.300 460.200 ;
        RECT 328.500 455.400 330.300 467.400 ;
        RECT 338.550 455.400 340.350 467.400 ;
        RECT 346.050 461.400 347.850 467.400 ;
        RECT 343.950 459.300 347.850 461.400 ;
        RECT 353.850 460.500 355.650 467.400 ;
        RECT 361.650 461.400 363.450 467.400 ;
        RECT 362.250 460.500 363.450 461.400 ;
        RECT 352.950 459.450 359.550 460.500 ;
        RECT 352.950 458.700 354.750 459.450 ;
        RECT 357.750 458.700 359.550 459.450 ;
        RECT 362.250 458.400 367.050 460.500 ;
        RECT 345.150 456.600 347.850 458.400 ;
        RECT 348.750 457.800 350.550 458.400 ;
        RECT 348.750 456.900 355.050 457.800 ;
        RECT 362.250 457.500 363.450 458.400 ;
        RECT 348.750 456.600 350.550 456.900 ;
        RECT 346.950 455.700 347.850 456.600 ;
        RECT 305.100 453.150 306.900 453.900 ;
        RECT 313.950 453.450 316.050 454.050 ;
        RECT 318.000 453.450 322.050 454.050 ;
        RECT 308.100 452.100 309.900 452.850 ;
        RECT 313.950 452.550 322.050 453.450 ;
        RECT 313.950 451.950 316.050 452.550 ;
        RECT 318.000 451.950 322.050 452.550 ;
        RECT 328.950 452.100 330.150 455.400 ;
        RECT 289.950 448.950 292.050 451.050 ;
        RECT 295.950 448.950 298.050 451.050 ;
        RECT 307.950 448.950 310.050 451.050 ;
        RECT 290.100 447.150 291.900 447.900 ;
        RECT 296.100 447.150 297.900 447.900 ;
        RECT 293.100 446.100 294.900 446.850 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 268.950 442.950 276.900 445.050 ;
        RECT 277.950 444.450 280.050 445.050 ;
        RECT 286.950 444.450 289.050 445.050 ;
        RECT 277.950 443.550 289.050 444.450 ;
        RECT 277.950 442.950 280.050 443.550 ;
        RECT 286.950 442.950 289.050 443.550 ;
        RECT 292.950 444.450 295.050 445.050 ;
        RECT 304.950 444.450 307.050 445.050 ;
        RECT 292.950 443.550 307.050 444.450 ;
        RECT 311.100 444.150 312.900 444.900 ;
        RECT 292.950 442.950 295.050 443.550 ;
        RECT 304.950 442.950 307.050 443.550 ;
        RECT 314.400 442.650 315.300 450.900 ;
        RECT 325.950 448.800 328.050 451.050 ;
        RECT 329.100 447.900 330.150 452.100 ;
        RECT 331.950 448.950 334.050 451.050 ;
        RECT 326.100 447.150 327.900 447.900 ;
        RECT 323.100 446.100 324.900 446.850 ;
        RECT 328.950 446.100 330.150 447.900 ;
        RECT 332.100 447.150 333.900 447.900 ;
        RECT 338.550 445.050 339.750 455.400 ;
        RECT 343.950 454.800 346.050 455.700 ;
        RECT 346.950 454.800 352.950 455.700 ;
        RECT 341.850 453.600 346.050 454.800 ;
        RECT 340.950 451.800 342.750 453.600 ;
        RECT 352.050 449.100 352.950 454.800 ;
        RECT 354.150 454.800 355.050 456.900 ;
        RECT 355.950 456.300 363.450 457.500 ;
        RECT 355.950 455.700 357.750 456.300 ;
        RECT 370.050 455.400 371.850 467.400 ;
        RECT 354.150 454.500 362.550 454.800 ;
        RECT 370.950 454.500 371.850 455.400 ;
        RECT 354.150 453.900 371.850 454.500 ;
        RECT 360.750 453.300 371.850 453.900 ;
        RECT 377.400 461.400 379.200 467.400 ;
        RECT 377.400 454.500 378.600 461.400 ;
        RECT 383.700 455.400 385.500 467.400 ;
        RECT 390.150 455.400 391.950 467.400 ;
        RECT 398.550 461.400 400.350 467.400 ;
        RECT 398.550 460.500 399.750 461.400 ;
        RECT 406.350 460.500 408.150 467.400 ;
        RECT 414.150 461.400 415.950 467.400 ;
        RECT 394.950 458.400 399.750 460.500 ;
        RECT 402.450 459.450 409.050 460.500 ;
        RECT 402.450 458.700 404.250 459.450 ;
        RECT 407.250 458.700 409.050 459.450 ;
        RECT 414.150 459.300 418.050 461.400 ;
        RECT 398.550 457.500 399.750 458.400 ;
        RECT 411.450 457.800 413.250 458.400 ;
        RECT 398.550 456.300 406.050 457.500 ;
        RECT 404.250 455.700 406.050 456.300 ;
        RECT 406.950 456.900 413.250 457.800 ;
        RECT 377.400 453.600 383.100 454.500 ;
        RECT 360.750 453.000 362.550 453.300 ;
        RECT 358.950 448.950 361.050 451.050 ;
        RECT 362.100 448.200 366.900 449.400 ;
        RECT 352.950 445.950 355.050 448.050 ;
        RECT 365.100 447.600 366.900 448.200 ;
        RECT 322.950 442.950 325.050 445.050 ;
        RECT 328.950 442.950 331.050 445.050 ;
        RECT 338.550 442.950 339.900 445.050 ;
        RECT 340.950 442.950 343.050 445.050 ;
        RECT 344.100 442.950 344.850 444.750 ;
        RECT 352.050 444.000 352.950 444.900 ;
        RECT 368.100 444.150 369.900 445.950 ;
        RECT 351.150 443.400 352.950 444.000 ;
        RECT 362.100 443.400 363.900 444.000 ;
        RECT 368.100 443.400 369.000 444.150 ;
        RECT 253.800 432.600 255.600 435.600 ;
        RECT 263.400 440.400 270.900 441.300 ;
        RECT 263.400 432.600 265.200 440.400 ;
        RECT 269.100 439.500 270.900 440.400 ;
        RECT 271.950 438.600 272.850 441.900 ;
        RECT 270.900 436.800 272.850 438.600 ;
        RECT 287.400 438.600 288.300 441.900 ;
        RECT 311.100 441.000 315.300 442.650 ;
        RECT 329.850 441.750 331.050 441.900 ;
        RECT 287.400 436.950 292.800 438.600 ;
        RECT 270.900 432.600 272.700 436.800 ;
        RECT 291.000 432.600 292.800 436.950 ;
        RECT 311.100 432.600 312.900 441.000 ;
        RECT 329.850 440.700 333.600 441.750 ;
        RECT 323.400 437.700 331.200 439.050 ;
        RECT 323.400 432.600 325.200 437.700 ;
        RECT 329.400 432.600 331.200 437.700 ;
        RECT 332.400 438.600 333.600 440.700 ;
        RECT 338.550 438.600 339.750 442.950 ;
        RECT 351.150 442.200 369.000 443.400 ;
        RECT 362.100 439.200 363.150 442.200 ;
        RECT 332.400 432.600 334.200 438.600 ;
        RECT 338.550 432.600 340.350 438.600 ;
        RECT 343.950 437.700 346.050 438.600 ;
        RECT 358.350 438.450 360.150 439.200 ;
        RECT 343.950 436.500 347.700 437.700 ;
        RECT 346.650 435.600 347.700 436.500 ;
        RECT 355.200 437.400 360.150 438.450 ;
        RECT 361.650 437.400 363.450 439.200 ;
        RECT 370.950 438.600 371.850 453.300 ;
        RECT 381.150 452.700 383.100 453.600 ;
        RECT 377.100 449.100 378.900 449.850 ;
        RECT 376.950 445.950 379.050 448.050 ;
        RECT 381.150 446.100 382.050 452.700 ;
        RECT 384.000 446.100 385.200 455.400 ;
        RECT 390.150 454.500 391.050 455.400 ;
        RECT 406.950 454.800 407.850 456.900 ;
        RECT 411.450 456.600 413.250 456.900 ;
        RECT 414.150 456.600 416.850 458.400 ;
        RECT 414.150 455.700 415.050 456.600 ;
        RECT 399.450 454.500 407.850 454.800 ;
        RECT 390.150 453.900 407.850 454.500 ;
        RECT 409.050 454.800 415.050 455.700 ;
        RECT 415.950 454.800 418.050 455.700 ;
        RECT 421.650 455.400 423.450 467.400 ;
        RECT 390.150 453.300 401.250 453.900 ;
        RECT 381.150 441.900 381.900 446.100 ;
        RECT 382.950 442.950 385.050 445.050 ;
        RECT 381.150 441.300 382.050 441.900 ;
        RECT 381.150 440.400 383.100 441.300 ;
        RECT 355.200 435.600 356.250 437.400 ;
        RECT 364.950 436.500 367.050 438.600 ;
        RECT 364.950 435.600 366.000 436.500 ;
        RECT 346.650 432.600 348.450 435.600 ;
        RECT 354.450 432.600 356.250 435.600 ;
        RECT 362.250 434.700 366.000 435.600 ;
        RECT 362.250 432.600 364.050 434.700 ;
        RECT 370.050 432.600 371.850 438.600 ;
        RECT 378.000 439.500 383.100 440.400 ;
        RECT 378.000 435.600 379.200 439.500 ;
        RECT 384.000 438.600 385.200 441.900 ;
        RECT 390.150 438.600 391.050 453.300 ;
        RECT 399.450 453.000 401.250 453.300 ;
        RECT 395.100 448.200 399.900 449.400 ;
        RECT 400.950 448.950 403.050 451.050 ;
        RECT 409.050 449.100 409.950 454.800 ;
        RECT 415.950 453.600 420.150 454.800 ;
        RECT 419.250 451.800 421.050 453.600 ;
        RECT 395.100 447.600 396.900 448.200 ;
        RECT 406.950 445.950 412.050 448.050 ;
        RECT 392.100 444.150 393.900 445.950 ;
        RECT 422.250 445.050 423.450 455.400 ;
        RECT 431.400 461.400 433.200 467.400 ;
        RECT 431.400 454.500 432.600 461.400 ;
        RECT 437.700 455.400 439.500 467.400 ;
        RECT 444.150 455.400 445.950 467.400 ;
        RECT 452.550 461.400 454.350 467.400 ;
        RECT 452.550 460.500 453.750 461.400 ;
        RECT 460.350 460.500 462.150 467.400 ;
        RECT 468.150 461.400 469.950 467.400 ;
        RECT 448.950 458.400 453.750 460.500 ;
        RECT 456.450 459.450 463.050 460.500 ;
        RECT 456.450 458.700 458.250 459.450 ;
        RECT 461.250 458.700 463.050 459.450 ;
        RECT 468.150 459.300 472.050 461.400 ;
        RECT 452.550 457.500 453.750 458.400 ;
        RECT 465.450 457.800 467.250 458.400 ;
        RECT 452.550 456.300 460.050 457.500 ;
        RECT 458.250 455.700 460.050 456.300 ;
        RECT 460.950 456.900 467.250 457.800 ;
        RECT 431.400 453.600 437.100 454.500 ;
        RECT 435.150 452.700 437.100 453.600 ;
        RECT 431.100 449.100 432.900 449.850 ;
        RECT 430.950 445.950 433.050 448.050 ;
        RECT 435.150 446.100 436.050 452.700 ;
        RECT 438.000 446.100 439.200 455.400 ;
        RECT 444.150 454.500 445.050 455.400 ;
        RECT 460.950 454.800 461.850 456.900 ;
        RECT 465.450 456.600 467.250 456.900 ;
        RECT 468.150 456.600 470.850 458.400 ;
        RECT 468.150 455.700 469.050 456.600 ;
        RECT 453.450 454.500 461.850 454.800 ;
        RECT 444.150 453.900 461.850 454.500 ;
        RECT 463.050 454.800 469.050 455.700 ;
        RECT 469.950 454.800 472.050 455.700 ;
        RECT 475.650 455.400 477.450 467.400 ;
        RECT 490.800 461.400 492.600 467.400 ;
        RECT 444.150 453.300 455.250 453.900 ;
        RECT 393.000 443.400 393.900 444.150 ;
        RECT 409.050 444.000 409.950 444.900 ;
        RECT 398.100 443.400 399.900 444.000 ;
        RECT 409.050 443.400 410.850 444.000 ;
        RECT 393.000 442.200 410.850 443.400 ;
        RECT 417.150 442.950 417.900 444.750 ;
        RECT 418.950 442.950 421.050 445.050 ;
        RECT 422.100 442.950 423.450 445.050 ;
        RECT 398.850 439.200 399.900 442.200 ;
        RECT 377.400 432.600 379.200 435.600 ;
        RECT 383.700 432.600 385.500 438.600 ;
        RECT 390.150 432.600 391.950 438.600 ;
        RECT 394.950 436.500 397.050 438.600 ;
        RECT 398.550 437.400 400.350 439.200 ;
        RECT 401.850 438.450 403.650 439.200 ;
        RECT 422.250 438.600 423.450 442.950 ;
        RECT 435.150 441.900 435.900 446.100 ;
        RECT 436.950 442.950 439.050 445.050 ;
        RECT 435.150 441.300 436.050 441.900 ;
        RECT 435.150 440.400 437.100 441.300 ;
        RECT 401.850 437.400 406.800 438.450 ;
        RECT 415.950 437.700 418.050 438.600 ;
        RECT 396.000 435.600 397.050 436.500 ;
        RECT 405.750 435.600 406.800 437.400 ;
        RECT 414.300 436.500 418.050 437.700 ;
        RECT 414.300 435.600 415.350 436.500 ;
        RECT 396.000 434.700 399.750 435.600 ;
        RECT 397.950 432.600 399.750 434.700 ;
        RECT 405.750 432.600 407.550 435.600 ;
        RECT 413.550 432.600 415.350 435.600 ;
        RECT 421.650 432.600 423.450 438.600 ;
        RECT 432.000 439.500 437.100 440.400 ;
        RECT 432.000 435.600 433.200 439.500 ;
        RECT 438.000 438.600 439.200 441.900 ;
        RECT 444.150 438.600 445.050 453.300 ;
        RECT 453.450 453.000 455.250 453.300 ;
        RECT 449.100 448.200 453.900 449.400 ;
        RECT 449.100 447.600 450.900 448.200 ;
        RECT 454.950 445.950 457.050 451.050 ;
        RECT 463.050 449.100 463.950 454.800 ;
        RECT 469.950 453.600 474.150 454.800 ;
        RECT 473.250 451.800 475.050 453.600 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 446.100 444.150 447.900 445.950 ;
        RECT 476.250 445.050 477.450 455.400 ;
        RECT 487.950 451.950 490.050 454.050 ;
        RECT 488.100 450.150 489.900 450.900 ;
        RECT 491.400 449.100 492.600 461.400 ;
        RECT 508.500 455.400 510.300 467.400 ;
        RECT 524.400 455.400 526.200 467.400 ;
        RECT 531.150 455.400 532.950 467.400 ;
        RECT 539.550 461.400 541.350 467.400 ;
        RECT 539.550 460.500 540.750 461.400 ;
        RECT 547.350 460.500 549.150 467.400 ;
        RECT 555.150 461.400 556.950 467.400 ;
        RECT 535.950 458.400 540.750 460.500 ;
        RECT 543.450 459.450 550.050 460.500 ;
        RECT 543.450 458.700 545.250 459.450 ;
        RECT 548.250 458.700 550.050 459.450 ;
        RECT 555.150 459.300 559.050 461.400 ;
        RECT 539.550 457.500 540.750 458.400 ;
        RECT 552.450 457.800 554.250 458.400 ;
        RECT 539.550 456.300 547.050 457.500 ;
        RECT 545.250 455.700 547.050 456.300 ;
        RECT 547.950 456.900 554.250 457.800 ;
        RECT 493.950 451.950 496.050 454.050 ;
        RECT 508.950 452.100 510.150 455.400 ;
        RECT 494.100 450.150 495.900 450.900 ;
        RECT 505.950 448.950 508.050 451.050 ;
        RECT 484.950 447.450 489.000 448.050 ;
        RECT 490.950 447.450 493.050 448.050 ;
        RECT 509.100 447.900 510.150 452.100 ;
        RECT 511.950 448.950 514.050 451.050 ;
        RECT 520.950 448.950 523.050 451.050 ;
        RECT 484.950 446.550 493.050 447.450 ;
        RECT 506.100 447.150 507.900 447.900 ;
        RECT 484.950 445.950 489.000 446.550 ;
        RECT 490.950 445.950 493.050 446.550 ;
        RECT 503.100 446.100 504.900 446.850 ;
        RECT 508.950 446.100 510.150 447.900 ;
        RECT 512.100 447.150 513.900 447.900 ;
        RECT 521.100 447.150 522.900 447.900 ;
        RECT 524.400 446.100 525.600 455.400 ;
        RECT 531.150 454.500 532.050 455.400 ;
        RECT 547.950 454.800 548.850 456.900 ;
        RECT 552.450 456.600 554.250 456.900 ;
        RECT 555.150 456.600 557.850 458.400 ;
        RECT 555.150 455.700 556.050 456.600 ;
        RECT 540.450 454.500 548.850 454.800 ;
        RECT 531.150 453.900 548.850 454.500 ;
        RECT 550.050 454.800 556.050 455.700 ;
        RECT 556.950 454.800 559.050 455.700 ;
        RECT 562.650 455.400 564.450 467.400 ;
        RECT 577.500 455.400 579.300 467.400 ;
        RECT 531.150 453.300 542.250 453.900 ;
        RECT 447.000 443.400 447.900 444.150 ;
        RECT 463.050 444.000 463.950 444.900 ;
        RECT 452.100 443.400 453.900 444.000 ;
        RECT 463.050 443.400 464.850 444.000 ;
        RECT 447.000 442.200 464.850 443.400 ;
        RECT 471.150 442.950 471.900 444.750 ;
        RECT 472.950 442.950 475.050 445.050 ;
        RECT 476.100 442.950 477.450 445.050 ;
        RECT 452.850 439.200 453.900 442.200 ;
        RECT 431.400 432.600 433.200 435.600 ;
        RECT 437.700 432.600 439.500 438.600 ;
        RECT 444.150 432.600 445.950 438.600 ;
        RECT 448.950 436.500 451.050 438.600 ;
        RECT 452.550 437.400 454.350 439.200 ;
        RECT 455.850 438.450 457.650 439.200 ;
        RECT 476.250 438.600 477.450 442.950 ;
        RECT 491.400 440.700 492.600 444.900 ;
        RECT 502.950 442.950 505.050 445.050 ;
        RECT 508.950 442.950 511.050 445.050 ;
        RECT 523.950 442.950 526.050 445.050 ;
        RECT 509.850 441.750 511.050 441.900 ;
        RECT 509.850 440.700 513.600 441.750 ;
        RECT 455.850 437.400 460.800 438.450 ;
        RECT 469.950 437.700 472.050 438.600 ;
        RECT 450.000 435.600 451.050 436.500 ;
        RECT 459.750 435.600 460.800 437.400 ;
        RECT 468.300 436.500 472.050 437.700 ;
        RECT 468.300 435.600 469.350 436.500 ;
        RECT 450.000 434.700 453.750 435.600 ;
        RECT 451.950 432.600 453.750 434.700 ;
        RECT 459.750 432.600 461.550 435.600 ;
        RECT 467.550 432.600 469.350 435.600 ;
        RECT 475.650 432.600 477.450 438.600 ;
        RECT 489.000 439.800 492.600 440.700 ;
        RECT 489.000 432.600 490.800 439.800 ;
        RECT 503.400 437.700 511.200 439.050 ;
        RECT 503.400 432.600 505.200 437.700 ;
        RECT 509.400 432.600 511.200 437.700 ;
        RECT 512.400 438.600 513.600 440.700 ;
        RECT 524.400 438.600 525.600 441.900 ;
        RECT 531.150 438.600 532.050 453.300 ;
        RECT 540.450 453.000 542.250 453.300 ;
        RECT 536.100 448.200 540.900 449.400 ;
        RECT 541.950 448.950 544.050 451.050 ;
        RECT 550.050 449.100 550.950 454.800 ;
        RECT 556.950 453.600 561.150 454.800 ;
        RECT 560.250 451.800 562.050 453.600 ;
        RECT 536.100 447.600 537.900 448.200 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 533.100 444.150 534.900 445.950 ;
        RECT 563.250 445.050 564.450 455.400 ;
        RECT 577.950 452.100 579.150 455.400 ;
        RECT 596.400 454.500 598.200 467.400 ;
        RECT 602.400 454.500 604.200 467.400 ;
        RECT 608.400 454.500 610.200 467.400 ;
        RECT 614.400 454.500 616.200 467.400 ;
        RECT 635.700 455.400 637.500 467.400 ;
        RECT 652.800 461.400 654.600 467.400 ;
        RECT 596.400 453.300 600.300 454.500 ;
        RECT 602.400 453.300 606.300 454.500 ;
        RECT 608.400 453.300 612.300 454.500 ;
        RECT 614.400 453.300 617.100 454.500 ;
        RECT 574.950 448.950 577.050 451.050 ;
        RECT 578.100 447.900 579.150 452.100 ;
        RECT 580.950 448.950 583.050 451.050 ;
        RECT 575.100 447.150 576.900 447.900 ;
        RECT 572.100 446.100 573.900 446.850 ;
        RECT 577.950 446.100 579.150 447.900 ;
        RECT 581.100 447.150 582.900 447.900 ;
        RECT 534.000 443.400 534.900 444.150 ;
        RECT 550.050 444.000 550.950 444.900 ;
        RECT 539.100 443.400 540.900 444.000 ;
        RECT 550.050 443.400 551.850 444.000 ;
        RECT 534.000 442.200 551.850 443.400 ;
        RECT 558.150 442.950 558.900 444.750 ;
        RECT 559.950 442.950 562.050 445.050 ;
        RECT 563.100 442.950 564.450 445.050 ;
        RECT 571.950 442.950 574.050 445.050 ;
        RECT 577.950 442.950 580.050 445.050 ;
        RECT 596.100 444.150 597.900 444.900 ;
        RECT 539.850 439.200 540.900 442.200 ;
        RECT 512.400 432.600 514.200 438.600 ;
        RECT 524.400 432.600 526.200 438.600 ;
        RECT 531.150 432.600 532.950 438.600 ;
        RECT 535.950 436.500 538.050 438.600 ;
        RECT 539.550 437.400 541.350 439.200 ;
        RECT 542.850 438.450 544.650 439.200 ;
        RECT 563.250 438.600 564.450 442.950 ;
        RECT 599.100 442.800 600.300 453.300 ;
        RECT 601.500 442.800 603.300 443.400 ;
        RECT 578.850 441.750 580.050 441.900 ;
        RECT 578.850 440.700 582.600 441.750 ;
        RECT 599.100 441.600 603.300 442.800 ;
        RECT 605.100 442.800 606.300 453.300 ;
        RECT 607.500 442.800 609.300 443.400 ;
        RECT 605.100 441.600 609.300 442.800 ;
        RECT 611.100 442.800 612.300 453.300 ;
        RECT 616.200 449.100 617.100 453.300 ;
        RECT 635.850 452.100 637.050 455.400 ;
        RECT 653.400 452.100 654.600 461.400 ;
        RECT 665.400 461.400 667.200 467.400 ;
        RECT 683.400 461.400 685.200 467.400 ;
        RECT 631.950 448.950 634.050 451.050 ;
        RECT 613.950 445.950 619.050 448.050 ;
        RECT 635.850 447.900 636.900 452.100 ;
        RECT 661.950 451.950 664.050 454.050 ;
        RECT 637.950 448.950 640.050 451.050 ;
        RECT 649.950 448.950 655.050 451.050 ;
        RECT 662.100 450.150 663.900 450.900 ;
        RECT 665.400 449.100 666.600 461.400 ;
        RECT 667.950 451.950 670.050 454.050 ;
        RECT 679.950 451.950 682.050 454.050 ;
        RECT 668.100 450.150 669.900 450.900 ;
        RECT 680.100 450.150 681.900 450.900 ;
        RECT 683.400 449.100 684.600 461.400 ;
        RECT 695.400 455.400 697.200 467.400 ;
        RECT 702.900 456.900 704.700 467.400 ;
        RECT 719.400 461.400 721.200 467.400 ;
        RECT 702.900 455.400 705.300 456.900 ;
        RECT 695.400 454.200 696.600 455.400 ;
        RECT 685.950 451.950 688.050 454.050 ;
        RECT 695.400 453.000 702.600 454.200 ;
        RECT 700.800 452.400 702.600 453.000 ;
        RECT 686.100 450.150 687.900 450.900 ;
        RECT 694.950 448.950 697.050 451.050 ;
        RECT 662.550 447.900 667.050 448.050 ;
        RECT 632.100 447.150 633.900 447.900 ;
        RECT 635.850 446.100 637.050 447.900 ;
        RECT 638.100 447.150 639.900 447.900 ;
        RECT 641.100 446.100 642.900 446.850 ;
        RECT 613.500 442.800 615.300 443.400 ;
        RECT 611.100 441.600 615.300 442.800 ;
        RECT 599.100 440.700 600.300 441.600 ;
        RECT 605.100 440.700 606.300 441.600 ;
        RECT 611.100 440.700 612.300 441.600 ;
        RECT 616.200 440.700 617.100 444.900 ;
        RECT 634.950 442.950 637.050 445.050 ;
        RECT 640.950 442.950 643.050 445.050 ;
        RECT 634.950 441.750 636.150 441.900 ;
        RECT 542.850 437.400 547.800 438.450 ;
        RECT 556.950 437.700 559.050 438.600 ;
        RECT 537.000 435.600 538.050 436.500 ;
        RECT 546.750 435.600 547.800 437.400 ;
        RECT 555.300 436.500 559.050 437.700 ;
        RECT 555.300 435.600 556.350 436.500 ;
        RECT 537.000 434.700 540.750 435.600 ;
        RECT 538.950 432.600 540.750 434.700 ;
        RECT 546.750 432.600 548.550 435.600 ;
        RECT 554.550 432.600 556.350 435.600 ;
        RECT 562.650 432.600 564.450 438.600 ;
        RECT 572.400 437.700 580.200 439.050 ;
        RECT 572.400 432.600 574.200 437.700 ;
        RECT 578.400 432.600 580.200 437.700 ;
        RECT 581.400 438.600 582.600 440.700 ;
        RECT 596.400 439.500 600.300 440.700 ;
        RECT 602.400 439.500 606.300 440.700 ;
        RECT 608.400 439.500 612.300 440.700 ;
        RECT 614.400 439.500 617.100 440.700 ;
        RECT 632.400 440.700 636.150 441.750 ;
        RECT 581.400 432.600 583.200 438.600 ;
        RECT 596.400 432.600 598.200 439.500 ;
        RECT 602.400 432.600 604.200 439.500 ;
        RECT 608.400 432.600 610.200 439.500 ;
        RECT 614.400 432.600 616.200 439.500 ;
        RECT 632.400 438.600 633.600 440.700 ;
        RECT 631.800 432.600 633.600 438.600 ;
        RECT 634.800 437.700 642.600 439.050 ;
        RECT 634.800 432.600 636.600 437.700 ;
        RECT 640.800 432.600 642.600 437.700 ;
        RECT 653.400 435.600 654.600 447.900 ;
        RECT 656.100 446.100 657.900 446.850 ;
        RECT 661.950 445.950 667.050 447.900 ;
        RECT 682.950 447.450 685.050 448.050 ;
        RECT 687.000 447.450 691.050 448.050 ;
        RECT 682.950 446.550 691.050 447.450 ;
        RECT 695.100 447.150 696.900 447.900 ;
        RECT 682.950 445.950 685.050 446.550 ;
        RECT 687.000 445.950 691.050 446.550 ;
        RECT 698.100 446.100 699.900 446.850 ;
        RECT 661.950 445.800 664.050 445.950 ;
        RECT 655.950 442.950 658.050 445.050 ;
        RECT 665.400 440.700 666.600 444.900 ;
        RECT 683.400 440.700 684.600 444.900 ;
        RECT 697.950 442.950 700.050 445.050 ;
        RECT 701.700 441.600 702.600 452.400 ;
        RECT 703.950 449.100 705.300 455.400 ;
        RECT 719.400 452.100 720.600 461.400 ;
        RECT 735.600 455.400 737.400 467.400 ;
        RECT 734.700 454.350 737.400 455.400 ;
        RECT 750.600 455.400 752.400 467.400 ;
        RECT 761.400 456.300 763.200 467.400 ;
        RECT 767.400 456.300 769.200 467.400 ;
        RECT 761.400 455.400 769.200 456.300 ;
        RECT 770.400 455.400 772.200 467.400 ;
        RECT 785.400 461.400 787.200 467.400 ;
        RECT 800.400 461.400 802.200 467.400 ;
        RECT 750.600 454.350 753.300 455.400 ;
        RECT 731.100 452.100 732.900 452.850 ;
        RECT 718.950 450.450 721.050 451.050 ;
        RECT 723.000 450.450 727.050 451.050 ;
        RECT 718.950 449.550 727.050 450.450 ;
        RECT 718.950 448.950 721.050 449.550 ;
        RECT 723.000 448.950 727.050 449.550 ;
        RECT 730.950 448.950 733.050 451.050 ;
        RECT 734.700 449.100 736.050 454.350 ;
        RECT 737.100 449.100 738.900 449.850 ;
        RECT 749.100 449.100 750.900 449.850 ;
        RECT 751.950 449.100 753.300 454.350 ;
        RECT 755.100 452.100 756.900 452.850 ;
        RECT 703.950 447.450 706.050 448.050 ;
        RECT 708.000 447.450 712.050 448.050 ;
        RECT 703.950 446.550 712.050 447.450 ;
        RECT 703.950 445.950 706.050 446.550 ;
        RECT 708.000 445.950 712.050 446.550 ;
        RECT 716.100 446.100 717.900 446.850 ;
        RECT 700.950 440.700 702.750 441.600 ;
        RECT 665.400 439.800 669.000 440.700 ;
        RECT 683.400 439.800 687.000 440.700 ;
        RECT 652.800 432.600 654.600 435.600 ;
        RECT 667.200 432.600 669.000 439.800 ;
        RECT 685.200 432.600 687.000 439.800 ;
        RECT 699.300 439.800 702.750 440.700 ;
        RECT 699.300 435.600 700.200 439.800 ;
        RECT 705.000 438.600 706.050 444.900 ;
        RECT 715.950 442.950 718.050 445.050 ;
        RECT 698.400 432.600 700.200 435.600 ;
        RECT 704.400 432.600 706.200 438.600 ;
        RECT 719.400 435.600 720.600 447.900 ;
        RECT 734.700 444.900 735.900 449.100 ;
        RECT 736.950 445.950 739.050 448.050 ;
        RECT 748.950 445.950 751.050 448.050 ;
        RECT 752.100 444.900 753.300 449.100 ;
        RECT 754.950 448.950 757.050 451.050 ;
        RECT 760.950 448.950 763.050 451.050 ;
        RECT 766.950 448.950 769.050 451.050 ;
        RECT 761.100 447.150 762.900 447.900 ;
        RECT 767.100 447.150 768.900 447.900 ;
        RECT 764.100 446.100 765.900 446.850 ;
        RECT 770.700 446.100 771.600 455.400 ;
        RECT 785.400 452.100 786.600 461.400 ;
        RECT 800.700 461.100 802.200 461.400 ;
        RECT 806.400 461.400 808.200 467.400 ;
        RECT 818.400 461.400 820.200 467.400 ;
        RECT 806.400 461.100 807.300 461.400 ;
        RECT 800.700 460.200 807.300 461.100 ;
        RECT 796.950 454.950 799.050 457.050 ;
        RECT 806.400 455.100 807.300 460.200 ;
        RECT 818.400 454.500 819.600 461.400 ;
        RECT 824.700 455.400 826.500 467.400 ;
        RECT 797.100 453.150 798.900 453.900 ;
        RECT 800.100 452.100 801.900 452.850 ;
        RECT 805.950 451.950 808.050 454.050 ;
        RECT 818.400 453.600 824.100 454.500 ;
        RECT 822.150 452.700 824.100 453.600 ;
        RECT 772.950 450.450 775.050 451.050 ;
        RECT 784.950 450.450 787.050 451.050 ;
        RECT 772.950 449.550 787.050 450.450 ;
        RECT 772.950 448.950 775.050 449.550 ;
        RECT 784.950 448.950 787.050 449.550 ;
        RECT 799.950 448.950 802.050 451.050 ;
        RECT 782.100 446.100 783.900 446.850 ;
        RECT 734.700 443.100 736.050 444.900 ;
        RECT 751.950 443.100 753.300 444.900 ;
        RECT 757.950 444.450 762.000 445.050 ;
        RECT 763.950 444.450 766.050 445.050 ;
        RECT 757.950 443.550 766.050 444.450 ;
        RECT 757.950 442.950 762.000 443.550 ;
        RECT 763.950 442.950 766.050 443.550 ;
        RECT 769.950 442.950 772.050 445.050 ;
        RECT 781.950 442.950 784.050 445.050 ;
        RECT 730.950 439.950 736.050 442.050 ;
        RECT 742.950 441.450 745.050 442.050 ;
        RECT 751.950 441.450 754.050 442.050 ;
        RECT 742.950 440.550 754.050 441.450 ;
        RECT 742.950 439.950 745.050 440.550 ;
        RECT 751.950 439.950 754.050 440.550 ;
        RECT 734.400 435.600 735.600 438.900 ;
        RECT 752.400 435.600 753.600 438.900 ;
        RECT 770.700 438.600 771.600 441.900 ;
        RECT 719.400 432.600 721.200 435.600 ;
        RECT 734.400 432.600 736.200 435.600 ;
        RECT 751.800 432.600 753.600 435.600 ;
        RECT 766.200 436.950 771.600 438.600 ;
        RECT 766.200 432.600 768.000 436.950 ;
        RECT 785.400 435.600 786.600 447.900 ;
        RECT 802.950 445.950 805.050 448.050 ;
        RECT 803.100 444.150 804.900 444.900 ;
        RECT 806.400 442.650 807.300 450.900 ;
        RECT 818.100 449.100 819.900 449.850 ;
        RECT 817.950 442.950 820.050 448.050 ;
        RECT 822.150 446.100 823.050 452.700 ;
        RECT 825.000 446.100 826.200 455.400 ;
        RECT 803.100 441.000 807.300 442.650 ;
        RECT 822.150 441.900 822.900 446.100 ;
        RECT 822.150 441.300 823.050 441.900 ;
        RECT 785.400 432.600 787.200 435.600 ;
        RECT 803.100 432.600 804.900 441.000 ;
        RECT 822.150 440.400 824.100 441.300 ;
        RECT 819.000 439.500 824.100 440.400 ;
        RECT 819.000 435.600 820.200 439.500 ;
        RECT 825.000 438.600 826.200 441.900 ;
        RECT 818.400 432.600 820.200 435.600 ;
        RECT 824.700 432.600 826.500 438.600 ;
        RECT 10.800 425.400 12.600 428.400 ;
        RECT 11.400 413.100 12.600 425.400 ;
        RECT 27.000 424.050 28.800 428.400 ;
        RECT 23.400 422.400 28.800 424.050 ;
        RECT 23.400 419.100 24.300 422.400 ;
        RECT 44.100 420.000 45.900 428.400 ;
        RECT 41.700 418.350 45.900 420.000 ;
        RECT 69.000 422.400 70.800 428.400 ;
        RECT 69.000 419.100 70.050 422.400 ;
        RECT 85.200 421.200 87.000 428.400 ;
        RECT 83.400 420.300 87.000 421.200 ;
        RECT 13.950 415.950 16.050 418.050 ;
        RECT 19.950 415.950 25.050 418.050 ;
        RECT 28.950 415.950 31.050 418.050 ;
        RECT 14.100 414.150 15.900 414.900 ;
        RECT 10.950 411.450 13.050 412.050 ;
        RECT 15.000 411.450 19.050 412.050 ;
        RECT 10.950 410.550 19.050 411.450 ;
        RECT 10.950 409.950 13.050 410.550 ;
        RECT 15.000 409.950 19.050 410.550 ;
        RECT 11.400 399.600 12.600 408.900 ;
        RECT 23.400 405.600 24.300 414.900 ;
        RECT 29.100 414.150 30.900 414.900 ;
        RECT 26.100 413.100 27.900 413.850 ;
        RECT 32.100 413.100 33.900 413.850 ;
        RECT 25.950 409.950 28.050 412.050 ;
        RECT 31.950 409.950 34.050 412.050 ;
        RECT 41.700 410.100 42.600 418.350 ;
        RECT 44.100 416.100 45.900 416.850 ;
        RECT 58.950 415.950 64.050 418.050 ;
        RECT 67.950 415.950 70.050 418.050 ;
        RECT 73.950 415.950 79.050 418.050 ;
        RECT 83.400 416.100 84.600 420.300 ;
        RECT 101.100 420.000 102.900 428.400 ;
        RECT 120.000 424.050 121.800 428.400 ;
        RECT 136.800 425.400 138.600 428.400 ;
        RECT 98.700 418.350 102.900 420.000 ;
        RECT 116.400 422.400 121.800 424.050 ;
        RECT 116.400 419.100 117.300 422.400 ;
        RECT 61.950 415.800 64.050 415.950 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 62.100 414.150 63.900 414.900 ;
        RECT 65.250 413.100 67.050 413.850 ;
        RECT 67.950 413.100 68.850 414.900 ;
        RECT 73.950 414.150 75.750 414.900 ;
        RECT 70.950 413.100 72.750 413.850 ;
        RECT 46.950 409.950 49.050 412.050 ;
        RECT 64.950 409.950 67.050 412.050 ;
        RECT 40.950 406.950 43.050 409.050 ;
        RECT 68.100 408.900 68.850 413.100 ;
        RECT 82.950 412.950 85.050 415.050 ;
        RECT 47.100 408.150 48.900 408.900 ;
        RECT 50.100 407.100 51.900 407.850 ;
        RECT 67.950 407.400 68.850 408.900 ;
        RECT 64.800 406.500 68.850 407.400 ;
        RECT 70.950 406.950 73.050 412.050 ;
        RECT 80.100 410.100 81.900 410.850 ;
        RECT 79.950 406.950 82.050 409.050 ;
        RECT 10.800 393.600 12.600 399.600 ;
        RECT 22.800 393.600 24.600 405.600 ;
        RECT 25.800 404.700 33.600 405.600 ;
        RECT 25.800 393.600 27.600 404.700 ;
        RECT 31.800 393.600 33.600 404.700 ;
        RECT 41.700 400.800 42.600 405.900 ;
        RECT 49.950 403.950 52.050 406.050 ;
        RECT 41.700 399.900 48.300 400.800 ;
        RECT 41.700 399.600 42.600 399.900 ;
        RECT 40.800 393.600 42.600 399.600 ;
        RECT 46.800 399.600 48.300 399.900 ;
        RECT 46.800 393.600 48.600 399.600 ;
        RECT 61.800 394.500 63.600 405.600 ;
        RECT 64.800 395.400 66.600 406.500 ;
        RECT 67.800 404.400 75.600 405.300 ;
        RECT 67.800 394.500 69.600 404.400 ;
        RECT 61.800 393.600 69.600 394.500 ;
        RECT 73.800 393.600 75.600 404.400 ;
        RECT 83.400 399.600 84.600 411.900 ;
        RECT 86.100 410.100 87.900 410.850 ;
        RECT 98.700 410.100 99.600 418.350 ;
        RECT 109.950 417.450 114.000 418.050 ;
        RECT 115.950 417.450 118.050 418.050 ;
        RECT 101.100 416.100 102.900 416.850 ;
        RECT 109.950 416.550 118.050 417.450 ;
        RECT 109.950 415.950 114.000 416.550 ;
        RECT 115.950 415.950 118.050 416.550 ;
        RECT 121.950 415.950 124.050 418.050 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 103.950 409.950 106.050 412.050 ;
        RECT 85.950 406.950 88.050 409.050 ;
        RECT 94.950 406.950 100.050 409.050 ;
        RECT 104.100 408.150 105.900 408.900 ;
        RECT 107.100 407.100 108.900 407.850 ;
        RECT 98.700 400.800 99.600 405.900 ;
        RECT 106.950 403.950 109.050 406.050 ;
        RECT 116.400 405.600 117.300 414.900 ;
        RECT 122.100 414.150 123.900 414.900 ;
        RECT 119.100 413.100 120.900 413.850 ;
        RECT 125.100 413.100 126.900 413.850 ;
        RECT 118.950 409.950 121.050 412.050 ;
        RECT 124.950 409.950 127.050 412.050 ;
        RECT 130.950 411.450 133.050 415.050 ;
        RECT 137.400 413.100 138.600 425.400 ;
        RECT 148.800 422.400 150.600 428.400 ;
        RECT 149.400 420.300 150.600 422.400 ;
        RECT 151.800 423.300 153.600 428.400 ;
        RECT 157.800 423.300 159.600 428.400 ;
        RECT 169.800 425.400 171.600 428.400 ;
        RECT 151.800 421.950 159.600 423.300 ;
        RECT 170.400 422.100 171.600 425.400 ;
        RECT 184.200 421.200 186.000 428.400 ;
        RECT 199.800 422.400 201.600 428.400 ;
        RECT 149.400 419.250 153.150 420.300 ;
        RECT 151.950 419.100 153.150 419.250 ;
        RECT 169.950 418.950 172.050 421.050 ;
        RECT 182.400 420.300 186.000 421.200 ;
        RECT 200.400 420.300 201.600 422.400 ;
        RECT 202.800 423.300 204.600 428.400 ;
        RECT 208.800 423.300 210.600 428.400 ;
        RECT 202.800 421.950 210.600 423.300 ;
        RECT 221.400 425.400 223.200 428.400 ;
        RECT 236.400 425.400 238.200 428.400 ;
        RECT 221.400 422.100 222.600 425.400 ;
        RECT 139.950 415.800 142.050 418.050 ;
        RECT 145.950 417.450 150.000 418.050 ;
        RECT 151.950 417.450 154.050 418.050 ;
        RECT 145.950 416.550 154.050 417.450 ;
        RECT 145.950 415.950 150.000 416.550 ;
        RECT 151.950 415.950 154.050 416.550 ;
        RECT 157.950 415.950 160.050 418.050 ;
        RECT 169.950 416.100 171.300 417.900 ;
        RECT 182.400 416.100 183.600 420.300 ;
        RECT 200.400 419.250 204.150 420.300 ;
        RECT 202.950 419.100 204.150 419.250 ;
        RECT 220.950 418.950 223.050 421.050 ;
        RECT 190.950 417.450 193.050 418.050 ;
        RECT 202.950 417.450 205.050 418.050 ;
        RECT 190.950 416.550 205.050 417.450 ;
        RECT 140.100 414.150 141.900 414.900 ;
        RECT 149.100 413.100 150.900 413.850 ;
        RECT 152.850 413.100 154.050 414.900 ;
        RECT 158.100 414.150 159.900 414.900 ;
        RECT 155.100 413.100 156.900 413.850 ;
        RECT 136.950 411.450 139.050 412.050 ;
        RECT 130.950 411.000 139.050 411.450 ;
        RECT 131.550 410.550 139.050 411.000 ;
        RECT 136.950 409.950 139.050 410.550 ;
        RECT 148.950 409.950 151.050 412.050 ;
        RECT 152.850 408.900 153.900 413.100 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 154.950 409.950 157.050 412.050 ;
        RECT 170.100 411.900 171.300 416.100 ;
        RECT 190.950 415.950 193.050 416.550 ;
        RECT 202.950 415.950 205.050 416.550 ;
        RECT 208.950 415.950 211.050 418.050 ;
        RECT 221.700 416.100 223.050 417.900 ;
        RECT 178.950 412.950 184.050 415.050 ;
        RECT 200.100 413.100 201.900 413.850 ;
        RECT 203.850 413.100 205.050 414.900 ;
        RECT 209.100 414.150 210.900 414.900 ;
        RECT 206.100 413.100 207.900 413.850 ;
        RECT 167.100 411.150 168.900 411.900 ;
        RECT 98.700 399.900 105.300 400.800 ;
        RECT 98.700 399.600 99.600 399.900 ;
        RECT 83.400 393.600 85.200 399.600 ;
        RECT 97.800 393.600 99.600 399.600 ;
        RECT 103.800 399.600 105.300 399.900 ;
        RECT 103.800 393.600 105.600 399.600 ;
        RECT 115.800 393.600 117.600 405.600 ;
        RECT 118.800 404.700 126.600 405.600 ;
        RECT 118.800 393.600 120.600 404.700 ;
        RECT 124.800 393.600 126.600 404.700 ;
        RECT 137.400 399.600 138.600 408.900 ;
        RECT 152.850 405.600 154.050 408.900 ;
        RECT 169.950 406.650 171.300 411.900 ;
        RECT 172.950 409.950 175.050 412.050 ;
        RECT 179.100 410.100 180.900 410.850 ;
        RECT 173.100 408.150 174.900 408.900 ;
        RECT 178.950 406.950 181.050 409.050 ;
        RECT 168.600 405.600 171.300 406.650 ;
        RECT 136.800 393.600 138.600 399.600 ;
        RECT 152.700 393.600 154.500 405.600 ;
        RECT 168.600 393.600 170.400 405.600 ;
        RECT 182.400 399.600 183.600 411.900 ;
        RECT 185.100 410.100 186.900 410.850 ;
        RECT 199.950 409.950 202.050 412.050 ;
        RECT 184.950 406.950 187.050 409.050 ;
        RECT 203.850 408.900 204.900 413.100 ;
        RECT 205.950 409.800 208.050 412.050 ;
        RECT 217.950 409.950 220.050 412.050 ;
        RECT 221.700 411.900 222.900 416.100 ;
        RECT 232.950 415.950 235.050 418.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 233.100 414.150 234.900 414.900 ;
        RECT 236.400 413.100 237.600 425.400 ;
        RECT 245.400 423.300 247.200 428.400 ;
        RECT 251.400 423.300 253.200 428.400 ;
        RECT 245.400 421.950 253.200 423.300 ;
        RECT 254.400 422.400 256.200 428.400 ;
        RECT 268.800 422.400 270.600 428.400 ;
        RECT 254.400 420.300 255.600 422.400 ;
        RECT 251.850 419.250 255.600 420.300 ;
        RECT 269.400 420.300 270.600 422.400 ;
        RECT 271.800 423.300 273.600 428.400 ;
        RECT 277.800 423.300 279.600 428.400 ;
        RECT 290.400 425.400 292.200 428.400 ;
        RECT 271.800 421.950 279.600 423.300 ;
        RECT 283.950 420.450 286.050 424.050 ;
        RECT 290.400 422.100 291.600 425.400 ;
        RECT 302.400 423.300 304.200 428.400 ;
        RECT 308.400 423.300 310.200 428.400 ;
        RECT 302.400 421.950 310.200 423.300 ;
        RECT 311.400 422.400 313.200 428.400 ;
        RECT 289.950 420.450 292.050 421.050 ;
        RECT 269.400 419.250 273.150 420.300 ;
        RECT 283.950 420.000 292.050 420.450 ;
        RECT 311.400 420.300 312.600 422.400 ;
        RECT 328.200 421.200 330.000 428.400 ;
        RECT 284.550 419.550 292.050 420.000 ;
        RECT 251.850 419.100 253.050 419.250 ;
        RECT 271.950 419.100 273.150 419.250 ;
        RECT 289.950 418.950 292.050 419.550 ;
        RECT 308.850 419.250 312.600 420.300 ;
        RECT 308.850 419.100 310.050 419.250 ;
        RECT 244.950 415.800 247.050 418.050 ;
        RECT 250.950 417.450 253.050 418.050 ;
        RECT 262.950 417.450 265.050 418.050 ;
        RECT 250.950 416.550 265.050 417.450 ;
        RECT 250.950 415.950 253.050 416.550 ;
        RECT 262.950 415.950 265.050 416.550 ;
        RECT 268.950 415.950 274.050 418.050 ;
        RECT 277.950 415.950 280.050 418.050 ;
        RECT 290.700 416.100 292.050 417.900 ;
        RECT 245.100 414.150 246.900 414.900 ;
        RECT 248.100 413.100 249.900 413.850 ;
        RECT 250.950 413.100 252.150 414.900 ;
        RECT 254.100 413.100 255.900 413.850 ;
        RECT 269.100 413.100 270.900 413.850 ;
        RECT 272.850 413.100 274.050 414.900 ;
        RECT 278.100 414.150 279.900 414.900 ;
        RECT 275.100 413.100 276.900 413.850 ;
        RECT 203.850 405.600 205.050 408.900 ;
        RECT 218.100 408.150 219.900 408.900 ;
        RECT 221.700 406.650 223.050 411.900 ;
        RECT 224.100 411.150 225.900 411.900 ;
        RECT 235.950 411.450 238.050 412.050 ;
        RECT 235.950 411.000 243.450 411.450 ;
        RECT 235.950 410.550 244.050 411.000 ;
        RECT 235.950 409.950 238.050 410.550 ;
        RECT 221.700 405.600 224.400 406.650 ;
        RECT 182.400 393.600 184.200 399.600 ;
        RECT 203.700 393.600 205.500 405.600 ;
        RECT 222.600 393.600 224.400 405.600 ;
        RECT 236.400 399.600 237.600 408.900 ;
        RECT 241.950 406.950 244.050 410.550 ;
        RECT 247.950 409.950 250.050 412.050 ;
        RECT 251.100 408.900 252.150 413.100 ;
        RECT 253.950 409.950 256.050 412.050 ;
        RECT 268.950 409.950 271.050 412.050 ;
        RECT 250.950 405.600 252.150 408.900 ;
        RECT 272.850 408.900 273.900 413.100 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 286.950 409.950 289.050 412.050 ;
        RECT 290.700 411.900 291.900 416.100 ;
        RECT 301.950 415.950 304.050 418.050 ;
        RECT 307.950 417.450 310.050 418.050 ;
        RECT 319.950 417.450 322.050 421.050 ;
        RECT 307.950 417.000 322.050 417.450 ;
        RECT 326.400 420.300 330.000 421.200 ;
        RECT 336.150 422.400 337.950 428.400 ;
        RECT 343.950 426.300 345.750 428.400 ;
        RECT 342.000 425.400 345.750 426.300 ;
        RECT 351.750 425.400 353.550 428.400 ;
        RECT 359.550 425.400 361.350 428.400 ;
        RECT 342.000 424.500 343.050 425.400 ;
        RECT 340.950 422.400 343.050 424.500 ;
        RECT 351.750 423.600 352.800 425.400 ;
        RECT 307.950 416.550 321.450 417.000 ;
        RECT 307.950 415.950 310.050 416.550 ;
        RECT 326.400 416.100 327.600 420.300 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 302.100 414.150 303.900 414.900 ;
        RECT 305.100 413.100 306.900 413.850 ;
        RECT 307.950 413.100 309.150 414.900 ;
        RECT 316.950 414.450 319.050 415.050 ;
        RECT 325.950 414.450 328.050 415.050 ;
        RECT 311.100 413.100 312.900 413.850 ;
        RECT 316.950 413.550 328.050 414.450 ;
        RECT 272.850 405.600 274.050 408.900 ;
        RECT 287.100 408.150 288.900 408.900 ;
        RECT 290.700 406.650 292.050 411.900 ;
        RECT 293.100 411.150 294.900 411.900 ;
        RECT 298.950 411.450 303.000 412.050 ;
        RECT 304.950 411.450 307.050 412.050 ;
        RECT 298.950 410.550 307.050 411.450 ;
        RECT 298.950 409.950 303.000 410.550 ;
        RECT 304.950 409.950 307.050 410.550 ;
        RECT 308.100 408.900 309.150 413.100 ;
        RECT 316.950 412.950 319.050 413.550 ;
        RECT 325.950 412.950 328.050 413.550 ;
        RECT 310.950 409.950 313.050 412.050 ;
        RECT 323.100 410.100 324.900 410.850 ;
        RECT 290.700 405.600 293.400 406.650 ;
        RECT 307.950 405.600 309.150 408.900 ;
        RECT 322.950 406.950 325.050 409.050 ;
        RECT 236.400 393.600 238.200 399.600 ;
        RECT 250.500 393.600 252.300 405.600 ;
        RECT 272.700 393.600 274.500 405.600 ;
        RECT 291.600 393.600 293.400 405.600 ;
        RECT 307.500 393.600 309.300 405.600 ;
        RECT 326.400 399.600 327.600 411.900 ;
        RECT 329.100 410.100 330.900 410.850 ;
        RECT 336.150 407.700 337.050 422.400 ;
        RECT 344.550 421.800 346.350 423.600 ;
        RECT 347.850 422.550 352.800 423.600 ;
        RECT 360.300 424.500 361.350 425.400 ;
        RECT 360.300 423.300 364.050 424.500 ;
        RECT 347.850 421.800 349.650 422.550 ;
        RECT 361.950 422.400 364.050 423.300 ;
        RECT 367.650 422.400 369.450 428.400 ;
        RECT 344.850 418.800 345.900 421.800 ;
        RECT 339.000 417.600 356.850 418.800 ;
        RECT 339.000 416.850 339.900 417.600 ;
        RECT 344.100 417.000 345.900 417.600 ;
        RECT 355.050 417.000 356.850 417.600 ;
        RECT 338.100 415.050 339.900 416.850 ;
        RECT 355.050 416.100 355.950 417.000 ;
        RECT 363.150 416.250 363.900 418.050 ;
        RECT 364.950 415.950 367.050 421.050 ;
        RECT 368.250 418.050 369.450 422.400 ;
        RECT 379.800 421.500 381.600 428.400 ;
        RECT 385.800 421.500 387.600 428.400 ;
        RECT 391.800 421.500 393.600 428.400 ;
        RECT 397.800 421.500 399.600 428.400 ;
        RECT 368.100 415.950 369.450 418.050 ;
        RECT 378.900 420.300 381.600 421.500 ;
        RECT 383.700 420.300 387.600 421.500 ;
        RECT 389.700 420.300 393.600 421.500 ;
        RECT 395.700 420.300 399.600 421.500 ;
        RECT 412.200 421.200 414.000 428.400 ;
        RECT 427.800 422.400 429.600 428.400 ;
        RECT 410.400 420.300 414.000 421.200 ;
        RECT 428.400 420.300 429.600 422.400 ;
        RECT 430.800 423.300 432.600 428.400 ;
        RECT 436.800 423.300 438.600 428.400 ;
        RECT 430.800 421.950 438.600 423.300 ;
        RECT 447.000 421.200 448.800 428.400 ;
        RECT 463.500 422.400 465.300 428.400 ;
        RECT 469.800 425.400 471.600 428.400 ;
        RECT 447.000 420.300 450.600 421.200 ;
        RECT 378.900 416.100 379.800 420.300 ;
        RECT 383.700 419.400 384.900 420.300 ;
        RECT 389.700 419.400 390.900 420.300 ;
        RECT 395.700 419.400 396.900 420.300 ;
        RECT 380.700 418.200 384.900 419.400 ;
        RECT 380.700 417.600 382.500 418.200 ;
        RECT 341.100 412.800 342.900 413.400 ;
        RECT 352.950 412.950 355.050 415.050 ;
        RECT 341.100 411.600 345.900 412.800 ;
        RECT 346.950 409.950 349.050 412.050 ;
        RECT 345.450 407.700 347.250 408.000 ;
        RECT 336.150 407.100 347.250 407.700 ;
        RECT 336.150 406.500 353.850 407.100 ;
        RECT 336.150 405.600 337.050 406.500 ;
        RECT 345.450 406.200 353.850 406.500 ;
        RECT 326.400 393.600 328.200 399.600 ;
        RECT 336.150 393.600 337.950 405.600 ;
        RECT 350.250 404.700 352.050 405.300 ;
        RECT 344.550 403.500 352.050 404.700 ;
        RECT 352.950 404.100 353.850 406.200 ;
        RECT 355.050 406.200 355.950 411.900 ;
        RECT 365.250 407.400 367.050 409.200 ;
        RECT 361.950 406.200 366.150 407.400 ;
        RECT 355.050 405.300 361.050 406.200 ;
        RECT 361.950 405.300 364.050 406.200 ;
        RECT 368.250 405.600 369.450 415.950 ;
        RECT 373.950 412.950 379.050 415.050 ;
        RECT 378.900 407.700 379.800 411.900 ;
        RECT 383.700 407.700 384.900 418.200 ;
        RECT 386.700 418.200 390.900 419.400 ;
        RECT 386.700 417.600 388.500 418.200 ;
        RECT 389.700 407.700 390.900 418.200 ;
        RECT 392.700 418.200 396.900 419.400 ;
        RECT 392.700 417.600 394.500 418.200 ;
        RECT 395.700 407.700 396.900 418.200 ;
        RECT 398.100 416.100 399.900 416.850 ;
        RECT 410.400 416.100 411.600 420.300 ;
        RECT 428.400 419.250 432.150 420.300 ;
        RECT 430.950 419.100 432.150 419.250 ;
        RECT 430.950 415.950 433.050 418.050 ;
        RECT 436.950 415.950 439.050 418.050 ;
        RECT 449.400 416.100 450.600 420.300 ;
        RECT 463.800 419.100 465.000 422.400 ;
        RECT 469.800 421.500 471.000 425.400 ;
        RECT 481.800 422.400 483.600 428.400 ;
        RECT 465.900 420.600 471.000 421.500 ;
        RECT 465.900 419.700 467.850 420.600 ;
        RECT 466.950 419.100 467.850 419.700 ;
        RECT 482.400 420.300 483.600 422.400 ;
        RECT 484.800 423.300 486.600 428.400 ;
        RECT 490.800 423.300 492.600 428.400 ;
        RECT 484.800 421.950 492.600 423.300 ;
        RECT 495.150 422.400 496.950 428.400 ;
        RECT 502.950 426.300 504.750 428.400 ;
        RECT 501.000 425.400 504.750 426.300 ;
        RECT 510.750 425.400 512.550 428.400 ;
        RECT 518.550 425.400 520.350 428.400 ;
        RECT 501.000 424.500 502.050 425.400 ;
        RECT 499.950 422.400 502.050 424.500 ;
        RECT 510.750 423.600 511.800 425.400 ;
        RECT 482.400 419.250 486.150 420.300 ;
        RECT 484.950 419.100 486.150 419.250 ;
        RECT 454.950 417.450 457.050 417.900 ;
        RECT 463.950 417.450 466.050 418.050 ;
        RECT 454.950 416.550 466.050 417.450 ;
        RECT 454.950 415.800 457.050 416.550 ;
        RECT 463.950 415.950 466.050 416.550 ;
        RECT 409.950 414.450 412.050 415.050 ;
        RECT 409.950 413.550 423.450 414.450 ;
        RECT 409.950 412.950 412.050 413.550 ;
        RECT 407.100 410.100 408.900 410.850 ;
        RECT 378.900 406.500 381.600 407.700 ;
        RECT 383.700 406.500 387.600 407.700 ;
        RECT 389.700 406.500 393.600 407.700 ;
        RECT 395.700 406.500 399.600 407.700 ;
        RECT 360.150 404.400 361.050 405.300 ;
        RECT 357.450 404.100 359.250 404.400 ;
        RECT 344.550 402.600 345.750 403.500 ;
        RECT 352.950 403.200 359.250 404.100 ;
        RECT 357.450 402.600 359.250 403.200 ;
        RECT 360.150 402.600 362.850 404.400 ;
        RECT 340.950 400.500 345.750 402.600 ;
        RECT 348.450 401.550 350.250 402.300 ;
        RECT 353.250 401.550 355.050 402.300 ;
        RECT 348.450 400.500 355.050 401.550 ;
        RECT 344.550 399.600 345.750 400.500 ;
        RECT 344.550 393.600 346.350 399.600 ;
        RECT 352.350 393.600 354.150 400.500 ;
        RECT 360.150 399.600 364.050 401.700 ;
        RECT 360.150 393.600 361.950 399.600 ;
        RECT 367.650 393.600 369.450 405.600 ;
        RECT 379.800 393.600 381.600 406.500 ;
        RECT 385.800 393.600 387.600 406.500 ;
        RECT 391.800 393.600 393.600 406.500 ;
        RECT 397.800 393.600 399.600 406.500 ;
        RECT 410.400 399.600 411.600 411.900 ;
        RECT 422.550 411.450 423.450 413.550 ;
        RECT 428.100 413.100 429.900 413.850 ;
        RECT 431.850 413.100 433.050 414.900 ;
        RECT 437.100 414.150 438.900 414.900 ;
        RECT 448.950 414.450 451.050 415.050 ;
        RECT 457.950 414.450 460.050 415.050 ;
        RECT 467.100 414.900 467.850 419.100 ;
        RECT 484.950 415.950 487.050 418.050 ;
        RECT 490.950 415.950 493.050 418.050 ;
        RECT 434.100 413.100 435.900 413.850 ;
        RECT 448.950 413.550 460.050 414.450 ;
        RECT 427.950 411.450 430.050 412.050 ;
        RECT 413.100 410.100 414.900 410.850 ;
        RECT 422.550 410.550 430.050 411.450 ;
        RECT 427.950 409.950 430.050 410.550 ;
        RECT 412.950 406.950 415.050 409.050 ;
        RECT 431.850 408.900 432.900 413.100 ;
        RECT 448.950 412.950 451.050 413.550 ;
        RECT 457.950 412.950 460.050 413.550 ;
        RECT 433.950 409.950 436.050 412.050 ;
        RECT 446.100 410.100 447.900 410.850 ;
        RECT 431.850 405.600 433.050 408.900 ;
        RECT 445.950 406.950 448.050 409.050 ;
        RECT 410.400 393.600 412.200 399.600 ;
        RECT 431.700 393.600 433.500 405.600 ;
        RECT 449.400 399.600 450.600 411.900 ;
        RECT 452.100 410.100 453.900 410.850 ;
        RECT 451.950 406.950 454.050 409.050 ;
        RECT 463.800 405.600 465.000 414.900 ;
        RECT 466.950 408.300 467.850 414.900 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 482.100 413.100 483.900 413.850 ;
        RECT 485.850 413.100 487.050 414.900 ;
        RECT 491.100 414.150 492.900 414.900 ;
        RECT 488.100 413.100 489.900 413.850 ;
        RECT 470.100 411.150 471.900 411.900 ;
        RECT 481.950 409.950 484.050 412.050 ;
        RECT 465.900 407.400 467.850 408.300 ;
        RECT 485.850 408.900 486.900 413.100 ;
        RECT 487.950 409.950 490.050 412.050 ;
        RECT 465.900 406.500 471.600 407.400 ;
        RECT 448.800 393.600 450.600 399.600 ;
        RECT 463.500 393.600 465.300 405.600 ;
        RECT 470.400 399.600 471.600 406.500 ;
        RECT 485.850 405.600 487.050 408.900 ;
        RECT 495.150 407.700 496.050 422.400 ;
        RECT 503.550 421.800 505.350 423.600 ;
        RECT 506.850 422.550 511.800 423.600 ;
        RECT 519.300 424.500 520.350 425.400 ;
        RECT 519.300 423.300 523.050 424.500 ;
        RECT 506.850 421.800 508.650 422.550 ;
        RECT 520.950 422.400 523.050 423.300 ;
        RECT 526.650 422.400 528.450 428.400 ;
        RECT 538.800 425.400 540.600 428.400 ;
        RECT 503.850 418.800 504.900 421.800 ;
        RECT 498.000 417.600 515.850 418.800 ;
        RECT 527.250 418.050 528.450 422.400 ;
        RECT 498.000 416.850 498.900 417.600 ;
        RECT 503.100 417.000 504.900 417.600 ;
        RECT 514.050 417.000 515.850 417.600 ;
        RECT 497.100 415.050 498.900 416.850 ;
        RECT 514.050 416.100 514.950 417.000 ;
        RECT 522.150 416.250 522.900 418.050 ;
        RECT 523.950 415.950 526.050 418.050 ;
        RECT 527.100 415.950 528.450 418.050 ;
        RECT 500.100 412.800 501.900 413.400 ;
        RECT 500.100 411.600 504.900 412.800 ;
        RECT 505.950 409.950 508.050 415.050 ;
        RECT 511.950 412.950 514.050 415.050 ;
        RECT 504.450 407.700 506.250 408.000 ;
        RECT 495.150 407.100 506.250 407.700 ;
        RECT 495.150 406.500 512.850 407.100 ;
        RECT 495.150 405.600 496.050 406.500 ;
        RECT 504.450 406.200 512.850 406.500 ;
        RECT 469.800 393.600 471.600 399.600 ;
        RECT 485.700 393.600 487.500 405.600 ;
        RECT 495.150 393.600 496.950 405.600 ;
        RECT 509.250 404.700 511.050 405.300 ;
        RECT 503.550 403.500 511.050 404.700 ;
        RECT 511.950 404.100 512.850 406.200 ;
        RECT 514.050 406.200 514.950 411.900 ;
        RECT 524.250 407.400 526.050 409.200 ;
        RECT 520.950 406.200 525.150 407.400 ;
        RECT 514.050 405.300 520.050 406.200 ;
        RECT 520.950 405.300 523.050 406.200 ;
        RECT 527.250 405.600 528.450 415.950 ;
        RECT 539.400 413.100 540.600 425.400 ;
        RECT 551.400 425.400 553.200 428.400 ;
        RECT 568.800 425.400 570.600 428.400 ;
        RECT 551.400 422.100 552.600 425.400 ;
        RECT 550.950 420.450 553.050 421.050 ;
        RECT 562.950 420.450 565.050 421.050 ;
        RECT 550.950 419.550 565.050 420.450 ;
        RECT 550.950 418.950 553.050 419.550 ;
        RECT 562.950 418.950 565.050 419.550 ;
        RECT 541.950 415.950 544.050 418.050 ;
        RECT 551.700 416.100 553.050 417.900 ;
        RECT 542.100 414.150 543.900 414.900 ;
        RECT 538.950 409.950 541.050 412.050 ;
        RECT 544.950 409.950 550.050 412.050 ;
        RECT 551.700 411.900 552.900 416.100 ;
        RECT 553.950 412.950 556.050 415.050 ;
        RECT 569.400 413.100 570.600 425.400 ;
        RECT 584.400 425.400 586.200 428.400 ;
        RECT 584.400 422.100 585.600 425.400 ;
        RECT 594.150 422.400 595.950 428.400 ;
        RECT 601.950 426.300 603.750 428.400 ;
        RECT 600.000 425.400 603.750 426.300 ;
        RECT 609.750 425.400 611.550 428.400 ;
        RECT 617.550 425.400 619.350 428.400 ;
        RECT 600.000 424.500 601.050 425.400 ;
        RECT 598.950 422.400 601.050 424.500 ;
        RECT 609.750 423.600 610.800 425.400 ;
        RECT 571.950 417.450 574.050 418.050 ;
        RECT 577.950 417.450 580.050 421.050 ;
        RECT 583.950 420.450 586.050 421.050 ;
        RECT 588.000 420.450 592.050 421.050 ;
        RECT 583.950 419.550 592.050 420.450 ;
        RECT 583.950 418.950 586.050 419.550 ;
        RECT 588.000 418.950 592.050 419.550 ;
        RECT 571.950 417.000 580.050 417.450 ;
        RECT 571.950 416.550 579.450 417.000 ;
        RECT 571.950 415.950 574.050 416.550 ;
        RECT 584.700 416.100 586.050 417.900 ;
        RECT 572.100 414.150 573.900 414.900 ;
        RECT 519.150 404.400 520.050 405.300 ;
        RECT 516.450 404.100 518.250 404.400 ;
        RECT 503.550 402.600 504.750 403.500 ;
        RECT 511.950 403.200 518.250 404.100 ;
        RECT 516.450 402.600 518.250 403.200 ;
        RECT 519.150 402.600 521.850 404.400 ;
        RECT 499.950 400.500 504.750 402.600 ;
        RECT 507.450 401.550 509.250 402.300 ;
        RECT 512.250 401.550 514.050 402.300 ;
        RECT 507.450 400.500 514.050 401.550 ;
        RECT 503.550 399.600 504.750 400.500 ;
        RECT 503.550 393.600 505.350 399.600 ;
        RECT 511.350 393.600 513.150 400.500 ;
        RECT 519.150 399.600 523.050 401.700 ;
        RECT 519.150 393.600 520.950 399.600 ;
        RECT 526.650 393.600 528.450 405.600 ;
        RECT 539.400 399.600 540.600 408.900 ;
        RECT 548.100 408.150 549.900 408.900 ;
        RECT 551.700 406.650 553.050 411.900 ;
        RECT 554.100 411.150 555.900 411.900 ;
        RECT 568.950 409.950 574.050 412.050 ;
        RECT 577.950 409.950 583.050 412.050 ;
        RECT 584.700 411.900 585.900 416.100 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 551.700 405.600 554.400 406.650 ;
        RECT 538.800 393.600 540.600 399.600 ;
        RECT 552.600 393.600 554.400 405.600 ;
        RECT 569.400 399.600 570.600 408.900 ;
        RECT 581.100 408.150 582.900 408.900 ;
        RECT 584.700 406.650 586.050 411.900 ;
        RECT 587.100 411.150 588.900 411.900 ;
        RECT 594.150 407.700 595.050 422.400 ;
        RECT 602.550 421.800 604.350 423.600 ;
        RECT 605.850 422.550 610.800 423.600 ;
        RECT 618.300 424.500 619.350 425.400 ;
        RECT 618.300 423.300 622.050 424.500 ;
        RECT 605.850 421.800 607.650 422.550 ;
        RECT 619.950 422.400 622.050 423.300 ;
        RECT 625.650 422.400 627.450 428.400 ;
        RECT 634.800 427.500 642.600 428.400 ;
        RECT 634.800 422.400 636.600 427.500 ;
        RECT 637.800 422.400 639.600 426.600 ;
        RECT 640.800 423.000 642.600 427.500 ;
        RECT 646.800 423.000 648.600 428.400 ;
        RECT 658.800 425.400 660.600 428.400 ;
        RECT 602.850 418.800 603.900 421.800 ;
        RECT 597.000 417.600 614.850 418.800 ;
        RECT 626.250 418.050 627.450 422.400 ;
        RECT 638.400 420.900 639.300 422.400 ;
        RECT 640.800 422.100 648.600 423.000 ;
        RECT 638.400 419.700 642.600 420.900 ;
        RECT 641.400 419.100 642.600 419.700 ;
        RECT 646.950 419.100 648.750 419.850 ;
        RECT 597.000 416.850 597.900 417.600 ;
        RECT 602.100 417.000 603.900 417.600 ;
        RECT 613.050 417.000 614.850 417.600 ;
        RECT 596.100 415.050 597.900 416.850 ;
        RECT 613.050 416.100 613.950 417.000 ;
        RECT 621.150 416.250 621.900 418.050 ;
        RECT 622.950 415.950 625.050 418.050 ;
        RECT 626.100 415.950 627.450 418.050 ;
        RECT 634.950 415.950 637.050 418.200 ;
        RECT 640.950 415.950 643.050 418.050 ;
        RECT 646.950 415.950 649.050 418.050 ;
        RECT 599.100 412.800 600.900 413.400 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 599.100 411.600 603.900 412.800 ;
        RECT 604.950 409.950 610.050 412.050 ;
        RECT 603.450 407.700 605.250 408.000 ;
        RECT 594.150 407.100 605.250 407.700 ;
        RECT 584.700 405.600 587.400 406.650 ;
        RECT 568.800 393.600 570.600 399.600 ;
        RECT 585.600 393.600 587.400 405.600 ;
        RECT 594.150 406.500 611.850 407.100 ;
        RECT 594.150 405.600 595.050 406.500 ;
        RECT 603.450 406.200 611.850 406.500 ;
        RECT 594.150 393.600 595.950 405.600 ;
        RECT 608.250 404.700 610.050 405.300 ;
        RECT 602.550 403.500 610.050 404.700 ;
        RECT 610.950 404.100 611.850 406.200 ;
        RECT 613.050 406.200 613.950 411.900 ;
        RECT 623.250 407.400 625.050 409.200 ;
        RECT 619.950 406.200 624.150 407.400 ;
        RECT 613.050 405.300 619.050 406.200 ;
        RECT 619.950 405.300 622.050 406.200 ;
        RECT 626.250 405.600 627.450 415.950 ;
        RECT 635.250 414.150 637.050 414.900 ;
        RECT 638.700 413.100 640.500 413.850 ;
        RECT 637.950 409.950 640.050 412.050 ;
        RECT 641.400 405.600 642.600 414.900 ;
        RECT 644.100 413.100 645.900 413.850 ;
        RECT 659.400 413.100 660.600 425.400 ;
        RECT 665.550 422.400 667.350 428.400 ;
        RECT 673.650 425.400 675.450 428.400 ;
        RECT 681.450 425.400 683.250 428.400 ;
        RECT 689.250 426.300 691.050 428.400 ;
        RECT 689.250 425.400 693.000 426.300 ;
        RECT 673.650 424.500 674.700 425.400 ;
        RECT 670.950 423.300 674.700 424.500 ;
        RECT 682.200 423.600 683.250 425.400 ;
        RECT 691.950 424.500 693.000 425.400 ;
        RECT 670.950 422.400 673.050 423.300 ;
        RECT 682.200 422.550 687.150 423.600 ;
        RECT 665.550 418.050 666.750 422.400 ;
        RECT 685.350 421.800 687.150 422.550 ;
        RECT 688.650 421.800 690.450 423.600 ;
        RECT 691.950 422.400 694.050 424.500 ;
        RECT 697.050 422.400 698.850 428.400 ;
        RECT 709.800 422.400 711.600 428.400 ;
        RECT 689.100 418.800 690.150 421.800 ;
        RECT 661.950 415.950 664.050 418.050 ;
        RECT 665.550 415.950 666.900 418.050 ;
        RECT 667.950 415.950 670.050 418.050 ;
        RECT 671.100 416.250 671.850 418.050 ;
        RECT 678.150 417.600 696.000 418.800 ;
        RECT 678.150 417.000 679.950 417.600 ;
        RECT 689.100 417.000 690.900 417.600 ;
        RECT 679.050 416.100 679.950 417.000 ;
        RECT 695.100 416.850 696.000 417.600 ;
        RECT 662.100 414.150 663.900 414.900 ;
        RECT 643.950 409.950 646.050 412.050 ;
        RECT 649.950 411.450 652.050 412.050 ;
        RECT 658.950 411.450 661.050 412.050 ;
        RECT 649.950 410.550 661.050 411.450 ;
        RECT 649.950 409.950 652.050 410.550 ;
        RECT 658.950 409.950 661.050 410.550 ;
        RECT 618.150 404.400 619.050 405.300 ;
        RECT 615.450 404.100 617.250 404.400 ;
        RECT 602.550 402.600 603.750 403.500 ;
        RECT 610.950 403.200 617.250 404.100 ;
        RECT 615.450 402.600 617.250 403.200 ;
        RECT 618.150 402.600 620.850 404.400 ;
        RECT 598.950 400.500 603.750 402.600 ;
        RECT 606.450 401.550 608.250 402.300 ;
        RECT 611.250 401.550 613.050 402.300 ;
        RECT 606.450 400.500 613.050 401.550 ;
        RECT 602.550 399.600 603.750 400.500 ;
        RECT 602.550 393.600 604.350 399.600 ;
        RECT 610.350 393.600 612.150 400.500 ;
        RECT 618.150 399.600 622.050 401.700 ;
        RECT 618.150 393.600 619.950 399.600 ;
        RECT 625.650 393.600 627.450 405.600 ;
        RECT 640.800 393.600 644.100 405.600 ;
        RECT 659.400 399.600 660.600 408.900 ;
        RECT 658.800 393.600 660.600 399.600 ;
        RECT 665.550 405.600 666.750 415.950 ;
        RECT 695.100 415.050 696.900 416.850 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 692.100 412.800 693.900 413.400 ;
        RECT 667.950 407.400 669.750 409.200 ;
        RECT 668.850 406.200 673.050 407.400 ;
        RECT 679.050 406.200 679.950 411.900 ;
        RECT 685.950 409.950 688.050 412.050 ;
        RECT 689.100 411.600 693.900 412.800 ;
        RECT 687.750 407.700 689.550 408.000 ;
        RECT 697.950 407.700 698.850 422.400 ;
        RECT 710.400 420.300 711.600 422.400 ;
        RECT 712.800 423.300 714.600 428.400 ;
        RECT 718.800 423.300 720.600 428.400 ;
        RECT 730.800 425.400 732.600 428.400 ;
        RECT 712.800 421.950 720.600 423.300 ;
        RECT 710.400 419.250 714.150 420.300 ;
        RECT 712.950 419.100 714.150 419.250 ;
        RECT 700.950 417.450 703.050 418.050 ;
        RECT 712.950 417.450 715.050 418.050 ;
        RECT 700.950 416.550 715.050 417.450 ;
        RECT 700.950 415.950 703.050 416.550 ;
        RECT 712.950 415.950 715.050 416.550 ;
        RECT 718.950 415.950 721.050 418.050 ;
        RECT 703.950 411.450 706.050 415.050 ;
        RECT 710.100 413.100 711.900 413.850 ;
        RECT 713.850 413.100 715.050 414.900 ;
        RECT 719.100 414.150 720.900 414.900 ;
        RECT 716.100 413.100 717.900 413.850 ;
        RECT 731.400 413.100 732.600 425.400 ;
        RECT 753.000 422.400 754.800 428.400 ;
        RECT 762.150 422.400 763.950 428.400 ;
        RECT 769.950 426.300 771.750 428.400 ;
        RECT 768.000 425.400 771.750 426.300 ;
        RECT 777.750 425.400 779.550 428.400 ;
        RECT 785.550 425.400 787.350 428.400 ;
        RECT 768.000 424.500 769.050 425.400 ;
        RECT 766.950 422.400 769.050 424.500 ;
        RECT 777.750 423.600 778.800 425.400 ;
        RECT 753.000 419.100 754.050 422.400 ;
        RECT 733.950 415.950 736.050 418.050 ;
        RECT 745.950 415.950 748.050 418.050 ;
        RECT 751.950 415.950 754.050 418.050 ;
        RECT 757.950 415.950 760.050 418.050 ;
        RECT 734.100 414.150 735.900 414.900 ;
        RECT 746.100 414.150 747.900 414.900 ;
        RECT 749.250 413.100 751.050 413.850 ;
        RECT 751.950 413.100 752.850 414.900 ;
        RECT 757.950 414.150 759.750 414.900 ;
        RECT 754.950 413.100 756.750 413.850 ;
        RECT 709.950 411.450 712.050 412.050 ;
        RECT 703.950 411.000 712.050 411.450 ;
        RECT 704.550 410.550 712.050 411.000 ;
        RECT 709.950 409.950 712.050 410.550 ;
        RECT 687.750 407.100 698.850 407.700 ;
        RECT 665.550 393.600 667.350 405.600 ;
        RECT 670.950 405.300 673.050 406.200 ;
        RECT 673.950 405.300 679.950 406.200 ;
        RECT 681.150 406.500 698.850 407.100 ;
        RECT 681.150 406.200 689.550 406.500 ;
        RECT 673.950 404.400 674.850 405.300 ;
        RECT 672.150 402.600 674.850 404.400 ;
        RECT 675.750 404.100 677.550 404.400 ;
        RECT 681.150 404.100 682.050 406.200 ;
        RECT 697.950 405.600 698.850 406.500 ;
        RECT 713.850 408.900 714.900 413.100 ;
        RECT 715.950 409.950 718.050 412.050 ;
        RECT 730.950 411.450 733.050 412.050 ;
        RECT 722.550 411.000 733.050 411.450 ;
        RECT 721.950 410.550 733.050 411.000 ;
        RECT 713.850 405.600 715.050 408.900 ;
        RECT 721.950 406.950 724.050 410.550 ;
        RECT 730.950 409.950 733.050 410.550 ;
        RECT 748.950 409.950 751.050 412.050 ;
        RECT 752.100 408.900 752.850 413.100 ;
        RECT 754.950 409.950 757.050 412.050 ;
        RECT 675.750 403.200 682.050 404.100 ;
        RECT 682.950 404.700 684.750 405.300 ;
        RECT 682.950 403.500 690.450 404.700 ;
        RECT 675.750 402.600 677.550 403.200 ;
        RECT 689.250 402.600 690.450 403.500 ;
        RECT 670.950 399.600 674.850 401.700 ;
        RECT 679.950 401.550 681.750 402.300 ;
        RECT 684.750 401.550 686.550 402.300 ;
        RECT 679.950 400.500 686.550 401.550 ;
        RECT 689.250 400.500 694.050 402.600 ;
        RECT 673.050 393.600 674.850 399.600 ;
        RECT 680.850 393.600 682.650 400.500 ;
        RECT 689.250 399.600 690.450 400.500 ;
        RECT 688.650 393.600 690.450 399.600 ;
        RECT 697.050 393.600 698.850 405.600 ;
        RECT 713.700 393.600 715.500 405.600 ;
        RECT 731.400 399.600 732.600 408.900 ;
        RECT 751.950 407.400 752.850 408.900 ;
        RECT 748.800 406.500 752.850 407.400 ;
        RECT 762.150 407.700 763.050 422.400 ;
        RECT 770.550 421.800 772.350 423.600 ;
        RECT 773.850 422.550 778.800 423.600 ;
        RECT 786.300 424.500 787.350 425.400 ;
        RECT 786.300 423.300 790.050 424.500 ;
        RECT 773.850 421.800 775.650 422.550 ;
        RECT 787.950 422.400 790.050 423.300 ;
        RECT 793.650 422.400 795.450 428.400 ;
        RECT 770.850 418.800 771.900 421.800 ;
        RECT 765.000 417.600 782.850 418.800 ;
        RECT 794.250 418.050 795.450 422.400 ;
        RECT 806.400 425.400 808.200 428.400 ;
        RECT 765.000 416.850 765.900 417.600 ;
        RECT 770.100 417.000 771.900 417.600 ;
        RECT 781.050 417.000 782.850 417.600 ;
        RECT 764.100 415.050 765.900 416.850 ;
        RECT 781.050 416.100 781.950 417.000 ;
        RECT 789.150 416.250 789.900 418.050 ;
        RECT 790.950 415.950 793.050 418.050 ;
        RECT 794.100 415.950 795.450 418.050 ;
        RECT 799.950 415.950 805.050 418.050 ;
        RECT 767.100 412.800 768.900 413.400 ;
        RECT 778.950 412.950 781.050 415.050 ;
        RECT 767.100 411.600 771.900 412.800 ;
        RECT 772.950 409.950 775.050 412.050 ;
        RECT 771.450 407.700 773.250 408.000 ;
        RECT 762.150 407.100 773.250 407.700 ;
        RECT 762.150 406.500 779.850 407.100 ;
        RECT 730.800 393.600 732.600 399.600 ;
        RECT 745.800 394.500 747.600 405.600 ;
        RECT 748.800 395.400 750.600 406.500 ;
        RECT 762.150 405.600 763.050 406.500 ;
        RECT 771.450 406.200 779.850 406.500 ;
        RECT 751.800 404.400 759.600 405.300 ;
        RECT 751.800 394.500 753.600 404.400 ;
        RECT 745.800 393.600 753.600 394.500 ;
        RECT 757.800 393.600 759.600 404.400 ;
        RECT 762.150 393.600 763.950 405.600 ;
        RECT 776.250 404.700 778.050 405.300 ;
        RECT 770.550 403.500 778.050 404.700 ;
        RECT 778.950 404.100 779.850 406.200 ;
        RECT 781.050 406.200 781.950 411.900 ;
        RECT 791.250 407.400 793.050 409.200 ;
        RECT 787.950 406.200 792.150 407.400 ;
        RECT 781.050 405.300 787.050 406.200 ;
        RECT 787.950 405.300 790.050 406.200 ;
        RECT 794.250 405.600 795.450 415.950 ;
        RECT 803.100 414.150 804.900 414.900 ;
        RECT 806.400 413.100 807.600 425.400 ;
        RECT 823.200 421.200 825.000 428.400 ;
        RECT 821.400 420.300 825.000 421.200 ;
        RECT 821.400 416.100 822.600 420.300 ;
        RECT 820.950 414.450 823.050 415.050 ;
        RECT 825.000 414.450 829.050 415.050 ;
        RECT 820.950 413.550 829.050 414.450 ;
        RECT 820.950 412.950 823.050 413.550 ;
        RECT 825.000 412.950 829.050 413.550 ;
        RECT 802.950 409.950 808.050 412.050 ;
        RECT 818.100 410.100 819.900 410.850 ;
        RECT 786.150 404.400 787.050 405.300 ;
        RECT 783.450 404.100 785.250 404.400 ;
        RECT 770.550 402.600 771.750 403.500 ;
        RECT 778.950 403.200 785.250 404.100 ;
        RECT 783.450 402.600 785.250 403.200 ;
        RECT 786.150 402.600 788.850 404.400 ;
        RECT 766.950 400.500 771.750 402.600 ;
        RECT 774.450 401.550 776.250 402.300 ;
        RECT 779.250 401.550 781.050 402.300 ;
        RECT 774.450 400.500 781.050 401.550 ;
        RECT 770.550 399.600 771.750 400.500 ;
        RECT 770.550 393.600 772.350 399.600 ;
        RECT 778.350 393.600 780.150 400.500 ;
        RECT 786.150 399.600 790.050 401.700 ;
        RECT 786.150 393.600 787.950 399.600 ;
        RECT 793.650 393.600 795.450 405.600 ;
        RECT 806.400 399.600 807.600 408.900 ;
        RECT 817.950 406.950 820.050 409.050 ;
        RECT 821.400 399.600 822.600 411.900 ;
        RECT 824.100 410.100 825.900 410.850 ;
        RECT 823.950 406.950 826.050 409.050 ;
        RECT 806.400 393.600 808.200 399.600 ;
        RECT 821.400 393.600 823.200 399.600 ;
        RECT 10.800 377.400 12.600 389.400 ;
        RECT 13.800 378.300 15.600 389.400 ;
        RECT 19.800 378.300 21.600 389.400 ;
        RECT 31.800 383.400 33.600 389.400 ;
        RECT 13.800 377.400 21.600 378.300 ;
        RECT 32.700 383.100 33.600 383.400 ;
        RECT 37.800 383.400 39.600 389.400 ;
        RECT 37.800 383.100 39.300 383.400 ;
        RECT 32.700 382.200 39.300 383.100 ;
        RECT 11.400 368.100 12.300 377.400 ;
        RECT 32.700 377.100 33.600 382.200 ;
        RECT 40.950 376.800 43.050 379.050 ;
        RECT 51.600 377.400 53.400 389.400 ;
        RECT 64.800 383.400 66.600 389.400 ;
        RECT 51.600 376.350 54.300 377.400 ;
        RECT 25.950 375.450 30.000 376.050 ;
        RECT 31.950 375.450 34.050 376.050 ;
        RECT 25.950 374.550 34.050 375.450 ;
        RECT 41.100 375.150 42.900 375.900 ;
        RECT 25.950 373.950 30.000 374.550 ;
        RECT 31.950 373.950 34.050 374.550 ;
        RECT 38.100 374.100 39.900 374.850 ;
        RECT 13.950 370.950 16.050 373.050 ;
        RECT 19.950 370.950 22.050 373.050 ;
        RECT 14.100 369.150 15.900 369.900 ;
        RECT 20.100 369.150 21.900 369.900 ;
        RECT 17.100 368.100 18.900 368.850 ;
        RECT 1.950 366.450 4.050 367.050 ;
        RECT 10.950 366.450 13.050 367.050 ;
        RECT 1.950 365.550 13.050 366.450 ;
        RECT 1.950 364.950 4.050 365.550 ;
        RECT 10.950 364.950 13.050 365.550 ;
        RECT 16.950 364.950 19.050 367.050 ;
        RECT 32.700 364.650 33.600 372.900 ;
        RECT 37.950 370.950 40.050 373.050 ;
        RECT 50.100 371.100 51.900 371.850 ;
        RECT 52.950 371.100 54.300 376.350 ;
        RECT 56.100 374.100 57.900 374.850 ;
        RECT 65.400 374.100 66.600 383.400 ;
        RECT 79.800 377.400 81.600 389.400 ;
        RECT 82.800 378.300 84.600 389.400 ;
        RECT 88.800 378.300 90.600 389.400 ;
        RECT 100.800 383.400 102.600 389.400 ;
        RECT 82.800 377.400 90.600 378.300 ;
        RECT 101.700 383.100 102.600 383.400 ;
        RECT 106.800 383.400 108.600 389.400 ;
        RECT 122.400 383.400 124.200 389.400 ;
        RECT 133.800 383.400 135.600 389.400 ;
        RECT 106.800 383.100 108.300 383.400 ;
        RECT 101.700 382.200 108.300 383.100 ;
        RECT 34.950 367.950 37.050 370.050 ;
        RECT 49.950 367.950 52.050 370.050 ;
        RECT 53.100 366.900 54.300 371.100 ;
        RECT 55.950 370.950 58.050 373.050 ;
        RECT 61.950 370.950 67.050 373.050 ;
        RECT 35.100 366.150 36.900 366.900 ;
        RECT 52.950 365.100 54.300 366.900 ;
        RECT 11.400 360.600 12.300 363.900 ;
        RECT 32.700 363.000 36.900 364.650 ;
        RECT 11.400 358.950 16.800 360.600 ;
        RECT 15.000 354.600 16.800 358.950 ;
        RECT 35.100 354.600 36.900 363.000 ;
        RECT 43.950 363.450 46.050 364.050 ;
        RECT 52.950 363.450 55.050 364.050 ;
        RECT 43.950 362.550 55.050 363.450 ;
        RECT 43.950 361.950 46.050 362.550 ;
        RECT 52.950 361.950 55.050 362.550 ;
        RECT 53.400 357.600 54.600 360.900 ;
        RECT 65.400 357.600 66.600 369.900 ;
        RECT 68.100 368.100 69.900 368.850 ;
        RECT 80.400 368.100 81.300 377.400 ;
        RECT 101.700 377.100 102.600 382.200 ;
        RECT 109.950 376.950 112.050 379.050 ;
        RECT 97.950 373.950 103.050 376.050 ;
        RECT 110.100 375.150 111.900 375.900 ;
        RECT 107.100 374.100 108.900 374.850 ;
        RECT 122.400 374.100 123.600 383.400 ;
        RECT 134.700 383.100 135.600 383.400 ;
        RECT 139.800 383.400 141.600 389.400 ;
        RECT 152.400 383.400 154.200 389.400 ;
        RECT 139.800 383.100 141.300 383.400 ;
        RECT 134.700 382.200 141.300 383.100 ;
        RECT 134.700 377.100 135.600 382.200 ;
        RECT 142.950 376.950 145.050 379.050 ;
        RECT 152.400 376.500 153.600 383.400 ;
        RECT 158.700 377.400 160.500 389.400 ;
        RECT 172.800 383.400 174.600 389.400 ;
        RECT 173.700 383.100 174.600 383.400 ;
        RECT 178.800 383.400 180.600 389.400 ;
        RECT 178.800 383.100 180.300 383.400 ;
        RECT 173.700 382.200 180.300 383.100 ;
        RECT 130.950 373.950 136.050 376.050 ;
        RECT 143.100 375.150 144.900 375.900 ;
        RECT 152.400 375.600 158.100 376.500 ;
        RECT 140.100 374.100 141.900 374.850 ;
        RECT 156.150 374.700 158.100 375.600 ;
        RECT 82.950 370.950 85.050 373.050 ;
        RECT 88.950 370.950 91.050 373.050 ;
        RECT 83.100 369.150 84.900 369.900 ;
        RECT 89.100 369.150 90.900 369.900 ;
        RECT 86.100 368.100 87.900 368.850 ;
        RECT 67.950 364.950 70.050 367.050 ;
        RECT 76.950 364.950 82.050 367.050 ;
        RECT 85.950 364.950 88.050 367.050 ;
        RECT 101.700 364.650 102.600 372.900 ;
        RECT 106.950 370.950 109.050 373.050 ;
        RECT 121.950 372.450 124.050 373.050 ;
        RECT 126.000 372.450 130.050 373.050 ;
        RECT 121.950 371.550 130.050 372.450 ;
        RECT 121.950 370.950 124.050 371.550 ;
        RECT 126.000 370.950 130.050 371.550 ;
        RECT 103.950 367.950 106.050 370.050 ;
        RECT 119.100 368.100 120.900 368.850 ;
        RECT 104.100 366.150 105.900 366.900 ;
        RECT 118.950 364.950 121.050 367.050 ;
        RECT 80.400 360.600 81.300 363.900 ;
        RECT 101.700 363.000 105.900 364.650 ;
        RECT 80.400 358.950 85.800 360.600 ;
        RECT 52.800 354.600 54.600 357.600 ;
        RECT 64.800 354.600 66.600 357.600 ;
        RECT 84.000 354.600 85.800 358.950 ;
        RECT 104.100 354.600 105.900 363.000 ;
        RECT 122.400 357.600 123.600 369.900 ;
        RECT 134.700 364.650 135.600 372.900 ;
        RECT 139.950 370.950 142.050 373.050 ;
        RECT 152.100 371.100 153.900 371.850 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 151.950 367.950 154.050 370.050 ;
        RECT 156.150 368.100 157.050 374.700 ;
        RECT 159.000 368.100 160.200 377.400 ;
        RECT 173.700 377.100 174.600 382.200 ;
        RECT 181.950 376.950 184.050 379.050 ;
        RECT 197.700 377.400 199.500 389.400 ;
        RECT 220.800 377.400 224.100 389.400 ;
        RECT 239.700 377.400 241.500 389.400 ;
        RECT 166.950 375.450 171.000 376.050 ;
        RECT 172.950 375.450 175.050 376.050 ;
        RECT 166.950 374.550 175.050 375.450 ;
        RECT 182.100 375.150 183.900 375.900 ;
        RECT 166.950 373.950 171.000 374.550 ;
        RECT 172.950 373.950 175.050 374.550 ;
        RECT 179.100 374.100 180.900 374.850 ;
        RECT 197.850 374.100 199.050 377.400 ;
        RECT 137.100 366.150 138.900 366.900 ;
        RECT 134.700 363.000 138.900 364.650 ;
        RECT 122.400 354.600 124.200 357.600 ;
        RECT 137.100 354.600 138.900 363.000 ;
        RECT 156.150 363.900 156.900 368.100 ;
        RECT 157.950 364.950 163.050 367.050 ;
        RECT 173.700 364.650 174.600 372.900 ;
        RECT 178.950 370.950 181.050 373.050 ;
        RECT 193.950 370.950 196.050 373.050 ;
        RECT 175.950 367.950 178.050 370.050 ;
        RECT 197.850 369.900 198.900 374.100 ;
        RECT 199.950 370.950 202.050 373.050 ;
        RECT 217.950 370.950 220.050 373.050 ;
        RECT 194.100 369.150 195.900 369.900 ;
        RECT 197.850 368.100 199.050 369.900 ;
        RECT 200.100 369.150 201.900 369.900 ;
        RECT 218.700 369.150 220.500 369.900 ;
        RECT 203.100 368.100 204.900 368.850 ;
        RECT 215.250 368.100 217.050 368.850 ;
        RECT 221.400 368.100 222.600 377.400 ;
        RECT 239.850 374.100 241.050 377.400 ;
        RECT 256.800 376.500 258.600 389.400 ;
        RECT 262.800 376.500 264.600 389.400 ;
        RECT 268.800 376.500 270.600 389.400 ;
        RECT 274.800 376.500 276.600 389.400 ;
        RECT 255.900 375.300 258.600 376.500 ;
        RECT 260.700 375.300 264.600 376.500 ;
        RECT 266.700 375.300 270.600 376.500 ;
        RECT 272.700 375.300 276.600 376.500 ;
        RECT 288.600 377.400 290.400 389.400 ;
        RECT 296.550 377.400 298.350 389.400 ;
        RECT 304.050 383.400 305.850 389.400 ;
        RECT 301.950 381.300 305.850 383.400 ;
        RECT 311.850 382.500 313.650 389.400 ;
        RECT 319.650 383.400 321.450 389.400 ;
        RECT 320.250 382.500 321.450 383.400 ;
        RECT 310.950 381.450 317.550 382.500 ;
        RECT 310.950 380.700 312.750 381.450 ;
        RECT 315.750 380.700 317.550 381.450 ;
        RECT 320.250 380.400 325.050 382.500 ;
        RECT 303.150 378.600 305.850 380.400 ;
        RECT 306.750 379.800 308.550 380.400 ;
        RECT 306.750 378.900 313.050 379.800 ;
        RECT 320.250 379.500 321.450 380.400 ;
        RECT 306.750 378.600 308.550 378.900 ;
        RECT 304.950 377.700 305.850 378.600 ;
        RECT 288.600 376.350 291.300 377.400 ;
        RECT 223.950 370.950 226.050 373.050 ;
        RECT 235.950 370.950 238.050 373.050 ;
        RECT 239.850 369.900 240.900 374.100 ;
        RECT 241.950 370.950 244.050 373.050 ;
        RECT 255.900 371.100 256.800 375.300 ;
        RECT 224.100 369.150 225.900 369.900 ;
        RECT 236.100 369.150 237.900 369.900 ;
        RECT 239.850 368.100 241.050 369.900 ;
        RECT 242.100 369.150 243.900 369.900 ;
        RECT 245.100 368.100 246.900 368.850 ;
        RECT 250.950 367.950 256.050 370.050 ;
        RECT 176.100 366.150 177.900 366.900 ;
        RECT 196.950 364.950 199.050 367.050 ;
        RECT 202.950 364.950 205.050 367.050 ;
        RECT 214.950 364.950 217.050 367.050 ;
        RECT 220.950 364.950 223.050 367.050 ;
        RECT 226.950 364.950 229.050 367.050 ;
        RECT 232.950 366.450 237.000 367.050 ;
        RECT 238.950 366.450 241.050 367.050 ;
        RECT 232.950 365.550 241.050 366.450 ;
        RECT 232.950 364.950 237.000 365.550 ;
        RECT 238.950 364.950 241.050 365.550 ;
        RECT 244.950 364.950 247.050 367.050 ;
        RECT 156.150 363.300 157.050 363.900 ;
        RECT 156.150 362.400 158.100 363.300 ;
        RECT 153.000 361.500 158.100 362.400 ;
        RECT 153.000 357.600 154.200 361.500 ;
        RECT 159.000 360.600 160.200 363.900 ;
        RECT 173.700 363.000 177.900 364.650 ;
        RECT 196.950 363.750 198.150 363.900 ;
        RECT 152.400 354.600 154.200 357.600 ;
        RECT 158.700 354.600 160.500 360.600 ;
        RECT 176.100 354.600 177.900 363.000 ;
        RECT 194.400 362.700 198.150 363.750 ;
        RECT 221.400 363.300 222.600 363.900 ;
        RECT 194.400 360.600 195.600 362.700 ;
        RECT 218.400 362.100 222.600 363.300 ;
        RECT 226.950 363.150 228.750 363.900 ;
        RECT 238.950 363.750 240.150 363.900 ;
        RECT 236.400 362.700 240.150 363.750 ;
        RECT 255.900 362.700 256.800 366.900 ;
        RECT 257.700 364.800 259.500 365.400 ;
        RECT 260.700 364.800 261.900 375.300 ;
        RECT 257.700 363.600 261.900 364.800 ;
        RECT 263.700 364.800 265.500 365.400 ;
        RECT 266.700 364.800 267.900 375.300 ;
        RECT 263.700 363.600 267.900 364.800 ;
        RECT 269.700 364.800 271.500 365.400 ;
        RECT 272.700 364.800 273.900 375.300 ;
        RECT 287.100 371.100 288.900 371.850 ;
        RECT 289.950 371.100 291.300 376.350 ;
        RECT 293.100 374.100 294.900 374.850 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 290.100 366.900 291.300 371.100 ;
        RECT 292.950 370.950 295.050 373.050 ;
        RECT 275.100 366.150 276.900 366.900 ;
        RECT 289.950 365.100 291.300 366.900 ;
        RECT 296.550 367.050 297.750 377.400 ;
        RECT 301.950 376.800 304.050 377.700 ;
        RECT 304.950 376.800 310.950 377.700 ;
        RECT 299.850 375.600 304.050 376.800 ;
        RECT 298.950 373.800 300.750 375.600 ;
        RECT 310.050 371.100 310.950 376.800 ;
        RECT 312.150 376.800 313.050 378.900 ;
        RECT 313.950 378.300 321.450 379.500 ;
        RECT 313.950 377.700 315.750 378.300 ;
        RECT 328.050 377.400 329.850 389.400 ;
        RECT 340.800 377.400 342.600 389.400 ;
        RECT 343.800 378.300 345.600 389.400 ;
        RECT 349.800 378.300 351.600 389.400 ;
        RECT 343.800 377.400 351.600 378.300 ;
        RECT 312.150 376.500 320.550 376.800 ;
        RECT 328.950 376.500 329.850 377.400 ;
        RECT 312.150 375.900 329.850 376.500 ;
        RECT 318.750 375.300 329.850 375.900 ;
        RECT 318.750 375.000 320.550 375.300 ;
        RECT 316.950 370.950 319.050 373.050 ;
        RECT 320.100 370.200 324.900 371.400 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 323.100 369.600 324.900 370.200 ;
        RECT 269.700 363.600 273.900 364.800 ;
        RECT 296.550 364.950 297.900 367.050 ;
        RECT 298.950 364.950 301.050 367.050 ;
        RECT 302.100 364.950 302.850 366.750 ;
        RECT 310.050 366.000 310.950 366.900 ;
        RECT 326.100 366.150 327.900 367.950 ;
        RECT 309.150 365.400 310.950 366.000 ;
        RECT 320.100 365.400 321.900 366.000 ;
        RECT 326.100 365.400 327.000 366.150 ;
        RECT 260.700 362.700 261.900 363.600 ;
        RECT 266.700 362.700 267.900 363.600 ;
        RECT 272.700 362.700 273.900 363.600 ;
        RECT 193.800 354.600 195.600 360.600 ;
        RECT 196.800 359.700 204.600 361.050 ;
        RECT 218.400 360.600 219.300 362.100 ;
        RECT 196.800 354.600 198.600 359.700 ;
        RECT 202.800 354.600 204.600 359.700 ;
        RECT 214.800 355.500 216.600 360.600 ;
        RECT 217.800 356.400 219.600 360.600 ;
        RECT 220.800 360.000 228.600 360.900 ;
        RECT 236.400 360.600 237.600 362.700 ;
        RECT 255.900 361.500 258.600 362.700 ;
        RECT 260.700 361.500 264.600 362.700 ;
        RECT 266.700 361.500 270.600 362.700 ;
        RECT 272.700 361.500 276.600 362.700 ;
        RECT 289.950 361.950 295.050 364.050 ;
        RECT 220.800 355.500 222.600 360.000 ;
        RECT 214.800 354.600 222.600 355.500 ;
        RECT 226.800 354.600 228.600 360.000 ;
        RECT 235.800 354.600 237.600 360.600 ;
        RECT 238.800 359.700 246.600 361.050 ;
        RECT 238.800 354.600 240.600 359.700 ;
        RECT 244.800 354.600 246.600 359.700 ;
        RECT 256.800 354.600 258.600 361.500 ;
        RECT 262.800 354.600 264.600 361.500 ;
        RECT 268.800 354.600 270.600 361.500 ;
        RECT 274.800 354.600 276.600 361.500 ;
        RECT 290.400 357.600 291.600 360.900 ;
        RECT 289.800 354.600 291.600 357.600 ;
        RECT 296.550 360.600 297.750 364.950 ;
        RECT 309.150 364.200 327.000 365.400 ;
        RECT 320.100 361.200 321.150 364.200 ;
        RECT 296.550 354.600 298.350 360.600 ;
        RECT 301.950 359.700 304.050 360.600 ;
        RECT 316.350 360.450 318.150 361.200 ;
        RECT 301.950 358.500 305.700 359.700 ;
        RECT 304.650 357.600 305.700 358.500 ;
        RECT 313.200 359.400 318.150 360.450 ;
        RECT 319.650 359.400 321.450 361.200 ;
        RECT 328.950 360.600 329.850 375.300 ;
        RECT 341.400 368.100 342.300 377.400 ;
        RECT 359.400 376.500 361.200 389.400 ;
        RECT 365.400 376.500 367.200 389.400 ;
        RECT 371.400 376.500 373.200 389.400 ;
        RECT 377.400 376.500 379.200 389.400 ;
        RECT 387.150 377.400 388.950 389.400 ;
        RECT 395.550 383.400 397.350 389.400 ;
        RECT 395.550 382.500 396.750 383.400 ;
        RECT 403.350 382.500 405.150 389.400 ;
        RECT 411.150 383.400 412.950 389.400 ;
        RECT 391.950 380.400 396.750 382.500 ;
        RECT 399.450 381.450 406.050 382.500 ;
        RECT 399.450 380.700 401.250 381.450 ;
        RECT 404.250 380.700 406.050 381.450 ;
        RECT 411.150 381.300 415.050 383.400 ;
        RECT 395.550 379.500 396.750 380.400 ;
        RECT 408.450 379.800 410.250 380.400 ;
        RECT 395.550 378.300 403.050 379.500 ;
        RECT 401.250 377.700 403.050 378.300 ;
        RECT 403.950 378.900 410.250 379.800 ;
        RECT 387.150 376.500 388.050 377.400 ;
        RECT 403.950 376.800 404.850 378.900 ;
        RECT 408.450 378.600 410.250 378.900 ;
        RECT 411.150 378.600 413.850 380.400 ;
        RECT 411.150 377.700 412.050 378.600 ;
        RECT 396.450 376.500 404.850 376.800 ;
        RECT 359.400 375.300 363.300 376.500 ;
        RECT 365.400 375.300 369.300 376.500 ;
        RECT 371.400 375.300 375.300 376.500 ;
        RECT 377.400 375.300 380.100 376.500 ;
        RECT 343.950 370.950 346.050 373.050 ;
        RECT 349.950 370.950 352.050 373.050 ;
        RECT 344.100 369.150 345.900 369.900 ;
        RECT 350.100 369.150 351.900 369.900 ;
        RECT 347.100 368.100 348.900 368.850 ;
        RECT 331.950 366.450 334.050 367.050 ;
        RECT 340.950 366.450 343.050 367.050 ;
        RECT 331.950 365.550 343.050 366.450 ;
        RECT 331.950 364.950 334.050 365.550 ;
        RECT 340.950 364.950 343.050 365.550 ;
        RECT 346.950 364.950 349.050 367.050 ;
        RECT 359.100 366.150 360.900 366.900 ;
        RECT 362.100 364.800 363.300 375.300 ;
        RECT 364.500 364.800 366.300 365.400 ;
        RECT 313.200 357.600 314.250 359.400 ;
        RECT 322.950 358.500 325.050 360.600 ;
        RECT 322.950 357.600 324.000 358.500 ;
        RECT 304.650 354.600 306.450 357.600 ;
        RECT 312.450 354.600 314.250 357.600 ;
        RECT 320.250 356.700 324.000 357.600 ;
        RECT 320.250 354.600 322.050 356.700 ;
        RECT 328.050 354.600 329.850 360.600 ;
        RECT 341.400 360.600 342.300 363.900 ;
        RECT 362.100 363.600 366.300 364.800 ;
        RECT 368.100 364.800 369.300 375.300 ;
        RECT 370.500 364.800 372.300 365.400 ;
        RECT 368.100 363.600 372.300 364.800 ;
        RECT 374.100 364.800 375.300 375.300 ;
        RECT 379.200 371.100 380.100 375.300 ;
        RECT 387.150 375.900 404.850 376.500 ;
        RECT 406.050 376.800 412.050 377.700 ;
        RECT 412.950 376.800 415.050 377.700 ;
        RECT 418.650 377.400 420.450 389.400 ;
        RECT 427.800 377.400 429.600 389.400 ;
        RECT 430.800 378.300 432.600 389.400 ;
        RECT 436.800 378.300 438.600 389.400 ;
        RECT 430.800 377.400 438.600 378.300 ;
        RECT 450.600 377.400 452.400 389.400 ;
        RECT 461.400 378.300 463.200 389.400 ;
        RECT 467.400 378.300 469.200 389.400 ;
        RECT 461.400 377.400 469.200 378.300 ;
        RECT 470.400 377.400 472.200 389.400 ;
        RECT 477.150 377.400 478.950 389.400 ;
        RECT 485.550 383.400 487.350 389.400 ;
        RECT 485.550 382.500 486.750 383.400 ;
        RECT 493.350 382.500 495.150 389.400 ;
        RECT 501.150 383.400 502.950 389.400 ;
        RECT 481.950 380.400 486.750 382.500 ;
        RECT 489.450 381.450 496.050 382.500 ;
        RECT 489.450 380.700 491.250 381.450 ;
        RECT 494.250 380.700 496.050 381.450 ;
        RECT 501.150 381.300 505.050 383.400 ;
        RECT 485.550 379.500 486.750 380.400 ;
        RECT 498.450 379.800 500.250 380.400 ;
        RECT 485.550 378.300 493.050 379.500 ;
        RECT 491.250 377.700 493.050 378.300 ;
        RECT 493.950 378.900 500.250 379.800 ;
        RECT 387.150 375.300 398.250 375.900 ;
        RECT 379.950 367.950 385.050 370.050 ;
        RECT 376.500 364.800 378.300 365.400 ;
        RECT 374.100 363.600 378.300 364.800 ;
        RECT 362.100 362.700 363.300 363.600 ;
        RECT 368.100 362.700 369.300 363.600 ;
        RECT 374.100 362.700 375.300 363.600 ;
        RECT 379.200 362.700 380.100 366.900 ;
        RECT 359.400 361.500 363.300 362.700 ;
        RECT 365.400 361.500 369.300 362.700 ;
        RECT 371.400 361.500 375.300 362.700 ;
        RECT 377.400 361.500 380.100 362.700 ;
        RECT 341.400 358.950 346.800 360.600 ;
        RECT 345.000 354.600 346.800 358.950 ;
        RECT 359.400 354.600 361.200 361.500 ;
        RECT 365.400 354.600 367.200 361.500 ;
        RECT 371.400 354.600 373.200 361.500 ;
        RECT 377.400 354.600 379.200 361.500 ;
        RECT 387.150 360.600 388.050 375.300 ;
        RECT 396.450 375.000 398.250 375.300 ;
        RECT 392.100 370.200 396.900 371.400 ;
        RECT 397.950 370.950 400.050 373.050 ;
        RECT 406.050 371.100 406.950 376.800 ;
        RECT 412.950 375.600 417.150 376.800 ;
        RECT 416.250 373.800 418.050 375.600 ;
        RECT 392.100 369.600 393.900 370.200 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 389.100 366.150 390.900 367.950 ;
        RECT 419.250 367.050 420.450 377.400 ;
        RECT 428.400 368.100 429.300 377.400 ;
        RECT 449.700 376.350 452.400 377.400 ;
        RECT 446.100 374.100 447.900 374.850 ;
        RECT 430.950 370.950 433.050 373.050 ;
        RECT 436.950 370.950 439.050 373.050 ;
        RECT 442.950 370.950 448.050 373.050 ;
        RECT 449.700 371.100 451.050 376.350 ;
        RECT 452.100 371.100 453.900 371.850 ;
        RECT 431.100 369.150 432.900 369.900 ;
        RECT 437.100 369.150 438.900 369.900 ;
        RECT 434.100 368.100 435.900 368.850 ;
        RECT 390.000 365.400 390.900 366.150 ;
        RECT 406.050 366.000 406.950 366.900 ;
        RECT 395.100 365.400 396.900 366.000 ;
        RECT 406.050 365.400 407.850 366.000 ;
        RECT 390.000 364.200 407.850 365.400 ;
        RECT 414.150 364.950 414.900 366.750 ;
        RECT 415.950 364.950 418.050 367.050 ;
        RECT 419.100 364.950 420.450 367.050 ;
        RECT 421.950 366.450 426.000 367.050 ;
        RECT 427.950 366.450 430.050 367.050 ;
        RECT 421.950 365.550 430.050 366.450 ;
        RECT 421.950 364.950 426.000 365.550 ;
        RECT 427.950 364.950 430.050 365.550 ;
        RECT 433.950 364.950 436.050 367.050 ;
        RECT 449.700 366.900 450.900 371.100 ;
        RECT 460.950 370.950 463.050 373.050 ;
        RECT 466.950 370.950 469.050 373.050 ;
        RECT 451.950 367.950 454.050 370.050 ;
        RECT 461.100 369.150 462.900 369.900 ;
        RECT 467.100 369.150 468.900 369.900 ;
        RECT 464.100 368.100 465.900 368.850 ;
        RECT 470.700 368.100 471.600 377.400 ;
        RECT 477.150 376.500 478.050 377.400 ;
        RECT 493.950 376.800 494.850 378.900 ;
        RECT 498.450 378.600 500.250 378.900 ;
        RECT 501.150 378.600 503.850 380.400 ;
        RECT 501.150 377.700 502.050 378.600 ;
        RECT 486.450 376.500 494.850 376.800 ;
        RECT 477.150 375.900 494.850 376.500 ;
        RECT 496.050 376.800 502.050 377.700 ;
        RECT 502.950 376.800 505.050 377.700 ;
        RECT 508.650 377.400 510.450 389.400 ;
        RECT 477.150 375.300 488.250 375.900 ;
        RECT 449.700 365.100 451.050 366.900 ;
        RECT 463.950 364.950 466.050 367.050 ;
        RECT 469.950 364.950 475.050 367.050 ;
        RECT 395.850 361.200 396.900 364.200 ;
        RECT 387.150 354.600 388.950 360.600 ;
        RECT 391.950 358.500 394.050 360.600 ;
        RECT 395.550 359.400 397.350 361.200 ;
        RECT 398.850 360.450 400.650 361.200 ;
        RECT 419.250 360.600 420.450 364.950 ;
        RECT 398.850 359.400 403.800 360.450 ;
        RECT 412.950 359.700 415.050 360.600 ;
        RECT 393.000 357.600 394.050 358.500 ;
        RECT 402.750 357.600 403.800 359.400 ;
        RECT 411.300 358.500 415.050 359.700 ;
        RECT 411.300 357.600 412.350 358.500 ;
        RECT 393.000 356.700 396.750 357.600 ;
        RECT 394.950 354.600 396.750 356.700 ;
        RECT 402.750 354.600 404.550 357.600 ;
        RECT 410.550 354.600 412.350 357.600 ;
        RECT 418.650 354.600 420.450 360.600 ;
        RECT 428.400 360.600 429.300 363.900 ;
        RECT 442.950 363.450 447.000 364.050 ;
        RECT 448.950 363.450 451.050 364.050 ;
        RECT 442.950 362.550 451.050 363.450 ;
        RECT 442.950 361.950 447.000 362.550 ;
        RECT 448.950 361.950 451.050 362.550 ;
        RECT 428.400 358.950 433.800 360.600 ;
        RECT 432.000 354.600 433.800 358.950 ;
        RECT 449.400 357.600 450.600 360.900 ;
        RECT 470.700 360.600 471.600 363.900 ;
        RECT 466.200 358.950 471.600 360.600 ;
        RECT 477.150 360.600 478.050 375.300 ;
        RECT 486.450 375.000 488.250 375.300 ;
        RECT 482.100 370.200 486.900 371.400 ;
        RECT 487.950 370.950 490.050 373.050 ;
        RECT 496.050 371.100 496.950 376.800 ;
        RECT 502.950 375.600 507.150 376.800 ;
        RECT 506.250 373.800 508.050 375.600 ;
        RECT 482.100 369.600 483.900 370.200 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 479.100 366.150 480.900 367.950 ;
        RECT 509.250 367.050 510.450 377.400 ;
        RECT 480.000 365.400 480.900 366.150 ;
        RECT 496.050 366.000 496.950 366.900 ;
        RECT 485.100 365.400 486.900 366.000 ;
        RECT 496.050 365.400 497.850 366.000 ;
        RECT 480.000 364.200 497.850 365.400 ;
        RECT 504.150 364.950 504.900 366.750 ;
        RECT 505.950 364.950 508.050 367.050 ;
        RECT 509.100 364.950 510.450 367.050 ;
        RECT 485.850 361.200 486.900 364.200 ;
        RECT 449.400 354.600 451.200 357.600 ;
        RECT 466.200 354.600 468.000 358.950 ;
        RECT 477.150 354.600 478.950 360.600 ;
        RECT 481.950 358.500 484.050 360.600 ;
        RECT 485.550 359.400 487.350 361.200 ;
        RECT 488.850 360.450 490.650 361.200 ;
        RECT 509.250 360.600 510.450 364.950 ;
        RECT 488.850 359.400 493.800 360.450 ;
        RECT 502.950 359.700 505.050 360.600 ;
        RECT 483.000 357.600 484.050 358.500 ;
        RECT 492.750 357.600 493.800 359.400 ;
        RECT 501.300 358.500 505.050 359.700 ;
        RECT 501.300 357.600 502.350 358.500 ;
        RECT 483.000 356.700 486.750 357.600 ;
        RECT 484.950 354.600 486.750 356.700 ;
        RECT 492.750 354.600 494.550 357.600 ;
        RECT 500.550 354.600 502.350 357.600 ;
        RECT 508.650 354.600 510.450 360.600 ;
        RECT 513.150 377.400 514.950 389.400 ;
        RECT 521.550 383.400 523.350 389.400 ;
        RECT 521.550 382.500 522.750 383.400 ;
        RECT 529.350 382.500 531.150 389.400 ;
        RECT 537.150 383.400 538.950 389.400 ;
        RECT 517.950 380.400 522.750 382.500 ;
        RECT 525.450 381.450 532.050 382.500 ;
        RECT 525.450 380.700 527.250 381.450 ;
        RECT 530.250 380.700 532.050 381.450 ;
        RECT 537.150 381.300 541.050 383.400 ;
        RECT 521.550 379.500 522.750 380.400 ;
        RECT 534.450 379.800 536.250 380.400 ;
        RECT 521.550 378.300 529.050 379.500 ;
        RECT 527.250 377.700 529.050 378.300 ;
        RECT 529.950 378.900 536.250 379.800 ;
        RECT 513.150 376.500 514.050 377.400 ;
        RECT 529.950 376.800 530.850 378.900 ;
        RECT 534.450 378.600 536.250 378.900 ;
        RECT 537.150 378.600 539.850 380.400 ;
        RECT 537.150 377.700 538.050 378.600 ;
        RECT 522.450 376.500 530.850 376.800 ;
        RECT 513.150 375.900 530.850 376.500 ;
        RECT 532.050 376.800 538.050 377.700 ;
        RECT 538.950 376.800 541.050 377.700 ;
        RECT 544.650 377.400 546.450 389.400 ;
        RECT 555.600 377.400 557.400 389.400 ;
        RECT 571.800 383.400 573.600 389.400 ;
        RECT 513.150 375.300 524.250 375.900 ;
        RECT 513.150 360.600 514.050 375.300 ;
        RECT 522.450 375.000 524.250 375.300 ;
        RECT 518.100 370.200 522.900 371.400 ;
        RECT 518.100 369.600 519.900 370.200 ;
        RECT 523.950 367.950 526.050 373.050 ;
        RECT 532.050 371.100 532.950 376.800 ;
        RECT 538.950 375.600 543.150 376.800 ;
        RECT 542.250 373.800 544.050 375.600 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 515.100 366.150 516.900 367.950 ;
        RECT 545.250 367.050 546.450 377.400 ;
        RECT 554.700 376.350 557.400 377.400 ;
        RECT 551.100 374.100 552.900 374.850 ;
        RECT 547.950 370.950 553.050 373.050 ;
        RECT 554.700 371.100 556.050 376.350 ;
        RECT 572.400 374.100 573.600 383.400 ;
        RECT 578.550 377.400 580.350 389.400 ;
        RECT 586.050 383.400 587.850 389.400 ;
        RECT 583.950 381.300 587.850 383.400 ;
        RECT 593.850 382.500 595.650 389.400 ;
        RECT 601.650 383.400 603.450 389.400 ;
        RECT 602.250 382.500 603.450 383.400 ;
        RECT 592.950 381.450 599.550 382.500 ;
        RECT 592.950 380.700 594.750 381.450 ;
        RECT 597.750 380.700 599.550 381.450 ;
        RECT 602.250 380.400 607.050 382.500 ;
        RECT 585.150 378.600 587.850 380.400 ;
        RECT 588.750 379.800 590.550 380.400 ;
        RECT 588.750 378.900 595.050 379.800 ;
        RECT 602.250 379.500 603.450 380.400 ;
        RECT 588.750 378.600 590.550 378.900 ;
        RECT 586.950 377.700 587.850 378.600 ;
        RECT 557.100 371.100 558.900 371.850 ;
        RECT 516.000 365.400 516.900 366.150 ;
        RECT 532.050 366.000 532.950 366.900 ;
        RECT 521.100 365.400 522.900 366.000 ;
        RECT 532.050 365.400 533.850 366.000 ;
        RECT 516.000 364.200 533.850 365.400 ;
        RECT 540.150 364.950 540.900 366.750 ;
        RECT 541.950 364.950 544.050 367.050 ;
        RECT 545.100 364.950 546.450 367.050 ;
        RECT 554.700 366.900 555.900 371.100 ;
        RECT 571.950 370.950 574.050 373.050 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 554.700 365.100 556.050 366.900 ;
        RECT 521.850 361.200 522.900 364.200 ;
        RECT 513.150 354.600 514.950 360.600 ;
        RECT 517.950 358.500 520.050 360.600 ;
        RECT 521.550 359.400 523.350 361.200 ;
        RECT 524.850 360.450 526.650 361.200 ;
        RECT 545.250 360.600 546.450 364.950 ;
        RECT 550.950 361.950 556.050 364.050 ;
        RECT 524.850 359.400 529.800 360.450 ;
        RECT 538.950 359.700 541.050 360.600 ;
        RECT 519.000 357.600 520.050 358.500 ;
        RECT 528.750 357.600 529.800 359.400 ;
        RECT 537.300 358.500 541.050 359.700 ;
        RECT 537.300 357.600 538.350 358.500 ;
        RECT 519.000 356.700 522.750 357.600 ;
        RECT 520.950 354.600 522.750 356.700 ;
        RECT 528.750 354.600 530.550 357.600 ;
        RECT 536.550 354.600 538.350 357.600 ;
        RECT 544.650 354.600 546.450 360.600 ;
        RECT 554.400 357.600 555.600 360.900 ;
        RECT 572.400 357.600 573.600 369.900 ;
        RECT 575.100 368.100 576.900 368.850 ;
        RECT 578.550 367.050 579.750 377.400 ;
        RECT 583.950 376.800 586.050 377.700 ;
        RECT 586.950 376.800 592.950 377.700 ;
        RECT 581.850 375.600 586.050 376.800 ;
        RECT 580.950 373.800 582.750 375.600 ;
        RECT 592.050 371.100 592.950 376.800 ;
        RECT 594.150 376.800 595.050 378.900 ;
        RECT 595.950 378.300 603.450 379.500 ;
        RECT 595.950 377.700 597.750 378.300 ;
        RECT 610.050 377.400 611.850 389.400 ;
        RECT 623.700 377.400 625.500 389.400 ;
        RECT 638.400 383.400 640.200 389.400 ;
        RECT 594.150 376.500 602.550 376.800 ;
        RECT 610.950 376.500 611.850 377.400 ;
        RECT 594.150 375.900 611.850 376.500 ;
        RECT 600.750 375.300 611.850 375.900 ;
        RECT 600.750 375.000 602.550 375.300 ;
        RECT 598.950 370.950 601.050 373.050 ;
        RECT 602.100 370.200 606.900 371.400 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 605.100 369.600 606.900 370.200 ;
        RECT 574.950 364.950 577.050 367.050 ;
        RECT 578.550 364.950 579.900 367.050 ;
        RECT 580.950 364.950 583.050 367.050 ;
        RECT 584.100 364.950 584.850 366.750 ;
        RECT 592.050 366.000 592.950 366.900 ;
        RECT 608.100 366.150 609.900 367.950 ;
        RECT 591.150 365.400 592.950 366.000 ;
        RECT 602.100 365.400 603.900 366.000 ;
        RECT 608.100 365.400 609.000 366.150 ;
        RECT 554.400 354.600 556.200 357.600 ;
        RECT 571.800 354.600 573.600 357.600 ;
        RECT 578.550 360.600 579.750 364.950 ;
        RECT 591.150 364.200 609.000 365.400 ;
        RECT 602.100 361.200 603.150 364.200 ;
        RECT 578.550 354.600 580.350 360.600 ;
        RECT 583.950 359.700 586.050 360.600 ;
        RECT 598.350 360.450 600.150 361.200 ;
        RECT 583.950 358.500 587.700 359.700 ;
        RECT 586.650 357.600 587.700 358.500 ;
        RECT 595.200 359.400 600.150 360.450 ;
        RECT 601.650 359.400 603.450 361.200 ;
        RECT 610.950 360.600 611.850 375.300 ;
        RECT 623.850 374.100 625.050 377.400 ;
        RECT 638.400 374.100 639.600 383.400 ;
        RECT 651.600 377.400 653.400 389.400 ;
        RECT 669.600 377.400 671.400 389.400 ;
        RECT 684.900 377.400 688.200 389.400 ;
        RECT 703.800 377.400 705.600 389.400 ;
        RECT 706.800 378.300 708.600 389.400 ;
        RECT 712.800 378.300 714.600 389.400 ;
        RECT 706.800 377.400 714.600 378.300 ;
        RECT 722.400 377.400 724.200 389.400 ;
        RECT 729.900 378.900 731.700 389.400 ;
        RECT 729.900 377.400 732.300 378.900 ;
        RECT 650.700 376.350 653.400 377.400 ;
        RECT 668.700 376.350 671.400 377.400 ;
        RECT 647.100 374.100 648.900 374.850 ;
        RECT 619.950 370.950 622.050 373.050 ;
        RECT 623.850 369.900 624.900 374.100 ;
        RECT 625.950 370.950 628.050 373.050 ;
        RECT 637.950 370.950 640.050 373.050 ;
        RECT 640.950 372.450 645.000 373.050 ;
        RECT 646.950 372.450 649.050 373.050 ;
        RECT 640.950 371.550 649.050 372.450 ;
        RECT 640.950 370.950 645.000 371.550 ;
        RECT 646.950 370.950 649.050 371.550 ;
        RECT 650.700 371.100 652.050 376.350 ;
        RECT 665.100 374.100 666.900 374.850 ;
        RECT 653.100 371.100 654.900 371.850 ;
        RECT 620.100 369.150 621.900 369.900 ;
        RECT 623.850 368.100 625.050 369.900 ;
        RECT 626.100 369.150 627.900 369.900 ;
        RECT 629.100 368.100 630.900 368.850 ;
        RECT 635.100 368.100 636.900 368.850 ;
        RECT 622.950 364.950 625.050 367.050 ;
        RECT 628.950 364.950 631.050 367.050 ;
        RECT 634.950 364.950 637.050 367.050 ;
        RECT 622.950 363.750 624.150 363.900 ;
        RECT 620.400 362.700 624.150 363.750 ;
        RECT 620.400 360.600 621.600 362.700 ;
        RECT 595.200 357.600 596.250 359.400 ;
        RECT 604.950 358.500 607.050 360.600 ;
        RECT 604.950 357.600 606.000 358.500 ;
        RECT 586.650 354.600 588.450 357.600 ;
        RECT 594.450 354.600 596.250 357.600 ;
        RECT 602.250 356.700 606.000 357.600 ;
        RECT 602.250 354.600 604.050 356.700 ;
        RECT 610.050 354.600 611.850 360.600 ;
        RECT 619.800 354.600 621.600 360.600 ;
        RECT 622.800 359.700 630.600 361.050 ;
        RECT 622.800 354.600 624.600 359.700 ;
        RECT 628.800 354.600 630.600 359.700 ;
        RECT 638.400 357.600 639.600 369.900 ;
        RECT 650.700 366.900 651.900 371.100 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 664.950 367.950 667.050 373.050 ;
        RECT 668.700 371.100 670.050 376.350 ;
        RECT 671.100 371.100 672.900 371.850 ;
        RECT 668.700 366.900 669.900 371.100 ;
        RECT 682.950 370.950 685.050 373.050 ;
        RECT 670.950 367.950 673.050 370.050 ;
        RECT 683.100 369.150 684.900 369.900 ;
        RECT 686.400 368.100 687.600 377.400 ;
        RECT 688.950 370.950 691.050 373.050 ;
        RECT 688.500 369.150 690.300 369.900 ;
        RECT 691.950 368.100 693.750 368.850 ;
        RECT 704.400 368.100 705.300 377.400 ;
        RECT 722.400 376.200 723.600 377.400 ;
        RECT 722.400 375.000 729.600 376.200 ;
        RECT 727.800 374.400 729.600 375.000 ;
        RECT 706.950 370.950 709.050 373.050 ;
        RECT 712.950 370.950 715.050 373.050 ;
        RECT 721.950 370.950 724.050 373.050 ;
        RECT 707.100 369.150 708.900 369.900 ;
        RECT 713.100 369.150 714.900 369.900 ;
        RECT 722.100 369.150 723.900 369.900 ;
        RECT 710.100 368.100 711.900 368.850 ;
        RECT 725.100 368.100 726.900 368.850 ;
        RECT 650.700 365.100 652.050 366.900 ;
        RECT 668.700 365.100 670.050 366.900 ;
        RECT 679.950 364.950 682.050 367.050 ;
        RECT 685.950 364.950 688.050 367.050 ;
        RECT 691.950 364.950 694.050 367.050 ;
        RECT 703.950 364.950 706.050 367.050 ;
        RECT 709.950 364.950 712.050 367.050 ;
        RECT 724.950 364.950 727.050 367.050 ;
        RECT 649.950 363.450 652.050 364.050 ;
        RECT 654.000 363.450 658.050 364.050 ;
        RECT 649.950 362.550 658.050 363.450 ;
        RECT 649.950 361.950 652.050 362.550 ;
        RECT 654.000 361.950 658.050 362.550 ;
        RECT 667.950 363.450 670.050 364.050 ;
        RECT 667.950 362.550 675.450 363.450 ;
        RECT 680.250 363.150 682.050 363.900 ;
        RECT 686.400 363.300 687.600 363.900 ;
        RECT 667.950 361.950 670.050 362.550 ;
        RECT 674.550 361.050 675.450 362.550 ;
        RECT 686.400 362.100 690.600 363.300 ;
        RECT 650.400 357.600 651.600 360.900 ;
        RECT 668.400 357.600 669.600 360.900 ;
        RECT 674.550 359.550 679.050 361.050 ;
        RECT 675.000 358.950 679.050 359.550 ;
        RECT 680.400 360.000 688.200 360.900 ;
        RECT 689.700 360.600 690.600 362.100 ;
        RECT 704.400 360.600 705.300 363.900 ;
        RECT 728.700 363.600 729.600 374.400 ;
        RECT 730.950 371.100 732.300 377.400 ;
        RECT 738.150 377.400 739.950 389.400 ;
        RECT 746.550 383.400 748.350 389.400 ;
        RECT 746.550 382.500 747.750 383.400 ;
        RECT 754.350 382.500 756.150 389.400 ;
        RECT 762.150 383.400 763.950 389.400 ;
        RECT 742.950 380.400 747.750 382.500 ;
        RECT 750.450 381.450 757.050 382.500 ;
        RECT 750.450 380.700 752.250 381.450 ;
        RECT 755.250 380.700 757.050 381.450 ;
        RECT 762.150 381.300 766.050 383.400 ;
        RECT 746.550 379.500 747.750 380.400 ;
        RECT 759.450 379.800 761.250 380.400 ;
        RECT 746.550 378.300 754.050 379.500 ;
        RECT 752.250 377.700 754.050 378.300 ;
        RECT 754.950 378.900 761.250 379.800 ;
        RECT 738.150 376.500 739.050 377.400 ;
        RECT 754.950 376.800 755.850 378.900 ;
        RECT 759.450 378.600 761.250 378.900 ;
        RECT 762.150 378.600 764.850 380.400 ;
        RECT 762.150 377.700 763.050 378.600 ;
        RECT 747.450 376.500 755.850 376.800 ;
        RECT 738.150 375.900 755.850 376.500 ;
        RECT 757.050 376.800 763.050 377.700 ;
        RECT 763.950 376.800 766.050 377.700 ;
        RECT 769.650 377.400 771.450 389.400 ;
        RECT 738.150 375.300 749.250 375.900 ;
        RECT 730.950 367.950 736.050 370.050 ;
        RECT 727.950 362.700 729.750 363.600 ;
        RECT 726.300 361.800 729.750 362.700 ;
        RECT 638.400 354.600 640.200 357.600 ;
        RECT 650.400 354.600 652.200 357.600 ;
        RECT 668.400 354.600 670.200 357.600 ;
        RECT 680.400 354.600 682.200 360.000 ;
        RECT 686.400 355.500 688.200 360.000 ;
        RECT 689.400 356.400 691.200 360.600 ;
        RECT 692.400 355.500 694.200 360.600 ;
        RECT 704.400 358.950 709.800 360.600 ;
        RECT 686.400 354.600 694.200 355.500 ;
        RECT 708.000 354.600 709.800 358.950 ;
        RECT 726.300 357.600 727.200 361.800 ;
        RECT 732.000 360.600 733.050 366.900 ;
        RECT 738.150 360.600 739.050 375.300 ;
        RECT 747.450 375.000 749.250 375.300 ;
        RECT 743.100 370.200 747.900 371.400 ;
        RECT 743.100 369.600 744.900 370.200 ;
        RECT 748.950 367.950 751.050 373.050 ;
        RECT 757.050 371.100 757.950 376.800 ;
        RECT 763.950 375.600 768.150 376.800 ;
        RECT 767.250 373.800 769.050 375.600 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 740.100 366.150 741.900 367.950 ;
        RECT 770.250 367.050 771.450 377.400 ;
        RECT 783.600 377.400 785.400 389.400 ;
        RECT 799.800 383.400 801.600 389.400 ;
        RECT 783.600 376.350 786.300 377.400 ;
        RECT 782.100 371.100 783.900 371.850 ;
        RECT 784.950 371.100 786.300 376.350 ;
        RECT 788.100 374.100 789.900 374.850 ;
        RECT 800.400 374.100 801.600 383.400 ;
        RECT 814.500 377.400 816.300 389.400 ;
        RECT 817.950 378.450 820.050 379.050 ;
        RECT 823.950 378.450 826.050 379.050 ;
        RECT 817.950 377.550 826.050 378.450 ;
        RECT 814.950 374.100 816.150 377.400 ;
        RECT 817.950 376.950 820.050 377.550 ;
        RECT 823.950 376.950 826.050 377.550 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 741.000 365.400 741.900 366.150 ;
        RECT 757.050 366.000 757.950 366.900 ;
        RECT 746.100 365.400 747.900 366.000 ;
        RECT 757.050 365.400 758.850 366.000 ;
        RECT 741.000 364.200 758.850 365.400 ;
        RECT 765.150 364.950 765.900 366.750 ;
        RECT 766.950 364.950 769.050 367.050 ;
        RECT 770.100 364.950 771.450 367.050 ;
        RECT 785.100 366.900 786.300 371.100 ;
        RECT 787.950 370.950 793.050 373.050 ;
        RECT 799.950 370.800 802.050 373.050 ;
        RECT 811.950 370.950 814.050 373.050 ;
        RECT 815.100 369.900 816.150 374.100 ;
        RECT 817.950 370.950 820.050 373.050 ;
        RECT 784.950 365.100 786.300 366.900 ;
        RECT 746.850 361.200 747.900 364.200 ;
        RECT 725.400 354.600 727.200 357.600 ;
        RECT 731.400 354.600 733.200 360.600 ;
        RECT 738.150 354.600 739.950 360.600 ;
        RECT 742.950 358.500 745.050 360.600 ;
        RECT 746.550 359.400 748.350 361.200 ;
        RECT 749.850 360.450 751.650 361.200 ;
        RECT 770.250 360.600 771.450 364.950 ;
        RECT 784.950 363.450 787.050 364.050 ;
        RECT 789.000 363.450 793.050 364.050 ;
        RECT 784.950 362.550 793.050 363.450 ;
        RECT 784.950 361.950 787.050 362.550 ;
        RECT 789.000 361.950 793.050 362.550 ;
        RECT 749.850 359.400 754.800 360.450 ;
        RECT 763.950 359.700 766.050 360.600 ;
        RECT 744.000 357.600 745.050 358.500 ;
        RECT 753.750 357.600 754.800 359.400 ;
        RECT 762.300 358.500 766.050 359.700 ;
        RECT 762.300 357.600 763.350 358.500 ;
        RECT 744.000 356.700 747.750 357.600 ;
        RECT 745.950 354.600 747.750 356.700 ;
        RECT 753.750 354.600 755.550 357.600 ;
        RECT 761.550 354.600 763.350 357.600 ;
        RECT 769.650 354.600 771.450 360.600 ;
        RECT 785.400 357.600 786.600 360.900 ;
        RECT 800.400 357.600 801.600 369.900 ;
        RECT 812.100 369.150 813.900 369.900 ;
        RECT 803.100 368.100 804.900 368.850 ;
        RECT 809.100 368.100 810.900 368.850 ;
        RECT 814.950 368.100 816.150 369.900 ;
        RECT 818.100 369.150 819.900 369.900 ;
        RECT 802.950 364.950 805.050 367.050 ;
        RECT 808.950 364.950 811.050 367.050 ;
        RECT 814.950 364.950 817.050 367.050 ;
        RECT 815.850 363.750 817.050 363.900 ;
        RECT 815.850 362.700 819.600 363.750 ;
        RECT 784.800 354.600 786.600 357.600 ;
        RECT 799.800 354.600 801.600 357.600 ;
        RECT 809.400 359.700 817.200 361.050 ;
        RECT 809.400 354.600 811.200 359.700 ;
        RECT 815.400 354.600 817.200 359.700 ;
        RECT 818.400 360.600 819.600 362.700 ;
        RECT 818.400 354.600 820.200 360.600 ;
        RECT 9.000 343.200 10.800 350.400 ;
        RECT 25.800 347.400 27.600 350.400 ;
        RECT 9.000 342.300 12.600 343.200 ;
        RECT 11.400 338.100 12.600 342.300 ;
        RECT 4.950 336.450 9.000 337.050 ;
        RECT 10.950 336.450 13.050 337.050 ;
        RECT 4.950 335.550 13.050 336.450 ;
        RECT 4.950 334.950 9.000 335.550 ;
        RECT 10.950 334.950 13.050 335.550 ;
        RECT 26.400 335.100 27.600 347.400 ;
        RECT 45.000 346.050 46.800 350.400 ;
        RECT 41.400 344.400 46.800 346.050 ;
        RECT 41.400 341.100 42.300 344.400 ;
        RECT 62.100 342.000 63.900 350.400 ;
        RECT 79.200 343.200 81.000 350.400 ;
        RECT 95.400 347.400 97.200 350.400 ;
        RECT 77.400 342.300 81.000 343.200 ;
        RECT 96.300 343.200 97.200 347.400 ;
        RECT 101.400 344.400 103.200 350.400 ;
        RECT 96.300 342.300 99.750 343.200 ;
        RECT 62.100 340.350 66.300 342.000 ;
        RECT 28.950 337.950 31.050 340.050 ;
        RECT 37.950 337.950 43.050 340.050 ;
        RECT 46.950 337.950 49.050 340.050 ;
        RECT 62.100 338.100 63.900 338.850 ;
        RECT 29.100 336.150 30.900 336.900 ;
        RECT 8.100 332.100 9.900 332.850 ;
        RECT 7.950 328.950 10.050 331.050 ;
        RECT 11.400 321.600 12.600 333.900 ;
        RECT 25.950 333.450 28.050 334.050 ;
        RECT 37.950 333.450 40.050 334.050 ;
        RECT 14.100 332.100 15.900 332.850 ;
        RECT 25.950 332.550 40.050 333.450 ;
        RECT 25.950 331.950 28.050 332.550 ;
        RECT 37.950 331.950 40.050 332.550 ;
        RECT 13.950 328.950 16.050 331.050 ;
        RECT 26.400 321.600 27.600 330.900 ;
        RECT 41.400 327.600 42.300 336.900 ;
        RECT 47.100 336.150 48.900 336.900 ;
        RECT 44.100 335.100 45.900 335.850 ;
        RECT 50.100 335.100 51.900 335.850 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 43.950 331.950 46.050 334.050 ;
        RECT 49.950 331.950 52.050 334.050 ;
        RECT 58.950 331.950 61.050 334.050 ;
        RECT 65.400 332.100 66.300 340.350 ;
        RECT 77.400 338.100 78.600 342.300 ;
        RECT 97.950 341.400 99.750 342.300 ;
        RECT 82.950 339.450 85.050 340.200 ;
        RECT 94.950 339.450 97.050 340.050 ;
        RECT 82.950 338.550 97.050 339.450 ;
        RECT 82.950 338.100 85.050 338.550 ;
        RECT 94.950 337.950 97.050 338.550 ;
        RECT 76.950 336.450 79.050 337.050 ;
        RECT 81.000 336.900 84.000 337.050 ;
        RECT 81.000 336.450 85.050 336.900 ;
        RECT 76.950 335.550 85.050 336.450 ;
        RECT 95.100 336.150 96.900 336.900 ;
        RECT 76.950 334.950 79.050 335.550 ;
        RECT 81.000 334.950 85.050 335.550 ;
        RECT 92.100 335.100 93.900 335.850 ;
        RECT 82.950 334.800 85.050 334.950 ;
        RECT 74.100 332.100 75.900 332.850 ;
        RECT 59.100 330.150 60.900 330.900 ;
        RECT 56.100 329.100 57.900 329.850 ;
        RECT 64.950 328.950 67.050 331.050 ;
        RECT 73.950 328.950 76.050 331.050 ;
        RECT 10.800 315.600 12.600 321.600 ;
        RECT 25.800 315.600 27.600 321.600 ;
        RECT 40.800 315.600 42.600 327.600 ;
        RECT 43.800 326.700 51.600 327.600 ;
        RECT 43.800 315.600 45.600 326.700 ;
        RECT 49.800 315.600 51.600 326.700 ;
        RECT 55.950 325.950 58.050 328.050 ;
        RECT 65.400 322.800 66.300 327.900 ;
        RECT 74.550 327.000 75.450 328.950 ;
        RECT 73.950 322.950 76.050 327.000 ;
        RECT 59.700 321.900 66.300 322.800 ;
        RECT 59.700 321.600 61.200 321.900 ;
        RECT 59.400 315.600 61.200 321.600 ;
        RECT 65.400 321.600 66.300 321.900 ;
        RECT 77.400 321.600 78.600 333.900 ;
        RECT 80.100 332.100 81.900 332.850 ;
        RECT 91.950 331.950 94.050 334.050 ;
        RECT 79.950 328.950 82.050 331.050 ;
        RECT 98.700 330.600 99.600 341.400 ;
        RECT 102.000 338.100 103.050 344.400 ;
        RECT 119.100 342.000 120.900 350.400 ;
        RECT 138.000 343.200 139.800 350.400 ;
        RECT 149.400 345.300 151.200 350.400 ;
        RECT 155.400 345.300 157.200 350.400 ;
        RECT 149.400 343.950 157.200 345.300 ;
        RECT 158.400 344.400 160.200 350.400 ;
        RECT 172.500 344.400 174.300 350.400 ;
        RECT 178.800 347.400 180.600 350.400 ;
        RECT 187.800 349.500 195.600 350.400 ;
        RECT 138.000 342.300 141.600 343.200 ;
        RECT 158.400 342.300 159.600 344.400 ;
        RECT 116.700 340.350 120.900 342.000 ;
        RECT 100.950 336.450 103.050 337.050 ;
        RECT 109.950 336.450 112.050 337.050 ;
        RECT 100.950 335.550 112.050 336.450 ;
        RECT 100.950 334.950 103.050 335.550 ;
        RECT 109.950 334.950 112.050 335.550 ;
        RECT 97.800 330.000 99.600 330.600 ;
        RECT 92.400 328.800 99.600 330.000 ;
        RECT 92.400 327.600 93.600 328.800 ;
        RECT 100.950 327.600 102.300 333.900 ;
        RECT 116.700 332.100 117.600 340.350 ;
        RECT 119.100 338.100 120.900 338.850 ;
        RECT 140.400 338.100 141.600 342.300 ;
        RECT 155.850 341.250 159.600 342.300 ;
        RECT 155.850 341.100 157.050 341.250 ;
        RECT 172.800 341.100 174.000 344.400 ;
        RECT 178.800 343.500 180.000 347.400 ;
        RECT 187.800 344.400 189.600 349.500 ;
        RECT 190.800 344.400 192.600 348.600 ;
        RECT 193.800 345.000 195.600 349.500 ;
        RECT 199.800 345.000 201.600 350.400 ;
        RECT 174.900 342.600 180.000 343.500 ;
        RECT 191.400 342.900 192.300 344.400 ;
        RECT 193.800 344.100 201.600 345.000 ;
        RECT 204.150 344.400 205.950 350.400 ;
        RECT 211.950 348.300 213.750 350.400 ;
        RECT 210.000 347.400 213.750 348.300 ;
        RECT 219.750 347.400 221.550 350.400 ;
        RECT 227.550 347.400 229.350 350.400 ;
        RECT 210.000 346.500 211.050 347.400 ;
        RECT 208.950 344.400 211.050 346.500 ;
        RECT 219.750 345.600 220.800 347.400 ;
        RECT 174.900 341.700 176.850 342.600 ;
        RECT 191.400 341.700 195.600 342.900 ;
        RECT 175.950 341.100 176.850 341.700 ;
        RECT 194.400 341.100 195.600 341.700 ;
        RECT 199.950 341.100 201.750 341.850 ;
        RECT 148.950 337.950 151.050 340.050 ;
        RECT 154.950 337.950 157.050 340.050 ;
        RECT 172.950 337.950 175.050 340.050 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 133.950 336.450 138.000 337.050 ;
        RECT 139.950 336.450 142.050 337.050 ;
        RECT 176.100 336.900 176.850 341.100 ;
        RECT 133.950 335.550 142.050 336.450 ;
        RECT 149.100 336.150 150.900 336.900 ;
        RECT 133.950 334.950 138.000 335.550 ;
        RECT 139.950 334.950 142.050 335.550 ;
        RECT 152.100 335.100 153.900 335.850 ;
        RECT 154.950 335.100 156.150 336.900 ;
        RECT 158.100 335.100 159.900 335.850 ;
        RECT 121.950 331.950 124.050 334.050 ;
        RECT 137.100 332.100 138.900 332.850 ;
        RECT 115.950 328.950 118.050 331.050 ;
        RECT 122.100 330.150 123.900 330.900 ;
        RECT 125.100 329.100 126.900 329.850 ;
        RECT 136.950 328.950 139.050 331.050 ;
        RECT 65.400 315.600 67.200 321.600 ;
        RECT 77.400 315.600 79.200 321.600 ;
        RECT 92.400 315.600 94.200 327.600 ;
        RECT 99.900 326.100 102.300 327.600 ;
        RECT 99.900 315.600 101.700 326.100 ;
        RECT 116.700 322.800 117.600 327.900 ;
        RECT 124.950 325.950 127.050 328.050 ;
        RECT 116.700 321.900 123.300 322.800 ;
        RECT 116.700 321.600 117.600 321.900 ;
        RECT 115.800 315.600 117.600 321.600 ;
        RECT 121.800 321.600 123.300 321.900 ;
        RECT 140.400 321.600 141.600 333.900 ;
        RECT 143.100 332.100 144.900 332.850 ;
        RECT 151.950 331.950 154.050 334.050 ;
        RECT 142.950 328.950 145.050 331.050 ;
        RECT 155.100 330.900 156.150 335.100 ;
        RECT 157.950 331.950 160.050 334.050 ;
        RECT 154.950 327.600 156.150 330.900 ;
        RECT 172.800 327.600 174.000 336.900 ;
        RECT 175.950 330.300 176.850 336.900 ;
        RECT 178.950 334.950 181.050 340.050 ;
        RECT 187.950 337.950 190.050 340.050 ;
        RECT 193.950 337.950 196.050 340.050 ;
        RECT 199.950 337.950 202.050 340.050 ;
        RECT 188.250 336.150 190.050 336.900 ;
        RECT 191.700 335.100 193.500 335.850 ;
        RECT 179.100 333.150 180.900 333.900 ;
        RECT 190.950 331.950 193.050 334.050 ;
        RECT 174.900 329.400 176.850 330.300 ;
        RECT 174.900 328.500 180.600 329.400 ;
        RECT 121.800 315.600 123.600 321.600 ;
        RECT 139.800 315.600 141.600 321.600 ;
        RECT 154.500 315.600 156.300 327.600 ;
        RECT 172.500 315.600 174.300 327.600 ;
        RECT 179.400 321.600 180.600 328.500 ;
        RECT 194.400 327.600 195.600 336.900 ;
        RECT 197.100 335.100 198.900 335.850 ;
        RECT 196.950 331.950 199.050 334.050 ;
        RECT 204.150 329.700 205.050 344.400 ;
        RECT 212.550 343.800 214.350 345.600 ;
        RECT 215.850 344.550 220.800 345.600 ;
        RECT 228.300 346.500 229.350 347.400 ;
        RECT 228.300 345.300 232.050 346.500 ;
        RECT 215.850 343.800 217.650 344.550 ;
        RECT 229.950 344.400 232.050 345.300 ;
        RECT 235.650 344.400 237.450 350.400 ;
        RECT 212.850 340.800 213.900 343.800 ;
        RECT 207.000 339.600 224.850 340.800 ;
        RECT 236.250 340.050 237.450 344.400 ;
        RECT 245.400 347.400 247.200 350.400 ;
        RECT 262.800 347.400 264.600 350.400 ;
        RECT 277.800 347.400 279.600 350.400 ;
        RECT 207.000 338.850 207.900 339.600 ;
        RECT 212.100 339.000 213.900 339.600 ;
        RECT 223.050 339.000 224.850 339.600 ;
        RECT 206.100 337.050 207.900 338.850 ;
        RECT 223.050 338.100 223.950 339.000 ;
        RECT 231.150 338.250 231.900 340.050 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 236.100 337.950 237.450 340.050 ;
        RECT 238.950 337.950 244.050 340.050 ;
        RECT 209.100 334.800 210.900 335.400 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 209.100 333.600 213.900 334.800 ;
        RECT 214.950 331.950 217.050 334.050 ;
        RECT 213.450 329.700 215.250 330.000 ;
        RECT 204.150 329.100 215.250 329.700 ;
        RECT 204.150 328.500 221.850 329.100 ;
        RECT 204.150 327.600 205.050 328.500 ;
        RECT 213.450 328.200 221.850 328.500 ;
        RECT 178.800 315.600 180.600 321.600 ;
        RECT 193.800 315.600 197.100 327.600 ;
        RECT 204.150 315.600 205.950 327.600 ;
        RECT 218.250 326.700 220.050 327.300 ;
        RECT 212.550 325.500 220.050 326.700 ;
        RECT 220.950 326.100 221.850 328.200 ;
        RECT 223.050 328.200 223.950 333.900 ;
        RECT 233.250 329.400 235.050 331.200 ;
        RECT 229.950 328.200 234.150 329.400 ;
        RECT 223.050 327.300 229.050 328.200 ;
        RECT 229.950 327.300 232.050 328.200 ;
        RECT 236.250 327.600 237.450 337.950 ;
        RECT 242.100 336.150 243.900 336.900 ;
        RECT 245.400 335.100 246.600 347.400 ;
        RECT 263.400 344.100 264.600 347.400 ;
        RECT 262.950 340.950 268.050 343.050 ;
        RECT 262.950 338.100 264.300 339.900 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 244.950 331.950 247.050 334.050 ;
        RECT 263.100 333.900 264.300 338.100 ;
        RECT 260.100 333.150 261.900 333.900 ;
        RECT 228.150 326.400 229.050 327.300 ;
        RECT 225.450 326.100 227.250 326.400 ;
        RECT 212.550 324.600 213.750 325.500 ;
        RECT 220.950 325.200 227.250 326.100 ;
        RECT 225.450 324.600 227.250 325.200 ;
        RECT 228.150 324.600 230.850 326.400 ;
        RECT 208.950 322.500 213.750 324.600 ;
        RECT 216.450 323.550 218.250 324.300 ;
        RECT 221.250 323.550 223.050 324.300 ;
        RECT 216.450 322.500 223.050 323.550 ;
        RECT 212.550 321.600 213.750 322.500 ;
        RECT 212.550 315.600 214.350 321.600 ;
        RECT 220.350 315.600 222.150 322.500 ;
        RECT 228.150 321.600 232.050 323.700 ;
        RECT 228.150 315.600 229.950 321.600 ;
        RECT 235.650 315.600 237.450 327.600 ;
        RECT 245.400 321.600 246.600 330.900 ;
        RECT 262.950 328.650 264.300 333.900 ;
        RECT 265.950 333.450 268.050 334.050 ;
        RECT 271.950 333.450 274.050 337.050 ;
        RECT 278.400 335.100 279.600 347.400 ;
        RECT 284.550 344.400 286.350 350.400 ;
        RECT 292.650 347.400 294.450 350.400 ;
        RECT 300.450 347.400 302.250 350.400 ;
        RECT 308.250 348.300 310.050 350.400 ;
        RECT 308.250 347.400 312.000 348.300 ;
        RECT 292.650 346.500 293.700 347.400 ;
        RECT 289.950 345.300 293.700 346.500 ;
        RECT 301.200 345.600 302.250 347.400 ;
        RECT 310.950 346.500 312.000 347.400 ;
        RECT 289.950 344.400 292.050 345.300 ;
        RECT 301.200 344.550 306.150 345.600 ;
        RECT 284.550 340.050 285.750 344.400 ;
        RECT 304.350 343.800 306.150 344.550 ;
        RECT 307.650 343.800 309.450 345.600 ;
        RECT 310.950 344.400 313.050 346.500 ;
        RECT 316.050 344.400 317.850 350.400 ;
        RECT 328.800 344.400 330.600 350.400 ;
        RECT 308.100 340.800 309.150 343.800 ;
        RECT 280.950 337.950 283.050 340.050 ;
        RECT 284.550 337.950 285.900 340.050 ;
        RECT 286.950 337.950 289.050 340.050 ;
        RECT 290.100 338.250 290.850 340.050 ;
        RECT 297.150 339.600 315.000 340.800 ;
        RECT 297.150 339.000 298.950 339.600 ;
        RECT 308.100 339.000 309.900 339.600 ;
        RECT 298.050 338.100 298.950 339.000 ;
        RECT 314.100 338.850 315.000 339.600 ;
        RECT 281.100 336.150 282.900 336.900 ;
        RECT 265.950 333.000 274.050 333.450 ;
        RECT 265.950 332.550 273.450 333.000 ;
        RECT 265.950 331.950 268.050 332.550 ;
        RECT 277.950 331.950 280.050 334.050 ;
        RECT 266.100 330.150 267.900 330.900 ;
        RECT 261.600 327.600 264.300 328.650 ;
        RECT 245.400 315.600 247.200 321.600 ;
        RECT 261.600 315.600 263.400 327.600 ;
        RECT 278.400 321.600 279.600 330.900 ;
        RECT 277.800 315.600 279.600 321.600 ;
        RECT 284.550 327.600 285.750 337.950 ;
        RECT 314.100 337.050 315.900 338.850 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 286.950 329.400 288.750 331.200 ;
        RECT 287.850 328.200 292.050 329.400 ;
        RECT 298.050 328.200 298.950 333.900 ;
        RECT 304.950 331.950 307.050 337.050 ;
        RECT 311.100 334.800 312.900 335.400 ;
        RECT 308.100 333.600 312.900 334.800 ;
        RECT 306.750 329.700 308.550 330.000 ;
        RECT 316.950 329.700 317.850 344.400 ;
        RECT 329.400 342.300 330.600 344.400 ;
        RECT 331.800 345.300 333.600 350.400 ;
        RECT 337.800 345.300 339.600 350.400 ;
        RECT 331.800 343.950 339.600 345.300 ;
        RECT 349.500 344.400 351.300 350.400 ;
        RECT 355.800 347.400 357.600 350.400 ;
        RECT 329.400 341.250 333.150 342.300 ;
        RECT 331.950 341.100 333.150 341.250 ;
        RECT 331.950 337.950 334.050 340.050 ;
        RECT 337.950 337.950 340.050 340.050 ;
        RECT 343.950 339.450 346.050 343.050 ;
        RECT 349.800 341.100 351.000 344.400 ;
        RECT 355.800 343.500 357.000 347.400 ;
        RECT 351.900 342.600 357.000 343.500 ;
        RECT 367.200 343.200 369.000 350.400 ;
        RECT 351.900 341.700 353.850 342.600 ;
        RECT 352.950 341.100 353.850 341.700 ;
        RECT 349.950 339.450 352.050 340.050 ;
        RECT 343.950 339.000 352.050 339.450 ;
        RECT 344.550 338.550 352.050 339.000 ;
        RECT 349.950 337.950 352.050 338.550 ;
        RECT 353.100 336.900 353.850 341.100 ;
        RECT 365.400 342.300 369.000 343.200 ;
        RECT 374.550 344.400 376.350 350.400 ;
        RECT 382.650 347.400 384.450 350.400 ;
        RECT 390.450 347.400 392.250 350.400 ;
        RECT 398.250 348.300 400.050 350.400 ;
        RECT 398.250 347.400 402.000 348.300 ;
        RECT 382.650 346.500 383.700 347.400 ;
        RECT 379.950 345.300 383.700 346.500 ;
        RECT 391.200 345.600 392.250 347.400 ;
        RECT 400.950 346.500 402.000 347.400 ;
        RECT 379.950 344.400 382.050 345.300 ;
        RECT 391.200 344.550 396.150 345.600 ;
        RECT 365.400 338.100 366.600 342.300 ;
        RECT 374.550 340.050 375.750 344.400 ;
        RECT 394.350 343.800 396.150 344.550 ;
        RECT 397.650 343.800 399.450 345.600 ;
        RECT 400.950 344.400 403.050 346.500 ;
        RECT 406.050 344.400 407.850 350.400 ;
        RECT 398.100 340.800 399.150 343.800 ;
        RECT 374.550 337.950 375.900 340.050 ;
        RECT 376.950 337.950 379.050 340.050 ;
        RECT 380.100 338.250 380.850 340.050 ;
        RECT 387.150 339.600 405.000 340.800 ;
        RECT 387.150 339.000 388.950 339.600 ;
        RECT 398.100 339.000 399.900 339.600 ;
        RECT 388.050 338.100 388.950 339.000 ;
        RECT 404.100 338.850 405.000 339.600 ;
        RECT 329.100 335.100 330.900 335.850 ;
        RECT 332.850 335.100 334.050 336.900 ;
        RECT 338.100 336.150 339.900 336.900 ;
        RECT 335.100 335.100 336.900 335.850 ;
        RECT 328.950 331.950 331.050 334.050 ;
        RECT 306.750 329.100 317.850 329.700 ;
        RECT 284.550 315.600 286.350 327.600 ;
        RECT 289.950 327.300 292.050 328.200 ;
        RECT 292.950 327.300 298.950 328.200 ;
        RECT 300.150 328.500 317.850 329.100 ;
        RECT 300.150 328.200 308.550 328.500 ;
        RECT 292.950 326.400 293.850 327.300 ;
        RECT 291.150 324.600 293.850 326.400 ;
        RECT 294.750 326.100 296.550 326.400 ;
        RECT 300.150 326.100 301.050 328.200 ;
        RECT 316.950 327.600 317.850 328.500 ;
        RECT 332.850 330.900 333.900 335.100 ;
        RECT 334.950 331.950 337.050 334.050 ;
        RECT 332.850 327.600 334.050 330.900 ;
        RECT 349.800 327.600 351.000 336.900 ;
        RECT 352.950 330.300 353.850 336.900 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 361.950 334.950 367.050 337.050 ;
        RECT 356.100 333.150 357.900 333.900 ;
        RECT 362.100 332.100 363.900 332.850 ;
        RECT 351.900 329.400 353.850 330.300 ;
        RECT 351.900 328.500 357.600 329.400 ;
        RECT 361.950 328.950 364.050 331.050 ;
        RECT 294.750 325.200 301.050 326.100 ;
        RECT 301.950 326.700 303.750 327.300 ;
        RECT 301.950 325.500 309.450 326.700 ;
        RECT 294.750 324.600 296.550 325.200 ;
        RECT 308.250 324.600 309.450 325.500 ;
        RECT 289.950 321.600 293.850 323.700 ;
        RECT 298.950 323.550 300.750 324.300 ;
        RECT 303.750 323.550 305.550 324.300 ;
        RECT 298.950 322.500 305.550 323.550 ;
        RECT 308.250 322.500 313.050 324.600 ;
        RECT 292.050 315.600 293.850 321.600 ;
        RECT 299.850 315.600 301.650 322.500 ;
        RECT 308.250 321.600 309.450 322.500 ;
        RECT 307.650 315.600 309.450 321.600 ;
        RECT 316.050 315.600 317.850 327.600 ;
        RECT 332.700 315.600 334.500 327.600 ;
        RECT 349.500 315.600 351.300 327.600 ;
        RECT 356.400 321.600 357.600 328.500 ;
        RECT 355.800 315.600 357.600 321.600 ;
        RECT 365.400 321.600 366.600 333.900 ;
        RECT 368.100 332.100 369.900 332.850 ;
        RECT 367.950 328.950 370.050 331.050 ;
        RECT 374.550 327.600 375.750 337.950 ;
        RECT 404.100 337.050 405.900 338.850 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 401.100 334.800 402.900 335.400 ;
        RECT 376.950 329.400 378.750 331.200 ;
        RECT 377.850 328.200 382.050 329.400 ;
        RECT 388.050 328.200 388.950 333.900 ;
        RECT 394.950 331.950 397.050 334.050 ;
        RECT 398.100 333.600 402.900 334.800 ;
        RECT 396.750 329.700 398.550 330.000 ;
        RECT 406.950 329.700 407.850 344.400 ;
        RECT 396.750 329.100 407.850 329.700 ;
        RECT 365.400 315.600 367.200 321.600 ;
        RECT 374.550 315.600 376.350 327.600 ;
        RECT 379.950 327.300 382.050 328.200 ;
        RECT 382.950 327.300 388.950 328.200 ;
        RECT 390.150 328.500 407.850 329.100 ;
        RECT 390.150 328.200 398.550 328.500 ;
        RECT 382.950 326.400 383.850 327.300 ;
        RECT 381.150 324.600 383.850 326.400 ;
        RECT 384.750 326.100 386.550 326.400 ;
        RECT 390.150 326.100 391.050 328.200 ;
        RECT 406.950 327.600 407.850 328.500 ;
        RECT 384.750 325.200 391.050 326.100 ;
        RECT 391.950 326.700 393.750 327.300 ;
        RECT 391.950 325.500 399.450 326.700 ;
        RECT 384.750 324.600 386.550 325.200 ;
        RECT 398.250 324.600 399.450 325.500 ;
        RECT 379.950 321.600 383.850 323.700 ;
        RECT 388.950 323.550 390.750 324.300 ;
        RECT 393.750 323.550 395.550 324.300 ;
        RECT 388.950 322.500 395.550 323.550 ;
        RECT 398.250 322.500 403.050 324.600 ;
        RECT 382.050 315.600 383.850 321.600 ;
        RECT 389.850 315.600 391.650 322.500 ;
        RECT 398.250 321.600 399.450 322.500 ;
        RECT 397.650 315.600 399.450 321.600 ;
        RECT 406.050 315.600 407.850 327.600 ;
        RECT 411.150 344.400 412.950 350.400 ;
        RECT 418.950 348.300 420.750 350.400 ;
        RECT 417.000 347.400 420.750 348.300 ;
        RECT 426.750 347.400 428.550 350.400 ;
        RECT 434.550 347.400 436.350 350.400 ;
        RECT 417.000 346.500 418.050 347.400 ;
        RECT 415.950 344.400 418.050 346.500 ;
        RECT 426.750 345.600 427.800 347.400 ;
        RECT 411.150 329.700 412.050 344.400 ;
        RECT 419.550 343.800 421.350 345.600 ;
        RECT 422.850 344.550 427.800 345.600 ;
        RECT 435.300 346.500 436.350 347.400 ;
        RECT 435.300 345.300 439.050 346.500 ;
        RECT 422.850 343.800 424.650 344.550 ;
        RECT 436.950 344.400 439.050 345.300 ;
        RECT 442.650 344.400 444.450 350.400 ;
        RECT 456.000 346.050 457.800 350.400 ;
        RECT 419.850 340.800 420.900 343.800 ;
        RECT 414.000 339.600 431.850 340.800 ;
        RECT 443.250 340.050 444.450 344.400 ;
        RECT 452.400 344.400 457.800 346.050 ;
        RECT 473.400 347.400 475.200 350.400 ;
        RECT 493.800 347.400 495.600 350.400 ;
        RECT 452.400 341.100 453.300 344.400 ;
        RECT 473.400 344.100 474.600 347.400 ;
        RECT 494.400 344.100 495.600 347.400 ;
        RECT 510.000 343.200 511.800 350.400 ;
        RECT 526.800 344.400 528.600 350.400 ;
        RECT 466.950 342.450 471.000 343.050 ;
        RECT 472.950 342.450 475.050 343.050 ;
        RECT 466.950 341.550 475.050 342.450 ;
        RECT 466.950 340.950 471.000 341.550 ;
        RECT 472.950 340.950 475.050 341.550 ;
        RECT 478.950 342.450 481.050 343.050 ;
        RECT 493.950 342.450 496.050 343.050 ;
        RECT 478.950 341.550 496.050 342.450 ;
        RECT 510.000 342.300 513.600 343.200 ;
        RECT 478.950 340.950 481.050 341.550 ;
        RECT 493.950 340.950 496.050 341.550 ;
        RECT 414.000 338.850 414.900 339.600 ;
        RECT 419.100 339.000 420.900 339.600 ;
        RECT 430.050 339.000 431.850 339.600 ;
        RECT 413.100 337.050 414.900 338.850 ;
        RECT 430.050 338.100 430.950 339.000 ;
        RECT 438.150 338.250 438.900 340.050 ;
        RECT 439.950 337.950 442.050 340.050 ;
        RECT 443.100 337.950 444.450 340.050 ;
        RECT 445.950 339.450 450.000 340.050 ;
        RECT 451.950 339.450 454.050 340.050 ;
        RECT 445.950 338.550 454.050 339.450 ;
        RECT 445.950 337.950 450.000 338.550 ;
        RECT 451.950 337.950 454.050 338.550 ;
        RECT 457.950 337.950 460.050 340.050 ;
        RECT 473.700 338.100 475.050 339.900 ;
        RECT 493.950 338.100 495.300 339.900 ;
        RECT 512.400 338.100 513.600 342.300 ;
        RECT 527.400 342.300 528.600 344.400 ;
        RECT 529.800 345.300 531.600 350.400 ;
        RECT 535.800 345.300 537.600 350.400 ;
        RECT 544.800 347.400 546.600 350.400 ;
        RECT 529.800 343.950 537.600 345.300 ;
        RECT 527.400 341.250 531.150 342.300 ;
        RECT 529.950 341.100 531.150 341.250 ;
        RECT 416.100 334.800 417.900 335.400 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 416.100 333.600 420.900 334.800 ;
        RECT 421.950 331.950 424.050 334.050 ;
        RECT 420.450 329.700 422.250 330.000 ;
        RECT 411.150 329.100 422.250 329.700 ;
        RECT 411.150 328.500 428.850 329.100 ;
        RECT 411.150 327.600 412.050 328.500 ;
        RECT 420.450 328.200 428.850 328.500 ;
        RECT 411.150 315.600 412.950 327.600 ;
        RECT 425.250 326.700 427.050 327.300 ;
        RECT 419.550 325.500 427.050 326.700 ;
        RECT 427.950 326.100 428.850 328.200 ;
        RECT 430.050 328.200 430.950 333.900 ;
        RECT 440.250 329.400 442.050 331.200 ;
        RECT 436.950 328.200 441.150 329.400 ;
        RECT 430.050 327.300 436.050 328.200 ;
        RECT 436.950 327.300 439.050 328.200 ;
        RECT 443.250 327.600 444.450 337.950 ;
        RECT 452.400 327.600 453.300 336.900 ;
        RECT 458.100 336.150 459.900 336.900 ;
        RECT 455.100 335.100 456.900 335.850 ;
        RECT 461.100 335.100 462.900 335.850 ;
        RECT 454.950 331.950 457.050 334.050 ;
        RECT 460.950 331.950 463.050 334.050 ;
        RECT 469.950 331.950 472.050 334.050 ;
        RECT 473.700 333.900 474.900 338.100 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 490.950 334.950 493.050 337.050 ;
        RECT 494.100 333.900 495.300 338.100 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 535.950 337.950 538.050 340.050 ;
        RECT 470.100 330.150 471.900 330.900 ;
        RECT 473.700 328.650 475.050 333.900 ;
        RECT 476.100 333.150 477.900 333.900 ;
        RECT 491.100 333.150 492.900 333.900 ;
        RECT 493.950 328.650 495.300 333.900 ;
        RECT 496.950 331.950 499.050 337.050 ;
        RECT 511.950 336.450 514.050 337.050 ;
        RECT 520.950 336.450 523.050 337.050 ;
        RECT 511.950 335.550 523.050 336.450 ;
        RECT 511.950 334.950 514.050 335.550 ;
        RECT 520.950 334.950 523.050 335.550 ;
        RECT 527.100 335.100 528.900 335.850 ;
        RECT 530.850 335.100 532.050 336.900 ;
        RECT 536.100 336.150 537.900 336.900 ;
        RECT 533.100 335.100 534.900 335.850 ;
        RECT 545.400 335.100 546.600 347.400 ;
        RECT 552.150 344.400 553.950 350.400 ;
        RECT 559.950 348.300 561.750 350.400 ;
        RECT 558.000 347.400 561.750 348.300 ;
        RECT 567.750 347.400 569.550 350.400 ;
        RECT 575.550 347.400 577.350 350.400 ;
        RECT 558.000 346.500 559.050 347.400 ;
        RECT 556.950 344.400 559.050 346.500 ;
        RECT 567.750 345.600 568.800 347.400 ;
        RECT 547.950 337.950 550.050 340.050 ;
        RECT 548.100 336.150 549.900 336.900 ;
        RECT 509.100 332.100 510.900 332.850 ;
        RECT 497.100 330.150 498.900 330.900 ;
        RECT 508.950 328.950 511.050 331.050 ;
        RECT 473.700 327.600 476.400 328.650 ;
        RECT 435.150 326.400 436.050 327.300 ;
        RECT 432.450 326.100 434.250 326.400 ;
        RECT 419.550 324.600 420.750 325.500 ;
        RECT 427.950 325.200 434.250 326.100 ;
        RECT 432.450 324.600 434.250 325.200 ;
        RECT 435.150 324.600 437.850 326.400 ;
        RECT 415.950 322.500 420.750 324.600 ;
        RECT 423.450 323.550 425.250 324.300 ;
        RECT 428.250 323.550 430.050 324.300 ;
        RECT 423.450 322.500 430.050 323.550 ;
        RECT 419.550 321.600 420.750 322.500 ;
        RECT 419.550 315.600 421.350 321.600 ;
        RECT 427.350 315.600 429.150 322.500 ;
        RECT 435.150 321.600 439.050 323.700 ;
        RECT 435.150 315.600 436.950 321.600 ;
        RECT 442.650 315.600 444.450 327.600 ;
        RECT 451.800 315.600 453.600 327.600 ;
        RECT 454.800 326.700 462.600 327.600 ;
        RECT 454.800 315.600 456.600 326.700 ;
        RECT 460.800 315.600 462.600 326.700 ;
        RECT 474.600 315.600 476.400 327.600 ;
        RECT 492.600 327.600 495.300 328.650 ;
        RECT 492.600 315.600 494.400 327.600 ;
        RECT 512.400 321.600 513.600 333.900 ;
        RECT 515.100 332.100 516.900 332.850 ;
        RECT 526.950 331.950 529.050 334.050 ;
        RECT 514.950 328.950 517.050 331.050 ;
        RECT 530.850 330.900 531.900 335.100 ;
        RECT 532.950 331.950 535.050 334.050 ;
        RECT 544.950 331.950 547.050 334.050 ;
        RECT 530.850 327.600 532.050 330.900 ;
        RECT 511.800 315.600 513.600 321.600 ;
        RECT 530.700 315.600 532.500 327.600 ;
        RECT 545.400 321.600 546.600 330.900 ;
        RECT 544.800 315.600 546.600 321.600 ;
        RECT 552.150 329.700 553.050 344.400 ;
        RECT 560.550 343.800 562.350 345.600 ;
        RECT 563.850 344.550 568.800 345.600 ;
        RECT 576.300 346.500 577.350 347.400 ;
        RECT 576.300 345.300 580.050 346.500 ;
        RECT 563.850 343.800 565.650 344.550 ;
        RECT 577.950 344.400 580.050 345.300 ;
        RECT 583.650 344.400 585.450 350.400 ;
        RECT 560.850 340.800 561.900 343.800 ;
        RECT 555.000 339.600 572.850 340.800 ;
        RECT 584.250 340.050 585.450 344.400 ;
        RECT 596.400 347.400 598.200 350.400 ;
        RECT 596.400 344.100 597.600 347.400 ;
        RECT 615.000 343.200 616.800 350.400 ;
        RECT 633.000 343.200 634.800 350.400 ;
        RECT 647.400 347.400 649.200 350.400 ;
        RECT 648.000 343.500 649.200 347.400 ;
        RECT 653.700 344.400 655.500 350.400 ;
        RECT 664.800 344.400 666.600 350.400 ;
        RECT 595.950 342.450 598.050 343.050 ;
        RECT 604.950 342.450 607.050 343.050 ;
        RECT 595.950 341.550 607.050 342.450 ;
        RECT 615.000 342.300 618.600 343.200 ;
        RECT 633.000 342.300 636.600 343.200 ;
        RECT 648.000 342.600 653.100 343.500 ;
        RECT 595.950 340.950 598.050 341.550 ;
        RECT 604.950 340.950 607.050 341.550 ;
        RECT 555.000 338.850 555.900 339.600 ;
        RECT 560.100 339.000 561.900 339.600 ;
        RECT 571.050 339.000 572.850 339.600 ;
        RECT 554.100 337.050 555.900 338.850 ;
        RECT 571.050 338.100 571.950 339.000 ;
        RECT 579.150 338.250 579.900 340.050 ;
        RECT 580.950 337.950 583.050 340.050 ;
        RECT 584.100 337.950 585.450 340.050 ;
        RECT 557.100 334.800 558.900 335.400 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 557.100 333.600 561.900 334.800 ;
        RECT 562.950 331.950 565.050 334.050 ;
        RECT 561.450 329.700 563.250 330.000 ;
        RECT 552.150 329.100 563.250 329.700 ;
        RECT 552.150 328.500 569.850 329.100 ;
        RECT 552.150 327.600 553.050 328.500 ;
        RECT 561.450 328.200 569.850 328.500 ;
        RECT 552.150 315.600 553.950 327.600 ;
        RECT 566.250 326.700 568.050 327.300 ;
        RECT 560.550 325.500 568.050 326.700 ;
        RECT 568.950 326.100 569.850 328.200 ;
        RECT 571.050 328.200 571.950 333.900 ;
        RECT 581.250 329.400 583.050 331.200 ;
        RECT 577.950 328.200 582.150 329.400 ;
        RECT 571.050 327.300 577.050 328.200 ;
        RECT 577.950 327.300 580.050 328.200 ;
        RECT 584.250 327.600 585.450 337.950 ;
        RECT 596.700 338.100 598.050 339.900 ;
        RECT 617.400 338.100 618.600 342.300 ;
        RECT 635.400 338.100 636.600 342.300 ;
        RECT 651.150 341.700 653.100 342.600 ;
        RECT 651.150 341.100 652.050 341.700 ;
        RECT 654.000 341.100 655.200 344.400 ;
        RECT 665.400 342.300 666.600 344.400 ;
        RECT 667.800 345.300 669.600 350.400 ;
        RECT 673.800 345.300 675.600 350.400 ;
        RECT 667.800 343.950 675.600 345.300 ;
        RECT 678.150 344.400 679.950 350.400 ;
        RECT 685.950 348.300 687.750 350.400 ;
        RECT 684.000 347.400 687.750 348.300 ;
        RECT 693.750 347.400 695.550 350.400 ;
        RECT 701.550 347.400 703.350 350.400 ;
        RECT 684.000 346.500 685.050 347.400 ;
        RECT 682.950 344.400 685.050 346.500 ;
        RECT 693.750 345.600 694.800 347.400 ;
        RECT 665.400 341.250 669.150 342.300 ;
        RECT 667.950 341.100 669.150 341.250 ;
        RECT 586.950 333.450 591.000 334.050 ;
        RECT 592.950 333.450 595.050 334.050 ;
        RECT 586.950 332.550 595.050 333.450 ;
        RECT 586.950 331.950 591.000 332.550 ;
        RECT 592.950 331.950 595.050 332.550 ;
        RECT 596.700 333.900 597.900 338.100 ;
        RECT 619.950 337.050 622.050 337.200 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 616.950 335.100 622.050 337.050 ;
        RECT 634.950 336.450 637.050 337.050 ;
        RECT 639.000 336.450 643.050 337.050 ;
        RECT 634.950 335.550 643.050 336.450 ;
        RECT 616.950 334.950 621.450 335.100 ;
        RECT 634.950 334.950 637.050 335.550 ;
        RECT 639.000 334.950 643.050 335.550 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 651.150 336.900 651.900 341.100 ;
        RECT 652.950 339.450 655.050 340.050 ;
        RECT 657.000 339.450 661.050 340.050 ;
        RECT 652.950 338.550 661.050 339.450 ;
        RECT 652.950 337.950 655.050 338.550 ;
        RECT 657.000 337.950 661.050 338.550 ;
        RECT 667.950 337.950 670.050 340.050 ;
        RECT 673.950 337.950 676.050 340.050 ;
        RECT 593.100 330.150 594.900 330.900 ;
        RECT 596.700 328.650 598.050 333.900 ;
        RECT 599.100 333.150 600.900 333.900 ;
        RECT 614.100 332.100 615.900 332.850 ;
        RECT 613.950 328.950 616.050 331.050 ;
        RECT 596.700 327.600 599.400 328.650 ;
        RECT 576.150 326.400 577.050 327.300 ;
        RECT 573.450 326.100 575.250 326.400 ;
        RECT 560.550 324.600 561.750 325.500 ;
        RECT 568.950 325.200 575.250 326.100 ;
        RECT 573.450 324.600 575.250 325.200 ;
        RECT 576.150 324.600 578.850 326.400 ;
        RECT 556.950 322.500 561.750 324.600 ;
        RECT 564.450 323.550 566.250 324.300 ;
        RECT 569.250 323.550 571.050 324.300 ;
        RECT 564.450 322.500 571.050 323.550 ;
        RECT 560.550 321.600 561.750 322.500 ;
        RECT 560.550 315.600 562.350 321.600 ;
        RECT 568.350 315.600 570.150 322.500 ;
        RECT 576.150 321.600 580.050 323.700 ;
        RECT 576.150 315.600 577.950 321.600 ;
        RECT 583.650 315.600 585.450 327.600 ;
        RECT 597.600 315.600 599.400 327.600 ;
        RECT 617.400 321.600 618.600 333.900 ;
        RECT 620.100 332.100 621.900 332.850 ;
        RECT 632.100 332.100 633.900 332.850 ;
        RECT 619.950 328.950 622.050 331.050 ;
        RECT 631.950 328.950 634.050 331.050 ;
        RECT 635.400 321.600 636.600 333.900 ;
        RECT 647.100 333.150 648.900 333.900 ;
        RECT 638.100 332.100 639.900 332.850 ;
        RECT 637.950 328.950 640.050 331.050 ;
        RECT 651.150 330.300 652.050 336.900 ;
        RECT 651.150 329.400 653.100 330.300 ;
        RECT 616.800 315.600 618.600 321.600 ;
        RECT 634.800 315.600 636.600 321.600 ;
        RECT 647.400 328.500 653.100 329.400 ;
        RECT 647.400 321.600 648.600 328.500 ;
        RECT 654.000 327.600 655.200 336.900 ;
        RECT 665.100 335.100 666.900 335.850 ;
        RECT 668.850 335.100 670.050 336.900 ;
        RECT 674.100 336.150 675.900 336.900 ;
        RECT 671.100 335.100 672.900 335.850 ;
        RECT 664.950 331.950 667.050 334.050 ;
        RECT 668.850 330.900 669.900 335.100 ;
        RECT 670.950 331.950 673.050 334.050 ;
        RECT 668.850 327.600 670.050 330.900 ;
        RECT 678.150 329.700 679.050 344.400 ;
        RECT 686.550 343.800 688.350 345.600 ;
        RECT 689.850 344.550 694.800 345.600 ;
        RECT 702.300 346.500 703.350 347.400 ;
        RECT 702.300 345.300 706.050 346.500 ;
        RECT 689.850 343.800 691.650 344.550 ;
        RECT 703.950 344.400 706.050 345.300 ;
        RECT 709.650 344.400 711.450 350.400 ;
        RECT 686.850 340.800 687.900 343.800 ;
        RECT 681.000 339.600 698.850 340.800 ;
        RECT 710.250 340.050 711.450 344.400 ;
        RECT 719.400 347.400 721.200 350.400 ;
        RECT 681.000 338.850 681.900 339.600 ;
        RECT 686.100 339.000 687.900 339.600 ;
        RECT 697.050 339.000 698.850 339.600 ;
        RECT 680.100 337.050 681.900 338.850 ;
        RECT 697.050 338.100 697.950 339.000 ;
        RECT 705.150 338.250 705.900 340.050 ;
        RECT 706.950 337.950 709.050 340.050 ;
        RECT 710.100 337.950 711.450 340.050 ;
        RECT 715.950 337.950 718.050 340.050 ;
        RECT 683.100 334.800 684.900 335.400 ;
        RECT 683.100 333.600 687.900 334.800 ;
        RECT 688.950 331.950 691.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 687.450 329.700 689.250 330.000 ;
        RECT 678.150 329.100 689.250 329.700 ;
        RECT 678.150 328.500 695.850 329.100 ;
        RECT 678.150 327.600 679.050 328.500 ;
        RECT 687.450 328.200 695.850 328.500 ;
        RECT 647.400 315.600 649.200 321.600 ;
        RECT 653.700 315.600 655.500 327.600 ;
        RECT 668.700 315.600 670.500 327.600 ;
        RECT 678.150 315.600 679.950 327.600 ;
        RECT 692.250 326.700 694.050 327.300 ;
        RECT 686.550 325.500 694.050 326.700 ;
        RECT 694.950 326.100 695.850 328.200 ;
        RECT 697.050 328.200 697.950 333.900 ;
        RECT 707.250 329.400 709.050 331.200 ;
        RECT 703.950 328.200 708.150 329.400 ;
        RECT 697.050 327.300 703.050 328.200 ;
        RECT 703.950 327.300 706.050 328.200 ;
        RECT 710.250 327.600 711.450 337.950 ;
        RECT 716.100 336.150 717.900 336.900 ;
        RECT 719.400 335.100 720.600 347.400 ;
        RECT 741.000 344.400 742.800 350.400 ;
        RECT 750.150 344.400 751.950 350.400 ;
        RECT 757.950 348.300 759.750 350.400 ;
        RECT 756.000 347.400 759.750 348.300 ;
        RECT 765.750 347.400 767.550 350.400 ;
        RECT 773.550 347.400 775.350 350.400 ;
        RECT 756.000 346.500 757.050 347.400 ;
        RECT 754.950 344.400 757.050 346.500 ;
        RECT 765.750 345.600 766.800 347.400 ;
        RECT 741.000 341.100 742.050 344.400 ;
        RECT 733.950 337.950 736.050 340.050 ;
        RECT 739.950 337.950 742.050 340.050 ;
        RECT 745.950 337.950 748.050 340.050 ;
        RECT 734.100 336.150 735.900 336.900 ;
        RECT 737.250 335.100 739.050 335.850 ;
        RECT 739.950 335.100 740.850 336.900 ;
        RECT 745.950 336.150 747.750 336.900 ;
        RECT 742.950 335.100 744.750 335.850 ;
        RECT 718.950 331.950 721.050 334.050 ;
        RECT 736.950 331.950 739.050 334.050 ;
        RECT 740.100 330.900 740.850 335.100 ;
        RECT 742.950 331.950 745.050 334.050 ;
        RECT 702.150 326.400 703.050 327.300 ;
        RECT 699.450 326.100 701.250 326.400 ;
        RECT 686.550 324.600 687.750 325.500 ;
        RECT 694.950 325.200 701.250 326.100 ;
        RECT 699.450 324.600 701.250 325.200 ;
        RECT 702.150 324.600 704.850 326.400 ;
        RECT 682.950 322.500 687.750 324.600 ;
        RECT 690.450 323.550 692.250 324.300 ;
        RECT 695.250 323.550 697.050 324.300 ;
        RECT 690.450 322.500 697.050 323.550 ;
        RECT 686.550 321.600 687.750 322.500 ;
        RECT 686.550 315.600 688.350 321.600 ;
        RECT 694.350 315.600 696.150 322.500 ;
        RECT 702.150 321.600 706.050 323.700 ;
        RECT 702.150 315.600 703.950 321.600 ;
        RECT 709.650 315.600 711.450 327.600 ;
        RECT 719.400 321.600 720.600 330.900 ;
        RECT 739.950 329.400 740.850 330.900 ;
        RECT 736.800 328.500 740.850 329.400 ;
        RECT 750.150 329.700 751.050 344.400 ;
        RECT 758.550 343.800 760.350 345.600 ;
        RECT 761.850 344.550 766.800 345.600 ;
        RECT 774.300 346.500 775.350 347.400 ;
        RECT 774.300 345.300 778.050 346.500 ;
        RECT 761.850 343.800 763.650 344.550 ;
        RECT 775.950 344.400 778.050 345.300 ;
        RECT 781.650 344.400 783.450 350.400 ;
        RECT 758.850 340.800 759.900 343.800 ;
        RECT 753.000 339.600 770.850 340.800 ;
        RECT 782.250 340.050 783.450 344.400 ;
        RECT 791.400 347.400 793.200 350.400 ;
        RECT 809.400 347.400 811.200 350.400 ;
        RECT 791.400 344.100 792.600 347.400 ;
        RECT 809.400 344.100 810.600 347.400 ;
        RECT 784.950 342.450 789.000 343.050 ;
        RECT 790.950 342.450 793.050 343.050 ;
        RECT 784.950 341.550 793.050 342.450 ;
        RECT 784.950 340.950 789.000 341.550 ;
        RECT 790.950 340.950 793.050 341.550 ;
        RECT 805.950 340.950 811.050 343.050 ;
        RECT 753.000 338.850 753.900 339.600 ;
        RECT 758.100 339.000 759.900 339.600 ;
        RECT 769.050 339.000 770.850 339.600 ;
        RECT 752.100 337.050 753.900 338.850 ;
        RECT 769.050 338.100 769.950 339.000 ;
        RECT 777.150 338.250 777.900 340.050 ;
        RECT 778.950 337.950 781.050 340.050 ;
        RECT 782.100 337.950 783.450 340.050 ;
        RECT 755.100 334.800 756.900 335.400 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 755.100 333.600 759.900 334.800 ;
        RECT 760.950 331.950 763.050 334.050 ;
        RECT 759.450 329.700 761.250 330.000 ;
        RECT 750.150 329.100 761.250 329.700 ;
        RECT 750.150 328.500 767.850 329.100 ;
        RECT 719.400 315.600 721.200 321.600 ;
        RECT 733.800 316.500 735.600 327.600 ;
        RECT 736.800 317.400 738.600 328.500 ;
        RECT 750.150 327.600 751.050 328.500 ;
        RECT 759.450 328.200 767.850 328.500 ;
        RECT 739.800 326.400 747.600 327.300 ;
        RECT 739.800 316.500 741.600 326.400 ;
        RECT 733.800 315.600 741.600 316.500 ;
        RECT 745.800 315.600 747.600 326.400 ;
        RECT 750.150 315.600 751.950 327.600 ;
        RECT 764.250 326.700 766.050 327.300 ;
        RECT 758.550 325.500 766.050 326.700 ;
        RECT 766.950 326.100 767.850 328.200 ;
        RECT 769.050 328.200 769.950 333.900 ;
        RECT 779.250 329.400 781.050 331.200 ;
        RECT 775.950 328.200 780.150 329.400 ;
        RECT 769.050 327.300 775.050 328.200 ;
        RECT 775.950 327.300 778.050 328.200 ;
        RECT 782.250 327.600 783.450 337.950 ;
        RECT 791.700 338.100 793.050 339.900 ;
        RECT 809.700 338.100 811.050 339.900 ;
        RECT 787.950 331.950 790.050 334.050 ;
        RECT 791.700 333.900 792.900 338.100 ;
        RECT 793.950 334.950 796.050 337.050 ;
        RECT 788.100 330.150 789.900 330.900 ;
        RECT 791.700 328.650 793.050 333.900 ;
        RECT 794.100 333.150 795.900 333.900 ;
        RECT 802.950 331.950 808.050 334.050 ;
        RECT 809.700 333.900 810.900 338.100 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 806.100 330.150 807.900 330.900 ;
        RECT 809.700 328.650 811.050 333.900 ;
        RECT 812.100 333.150 813.900 333.900 ;
        RECT 791.700 327.600 794.400 328.650 ;
        RECT 809.700 327.600 812.400 328.650 ;
        RECT 774.150 326.400 775.050 327.300 ;
        RECT 771.450 326.100 773.250 326.400 ;
        RECT 758.550 324.600 759.750 325.500 ;
        RECT 766.950 325.200 773.250 326.100 ;
        RECT 771.450 324.600 773.250 325.200 ;
        RECT 774.150 324.600 776.850 326.400 ;
        RECT 754.950 322.500 759.750 324.600 ;
        RECT 762.450 323.550 764.250 324.300 ;
        RECT 767.250 323.550 769.050 324.300 ;
        RECT 762.450 322.500 769.050 323.550 ;
        RECT 758.550 321.600 759.750 322.500 ;
        RECT 758.550 315.600 760.350 321.600 ;
        RECT 766.350 315.600 768.150 322.500 ;
        RECT 774.150 321.600 778.050 323.700 ;
        RECT 774.150 315.600 775.950 321.600 ;
        RECT 781.650 315.600 783.450 327.600 ;
        RECT 792.600 315.600 794.400 327.600 ;
        RECT 810.600 315.600 812.400 327.600 ;
        RECT 3.150 299.400 4.950 311.400 ;
        RECT 11.550 305.400 13.350 311.400 ;
        RECT 11.550 304.500 12.750 305.400 ;
        RECT 19.350 304.500 21.150 311.400 ;
        RECT 27.150 305.400 28.950 311.400 ;
        RECT 7.950 302.400 12.750 304.500 ;
        RECT 15.450 303.450 22.050 304.500 ;
        RECT 15.450 302.700 17.250 303.450 ;
        RECT 20.250 302.700 22.050 303.450 ;
        RECT 27.150 303.300 31.050 305.400 ;
        RECT 11.550 301.500 12.750 302.400 ;
        RECT 24.450 301.800 26.250 302.400 ;
        RECT 11.550 300.300 19.050 301.500 ;
        RECT 17.250 299.700 19.050 300.300 ;
        RECT 19.950 300.900 26.250 301.800 ;
        RECT 3.150 298.500 4.050 299.400 ;
        RECT 19.950 298.800 20.850 300.900 ;
        RECT 24.450 300.600 26.250 300.900 ;
        RECT 27.150 300.600 29.850 302.400 ;
        RECT 27.150 299.700 28.050 300.600 ;
        RECT 12.450 298.500 20.850 298.800 ;
        RECT 3.150 297.900 20.850 298.500 ;
        RECT 22.050 298.800 28.050 299.700 ;
        RECT 28.950 298.800 31.050 299.700 ;
        RECT 34.650 299.400 36.450 311.400 ;
        RECT 3.150 297.300 14.250 297.900 ;
        RECT 3.150 282.600 4.050 297.300 ;
        RECT 12.450 297.000 14.250 297.300 ;
        RECT 8.100 292.200 12.900 293.400 ;
        RECT 22.050 293.100 22.950 298.800 ;
        RECT 28.950 297.600 33.150 298.800 ;
        RECT 32.250 295.800 34.050 297.600 ;
        RECT 8.100 291.600 9.900 292.200 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 5.100 288.150 6.900 289.950 ;
        RECT 35.250 289.050 36.450 299.400 ;
        RECT 44.400 305.400 46.200 311.400 ;
        RECT 40.950 295.800 43.050 298.050 ;
        RECT 41.100 294.150 42.900 294.900 ;
        RECT 44.400 293.100 45.600 305.400 ;
        RECT 53.550 299.400 55.350 311.400 ;
        RECT 61.050 305.400 62.850 311.400 ;
        RECT 58.950 303.300 62.850 305.400 ;
        RECT 68.850 304.500 70.650 311.400 ;
        RECT 76.650 305.400 78.450 311.400 ;
        RECT 77.250 304.500 78.450 305.400 ;
        RECT 67.950 303.450 74.550 304.500 ;
        RECT 67.950 302.700 69.750 303.450 ;
        RECT 72.750 302.700 74.550 303.450 ;
        RECT 77.250 302.400 82.050 304.500 ;
        RECT 60.150 300.600 62.850 302.400 ;
        RECT 63.750 301.800 65.550 302.400 ;
        RECT 63.750 300.900 70.050 301.800 ;
        RECT 77.250 301.500 78.450 302.400 ;
        RECT 63.750 300.600 65.550 300.900 ;
        RECT 61.950 299.700 62.850 300.600 ;
        RECT 46.950 295.950 49.050 298.050 ;
        RECT 47.100 294.150 48.900 294.900 ;
        RECT 40.950 289.950 46.050 292.050 ;
        RECT 6.000 287.400 6.900 288.150 ;
        RECT 22.050 288.000 22.950 288.900 ;
        RECT 11.100 287.400 12.900 288.000 ;
        RECT 22.050 287.400 23.850 288.000 ;
        RECT 6.000 286.200 23.850 287.400 ;
        RECT 30.150 286.950 30.900 288.750 ;
        RECT 31.950 286.950 34.050 289.050 ;
        RECT 35.100 286.950 36.450 289.050 ;
        RECT 53.550 289.050 54.750 299.400 ;
        RECT 58.950 298.800 61.050 299.700 ;
        RECT 61.950 298.800 67.950 299.700 ;
        RECT 56.850 297.600 61.050 298.800 ;
        RECT 55.950 295.800 57.750 297.600 ;
        RECT 67.050 293.100 67.950 298.800 ;
        RECT 69.150 298.800 70.050 300.900 ;
        RECT 70.950 300.300 78.450 301.500 ;
        RECT 70.950 299.700 72.750 300.300 ;
        RECT 85.050 299.400 86.850 311.400 ;
        RECT 100.500 299.400 102.300 311.400 ;
        RECT 119.700 299.400 121.500 311.400 ;
        RECT 133.800 305.400 135.600 311.400 ;
        RECT 69.150 298.500 77.550 298.800 ;
        RECT 85.950 298.500 86.850 299.400 ;
        RECT 69.150 297.900 86.850 298.500 ;
        RECT 75.750 297.300 86.850 297.900 ;
        RECT 75.750 297.000 77.550 297.300 ;
        RECT 67.950 289.950 70.050 292.050 ;
        RECT 73.950 289.950 76.050 295.050 ;
        RECT 77.100 292.200 81.900 293.400 ;
        RECT 80.100 291.600 81.900 292.200 ;
        RECT 11.850 283.200 12.900 286.200 ;
        RECT 3.150 276.600 4.950 282.600 ;
        RECT 7.950 280.500 10.050 282.600 ;
        RECT 11.550 281.400 13.350 283.200 ;
        RECT 14.850 282.450 16.650 283.200 ;
        RECT 35.250 282.600 36.450 286.950 ;
        RECT 44.400 284.700 45.600 288.900 ;
        RECT 53.550 286.950 54.900 289.050 ;
        RECT 55.950 286.950 58.050 289.050 ;
        RECT 59.100 286.950 59.850 288.750 ;
        RECT 67.050 288.000 67.950 288.900 ;
        RECT 83.100 288.150 84.900 289.950 ;
        RECT 66.150 287.400 67.950 288.000 ;
        RECT 77.100 287.400 78.900 288.000 ;
        RECT 83.100 287.400 84.000 288.150 ;
        RECT 44.400 283.800 48.000 284.700 ;
        RECT 14.850 281.400 19.800 282.450 ;
        RECT 28.950 281.700 31.050 282.600 ;
        RECT 9.000 279.600 10.050 280.500 ;
        RECT 18.750 279.600 19.800 281.400 ;
        RECT 27.300 280.500 31.050 281.700 ;
        RECT 27.300 279.600 28.350 280.500 ;
        RECT 9.000 278.700 12.750 279.600 ;
        RECT 10.950 276.600 12.750 278.700 ;
        RECT 18.750 276.600 20.550 279.600 ;
        RECT 26.550 276.600 28.350 279.600 ;
        RECT 34.650 276.600 36.450 282.600 ;
        RECT 46.200 276.600 48.000 283.800 ;
        RECT 53.550 282.600 54.750 286.950 ;
        RECT 66.150 286.200 84.000 287.400 ;
        RECT 77.100 283.200 78.150 286.200 ;
        RECT 53.550 276.600 55.350 282.600 ;
        RECT 58.950 281.700 61.050 282.600 ;
        RECT 73.350 282.450 75.150 283.200 ;
        RECT 58.950 280.500 62.700 281.700 ;
        RECT 61.650 279.600 62.700 280.500 ;
        RECT 70.200 281.400 75.150 282.450 ;
        RECT 76.650 281.400 78.450 283.200 ;
        RECT 85.950 282.600 86.850 297.300 ;
        RECT 100.950 296.100 102.150 299.400 ;
        RECT 97.950 292.950 100.050 295.050 ;
        RECT 101.100 291.900 102.150 296.100 ;
        RECT 119.850 296.100 121.050 299.400 ;
        RECT 134.400 296.100 135.600 305.400 ;
        RECT 140.550 299.400 142.350 311.400 ;
        RECT 148.050 305.400 149.850 311.400 ;
        RECT 145.950 303.300 149.850 305.400 ;
        RECT 155.850 304.500 157.650 311.400 ;
        RECT 163.650 305.400 165.450 311.400 ;
        RECT 164.250 304.500 165.450 305.400 ;
        RECT 154.950 303.450 161.550 304.500 ;
        RECT 154.950 302.700 156.750 303.450 ;
        RECT 159.750 302.700 161.550 303.450 ;
        RECT 164.250 302.400 169.050 304.500 ;
        RECT 147.150 300.600 149.850 302.400 ;
        RECT 150.750 301.800 152.550 302.400 ;
        RECT 150.750 300.900 157.050 301.800 ;
        RECT 164.250 301.500 165.450 302.400 ;
        RECT 150.750 300.600 152.550 300.900 ;
        RECT 148.950 299.700 149.850 300.600 ;
        RECT 103.950 292.950 106.050 295.050 ;
        RECT 115.950 292.950 118.050 295.050 ;
        RECT 119.850 291.900 120.900 296.100 ;
        RECT 121.950 292.950 127.050 295.050 ;
        RECT 130.950 292.950 136.050 295.050 ;
        RECT 98.100 291.150 99.900 291.900 ;
        RECT 95.100 290.100 96.900 290.850 ;
        RECT 100.950 290.100 102.150 291.900 ;
        RECT 104.100 291.150 105.900 291.900 ;
        RECT 116.100 291.150 117.900 291.900 ;
        RECT 119.850 290.100 121.050 291.900 ;
        RECT 122.100 291.150 123.900 291.900 ;
        RECT 125.100 290.100 126.900 290.850 ;
        RECT 94.950 286.950 97.050 289.050 ;
        RECT 100.950 286.950 103.050 289.050 ;
        RECT 106.950 288.450 109.050 289.050 ;
        RECT 118.950 288.450 121.050 289.050 ;
        RECT 106.950 287.550 121.050 288.450 ;
        RECT 106.950 286.950 109.050 287.550 ;
        RECT 118.950 286.950 121.050 287.550 ;
        RECT 124.950 286.950 127.050 289.050 ;
        RECT 101.850 285.750 103.050 285.900 ;
        RECT 118.950 285.750 120.150 285.900 ;
        RECT 101.850 284.700 105.600 285.750 ;
        RECT 70.200 279.600 71.250 281.400 ;
        RECT 79.950 280.500 82.050 282.600 ;
        RECT 79.950 279.600 81.000 280.500 ;
        RECT 61.650 276.600 63.450 279.600 ;
        RECT 69.450 276.600 71.250 279.600 ;
        RECT 77.250 278.700 81.000 279.600 ;
        RECT 77.250 276.600 79.050 278.700 ;
        RECT 85.050 276.600 86.850 282.600 ;
        RECT 95.400 281.700 103.200 283.050 ;
        RECT 95.400 276.600 97.200 281.700 ;
        RECT 101.400 276.600 103.200 281.700 ;
        RECT 104.400 282.600 105.600 284.700 ;
        RECT 116.400 284.700 120.150 285.750 ;
        RECT 116.400 282.600 117.600 284.700 ;
        RECT 104.400 276.600 106.200 282.600 ;
        RECT 115.800 276.600 117.600 282.600 ;
        RECT 118.800 281.700 126.600 283.050 ;
        RECT 118.800 276.600 120.600 281.700 ;
        RECT 124.800 276.600 126.600 281.700 ;
        RECT 134.400 279.600 135.600 291.900 ;
        RECT 137.100 290.100 138.900 290.850 ;
        RECT 140.550 289.050 141.750 299.400 ;
        RECT 145.950 298.800 148.050 299.700 ;
        RECT 148.950 298.800 154.950 299.700 ;
        RECT 143.850 297.600 148.050 298.800 ;
        RECT 142.950 295.800 144.750 297.600 ;
        RECT 154.050 293.100 154.950 298.800 ;
        RECT 156.150 298.800 157.050 300.900 ;
        RECT 157.950 300.300 165.450 301.500 ;
        RECT 157.950 299.700 159.750 300.300 ;
        RECT 172.050 299.400 173.850 311.400 ;
        RECT 156.150 298.500 164.550 298.800 ;
        RECT 172.950 298.500 173.850 299.400 ;
        RECT 156.150 297.900 173.850 298.500 ;
        RECT 162.750 297.300 173.850 297.900 ;
        RECT 162.750 297.000 164.550 297.300 ;
        RECT 160.950 292.950 163.050 295.050 ;
        RECT 164.100 292.200 168.900 293.400 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 167.100 291.600 168.900 292.200 ;
        RECT 136.950 286.950 139.050 289.050 ;
        RECT 140.550 286.950 141.900 289.050 ;
        RECT 142.950 286.950 145.050 289.050 ;
        RECT 146.100 286.950 146.850 288.750 ;
        RECT 154.050 288.000 154.950 288.900 ;
        RECT 170.100 288.150 171.900 289.950 ;
        RECT 153.150 287.400 154.950 288.000 ;
        RECT 164.100 287.400 165.900 288.000 ;
        RECT 170.100 287.400 171.000 288.150 ;
        RECT 133.800 276.600 135.600 279.600 ;
        RECT 140.550 282.600 141.750 286.950 ;
        RECT 153.150 286.200 171.000 287.400 ;
        RECT 164.100 283.200 165.150 286.200 ;
        RECT 140.550 276.600 142.350 282.600 ;
        RECT 145.950 281.700 148.050 282.600 ;
        RECT 160.350 282.450 162.150 283.200 ;
        RECT 145.950 280.500 149.700 281.700 ;
        RECT 148.650 279.600 149.700 280.500 ;
        RECT 157.200 281.400 162.150 282.450 ;
        RECT 163.650 281.400 165.450 283.200 ;
        RECT 172.950 282.600 173.850 297.300 ;
        RECT 157.200 279.600 158.250 281.400 ;
        RECT 166.950 280.500 169.050 282.600 ;
        RECT 166.950 279.600 168.000 280.500 ;
        RECT 148.650 276.600 150.450 279.600 ;
        RECT 156.450 276.600 158.250 279.600 ;
        RECT 164.250 278.700 168.000 279.600 ;
        RECT 164.250 276.600 166.050 278.700 ;
        RECT 172.050 276.600 173.850 282.600 ;
        RECT 177.150 299.400 178.950 311.400 ;
        RECT 185.550 305.400 187.350 311.400 ;
        RECT 185.550 304.500 186.750 305.400 ;
        RECT 193.350 304.500 195.150 311.400 ;
        RECT 201.150 305.400 202.950 311.400 ;
        RECT 181.950 302.400 186.750 304.500 ;
        RECT 189.450 303.450 196.050 304.500 ;
        RECT 189.450 302.700 191.250 303.450 ;
        RECT 194.250 302.700 196.050 303.450 ;
        RECT 201.150 303.300 205.050 305.400 ;
        RECT 185.550 301.500 186.750 302.400 ;
        RECT 198.450 301.800 200.250 302.400 ;
        RECT 185.550 300.300 193.050 301.500 ;
        RECT 191.250 299.700 193.050 300.300 ;
        RECT 193.950 300.900 200.250 301.800 ;
        RECT 177.150 298.500 178.050 299.400 ;
        RECT 193.950 298.800 194.850 300.900 ;
        RECT 198.450 300.600 200.250 300.900 ;
        RECT 201.150 300.600 203.850 302.400 ;
        RECT 201.150 299.700 202.050 300.600 ;
        RECT 186.450 298.500 194.850 298.800 ;
        RECT 177.150 297.900 194.850 298.500 ;
        RECT 196.050 298.800 202.050 299.700 ;
        RECT 202.950 298.800 205.050 299.700 ;
        RECT 208.650 299.400 210.450 311.400 ;
        RECT 177.150 297.300 188.250 297.900 ;
        RECT 177.150 282.600 178.050 297.300 ;
        RECT 186.450 297.000 188.250 297.300 ;
        RECT 182.100 292.200 186.900 293.400 ;
        RECT 187.950 292.950 193.050 295.050 ;
        RECT 196.050 293.100 196.950 298.800 ;
        RECT 202.950 297.600 207.150 298.800 ;
        RECT 206.250 295.800 208.050 297.600 ;
        RECT 182.100 291.600 183.900 292.200 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 179.100 288.150 180.900 289.950 ;
        RECT 209.250 289.050 210.450 299.400 ;
        RECT 180.000 287.400 180.900 288.150 ;
        RECT 196.050 288.000 196.950 288.900 ;
        RECT 185.100 287.400 186.900 288.000 ;
        RECT 196.050 287.400 197.850 288.000 ;
        RECT 180.000 286.200 197.850 287.400 ;
        RECT 204.150 286.950 204.900 288.750 ;
        RECT 205.950 286.950 208.050 289.050 ;
        RECT 209.100 286.950 210.450 289.050 ;
        RECT 185.850 283.200 186.900 286.200 ;
        RECT 177.150 276.600 178.950 282.600 ;
        RECT 181.950 280.500 184.050 282.600 ;
        RECT 185.550 281.400 187.350 283.200 ;
        RECT 188.850 282.450 190.650 283.200 ;
        RECT 209.250 282.600 210.450 286.950 ;
        RECT 188.850 281.400 193.800 282.450 ;
        RECT 202.950 281.700 205.050 282.600 ;
        RECT 183.000 279.600 184.050 280.500 ;
        RECT 192.750 279.600 193.800 281.400 ;
        RECT 201.300 280.500 205.050 281.700 ;
        RECT 201.300 279.600 202.350 280.500 ;
        RECT 183.000 278.700 186.750 279.600 ;
        RECT 184.950 276.600 186.750 278.700 ;
        RECT 192.750 276.600 194.550 279.600 ;
        RECT 200.550 276.600 202.350 279.600 ;
        RECT 208.650 276.600 210.450 282.600 ;
        RECT 213.150 299.400 214.950 311.400 ;
        RECT 221.550 305.400 223.350 311.400 ;
        RECT 221.550 304.500 222.750 305.400 ;
        RECT 229.350 304.500 231.150 311.400 ;
        RECT 237.150 305.400 238.950 311.400 ;
        RECT 217.950 302.400 222.750 304.500 ;
        RECT 225.450 303.450 232.050 304.500 ;
        RECT 225.450 302.700 227.250 303.450 ;
        RECT 230.250 302.700 232.050 303.450 ;
        RECT 237.150 303.300 241.050 305.400 ;
        RECT 221.550 301.500 222.750 302.400 ;
        RECT 234.450 301.800 236.250 302.400 ;
        RECT 221.550 300.300 229.050 301.500 ;
        RECT 227.250 299.700 229.050 300.300 ;
        RECT 229.950 300.900 236.250 301.800 ;
        RECT 213.150 298.500 214.050 299.400 ;
        RECT 229.950 298.800 230.850 300.900 ;
        RECT 234.450 300.600 236.250 300.900 ;
        RECT 237.150 300.600 239.850 302.400 ;
        RECT 237.150 299.700 238.050 300.600 ;
        RECT 222.450 298.500 230.850 298.800 ;
        RECT 213.150 297.900 230.850 298.500 ;
        RECT 232.050 298.800 238.050 299.700 ;
        RECT 238.950 298.800 241.050 299.700 ;
        RECT 244.650 299.400 246.450 311.400 ;
        RECT 213.150 297.300 224.250 297.900 ;
        RECT 213.150 282.600 214.050 297.300 ;
        RECT 222.450 297.000 224.250 297.300 ;
        RECT 218.100 292.200 222.900 293.400 ;
        RECT 223.950 292.800 226.050 295.050 ;
        RECT 232.050 293.100 232.950 298.800 ;
        RECT 238.950 297.600 243.150 298.800 ;
        RECT 242.250 295.800 244.050 297.600 ;
        RECT 218.100 291.600 219.900 292.200 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 215.100 288.150 216.900 289.950 ;
        RECT 245.250 289.050 246.450 299.400 ;
        RECT 254.400 305.400 256.200 311.400 ;
        RECT 254.400 296.100 255.600 305.400 ;
        RECT 270.600 299.400 272.400 311.400 ;
        RECT 285.600 299.400 287.400 311.400 ;
        RECT 303.600 299.400 305.400 311.400 ;
        RECT 319.800 305.400 321.600 311.400 ;
        RECT 270.600 298.350 273.300 299.400 ;
        RECT 285.600 298.350 288.300 299.400 ;
        RECT 303.600 298.350 306.300 299.400 ;
        RECT 253.950 292.950 256.050 295.050 ;
        RECT 269.100 293.100 270.900 293.850 ;
        RECT 271.950 293.100 273.300 298.350 ;
        RECT 275.100 296.100 276.900 296.850 ;
        RECT 251.100 290.100 252.900 290.850 ;
        RECT 216.000 287.400 216.900 288.150 ;
        RECT 232.050 288.000 232.950 288.900 ;
        RECT 221.100 287.400 222.900 288.000 ;
        RECT 232.050 287.400 233.850 288.000 ;
        RECT 216.000 286.200 233.850 287.400 ;
        RECT 240.150 286.950 240.900 288.750 ;
        RECT 241.950 286.950 244.050 289.050 ;
        RECT 245.100 286.950 246.450 289.050 ;
        RECT 250.950 286.950 253.050 289.050 ;
        RECT 221.850 283.200 222.900 286.200 ;
        RECT 213.150 276.600 214.950 282.600 ;
        RECT 217.950 280.500 220.050 282.600 ;
        RECT 221.550 281.400 223.350 283.200 ;
        RECT 224.850 282.450 226.650 283.200 ;
        RECT 245.250 282.600 246.450 286.950 ;
        RECT 224.850 281.400 229.800 282.450 ;
        RECT 238.950 281.700 241.050 282.600 ;
        RECT 219.000 279.600 220.050 280.500 ;
        RECT 228.750 279.600 229.800 281.400 ;
        RECT 237.300 280.500 241.050 281.700 ;
        RECT 237.300 279.600 238.350 280.500 ;
        RECT 219.000 278.700 222.750 279.600 ;
        RECT 220.950 276.600 222.750 278.700 ;
        RECT 228.750 276.600 230.550 279.600 ;
        RECT 236.550 276.600 238.350 279.600 ;
        RECT 244.650 276.600 246.450 282.600 ;
        RECT 254.400 279.600 255.600 291.900 ;
        RECT 259.950 291.450 262.050 292.050 ;
        RECT 268.950 291.450 271.050 292.050 ;
        RECT 259.950 290.550 271.050 291.450 ;
        RECT 259.950 289.950 262.050 290.550 ;
        RECT 268.950 289.950 271.050 290.550 ;
        RECT 272.100 288.900 273.300 293.100 ;
        RECT 274.950 292.950 280.050 295.050 ;
        RECT 284.100 293.100 285.900 293.850 ;
        RECT 286.950 293.100 288.300 298.350 ;
        RECT 290.100 296.100 291.900 296.850 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 287.100 288.900 288.300 293.100 ;
        RECT 289.950 292.950 292.050 295.050 ;
        RECT 302.100 293.100 303.900 293.850 ;
        RECT 304.950 293.100 306.300 298.350 ;
        RECT 308.100 296.100 309.900 296.850 ;
        RECT 320.400 296.100 321.600 305.400 ;
        RECT 326.550 299.400 328.350 311.400 ;
        RECT 334.050 305.400 335.850 311.400 ;
        RECT 331.950 303.300 335.850 305.400 ;
        RECT 341.850 304.500 343.650 311.400 ;
        RECT 349.650 305.400 351.450 311.400 ;
        RECT 350.250 304.500 351.450 305.400 ;
        RECT 340.950 303.450 347.550 304.500 ;
        RECT 340.950 302.700 342.750 303.450 ;
        RECT 345.750 302.700 347.550 303.450 ;
        RECT 350.250 302.400 355.050 304.500 ;
        RECT 333.150 300.600 335.850 302.400 ;
        RECT 336.750 301.800 338.550 302.400 ;
        RECT 336.750 300.900 343.050 301.800 ;
        RECT 350.250 301.500 351.450 302.400 ;
        RECT 336.750 300.600 338.550 300.900 ;
        RECT 334.950 299.700 335.850 300.600 ;
        RECT 295.950 291.450 300.000 292.050 ;
        RECT 301.950 291.450 304.050 292.050 ;
        RECT 295.950 290.550 304.050 291.450 ;
        RECT 295.950 289.950 300.000 290.550 ;
        RECT 301.950 289.950 304.050 290.550 ;
        RECT 305.100 288.900 306.300 293.100 ;
        RECT 307.950 294.450 310.050 295.050 ;
        RECT 312.000 294.450 316.050 295.050 ;
        RECT 307.950 293.550 316.050 294.450 ;
        RECT 307.950 292.950 310.050 293.550 ;
        RECT 312.000 292.950 316.050 293.550 ;
        RECT 319.950 292.950 322.050 295.050 ;
        RECT 271.950 287.100 273.300 288.900 ;
        RECT 286.950 287.100 288.300 288.900 ;
        RECT 304.950 287.100 306.300 288.900 ;
        RECT 256.950 285.450 259.050 286.050 ;
        RECT 271.950 285.450 274.050 286.050 ;
        RECT 256.950 284.550 274.050 285.450 ;
        RECT 256.950 283.950 259.050 284.550 ;
        RECT 271.950 283.950 274.050 284.550 ;
        RECT 286.950 285.450 289.050 286.050 ;
        RECT 291.000 285.450 295.050 286.050 ;
        RECT 286.950 284.550 295.050 285.450 ;
        RECT 286.950 283.950 289.050 284.550 ;
        RECT 291.000 283.950 295.050 284.550 ;
        RECT 304.950 283.950 310.050 286.050 ;
        RECT 272.400 279.600 273.600 282.900 ;
        RECT 287.400 279.600 288.600 282.900 ;
        RECT 305.400 279.600 306.600 282.900 ;
        RECT 320.400 279.600 321.600 291.900 ;
        RECT 323.100 290.100 324.900 290.850 ;
        RECT 326.550 289.050 327.750 299.400 ;
        RECT 331.950 298.800 334.050 299.700 ;
        RECT 334.950 298.800 340.950 299.700 ;
        RECT 329.850 297.600 334.050 298.800 ;
        RECT 328.950 295.800 330.750 297.600 ;
        RECT 340.050 293.100 340.950 298.800 ;
        RECT 342.150 298.800 343.050 300.900 ;
        RECT 343.950 300.300 351.450 301.500 ;
        RECT 343.950 299.700 345.750 300.300 ;
        RECT 358.050 299.400 359.850 311.400 ;
        RECT 373.500 299.400 375.300 311.400 ;
        RECT 394.500 299.400 396.300 311.400 ;
        RECT 416.700 299.400 418.500 311.400 ;
        RECT 431.400 305.400 433.200 311.400 ;
        RECT 342.150 298.500 350.550 298.800 ;
        RECT 358.950 298.500 359.850 299.400 ;
        RECT 342.150 297.900 359.850 298.500 ;
        RECT 348.750 297.300 359.850 297.900 ;
        RECT 348.750 297.000 350.550 297.300 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 346.950 289.950 349.050 295.050 ;
        RECT 350.100 292.200 354.900 293.400 ;
        RECT 353.100 291.600 354.900 292.200 ;
        RECT 322.950 286.950 325.050 289.050 ;
        RECT 326.550 286.950 327.900 289.050 ;
        RECT 328.950 286.950 331.050 289.050 ;
        RECT 332.100 286.950 332.850 288.750 ;
        RECT 340.050 288.000 340.950 288.900 ;
        RECT 356.100 288.150 357.900 289.950 ;
        RECT 339.150 287.400 340.950 288.000 ;
        RECT 350.100 287.400 351.900 288.000 ;
        RECT 356.100 287.400 357.000 288.150 ;
        RECT 254.400 276.600 256.200 279.600 ;
        RECT 271.800 276.600 273.600 279.600 ;
        RECT 286.800 276.600 288.600 279.600 ;
        RECT 304.800 276.600 306.600 279.600 ;
        RECT 319.800 276.600 321.600 279.600 ;
        RECT 326.550 282.600 327.750 286.950 ;
        RECT 339.150 286.200 357.000 287.400 ;
        RECT 350.100 283.200 351.150 286.200 ;
        RECT 326.550 276.600 328.350 282.600 ;
        RECT 331.950 281.700 334.050 282.600 ;
        RECT 346.350 282.450 348.150 283.200 ;
        RECT 331.950 280.500 335.700 281.700 ;
        RECT 334.650 279.600 335.700 280.500 ;
        RECT 343.200 281.400 348.150 282.450 ;
        RECT 349.650 281.400 351.450 283.200 ;
        RECT 358.950 282.600 359.850 297.300 ;
        RECT 373.950 296.100 375.150 299.400 ;
        RECT 394.950 296.100 396.150 299.400 ;
        RECT 370.950 292.950 373.050 295.050 ;
        RECT 374.100 291.900 375.150 296.100 ;
        RECT 376.950 292.950 379.050 295.050 ;
        RECT 391.950 292.950 394.050 295.050 ;
        RECT 395.100 291.900 396.150 296.100 ;
        RECT 397.950 292.950 400.050 298.050 ;
        RECT 416.850 296.100 418.050 299.400 ;
        RECT 412.950 292.950 415.050 295.050 ;
        RECT 416.850 291.900 417.900 296.100 ;
        RECT 427.950 295.950 430.050 298.050 ;
        RECT 418.950 292.950 421.050 295.050 ;
        RECT 428.100 294.150 429.900 294.900 ;
        RECT 431.400 293.100 432.600 305.400 ;
        RECT 448.500 299.400 450.300 311.400 ;
        RECT 458.550 299.400 460.350 311.400 ;
        RECT 466.050 305.400 467.850 311.400 ;
        RECT 463.950 303.300 467.850 305.400 ;
        RECT 473.850 304.500 475.650 311.400 ;
        RECT 481.650 305.400 483.450 311.400 ;
        RECT 482.250 304.500 483.450 305.400 ;
        RECT 472.950 303.450 479.550 304.500 ;
        RECT 472.950 302.700 474.750 303.450 ;
        RECT 477.750 302.700 479.550 303.450 ;
        RECT 482.250 302.400 487.050 304.500 ;
        RECT 465.150 300.600 467.850 302.400 ;
        RECT 468.750 301.800 470.550 302.400 ;
        RECT 468.750 300.900 475.050 301.800 ;
        RECT 482.250 301.500 483.450 302.400 ;
        RECT 468.750 300.600 470.550 300.900 ;
        RECT 466.950 299.700 467.850 300.600 ;
        RECT 433.950 295.950 436.050 298.050 ;
        RECT 448.950 296.100 450.150 299.400 ;
        RECT 434.100 294.150 435.900 294.900 ;
        RECT 445.950 292.950 448.050 295.050 ;
        RECT 371.100 291.150 372.900 291.900 ;
        RECT 368.100 290.100 369.900 290.850 ;
        RECT 373.950 290.100 375.150 291.900 ;
        RECT 377.100 291.150 378.900 291.900 ;
        RECT 392.100 291.150 393.900 291.900 ;
        RECT 389.100 290.100 390.900 290.850 ;
        RECT 394.950 290.100 396.150 291.900 ;
        RECT 398.100 291.150 399.900 291.900 ;
        RECT 413.100 291.150 414.900 291.900 ;
        RECT 416.850 290.100 418.050 291.900 ;
        RECT 419.100 291.150 420.900 291.900 ;
        RECT 422.100 290.100 423.900 290.850 ;
        RECT 427.950 289.950 433.050 292.050 ;
        RECT 449.100 291.900 450.150 296.100 ;
        RECT 451.950 292.950 454.050 295.200 ;
        RECT 446.100 291.150 447.900 291.900 ;
        RECT 443.100 290.100 444.900 290.850 ;
        RECT 448.950 290.100 450.150 291.900 ;
        RECT 452.100 291.150 453.900 291.900 ;
        RECT 451.950 289.050 454.050 289.200 ;
        RECT 367.950 286.950 370.050 289.050 ;
        RECT 373.950 286.950 376.050 289.050 ;
        RECT 388.950 286.950 391.050 289.050 ;
        RECT 394.950 288.450 397.050 289.050 ;
        RECT 399.000 288.450 402.900 289.050 ;
        RECT 394.950 287.550 402.900 288.450 ;
        RECT 394.950 286.950 397.050 287.550 ;
        RECT 399.000 286.950 402.900 287.550 ;
        RECT 403.950 288.450 406.050 289.050 ;
        RECT 415.950 288.450 418.050 289.050 ;
        RECT 403.950 287.550 418.050 288.450 ;
        RECT 403.950 286.950 406.050 287.550 ;
        RECT 415.950 286.950 418.050 287.550 ;
        RECT 421.950 286.950 424.050 289.050 ;
        RECT 374.850 285.750 376.050 285.900 ;
        RECT 395.850 285.750 397.050 285.900 ;
        RECT 415.950 285.750 417.150 285.900 ;
        RECT 374.850 284.700 378.600 285.750 ;
        RECT 395.850 284.700 399.600 285.750 ;
        RECT 343.200 279.600 344.250 281.400 ;
        RECT 352.950 280.500 355.050 282.600 ;
        RECT 352.950 279.600 354.000 280.500 ;
        RECT 334.650 276.600 336.450 279.600 ;
        RECT 342.450 276.600 344.250 279.600 ;
        RECT 350.250 278.700 354.000 279.600 ;
        RECT 350.250 276.600 352.050 278.700 ;
        RECT 358.050 276.600 359.850 282.600 ;
        RECT 368.400 281.700 376.200 283.050 ;
        RECT 368.400 276.600 370.200 281.700 ;
        RECT 374.400 276.600 376.200 281.700 ;
        RECT 377.400 282.600 378.600 284.700 ;
        RECT 377.400 276.600 379.200 282.600 ;
        RECT 389.400 281.700 397.200 283.050 ;
        RECT 389.400 276.600 391.200 281.700 ;
        RECT 395.400 276.600 397.200 281.700 ;
        RECT 398.400 282.600 399.600 284.700 ;
        RECT 413.400 284.700 417.150 285.750 ;
        RECT 431.400 284.700 432.600 288.900 ;
        RECT 442.950 286.950 445.050 289.050 ;
        RECT 448.950 287.100 454.050 289.050 ;
        RECT 458.550 289.050 459.750 299.400 ;
        RECT 463.950 298.800 466.050 299.700 ;
        RECT 466.950 298.800 472.950 299.700 ;
        RECT 461.850 297.600 466.050 298.800 ;
        RECT 460.950 295.800 462.750 297.600 ;
        RECT 472.050 293.100 472.950 298.800 ;
        RECT 474.150 298.800 475.050 300.900 ;
        RECT 475.950 300.300 483.450 301.500 ;
        RECT 475.950 299.700 477.750 300.300 ;
        RECT 490.050 299.400 491.850 311.400 ;
        RECT 474.150 298.500 482.550 298.800 ;
        RECT 490.950 298.500 491.850 299.400 ;
        RECT 474.150 297.900 491.850 298.500 ;
        RECT 500.400 305.400 502.200 311.400 ;
        RECT 480.750 297.300 491.850 297.900 ;
        RECT 480.750 297.000 482.550 297.300 ;
        RECT 478.950 292.950 481.050 295.050 ;
        RECT 482.100 292.200 486.900 293.400 ;
        RECT 472.950 289.950 475.050 292.050 ;
        RECT 485.100 291.600 486.900 292.200 ;
        RECT 448.950 286.950 453.450 287.100 ;
        RECT 458.550 286.950 459.900 289.050 ;
        RECT 460.950 286.950 463.050 289.050 ;
        RECT 464.100 286.950 464.850 288.750 ;
        RECT 472.050 288.000 472.950 288.900 ;
        RECT 488.100 288.150 489.900 289.950 ;
        RECT 471.150 287.400 472.950 288.000 ;
        RECT 482.100 287.400 483.900 288.000 ;
        RECT 488.100 287.400 489.000 288.150 ;
        RECT 449.850 285.750 451.050 285.900 ;
        RECT 449.850 284.700 453.600 285.750 ;
        RECT 413.400 282.600 414.600 284.700 ;
        RECT 431.400 283.800 435.000 284.700 ;
        RECT 398.400 276.600 400.200 282.600 ;
        RECT 412.800 276.600 414.600 282.600 ;
        RECT 415.800 281.700 423.600 283.050 ;
        RECT 415.800 276.600 417.600 281.700 ;
        RECT 421.800 276.600 423.600 281.700 ;
        RECT 433.200 276.600 435.000 283.800 ;
        RECT 443.400 281.700 451.200 283.050 ;
        RECT 443.400 276.600 445.200 281.700 ;
        RECT 449.400 276.600 451.200 281.700 ;
        RECT 452.400 282.600 453.600 284.700 ;
        RECT 458.550 282.600 459.750 286.950 ;
        RECT 471.150 286.200 489.000 287.400 ;
        RECT 482.100 283.200 483.150 286.200 ;
        RECT 452.400 276.600 454.200 282.600 ;
        RECT 458.550 276.600 460.350 282.600 ;
        RECT 463.950 281.700 466.050 282.600 ;
        RECT 478.350 282.450 480.150 283.200 ;
        RECT 463.950 280.500 467.700 281.700 ;
        RECT 466.650 279.600 467.700 280.500 ;
        RECT 475.200 281.400 480.150 282.450 ;
        RECT 481.650 281.400 483.450 283.200 ;
        RECT 490.950 282.600 491.850 297.300 ;
        RECT 496.950 295.950 499.050 298.050 ;
        RECT 497.100 294.150 498.900 294.900 ;
        RECT 500.400 293.100 501.600 305.400 ;
        RECT 519.600 299.400 521.400 311.400 ;
        RECT 530.400 300.300 532.200 311.400 ;
        RECT 536.400 300.300 538.200 311.400 ;
        RECT 530.400 299.400 538.200 300.300 ;
        RECT 539.400 299.400 541.200 311.400 ;
        RECT 548.400 305.400 550.200 311.400 ;
        RECT 519.600 298.350 522.300 299.400 ;
        RECT 502.950 295.950 505.050 298.050 ;
        RECT 503.100 294.150 504.900 294.900 ;
        RECT 518.100 293.100 519.900 293.850 ;
        RECT 520.950 293.100 522.300 298.350 ;
        RECT 524.100 296.100 525.900 296.850 ;
        RECT 493.950 291.450 498.000 292.050 ;
        RECT 499.950 291.450 502.050 292.050 ;
        RECT 493.950 290.550 502.050 291.450 ;
        RECT 493.950 289.950 498.000 290.550 ;
        RECT 499.950 289.950 502.050 290.550 ;
        RECT 517.950 289.950 520.050 292.050 ;
        RECT 521.100 288.900 522.300 293.100 ;
        RECT 523.950 292.950 526.050 295.050 ;
        RECT 529.950 292.950 532.050 295.050 ;
        RECT 535.950 292.950 538.050 295.050 ;
        RECT 530.100 291.150 531.900 291.900 ;
        RECT 536.100 291.150 537.900 291.900 ;
        RECT 533.100 290.100 534.900 290.850 ;
        RECT 539.700 290.100 540.600 299.400 ;
        RECT 548.400 298.500 549.600 305.400 ;
        RECT 554.700 299.400 556.500 311.400 ;
        RECT 569.700 299.400 571.500 311.400 ;
        RECT 587.400 305.400 589.200 311.400 ;
        RECT 548.400 297.600 554.100 298.500 ;
        RECT 552.150 296.700 554.100 297.600 ;
        RECT 548.100 293.100 549.900 293.850 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 552.150 290.100 553.050 296.700 ;
        RECT 555.000 290.100 556.200 299.400 ;
        RECT 569.850 296.100 571.050 299.400 ;
        RECT 565.950 292.950 568.050 295.050 ;
        RECT 569.850 291.900 570.900 296.100 ;
        RECT 583.950 295.950 586.050 301.050 ;
        RECT 571.950 292.950 574.050 295.050 ;
        RECT 584.100 294.150 585.900 294.900 ;
        RECT 587.400 293.100 588.600 305.400 ;
        RECT 603.600 299.400 605.400 311.400 ;
        RECT 621.600 299.400 623.400 311.400 ;
        RECT 632.400 300.300 634.200 311.400 ;
        RECT 638.400 300.300 640.200 311.400 ;
        RECT 632.400 299.400 640.200 300.300 ;
        RECT 641.400 299.400 643.200 311.400 ;
        RECT 659.700 299.400 661.500 311.400 ;
        RECT 673.200 299.400 675.000 311.400 ;
        RECT 679.800 305.400 681.600 311.400 ;
        RECT 602.700 298.350 605.400 299.400 ;
        RECT 620.700 298.350 623.400 299.400 ;
        RECT 589.950 295.950 592.050 298.050 ;
        RECT 599.100 296.100 600.900 296.850 ;
        RECT 590.100 294.150 591.900 294.900 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 602.700 293.100 604.050 298.350 ;
        RECT 617.100 296.100 618.900 296.850 ;
        RECT 605.100 293.100 606.900 293.850 ;
        RECT 566.100 291.150 567.900 291.900 ;
        RECT 569.850 290.100 571.050 291.900 ;
        RECT 572.100 291.150 573.900 291.900 ;
        RECT 580.950 291.450 585.000 292.050 ;
        RECT 586.950 291.450 589.050 292.050 ;
        RECT 575.100 290.100 576.900 290.850 ;
        RECT 580.950 290.550 589.050 291.450 ;
        RECT 500.400 284.700 501.600 288.900 ;
        RECT 520.950 287.100 522.300 288.900 ;
        RECT 532.950 286.950 535.050 289.050 ;
        RECT 538.950 286.950 541.050 289.050 ;
        RECT 520.950 285.450 523.050 286.050 ;
        RECT 525.000 285.450 529.050 286.050 ;
        RECT 552.150 285.900 552.900 290.100 ;
        RECT 580.950 289.950 585.000 290.550 ;
        RECT 586.950 289.950 589.050 290.550 ;
        RECT 553.950 286.950 556.050 289.050 ;
        RECT 562.950 288.450 567.000 289.050 ;
        RECT 568.950 288.450 571.050 289.050 ;
        RECT 562.950 287.550 571.050 288.450 ;
        RECT 562.950 286.950 567.000 287.550 ;
        RECT 568.950 286.950 571.050 287.550 ;
        RECT 574.950 286.950 577.050 289.050 ;
        RECT 602.700 288.900 603.900 293.100 ;
        RECT 616.950 292.950 619.050 295.050 ;
        RECT 620.700 293.100 622.050 298.350 ;
        RECT 623.100 293.100 624.900 293.850 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 620.700 288.900 621.900 293.100 ;
        RECT 631.950 292.950 634.050 295.050 ;
        RECT 637.950 292.950 640.050 295.050 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 632.100 291.150 633.900 291.900 ;
        RECT 638.100 291.150 639.900 291.900 ;
        RECT 635.100 290.100 636.900 290.850 ;
        RECT 641.700 290.100 642.600 299.400 ;
        RECT 659.850 296.100 661.050 299.400 ;
        RECT 655.950 292.950 658.050 295.050 ;
        RECT 659.850 291.900 660.900 296.100 ;
        RECT 661.950 292.950 664.050 295.050 ;
        RECT 656.100 291.150 657.900 291.900 ;
        RECT 659.850 290.100 661.050 291.900 ;
        RECT 662.100 291.150 663.900 291.900 ;
        RECT 665.100 290.100 666.900 290.850 ;
        RECT 673.950 290.100 675.000 299.400 ;
        RECT 676.950 292.950 679.050 295.050 ;
        RECT 677.100 291.150 678.900 291.900 ;
        RECT 500.400 283.800 504.000 284.700 ;
        RECT 520.950 284.550 529.050 285.450 ;
        RECT 520.950 283.950 523.050 284.550 ;
        RECT 525.000 283.950 529.050 284.550 ;
        RECT 475.200 279.600 476.250 281.400 ;
        RECT 484.950 280.500 487.050 282.600 ;
        RECT 484.950 279.600 486.000 280.500 ;
        RECT 466.650 276.600 468.450 279.600 ;
        RECT 474.450 276.600 476.250 279.600 ;
        RECT 482.250 278.700 486.000 279.600 ;
        RECT 482.250 276.600 484.050 278.700 ;
        RECT 490.050 276.600 491.850 282.600 ;
        RECT 502.200 276.600 504.000 283.800 ;
        RECT 521.400 279.600 522.600 282.900 ;
        RECT 539.700 282.600 540.600 285.900 ;
        RECT 552.150 285.300 553.050 285.900 ;
        RECT 552.150 284.400 554.100 285.300 ;
        RECT 520.800 276.600 522.600 279.600 ;
        RECT 535.200 280.950 540.600 282.600 ;
        RECT 549.000 283.500 554.100 284.400 ;
        RECT 535.200 276.600 537.000 280.950 ;
        RECT 549.000 279.600 550.200 283.500 ;
        RECT 555.000 282.600 556.200 285.900 ;
        RECT 568.950 285.750 570.150 285.900 ;
        RECT 566.400 284.700 570.150 285.750 ;
        RECT 587.400 284.700 588.600 288.900 ;
        RECT 602.700 287.100 604.050 288.900 ;
        RECT 620.700 287.100 622.050 288.900 ;
        RECT 634.950 286.950 637.050 289.050 ;
        RECT 640.950 288.450 643.050 289.050 ;
        RECT 652.800 288.450 654.900 289.050 ;
        RECT 640.950 287.550 654.900 288.450 ;
        RECT 640.950 286.950 643.050 287.550 ;
        RECT 652.800 286.950 654.900 287.550 ;
        RECT 655.950 286.950 661.050 289.050 ;
        RECT 664.950 286.950 667.050 289.050 ;
        RECT 670.950 286.950 676.050 289.050 ;
        RECT 601.950 285.450 604.050 286.050 ;
        RECT 613.950 285.450 616.050 286.050 ;
        RECT 566.400 282.600 567.600 284.700 ;
        RECT 587.400 283.800 591.000 284.700 ;
        RECT 601.950 284.550 616.050 285.450 ;
        RECT 601.950 283.950 604.050 284.550 ;
        RECT 613.950 283.950 616.050 284.550 ;
        RECT 619.950 285.450 622.050 286.050 ;
        RECT 624.000 285.450 628.050 286.050 ;
        RECT 619.950 284.550 628.050 285.450 ;
        RECT 619.950 283.950 622.050 284.550 ;
        RECT 624.000 283.950 628.050 284.550 ;
        RECT 548.400 276.600 550.200 279.600 ;
        RECT 554.700 276.600 556.500 282.600 ;
        RECT 565.800 276.600 567.600 282.600 ;
        RECT 568.800 281.700 576.600 283.050 ;
        RECT 568.800 276.600 570.600 281.700 ;
        RECT 574.800 276.600 576.600 281.700 ;
        RECT 589.200 276.600 591.000 283.800 ;
        RECT 602.400 279.600 603.600 282.900 ;
        RECT 620.400 279.600 621.600 282.900 ;
        RECT 641.700 282.600 642.600 285.900 ;
        RECT 658.950 285.750 660.150 285.900 ;
        RECT 656.400 284.700 660.150 285.750 ;
        RECT 656.400 282.600 657.600 284.700 ;
        RECT 637.200 280.950 642.600 282.600 ;
        RECT 602.400 276.600 604.200 279.600 ;
        RECT 620.400 276.600 622.200 279.600 ;
        RECT 637.200 276.600 639.000 280.950 ;
        RECT 655.800 276.600 657.600 282.600 ;
        RECT 658.800 281.700 666.600 283.050 ;
        RECT 658.800 276.600 660.600 281.700 ;
        RECT 664.800 276.600 666.600 281.700 ;
        RECT 675.150 282.600 676.050 285.900 ;
        RECT 680.550 285.300 681.600 305.400 ;
        RECT 696.600 299.400 698.400 311.400 ;
        RECT 711.600 299.400 713.400 311.400 ;
        RECT 727.500 299.400 729.300 311.400 ;
        RECT 749.700 299.400 751.500 311.400 ;
        RECT 768.600 299.400 770.400 311.400 ;
        RECT 696.600 298.350 699.300 299.400 ;
        RECT 683.100 293.100 684.900 293.850 ;
        RECT 695.100 293.100 696.900 293.850 ;
        RECT 697.950 293.100 699.300 298.350 ;
        RECT 710.700 298.350 713.400 299.400 ;
        RECT 701.100 296.100 702.900 296.850 ;
        RECT 707.100 296.100 708.900 296.850 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 694.950 289.950 697.050 292.050 ;
        RECT 698.100 288.900 699.300 293.100 ;
        RECT 700.950 292.950 703.050 295.050 ;
        RECT 706.950 292.950 709.050 295.050 ;
        RECT 710.700 293.100 712.050 298.350 ;
        RECT 727.950 296.100 729.150 299.400 ;
        RECT 713.100 293.100 714.900 293.850 ;
        RECT 697.950 287.100 699.300 288.900 ;
        RECT 710.700 288.900 711.900 293.100 ;
        RECT 724.950 292.950 727.050 295.050 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 728.100 291.900 729.150 296.100 ;
        RECT 749.850 296.100 751.050 299.400 ;
        RECT 767.700 298.350 770.400 299.400 ;
        RECT 785.400 305.400 787.200 311.400 ;
        RECT 799.800 305.400 801.600 311.400 ;
        RECT 764.100 296.100 765.900 296.850 ;
        RECT 730.950 292.950 733.050 295.050 ;
        RECT 745.950 292.950 748.050 295.050 ;
        RECT 749.850 291.900 750.900 296.100 ;
        RECT 751.950 292.950 754.050 295.050 ;
        RECT 757.950 294.450 762.000 295.050 ;
        RECT 763.950 294.450 766.050 295.050 ;
        RECT 757.950 293.550 766.050 294.450 ;
        RECT 757.950 292.950 762.000 293.550 ;
        RECT 763.950 292.950 766.050 293.550 ;
        RECT 767.700 293.100 769.050 298.350 ;
        RECT 785.400 296.100 786.600 305.400 ;
        RECT 796.950 295.950 799.050 298.050 ;
        RECT 775.950 294.450 778.050 295.200 ;
        RECT 784.950 294.450 787.050 295.050 ;
        RECT 770.100 293.100 771.900 293.850 ;
        RECT 775.950 293.550 787.050 294.450 ;
        RECT 797.100 294.150 798.900 294.900 ;
        RECT 775.950 293.100 778.050 293.550 ;
        RECT 725.100 291.150 726.900 291.900 ;
        RECT 722.100 290.100 723.900 290.850 ;
        RECT 727.950 290.100 729.150 291.900 ;
        RECT 731.100 291.150 732.900 291.900 ;
        RECT 746.100 291.150 747.900 291.900 ;
        RECT 749.850 290.100 751.050 291.900 ;
        RECT 752.100 291.150 753.900 291.900 ;
        RECT 755.100 290.100 756.900 290.850 ;
        RECT 710.700 287.100 712.050 288.900 ;
        RECT 721.950 286.950 724.050 289.050 ;
        RECT 727.950 286.950 730.050 289.050 ;
        RECT 733.950 288.450 736.050 289.050 ;
        RECT 748.950 288.450 751.050 289.050 ;
        RECT 733.950 287.550 751.050 288.450 ;
        RECT 733.950 286.950 736.050 287.550 ;
        RECT 748.950 286.950 751.050 287.550 ;
        RECT 754.950 286.950 757.050 289.050 ;
        RECT 767.700 288.900 768.900 293.100 ;
        RECT 784.950 292.950 787.050 293.550 ;
        RECT 800.400 293.100 801.600 305.400 ;
        RECT 802.950 297.450 805.050 298.050 ;
        RECT 808.950 297.450 811.050 301.050 ;
        RECT 817.500 299.400 819.300 311.400 ;
        RECT 802.950 297.000 811.050 297.450 ;
        RECT 802.950 296.550 810.450 297.000 ;
        RECT 802.950 295.950 805.050 296.550 ;
        RECT 817.950 296.100 819.150 299.400 ;
        RECT 803.100 294.150 804.900 294.900 ;
        RECT 814.950 292.950 817.050 295.050 ;
        RECT 805.950 292.050 808.050 292.200 ;
        RECT 769.950 289.950 772.050 292.050 ;
        RECT 782.100 290.100 783.900 290.850 ;
        RECT 767.700 287.100 769.050 288.900 ;
        RECT 775.950 288.450 780.000 289.050 ;
        RECT 781.950 288.450 784.050 289.050 ;
        RECT 775.950 287.550 784.050 288.450 ;
        RECT 775.950 286.950 780.000 287.550 ;
        RECT 781.950 286.950 784.050 287.550 ;
        RECT 697.950 285.450 700.050 286.050 ;
        RECT 677.100 284.400 684.600 285.300 ;
        RECT 686.550 285.000 700.050 285.450 ;
        RECT 677.100 283.500 678.900 284.400 ;
        RECT 675.150 280.800 677.100 282.600 ;
        RECT 675.300 276.600 677.100 280.800 ;
        RECT 682.800 276.600 684.600 284.400 ;
        RECT 685.950 284.550 700.050 285.000 ;
        RECT 685.950 280.950 688.050 284.550 ;
        RECT 697.950 283.950 700.050 284.550 ;
        RECT 709.950 285.450 712.050 286.050 ;
        RECT 714.000 285.900 717.000 286.050 ;
        RECT 714.000 285.450 718.050 285.900 ;
        RECT 709.950 284.550 718.050 285.450 ;
        RECT 728.850 285.750 730.050 285.900 ;
        RECT 748.950 285.750 750.150 285.900 ;
        RECT 728.850 284.700 732.600 285.750 ;
        RECT 709.950 283.950 712.050 284.550 ;
        RECT 714.000 283.950 718.050 284.550 ;
        RECT 715.950 283.800 718.050 283.950 ;
        RECT 698.400 279.600 699.600 282.900 ;
        RECT 697.800 276.600 699.600 279.600 ;
        RECT 710.400 279.600 711.600 282.900 ;
        RECT 722.400 281.700 730.200 283.050 ;
        RECT 710.400 276.600 712.200 279.600 ;
        RECT 722.400 276.600 724.200 281.700 ;
        RECT 728.400 276.600 730.200 281.700 ;
        RECT 731.400 282.600 732.600 284.700 ;
        RECT 746.400 284.700 750.150 285.750 ;
        RECT 746.400 282.600 747.600 284.700 ;
        RECT 766.950 283.950 772.050 286.050 ;
        RECT 731.400 276.600 733.200 282.600 ;
        RECT 745.800 276.600 747.600 282.600 ;
        RECT 748.800 281.700 756.600 283.050 ;
        RECT 748.800 276.600 750.600 281.700 ;
        RECT 754.800 276.600 756.600 281.700 ;
        RECT 767.400 279.600 768.600 282.900 ;
        RECT 785.400 279.600 786.600 291.900 ;
        RECT 799.950 291.450 802.050 292.050 ;
        RECT 804.000 291.450 808.050 292.050 ;
        RECT 818.100 291.900 819.150 296.100 ;
        RECT 820.950 292.950 823.050 295.050 ;
        RECT 799.950 290.550 808.050 291.450 ;
        RECT 815.100 291.150 816.900 291.900 ;
        RECT 799.950 289.950 802.050 290.550 ;
        RECT 804.000 290.100 808.050 290.550 ;
        RECT 812.100 290.100 813.900 290.850 ;
        RECT 817.950 290.100 819.150 291.900 ;
        RECT 821.100 291.150 822.900 291.900 ;
        RECT 804.000 289.950 807.000 290.100 ;
        RECT 800.400 284.700 801.600 288.900 ;
        RECT 811.950 286.950 814.050 289.050 ;
        RECT 817.950 286.950 820.050 289.050 ;
        RECT 818.850 285.750 820.050 285.900 ;
        RECT 818.850 284.700 822.600 285.750 ;
        RECT 798.000 283.800 801.600 284.700 ;
        RECT 767.400 276.600 769.200 279.600 ;
        RECT 785.400 276.600 787.200 279.600 ;
        RECT 798.000 276.600 799.800 283.800 ;
        RECT 812.400 281.700 820.200 283.050 ;
        RECT 812.400 276.600 814.200 281.700 ;
        RECT 818.400 276.600 820.200 281.700 ;
        RECT 821.400 282.600 822.600 284.700 ;
        RECT 821.400 276.600 823.200 282.600 ;
        RECT 3.150 266.400 4.950 272.400 ;
        RECT 10.950 270.300 12.750 272.400 ;
        RECT 9.000 269.400 12.750 270.300 ;
        RECT 18.750 269.400 20.550 272.400 ;
        RECT 26.550 269.400 28.350 272.400 ;
        RECT 9.000 268.500 10.050 269.400 ;
        RECT 7.950 266.400 10.050 268.500 ;
        RECT 18.750 267.600 19.800 269.400 ;
        RECT 3.150 251.700 4.050 266.400 ;
        RECT 11.550 265.800 13.350 267.600 ;
        RECT 14.850 266.550 19.800 267.600 ;
        RECT 27.300 268.500 28.350 269.400 ;
        RECT 27.300 267.300 31.050 268.500 ;
        RECT 14.850 265.800 16.650 266.550 ;
        RECT 28.950 266.400 31.050 267.300 ;
        RECT 34.650 266.400 36.450 272.400 ;
        RECT 46.800 266.400 48.600 272.400 ;
        RECT 11.850 262.800 12.900 265.800 ;
        RECT 6.000 261.600 23.850 262.800 ;
        RECT 35.250 262.050 36.450 266.400 ;
        RECT 47.400 264.300 48.600 266.400 ;
        RECT 49.800 267.300 51.600 272.400 ;
        RECT 55.800 267.300 57.600 272.400 ;
        RECT 49.800 265.950 57.600 267.300 ;
        RECT 68.400 269.400 70.200 272.400 ;
        RECT 83.400 269.400 85.200 272.400 ;
        RECT 47.400 263.250 51.150 264.300 ;
        RECT 49.950 263.100 51.150 263.250 ;
        RECT 6.000 260.850 6.900 261.600 ;
        RECT 11.100 261.000 12.900 261.600 ;
        RECT 22.050 261.000 23.850 261.600 ;
        RECT 5.100 259.050 6.900 260.850 ;
        RECT 22.050 260.100 22.950 261.000 ;
        RECT 30.150 260.250 30.900 262.050 ;
        RECT 31.950 259.950 34.050 262.050 ;
        RECT 35.100 259.950 36.450 262.050 ;
        RECT 43.800 261.450 45.900 262.050 ;
        RECT 8.100 256.800 9.900 257.400 ;
        RECT 8.100 255.600 12.900 256.800 ;
        RECT 13.950 253.950 16.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 12.450 251.700 14.250 252.000 ;
        RECT 3.150 251.100 14.250 251.700 ;
        RECT 3.150 250.500 20.850 251.100 ;
        RECT 3.150 249.600 4.050 250.500 ;
        RECT 12.450 250.200 20.850 250.500 ;
        RECT 3.150 237.600 4.950 249.600 ;
        RECT 17.250 248.700 19.050 249.300 ;
        RECT 11.550 247.500 19.050 248.700 ;
        RECT 19.950 248.100 20.850 250.200 ;
        RECT 22.050 250.200 22.950 255.900 ;
        RECT 32.250 251.400 34.050 253.200 ;
        RECT 28.950 250.200 33.150 251.400 ;
        RECT 22.050 249.300 28.050 250.200 ;
        RECT 28.950 249.300 31.050 250.200 ;
        RECT 35.250 249.600 36.450 259.950 ;
        RECT 38.550 260.550 45.900 261.450 ;
        RECT 38.550 252.900 39.450 260.550 ;
        RECT 43.800 259.950 45.900 260.550 ;
        RECT 46.950 259.950 52.050 262.050 ;
        RECT 55.950 259.950 58.050 262.050 ;
        RECT 64.950 259.950 67.050 262.050 ;
        RECT 47.100 257.100 48.900 257.850 ;
        RECT 50.850 257.100 52.050 258.900 ;
        RECT 56.100 258.150 57.900 258.900 ;
        RECT 65.100 258.150 66.900 258.900 ;
        RECT 53.100 257.100 54.900 257.850 ;
        RECT 68.400 257.100 69.600 269.400 ;
        RECT 79.950 259.950 82.050 262.050 ;
        RECT 80.100 258.150 81.900 258.900 ;
        RECT 83.400 257.100 84.600 269.400 ;
        RECT 90.150 266.400 91.950 272.400 ;
        RECT 97.950 270.300 99.750 272.400 ;
        RECT 96.000 269.400 99.750 270.300 ;
        RECT 105.750 269.400 107.550 272.400 ;
        RECT 113.550 269.400 115.350 272.400 ;
        RECT 96.000 268.500 97.050 269.400 ;
        RECT 94.950 266.400 97.050 268.500 ;
        RECT 105.750 267.600 106.800 269.400 ;
        RECT 46.950 253.950 49.050 256.050 ;
        RECT 50.850 252.900 51.900 257.100 ;
        RECT 52.950 253.950 55.050 256.050 ;
        RECT 67.950 253.950 70.050 256.050 ;
        RECT 82.950 253.950 85.050 256.050 ;
        RECT 37.950 250.800 40.050 252.900 ;
        RECT 50.850 249.600 52.050 252.900 ;
        RECT 27.150 248.400 28.050 249.300 ;
        RECT 24.450 248.100 26.250 248.400 ;
        RECT 11.550 246.600 12.750 247.500 ;
        RECT 19.950 247.200 26.250 248.100 ;
        RECT 24.450 246.600 26.250 247.200 ;
        RECT 27.150 246.600 29.850 248.400 ;
        RECT 7.950 244.500 12.750 246.600 ;
        RECT 15.450 245.550 17.250 246.300 ;
        RECT 20.250 245.550 22.050 246.300 ;
        RECT 15.450 244.500 22.050 245.550 ;
        RECT 11.550 243.600 12.750 244.500 ;
        RECT 11.550 237.600 13.350 243.600 ;
        RECT 19.350 237.600 21.150 244.500 ;
        RECT 27.150 243.600 31.050 245.700 ;
        RECT 27.150 237.600 28.950 243.600 ;
        RECT 34.650 237.600 36.450 249.600 ;
        RECT 50.700 237.600 52.500 249.600 ;
        RECT 68.400 243.600 69.600 252.900 ;
        RECT 83.400 243.600 84.600 252.900 ;
        RECT 90.150 251.700 91.050 266.400 ;
        RECT 98.550 265.800 100.350 267.600 ;
        RECT 101.850 266.550 106.800 267.600 ;
        RECT 114.300 268.500 115.350 269.400 ;
        RECT 114.300 267.300 118.050 268.500 ;
        RECT 101.850 265.800 103.650 266.550 ;
        RECT 115.950 266.400 118.050 267.300 ;
        RECT 121.650 266.400 123.450 272.400 ;
        RECT 98.850 262.800 99.900 265.800 ;
        RECT 93.000 261.600 110.850 262.800 ;
        RECT 122.250 262.050 123.450 266.400 ;
        RECT 134.400 269.400 136.200 272.400 ;
        RECT 93.000 260.850 93.900 261.600 ;
        RECT 98.100 261.000 99.900 261.600 ;
        RECT 109.050 261.000 110.850 261.600 ;
        RECT 92.100 259.050 93.900 260.850 ;
        RECT 109.050 260.100 109.950 261.000 ;
        RECT 117.150 260.250 117.900 262.050 ;
        RECT 118.950 259.950 121.050 262.050 ;
        RECT 122.100 259.950 123.450 262.050 ;
        RECT 130.950 259.950 133.050 262.050 ;
        RECT 95.100 256.800 96.900 257.400 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 95.100 255.600 99.900 256.800 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 99.450 251.700 101.250 252.000 ;
        RECT 90.150 251.100 101.250 251.700 ;
        RECT 90.150 250.500 107.850 251.100 ;
        RECT 90.150 249.600 91.050 250.500 ;
        RECT 99.450 250.200 107.850 250.500 ;
        RECT 68.400 237.600 70.200 243.600 ;
        RECT 83.400 237.600 85.200 243.600 ;
        RECT 90.150 237.600 91.950 249.600 ;
        RECT 104.250 248.700 106.050 249.300 ;
        RECT 98.550 247.500 106.050 248.700 ;
        RECT 106.950 248.100 107.850 250.200 ;
        RECT 109.050 250.200 109.950 255.900 ;
        RECT 119.250 251.400 121.050 253.200 ;
        RECT 115.950 250.200 120.150 251.400 ;
        RECT 109.050 249.300 115.050 250.200 ;
        RECT 115.950 249.300 118.050 250.200 ;
        RECT 122.250 249.600 123.450 259.950 ;
        RECT 131.100 258.150 132.900 258.900 ;
        RECT 134.400 257.100 135.600 269.400 ;
        RECT 141.150 266.400 142.950 272.400 ;
        RECT 148.950 270.300 150.750 272.400 ;
        RECT 147.000 269.400 150.750 270.300 ;
        RECT 156.750 269.400 158.550 272.400 ;
        RECT 164.550 269.400 166.350 272.400 ;
        RECT 147.000 268.500 148.050 269.400 ;
        RECT 145.950 266.400 148.050 268.500 ;
        RECT 156.750 267.600 157.800 269.400 ;
        RECT 133.950 253.950 136.050 256.050 ;
        RECT 114.150 248.400 115.050 249.300 ;
        RECT 111.450 248.100 113.250 248.400 ;
        RECT 98.550 246.600 99.750 247.500 ;
        RECT 106.950 247.200 113.250 248.100 ;
        RECT 111.450 246.600 113.250 247.200 ;
        RECT 114.150 246.600 116.850 248.400 ;
        RECT 94.950 244.500 99.750 246.600 ;
        RECT 102.450 245.550 104.250 246.300 ;
        RECT 107.250 245.550 109.050 246.300 ;
        RECT 102.450 244.500 109.050 245.550 ;
        RECT 98.550 243.600 99.750 244.500 ;
        RECT 98.550 237.600 100.350 243.600 ;
        RECT 106.350 237.600 108.150 244.500 ;
        RECT 114.150 243.600 118.050 245.700 ;
        RECT 114.150 237.600 115.950 243.600 ;
        RECT 121.650 237.600 123.450 249.600 ;
        RECT 134.400 243.600 135.600 252.900 ;
        RECT 141.150 251.700 142.050 266.400 ;
        RECT 149.550 265.800 151.350 267.600 ;
        RECT 152.850 266.550 157.800 267.600 ;
        RECT 165.300 268.500 166.350 269.400 ;
        RECT 165.300 267.300 169.050 268.500 ;
        RECT 152.850 265.800 154.650 266.550 ;
        RECT 166.950 266.400 169.050 267.300 ;
        RECT 172.650 266.400 174.450 272.400 ;
        RECT 149.850 262.800 150.900 265.800 ;
        RECT 144.000 261.600 161.850 262.800 ;
        RECT 173.250 262.050 174.450 266.400 ;
        RECT 179.400 267.300 181.200 272.400 ;
        RECT 185.400 267.300 187.200 272.400 ;
        RECT 179.400 265.950 187.200 267.300 ;
        RECT 188.400 266.400 190.200 272.400 ;
        RECT 202.800 269.400 204.600 272.400 ;
        RECT 188.400 264.300 189.600 266.400 ;
        RECT 185.850 263.250 189.600 264.300 ;
        RECT 185.850 263.100 187.050 263.250 ;
        RECT 144.000 260.850 144.900 261.600 ;
        RECT 149.100 261.000 150.900 261.600 ;
        RECT 160.050 261.000 161.850 261.600 ;
        RECT 143.100 259.050 144.900 260.850 ;
        RECT 160.050 260.100 160.950 261.000 ;
        RECT 168.150 260.250 168.900 262.050 ;
        RECT 169.950 259.950 172.050 262.050 ;
        RECT 173.100 259.950 174.450 262.050 ;
        RECT 178.950 259.950 181.050 262.050 ;
        RECT 184.950 259.950 187.050 262.050 ;
        RECT 146.100 256.800 147.900 257.400 ;
        RECT 146.100 255.600 150.900 256.800 ;
        RECT 151.950 253.950 154.050 259.050 ;
        RECT 157.950 256.950 160.050 259.050 ;
        RECT 150.450 251.700 152.250 252.000 ;
        RECT 141.150 251.100 152.250 251.700 ;
        RECT 141.150 250.500 158.850 251.100 ;
        RECT 141.150 249.600 142.050 250.500 ;
        RECT 150.450 250.200 158.850 250.500 ;
        RECT 134.400 237.600 136.200 243.600 ;
        RECT 141.150 237.600 142.950 249.600 ;
        RECT 155.250 248.700 157.050 249.300 ;
        RECT 149.550 247.500 157.050 248.700 ;
        RECT 157.950 248.100 158.850 250.200 ;
        RECT 160.050 250.200 160.950 255.900 ;
        RECT 170.250 251.400 172.050 253.200 ;
        RECT 166.950 250.200 171.150 251.400 ;
        RECT 160.050 249.300 166.050 250.200 ;
        RECT 166.950 249.300 169.050 250.200 ;
        RECT 173.250 249.600 174.450 259.950 ;
        RECT 179.100 258.150 180.900 258.900 ;
        RECT 182.100 257.100 183.900 257.850 ;
        RECT 184.950 257.100 186.150 258.900 ;
        RECT 188.100 257.100 189.900 257.850 ;
        RECT 203.400 257.100 204.600 269.400 ;
        RECT 218.400 269.400 220.200 272.400 ;
        RECT 235.800 269.400 237.600 272.400 ;
        RECT 218.400 266.100 219.600 269.400 ;
        RECT 217.950 264.450 220.050 265.050 ;
        RECT 232.950 264.450 235.050 265.050 ;
        RECT 217.950 263.550 235.050 264.450 ;
        RECT 217.950 262.950 220.050 263.550 ;
        RECT 232.950 262.950 235.050 263.550 ;
        RECT 205.950 259.950 208.050 262.050 ;
        RECT 218.700 260.100 220.050 261.900 ;
        RECT 206.100 258.150 207.900 258.900 ;
        RECT 181.950 253.950 184.050 256.050 ;
        RECT 185.100 252.900 186.150 257.100 ;
        RECT 187.950 253.950 190.050 256.050 ;
        RECT 202.950 253.950 205.050 256.050 ;
        RECT 211.950 253.950 217.050 256.050 ;
        RECT 218.700 255.900 219.900 260.100 ;
        RECT 220.950 256.950 223.050 259.050 ;
        RECT 236.400 257.100 237.600 269.400 ;
        RECT 251.400 269.400 253.200 272.400 ;
        RECT 266.400 269.400 268.200 272.400 ;
        RECT 284.400 269.400 286.200 272.400 ;
        RECT 296.400 269.400 298.200 272.400 ;
        RECT 251.400 266.100 252.600 269.400 ;
        RECT 266.400 266.100 267.600 269.400 ;
        RECT 250.950 264.450 253.050 265.050 ;
        RECT 259.950 264.450 262.050 265.050 ;
        RECT 250.950 263.550 262.050 264.450 ;
        RECT 250.950 262.950 253.050 263.550 ;
        RECT 259.950 262.950 262.050 263.550 ;
        RECT 265.950 262.950 268.050 265.050 ;
        RECT 238.950 261.450 241.050 262.050 ;
        RECT 243.000 261.450 247.050 262.050 ;
        RECT 238.950 260.550 247.050 261.450 ;
        RECT 238.950 259.950 241.050 260.550 ;
        RECT 243.000 259.950 247.050 260.550 ;
        RECT 251.700 260.100 253.050 261.900 ;
        RECT 266.700 260.100 268.050 261.900 ;
        RECT 239.100 258.150 240.900 258.900 ;
        RECT 184.950 249.600 186.150 252.900 ;
        RECT 165.150 248.400 166.050 249.300 ;
        RECT 162.450 248.100 164.250 248.400 ;
        RECT 149.550 246.600 150.750 247.500 ;
        RECT 157.950 247.200 164.250 248.100 ;
        RECT 162.450 246.600 164.250 247.200 ;
        RECT 165.150 246.600 167.850 248.400 ;
        RECT 145.950 244.500 150.750 246.600 ;
        RECT 153.450 245.550 155.250 246.300 ;
        RECT 158.250 245.550 160.050 246.300 ;
        RECT 153.450 244.500 160.050 245.550 ;
        RECT 149.550 243.600 150.750 244.500 ;
        RECT 149.550 237.600 151.350 243.600 ;
        RECT 157.350 237.600 159.150 244.500 ;
        RECT 165.150 243.600 169.050 245.700 ;
        RECT 165.150 237.600 166.950 243.600 ;
        RECT 172.650 237.600 174.450 249.600 ;
        RECT 184.500 237.600 186.300 249.600 ;
        RECT 203.400 243.600 204.600 252.900 ;
        RECT 215.100 252.150 216.900 252.900 ;
        RECT 218.700 250.650 220.050 255.900 ;
        RECT 221.100 255.150 222.900 255.900 ;
        RECT 226.950 255.450 229.050 256.050 ;
        RECT 235.950 255.450 238.050 256.050 ;
        RECT 226.950 254.550 238.050 255.450 ;
        RECT 226.950 253.950 229.050 254.550 ;
        RECT 235.950 253.950 238.050 254.550 ;
        RECT 241.950 255.450 246.000 256.050 ;
        RECT 247.950 255.450 250.050 256.050 ;
        RECT 241.950 254.550 250.050 255.450 ;
        RECT 241.950 253.950 246.000 254.550 ;
        RECT 247.950 253.950 250.050 254.550 ;
        RECT 251.700 255.900 252.900 260.100 ;
        RECT 253.950 256.950 256.050 259.050 ;
        RECT 205.950 249.450 208.050 250.050 ;
        RECT 211.950 249.450 214.050 250.050 ;
        RECT 218.700 249.600 221.400 250.650 ;
        RECT 205.950 248.550 214.050 249.450 ;
        RECT 205.950 247.950 208.050 248.550 ;
        RECT 211.950 247.950 214.050 248.550 ;
        RECT 202.800 237.600 204.600 243.600 ;
        RECT 219.600 237.600 221.400 249.600 ;
        RECT 236.400 243.600 237.600 252.900 ;
        RECT 248.100 252.150 249.900 252.900 ;
        RECT 251.700 250.650 253.050 255.900 ;
        RECT 254.100 255.150 255.900 255.900 ;
        RECT 262.950 253.950 265.050 256.050 ;
        RECT 266.700 255.900 267.900 260.100 ;
        RECT 280.950 259.950 283.050 262.050 ;
        RECT 268.950 256.950 271.050 259.050 ;
        RECT 281.100 258.150 282.900 258.900 ;
        RECT 284.400 257.100 285.600 269.400 ;
        RECT 296.400 266.100 297.600 269.400 ;
        RECT 311.400 267.300 313.200 272.400 ;
        RECT 317.400 267.300 319.200 272.400 ;
        RECT 311.400 265.950 319.200 267.300 ;
        RECT 320.400 266.400 322.200 272.400 ;
        RECT 332.400 269.400 334.200 272.400 ;
        RECT 286.950 264.450 289.050 265.050 ;
        RECT 295.950 264.450 298.050 265.050 ;
        RECT 286.950 263.550 298.050 264.450 ;
        RECT 320.400 264.300 321.600 266.400 ;
        RECT 286.950 262.950 289.050 263.550 ;
        RECT 295.950 262.950 298.050 263.550 ;
        RECT 317.850 263.250 321.600 264.300 ;
        RECT 317.850 263.100 319.050 263.250 ;
        RECT 296.700 260.100 298.050 261.900 ;
        RECT 263.100 252.150 264.900 252.900 ;
        RECT 266.700 250.650 268.050 255.900 ;
        RECT 269.100 255.150 270.900 255.900 ;
        RECT 283.950 253.950 286.050 256.050 ;
        RECT 292.950 253.950 295.050 256.050 ;
        RECT 296.700 255.900 297.900 260.100 ;
        RECT 310.950 259.950 313.050 262.050 ;
        RECT 316.950 261.450 319.050 262.050 ;
        RECT 321.000 261.450 325.050 262.050 ;
        RECT 316.950 260.550 325.050 261.450 ;
        RECT 316.950 259.950 319.050 260.550 ;
        RECT 321.000 259.950 325.050 260.550 ;
        RECT 328.950 259.950 331.050 262.200 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 311.100 258.150 312.900 258.900 ;
        RECT 314.100 257.100 315.900 257.850 ;
        RECT 316.950 257.100 318.150 258.900 ;
        RECT 329.100 258.150 330.900 258.900 ;
        RECT 320.100 257.100 321.900 257.850 ;
        RECT 332.400 257.100 333.600 269.400 ;
        RECT 349.200 265.200 351.000 272.400 ;
        RECT 347.400 264.300 351.000 265.200 ;
        RECT 356.550 266.400 358.350 272.400 ;
        RECT 364.650 269.400 366.450 272.400 ;
        RECT 372.450 269.400 374.250 272.400 ;
        RECT 380.250 270.300 382.050 272.400 ;
        RECT 380.250 269.400 384.000 270.300 ;
        RECT 364.650 268.500 365.700 269.400 ;
        RECT 361.950 267.300 365.700 268.500 ;
        RECT 373.200 267.600 374.250 269.400 ;
        RECT 382.950 268.500 384.000 269.400 ;
        RECT 361.950 266.400 364.050 267.300 ;
        RECT 373.200 266.550 378.150 267.600 ;
        RECT 347.400 260.100 348.600 264.300 ;
        RECT 356.550 262.050 357.750 266.400 ;
        RECT 376.350 265.800 378.150 266.550 ;
        RECT 379.650 265.800 381.450 267.600 ;
        RECT 382.950 266.400 385.050 268.500 ;
        RECT 388.050 266.400 389.850 272.400 ;
        RECT 400.800 266.400 402.600 272.400 ;
        RECT 380.100 262.800 381.150 265.800 ;
        RECT 356.550 259.950 357.900 262.050 ;
        RECT 358.950 259.950 361.050 262.050 ;
        RECT 362.100 260.250 362.850 262.050 ;
        RECT 369.150 261.600 387.000 262.800 ;
        RECT 369.150 261.000 370.950 261.600 ;
        RECT 380.100 261.000 381.900 261.600 ;
        RECT 370.050 260.100 370.950 261.000 ;
        RECT 386.100 260.850 387.000 261.600 ;
        RECT 337.950 258.450 340.050 259.050 ;
        RECT 346.950 258.450 349.050 259.050 ;
        RECT 337.950 257.550 349.050 258.450 ;
        RECT 251.700 249.600 254.400 250.650 ;
        RECT 266.700 249.600 269.400 250.650 ;
        RECT 235.800 237.600 237.600 243.600 ;
        RECT 252.600 237.600 254.400 249.600 ;
        RECT 267.600 237.600 269.400 249.600 ;
        RECT 284.400 243.600 285.600 252.900 ;
        RECT 293.100 252.150 294.900 252.900 ;
        RECT 296.700 250.650 298.050 255.900 ;
        RECT 299.100 255.150 300.900 255.900 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 317.100 252.900 318.150 257.100 ;
        RECT 337.950 256.950 340.050 257.550 ;
        RECT 346.950 256.950 349.050 257.550 ;
        RECT 319.950 253.950 322.050 256.050 ;
        RECT 331.950 255.450 334.050 256.050 ;
        RECT 326.550 255.000 334.050 255.450 ;
        RECT 325.950 254.550 334.050 255.000 ;
        RECT 296.700 249.600 299.400 250.650 ;
        RECT 316.950 249.600 318.150 252.900 ;
        RECT 325.950 250.950 328.050 254.550 ;
        RECT 331.950 253.950 334.050 254.550 ;
        RECT 344.100 254.100 345.900 254.850 ;
        RECT 284.400 237.600 286.200 243.600 ;
        RECT 297.600 237.600 299.400 249.600 ;
        RECT 316.500 237.600 318.300 249.600 ;
        RECT 332.400 243.600 333.600 252.900 ;
        RECT 343.950 250.950 346.050 253.050 ;
        RECT 347.400 243.600 348.600 255.900 ;
        RECT 350.100 254.100 351.900 254.850 ;
        RECT 349.950 250.950 352.050 253.050 ;
        RECT 356.550 249.600 357.750 259.950 ;
        RECT 386.100 259.050 387.900 260.850 ;
        RECT 370.950 256.950 373.050 259.050 ;
        RECT 383.100 256.800 384.900 257.400 ;
        RECT 358.950 251.400 360.750 253.200 ;
        RECT 359.850 250.200 364.050 251.400 ;
        RECT 370.050 250.200 370.950 255.900 ;
        RECT 376.950 253.950 379.050 256.050 ;
        RECT 380.100 255.600 384.900 256.800 ;
        RECT 378.750 251.700 380.550 252.000 ;
        RECT 388.950 251.700 389.850 266.400 ;
        RECT 401.400 264.300 402.600 266.400 ;
        RECT 403.800 267.300 405.600 272.400 ;
        RECT 409.800 267.300 411.600 272.400 ;
        RECT 403.800 265.950 411.600 267.300 ;
        RECT 418.800 266.400 420.600 272.400 ;
        RECT 419.400 264.300 420.600 266.400 ;
        RECT 421.800 267.300 423.600 272.400 ;
        RECT 427.800 267.300 429.600 272.400 ;
        RECT 440.400 269.400 442.200 272.400 ;
        RECT 421.800 265.950 429.600 267.300 ;
        RECT 401.400 263.250 405.150 264.300 ;
        RECT 419.400 263.250 423.150 264.300 ;
        RECT 436.950 264.000 439.050 268.050 ;
        RECT 403.950 263.100 405.150 263.250 ;
        RECT 421.950 263.100 423.150 263.250 ;
        RECT 437.550 262.050 438.450 264.000 ;
        RECT 403.950 259.950 406.050 262.050 ;
        RECT 409.950 259.950 412.050 262.050 ;
        RECT 415.950 261.450 420.000 262.050 ;
        RECT 421.950 261.450 424.050 262.050 ;
        RECT 415.950 260.550 424.050 261.450 ;
        RECT 415.950 259.950 420.000 260.550 ;
        RECT 421.950 259.950 424.050 260.550 ;
        RECT 427.950 259.950 430.050 262.050 ;
        RECT 436.950 259.950 439.050 262.050 ;
        RECT 401.100 257.100 402.900 257.850 ;
        RECT 404.850 257.100 406.050 258.900 ;
        RECT 410.100 258.150 411.900 258.900 ;
        RECT 407.100 257.100 408.900 257.850 ;
        RECT 419.100 257.100 420.900 257.850 ;
        RECT 422.850 257.100 424.050 258.900 ;
        RECT 428.100 258.150 429.900 258.900 ;
        RECT 437.100 258.150 438.900 258.900 ;
        RECT 425.100 257.100 426.900 257.850 ;
        RECT 440.400 257.100 441.600 269.400 ;
        RECT 454.800 266.400 456.600 272.400 ;
        RECT 455.400 264.300 456.600 266.400 ;
        RECT 457.800 267.300 459.600 272.400 ;
        RECT 463.800 267.300 465.600 272.400 ;
        RECT 457.800 265.950 465.600 267.300 ;
        RECT 473.400 269.400 475.200 272.400 ;
        RECT 473.400 266.100 474.600 269.400 ;
        RECT 490.800 266.400 492.600 272.400 ;
        RECT 455.400 263.250 459.150 264.300 ;
        RECT 457.950 263.100 459.150 263.250 ;
        RECT 472.950 262.950 475.050 265.050 ;
        RECT 491.400 264.300 492.600 266.400 ;
        RECT 493.800 267.300 495.600 272.400 ;
        RECT 499.800 267.300 501.600 272.400 ;
        RECT 511.800 269.400 513.600 272.400 ;
        RECT 493.800 265.950 501.600 267.300 ;
        RECT 491.400 263.250 495.150 264.300 ;
        RECT 493.950 263.100 495.150 263.250 ;
        RECT 457.950 259.950 460.050 262.050 ;
        RECT 463.950 259.950 466.050 262.050 ;
        RECT 473.700 260.100 475.050 261.900 ;
        RECT 455.100 257.100 456.900 257.850 ;
        RECT 458.850 257.100 460.050 258.900 ;
        RECT 464.100 258.150 465.900 258.900 ;
        RECT 461.100 257.100 462.900 257.850 ;
        RECT 391.950 255.450 394.050 256.050 ;
        RECT 400.950 255.450 403.050 256.050 ;
        RECT 391.950 254.550 403.050 255.450 ;
        RECT 391.950 253.950 394.050 254.550 ;
        RECT 400.950 253.950 403.050 254.550 ;
        RECT 378.750 251.100 389.850 251.700 ;
        RECT 332.400 237.600 334.200 243.600 ;
        RECT 347.400 237.600 349.200 243.600 ;
        RECT 356.550 237.600 358.350 249.600 ;
        RECT 361.950 249.300 364.050 250.200 ;
        RECT 364.950 249.300 370.950 250.200 ;
        RECT 372.150 250.500 389.850 251.100 ;
        RECT 372.150 250.200 380.550 250.500 ;
        RECT 364.950 248.400 365.850 249.300 ;
        RECT 363.150 246.600 365.850 248.400 ;
        RECT 366.750 248.100 368.550 248.400 ;
        RECT 372.150 248.100 373.050 250.200 ;
        RECT 388.950 249.600 389.850 250.500 ;
        RECT 404.850 252.900 405.900 257.100 ;
        RECT 406.950 253.950 409.050 256.050 ;
        RECT 418.950 253.950 421.050 256.050 ;
        RECT 422.850 252.900 423.900 257.100 ;
        RECT 424.950 253.950 427.050 256.050 ;
        RECT 436.950 253.950 442.050 256.050 ;
        RECT 451.950 253.950 457.050 256.050 ;
        RECT 458.850 252.900 459.900 257.100 ;
        RECT 460.950 255.900 465.450 256.050 ;
        RECT 460.950 253.950 466.050 255.900 ;
        RECT 469.950 253.950 472.050 256.050 ;
        RECT 473.700 255.900 474.900 260.100 ;
        RECT 493.950 259.950 496.050 262.050 ;
        RECT 499.950 261.450 502.050 262.200 ;
        RECT 508.950 261.450 511.050 262.050 ;
        RECT 499.950 260.550 511.050 261.450 ;
        RECT 499.950 259.950 502.050 260.550 ;
        RECT 508.950 259.950 511.050 260.550 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 491.100 257.100 492.900 257.850 ;
        RECT 494.850 257.100 496.050 258.900 ;
        RECT 500.100 258.150 501.900 258.900 ;
        RECT 497.100 257.100 498.900 257.850 ;
        RECT 512.400 257.100 513.600 269.400 ;
        RECT 518.550 266.400 520.350 272.400 ;
        RECT 526.650 269.400 528.450 272.400 ;
        RECT 534.450 269.400 536.250 272.400 ;
        RECT 542.250 270.300 544.050 272.400 ;
        RECT 542.250 269.400 546.000 270.300 ;
        RECT 526.650 268.500 527.700 269.400 ;
        RECT 523.950 267.300 527.700 268.500 ;
        RECT 535.200 267.600 536.250 269.400 ;
        RECT 544.950 268.500 546.000 269.400 ;
        RECT 523.950 266.400 526.050 267.300 ;
        RECT 535.200 266.550 540.150 267.600 ;
        RECT 518.550 262.050 519.750 266.400 ;
        RECT 538.350 265.800 540.150 266.550 ;
        RECT 541.650 265.800 543.450 267.600 ;
        RECT 544.950 266.400 547.050 268.500 ;
        RECT 550.050 266.400 551.850 272.400 ;
        RECT 542.100 262.800 543.150 265.800 ;
        RECT 514.950 259.950 517.050 262.050 ;
        RECT 518.550 259.950 519.900 262.050 ;
        RECT 520.950 259.950 523.050 262.050 ;
        RECT 524.100 260.250 524.850 262.050 ;
        RECT 531.150 261.600 549.000 262.800 ;
        RECT 531.150 261.000 532.950 261.600 ;
        RECT 542.100 261.000 543.900 261.600 ;
        RECT 532.050 260.100 532.950 261.000 ;
        RECT 548.100 260.850 549.000 261.600 ;
        RECT 515.100 258.150 516.900 258.900 ;
        RECT 463.950 253.800 466.050 253.950 ;
        RECT 404.850 249.600 406.050 252.900 ;
        RECT 422.850 249.600 424.050 252.900 ;
        RECT 366.750 247.200 373.050 248.100 ;
        RECT 373.950 248.700 375.750 249.300 ;
        RECT 373.950 247.500 381.450 248.700 ;
        RECT 366.750 246.600 368.550 247.200 ;
        RECT 380.250 246.600 381.450 247.500 ;
        RECT 361.950 243.600 365.850 245.700 ;
        RECT 370.950 245.550 372.750 246.300 ;
        RECT 375.750 245.550 377.550 246.300 ;
        RECT 370.950 244.500 377.550 245.550 ;
        RECT 380.250 244.500 385.050 246.600 ;
        RECT 364.050 237.600 365.850 243.600 ;
        RECT 371.850 237.600 373.650 244.500 ;
        RECT 380.250 243.600 381.450 244.500 ;
        RECT 379.650 237.600 381.450 243.600 ;
        RECT 388.050 237.600 389.850 249.600 ;
        RECT 404.700 237.600 406.500 249.600 ;
        RECT 422.700 237.600 424.500 249.600 ;
        RECT 440.400 243.600 441.600 252.900 ;
        RECT 458.850 249.600 460.050 252.900 ;
        RECT 470.100 252.150 471.900 252.900 ;
        RECT 473.700 250.650 475.050 255.900 ;
        RECT 476.100 255.150 477.900 255.900 ;
        RECT 490.950 253.950 493.050 256.050 ;
        RECT 494.850 252.900 495.900 257.100 ;
        RECT 496.950 255.450 499.050 256.050 ;
        RECT 511.950 255.450 514.050 256.050 ;
        RECT 496.950 254.550 514.050 255.450 ;
        RECT 496.950 253.950 499.050 254.550 ;
        RECT 511.950 253.950 514.050 254.550 ;
        RECT 473.700 249.600 476.400 250.650 ;
        RECT 494.850 249.600 496.050 252.900 ;
        RECT 440.400 237.600 442.200 243.600 ;
        RECT 458.700 237.600 460.500 249.600 ;
        RECT 474.600 237.600 476.400 249.600 ;
        RECT 494.700 237.600 496.500 249.600 ;
        RECT 512.400 243.600 513.600 252.900 ;
        RECT 511.800 237.600 513.600 243.600 ;
        RECT 518.550 249.600 519.750 259.950 ;
        RECT 548.100 259.050 549.900 260.850 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 545.100 256.800 546.900 257.400 ;
        RECT 520.950 251.400 522.750 253.200 ;
        RECT 521.850 250.200 526.050 251.400 ;
        RECT 532.050 250.200 532.950 255.900 ;
        RECT 538.950 253.950 541.050 256.050 ;
        RECT 542.100 255.600 546.900 256.800 ;
        RECT 540.750 251.700 542.550 252.000 ;
        RECT 550.950 251.700 551.850 266.400 ;
        RECT 560.400 269.400 562.200 272.400 ;
        RECT 560.400 266.100 561.600 269.400 ;
        RECT 580.200 268.050 582.000 272.400 ;
        RECT 598.800 269.400 600.600 272.400 ;
        RECT 559.950 264.450 562.050 265.050 ;
        RECT 565.950 264.450 568.050 268.050 ;
        RECT 580.200 266.400 585.600 268.050 ;
        RECT 559.950 264.000 568.050 264.450 ;
        RECT 559.950 263.550 567.450 264.000 ;
        RECT 559.950 262.950 562.050 263.550 ;
        RECT 584.700 263.100 585.600 266.400 ;
        RECT 560.700 260.100 562.050 261.900 ;
        RECT 556.950 253.950 559.050 256.050 ;
        RECT 560.700 255.900 561.900 260.100 ;
        RECT 577.950 259.950 580.050 262.050 ;
        RECT 583.950 261.450 586.050 262.050 ;
        RECT 595.950 261.450 598.050 262.050 ;
        RECT 583.950 260.550 598.050 261.450 ;
        RECT 583.950 259.950 586.050 260.550 ;
        RECT 595.950 259.950 598.050 260.550 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 578.100 258.150 579.900 258.900 ;
        RECT 575.100 257.100 576.900 257.850 ;
        RECT 581.100 257.100 582.900 257.850 ;
        RECT 557.100 252.150 558.900 252.900 ;
        RECT 540.750 251.100 551.850 251.700 ;
        RECT 518.550 237.600 520.350 249.600 ;
        RECT 523.950 249.300 526.050 250.200 ;
        RECT 526.950 249.300 532.950 250.200 ;
        RECT 534.150 250.500 551.850 251.100 ;
        RECT 534.150 250.200 542.550 250.500 ;
        RECT 526.950 248.400 527.850 249.300 ;
        RECT 525.150 246.600 527.850 248.400 ;
        RECT 528.750 248.100 530.550 248.400 ;
        RECT 534.150 248.100 535.050 250.200 ;
        RECT 550.950 249.600 551.850 250.500 ;
        RECT 560.700 250.650 562.050 255.900 ;
        RECT 563.100 255.150 564.900 255.900 ;
        RECT 574.950 253.950 577.050 256.050 ;
        RECT 580.950 253.950 583.050 256.050 ;
        RECT 560.700 249.600 563.400 250.650 ;
        RECT 584.700 249.600 585.600 258.900 ;
        RECT 599.400 257.100 600.600 269.400 ;
        RECT 610.800 266.400 612.600 272.400 ;
        RECT 601.950 259.950 604.050 262.050 ;
        RECT 607.950 261.450 610.050 265.050 ;
        RECT 611.400 264.300 612.600 266.400 ;
        RECT 613.800 267.300 615.600 272.400 ;
        RECT 619.800 267.300 621.600 272.400 ;
        RECT 613.800 265.950 621.600 267.300 ;
        RECT 629.400 269.400 631.200 272.400 ;
        RECT 644.400 269.400 646.200 272.400 ;
        RECT 656.400 269.400 658.200 272.400 ;
        RECT 611.400 263.250 615.150 264.300 ;
        RECT 613.950 263.100 615.150 263.250 ;
        RECT 613.950 261.450 616.050 262.050 ;
        RECT 607.950 261.000 616.050 261.450 ;
        RECT 608.550 260.550 616.050 261.000 ;
        RECT 613.950 259.950 616.050 260.550 ;
        RECT 619.950 259.950 622.050 262.050 ;
        RECT 625.950 259.950 628.050 262.050 ;
        RECT 602.100 258.150 603.900 258.900 ;
        RECT 611.100 257.100 612.900 257.850 ;
        RECT 614.850 257.100 616.050 258.900 ;
        RECT 620.100 258.150 621.900 258.900 ;
        RECT 626.100 258.150 627.900 258.900 ;
        RECT 617.100 257.100 618.900 257.850 ;
        RECT 629.400 257.100 630.600 269.400 ;
        RECT 640.950 259.950 643.050 262.050 ;
        RECT 641.100 258.150 642.900 258.900 ;
        RECT 644.400 257.100 645.600 269.400 ;
        RECT 656.400 266.100 657.600 269.400 ;
        RECT 655.950 264.450 658.050 265.050 ;
        RECT 664.950 264.450 667.050 265.050 ;
        RECT 655.950 263.550 667.050 264.450 ;
        RECT 668.400 264.600 670.200 272.400 ;
        RECT 675.900 268.200 677.700 272.400 ;
        RECT 675.900 266.400 677.850 268.200 ;
        RECT 674.100 264.600 675.900 265.500 ;
        RECT 668.400 263.700 675.900 264.600 ;
        RECT 655.950 262.950 658.050 263.550 ;
        RECT 664.950 262.950 667.050 263.550 ;
        RECT 656.700 260.100 658.050 261.900 ;
        RECT 598.950 255.450 601.050 256.050 ;
        RECT 598.950 255.000 606.450 255.450 ;
        RECT 598.950 254.550 607.050 255.000 ;
        RECT 598.950 253.950 601.050 254.550 ;
        RECT 528.750 247.200 535.050 248.100 ;
        RECT 535.950 248.700 537.750 249.300 ;
        RECT 535.950 247.500 543.450 248.700 ;
        RECT 528.750 246.600 530.550 247.200 ;
        RECT 542.250 246.600 543.450 247.500 ;
        RECT 523.950 243.600 527.850 245.700 ;
        RECT 532.950 245.550 534.750 246.300 ;
        RECT 537.750 245.550 539.550 246.300 ;
        RECT 532.950 244.500 539.550 245.550 ;
        RECT 542.250 244.500 547.050 246.600 ;
        RECT 526.050 237.600 527.850 243.600 ;
        RECT 533.850 237.600 535.650 244.500 ;
        RECT 542.250 243.600 543.450 244.500 ;
        RECT 541.650 237.600 543.450 243.600 ;
        RECT 550.050 237.600 551.850 249.600 ;
        RECT 561.600 237.600 563.400 249.600 ;
        RECT 575.400 248.700 583.200 249.600 ;
        RECT 575.400 237.600 577.200 248.700 ;
        RECT 581.400 237.600 583.200 248.700 ;
        RECT 584.400 237.600 586.200 249.600 ;
        RECT 599.400 243.600 600.600 252.900 ;
        RECT 604.950 250.950 607.050 254.550 ;
        RECT 610.950 253.950 613.050 256.050 ;
        RECT 614.850 252.900 615.900 257.100 ;
        RECT 616.950 253.950 619.050 256.050 ;
        RECT 628.950 255.450 631.050 256.050 ;
        RECT 637.950 255.450 640.050 256.050 ;
        RECT 628.950 254.550 640.050 255.450 ;
        RECT 628.950 253.950 631.050 254.550 ;
        RECT 637.950 253.950 640.050 254.550 ;
        RECT 643.950 253.950 646.050 256.050 ;
        RECT 652.950 253.950 655.050 256.050 ;
        RECT 656.700 255.900 657.900 260.100 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 667.950 256.950 670.050 259.050 ;
        RECT 614.850 249.600 616.050 252.900 ;
        RECT 598.800 237.600 600.600 243.600 ;
        RECT 614.700 237.600 616.500 249.600 ;
        RECT 629.400 243.600 630.600 252.900 ;
        RECT 644.400 243.600 645.600 252.900 ;
        RECT 653.100 252.150 654.900 252.900 ;
        RECT 656.700 250.650 658.050 255.900 ;
        RECT 659.100 255.150 660.900 255.900 ;
        RECT 668.100 255.150 669.900 255.900 ;
        RECT 656.700 249.600 659.400 250.650 ;
        RECT 629.400 237.600 631.200 243.600 ;
        RECT 644.400 237.600 646.200 243.600 ;
        RECT 657.600 237.600 659.400 249.600 ;
        RECT 671.400 243.600 672.450 263.700 ;
        RECT 676.950 263.100 677.850 266.400 ;
        RECT 691.200 265.200 693.000 272.400 ;
        RECT 709.200 268.050 711.000 272.400 ;
        RECT 709.200 266.400 714.600 268.050 ;
        RECT 689.400 264.300 693.000 265.200 ;
        RECT 676.950 261.450 679.050 262.050 ;
        RECT 681.000 261.450 685.050 262.050 ;
        RECT 676.950 260.550 685.050 261.450 ;
        RECT 676.950 259.950 679.050 260.550 ;
        RECT 681.000 259.950 685.050 260.550 ;
        RECT 689.400 260.100 690.600 264.300 ;
        RECT 713.700 263.100 714.600 266.400 ;
        RECT 730.200 265.200 732.000 272.400 ;
        RECT 748.200 265.200 750.000 272.400 ;
        RECT 766.800 269.400 768.600 272.400 ;
        RECT 767.400 266.100 768.600 269.400 ;
        RECT 786.000 268.050 787.800 272.400 ;
        RECT 782.400 266.400 787.800 268.050 ;
        RECT 794.550 266.400 796.350 272.400 ;
        RECT 802.650 269.400 804.450 272.400 ;
        RECT 810.450 269.400 812.250 272.400 ;
        RECT 818.250 270.300 820.050 272.400 ;
        RECT 818.250 269.400 822.000 270.300 ;
        RECT 802.650 268.500 803.700 269.400 ;
        RECT 799.950 267.300 803.700 268.500 ;
        RECT 811.200 267.600 812.250 269.400 ;
        RECT 820.950 268.500 822.000 269.400 ;
        RECT 799.950 266.400 802.050 267.300 ;
        RECT 811.200 266.550 816.150 267.600 ;
        RECT 728.400 264.300 732.000 265.200 ;
        RECT 746.400 264.300 750.000 265.200 ;
        RECT 760.950 264.450 765.000 265.050 ;
        RECT 766.950 264.450 769.050 265.050 ;
        RECT 706.950 259.950 709.050 262.050 ;
        RECT 712.950 259.950 715.050 262.050 ;
        RECT 728.400 260.100 729.600 264.300 ;
        RECT 746.400 260.100 747.600 264.300 ;
        RECT 760.950 263.550 769.050 264.450 ;
        RECT 760.950 262.950 765.000 263.550 ;
        RECT 766.950 262.950 769.050 263.550 ;
        RECT 782.400 263.100 783.300 266.400 ;
        RECT 794.550 262.050 795.750 266.400 ;
        RECT 814.350 265.800 816.150 266.550 ;
        RECT 817.650 265.800 819.450 267.600 ;
        RECT 820.950 266.400 823.050 268.500 ;
        RECT 826.050 266.400 827.850 272.400 ;
        RECT 818.100 262.800 819.150 265.800 ;
        RECT 766.950 260.100 768.300 261.900 ;
        RECT 674.100 257.100 675.900 257.850 ;
        RECT 673.950 253.950 676.050 256.050 ;
        RECT 678.000 249.600 679.050 258.900 ;
        RECT 688.950 258.450 691.050 259.050 ;
        RECT 697.950 258.450 700.050 259.050 ;
        RECT 688.950 257.550 700.050 258.450 ;
        RECT 707.100 258.150 708.900 258.900 ;
        RECT 688.950 256.950 691.050 257.550 ;
        RECT 697.950 256.950 700.050 257.550 ;
        RECT 704.100 257.100 705.900 257.850 ;
        RECT 710.100 257.100 711.900 257.850 ;
        RECT 686.100 254.100 687.900 254.850 ;
        RECT 685.950 250.950 688.050 253.050 ;
        RECT 671.400 237.600 673.200 243.600 ;
        RECT 678.000 237.600 679.800 249.600 ;
        RECT 689.400 243.600 690.600 255.900 ;
        RECT 692.100 254.100 693.900 254.850 ;
        RECT 703.950 253.950 706.050 256.050 ;
        RECT 709.950 253.800 712.050 256.050 ;
        RECT 691.950 250.950 694.050 253.050 ;
        RECT 713.700 249.600 714.600 258.900 ;
        RECT 718.950 258.450 721.050 259.050 ;
        RECT 727.950 258.450 730.050 259.050 ;
        RECT 718.950 257.550 730.050 258.450 ;
        RECT 718.950 256.950 721.050 257.550 ;
        RECT 727.950 256.950 730.050 257.550 ;
        RECT 733.950 258.450 736.050 259.050 ;
        RECT 745.950 258.450 748.050 259.050 ;
        RECT 733.950 257.550 748.050 258.450 ;
        RECT 733.950 256.950 736.050 257.550 ;
        RECT 745.950 256.950 748.050 257.550 ;
        RECT 763.950 256.950 766.050 259.050 ;
        RECT 767.100 255.900 768.300 260.100 ;
        RECT 775.950 261.450 780.000 262.050 ;
        RECT 781.950 261.450 784.050 262.050 ;
        RECT 775.950 260.550 784.050 261.450 ;
        RECT 775.950 259.950 780.000 260.550 ;
        RECT 781.950 259.950 784.050 260.550 ;
        RECT 787.950 259.950 790.050 262.050 ;
        RECT 794.550 259.950 795.900 262.050 ;
        RECT 796.950 259.950 799.050 262.050 ;
        RECT 800.100 260.250 800.850 262.050 ;
        RECT 807.150 261.600 825.000 262.800 ;
        RECT 807.150 261.000 808.950 261.600 ;
        RECT 818.100 261.000 819.900 261.600 ;
        RECT 808.050 260.100 808.950 261.000 ;
        RECT 824.100 260.850 825.000 261.600 ;
        RECT 725.100 254.100 726.900 254.850 ;
        RECT 724.950 250.950 727.050 253.050 ;
        RECT 704.400 248.700 712.200 249.600 ;
        RECT 689.400 237.600 691.200 243.600 ;
        RECT 704.400 237.600 706.200 248.700 ;
        RECT 710.400 237.600 712.200 248.700 ;
        RECT 713.400 237.600 715.200 249.600 ;
        RECT 728.400 243.600 729.600 255.900 ;
        RECT 731.100 254.100 732.900 254.850 ;
        RECT 743.100 254.100 744.900 254.850 ;
        RECT 730.950 250.950 733.050 253.050 ;
        RECT 742.950 250.950 745.050 253.050 ;
        RECT 746.400 243.600 747.600 255.900 ;
        RECT 764.100 255.150 765.900 255.900 ;
        RECT 749.100 254.100 750.900 254.850 ;
        RECT 748.950 250.950 751.050 253.050 ;
        RECT 766.950 250.650 768.300 255.900 ;
        RECT 769.950 253.950 772.050 256.050 ;
        RECT 770.100 252.150 771.900 252.900 ;
        RECT 765.600 249.600 768.300 250.650 ;
        RECT 782.400 249.600 783.300 258.900 ;
        RECT 788.100 258.150 789.900 258.900 ;
        RECT 785.100 257.100 786.900 257.850 ;
        RECT 791.100 257.100 792.900 257.850 ;
        RECT 784.950 253.800 787.050 256.050 ;
        RECT 790.950 253.950 793.050 256.050 ;
        RECT 794.550 249.600 795.750 259.950 ;
        RECT 824.100 259.050 825.900 260.850 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 821.100 256.800 822.900 257.400 ;
        RECT 796.950 251.400 798.750 253.200 ;
        RECT 797.850 250.200 802.050 251.400 ;
        RECT 808.050 250.200 808.950 255.900 ;
        RECT 814.950 253.950 817.050 256.050 ;
        RECT 818.100 255.600 822.900 256.800 ;
        RECT 816.750 251.700 818.550 252.000 ;
        RECT 826.950 251.700 827.850 266.400 ;
        RECT 816.750 251.100 827.850 251.700 ;
        RECT 728.400 237.600 730.200 243.600 ;
        RECT 746.400 237.600 748.200 243.600 ;
        RECT 765.600 237.600 767.400 249.600 ;
        RECT 781.800 237.600 783.600 249.600 ;
        RECT 784.800 248.700 792.600 249.600 ;
        RECT 784.800 237.600 786.600 248.700 ;
        RECT 790.800 237.600 792.600 248.700 ;
        RECT 794.550 237.600 796.350 249.600 ;
        RECT 799.950 249.300 802.050 250.200 ;
        RECT 802.950 249.300 808.950 250.200 ;
        RECT 810.150 250.500 827.850 251.100 ;
        RECT 810.150 250.200 818.550 250.500 ;
        RECT 802.950 248.400 803.850 249.300 ;
        RECT 801.150 246.600 803.850 248.400 ;
        RECT 804.750 248.100 806.550 248.400 ;
        RECT 810.150 248.100 811.050 250.200 ;
        RECT 826.950 249.600 827.850 250.500 ;
        RECT 804.750 247.200 811.050 248.100 ;
        RECT 811.950 248.700 813.750 249.300 ;
        RECT 811.950 247.500 819.450 248.700 ;
        RECT 804.750 246.600 806.550 247.200 ;
        RECT 818.250 246.600 819.450 247.500 ;
        RECT 799.950 243.600 803.850 245.700 ;
        RECT 808.950 245.550 810.750 246.300 ;
        RECT 813.750 245.550 815.550 246.300 ;
        RECT 808.950 244.500 815.550 245.550 ;
        RECT 818.250 244.500 823.050 246.600 ;
        RECT 802.050 237.600 803.850 243.600 ;
        RECT 809.850 237.600 811.650 244.500 ;
        RECT 818.250 243.600 819.450 244.500 ;
        RECT 817.650 237.600 819.450 243.600 ;
        RECT 826.050 237.600 827.850 249.600 ;
        RECT 16.800 221.400 20.100 233.400 ;
        RECT 36.600 221.400 38.400 233.400 ;
        RECT 55.800 227.400 57.600 233.400 ;
        RECT 13.950 214.950 16.050 217.050 ;
        RECT 14.700 213.150 16.500 213.900 ;
        RECT 11.250 212.100 13.050 212.850 ;
        RECT 17.400 212.100 18.600 221.400 ;
        RECT 36.600 220.350 39.300 221.400 ;
        RECT 19.950 214.950 22.050 217.050 ;
        RECT 35.100 215.100 36.900 215.850 ;
        RECT 37.950 215.100 39.300 220.350 ;
        RECT 41.100 218.100 42.900 218.850 ;
        RECT 52.950 217.950 55.050 220.050 ;
        RECT 20.100 213.150 21.900 213.900 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 10.950 208.950 13.050 211.050 ;
        RECT 16.950 208.950 19.050 211.050 ;
        RECT 22.950 208.950 25.050 211.050 ;
        RECT 38.100 210.900 39.300 215.100 ;
        RECT 40.950 214.950 43.050 217.050 ;
        RECT 53.100 216.150 54.900 216.900 ;
        RECT 56.400 215.100 57.600 227.400 ;
        RECT 69.600 221.400 71.400 233.400 ;
        RECT 84.600 221.400 86.400 233.400 ;
        RECT 100.800 221.400 102.600 233.400 ;
        RECT 103.800 222.300 105.600 233.400 ;
        RECT 109.800 222.300 111.600 233.400 ;
        RECT 103.800 221.400 111.600 222.300 ;
        RECT 121.500 221.400 123.300 233.400 ;
        RECT 127.800 227.400 129.600 233.400 ;
        RECT 69.600 220.350 72.300 221.400 ;
        RECT 84.600 220.350 87.300 221.400 ;
        RECT 58.950 217.950 61.050 220.050 ;
        RECT 59.100 216.150 60.900 216.900 ;
        RECT 68.100 215.100 69.900 215.850 ;
        RECT 70.950 215.100 72.300 220.350 ;
        RECT 74.100 218.100 75.900 218.850 ;
        RECT 52.950 211.950 58.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 71.100 210.900 72.300 215.100 ;
        RECT 73.950 214.950 76.050 217.050 ;
        RECT 83.100 215.100 84.900 215.850 ;
        RECT 85.950 215.100 87.300 220.350 ;
        RECT 89.100 218.100 90.900 218.850 ;
        RECT 82.950 211.800 85.050 214.050 ;
        RECT 86.100 210.900 87.300 215.100 ;
        RECT 88.950 214.950 91.050 217.050 ;
        RECT 101.400 212.100 102.300 221.400 ;
        RECT 103.950 214.950 106.050 217.050 ;
        RECT 109.950 214.950 112.050 217.050 ;
        RECT 104.100 213.150 105.900 213.900 ;
        RECT 110.100 213.150 111.900 213.900 ;
        RECT 107.100 212.100 108.900 212.850 ;
        RECT 121.800 212.100 123.000 221.400 ;
        RECT 128.400 220.500 129.600 227.400 ;
        RECT 123.900 219.600 129.600 220.500 ;
        RECT 138.600 221.400 140.400 233.400 ;
        RECT 153.600 221.400 155.400 233.400 ;
        RECT 171.600 221.400 173.400 233.400 ;
        RECT 187.500 221.400 189.300 233.400 ;
        RECT 208.800 227.400 210.600 233.400 ;
        RECT 138.600 220.350 141.300 221.400 ;
        RECT 123.900 218.700 125.850 219.600 ;
        RECT 124.950 212.100 125.850 218.700 ;
        RECT 128.100 215.100 129.900 215.850 ;
        RECT 137.100 215.100 138.900 215.850 ;
        RECT 139.950 215.100 141.300 220.350 ;
        RECT 152.700 220.350 155.400 221.400 ;
        RECT 170.700 220.350 173.400 221.400 ;
        RECT 143.100 218.100 144.900 218.850 ;
        RECT 149.100 218.100 150.900 218.850 ;
        RECT 37.950 209.100 39.300 210.900 ;
        RECT 17.400 207.300 18.600 207.900 ;
        RECT 14.400 206.100 18.600 207.300 ;
        RECT 22.950 207.150 24.750 207.900 ;
        RECT 37.950 207.450 40.050 208.050 ;
        RECT 49.950 207.450 52.050 208.050 ;
        RECT 37.950 206.550 52.050 207.450 ;
        RECT 56.400 206.700 57.600 210.900 ;
        RECT 70.950 209.100 72.300 210.900 ;
        RECT 85.950 209.100 87.300 210.900 ;
        RECT 100.950 208.950 103.050 211.050 ;
        RECT 106.950 208.950 109.050 211.050 ;
        RECT 121.950 208.950 124.050 211.050 ;
        RECT 14.400 204.600 15.300 206.100 ;
        RECT 37.950 205.950 40.050 206.550 ;
        RECT 49.950 205.950 52.050 206.550 ;
        RECT 54.000 205.800 57.600 206.700 ;
        RECT 70.950 207.450 73.050 208.050 ;
        RECT 79.950 207.450 82.050 208.050 ;
        RECT 70.950 206.550 82.050 207.450 ;
        RECT 70.950 205.950 73.050 206.550 ;
        RECT 79.950 205.950 82.050 206.550 ;
        RECT 85.950 207.450 88.050 208.050 ;
        RECT 94.950 207.450 97.050 208.050 ;
        RECT 125.100 207.900 125.850 212.100 ;
        RECT 127.950 211.950 130.050 214.050 ;
        RECT 133.950 211.950 139.050 214.050 ;
        RECT 140.100 210.900 141.300 215.100 ;
        RECT 142.950 211.950 145.050 217.050 ;
        RECT 148.950 214.950 151.050 217.050 ;
        RECT 152.700 215.100 154.050 220.350 ;
        RECT 167.100 218.100 168.900 218.850 ;
        RECT 155.100 215.100 156.900 215.850 ;
        RECT 139.950 209.100 141.300 210.900 ;
        RECT 152.700 210.900 153.900 215.100 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 166.950 211.950 169.050 217.050 ;
        RECT 170.700 215.100 172.050 220.350 ;
        RECT 187.950 218.100 189.150 221.400 ;
        RECT 173.100 215.100 174.900 215.850 ;
        RECT 170.700 210.900 171.900 215.100 ;
        RECT 184.950 214.950 187.050 217.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 188.100 213.900 189.150 218.100 ;
        RECT 205.950 217.950 208.050 220.050 ;
        RECT 190.950 214.950 193.050 217.050 ;
        RECT 206.100 216.150 207.900 216.900 ;
        RECT 209.400 215.100 210.600 227.400 ;
        RECT 220.800 221.400 222.600 233.400 ;
        RECT 223.800 222.300 225.600 233.400 ;
        RECT 229.800 222.300 231.600 233.400 ;
        RECT 223.800 221.400 231.600 222.300 ;
        RECT 239.400 227.400 241.200 233.400 ;
        RECT 211.950 217.950 214.050 220.050 ;
        RECT 212.100 216.150 213.900 216.900 ;
        RECT 185.100 213.150 186.900 213.900 ;
        RECT 182.100 212.100 183.900 212.850 ;
        RECT 187.950 212.100 189.150 213.900 ;
        RECT 191.100 213.150 192.900 213.900 ;
        RECT 196.950 213.450 199.050 214.050 ;
        RECT 208.950 213.450 211.050 214.050 ;
        RECT 196.950 212.550 211.050 213.450 ;
        RECT 196.950 211.950 199.050 212.550 ;
        RECT 208.950 211.950 211.050 212.550 ;
        RECT 221.400 212.100 222.300 221.400 ;
        RECT 223.950 214.950 226.050 217.050 ;
        RECT 229.950 214.950 232.050 217.050 ;
        RECT 236.100 215.100 237.900 215.850 ;
        RECT 224.100 213.150 225.900 213.900 ;
        RECT 230.100 213.150 231.900 213.900 ;
        RECT 227.100 212.100 228.900 212.850 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 152.700 209.100 154.050 210.900 ;
        RECT 170.700 209.100 172.050 210.900 ;
        RECT 181.950 208.950 184.050 211.050 ;
        RECT 187.950 210.450 190.050 211.050 ;
        RECT 202.950 210.450 205.050 211.050 ;
        RECT 187.950 209.550 205.050 210.450 ;
        RECT 187.950 208.950 190.050 209.550 ;
        RECT 202.950 208.950 205.050 209.550 ;
        RECT 85.950 206.550 97.050 207.450 ;
        RECT 85.950 205.950 88.050 206.550 ;
        RECT 94.950 205.950 97.050 206.550 ;
        RECT 10.800 199.500 12.600 204.600 ;
        RECT 13.800 200.400 15.600 204.600 ;
        RECT 16.800 204.000 24.600 204.900 ;
        RECT 16.800 199.500 18.600 204.000 ;
        RECT 10.800 198.600 18.600 199.500 ;
        RECT 22.800 198.600 24.600 204.000 ;
        RECT 38.400 201.600 39.600 204.900 ;
        RECT 37.800 198.600 39.600 201.600 ;
        RECT 54.000 198.600 55.800 205.800 ;
        RECT 71.400 201.600 72.600 204.900 ;
        RECT 86.400 201.600 87.600 204.900 ;
        RECT 101.400 204.600 102.300 207.900 ;
        RECT 121.800 204.600 123.000 207.900 ;
        RECT 124.950 207.300 125.850 207.900 ;
        RECT 123.900 206.400 125.850 207.300 ;
        RECT 123.900 205.500 129.000 206.400 ;
        RECT 136.950 205.950 142.050 208.050 ;
        RECT 151.950 207.450 154.050 208.050 ;
        RECT 163.950 207.450 166.050 208.050 ;
        RECT 151.950 206.550 166.050 207.450 ;
        RECT 151.950 205.950 154.050 206.550 ;
        RECT 163.950 205.950 166.050 206.550 ;
        RECT 169.950 205.950 172.050 208.050 ;
        RECT 188.850 207.750 190.050 207.900 ;
        RECT 188.850 206.700 192.600 207.750 ;
        RECT 209.400 206.700 210.600 210.900 ;
        RECT 220.950 208.950 223.050 211.050 ;
        RECT 226.950 208.950 229.050 211.050 ;
        RECT 101.400 202.950 106.800 204.600 ;
        RECT 70.800 198.600 72.600 201.600 ;
        RECT 85.800 198.600 87.600 201.600 ;
        RECT 105.000 198.600 106.800 202.950 ;
        RECT 121.500 198.600 123.300 204.600 ;
        RECT 127.800 201.600 129.000 205.500 ;
        RECT 140.400 201.600 141.600 204.900 ;
        RECT 127.800 198.600 129.600 201.600 ;
        RECT 139.800 198.600 141.600 201.600 ;
        RECT 152.400 201.600 153.600 204.900 ;
        RECT 170.400 201.600 171.600 204.900 ;
        RECT 182.400 203.700 190.200 205.050 ;
        RECT 152.400 198.600 154.200 201.600 ;
        RECT 170.400 198.600 172.200 201.600 ;
        RECT 182.400 198.600 184.200 203.700 ;
        RECT 188.400 198.600 190.200 203.700 ;
        RECT 191.400 204.600 192.600 206.700 ;
        RECT 207.000 205.800 210.600 206.700 ;
        RECT 191.400 198.600 193.200 204.600 ;
        RECT 207.000 198.600 208.800 205.800 ;
        RECT 221.400 204.600 222.300 207.900 ;
        RECT 239.400 207.300 240.450 227.400 ;
        RECT 246.000 221.400 247.800 233.400 ;
        RECT 260.400 227.400 262.200 233.400 ;
        RECT 260.700 227.100 262.200 227.400 ;
        RECT 266.400 227.400 268.200 233.400 ;
        RECT 266.400 227.100 267.300 227.400 ;
        RECT 260.700 226.200 267.300 227.100 ;
        RECT 241.950 214.950 244.050 217.050 ;
        RECT 242.100 213.150 243.900 213.900 ;
        RECT 246.000 212.100 247.050 221.400 ;
        RECT 256.950 220.950 259.050 223.050 ;
        RECT 266.400 221.100 267.300 226.200 ;
        RECT 278.400 222.300 280.200 233.400 ;
        RECT 284.400 222.300 286.200 233.400 ;
        RECT 278.400 221.400 286.200 222.300 ;
        RECT 287.400 221.400 289.200 233.400 ;
        RECT 299.400 227.400 301.200 233.400 ;
        RECT 257.100 219.150 258.900 219.900 ;
        RECT 265.950 219.450 268.050 220.050 ;
        RECT 270.000 219.450 274.050 220.050 ;
        RECT 260.100 218.100 261.900 218.850 ;
        RECT 265.950 218.550 274.050 219.450 ;
        RECT 265.950 217.950 268.050 218.550 ;
        RECT 270.000 217.950 274.050 218.550 ;
        RECT 259.950 214.950 262.050 217.050 ;
        RECT 262.950 211.950 265.050 214.050 ;
        RECT 244.950 210.450 247.050 211.050 ;
        RECT 256.950 210.450 259.050 211.050 ;
        RECT 244.950 209.550 259.050 210.450 ;
        RECT 263.100 210.150 264.900 210.900 ;
        RECT 244.950 208.950 247.050 209.550 ;
        RECT 256.950 208.950 259.050 209.550 ;
        RECT 266.400 208.650 267.300 216.900 ;
        RECT 277.950 214.950 280.050 217.050 ;
        RECT 283.950 214.950 286.050 217.200 ;
        RECT 278.100 213.150 279.900 213.900 ;
        RECT 284.100 213.150 285.900 213.900 ;
        RECT 281.100 212.100 282.900 212.850 ;
        RECT 287.700 212.100 288.600 221.400 ;
        RECT 296.100 215.100 297.900 215.850 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 280.950 208.950 283.050 211.050 ;
        RECT 286.950 210.900 291.450 211.050 ;
        RECT 286.950 208.950 292.050 210.900 ;
        RECT 289.950 208.800 292.050 208.950 ;
        RECT 236.400 206.400 243.900 207.300 ;
        RECT 221.400 202.950 226.800 204.600 ;
        RECT 225.000 198.600 226.800 202.950 ;
        RECT 236.400 198.600 238.200 206.400 ;
        RECT 242.100 205.500 243.900 206.400 ;
        RECT 244.950 204.600 245.850 207.900 ;
        RECT 243.900 202.800 245.850 204.600 ;
        RECT 263.100 207.000 267.300 208.650 ;
        RECT 243.900 198.600 245.700 202.800 ;
        RECT 263.100 198.600 264.900 207.000 ;
        RECT 287.700 204.600 288.600 207.900 ;
        RECT 299.400 207.300 300.450 227.400 ;
        RECT 306.000 221.400 307.800 233.400 ;
        RECT 312.150 221.400 313.950 233.400 ;
        RECT 320.550 227.400 322.350 233.400 ;
        RECT 320.550 226.500 321.750 227.400 ;
        RECT 328.350 226.500 330.150 233.400 ;
        RECT 336.150 227.400 337.950 233.400 ;
        RECT 316.950 224.400 321.750 226.500 ;
        RECT 324.450 225.450 331.050 226.500 ;
        RECT 324.450 224.700 326.250 225.450 ;
        RECT 329.250 224.700 331.050 225.450 ;
        RECT 336.150 225.300 340.050 227.400 ;
        RECT 320.550 223.500 321.750 224.400 ;
        RECT 333.450 223.800 335.250 224.400 ;
        RECT 320.550 222.300 328.050 223.500 ;
        RECT 326.250 221.700 328.050 222.300 ;
        RECT 328.950 222.900 335.250 223.800 ;
        RECT 301.950 214.950 304.050 217.050 ;
        RECT 302.100 213.150 303.900 213.900 ;
        RECT 306.000 212.100 307.050 221.400 ;
        RECT 312.150 220.500 313.050 221.400 ;
        RECT 328.950 220.800 329.850 222.900 ;
        RECT 333.450 222.600 335.250 222.900 ;
        RECT 336.150 222.600 338.850 224.400 ;
        RECT 336.150 221.700 337.050 222.600 ;
        RECT 321.450 220.500 329.850 220.800 ;
        RECT 312.150 219.900 329.850 220.500 ;
        RECT 331.050 220.800 337.050 221.700 ;
        RECT 337.950 220.800 340.050 221.700 ;
        RECT 343.650 221.400 345.450 233.400 ;
        RECT 358.800 227.400 360.600 233.400 ;
        RECT 312.150 219.300 323.250 219.900 ;
        RECT 304.950 208.950 310.050 211.050 ;
        RECT 283.200 202.950 288.600 204.600 ;
        RECT 296.400 206.400 303.900 207.300 ;
        RECT 283.200 198.600 285.000 202.950 ;
        RECT 296.400 198.600 298.200 206.400 ;
        RECT 302.100 205.500 303.900 206.400 ;
        RECT 304.950 204.600 305.850 207.900 ;
        RECT 303.900 202.800 305.850 204.600 ;
        RECT 312.150 204.600 313.050 219.300 ;
        RECT 321.450 219.000 323.250 219.300 ;
        RECT 317.100 214.200 321.900 215.400 ;
        RECT 322.950 214.950 325.050 217.050 ;
        RECT 331.050 215.100 331.950 220.800 ;
        RECT 337.950 219.600 342.150 220.800 ;
        RECT 341.250 217.800 343.050 219.600 ;
        RECT 317.100 213.600 318.900 214.200 ;
        RECT 328.950 211.950 331.050 214.050 ;
        RECT 314.100 210.150 315.900 211.950 ;
        RECT 344.250 211.050 345.450 221.400 ;
        RECT 355.950 217.800 358.050 220.050 ;
        RECT 356.100 216.150 357.900 216.900 ;
        RECT 359.400 215.100 360.600 227.400 ;
        RECT 373.500 221.400 375.300 233.400 ;
        RECT 395.700 221.400 397.500 233.400 ;
        RECT 412.800 221.400 414.600 233.400 ;
        RECT 361.950 217.950 364.050 220.050 ;
        RECT 373.950 218.100 375.150 221.400 ;
        RECT 362.100 216.150 363.900 216.900 ;
        RECT 370.950 214.950 373.050 217.050 ;
        RECT 352.950 213.450 357.000 214.050 ;
        RECT 358.950 213.450 361.050 214.050 ;
        RECT 374.100 213.900 375.150 218.100 ;
        RECT 395.850 218.100 397.050 221.400 ;
        RECT 376.950 214.950 379.050 217.050 ;
        RECT 385.950 216.450 390.000 217.050 ;
        RECT 391.950 216.450 394.050 217.050 ;
        RECT 385.950 215.550 394.050 216.450 ;
        RECT 385.950 214.950 390.000 215.550 ;
        RECT 391.950 214.950 394.050 215.550 ;
        RECT 395.850 213.900 396.900 218.100 ;
        RECT 397.950 214.950 400.050 217.050 ;
        RECT 352.950 212.550 361.050 213.450 ;
        RECT 371.100 213.150 372.900 213.900 ;
        RECT 352.950 211.950 357.000 212.550 ;
        RECT 358.950 211.950 361.050 212.550 ;
        RECT 368.100 212.100 369.900 212.850 ;
        RECT 373.950 212.100 375.150 213.900 ;
        RECT 377.100 213.150 378.900 213.900 ;
        RECT 392.100 213.150 393.900 213.900 ;
        RECT 395.850 212.100 397.050 213.900 ;
        RECT 398.100 213.150 399.900 213.900 ;
        RECT 401.100 212.100 402.900 212.850 ;
        RECT 413.400 212.100 414.600 221.400 ;
        RECT 422.400 227.400 424.200 233.400 ;
        RECT 422.400 220.500 423.600 227.400 ;
        RECT 428.700 221.400 430.500 233.400 ;
        RECT 435.150 221.400 436.950 233.400 ;
        RECT 443.550 227.400 445.350 233.400 ;
        RECT 443.550 226.500 444.750 227.400 ;
        RECT 451.350 226.500 453.150 233.400 ;
        RECT 459.150 227.400 460.950 233.400 ;
        RECT 439.950 224.400 444.750 226.500 ;
        RECT 447.450 225.450 454.050 226.500 ;
        RECT 447.450 224.700 449.250 225.450 ;
        RECT 452.250 224.700 454.050 225.450 ;
        RECT 459.150 225.300 463.050 227.400 ;
        RECT 443.550 223.500 444.750 224.400 ;
        RECT 456.450 223.800 458.250 224.400 ;
        RECT 443.550 222.300 451.050 223.500 ;
        RECT 449.250 221.700 451.050 222.300 ;
        RECT 451.950 222.900 458.250 223.800 ;
        RECT 422.400 219.600 428.100 220.500 ;
        RECT 426.150 218.700 428.100 219.600 ;
        RECT 415.950 214.950 418.050 217.050 ;
        RECT 422.100 215.100 423.900 215.850 ;
        RECT 416.100 213.150 417.900 213.900 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 426.150 212.100 427.050 218.700 ;
        RECT 429.000 212.100 430.200 221.400 ;
        RECT 435.150 220.500 436.050 221.400 ;
        RECT 451.950 220.800 452.850 222.900 ;
        RECT 456.450 222.600 458.250 222.900 ;
        RECT 459.150 222.600 461.850 224.400 ;
        RECT 459.150 221.700 460.050 222.600 ;
        RECT 444.450 220.500 452.850 220.800 ;
        RECT 435.150 219.900 452.850 220.500 ;
        RECT 454.050 220.800 460.050 221.700 ;
        RECT 460.950 220.800 463.050 221.700 ;
        RECT 466.650 221.400 468.450 233.400 ;
        RECT 478.800 227.400 480.600 233.400 ;
        RECT 435.150 219.300 446.250 219.900 ;
        RECT 315.000 209.400 315.900 210.150 ;
        RECT 331.050 210.000 331.950 210.900 ;
        RECT 320.100 209.400 321.900 210.000 ;
        RECT 331.050 209.400 332.850 210.000 ;
        RECT 315.000 208.200 332.850 209.400 ;
        RECT 339.150 208.950 339.900 210.750 ;
        RECT 340.950 208.950 343.050 211.050 ;
        RECT 344.100 208.950 345.450 211.050 ;
        RECT 320.850 205.200 321.900 208.200 ;
        RECT 303.900 198.600 305.700 202.800 ;
        RECT 312.150 198.600 313.950 204.600 ;
        RECT 316.950 202.500 319.050 204.600 ;
        RECT 320.550 203.400 322.350 205.200 ;
        RECT 323.850 204.450 325.650 205.200 ;
        RECT 344.250 204.600 345.450 208.950 ;
        RECT 359.400 206.700 360.600 210.900 ;
        RECT 367.950 208.950 370.050 211.050 ;
        RECT 373.950 208.950 376.050 211.050 ;
        RECT 379.950 210.450 382.050 211.050 ;
        RECT 394.950 210.450 397.050 211.050 ;
        RECT 379.950 209.550 397.050 210.450 ;
        RECT 379.950 208.950 382.050 209.550 ;
        RECT 394.950 208.950 397.050 209.550 ;
        RECT 400.950 208.950 403.050 211.050 ;
        RECT 412.950 208.950 415.050 211.050 ;
        RECT 426.150 207.900 426.900 212.100 ;
        RECT 427.950 208.950 430.050 211.050 ;
        RECT 374.850 207.750 376.050 207.900 ;
        RECT 394.950 207.750 396.150 207.900 ;
        RECT 374.850 206.700 378.600 207.750 ;
        RECT 323.850 203.400 328.800 204.450 ;
        RECT 337.950 203.700 340.050 204.600 ;
        RECT 318.000 201.600 319.050 202.500 ;
        RECT 327.750 201.600 328.800 203.400 ;
        RECT 336.300 202.500 340.050 203.700 ;
        RECT 336.300 201.600 337.350 202.500 ;
        RECT 318.000 200.700 321.750 201.600 ;
        RECT 319.950 198.600 321.750 200.700 ;
        RECT 327.750 198.600 329.550 201.600 ;
        RECT 335.550 198.600 337.350 201.600 ;
        RECT 343.650 198.600 345.450 204.600 ;
        RECT 357.000 205.800 360.600 206.700 ;
        RECT 357.000 198.600 358.800 205.800 ;
        RECT 368.400 203.700 376.200 205.050 ;
        RECT 368.400 198.600 370.200 203.700 ;
        RECT 374.400 198.600 376.200 203.700 ;
        RECT 377.400 204.600 378.600 206.700 ;
        RECT 392.400 206.700 396.150 207.750 ;
        RECT 392.400 204.600 393.600 206.700 ;
        RECT 377.400 198.600 379.200 204.600 ;
        RECT 391.800 198.600 393.600 204.600 ;
        RECT 394.800 203.700 402.600 205.050 ;
        RECT 413.400 204.600 414.600 207.900 ;
        RECT 426.150 207.300 427.050 207.900 ;
        RECT 426.150 206.400 428.100 207.300 ;
        RECT 394.800 198.600 396.600 203.700 ;
        RECT 400.800 198.600 402.600 203.700 ;
        RECT 412.800 198.600 414.600 204.600 ;
        RECT 423.000 205.500 428.100 206.400 ;
        RECT 423.000 201.600 424.200 205.500 ;
        RECT 429.000 204.600 430.200 207.900 ;
        RECT 435.150 204.600 436.050 219.300 ;
        RECT 444.450 219.000 446.250 219.300 ;
        RECT 440.100 214.200 444.900 215.400 ;
        RECT 445.950 214.950 451.050 217.050 ;
        RECT 454.050 215.100 454.950 220.800 ;
        RECT 460.950 219.600 465.150 220.800 ;
        RECT 464.250 217.800 466.050 219.600 ;
        RECT 440.100 213.600 441.900 214.200 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 437.100 210.150 438.900 211.950 ;
        RECT 467.250 211.050 468.450 221.400 ;
        RECT 479.400 218.100 480.600 227.400 ;
        RECT 491.400 227.400 493.200 233.400 ;
        RECT 487.950 217.950 490.050 220.050 ;
        RECT 478.950 214.950 484.050 217.050 ;
        RECT 488.100 216.150 489.900 216.900 ;
        RECT 491.400 215.100 492.600 227.400 ;
        RECT 510.600 221.400 512.400 233.400 ;
        RECT 527.700 221.400 529.500 233.400 ;
        RECT 544.800 227.400 546.600 233.400 ;
        RECT 509.700 220.350 512.400 221.400 ;
        RECT 493.950 217.950 496.050 220.050 ;
        RECT 506.100 218.100 507.900 218.850 ;
        RECT 494.100 216.150 495.900 216.900 ;
        RECT 499.950 216.450 504.000 217.050 ;
        RECT 505.950 216.450 508.050 217.050 ;
        RECT 499.950 215.550 508.050 216.450 ;
        RECT 499.950 214.950 504.000 215.550 ;
        RECT 505.950 214.950 508.050 215.550 ;
        RECT 509.700 215.100 511.050 220.350 ;
        RECT 527.850 218.100 529.050 221.400 ;
        RECT 545.400 218.100 546.600 227.400 ;
        RECT 561.600 221.400 563.400 233.400 ;
        RECT 560.700 220.350 563.400 221.400 ;
        RECT 578.400 227.400 580.200 233.400 ;
        RECT 557.100 218.100 558.900 218.850 ;
        RECT 512.100 215.100 513.900 215.850 ;
        RECT 438.000 209.400 438.900 210.150 ;
        RECT 454.050 210.000 454.950 210.900 ;
        RECT 443.100 209.400 444.900 210.000 ;
        RECT 454.050 209.400 455.850 210.000 ;
        RECT 438.000 208.200 455.850 209.400 ;
        RECT 462.150 208.950 462.900 210.750 ;
        RECT 463.950 208.950 466.050 211.050 ;
        RECT 467.100 208.950 468.450 211.050 ;
        RECT 443.850 205.200 444.900 208.200 ;
        RECT 422.400 198.600 424.200 201.600 ;
        RECT 428.700 198.600 430.500 204.600 ;
        RECT 435.150 198.600 436.950 204.600 ;
        RECT 439.950 202.500 442.050 204.600 ;
        RECT 443.550 203.400 445.350 205.200 ;
        RECT 446.850 204.450 448.650 205.200 ;
        RECT 467.250 204.600 468.450 208.950 ;
        RECT 446.850 203.400 451.800 204.450 ;
        RECT 460.950 203.700 463.050 204.600 ;
        RECT 441.000 201.600 442.050 202.500 ;
        RECT 450.750 201.600 451.800 203.400 ;
        RECT 459.300 202.500 463.050 203.700 ;
        RECT 459.300 201.600 460.350 202.500 ;
        RECT 441.000 200.700 444.750 201.600 ;
        RECT 442.950 198.600 444.750 200.700 ;
        RECT 450.750 198.600 452.550 201.600 ;
        RECT 458.550 198.600 460.350 201.600 ;
        RECT 466.650 198.600 468.450 204.600 ;
        RECT 479.400 201.600 480.600 213.900 ;
        RECT 482.100 212.100 483.900 212.850 ;
        RECT 487.950 211.950 493.050 214.050 ;
        RECT 481.950 208.950 484.050 211.050 ;
        RECT 509.700 210.900 510.900 215.100 ;
        RECT 523.950 214.950 526.050 217.050 ;
        RECT 511.950 211.950 514.050 214.050 ;
        RECT 527.850 213.900 528.900 218.100 ;
        RECT 529.950 214.950 532.050 217.050 ;
        RECT 535.950 216.450 538.050 217.050 ;
        RECT 544.950 216.450 547.050 217.050 ;
        RECT 535.950 215.550 547.050 216.450 ;
        RECT 535.950 214.950 538.050 215.550 ;
        RECT 544.950 214.950 547.050 215.550 ;
        RECT 556.950 214.950 559.050 217.050 ;
        RECT 560.700 215.100 562.050 220.350 ;
        RECT 578.400 218.100 579.600 227.400 ;
        RECT 593.400 220.500 595.200 233.400 ;
        RECT 599.400 220.500 601.200 233.400 ;
        RECT 605.400 220.500 607.200 233.400 ;
        RECT 611.400 220.500 613.200 233.400 ;
        RECT 621.150 221.400 622.950 233.400 ;
        RECT 629.550 227.400 631.350 233.400 ;
        RECT 629.550 226.500 630.750 227.400 ;
        RECT 637.350 226.500 639.150 233.400 ;
        RECT 645.150 227.400 646.950 233.400 ;
        RECT 625.950 224.400 630.750 226.500 ;
        RECT 633.450 225.450 640.050 226.500 ;
        RECT 633.450 224.700 635.250 225.450 ;
        RECT 638.250 224.700 640.050 225.450 ;
        RECT 645.150 225.300 649.050 227.400 ;
        RECT 629.550 223.500 630.750 224.400 ;
        RECT 642.450 223.800 644.250 224.400 ;
        RECT 629.550 222.300 637.050 223.500 ;
        RECT 635.250 221.700 637.050 222.300 ;
        RECT 637.950 222.900 644.250 223.800 ;
        RECT 621.150 220.500 622.050 221.400 ;
        RECT 637.950 220.800 638.850 222.900 ;
        RECT 642.450 222.600 644.250 222.900 ;
        RECT 645.150 222.600 647.850 224.400 ;
        RECT 645.150 221.700 646.050 222.600 ;
        RECT 630.450 220.500 638.850 220.800 ;
        RECT 593.400 219.300 597.300 220.500 ;
        RECT 599.400 219.300 603.300 220.500 ;
        RECT 605.400 219.300 609.300 220.500 ;
        RECT 611.400 219.300 614.100 220.500 ;
        RECT 571.950 216.450 576.000 217.050 ;
        RECT 577.950 216.450 580.050 217.050 ;
        RECT 563.100 215.100 564.900 215.850 ;
        RECT 571.950 215.550 580.050 216.450 ;
        RECT 524.100 213.150 525.900 213.900 ;
        RECT 527.850 212.100 529.050 213.900 ;
        RECT 530.100 213.150 531.900 213.900 ;
        RECT 533.100 212.100 534.900 212.850 ;
        RECT 491.400 206.700 492.600 210.900 ;
        RECT 509.700 209.100 511.050 210.900 ;
        RECT 526.950 208.950 529.050 211.050 ;
        RECT 532.950 208.950 535.050 211.050 ;
        RECT 508.950 207.450 511.050 208.050 ;
        RECT 517.950 207.450 520.050 208.050 ;
        RECT 526.950 207.750 528.150 207.900 ;
        RECT 491.400 205.800 495.000 206.700 ;
        RECT 508.950 206.550 520.050 207.450 ;
        RECT 508.950 205.950 511.050 206.550 ;
        RECT 517.950 205.950 520.050 206.550 ;
        RECT 524.400 206.700 528.150 207.750 ;
        RECT 478.800 198.600 480.600 201.600 ;
        RECT 493.200 198.600 495.000 205.800 ;
        RECT 509.400 201.600 510.600 204.900 ;
        RECT 524.400 204.600 525.600 206.700 ;
        RECT 509.400 198.600 511.200 201.600 ;
        RECT 523.800 198.600 525.600 204.600 ;
        RECT 526.800 203.700 534.600 205.050 ;
        RECT 526.800 198.600 528.600 203.700 ;
        RECT 532.800 198.600 534.600 203.700 ;
        RECT 545.400 201.600 546.600 213.900 ;
        RECT 548.100 212.100 549.900 212.850 ;
        RECT 547.950 208.950 550.050 211.050 ;
        RECT 560.700 210.900 561.900 215.100 ;
        RECT 571.950 214.950 576.000 215.550 ;
        RECT 577.950 214.950 580.050 215.550 ;
        RECT 562.950 211.950 565.050 214.050 ;
        RECT 575.100 212.100 576.900 212.850 ;
        RECT 560.700 209.100 562.050 210.900 ;
        RECT 574.950 208.950 577.050 211.050 ;
        RECT 553.950 207.450 558.000 208.050 ;
        RECT 559.950 207.450 562.050 208.050 ;
        RECT 553.950 206.550 562.050 207.450 ;
        RECT 553.950 205.950 558.000 206.550 ;
        RECT 559.950 205.950 562.050 206.550 ;
        RECT 544.800 198.600 546.600 201.600 ;
        RECT 560.400 201.600 561.600 204.900 ;
        RECT 578.400 201.600 579.600 213.900 ;
        RECT 593.100 210.150 594.900 210.900 ;
        RECT 596.100 208.800 597.300 219.300 ;
        RECT 598.500 208.800 600.300 209.400 ;
        RECT 596.100 207.600 600.300 208.800 ;
        RECT 602.100 208.800 603.300 219.300 ;
        RECT 604.500 208.800 606.300 209.400 ;
        RECT 602.100 207.600 606.300 208.800 ;
        RECT 608.100 208.800 609.300 219.300 ;
        RECT 613.200 215.100 614.100 219.300 ;
        RECT 621.150 219.900 638.850 220.500 ;
        RECT 640.050 220.800 646.050 221.700 ;
        RECT 646.950 220.800 649.050 221.700 ;
        RECT 652.650 221.400 654.450 233.400 ;
        RECT 664.500 221.400 666.300 233.400 ;
        RECT 684.600 221.400 686.400 233.400 ;
        RECT 699.600 221.400 701.400 233.400 ;
        RECT 710.400 221.400 712.200 233.400 ;
        RECT 717.900 222.900 719.700 233.400 ;
        RECT 733.800 227.400 735.600 233.400 ;
        RECT 717.900 221.400 720.300 222.900 ;
        RECT 621.150 219.300 632.250 219.900 ;
        RECT 613.950 211.950 619.050 214.050 ;
        RECT 610.500 208.800 612.300 209.400 ;
        RECT 608.100 207.600 612.300 208.800 ;
        RECT 596.100 206.700 597.300 207.600 ;
        RECT 602.100 206.700 603.300 207.600 ;
        RECT 608.100 206.700 609.300 207.600 ;
        RECT 613.200 206.700 614.100 210.900 ;
        RECT 593.400 205.500 597.300 206.700 ;
        RECT 599.400 205.500 603.300 206.700 ;
        RECT 605.400 205.500 609.300 206.700 ;
        RECT 611.400 205.500 614.100 206.700 ;
        RECT 560.400 198.600 562.200 201.600 ;
        RECT 578.400 198.600 580.200 201.600 ;
        RECT 593.400 198.600 595.200 205.500 ;
        RECT 599.400 198.600 601.200 205.500 ;
        RECT 605.400 198.600 607.200 205.500 ;
        RECT 611.400 198.600 613.200 205.500 ;
        RECT 621.150 204.600 622.050 219.300 ;
        RECT 630.450 219.000 632.250 219.300 ;
        RECT 626.100 214.200 630.900 215.400 ;
        RECT 631.950 214.950 634.050 217.050 ;
        RECT 640.050 215.100 640.950 220.800 ;
        RECT 646.950 219.600 651.150 220.800 ;
        RECT 650.250 217.800 652.050 219.600 ;
        RECT 626.100 213.600 627.900 214.200 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 623.100 210.150 624.900 211.950 ;
        RECT 653.250 211.050 654.450 221.400 ;
        RECT 664.950 218.100 666.150 221.400 ;
        RECT 684.600 220.350 687.300 221.400 ;
        RECT 699.600 220.350 702.300 221.400 ;
        RECT 661.950 214.950 664.050 217.050 ;
        RECT 665.100 213.900 666.150 218.100 ;
        RECT 667.950 214.950 670.050 217.050 ;
        RECT 683.100 215.100 684.900 215.850 ;
        RECT 685.950 215.100 687.300 220.350 ;
        RECT 689.100 218.100 690.900 218.850 ;
        RECT 662.100 213.150 663.900 213.900 ;
        RECT 659.100 212.100 660.900 212.850 ;
        RECT 664.950 212.100 666.150 213.900 ;
        RECT 668.100 213.150 669.900 213.900 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 624.000 209.400 624.900 210.150 ;
        RECT 640.050 210.000 640.950 210.900 ;
        RECT 629.100 209.400 630.900 210.000 ;
        RECT 640.050 209.400 641.850 210.000 ;
        RECT 624.000 208.200 641.850 209.400 ;
        RECT 648.150 208.950 648.900 210.750 ;
        RECT 629.850 205.200 630.900 208.200 ;
        RECT 649.950 205.950 652.050 211.050 ;
        RECT 653.100 208.950 654.450 211.050 ;
        RECT 655.950 208.950 661.050 211.050 ;
        RECT 664.950 208.950 667.050 211.050 ;
        RECT 686.100 210.900 687.300 215.100 ;
        RECT 688.950 214.950 691.050 217.050 ;
        RECT 698.100 215.100 699.900 215.850 ;
        RECT 700.950 215.100 702.300 220.350 ;
        RECT 710.400 220.200 711.600 221.400 ;
        RECT 710.400 219.000 717.600 220.200 ;
        RECT 704.100 218.100 705.900 218.850 ;
        RECT 715.800 218.400 717.600 219.000 ;
        RECT 697.950 211.950 700.050 214.050 ;
        RECT 701.100 210.900 702.300 215.100 ;
        RECT 703.950 214.950 706.050 217.050 ;
        RECT 709.950 214.950 712.050 217.050 ;
        RECT 710.100 213.150 711.900 213.900 ;
        RECT 713.100 212.100 714.900 212.850 ;
        RECT 685.950 209.100 687.300 210.900 ;
        RECT 700.950 209.100 702.300 210.900 ;
        RECT 712.950 208.950 715.050 211.050 ;
        RECT 621.150 198.600 622.950 204.600 ;
        RECT 625.950 202.500 628.050 204.600 ;
        RECT 629.550 203.400 631.350 205.200 ;
        RECT 632.850 204.450 634.650 205.200 ;
        RECT 653.250 204.600 654.450 208.950 ;
        RECT 665.850 207.750 667.050 207.900 ;
        RECT 665.850 206.700 669.600 207.750 ;
        RECT 632.850 203.400 637.800 204.450 ;
        RECT 646.950 203.700 649.050 204.600 ;
        RECT 627.000 201.600 628.050 202.500 ;
        RECT 636.750 201.600 637.800 203.400 ;
        RECT 645.300 202.500 649.050 203.700 ;
        RECT 645.300 201.600 646.350 202.500 ;
        RECT 627.000 200.700 630.750 201.600 ;
        RECT 628.950 198.600 630.750 200.700 ;
        RECT 636.750 198.600 638.550 201.600 ;
        RECT 644.550 198.600 646.350 201.600 ;
        RECT 652.650 198.600 654.450 204.600 ;
        RECT 659.400 203.700 667.200 205.050 ;
        RECT 659.400 198.600 661.200 203.700 ;
        RECT 665.400 198.600 667.200 203.700 ;
        RECT 668.400 204.600 669.600 206.700 ;
        RECT 685.950 207.450 688.050 208.050 ;
        RECT 694.800 207.450 696.900 208.050 ;
        RECT 685.950 206.550 696.900 207.450 ;
        RECT 685.950 205.950 688.050 206.550 ;
        RECT 694.800 205.950 696.900 206.550 ;
        RECT 697.950 205.950 703.050 208.050 ;
        RECT 716.700 207.600 717.600 218.400 ;
        RECT 718.950 215.100 720.300 221.400 ;
        RECT 730.950 217.950 733.050 220.050 ;
        RECT 731.100 216.150 732.900 216.900 ;
        RECT 734.400 215.100 735.600 227.400 ;
        RECT 740.550 221.400 742.350 233.400 ;
        RECT 748.050 227.400 749.850 233.400 ;
        RECT 745.950 225.300 749.850 227.400 ;
        RECT 755.850 226.500 757.650 233.400 ;
        RECT 763.650 227.400 765.450 233.400 ;
        RECT 764.250 226.500 765.450 227.400 ;
        RECT 754.950 225.450 761.550 226.500 ;
        RECT 754.950 224.700 756.750 225.450 ;
        RECT 759.750 224.700 761.550 225.450 ;
        RECT 764.250 224.400 769.050 226.500 ;
        RECT 747.150 222.600 749.850 224.400 ;
        RECT 750.750 223.800 752.550 224.400 ;
        RECT 750.750 222.900 757.050 223.800 ;
        RECT 764.250 223.500 765.450 224.400 ;
        RECT 750.750 222.600 752.550 222.900 ;
        RECT 748.950 221.700 749.850 222.600 ;
        RECT 736.950 217.950 739.050 220.050 ;
        RECT 737.100 216.150 738.900 216.900 ;
        RECT 718.950 211.950 724.050 214.050 ;
        RECT 733.950 211.950 736.050 214.050 ;
        RECT 740.550 211.050 741.750 221.400 ;
        RECT 745.950 220.800 748.050 221.700 ;
        RECT 748.950 220.800 754.950 221.700 ;
        RECT 743.850 219.600 748.050 220.800 ;
        RECT 742.950 217.800 744.750 219.600 ;
        RECT 754.050 215.100 754.950 220.800 ;
        RECT 756.150 220.800 757.050 222.900 ;
        RECT 757.950 222.300 765.450 223.500 ;
        RECT 757.950 221.700 759.750 222.300 ;
        RECT 772.050 221.400 773.850 233.400 ;
        RECT 756.150 220.500 764.550 220.800 ;
        RECT 772.950 220.500 773.850 221.400 ;
        RECT 756.150 219.900 773.850 220.500 ;
        RECT 782.400 227.400 784.200 233.400 ;
        RECT 800.400 227.400 802.200 233.400 ;
        RECT 815.400 227.400 817.200 233.400 ;
        RECT 762.750 219.300 773.850 219.900 ;
        RECT 762.750 219.000 764.550 219.300 ;
        RECT 760.950 214.950 763.050 217.050 ;
        RECT 764.100 214.200 768.900 215.400 ;
        RECT 754.950 211.950 757.050 214.050 ;
        RECT 767.100 213.600 768.900 214.200 ;
        RECT 715.950 206.700 717.750 207.600 ;
        RECT 714.300 205.800 717.750 206.700 ;
        RECT 668.400 198.600 670.200 204.600 ;
        RECT 686.400 201.600 687.600 204.900 ;
        RECT 701.400 201.600 702.600 204.900 ;
        RECT 714.300 201.600 715.200 205.800 ;
        RECT 720.000 204.600 721.050 210.900 ;
        RECT 734.400 206.700 735.600 210.900 ;
        RECT 732.000 205.800 735.600 206.700 ;
        RECT 740.550 208.950 741.900 211.050 ;
        RECT 742.950 208.950 745.050 211.050 ;
        RECT 746.100 208.950 746.850 210.750 ;
        RECT 754.050 210.000 754.950 210.900 ;
        RECT 770.100 210.150 771.900 211.950 ;
        RECT 753.150 209.400 754.950 210.000 ;
        RECT 764.100 209.400 765.900 210.000 ;
        RECT 770.100 209.400 771.000 210.150 ;
        RECT 685.800 198.600 687.600 201.600 ;
        RECT 700.800 198.600 702.600 201.600 ;
        RECT 713.400 198.600 715.200 201.600 ;
        RECT 719.400 198.600 721.200 204.600 ;
        RECT 732.000 198.600 733.800 205.800 ;
        RECT 740.550 204.600 741.750 208.950 ;
        RECT 753.150 208.200 771.000 209.400 ;
        RECT 764.100 205.200 765.150 208.200 ;
        RECT 740.550 198.600 742.350 204.600 ;
        RECT 745.950 203.700 748.050 204.600 ;
        RECT 760.350 204.450 762.150 205.200 ;
        RECT 745.950 202.500 749.700 203.700 ;
        RECT 748.650 201.600 749.700 202.500 ;
        RECT 757.200 203.400 762.150 204.450 ;
        RECT 763.650 203.400 765.450 205.200 ;
        RECT 772.950 204.600 773.850 219.300 ;
        RECT 778.950 217.950 781.050 220.050 ;
        RECT 779.100 216.150 780.900 216.900 ;
        RECT 782.400 215.100 783.600 227.400 ;
        RECT 784.950 217.950 787.050 220.050 ;
        RECT 800.400 218.100 801.600 227.400 ;
        RECT 815.400 218.100 816.600 227.400 ;
        RECT 785.100 216.150 786.900 216.900 ;
        RECT 790.950 216.450 793.050 216.900 ;
        RECT 799.950 216.450 802.050 217.050 ;
        RECT 790.950 215.550 802.050 216.450 ;
        RECT 790.950 214.800 793.050 215.550 ;
        RECT 799.950 214.950 802.050 215.550 ;
        RECT 805.950 216.450 808.050 217.050 ;
        RECT 814.950 216.450 817.050 217.050 ;
        RECT 805.950 215.550 817.050 216.450 ;
        RECT 805.950 214.950 808.050 215.550 ;
        RECT 814.950 214.950 817.050 215.550 ;
        RECT 779.550 213.900 784.050 214.050 ;
        RECT 778.950 211.950 784.050 213.900 ;
        RECT 797.100 212.100 798.900 212.850 ;
        RECT 778.950 211.800 781.050 211.950 ;
        RECT 782.400 206.700 783.600 210.900 ;
        RECT 796.950 208.950 799.050 211.050 ;
        RECT 782.400 205.800 786.000 206.700 ;
        RECT 757.200 201.600 758.250 203.400 ;
        RECT 766.950 202.500 769.050 204.600 ;
        RECT 766.950 201.600 768.000 202.500 ;
        RECT 748.650 198.600 750.450 201.600 ;
        RECT 756.450 198.600 758.250 201.600 ;
        RECT 764.250 200.700 768.000 201.600 ;
        RECT 764.250 198.600 766.050 200.700 ;
        RECT 772.050 198.600 773.850 204.600 ;
        RECT 784.200 198.600 786.000 205.800 ;
        RECT 800.400 201.600 801.600 213.900 ;
        RECT 812.100 212.100 813.900 212.850 ;
        RECT 815.400 201.600 816.600 213.900 ;
        RECT 800.400 198.600 802.200 201.600 ;
        RECT 815.400 198.600 817.200 201.600 ;
        RECT 7.800 191.400 9.600 194.400 ;
        RECT 8.400 179.100 9.600 191.400 ;
        RECT 14.550 188.400 16.350 194.400 ;
        RECT 22.650 191.400 24.450 194.400 ;
        RECT 30.450 191.400 32.250 194.400 ;
        RECT 38.250 192.300 40.050 194.400 ;
        RECT 38.250 191.400 42.000 192.300 ;
        RECT 22.650 190.500 23.700 191.400 ;
        RECT 19.950 189.300 23.700 190.500 ;
        RECT 31.200 189.600 32.250 191.400 ;
        RECT 40.950 190.500 42.000 191.400 ;
        RECT 19.950 188.400 22.050 189.300 ;
        RECT 31.200 188.550 36.150 189.600 ;
        RECT 14.550 184.050 15.750 188.400 ;
        RECT 34.350 187.800 36.150 188.550 ;
        RECT 37.650 187.800 39.450 189.600 ;
        RECT 40.950 188.400 43.050 190.500 ;
        RECT 46.050 188.400 47.850 194.400 ;
        RECT 38.100 184.800 39.150 187.800 ;
        RECT 10.950 181.950 13.050 184.050 ;
        RECT 14.550 181.950 15.900 184.050 ;
        RECT 16.950 181.950 19.050 184.050 ;
        RECT 20.100 182.250 20.850 184.050 ;
        RECT 27.150 183.600 45.000 184.800 ;
        RECT 27.150 183.000 28.950 183.600 ;
        RECT 38.100 183.000 39.900 183.600 ;
        RECT 28.050 182.100 28.950 183.000 ;
        RECT 44.100 182.850 45.000 183.600 ;
        RECT 11.100 180.150 12.900 180.900 ;
        RECT 7.950 175.950 10.050 178.050 ;
        RECT 8.400 165.600 9.600 174.900 ;
        RECT 7.800 159.600 9.600 165.600 ;
        RECT 14.550 171.600 15.750 181.950 ;
        RECT 44.100 181.050 45.900 182.850 ;
        RECT 28.950 178.950 31.050 181.050 ;
        RECT 16.950 173.400 18.750 175.200 ;
        RECT 17.850 172.200 22.050 173.400 ;
        RECT 28.050 172.200 28.950 177.900 ;
        RECT 34.950 175.950 37.050 181.050 ;
        RECT 41.100 178.800 42.900 179.400 ;
        RECT 38.100 177.600 42.900 178.800 ;
        RECT 36.750 173.700 38.550 174.000 ;
        RECT 46.950 173.700 47.850 188.400 ;
        RECT 56.400 189.300 58.200 194.400 ;
        RECT 62.400 189.300 64.200 194.400 ;
        RECT 56.400 187.950 64.200 189.300 ;
        RECT 65.400 188.400 67.200 194.400 ;
        RECT 65.400 186.300 66.600 188.400 ;
        RECT 82.200 187.200 84.000 194.400 ;
        RECT 95.400 189.300 97.200 194.400 ;
        RECT 101.400 189.300 103.200 194.400 ;
        RECT 95.400 187.950 103.200 189.300 ;
        RECT 104.400 188.400 106.200 194.400 ;
        RECT 110.550 188.400 112.350 194.400 ;
        RECT 118.650 191.400 120.450 194.400 ;
        RECT 126.450 191.400 128.250 194.400 ;
        RECT 134.250 192.300 136.050 194.400 ;
        RECT 134.250 191.400 138.000 192.300 ;
        RECT 118.650 190.500 119.700 191.400 ;
        RECT 115.950 189.300 119.700 190.500 ;
        RECT 127.200 189.600 128.250 191.400 ;
        RECT 136.950 190.500 138.000 191.400 ;
        RECT 115.950 188.400 118.050 189.300 ;
        RECT 127.200 188.550 132.150 189.600 ;
        RECT 62.850 185.250 66.600 186.300 ;
        RECT 80.400 186.300 84.000 187.200 ;
        RECT 104.400 186.300 105.600 188.400 ;
        RECT 62.850 185.100 64.050 185.250 ;
        RECT 55.950 181.950 58.050 184.050 ;
        RECT 61.950 181.950 64.050 184.050 ;
        RECT 80.400 182.100 81.600 186.300 ;
        RECT 101.850 185.250 105.600 186.300 ;
        RECT 101.850 185.100 103.050 185.250 ;
        RECT 110.550 184.050 111.750 188.400 ;
        RECT 130.350 187.800 132.150 188.550 ;
        RECT 133.650 187.800 135.450 189.600 ;
        RECT 136.950 188.400 139.050 190.500 ;
        RECT 142.050 188.400 143.850 194.400 ;
        RECT 151.500 188.400 153.300 194.400 ;
        RECT 157.800 191.400 159.600 194.400 ;
        RECT 166.800 191.400 168.600 194.400 ;
        RECT 134.100 184.800 135.150 187.800 ;
        RECT 75.000 180.900 78.000 181.050 ;
        RECT 56.100 180.150 57.900 180.900 ;
        RECT 59.100 179.100 60.900 179.850 ;
        RECT 61.950 179.100 63.150 180.900 ;
        RECT 73.950 180.450 78.000 180.900 ;
        RECT 79.950 180.450 82.050 181.050 ;
        RECT 65.100 179.100 66.900 179.850 ;
        RECT 73.950 179.550 82.050 180.450 ;
        RECT 85.950 180.450 88.050 184.050 ;
        RECT 94.950 181.950 97.050 184.050 ;
        RECT 100.950 181.950 103.050 184.050 ;
        RECT 110.550 181.950 111.900 184.050 ;
        RECT 112.950 181.950 115.050 184.050 ;
        RECT 116.100 182.250 116.850 184.050 ;
        RECT 123.150 183.600 141.000 184.800 ;
        RECT 123.150 183.000 124.950 183.600 ;
        RECT 134.100 183.000 135.900 183.600 ;
        RECT 124.050 182.100 124.950 183.000 ;
        RECT 140.100 182.850 141.000 183.600 ;
        RECT 85.950 180.000 90.450 180.450 ;
        RECT 95.100 180.150 96.900 180.900 ;
        RECT 86.550 179.550 90.450 180.000 ;
        RECT 58.950 175.950 61.050 178.050 ;
        RECT 62.100 174.900 63.150 179.100 ;
        RECT 73.950 178.950 78.000 179.550 ;
        RECT 79.950 178.950 82.050 179.550 ;
        RECT 73.950 178.800 76.050 178.950 ;
        RECT 89.550 178.050 90.450 179.550 ;
        RECT 98.100 179.100 99.900 179.850 ;
        RECT 100.950 179.100 102.150 180.900 ;
        RECT 104.100 179.100 105.900 179.850 ;
        RECT 64.950 175.950 67.050 178.050 ;
        RECT 77.100 176.100 78.900 176.850 ;
        RECT 36.750 173.100 47.850 173.700 ;
        RECT 14.550 159.600 16.350 171.600 ;
        RECT 19.950 171.300 22.050 172.200 ;
        RECT 22.950 171.300 28.950 172.200 ;
        RECT 30.150 172.500 47.850 173.100 ;
        RECT 30.150 172.200 38.550 172.500 ;
        RECT 22.950 170.400 23.850 171.300 ;
        RECT 21.150 168.600 23.850 170.400 ;
        RECT 24.750 170.100 26.550 170.400 ;
        RECT 30.150 170.100 31.050 172.200 ;
        RECT 46.950 171.600 47.850 172.500 ;
        RECT 61.950 171.600 63.150 174.900 ;
        RECT 76.950 172.950 79.050 175.050 ;
        RECT 24.750 169.200 31.050 170.100 ;
        RECT 31.950 170.700 33.750 171.300 ;
        RECT 31.950 169.500 39.450 170.700 ;
        RECT 24.750 168.600 26.550 169.200 ;
        RECT 38.250 168.600 39.450 169.500 ;
        RECT 19.950 165.600 23.850 167.700 ;
        RECT 28.950 167.550 30.750 168.300 ;
        RECT 33.750 167.550 35.550 168.300 ;
        RECT 28.950 166.500 35.550 167.550 ;
        RECT 38.250 166.500 43.050 168.600 ;
        RECT 22.050 159.600 23.850 165.600 ;
        RECT 29.850 159.600 31.650 166.500 ;
        RECT 38.250 165.600 39.450 166.500 ;
        RECT 37.650 159.600 39.450 165.600 ;
        RECT 46.050 159.600 47.850 171.600 ;
        RECT 61.500 159.600 63.300 171.600 ;
        RECT 80.400 165.600 81.600 177.900 ;
        RECT 83.100 176.100 84.900 176.850 ;
        RECT 89.550 176.550 94.050 178.050 ;
        RECT 90.000 175.950 94.050 176.550 ;
        RECT 97.950 175.950 100.050 178.050 ;
        RECT 82.950 172.950 85.050 175.050 ;
        RECT 101.100 174.900 102.150 179.100 ;
        RECT 103.950 175.950 106.050 178.050 ;
        RECT 100.950 171.600 102.150 174.900 ;
        RECT 110.550 171.600 111.750 181.950 ;
        RECT 140.100 181.050 141.900 182.850 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 137.100 178.800 138.900 179.400 ;
        RECT 112.950 173.400 114.750 175.200 ;
        RECT 113.850 172.200 118.050 173.400 ;
        RECT 124.050 172.200 124.950 177.900 ;
        RECT 130.950 175.950 133.050 178.050 ;
        RECT 134.100 177.600 138.900 178.800 ;
        RECT 132.750 173.700 134.550 174.000 ;
        RECT 142.950 173.700 143.850 188.400 ;
        RECT 151.800 185.100 153.000 188.400 ;
        RECT 157.800 187.500 159.000 191.400 ;
        RECT 153.900 186.600 159.000 187.500 ;
        RECT 153.900 185.700 155.850 186.600 ;
        RECT 154.950 185.100 155.850 185.700 ;
        RECT 151.950 181.950 154.050 184.050 ;
        RECT 155.100 180.900 155.850 185.100 ;
        RECT 132.750 173.100 143.850 173.700 ;
        RECT 80.400 159.600 82.200 165.600 ;
        RECT 100.500 159.600 102.300 171.600 ;
        RECT 110.550 159.600 112.350 171.600 ;
        RECT 115.950 171.300 118.050 172.200 ;
        RECT 118.950 171.300 124.950 172.200 ;
        RECT 126.150 172.500 143.850 173.100 ;
        RECT 126.150 172.200 134.550 172.500 ;
        RECT 118.950 170.400 119.850 171.300 ;
        RECT 117.150 168.600 119.850 170.400 ;
        RECT 120.750 170.100 122.550 170.400 ;
        RECT 126.150 170.100 127.050 172.200 ;
        RECT 142.950 171.600 143.850 172.500 ;
        RECT 151.800 171.600 153.000 180.900 ;
        RECT 154.950 174.300 155.850 180.900 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 167.400 179.100 168.600 191.400 ;
        RECT 173.550 188.400 175.350 194.400 ;
        RECT 181.650 191.400 183.450 194.400 ;
        RECT 189.450 191.400 191.250 194.400 ;
        RECT 197.250 192.300 199.050 194.400 ;
        RECT 197.250 191.400 201.000 192.300 ;
        RECT 181.650 190.500 182.700 191.400 ;
        RECT 178.950 189.300 182.700 190.500 ;
        RECT 190.200 189.600 191.250 191.400 ;
        RECT 199.950 190.500 201.000 191.400 ;
        RECT 178.950 188.400 181.050 189.300 ;
        RECT 190.200 188.550 195.150 189.600 ;
        RECT 173.550 184.050 174.750 188.400 ;
        RECT 193.350 187.800 195.150 188.550 ;
        RECT 196.650 187.800 198.450 189.600 ;
        RECT 199.950 188.400 202.050 190.500 ;
        RECT 205.050 188.400 206.850 194.400 ;
        RECT 197.100 184.800 198.150 187.800 ;
        RECT 169.950 181.950 172.050 184.050 ;
        RECT 173.550 181.950 174.900 184.050 ;
        RECT 175.950 181.950 178.050 184.050 ;
        RECT 179.100 182.250 179.850 184.050 ;
        RECT 186.150 183.600 204.000 184.800 ;
        RECT 186.150 183.000 187.950 183.600 ;
        RECT 197.100 183.000 198.900 183.600 ;
        RECT 187.050 182.100 187.950 183.000 ;
        RECT 203.100 182.850 204.000 183.600 ;
        RECT 170.100 180.150 171.900 180.900 ;
        RECT 158.100 177.150 159.900 177.900 ;
        RECT 166.950 175.950 169.050 178.050 ;
        RECT 153.900 173.400 155.850 174.300 ;
        RECT 153.900 172.500 159.600 173.400 ;
        RECT 120.750 169.200 127.050 170.100 ;
        RECT 127.950 170.700 129.750 171.300 ;
        RECT 127.950 169.500 135.450 170.700 ;
        RECT 120.750 168.600 122.550 169.200 ;
        RECT 134.250 168.600 135.450 169.500 ;
        RECT 115.950 165.600 119.850 167.700 ;
        RECT 124.950 167.550 126.750 168.300 ;
        RECT 129.750 167.550 131.550 168.300 ;
        RECT 124.950 166.500 131.550 167.550 ;
        RECT 134.250 166.500 139.050 168.600 ;
        RECT 118.050 159.600 119.850 165.600 ;
        RECT 125.850 159.600 127.650 166.500 ;
        RECT 134.250 165.600 135.450 166.500 ;
        RECT 133.650 159.600 135.450 165.600 ;
        RECT 142.050 159.600 143.850 171.600 ;
        RECT 151.500 159.600 153.300 171.600 ;
        RECT 158.400 165.600 159.600 172.500 ;
        RECT 167.400 165.600 168.600 174.900 ;
        RECT 157.800 159.600 159.600 165.600 ;
        RECT 166.800 159.600 168.600 165.600 ;
        RECT 173.550 171.600 174.750 181.950 ;
        RECT 203.100 181.050 204.900 182.850 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 175.950 173.400 177.750 175.200 ;
        RECT 176.850 172.200 181.050 173.400 ;
        RECT 187.050 172.200 187.950 177.900 ;
        RECT 193.950 175.950 196.050 181.050 ;
        RECT 200.100 178.800 201.900 179.400 ;
        RECT 197.100 177.600 201.900 178.800 ;
        RECT 195.750 173.700 197.550 174.000 ;
        RECT 205.950 173.700 206.850 188.400 ;
        RECT 212.400 189.300 214.200 194.400 ;
        RECT 218.400 189.300 220.200 194.400 ;
        RECT 212.400 187.950 220.200 189.300 ;
        RECT 221.400 188.400 223.200 194.400 ;
        RECT 221.400 186.300 222.600 188.400 ;
        RECT 238.800 187.500 240.600 194.400 ;
        RECT 244.800 187.500 246.600 194.400 ;
        RECT 250.800 187.500 252.600 194.400 ;
        RECT 256.800 187.500 258.600 194.400 ;
        RECT 269.400 189.300 271.200 194.400 ;
        RECT 275.400 189.300 277.200 194.400 ;
        RECT 269.400 187.950 277.200 189.300 ;
        RECT 278.400 188.400 280.200 194.400 ;
        RECT 294.300 190.200 296.100 194.400 ;
        RECT 294.150 188.400 296.100 190.200 ;
        RECT 218.850 185.250 222.600 186.300 ;
        RECT 237.900 186.300 240.600 187.500 ;
        RECT 242.700 186.300 246.600 187.500 ;
        RECT 248.700 186.300 252.600 187.500 ;
        RECT 254.700 186.300 258.600 187.500 ;
        RECT 278.400 186.300 279.600 188.400 ;
        RECT 218.850 185.100 220.050 185.250 ;
        RECT 211.950 181.950 214.050 184.050 ;
        RECT 217.950 181.950 220.050 184.050 ;
        RECT 237.900 182.100 238.800 186.300 ;
        RECT 242.700 185.400 243.900 186.300 ;
        RECT 248.700 185.400 249.900 186.300 ;
        RECT 254.700 185.400 255.900 186.300 ;
        RECT 239.700 184.200 243.900 185.400 ;
        RECT 239.700 183.600 241.500 184.200 ;
        RECT 212.100 180.150 213.900 180.900 ;
        RECT 215.100 179.100 216.900 179.850 ;
        RECT 217.950 179.100 219.150 180.900 ;
        RECT 229.950 180.450 234.000 181.050 ;
        RECT 235.950 180.450 238.050 181.050 ;
        RECT 221.100 179.100 222.900 179.850 ;
        RECT 229.950 179.550 238.050 180.450 ;
        RECT 214.950 175.950 217.050 178.050 ;
        RECT 218.100 174.900 219.150 179.100 ;
        RECT 229.950 178.950 234.000 179.550 ;
        RECT 235.950 178.950 238.050 179.550 ;
        RECT 220.950 175.950 223.050 178.050 ;
        RECT 195.750 173.100 206.850 173.700 ;
        RECT 173.550 159.600 175.350 171.600 ;
        RECT 178.950 171.300 181.050 172.200 ;
        RECT 181.950 171.300 187.950 172.200 ;
        RECT 189.150 172.500 206.850 173.100 ;
        RECT 189.150 172.200 197.550 172.500 ;
        RECT 181.950 170.400 182.850 171.300 ;
        RECT 180.150 168.600 182.850 170.400 ;
        RECT 183.750 170.100 185.550 170.400 ;
        RECT 189.150 170.100 190.050 172.200 ;
        RECT 205.950 171.600 206.850 172.500 ;
        RECT 217.950 171.600 219.150 174.900 ;
        RECT 237.900 173.700 238.800 177.900 ;
        RECT 242.700 173.700 243.900 184.200 ;
        RECT 245.700 184.200 249.900 185.400 ;
        RECT 245.700 183.600 247.500 184.200 ;
        RECT 248.700 173.700 249.900 184.200 ;
        RECT 251.700 184.200 255.900 185.400 ;
        RECT 275.850 185.250 279.600 186.300 ;
        RECT 275.850 185.100 277.050 185.250 ;
        RECT 294.150 185.100 295.050 188.400 ;
        RECT 296.100 186.600 297.900 187.500 ;
        RECT 301.800 186.600 303.600 194.400 ;
        RECT 314.400 191.400 316.200 194.400 ;
        RECT 314.400 188.100 315.600 191.400 ;
        RECT 326.400 189.300 328.200 194.400 ;
        RECT 332.400 189.300 334.200 194.400 ;
        RECT 326.400 187.950 334.200 189.300 ;
        RECT 335.400 188.400 337.200 194.400 ;
        RECT 350.400 191.400 352.200 194.400 ;
        RECT 296.100 185.700 303.600 186.600 ;
        RECT 307.950 186.450 312.000 187.050 ;
        RECT 313.950 186.450 316.050 187.050 ;
        RECT 251.700 183.600 253.500 184.200 ;
        RECT 254.700 173.700 255.900 184.200 ;
        RECT 257.100 182.100 258.900 182.850 ;
        RECT 268.950 181.950 271.050 184.050 ;
        RECT 274.950 183.450 277.050 184.050 ;
        RECT 274.950 182.550 288.450 183.450 ;
        RECT 274.950 181.950 277.050 182.550 ;
        RECT 269.100 180.150 270.900 180.900 ;
        RECT 272.100 179.100 273.900 179.850 ;
        RECT 274.950 179.100 276.150 180.900 ;
        RECT 278.100 179.100 279.900 179.850 ;
        RECT 271.950 175.950 274.050 178.050 ;
        RECT 275.100 174.900 276.150 179.100 ;
        RECT 277.950 175.950 280.050 178.050 ;
        RECT 287.550 177.900 288.450 182.550 ;
        RECT 289.950 181.950 295.050 184.050 ;
        RECT 286.950 175.800 289.050 177.900 ;
        RECT 237.900 172.500 240.600 173.700 ;
        RECT 242.700 172.500 246.600 173.700 ;
        RECT 248.700 172.500 252.600 173.700 ;
        RECT 254.700 172.500 258.600 173.700 ;
        RECT 183.750 169.200 190.050 170.100 ;
        RECT 190.950 170.700 192.750 171.300 ;
        RECT 190.950 169.500 198.450 170.700 ;
        RECT 183.750 168.600 185.550 169.200 ;
        RECT 197.250 168.600 198.450 169.500 ;
        RECT 178.950 165.600 182.850 167.700 ;
        RECT 187.950 167.550 189.750 168.300 ;
        RECT 192.750 167.550 194.550 168.300 ;
        RECT 187.950 166.500 194.550 167.550 ;
        RECT 197.250 166.500 202.050 168.600 ;
        RECT 181.050 159.600 182.850 165.600 ;
        RECT 188.850 159.600 190.650 166.500 ;
        RECT 197.250 165.600 198.450 166.500 ;
        RECT 196.650 159.600 198.450 165.600 ;
        RECT 205.050 159.600 206.850 171.600 ;
        RECT 217.500 159.600 219.300 171.600 ;
        RECT 238.800 159.600 240.600 172.500 ;
        RECT 244.800 159.600 246.600 172.500 ;
        RECT 250.800 159.600 252.600 172.500 ;
        RECT 256.800 159.600 258.600 172.500 ;
        RECT 274.950 171.600 276.150 174.900 ;
        RECT 292.950 171.600 294.000 180.900 ;
        RECT 296.100 179.100 297.900 179.850 ;
        RECT 295.950 175.950 298.050 178.050 ;
        RECT 274.500 159.600 276.300 171.600 ;
        RECT 292.200 159.600 294.000 171.600 ;
        RECT 299.550 165.600 300.600 185.700 ;
        RECT 307.950 185.550 316.050 186.450 ;
        RECT 335.400 186.300 336.600 188.400 ;
        RECT 307.950 184.950 312.000 185.550 ;
        RECT 313.950 184.950 316.050 185.550 ;
        RECT 332.850 185.250 336.600 186.300 ;
        RECT 332.850 185.100 334.050 185.250 ;
        RECT 337.950 184.050 340.050 184.200 ;
        RECT 314.700 182.100 316.050 183.900 ;
        RECT 301.950 178.950 304.050 181.050 ;
        RECT 302.100 177.150 303.900 177.900 ;
        RECT 310.950 175.950 313.050 178.050 ;
        RECT 314.700 177.900 315.900 182.100 ;
        RECT 325.950 181.950 328.050 184.050 ;
        RECT 331.950 183.450 334.050 184.050 ;
        RECT 336.000 183.450 340.050 184.050 ;
        RECT 331.950 182.550 340.050 183.450 ;
        RECT 331.950 181.950 334.050 182.550 ;
        RECT 336.000 182.100 340.050 182.550 ;
        RECT 336.000 181.950 339.000 182.100 ;
        RECT 346.950 181.950 349.050 184.050 ;
        RECT 316.950 178.950 319.050 181.050 ;
        RECT 326.100 180.150 327.900 180.900 ;
        RECT 329.100 179.100 330.900 179.850 ;
        RECT 331.950 179.100 333.150 180.900 ;
        RECT 335.100 179.100 336.900 179.850 ;
        RECT 311.100 174.150 312.900 174.900 ;
        RECT 314.700 172.650 316.050 177.900 ;
        RECT 317.100 177.150 318.900 177.900 ;
        RECT 328.950 175.800 331.050 178.050 ;
        RECT 332.100 174.900 333.150 179.100 ;
        RECT 334.950 175.950 337.050 178.050 ;
        RECT 340.950 177.450 343.050 180.900 ;
        RECT 347.100 180.150 348.900 180.900 ;
        RECT 350.400 179.100 351.600 191.400 ;
        RECT 356.550 188.400 358.350 194.400 ;
        RECT 364.650 191.400 366.450 194.400 ;
        RECT 372.450 191.400 374.250 194.400 ;
        RECT 380.250 192.300 382.050 194.400 ;
        RECT 380.250 191.400 384.000 192.300 ;
        RECT 364.650 190.500 365.700 191.400 ;
        RECT 361.950 189.300 365.700 190.500 ;
        RECT 373.200 189.600 374.250 191.400 ;
        RECT 382.950 190.500 384.000 191.400 ;
        RECT 361.950 188.400 364.050 189.300 ;
        RECT 373.200 188.550 378.150 189.600 ;
        RECT 356.550 184.050 357.750 188.400 ;
        RECT 376.350 187.800 378.150 188.550 ;
        RECT 379.650 187.800 381.450 189.600 ;
        RECT 382.950 188.400 385.050 190.500 ;
        RECT 388.050 188.400 389.850 194.400 ;
        RECT 400.800 191.400 402.600 194.400 ;
        RECT 380.100 184.800 381.150 187.800 ;
        RECT 356.550 181.950 357.900 184.050 ;
        RECT 358.950 181.950 361.050 184.050 ;
        RECT 362.100 182.250 362.850 184.050 ;
        RECT 369.150 183.600 387.000 184.800 ;
        RECT 369.150 183.000 370.950 183.600 ;
        RECT 380.100 183.000 381.900 183.600 ;
        RECT 370.050 182.100 370.950 183.000 ;
        RECT 386.100 182.850 387.000 183.600 ;
        RECT 349.950 177.450 352.050 178.050 ;
        RECT 340.950 177.000 352.050 177.450 ;
        RECT 341.550 176.550 352.050 177.000 ;
        RECT 349.950 175.950 352.050 176.550 ;
        RECT 314.700 171.600 317.400 172.650 ;
        RECT 331.950 171.600 333.150 174.900 ;
        RECT 298.800 159.600 300.600 165.600 ;
        RECT 315.600 159.600 317.400 171.600 ;
        RECT 331.500 159.600 333.300 171.600 ;
        RECT 337.950 171.450 340.050 172.050 ;
        RECT 346.950 171.450 349.050 172.050 ;
        RECT 337.950 170.550 349.050 171.450 ;
        RECT 337.950 169.950 340.050 170.550 ;
        RECT 346.950 169.950 349.050 170.550 ;
        RECT 350.400 165.600 351.600 174.900 ;
        RECT 356.550 171.600 357.750 181.950 ;
        RECT 386.100 181.050 387.900 182.850 ;
        RECT 370.950 178.950 373.050 181.050 ;
        RECT 383.100 178.800 384.900 179.400 ;
        RECT 358.950 173.400 360.750 175.200 ;
        RECT 359.850 172.200 364.050 173.400 ;
        RECT 370.050 172.200 370.950 177.900 ;
        RECT 376.950 175.950 379.050 178.050 ;
        RECT 380.100 177.600 384.900 178.800 ;
        RECT 378.750 173.700 380.550 174.000 ;
        RECT 388.950 173.700 389.850 188.400 ;
        RECT 401.400 188.100 402.600 191.400 ;
        RECT 420.000 190.050 421.800 194.400 ;
        RECT 416.400 188.400 421.800 190.050 ;
        RECT 400.950 186.450 403.050 187.050 ;
        RECT 409.950 186.450 412.050 187.050 ;
        RECT 400.950 185.550 412.050 186.450 ;
        RECT 400.950 184.950 403.050 185.550 ;
        RECT 409.950 184.950 412.050 185.550 ;
        RECT 416.400 185.100 417.300 188.400 ;
        RECT 436.800 187.500 438.600 194.400 ;
        RECT 442.800 187.500 444.600 194.400 ;
        RECT 448.800 187.500 450.600 194.400 ;
        RECT 454.800 187.500 456.600 194.400 ;
        RECT 435.900 186.300 438.600 187.500 ;
        RECT 440.700 186.300 444.600 187.500 ;
        RECT 446.700 186.300 450.600 187.500 ;
        RECT 452.700 186.300 456.600 187.500 ;
        RECT 470.400 187.500 472.200 194.400 ;
        RECT 476.400 187.500 478.200 194.400 ;
        RECT 482.400 187.500 484.200 194.400 ;
        RECT 488.400 187.500 490.200 194.400 ;
        RECT 470.400 186.300 474.300 187.500 ;
        RECT 476.400 186.300 480.300 187.500 ;
        RECT 482.400 186.300 486.300 187.500 ;
        RECT 488.400 186.300 491.100 187.500 ;
        RECT 507.000 187.200 508.800 194.400 ;
        RECT 523.800 188.400 525.600 194.400 ;
        RECT 507.000 186.300 510.600 187.200 ;
        RECT 400.950 182.100 402.300 183.900 ;
        RECT 391.950 180.450 396.000 181.050 ;
        RECT 397.950 180.450 400.050 181.050 ;
        RECT 391.950 179.550 400.050 180.450 ;
        RECT 391.950 178.950 396.000 179.550 ;
        RECT 397.950 178.950 400.050 179.550 ;
        RECT 401.100 177.900 402.300 182.100 ;
        RECT 406.950 183.450 409.050 184.050 ;
        RECT 415.950 183.450 418.050 184.050 ;
        RECT 406.950 182.550 418.050 183.450 ;
        RECT 406.950 181.950 409.050 182.550 ;
        RECT 415.950 181.950 418.050 182.550 ;
        RECT 421.950 181.950 424.050 184.050 ;
        RECT 435.900 182.100 436.800 186.300 ;
        RECT 440.700 185.400 441.900 186.300 ;
        RECT 446.700 185.400 447.900 186.300 ;
        RECT 452.700 185.400 453.900 186.300 ;
        RECT 437.700 184.200 441.900 185.400 ;
        RECT 437.700 183.600 439.500 184.200 ;
        RECT 431.550 180.900 436.050 181.050 ;
        RECT 398.100 177.150 399.900 177.900 ;
        RECT 378.750 173.100 389.850 173.700 ;
        RECT 350.400 159.600 352.200 165.600 ;
        RECT 356.550 159.600 358.350 171.600 ;
        RECT 361.950 171.300 364.050 172.200 ;
        RECT 364.950 171.300 370.950 172.200 ;
        RECT 372.150 172.500 389.850 173.100 ;
        RECT 400.950 172.650 402.300 177.900 ;
        RECT 403.950 175.950 406.050 178.050 ;
        RECT 404.100 174.150 405.900 174.900 ;
        RECT 372.150 172.200 380.550 172.500 ;
        RECT 364.950 170.400 365.850 171.300 ;
        RECT 363.150 168.600 365.850 170.400 ;
        RECT 366.750 170.100 368.550 170.400 ;
        RECT 372.150 170.100 373.050 172.200 ;
        RECT 388.950 171.600 389.850 172.500 ;
        RECT 366.750 169.200 373.050 170.100 ;
        RECT 373.950 170.700 375.750 171.300 ;
        RECT 373.950 169.500 381.450 170.700 ;
        RECT 366.750 168.600 368.550 169.200 ;
        RECT 380.250 168.600 381.450 169.500 ;
        RECT 361.950 165.600 365.850 167.700 ;
        RECT 370.950 167.550 372.750 168.300 ;
        RECT 375.750 167.550 377.550 168.300 ;
        RECT 370.950 166.500 377.550 167.550 ;
        RECT 380.250 166.500 385.050 168.600 ;
        RECT 364.050 159.600 365.850 165.600 ;
        RECT 371.850 159.600 373.650 166.500 ;
        RECT 380.250 165.600 381.450 166.500 ;
        RECT 379.650 159.600 381.450 165.600 ;
        RECT 388.050 159.600 389.850 171.600 ;
        RECT 399.600 171.600 402.300 172.650 ;
        RECT 416.400 171.600 417.300 180.900 ;
        RECT 422.100 180.150 423.900 180.900 ;
        RECT 419.100 179.100 420.900 179.850 ;
        RECT 425.100 179.100 426.900 179.850 ;
        RECT 430.950 178.950 436.050 180.900 ;
        RECT 430.950 178.800 433.050 178.950 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 424.950 175.950 427.050 178.050 ;
        RECT 435.900 173.700 436.800 177.900 ;
        RECT 440.700 173.700 441.900 184.200 ;
        RECT 443.700 184.200 447.900 185.400 ;
        RECT 443.700 183.600 445.500 184.200 ;
        RECT 446.700 173.700 447.900 184.200 ;
        RECT 449.700 184.200 453.900 185.400 ;
        RECT 449.700 183.600 451.500 184.200 ;
        RECT 452.700 173.700 453.900 184.200 ;
        RECT 473.100 185.400 474.300 186.300 ;
        RECT 479.100 185.400 480.300 186.300 ;
        RECT 485.100 185.400 486.300 186.300 ;
        RECT 473.100 184.200 477.300 185.400 ;
        RECT 455.100 182.100 456.900 182.850 ;
        RECT 470.100 182.100 471.900 182.850 ;
        RECT 473.100 173.700 474.300 184.200 ;
        RECT 475.500 183.600 477.300 184.200 ;
        RECT 479.100 184.200 483.300 185.400 ;
        RECT 479.100 173.700 480.300 184.200 ;
        RECT 481.500 183.600 483.300 184.200 ;
        RECT 485.100 184.200 489.300 185.400 ;
        RECT 485.100 173.700 486.300 184.200 ;
        RECT 487.500 183.600 489.300 184.200 ;
        RECT 490.200 182.100 491.100 186.300 ;
        RECT 509.400 182.100 510.600 186.300 ;
        RECT 524.400 186.300 525.600 188.400 ;
        RECT 526.800 189.300 528.600 194.400 ;
        RECT 532.800 189.300 534.600 194.400 ;
        RECT 526.800 187.950 534.600 189.300 ;
        RECT 536.550 188.400 538.350 194.400 ;
        RECT 544.650 191.400 546.450 194.400 ;
        RECT 552.450 191.400 554.250 194.400 ;
        RECT 560.250 192.300 562.050 194.400 ;
        RECT 560.250 191.400 564.000 192.300 ;
        RECT 544.650 190.500 545.700 191.400 ;
        RECT 541.950 189.300 545.700 190.500 ;
        RECT 553.200 189.600 554.250 191.400 ;
        RECT 562.950 190.500 564.000 191.400 ;
        RECT 541.950 188.400 544.050 189.300 ;
        RECT 553.200 188.550 558.150 189.600 ;
        RECT 524.400 185.250 528.150 186.300 ;
        RECT 526.950 185.100 528.150 185.250 ;
        RECT 536.550 184.050 537.750 188.400 ;
        RECT 556.350 187.800 558.150 188.550 ;
        RECT 559.650 187.800 561.450 189.600 ;
        RECT 562.950 188.400 565.050 190.500 ;
        RECT 568.050 188.400 569.850 194.400 ;
        RECT 580.800 188.400 582.600 194.400 ;
        RECT 560.100 184.800 561.150 187.800 ;
        RECT 523.950 181.950 529.050 184.050 ;
        RECT 532.950 181.950 535.050 184.050 ;
        RECT 536.550 181.950 537.900 184.050 ;
        RECT 538.950 181.950 541.050 184.050 ;
        RECT 542.100 182.250 542.850 184.050 ;
        RECT 549.150 183.600 567.000 184.800 ;
        RECT 549.150 183.000 550.950 183.600 ;
        RECT 560.100 183.000 561.900 183.600 ;
        RECT 550.050 182.100 550.950 183.000 ;
        RECT 566.100 182.850 567.000 183.600 ;
        RECT 490.950 178.950 496.050 181.050 ;
        RECT 508.950 180.450 511.050 181.050 ;
        RECT 517.950 180.450 520.050 181.050 ;
        RECT 508.950 179.550 520.050 180.450 ;
        RECT 508.950 178.950 511.050 179.550 ;
        RECT 517.950 178.950 520.050 179.550 ;
        RECT 524.100 179.100 525.900 179.850 ;
        RECT 527.850 179.100 529.050 180.900 ;
        RECT 533.100 180.150 534.900 180.900 ;
        RECT 530.100 179.100 531.900 179.850 ;
        RECT 490.200 173.700 491.100 177.900 ;
        RECT 506.100 176.100 507.900 176.850 ;
        RECT 435.900 172.500 438.600 173.700 ;
        RECT 440.700 172.500 444.600 173.700 ;
        RECT 446.700 172.500 450.600 173.700 ;
        RECT 452.700 172.500 456.600 173.700 ;
        RECT 399.600 159.600 401.400 171.600 ;
        RECT 415.800 159.600 417.600 171.600 ;
        RECT 418.800 170.700 426.600 171.600 ;
        RECT 418.800 159.600 420.600 170.700 ;
        RECT 424.800 159.600 426.600 170.700 ;
        RECT 436.800 159.600 438.600 172.500 ;
        RECT 442.800 159.600 444.600 172.500 ;
        RECT 448.800 159.600 450.600 172.500 ;
        RECT 454.800 159.600 456.600 172.500 ;
        RECT 470.400 172.500 474.300 173.700 ;
        RECT 476.400 172.500 480.300 173.700 ;
        RECT 482.400 172.500 486.300 173.700 ;
        RECT 488.400 172.500 491.100 173.700 ;
        RECT 505.950 172.950 508.050 175.050 ;
        RECT 470.400 159.600 472.200 172.500 ;
        RECT 476.400 159.600 478.200 172.500 ;
        RECT 482.400 159.600 484.200 172.500 ;
        RECT 488.400 159.600 490.200 172.500 ;
        RECT 509.400 165.600 510.600 177.900 ;
        RECT 512.100 176.100 513.900 176.850 ;
        RECT 523.950 175.950 526.050 178.050 ;
        RECT 511.950 172.950 517.050 175.050 ;
        RECT 527.850 174.900 528.900 179.100 ;
        RECT 529.950 175.950 532.050 178.050 ;
        RECT 527.850 171.600 529.050 174.900 ;
        RECT 536.550 171.600 537.750 181.950 ;
        RECT 566.100 181.050 567.900 182.850 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 563.100 178.800 564.900 179.400 ;
        RECT 538.950 173.400 540.750 175.200 ;
        RECT 539.850 172.200 544.050 173.400 ;
        RECT 550.050 172.200 550.950 177.900 ;
        RECT 556.950 175.950 559.050 178.050 ;
        RECT 560.100 177.600 564.900 178.800 ;
        RECT 558.750 173.700 560.550 174.000 ;
        RECT 568.950 173.700 569.850 188.400 ;
        RECT 581.400 186.300 582.600 188.400 ;
        RECT 583.800 189.300 585.600 194.400 ;
        RECT 589.800 189.300 591.600 194.400 ;
        RECT 603.300 190.200 605.100 194.400 ;
        RECT 583.800 187.950 591.600 189.300 ;
        RECT 603.150 188.400 605.100 190.200 ;
        RECT 581.400 185.250 585.150 186.300 ;
        RECT 583.950 185.100 585.150 185.250 ;
        RECT 603.150 185.100 604.050 188.400 ;
        RECT 605.100 186.600 606.900 187.500 ;
        RECT 610.800 186.600 612.600 194.400 ;
        RECT 617.400 189.300 619.200 194.400 ;
        RECT 623.400 189.300 625.200 194.400 ;
        RECT 617.400 187.950 625.200 189.300 ;
        RECT 626.400 188.400 628.200 194.400 ;
        RECT 635.400 191.400 637.200 194.400 ;
        RECT 605.100 185.700 612.600 186.600 ;
        RECT 626.400 186.300 627.600 188.400 ;
        RECT 636.000 187.500 637.200 191.400 ;
        RECT 641.700 188.400 643.500 194.400 ;
        RECT 653.400 191.400 655.200 194.400 ;
        RECT 668.400 191.400 670.200 194.400 ;
        RECT 636.000 186.600 641.100 187.500 ;
        RECT 571.950 183.450 574.050 184.050 ;
        RECT 583.950 183.450 586.050 184.050 ;
        RECT 571.950 182.550 586.050 183.450 ;
        RECT 571.950 181.950 574.050 182.550 ;
        RECT 583.950 181.950 586.050 182.550 ;
        RECT 589.950 181.950 592.050 184.050 ;
        RECT 601.950 181.950 604.050 184.050 ;
        RECT 581.100 179.100 582.900 179.850 ;
        RECT 584.850 179.100 586.050 180.900 ;
        RECT 590.100 180.150 591.900 180.900 ;
        RECT 587.100 179.100 588.900 179.850 ;
        RECT 580.950 175.950 583.050 178.050 ;
        RECT 558.750 173.100 569.850 173.700 ;
        RECT 508.800 159.600 510.600 165.600 ;
        RECT 527.700 159.600 529.500 171.600 ;
        RECT 536.550 159.600 538.350 171.600 ;
        RECT 541.950 171.300 544.050 172.200 ;
        RECT 544.950 171.300 550.950 172.200 ;
        RECT 552.150 172.500 569.850 173.100 ;
        RECT 552.150 172.200 560.550 172.500 ;
        RECT 544.950 170.400 545.850 171.300 ;
        RECT 543.150 168.600 545.850 170.400 ;
        RECT 546.750 170.100 548.550 170.400 ;
        RECT 552.150 170.100 553.050 172.200 ;
        RECT 568.950 171.600 569.850 172.500 ;
        RECT 584.850 174.900 585.900 179.100 ;
        RECT 586.950 175.950 589.050 178.050 ;
        RECT 584.850 171.600 586.050 174.900 ;
        RECT 601.950 171.600 603.000 180.900 ;
        RECT 605.100 179.100 606.900 179.850 ;
        RECT 604.950 175.950 607.050 178.050 ;
        RECT 546.750 169.200 553.050 170.100 ;
        RECT 553.950 170.700 555.750 171.300 ;
        RECT 553.950 169.500 561.450 170.700 ;
        RECT 546.750 168.600 548.550 169.200 ;
        RECT 560.250 168.600 561.450 169.500 ;
        RECT 541.950 165.600 545.850 167.700 ;
        RECT 550.950 167.550 552.750 168.300 ;
        RECT 555.750 167.550 557.550 168.300 ;
        RECT 550.950 166.500 557.550 167.550 ;
        RECT 560.250 166.500 565.050 168.600 ;
        RECT 544.050 159.600 545.850 165.600 ;
        RECT 551.850 159.600 553.650 166.500 ;
        RECT 560.250 165.600 561.450 166.500 ;
        RECT 559.650 159.600 561.450 165.600 ;
        RECT 568.050 159.600 569.850 171.600 ;
        RECT 584.700 159.600 586.500 171.600 ;
        RECT 601.200 159.600 603.000 171.600 ;
        RECT 608.550 165.600 609.600 185.700 ;
        RECT 623.850 185.250 627.600 186.300 ;
        RECT 639.150 185.700 641.100 186.600 ;
        RECT 623.850 185.100 625.050 185.250 ;
        RECT 639.150 185.100 640.050 185.700 ;
        RECT 642.000 185.100 643.200 188.400 ;
        RECT 616.950 181.950 619.050 184.050 ;
        RECT 622.950 181.950 625.050 184.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 617.100 180.150 618.900 180.900 ;
        RECT 620.100 179.100 621.900 179.850 ;
        RECT 622.950 179.100 624.150 180.900 ;
        RECT 626.100 179.100 627.900 179.850 ;
        RECT 611.100 177.150 612.900 177.900 ;
        RECT 619.950 175.950 622.050 178.050 ;
        RECT 623.100 174.900 624.150 179.100 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 639.150 180.900 639.900 185.100 ;
        RECT 640.950 181.950 643.050 184.050 ;
        RECT 649.950 181.950 652.050 184.050 ;
        RECT 625.950 175.950 628.050 178.050 ;
        RECT 635.100 177.150 636.900 177.900 ;
        RECT 622.950 171.600 624.150 174.900 ;
        RECT 639.150 174.300 640.050 180.900 ;
        RECT 639.150 173.400 641.100 174.300 ;
        RECT 635.400 172.500 641.100 173.400 ;
        RECT 607.800 159.600 609.600 165.600 ;
        RECT 622.500 159.600 624.300 171.600 ;
        RECT 635.400 165.600 636.600 172.500 ;
        RECT 642.000 171.600 643.200 180.900 ;
        RECT 650.100 180.150 651.900 180.900 ;
        RECT 653.400 179.100 654.600 191.400 ;
        RECT 664.950 181.950 667.050 184.050 ;
        RECT 665.100 180.150 666.900 180.900 ;
        RECT 668.400 179.100 669.600 191.400 ;
        RECT 679.800 188.400 681.600 194.400 ;
        RECT 680.400 186.300 681.600 188.400 ;
        RECT 682.800 189.300 684.600 194.400 ;
        RECT 688.800 189.300 690.600 194.400 ;
        RECT 682.800 187.950 690.600 189.300 ;
        RECT 701.400 191.400 703.200 194.400 ;
        RECT 719.400 191.400 721.200 194.400 ;
        RECT 737.400 191.400 739.200 194.400 ;
        RECT 748.800 191.400 750.600 194.400 ;
        RECT 701.400 188.100 702.600 191.400 ;
        RECT 719.400 188.100 720.600 191.400 ;
        RECT 700.950 186.450 703.050 187.050 ;
        RECT 709.950 186.450 712.050 187.050 ;
        RECT 680.400 185.250 684.150 186.300 ;
        RECT 682.950 185.100 684.150 185.250 ;
        RECT 700.950 185.550 712.050 186.450 ;
        RECT 700.950 184.950 703.050 185.550 ;
        RECT 709.950 184.950 712.050 185.550 ;
        RECT 718.950 186.450 721.050 187.050 ;
        RECT 727.950 186.450 730.050 187.050 ;
        RECT 718.950 185.550 730.050 186.450 ;
        RECT 718.950 184.950 721.050 185.550 ;
        RECT 727.950 184.950 730.050 185.550 ;
        RECT 673.950 183.450 676.050 184.050 ;
        RECT 682.950 183.450 685.050 184.050 ;
        RECT 673.950 182.550 685.050 183.450 ;
        RECT 673.950 181.950 676.050 182.550 ;
        RECT 682.950 181.950 685.050 182.550 ;
        RECT 688.950 183.450 691.050 184.050 ;
        RECT 693.000 183.450 697.050 184.050 ;
        RECT 688.950 182.550 697.050 183.450 ;
        RECT 688.950 181.950 691.050 182.550 ;
        RECT 693.000 181.950 697.050 182.550 ;
        RECT 701.700 182.100 703.050 183.900 ;
        RECT 719.700 182.100 721.050 183.900 ;
        RECT 680.100 179.100 681.900 179.850 ;
        RECT 683.850 179.100 685.050 180.900 ;
        RECT 689.100 180.150 690.900 180.900 ;
        RECT 686.100 179.100 687.900 179.850 ;
        RECT 652.950 175.950 655.050 178.050 ;
        RECT 667.950 175.950 673.050 178.050 ;
        RECT 679.950 175.950 682.050 178.050 ;
        RECT 683.850 174.900 684.900 179.100 ;
        RECT 685.950 175.950 688.050 178.050 ;
        RECT 697.950 175.800 700.050 178.050 ;
        RECT 701.700 177.900 702.900 182.100 ;
        RECT 703.950 178.950 706.050 181.050 ;
        RECT 635.400 159.600 637.200 165.600 ;
        RECT 641.700 159.600 643.500 171.600 ;
        RECT 653.400 165.600 654.600 174.900 ;
        RECT 668.400 165.600 669.600 174.900 ;
        RECT 683.850 171.600 685.050 174.900 ;
        RECT 698.100 174.150 699.900 174.900 ;
        RECT 701.700 172.650 703.050 177.900 ;
        RECT 704.100 177.150 705.900 177.900 ;
        RECT 715.950 175.950 718.050 178.050 ;
        RECT 719.700 177.900 720.900 182.100 ;
        RECT 733.950 181.950 736.050 184.050 ;
        RECT 721.950 178.950 727.050 181.050 ;
        RECT 734.100 180.150 735.900 180.900 ;
        RECT 737.400 179.100 738.600 191.400 ;
        RECT 749.400 179.100 750.600 191.400 ;
        RECT 761.400 189.300 763.200 194.400 ;
        RECT 767.400 189.300 769.200 194.400 ;
        RECT 761.400 187.950 769.200 189.300 ;
        RECT 770.400 188.400 772.200 194.400 ;
        RECT 770.400 186.300 771.600 188.400 ;
        RECT 783.000 187.200 784.800 194.400 ;
        RECT 792.150 188.400 793.950 194.400 ;
        RECT 799.950 192.300 801.750 194.400 ;
        RECT 798.000 191.400 801.750 192.300 ;
        RECT 807.750 191.400 809.550 194.400 ;
        RECT 815.550 191.400 817.350 194.400 ;
        RECT 798.000 190.500 799.050 191.400 ;
        RECT 796.950 188.400 799.050 190.500 ;
        RECT 807.750 189.600 808.800 191.400 ;
        RECT 783.000 186.300 786.600 187.200 ;
        RECT 767.850 185.250 771.600 186.300 ;
        RECT 767.850 185.100 769.050 185.250 ;
        RECT 751.950 181.950 754.050 184.050 ;
        RECT 760.950 181.950 763.050 184.050 ;
        RECT 766.950 183.450 769.050 184.050 ;
        RECT 778.950 183.450 781.050 184.050 ;
        RECT 766.950 182.550 781.050 183.450 ;
        RECT 766.950 181.950 769.050 182.550 ;
        RECT 778.950 181.950 781.050 182.550 ;
        RECT 785.400 182.100 786.600 186.300 ;
        RECT 752.100 180.150 753.900 180.900 ;
        RECT 761.100 180.150 762.900 180.900 ;
        RECT 764.100 179.100 765.900 179.850 ;
        RECT 766.950 179.100 768.150 180.900 ;
        RECT 784.950 180.450 787.050 181.050 ;
        RECT 770.100 179.100 771.900 179.850 ;
        RECT 776.550 179.550 787.050 180.450 ;
        RECT 716.100 174.150 717.900 174.900 ;
        RECT 719.700 172.650 721.050 177.900 ;
        RECT 722.100 177.150 723.900 177.900 ;
        RECT 736.950 177.450 739.050 178.050 ;
        RECT 741.000 177.450 745.050 178.050 ;
        RECT 736.950 176.550 745.050 177.450 ;
        RECT 736.950 175.950 739.050 176.550 ;
        RECT 741.000 175.950 745.050 176.550 ;
        RECT 748.950 177.450 751.050 178.050 ;
        RECT 753.000 177.450 757.050 178.050 ;
        RECT 748.950 176.550 757.050 177.450 ;
        RECT 748.950 175.950 751.050 176.550 ;
        RECT 753.000 175.950 757.050 176.550 ;
        RECT 763.950 175.950 766.050 178.050 ;
        RECT 767.100 174.900 768.150 179.100 ;
        RECT 769.950 177.450 772.050 178.050 ;
        RECT 776.550 177.450 777.450 179.550 ;
        RECT 784.950 178.950 787.050 179.550 ;
        RECT 769.950 176.550 777.450 177.450 ;
        RECT 769.950 175.950 772.050 176.550 ;
        RECT 782.100 176.100 783.900 176.850 ;
        RECT 701.700 171.600 704.400 172.650 ;
        RECT 719.700 171.600 722.400 172.650 ;
        RECT 653.400 159.600 655.200 165.600 ;
        RECT 668.400 159.600 670.200 165.600 ;
        RECT 683.700 159.600 685.500 171.600 ;
        RECT 702.600 159.600 704.400 171.600 ;
        RECT 720.600 159.600 722.400 171.600 ;
        RECT 737.400 165.600 738.600 174.900 ;
        RECT 749.400 165.600 750.600 174.900 ;
        RECT 766.950 171.600 768.150 174.900 ;
        RECT 781.950 172.950 784.050 175.050 ;
        RECT 737.400 159.600 739.200 165.600 ;
        RECT 748.800 159.600 750.600 165.600 ;
        RECT 766.500 159.600 768.300 171.600 ;
        RECT 785.400 165.600 786.600 177.900 ;
        RECT 788.100 176.100 789.900 176.850 ;
        RECT 787.950 169.950 790.050 175.050 ;
        RECT 792.150 173.700 793.050 188.400 ;
        RECT 800.550 187.800 802.350 189.600 ;
        RECT 803.850 188.550 808.800 189.600 ;
        RECT 816.300 190.500 817.350 191.400 ;
        RECT 816.300 189.300 820.050 190.500 ;
        RECT 803.850 187.800 805.650 188.550 ;
        RECT 817.950 188.400 820.050 189.300 ;
        RECT 823.650 188.400 825.450 194.400 ;
        RECT 800.850 184.800 801.900 187.800 ;
        RECT 795.000 183.600 812.850 184.800 ;
        RECT 824.250 184.050 825.450 188.400 ;
        RECT 795.000 182.850 795.900 183.600 ;
        RECT 800.100 183.000 801.900 183.600 ;
        RECT 811.050 183.000 812.850 183.600 ;
        RECT 794.100 181.050 795.900 182.850 ;
        RECT 811.050 182.100 811.950 183.000 ;
        RECT 819.150 182.250 819.900 184.050 ;
        RECT 820.950 181.950 823.050 184.050 ;
        RECT 824.100 181.950 825.450 184.050 ;
        RECT 797.100 178.800 798.900 179.400 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 797.100 177.600 801.900 178.800 ;
        RECT 802.950 175.950 805.050 178.050 ;
        RECT 801.450 173.700 803.250 174.000 ;
        RECT 792.150 173.100 803.250 173.700 ;
        RECT 792.150 172.500 809.850 173.100 ;
        RECT 792.150 171.600 793.050 172.500 ;
        RECT 801.450 172.200 809.850 172.500 ;
        RECT 784.800 159.600 786.600 165.600 ;
        RECT 792.150 159.600 793.950 171.600 ;
        RECT 806.250 170.700 808.050 171.300 ;
        RECT 800.550 169.500 808.050 170.700 ;
        RECT 808.950 170.100 809.850 172.200 ;
        RECT 811.050 172.200 811.950 177.900 ;
        RECT 821.250 173.400 823.050 175.200 ;
        RECT 817.950 172.200 822.150 173.400 ;
        RECT 811.050 171.300 817.050 172.200 ;
        RECT 817.950 171.300 820.050 172.200 ;
        RECT 824.250 171.600 825.450 181.950 ;
        RECT 816.150 170.400 817.050 171.300 ;
        RECT 813.450 170.100 815.250 170.400 ;
        RECT 800.550 168.600 801.750 169.500 ;
        RECT 808.950 169.200 815.250 170.100 ;
        RECT 813.450 168.600 815.250 169.200 ;
        RECT 816.150 168.600 818.850 170.400 ;
        RECT 796.950 166.500 801.750 168.600 ;
        RECT 804.450 167.550 806.250 168.300 ;
        RECT 809.250 167.550 811.050 168.300 ;
        RECT 804.450 166.500 811.050 167.550 ;
        RECT 800.550 165.600 801.750 166.500 ;
        RECT 800.550 159.600 802.350 165.600 ;
        RECT 808.350 159.600 810.150 166.500 ;
        RECT 816.150 165.600 820.050 167.700 ;
        RECT 816.150 159.600 817.950 165.600 ;
        RECT 823.650 159.600 825.450 171.600 ;
        RECT 3.150 143.400 4.950 155.400 ;
        RECT 11.550 149.400 13.350 155.400 ;
        RECT 11.550 148.500 12.750 149.400 ;
        RECT 19.350 148.500 21.150 155.400 ;
        RECT 27.150 149.400 28.950 155.400 ;
        RECT 7.950 146.400 12.750 148.500 ;
        RECT 15.450 147.450 22.050 148.500 ;
        RECT 15.450 146.700 17.250 147.450 ;
        RECT 20.250 146.700 22.050 147.450 ;
        RECT 27.150 147.300 31.050 149.400 ;
        RECT 11.550 145.500 12.750 146.400 ;
        RECT 24.450 145.800 26.250 146.400 ;
        RECT 11.550 144.300 19.050 145.500 ;
        RECT 17.250 143.700 19.050 144.300 ;
        RECT 19.950 144.900 26.250 145.800 ;
        RECT 3.150 142.500 4.050 143.400 ;
        RECT 19.950 142.800 20.850 144.900 ;
        RECT 24.450 144.600 26.250 144.900 ;
        RECT 27.150 144.600 29.850 146.400 ;
        RECT 27.150 143.700 28.050 144.600 ;
        RECT 12.450 142.500 20.850 142.800 ;
        RECT 3.150 141.900 20.850 142.500 ;
        RECT 22.050 142.800 28.050 143.700 ;
        RECT 28.950 142.800 31.050 143.700 ;
        RECT 34.650 143.400 36.450 155.400 ;
        RECT 3.150 141.300 14.250 141.900 ;
        RECT 3.150 126.600 4.050 141.300 ;
        RECT 12.450 141.000 14.250 141.300 ;
        RECT 8.100 136.200 12.900 137.400 ;
        RECT 13.950 136.950 19.050 139.050 ;
        RECT 22.050 137.100 22.950 142.800 ;
        RECT 28.950 141.600 33.150 142.800 ;
        RECT 32.250 139.800 34.050 141.600 ;
        RECT 8.100 135.600 9.900 136.200 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 5.100 132.150 6.900 133.950 ;
        RECT 35.250 133.050 36.450 143.400 ;
        RECT 45.600 143.400 47.400 155.400 ;
        RECT 59.400 149.400 61.200 155.400 ;
        RECT 45.600 142.350 48.300 143.400 ;
        RECT 44.100 137.100 45.900 137.850 ;
        RECT 46.950 137.100 48.300 142.350 ;
        RECT 50.100 140.100 51.900 140.850 ;
        RECT 59.400 140.100 60.600 149.400 ;
        RECT 73.500 143.400 75.300 155.400 ;
        RECT 93.600 143.400 95.400 155.400 ;
        RECT 112.500 143.400 114.300 155.400 ;
        RECT 130.800 149.400 132.600 155.400 ;
        RECT 73.950 140.100 75.150 143.400 ;
        RECT 93.600 142.350 96.300 143.400 ;
        RECT 37.950 135.450 42.000 136.050 ;
        RECT 43.950 135.450 46.050 136.050 ;
        RECT 37.950 134.550 46.050 135.450 ;
        RECT 37.950 133.950 42.000 134.550 ;
        RECT 43.950 133.950 46.050 134.550 ;
        RECT 6.000 131.400 6.900 132.150 ;
        RECT 22.050 132.000 22.950 132.900 ;
        RECT 11.100 131.400 12.900 132.000 ;
        RECT 22.050 131.400 23.850 132.000 ;
        RECT 6.000 130.200 23.850 131.400 ;
        RECT 30.150 130.950 30.900 132.750 ;
        RECT 31.950 130.950 34.050 133.050 ;
        RECT 35.100 130.950 36.450 133.050 ;
        RECT 47.100 132.900 48.300 137.100 ;
        RECT 49.950 138.450 52.050 139.050 ;
        RECT 54.000 138.450 58.050 139.050 ;
        RECT 49.950 137.550 58.050 138.450 ;
        RECT 49.950 136.950 52.050 137.550 ;
        RECT 54.000 136.950 58.050 137.550 ;
        RECT 58.950 136.950 61.050 139.050 ;
        RECT 70.950 136.800 73.050 139.050 ;
        RECT 74.100 135.900 75.150 140.100 ;
        RECT 76.950 136.950 79.050 139.050 ;
        RECT 92.100 137.100 93.900 137.850 ;
        RECT 94.950 137.100 96.300 142.350 ;
        RECT 98.100 140.100 99.900 140.850 ;
        RECT 112.950 140.100 114.150 143.400 ;
        RECT 56.100 134.100 57.900 134.850 ;
        RECT 46.950 131.100 48.300 132.900 ;
        RECT 55.950 130.950 58.050 133.050 ;
        RECT 11.850 127.200 12.900 130.200 ;
        RECT 3.150 120.600 4.950 126.600 ;
        RECT 7.950 124.500 10.050 126.600 ;
        RECT 11.550 125.400 13.350 127.200 ;
        RECT 14.850 126.450 16.650 127.200 ;
        RECT 35.250 126.600 36.450 130.950 ;
        RECT 37.950 129.450 40.050 130.050 ;
        RECT 46.950 129.450 49.050 130.050 ;
        RECT 37.950 128.550 49.050 129.450 ;
        RECT 37.950 127.950 40.050 128.550 ;
        RECT 46.950 127.950 49.050 128.550 ;
        RECT 14.850 125.400 19.800 126.450 ;
        RECT 28.950 125.700 31.050 126.600 ;
        RECT 9.000 123.600 10.050 124.500 ;
        RECT 18.750 123.600 19.800 125.400 ;
        RECT 27.300 124.500 31.050 125.700 ;
        RECT 27.300 123.600 28.350 124.500 ;
        RECT 9.000 122.700 12.750 123.600 ;
        RECT 10.950 120.600 12.750 122.700 ;
        RECT 18.750 120.600 20.550 123.600 ;
        RECT 26.550 120.600 28.350 123.600 ;
        RECT 34.650 120.600 36.450 126.600 ;
        RECT 47.400 123.600 48.600 126.900 ;
        RECT 46.800 120.600 48.600 123.600 ;
        RECT 59.400 123.600 60.600 135.900 ;
        RECT 71.100 135.150 72.900 135.900 ;
        RECT 68.100 134.100 69.900 134.850 ;
        RECT 73.950 134.100 75.150 135.900 ;
        RECT 77.100 135.150 78.900 135.900 ;
        RECT 91.950 133.950 94.050 136.050 ;
        RECT 67.950 130.950 70.050 133.050 ;
        RECT 73.950 130.950 76.050 133.050 ;
        RECT 95.100 132.900 96.300 137.100 ;
        RECT 97.950 136.950 100.050 139.050 ;
        RECT 109.950 136.950 112.050 139.050 ;
        RECT 113.100 135.900 114.150 140.100 ;
        RECT 127.950 139.950 130.050 142.050 ;
        RECT 115.950 136.950 118.050 139.050 ;
        RECT 128.100 138.150 129.900 138.900 ;
        RECT 131.400 137.100 132.600 149.400 ;
        RECT 144.600 143.400 146.400 155.400 ;
        RECT 160.800 149.400 162.600 155.400 ;
        RECT 175.800 149.400 177.600 155.400 ;
        RECT 144.600 142.350 147.300 143.400 ;
        RECT 133.950 139.950 136.050 142.050 ;
        RECT 134.100 138.150 135.900 138.900 ;
        RECT 143.100 137.100 144.900 137.850 ;
        RECT 145.950 137.100 147.300 142.350 ;
        RECT 149.100 140.100 150.900 140.850 ;
        RECT 157.950 139.950 160.050 142.050 ;
        RECT 110.100 135.150 111.900 135.900 ;
        RECT 107.100 134.100 108.900 134.850 ;
        RECT 112.950 134.100 114.150 135.900 ;
        RECT 116.100 135.150 117.900 135.900 ;
        RECT 121.950 135.450 124.050 136.050 ;
        RECT 130.950 135.450 133.050 136.050 ;
        RECT 121.950 134.550 133.050 135.450 ;
        RECT 121.950 133.950 124.050 134.550 ;
        RECT 130.950 133.950 133.050 134.550 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 94.950 131.100 96.300 132.900 ;
        RECT 106.950 130.950 109.050 133.050 ;
        RECT 112.950 130.950 115.050 133.050 ;
        RECT 146.100 132.900 147.300 137.100 ;
        RECT 148.950 136.950 154.050 139.050 ;
        RECT 158.100 138.150 159.900 138.900 ;
        RECT 161.400 137.100 162.600 149.400 ;
        RECT 163.950 139.950 166.050 142.050 ;
        RECT 176.400 140.100 177.600 149.400 ;
        RECT 193.500 143.400 195.300 155.400 ;
        RECT 215.700 143.400 217.500 155.400 ;
        RECT 232.800 149.400 234.600 155.400 ;
        RECT 193.950 140.100 195.150 143.400 ;
        RECT 164.100 138.150 165.900 138.900 ;
        RECT 175.950 136.950 178.050 139.050 ;
        RECT 190.950 136.950 193.050 139.050 ;
        RECT 160.950 133.950 163.050 136.050 ;
        RECT 194.100 135.900 195.150 140.100 ;
        RECT 215.850 140.100 217.050 143.400 ;
        RECT 233.400 140.100 234.600 149.400 ;
        RECT 245.400 149.400 247.200 155.400 ;
        RECT 260.400 149.400 262.200 155.400 ;
        RECT 278.400 149.400 280.200 155.400 ;
        RECT 196.950 136.950 199.050 139.050 ;
        RECT 211.950 136.950 214.050 139.050 ;
        RECT 215.850 135.900 216.900 140.100 ;
        RECT 241.950 139.950 244.050 142.050 ;
        RECT 217.950 136.950 220.050 139.050 ;
        RECT 223.950 138.450 226.050 139.050 ;
        RECT 232.950 138.450 235.050 139.050 ;
        RECT 223.950 137.550 235.050 138.450 ;
        RECT 242.100 138.150 243.900 138.900 ;
        RECT 223.950 136.950 226.050 137.550 ;
        RECT 232.950 136.950 235.050 137.550 ;
        RECT 245.400 137.100 246.600 149.400 ;
        RECT 247.950 139.950 250.050 142.050 ;
        RECT 256.950 139.950 259.050 142.050 ;
        RECT 248.100 138.150 249.900 138.900 ;
        RECT 257.100 138.150 258.900 138.900 ;
        RECT 260.400 137.100 261.600 149.400 ;
        RECT 262.950 139.950 265.050 142.050 ;
        RECT 274.950 139.950 277.050 142.050 ;
        RECT 263.100 138.150 264.900 138.900 ;
        RECT 275.100 138.150 276.900 138.900 ;
        RECT 278.400 137.100 279.600 149.400 ;
        RECT 293.400 143.400 295.200 155.400 ;
        RECT 300.900 144.900 302.700 155.400 ;
        RECT 300.900 143.400 303.300 144.900 ;
        RECT 316.800 143.400 318.600 155.400 ;
        RECT 319.800 144.300 321.600 155.400 ;
        RECT 325.800 144.300 327.600 155.400 ;
        RECT 319.800 143.400 327.600 144.300 ;
        RECT 335.400 149.400 337.200 155.400 ;
        RECT 353.400 149.400 355.200 155.400 ;
        RECT 293.400 142.200 294.600 143.400 ;
        RECT 280.950 139.950 283.050 142.050 ;
        RECT 293.400 141.000 300.600 142.200 ;
        RECT 298.800 140.400 300.600 141.000 ;
        RECT 281.100 138.150 282.900 138.900 ;
        RECT 292.950 136.950 295.050 139.050 ;
        RECT 74.850 129.750 76.050 129.900 ;
        RECT 74.850 128.700 78.600 129.750 ;
        RECT 68.400 125.700 76.200 127.050 ;
        RECT 59.400 120.600 61.200 123.600 ;
        RECT 68.400 120.600 70.200 125.700 ;
        RECT 74.400 120.600 76.200 125.700 ;
        RECT 77.400 126.600 78.600 128.700 ;
        RECT 88.950 129.450 93.000 130.050 ;
        RECT 94.950 129.450 97.050 130.050 ;
        RECT 88.950 128.550 97.050 129.450 ;
        RECT 113.850 129.750 115.050 129.900 ;
        RECT 113.850 128.700 117.600 129.750 ;
        RECT 131.400 128.700 132.600 132.900 ;
        RECT 145.950 131.100 147.300 132.900 ;
        RECT 88.950 127.950 93.000 128.550 ;
        RECT 94.950 127.950 97.050 128.550 ;
        RECT 77.400 120.600 79.200 126.600 ;
        RECT 95.400 123.600 96.600 126.900 ;
        RECT 94.800 120.600 96.600 123.600 ;
        RECT 107.400 125.700 115.200 127.050 ;
        RECT 107.400 120.600 109.200 125.700 ;
        RECT 113.400 120.600 115.200 125.700 ;
        RECT 116.400 126.600 117.600 128.700 ;
        RECT 129.000 127.800 132.600 128.700 ;
        RECT 133.950 129.450 136.050 130.050 ;
        RECT 145.950 129.450 148.050 130.050 ;
        RECT 133.950 128.550 148.050 129.450 ;
        RECT 161.400 128.700 162.600 132.900 ;
        RECT 133.950 127.950 136.050 128.550 ;
        RECT 145.950 127.950 148.050 128.550 ;
        RECT 159.000 127.800 162.600 128.700 ;
        RECT 116.400 120.600 118.200 126.600 ;
        RECT 129.000 120.600 130.800 127.800 ;
        RECT 146.400 123.600 147.600 126.900 ;
        RECT 145.800 120.600 147.600 123.600 ;
        RECT 159.000 120.600 160.800 127.800 ;
        RECT 176.400 123.600 177.600 135.900 ;
        RECT 191.100 135.150 192.900 135.900 ;
        RECT 179.100 134.100 180.900 134.850 ;
        RECT 188.100 134.100 189.900 134.850 ;
        RECT 193.950 134.100 195.150 135.900 ;
        RECT 197.100 135.150 198.900 135.900 ;
        RECT 212.100 135.150 213.900 135.900 ;
        RECT 215.850 134.100 217.050 135.900 ;
        RECT 218.100 135.150 219.900 135.900 ;
        RECT 221.100 134.100 222.900 134.850 ;
        RECT 178.950 130.950 181.050 133.050 ;
        RECT 187.950 130.950 190.050 133.050 ;
        RECT 193.950 130.950 196.050 133.050 ;
        RECT 214.950 130.950 217.050 133.050 ;
        RECT 220.950 130.950 223.050 133.050 ;
        RECT 194.850 129.750 196.050 129.900 ;
        RECT 214.950 129.750 216.150 129.900 ;
        RECT 194.850 128.700 198.600 129.750 ;
        RECT 175.800 120.600 177.600 123.600 ;
        RECT 188.400 125.700 196.200 127.050 ;
        RECT 188.400 120.600 190.200 125.700 ;
        RECT 194.400 120.600 196.200 125.700 ;
        RECT 197.400 126.600 198.600 128.700 ;
        RECT 212.400 128.700 216.150 129.750 ;
        RECT 212.400 126.600 213.600 128.700 ;
        RECT 197.400 120.600 199.200 126.600 ;
        RECT 211.800 120.600 213.600 126.600 ;
        RECT 214.800 125.700 222.600 127.050 ;
        RECT 214.800 120.600 216.600 125.700 ;
        RECT 220.800 120.600 222.600 125.700 ;
        RECT 233.400 123.600 234.600 135.900 ;
        RECT 236.100 134.100 237.900 134.850 ;
        RECT 241.950 133.950 247.050 136.050 ;
        RECT 259.950 135.450 262.050 136.050 ;
        RECT 271.950 135.450 274.050 136.050 ;
        RECT 259.950 134.550 274.050 135.450 ;
        RECT 259.950 133.950 262.050 134.550 ;
        RECT 271.950 133.950 274.050 134.550 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 293.100 135.150 294.900 135.900 ;
        RECT 296.100 134.100 297.900 134.850 ;
        RECT 235.950 130.950 238.050 133.050 ;
        RECT 245.400 128.700 246.600 132.900 ;
        RECT 260.400 128.700 261.600 132.900 ;
        RECT 278.400 128.700 279.600 132.900 ;
        RECT 295.950 130.950 298.050 133.050 ;
        RECT 299.700 129.600 300.600 140.400 ;
        RECT 301.950 137.100 303.300 143.400 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 317.400 134.100 318.300 143.400 ;
        RECT 331.950 139.950 334.050 142.050 ;
        RECT 319.950 136.950 322.050 139.050 ;
        RECT 325.950 136.950 328.050 139.050 ;
        RECT 332.100 138.150 333.900 138.900 ;
        RECT 335.400 137.100 336.600 149.400 ;
        RECT 337.950 139.950 340.050 142.050 ;
        RECT 349.950 139.950 352.050 142.050 ;
        RECT 338.100 138.150 339.900 138.900 ;
        RECT 350.100 138.150 351.900 138.900 ;
        RECT 353.400 137.100 354.600 149.400 ;
        RECT 373.500 143.400 375.300 155.400 ;
        RECT 391.800 149.400 393.600 155.400 ;
        RECT 355.950 139.950 358.050 142.050 ;
        RECT 373.950 140.100 375.150 143.400 ;
        RECT 356.100 138.150 357.900 138.900 ;
        RECT 370.950 136.950 373.050 139.050 ;
        RECT 320.100 135.150 321.900 135.900 ;
        RECT 326.100 135.150 327.900 135.900 ;
        RECT 334.950 135.450 337.050 136.050 ;
        RECT 346.950 135.450 349.050 136.050 ;
        RECT 323.100 134.100 324.900 134.850 ;
        RECT 334.950 134.550 349.050 135.450 ;
        RECT 334.950 133.950 337.050 134.550 ;
        RECT 346.950 133.950 349.050 134.550 ;
        RECT 352.950 135.450 355.050 136.050 ;
        RECT 361.950 135.450 364.050 136.050 ;
        RECT 374.100 135.900 375.150 140.100 ;
        RECT 388.950 139.950 391.050 142.050 ;
        RECT 376.950 136.950 379.050 139.050 ;
        RECT 389.100 138.150 390.900 138.900 ;
        RECT 392.400 137.100 393.600 149.400 ;
        RECT 394.950 139.950 397.050 145.050 ;
        RECT 399.150 143.400 400.950 155.400 ;
        RECT 407.550 149.400 409.350 155.400 ;
        RECT 407.550 148.500 408.750 149.400 ;
        RECT 415.350 148.500 417.150 155.400 ;
        RECT 423.150 149.400 424.950 155.400 ;
        RECT 403.950 146.400 408.750 148.500 ;
        RECT 411.450 147.450 418.050 148.500 ;
        RECT 411.450 146.700 413.250 147.450 ;
        RECT 416.250 146.700 418.050 147.450 ;
        RECT 423.150 147.300 427.050 149.400 ;
        RECT 407.550 145.500 408.750 146.400 ;
        RECT 420.450 145.800 422.250 146.400 ;
        RECT 407.550 144.300 415.050 145.500 ;
        RECT 413.250 143.700 415.050 144.300 ;
        RECT 415.950 144.900 422.250 145.800 ;
        RECT 399.150 142.500 400.050 143.400 ;
        RECT 415.950 142.800 416.850 144.900 ;
        RECT 420.450 144.600 422.250 144.900 ;
        RECT 423.150 144.600 425.850 146.400 ;
        RECT 423.150 143.700 424.050 144.600 ;
        RECT 408.450 142.500 416.850 142.800 ;
        RECT 399.150 141.900 416.850 142.500 ;
        RECT 418.050 142.800 424.050 143.700 ;
        RECT 424.950 142.800 427.050 143.700 ;
        RECT 430.650 143.400 432.450 155.400 ;
        RECT 440.400 144.600 442.200 155.400 ;
        RECT 446.400 154.500 454.200 155.400 ;
        RECT 446.400 144.600 448.200 154.500 ;
        RECT 440.400 143.700 448.200 144.600 ;
        RECT 399.150 141.300 410.250 141.900 ;
        RECT 395.100 138.150 396.900 138.900 ;
        RECT 352.950 134.550 364.050 135.450 ;
        RECT 371.100 135.150 372.900 135.900 ;
        RECT 352.950 133.950 355.050 134.550 ;
        RECT 361.950 133.950 364.050 134.550 ;
        RECT 368.100 134.100 369.900 134.850 ;
        RECT 373.950 134.100 375.150 135.900 ;
        RECT 377.100 135.150 378.900 135.900 ;
        RECT 382.950 135.450 385.050 136.050 ;
        RECT 391.950 135.450 394.050 136.050 ;
        RECT 382.950 134.550 394.050 135.450 ;
        RECT 382.950 133.950 385.050 134.550 ;
        RECT 391.950 133.950 394.050 134.550 ;
        RECT 298.950 128.700 300.750 129.600 ;
        RECT 245.400 127.800 249.000 128.700 ;
        RECT 260.400 127.800 264.000 128.700 ;
        RECT 278.400 127.800 282.000 128.700 ;
        RECT 232.800 120.600 234.600 123.600 ;
        RECT 247.200 120.600 249.000 127.800 ;
        RECT 262.200 120.600 264.000 127.800 ;
        RECT 280.200 120.600 282.000 127.800 ;
        RECT 297.300 127.800 300.750 128.700 ;
        RECT 297.300 123.600 298.200 127.800 ;
        RECT 303.000 126.600 304.050 132.900 ;
        RECT 307.950 132.450 310.050 133.050 ;
        RECT 316.950 132.450 319.050 133.050 ;
        RECT 307.950 131.550 319.050 132.450 ;
        RECT 307.950 130.950 310.050 131.550 ;
        RECT 316.950 130.950 319.050 131.550 ;
        RECT 322.950 130.950 325.050 133.050 ;
        RECT 317.400 126.600 318.300 129.900 ;
        RECT 335.400 128.700 336.600 132.900 ;
        RECT 353.400 128.700 354.600 132.900 ;
        RECT 367.950 130.950 370.050 133.050 ;
        RECT 373.950 132.450 376.050 133.050 ;
        RECT 385.950 132.450 388.050 133.050 ;
        RECT 373.950 131.550 388.050 132.450 ;
        RECT 373.950 130.950 376.050 131.550 ;
        RECT 385.950 130.950 388.050 131.550 ;
        RECT 374.850 129.750 376.050 129.900 ;
        RECT 374.850 128.700 378.600 129.750 ;
        RECT 392.400 128.700 393.600 132.900 ;
        RECT 335.400 127.800 339.000 128.700 ;
        RECT 353.400 127.800 357.000 128.700 ;
        RECT 296.400 120.600 298.200 123.600 ;
        RECT 302.400 120.600 304.200 126.600 ;
        RECT 317.400 124.950 322.800 126.600 ;
        RECT 321.000 120.600 322.800 124.950 ;
        RECT 337.200 120.600 339.000 127.800 ;
        RECT 355.200 120.600 357.000 127.800 ;
        RECT 368.400 125.700 376.200 127.050 ;
        RECT 368.400 120.600 370.200 125.700 ;
        RECT 374.400 120.600 376.200 125.700 ;
        RECT 377.400 126.600 378.600 128.700 ;
        RECT 390.000 127.800 393.600 128.700 ;
        RECT 377.400 120.600 379.200 126.600 ;
        RECT 390.000 120.600 391.800 127.800 ;
        RECT 399.150 126.600 400.050 141.300 ;
        RECT 408.450 141.000 410.250 141.300 ;
        RECT 404.100 136.200 408.900 137.400 ;
        RECT 409.950 136.950 412.050 139.200 ;
        RECT 418.050 137.100 418.950 142.800 ;
        RECT 424.950 141.600 429.150 142.800 ;
        RECT 428.250 139.800 430.050 141.600 ;
        RECT 404.100 135.600 405.900 136.200 ;
        RECT 415.950 133.950 418.050 136.050 ;
        RECT 401.100 132.150 402.900 133.950 ;
        RECT 431.250 133.050 432.450 143.400 ;
        RECT 449.400 142.500 451.200 153.600 ;
        RECT 452.400 143.400 454.200 154.500 ;
        RECT 464.400 149.400 466.200 155.400 ;
        RECT 447.150 141.600 451.200 142.500 ;
        RECT 464.400 142.500 465.600 149.400 ;
        RECT 470.700 143.400 472.500 155.400 ;
        RECT 485.700 143.400 487.500 155.400 ;
        RECT 494.550 143.400 496.350 155.400 ;
        RECT 502.050 149.400 503.850 155.400 ;
        RECT 499.950 147.300 503.850 149.400 ;
        RECT 509.850 148.500 511.650 155.400 ;
        RECT 517.650 149.400 519.450 155.400 ;
        RECT 518.250 148.500 519.450 149.400 ;
        RECT 508.950 147.450 515.550 148.500 ;
        RECT 508.950 146.700 510.750 147.450 ;
        RECT 513.750 146.700 515.550 147.450 ;
        RECT 518.250 146.400 523.050 148.500 ;
        RECT 501.150 144.600 503.850 146.400 ;
        RECT 504.750 145.800 506.550 146.400 ;
        RECT 504.750 144.900 511.050 145.800 ;
        RECT 518.250 145.500 519.450 146.400 ;
        RECT 504.750 144.600 506.550 144.900 ;
        RECT 502.950 143.700 503.850 144.600 ;
        RECT 464.400 141.600 470.100 142.500 ;
        RECT 447.150 140.100 448.050 141.600 ;
        RECT 468.150 140.700 470.100 141.600 ;
        RECT 435.000 138.450 439.050 139.050 ;
        RECT 402.000 131.400 402.900 132.150 ;
        RECT 418.050 132.000 418.950 132.900 ;
        RECT 407.100 131.400 408.900 132.000 ;
        RECT 418.050 131.400 419.850 132.000 ;
        RECT 402.000 130.200 419.850 131.400 ;
        RECT 426.150 130.950 426.900 132.750 ;
        RECT 427.950 130.950 430.050 133.050 ;
        RECT 431.100 130.950 432.450 133.050 ;
        RECT 407.850 127.200 408.900 130.200 ;
        RECT 399.150 120.600 400.950 126.600 ;
        RECT 403.950 124.500 406.050 126.600 ;
        RECT 407.550 125.400 409.350 127.200 ;
        RECT 410.850 126.450 412.650 127.200 ;
        RECT 431.250 126.600 432.450 130.950 ;
        RECT 434.550 136.950 439.050 138.450 ;
        RECT 442.950 136.950 445.050 139.050 ;
        RECT 434.550 129.900 435.450 136.950 ;
        RECT 447.150 135.900 447.900 140.100 ;
        RECT 448.950 136.950 451.050 139.050 ;
        RECT 464.100 137.100 465.900 137.850 ;
        RECT 443.250 135.150 445.050 135.900 ;
        RECT 440.250 134.100 442.050 134.850 ;
        RECT 447.150 134.100 448.050 135.900 ;
        RECT 448.950 135.150 450.750 135.900 ;
        RECT 452.100 134.100 453.900 134.850 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 468.150 134.100 469.050 140.700 ;
        RECT 471.000 134.100 472.200 143.400 ;
        RECT 485.850 140.100 487.050 143.400 ;
        RECT 481.950 136.950 484.050 139.050 ;
        RECT 485.850 135.900 486.900 140.100 ;
        RECT 487.950 136.950 490.050 139.050 ;
        RECT 482.100 135.150 483.900 135.900 ;
        RECT 485.850 134.100 487.050 135.900 ;
        RECT 488.100 135.150 489.900 135.900 ;
        RECT 491.100 134.100 492.900 134.850 ;
        RECT 439.950 130.950 442.050 133.050 ;
        RECT 445.950 130.950 448.050 133.050 ;
        RECT 451.950 130.950 454.050 133.050 ;
        RECT 468.150 129.900 468.900 134.100 ;
        RECT 494.550 133.050 495.750 143.400 ;
        RECT 499.950 142.800 502.050 143.700 ;
        RECT 502.950 142.800 508.950 143.700 ;
        RECT 497.850 141.600 502.050 142.800 ;
        RECT 496.950 139.800 498.750 141.600 ;
        RECT 508.050 137.100 508.950 142.800 ;
        RECT 510.150 142.800 511.050 144.900 ;
        RECT 511.950 144.300 519.450 145.500 ;
        RECT 511.950 143.700 513.750 144.300 ;
        RECT 526.050 143.400 527.850 155.400 ;
        RECT 537.600 143.400 539.400 155.400 ;
        RECT 510.150 142.500 518.550 142.800 ;
        RECT 526.950 142.500 527.850 143.400 ;
        RECT 510.150 141.900 527.850 142.500 ;
        RECT 516.750 141.300 527.850 141.900 ;
        RECT 516.750 141.000 518.550 141.300 ;
        RECT 511.950 136.950 517.050 139.050 ;
        RECT 518.100 136.200 522.900 137.400 ;
        RECT 508.950 133.950 511.050 136.050 ;
        RECT 521.100 135.600 522.900 136.200 ;
        RECT 469.950 130.950 475.050 133.050 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 490.950 130.950 493.050 133.050 ;
        RECT 494.550 130.950 495.900 133.050 ;
        RECT 496.950 130.950 499.050 133.050 ;
        RECT 500.100 130.950 500.850 132.750 ;
        RECT 508.050 132.000 508.950 132.900 ;
        RECT 524.100 132.150 525.900 133.950 ;
        RECT 507.150 131.400 508.950 132.000 ;
        RECT 518.100 131.400 519.900 132.000 ;
        RECT 524.100 131.400 525.000 132.150 ;
        RECT 433.950 127.800 436.050 129.900 ;
        RECT 445.950 126.600 447.000 129.900 ;
        RECT 468.150 129.300 469.050 129.900 ;
        RECT 468.150 128.400 470.100 129.300 ;
        RECT 410.850 125.400 415.800 126.450 ;
        RECT 424.950 125.700 427.050 126.600 ;
        RECT 405.000 123.600 406.050 124.500 ;
        RECT 414.750 123.600 415.800 125.400 ;
        RECT 423.300 124.500 427.050 125.700 ;
        RECT 423.300 123.600 424.350 124.500 ;
        RECT 405.000 122.700 408.750 123.600 ;
        RECT 406.950 120.600 408.750 122.700 ;
        RECT 414.750 120.600 416.550 123.600 ;
        RECT 422.550 120.600 424.350 123.600 ;
        RECT 430.650 120.600 432.450 126.600 ;
        RECT 445.200 120.600 447.000 126.600 ;
        RECT 465.000 127.500 470.100 128.400 ;
        RECT 465.000 123.600 466.200 127.500 ;
        RECT 471.000 126.600 472.200 129.900 ;
        RECT 484.950 129.750 486.150 129.900 ;
        RECT 482.400 128.700 486.150 129.750 ;
        RECT 482.400 126.600 483.600 128.700 ;
        RECT 464.400 120.600 466.200 123.600 ;
        RECT 470.700 120.600 472.500 126.600 ;
        RECT 481.800 120.600 483.600 126.600 ;
        RECT 484.800 125.700 492.600 127.050 ;
        RECT 484.800 120.600 486.600 125.700 ;
        RECT 490.800 120.600 492.600 125.700 ;
        RECT 494.550 126.600 495.750 130.950 ;
        RECT 507.150 130.200 525.000 131.400 ;
        RECT 518.100 127.200 519.150 130.200 ;
        RECT 494.550 120.600 496.350 126.600 ;
        RECT 499.950 125.700 502.050 126.600 ;
        RECT 514.350 126.450 516.150 127.200 ;
        RECT 499.950 124.500 503.700 125.700 ;
        RECT 502.650 123.600 503.700 124.500 ;
        RECT 511.200 125.400 516.150 126.450 ;
        RECT 517.650 125.400 519.450 127.200 ;
        RECT 526.950 126.600 527.850 141.300 ;
        RECT 536.700 142.350 539.400 143.400 ;
        RECT 545.550 143.400 547.350 155.400 ;
        RECT 553.050 149.400 554.850 155.400 ;
        RECT 550.950 147.300 554.850 149.400 ;
        RECT 560.850 148.500 562.650 155.400 ;
        RECT 568.650 149.400 570.450 155.400 ;
        RECT 569.250 148.500 570.450 149.400 ;
        RECT 559.950 147.450 566.550 148.500 ;
        RECT 559.950 146.700 561.750 147.450 ;
        RECT 564.750 146.700 566.550 147.450 ;
        RECT 569.250 146.400 574.050 148.500 ;
        RECT 552.150 144.600 554.850 146.400 ;
        RECT 555.750 145.800 557.550 146.400 ;
        RECT 555.750 144.900 562.050 145.800 ;
        RECT 569.250 145.500 570.450 146.400 ;
        RECT 555.750 144.600 557.550 144.900 ;
        RECT 553.950 143.700 554.850 144.600 ;
        RECT 533.100 140.100 534.900 140.850 ;
        RECT 532.950 136.950 535.050 139.050 ;
        RECT 536.700 137.100 538.050 142.350 ;
        RECT 539.100 137.100 540.900 137.850 ;
        RECT 529.950 129.450 532.050 133.050 ;
        RECT 536.700 132.900 537.900 137.100 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 545.550 133.050 546.750 143.400 ;
        RECT 550.950 142.800 553.050 143.700 ;
        RECT 553.950 142.800 559.950 143.700 ;
        RECT 548.850 141.600 553.050 142.800 ;
        RECT 547.950 139.800 549.750 141.600 ;
        RECT 559.050 137.100 559.950 142.800 ;
        RECT 561.150 142.800 562.050 144.900 ;
        RECT 562.950 144.300 570.450 145.500 ;
        RECT 562.950 143.700 564.750 144.300 ;
        RECT 577.050 143.400 578.850 155.400 ;
        RECT 586.800 143.400 588.600 155.400 ;
        RECT 589.800 144.300 591.600 155.400 ;
        RECT 595.800 144.300 597.600 155.400 ;
        RECT 609.300 144.900 611.100 155.400 ;
        RECT 589.800 143.400 597.600 144.300 ;
        RECT 608.700 143.400 611.100 144.900 ;
        RECT 616.800 143.400 618.600 155.400 ;
        RECT 561.150 142.500 569.550 142.800 ;
        RECT 577.950 142.500 578.850 143.400 ;
        RECT 561.150 141.900 578.850 142.500 ;
        RECT 567.750 141.300 578.850 141.900 ;
        RECT 567.750 141.000 569.550 141.300 ;
        RECT 565.950 136.950 568.050 139.050 ;
        RECT 569.100 136.200 573.900 137.400 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 572.100 135.600 573.900 136.200 ;
        RECT 536.700 131.100 538.050 132.900 ;
        RECT 545.550 130.950 546.900 133.050 ;
        RECT 547.950 130.950 550.050 133.050 ;
        RECT 551.100 130.950 551.850 132.750 ;
        RECT 559.050 132.000 559.950 132.900 ;
        RECT 575.100 132.150 576.900 133.950 ;
        RECT 558.150 131.400 559.950 132.000 ;
        RECT 569.100 131.400 570.900 132.000 ;
        RECT 575.100 131.400 576.000 132.150 ;
        RECT 535.950 129.450 538.050 130.050 ;
        RECT 529.950 129.000 538.050 129.450 ;
        RECT 530.550 128.550 538.050 129.000 ;
        RECT 535.950 127.950 538.050 128.550 ;
        RECT 511.200 123.600 512.250 125.400 ;
        RECT 520.950 124.500 523.050 126.600 ;
        RECT 520.950 123.600 522.000 124.500 ;
        RECT 502.650 120.600 504.450 123.600 ;
        RECT 510.450 120.600 512.250 123.600 ;
        RECT 518.250 122.700 522.000 123.600 ;
        RECT 518.250 120.600 520.050 122.700 ;
        RECT 526.050 120.600 527.850 126.600 ;
        RECT 536.400 123.600 537.600 126.900 ;
        RECT 545.550 126.600 546.750 130.950 ;
        RECT 558.150 130.200 576.000 131.400 ;
        RECT 569.100 127.200 570.150 130.200 ;
        RECT 536.400 120.600 538.200 123.600 ;
        RECT 545.550 120.600 547.350 126.600 ;
        RECT 550.950 125.700 553.050 126.600 ;
        RECT 565.350 126.450 567.150 127.200 ;
        RECT 550.950 124.500 554.700 125.700 ;
        RECT 553.650 123.600 554.700 124.500 ;
        RECT 562.200 125.400 567.150 126.450 ;
        RECT 568.650 125.400 570.450 127.200 ;
        RECT 577.950 126.600 578.850 141.300 ;
        RECT 587.400 134.100 588.300 143.400 ;
        RECT 589.950 136.950 592.050 139.050 ;
        RECT 595.950 136.950 598.050 139.050 ;
        RECT 608.700 137.100 610.050 143.400 ;
        RECT 617.400 142.200 618.600 143.400 ;
        RECT 611.400 141.000 618.600 142.200 ;
        RECT 629.400 149.400 631.200 155.400 ;
        RECT 644.400 149.400 646.200 155.400 ;
        RECT 611.400 140.400 613.200 141.000 ;
        RECT 590.100 135.150 591.900 135.900 ;
        RECT 596.100 135.150 597.900 135.900 ;
        RECT 601.950 135.450 606.000 136.050 ;
        RECT 607.950 135.450 610.050 136.050 ;
        RECT 593.100 134.100 594.900 134.850 ;
        RECT 601.950 134.550 610.050 135.450 ;
        RECT 601.950 133.950 606.000 134.550 ;
        RECT 607.950 133.950 610.050 134.550 ;
        RECT 583.950 130.950 589.050 133.050 ;
        RECT 592.950 130.950 595.050 133.050 ;
        RECT 562.200 123.600 563.250 125.400 ;
        RECT 571.950 124.500 574.050 126.600 ;
        RECT 571.950 123.600 573.000 124.500 ;
        RECT 553.650 120.600 555.450 123.600 ;
        RECT 561.450 120.600 563.250 123.600 ;
        RECT 569.250 122.700 573.000 123.600 ;
        RECT 569.250 120.600 571.050 122.700 ;
        RECT 577.050 120.600 578.850 126.600 ;
        RECT 587.400 126.600 588.300 129.900 ;
        RECT 607.950 126.600 609.000 132.900 ;
        RECT 611.400 129.600 612.300 140.400 ;
        RECT 629.400 140.100 630.600 149.400 ;
        RECT 640.950 139.950 643.050 142.050 ;
        RECT 616.950 136.950 619.050 139.050 ;
        RECT 622.950 138.450 627.000 139.050 ;
        RECT 628.950 138.450 631.050 139.050 ;
        RECT 622.950 137.550 631.050 138.450 ;
        RECT 641.100 138.150 642.900 138.900 ;
        RECT 622.950 136.950 627.000 137.550 ;
        RECT 628.950 136.950 631.050 137.550 ;
        RECT 644.400 137.100 645.600 149.400 ;
        RECT 653.550 143.400 655.350 155.400 ;
        RECT 661.050 149.400 662.850 155.400 ;
        RECT 658.950 147.300 662.850 149.400 ;
        RECT 668.850 148.500 670.650 155.400 ;
        RECT 676.650 149.400 678.450 155.400 ;
        RECT 677.250 148.500 678.450 149.400 ;
        RECT 667.950 147.450 674.550 148.500 ;
        RECT 667.950 146.700 669.750 147.450 ;
        RECT 672.750 146.700 674.550 147.450 ;
        RECT 677.250 146.400 682.050 148.500 ;
        RECT 660.150 144.600 662.850 146.400 ;
        RECT 663.750 145.800 665.550 146.400 ;
        RECT 663.750 144.900 670.050 145.800 ;
        RECT 677.250 145.500 678.450 146.400 ;
        RECT 663.750 144.600 665.550 144.900 ;
        RECT 661.950 143.700 662.850 144.600 ;
        RECT 646.950 139.950 649.050 142.050 ;
        RECT 647.100 138.150 648.900 138.900 ;
        RECT 617.100 135.150 618.900 135.900 ;
        RECT 614.100 134.100 615.900 134.850 ;
        RECT 626.100 134.100 627.900 134.850 ;
        RECT 613.950 130.950 616.050 133.050 ;
        RECT 611.250 128.700 613.050 129.600 ;
        RECT 611.250 127.800 614.700 128.700 ;
        RECT 587.400 124.950 592.800 126.600 ;
        RECT 591.000 120.600 592.800 124.950 ;
        RECT 607.800 120.600 609.600 126.600 ;
        RECT 613.800 123.600 614.700 127.800 ;
        RECT 629.400 123.600 630.600 135.900 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 653.550 133.050 654.750 143.400 ;
        RECT 658.950 142.800 661.050 143.700 ;
        RECT 661.950 142.800 667.950 143.700 ;
        RECT 656.850 141.600 661.050 142.800 ;
        RECT 655.950 139.800 657.750 141.600 ;
        RECT 667.050 137.100 667.950 142.800 ;
        RECT 669.150 142.800 670.050 144.900 ;
        RECT 670.950 144.300 678.450 145.500 ;
        RECT 670.950 143.700 672.750 144.300 ;
        RECT 685.050 143.400 686.850 155.400 ;
        RECT 669.150 142.500 677.550 142.800 ;
        RECT 685.950 142.500 686.850 143.400 ;
        RECT 669.150 141.900 686.850 142.500 ;
        RECT 695.400 149.400 697.200 155.400 ;
        RECT 675.750 141.300 686.850 141.900 ;
        RECT 675.750 141.000 677.550 141.300 ;
        RECT 673.950 136.950 676.050 139.050 ;
        RECT 677.100 136.200 681.900 137.400 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 680.100 135.600 681.900 136.200 ;
        RECT 644.400 128.700 645.600 132.900 ;
        RECT 653.550 130.950 654.900 133.050 ;
        RECT 655.950 130.950 658.050 133.050 ;
        RECT 659.100 130.950 659.850 132.750 ;
        RECT 667.050 132.000 667.950 132.900 ;
        RECT 683.100 132.150 684.900 133.950 ;
        RECT 666.150 131.400 667.950 132.000 ;
        RECT 677.100 131.400 678.900 132.000 ;
        RECT 683.100 131.400 684.000 132.150 ;
        RECT 644.400 127.800 648.000 128.700 ;
        RECT 613.800 120.600 615.600 123.600 ;
        RECT 629.400 120.600 631.200 123.600 ;
        RECT 646.200 120.600 648.000 127.800 ;
        RECT 653.550 126.600 654.750 130.950 ;
        RECT 666.150 130.200 684.000 131.400 ;
        RECT 677.100 127.200 678.150 130.200 ;
        RECT 653.550 120.600 655.350 126.600 ;
        RECT 658.950 125.700 661.050 126.600 ;
        RECT 673.350 126.450 675.150 127.200 ;
        RECT 658.950 124.500 662.700 125.700 ;
        RECT 661.650 123.600 662.700 124.500 ;
        RECT 670.200 125.400 675.150 126.450 ;
        RECT 676.650 125.400 678.450 127.200 ;
        RECT 685.950 126.600 686.850 141.300 ;
        RECT 688.950 139.950 694.050 142.050 ;
        RECT 692.100 138.150 693.900 138.900 ;
        RECT 695.400 137.100 696.600 149.400 ;
        RECT 716.700 143.400 718.500 155.400 ;
        RECT 734.700 143.400 736.500 155.400 ;
        RECT 749.400 144.300 751.200 155.400 ;
        RECT 755.400 144.300 757.200 155.400 ;
        RECT 749.400 143.400 757.200 144.300 ;
        RECT 758.400 143.400 760.200 155.400 ;
        RECT 773.700 143.400 775.500 155.400 ;
        RECT 789.600 143.400 791.400 155.400 ;
        RECT 697.950 139.950 700.050 142.050 ;
        RECT 716.850 140.100 718.050 143.400 ;
        RECT 734.850 140.100 736.050 143.400 ;
        RECT 698.100 138.150 699.900 138.900 ;
        RECT 712.950 136.950 715.050 139.050 ;
        RECT 694.950 135.450 697.050 136.050 ;
        RECT 706.950 135.450 709.050 136.200 ;
        RECT 716.850 135.900 717.900 140.100 ;
        RECT 718.950 136.950 721.050 139.050 ;
        RECT 730.950 136.950 733.050 139.050 ;
        RECT 734.850 135.900 735.900 140.100 ;
        RECT 736.950 136.950 739.050 139.050 ;
        RECT 748.950 136.950 751.050 139.050 ;
        RECT 754.950 136.950 757.050 139.050 ;
        RECT 694.950 134.550 709.050 135.450 ;
        RECT 713.100 135.150 714.900 135.900 ;
        RECT 694.950 133.950 697.050 134.550 ;
        RECT 706.950 134.100 709.050 134.550 ;
        RECT 716.850 134.100 718.050 135.900 ;
        RECT 719.100 135.150 720.900 135.900 ;
        RECT 731.100 135.150 732.900 135.900 ;
        RECT 722.100 134.100 723.900 134.850 ;
        RECT 734.850 134.100 736.050 135.900 ;
        RECT 737.100 135.150 738.900 135.900 ;
        RECT 749.100 135.150 750.900 135.900 ;
        RECT 755.100 135.150 756.900 135.900 ;
        RECT 740.100 134.100 741.900 134.850 ;
        RECT 752.100 134.100 753.900 134.850 ;
        RECT 758.700 134.100 759.600 143.400 ;
        RECT 773.850 140.100 775.050 143.400 ;
        RECT 788.700 142.350 791.400 143.400 ;
        RECT 806.400 149.400 808.200 155.400 ;
        RECT 818.400 149.400 820.200 155.400 ;
        RECT 785.100 140.100 786.900 140.850 ;
        RECT 769.950 136.950 772.050 139.050 ;
        RECT 773.850 135.900 774.900 140.100 ;
        RECT 775.950 136.950 778.050 139.050 ;
        RECT 784.950 136.950 787.050 139.050 ;
        RECT 788.700 137.100 790.050 142.350 ;
        RECT 793.950 141.450 798.000 142.050 ;
        RECT 793.950 139.950 798.450 141.450 ;
        RECT 806.400 140.100 807.600 149.400 ;
        RECT 814.950 139.950 817.050 142.050 ;
        RECT 797.550 138.450 798.450 139.950 ;
        RECT 805.950 138.450 808.050 139.050 ;
        RECT 791.100 137.100 792.900 137.850 ;
        RECT 797.550 137.550 808.050 138.450 ;
        RECT 815.100 138.150 816.900 138.900 ;
        RECT 770.100 135.150 771.900 135.900 ;
        RECT 773.850 134.100 775.050 135.900 ;
        RECT 776.100 135.150 777.900 135.900 ;
        RECT 779.100 134.100 780.900 134.850 ;
        RECT 695.400 128.700 696.600 132.900 ;
        RECT 706.950 132.450 709.050 132.900 ;
        RECT 715.950 132.450 718.050 133.050 ;
        RECT 706.950 131.550 718.050 132.450 ;
        RECT 706.950 130.800 709.050 131.550 ;
        RECT 715.950 130.950 718.050 131.550 ;
        RECT 721.950 130.950 724.050 133.050 ;
        RECT 730.950 130.950 736.050 133.050 ;
        RECT 739.950 130.950 742.050 133.050 ;
        RECT 751.950 130.950 754.050 133.050 ;
        RECT 757.950 130.950 760.050 133.050 ;
        RECT 768.000 132.900 771.000 133.050 ;
        RECT 766.950 132.450 771.000 132.900 ;
        RECT 772.950 132.450 775.050 133.050 ;
        RECT 766.950 131.550 775.050 132.450 ;
        RECT 766.950 130.950 771.000 131.550 ;
        RECT 772.950 130.950 775.050 131.550 ;
        RECT 778.950 130.950 781.050 133.050 ;
        RECT 788.700 132.900 789.900 137.100 ;
        RECT 805.950 136.950 808.050 137.550 ;
        RECT 818.400 137.100 819.600 149.400 ;
        RECT 820.950 139.950 823.050 142.050 ;
        RECT 821.100 138.150 822.900 138.900 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 803.100 134.100 804.900 134.850 ;
        RECT 788.700 131.100 790.050 132.900 ;
        RECT 802.950 130.950 805.050 133.050 ;
        RECT 766.950 130.800 769.050 130.950 ;
        RECT 715.950 129.750 717.150 129.900 ;
        RECT 733.950 129.750 735.150 129.900 ;
        RECT 713.400 128.700 717.150 129.750 ;
        RECT 731.400 128.700 735.150 129.750 ;
        RECT 695.400 127.800 699.000 128.700 ;
        RECT 670.200 123.600 671.250 125.400 ;
        RECT 679.950 124.500 682.050 126.600 ;
        RECT 679.950 123.600 681.000 124.500 ;
        RECT 661.650 120.600 663.450 123.600 ;
        RECT 669.450 120.600 671.250 123.600 ;
        RECT 677.250 122.700 681.000 123.600 ;
        RECT 677.250 120.600 679.050 122.700 ;
        RECT 685.050 120.600 686.850 126.600 ;
        RECT 697.200 120.600 699.000 127.800 ;
        RECT 713.400 126.600 714.600 128.700 ;
        RECT 712.800 120.600 714.600 126.600 ;
        RECT 715.800 125.700 723.600 127.050 ;
        RECT 731.400 126.600 732.600 128.700 ;
        RECT 715.800 120.600 717.600 125.700 ;
        RECT 721.800 120.600 723.600 125.700 ;
        RECT 730.800 120.600 732.600 126.600 ;
        RECT 733.800 125.700 741.600 127.050 ;
        RECT 758.700 126.600 759.600 129.900 ;
        RECT 772.950 129.750 774.150 129.900 ;
        RECT 770.400 128.700 774.150 129.750 ;
        RECT 784.950 129.450 790.050 130.050 ;
        RECT 770.400 126.600 771.600 128.700 ;
        RECT 784.950 128.550 798.450 129.450 ;
        RECT 784.950 127.950 790.050 128.550 ;
        RECT 733.800 120.600 735.600 125.700 ;
        RECT 739.800 120.600 741.600 125.700 ;
        RECT 754.200 124.950 759.600 126.600 ;
        RECT 754.200 120.600 756.000 124.950 ;
        RECT 769.800 120.600 771.600 126.600 ;
        RECT 772.800 125.700 780.600 127.050 ;
        RECT 772.800 120.600 774.600 125.700 ;
        RECT 778.800 120.600 780.600 125.700 ;
        RECT 788.400 123.600 789.600 126.900 ;
        RECT 797.550 126.450 798.450 128.550 ;
        RECT 802.950 126.450 805.050 127.050 ;
        RECT 797.550 125.550 805.050 126.450 ;
        RECT 802.950 124.950 805.050 125.550 ;
        RECT 806.400 123.600 807.600 135.900 ;
        RECT 811.950 135.450 816.000 136.050 ;
        RECT 817.950 135.450 820.050 136.050 ;
        RECT 811.950 134.550 820.050 135.450 ;
        RECT 811.950 133.950 816.000 134.550 ;
        RECT 817.950 133.950 820.050 134.550 ;
        RECT 818.400 128.700 819.600 132.900 ;
        RECT 818.400 127.800 822.000 128.700 ;
        RECT 788.400 120.600 790.200 123.600 ;
        RECT 806.400 120.600 808.200 123.600 ;
        RECT 820.200 120.600 822.000 127.800 ;
        RECT 13.800 113.400 15.600 116.400 ;
        RECT 14.400 110.100 15.600 113.400 ;
        RECT 29.400 113.400 31.200 116.400 ;
        RECT 29.400 110.100 30.600 113.400 ;
        RECT 48.000 112.050 49.800 116.400 ;
        RECT 65.400 113.400 67.200 116.400 ;
        RECT 44.400 110.400 49.800 112.050 ;
        RECT 13.950 108.450 16.050 109.050 ;
        RECT 22.950 108.450 25.050 109.050 ;
        RECT 13.950 107.550 25.050 108.450 ;
        RECT 13.950 106.950 16.050 107.550 ;
        RECT 22.950 106.950 25.050 107.550 ;
        RECT 28.950 108.450 31.050 109.050 ;
        RECT 37.950 108.450 40.050 108.900 ;
        RECT 28.950 107.550 40.050 108.450 ;
        RECT 28.950 106.950 31.050 107.550 ;
        RECT 37.950 106.800 40.050 107.550 ;
        RECT 44.400 107.100 45.300 110.400 ;
        RECT 66.300 109.200 67.200 113.400 ;
        RECT 71.400 110.400 73.200 116.400 ;
        RECT 66.300 108.300 69.750 109.200 ;
        RECT 67.950 107.400 69.750 108.300 ;
        RECT 13.950 104.100 15.300 105.900 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 14.100 99.900 15.300 104.100 ;
        RECT 29.700 104.100 31.050 105.900 ;
        RECT 11.100 99.150 12.900 99.900 ;
        RECT 13.950 94.650 15.300 99.900 ;
        RECT 16.950 97.950 19.050 103.050 ;
        RECT 25.950 97.950 28.050 100.050 ;
        RECT 29.700 99.900 30.900 104.100 ;
        RECT 40.950 103.950 46.050 106.050 ;
        RECT 49.950 103.950 52.050 106.050 ;
        RECT 64.950 103.950 67.050 106.050 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 17.100 96.150 18.900 96.900 ;
        RECT 26.100 96.150 27.900 96.900 ;
        RECT 12.600 93.600 15.300 94.650 ;
        RECT 29.700 94.650 31.050 99.900 ;
        RECT 32.100 99.150 33.900 99.900 ;
        RECT 29.700 93.600 32.400 94.650 ;
        RECT 44.400 93.600 45.300 102.900 ;
        RECT 50.100 102.150 51.900 102.900 ;
        RECT 65.100 102.150 66.900 102.900 ;
        RECT 47.100 101.100 48.900 101.850 ;
        RECT 53.100 101.100 54.900 101.850 ;
        RECT 62.100 101.100 63.900 101.850 ;
        RECT 46.950 97.950 49.050 100.050 ;
        RECT 52.950 97.950 55.050 100.050 ;
        RECT 61.950 97.950 64.050 100.050 ;
        RECT 68.700 96.600 69.600 107.400 ;
        RECT 72.000 104.100 73.050 110.400 ;
        RECT 85.200 109.200 87.000 116.400 ;
        RECT 100.200 109.200 102.000 116.400 ;
        RECT 115.200 109.200 117.000 116.400 ;
        RECT 130.800 110.400 132.600 116.400 ;
        RECT 83.400 108.300 87.000 109.200 ;
        RECT 98.400 108.300 102.000 109.200 ;
        RECT 113.400 108.300 117.000 109.200 ;
        RECT 131.400 108.300 132.600 110.400 ;
        RECT 133.800 111.300 135.600 116.400 ;
        RECT 139.800 111.300 141.600 116.400 ;
        RECT 133.800 109.950 141.600 111.300 ;
        RECT 152.400 113.400 154.200 116.400 ;
        RECT 83.400 104.100 84.600 108.300 ;
        RECT 98.400 104.100 99.600 108.300 ;
        RECT 113.400 104.100 114.600 108.300 ;
        RECT 131.400 107.250 135.150 108.300 ;
        RECT 133.950 107.100 135.150 107.250 ;
        RECT 133.950 103.950 136.050 106.050 ;
        RECT 139.950 103.950 142.050 106.050 ;
        RECT 148.950 103.950 151.050 106.050 ;
        RECT 70.950 102.450 73.050 103.050 ;
        RECT 75.000 102.450 79.050 103.050 ;
        RECT 70.950 101.550 79.050 102.450 ;
        RECT 70.950 100.950 73.050 101.550 ;
        RECT 75.000 100.950 79.050 101.550 ;
        RECT 82.950 102.450 85.050 103.050 ;
        RECT 91.950 102.450 94.050 103.050 ;
        RECT 82.950 101.550 94.050 102.450 ;
        RECT 82.950 100.950 85.050 101.550 ;
        RECT 91.950 100.950 94.050 101.550 ;
        RECT 97.950 102.450 100.050 103.050 ;
        RECT 102.000 102.450 106.050 103.050 ;
        RECT 97.950 101.550 106.050 102.450 ;
        RECT 97.950 100.950 100.050 101.550 ;
        RECT 102.000 100.950 106.050 101.550 ;
        RECT 112.950 102.450 115.050 103.050 ;
        RECT 124.950 102.450 127.050 103.050 ;
        RECT 112.950 101.550 127.050 102.450 ;
        RECT 112.950 100.950 115.050 101.550 ;
        RECT 124.950 100.950 127.050 101.550 ;
        RECT 131.100 101.100 132.900 101.850 ;
        RECT 134.850 101.100 136.050 102.900 ;
        RECT 140.100 102.150 141.900 102.900 ;
        RECT 149.100 102.150 150.900 102.900 ;
        RECT 137.100 101.100 138.900 101.850 ;
        RECT 152.400 101.100 153.600 113.400 ;
        RECT 168.000 109.200 169.800 116.400 ;
        RECT 176.550 110.400 178.350 116.400 ;
        RECT 184.650 113.400 186.450 116.400 ;
        RECT 192.450 113.400 194.250 116.400 ;
        RECT 200.250 114.300 202.050 116.400 ;
        RECT 200.250 113.400 204.000 114.300 ;
        RECT 184.650 112.500 185.700 113.400 ;
        RECT 181.950 111.300 185.700 112.500 ;
        RECT 193.200 111.600 194.250 113.400 ;
        RECT 202.950 112.500 204.000 113.400 ;
        RECT 181.950 110.400 184.050 111.300 ;
        RECT 193.200 110.550 198.150 111.600 ;
        RECT 168.000 108.300 171.600 109.200 ;
        RECT 170.400 104.100 171.600 108.300 ;
        RECT 176.550 106.050 177.750 110.400 ;
        RECT 196.350 109.800 198.150 110.550 ;
        RECT 199.650 109.800 201.450 111.600 ;
        RECT 202.950 110.400 205.050 112.500 ;
        RECT 208.050 110.400 209.850 116.400 ;
        RECT 176.550 103.950 177.900 106.050 ;
        RECT 178.950 103.950 181.050 109.050 ;
        RECT 200.100 106.800 201.150 109.800 ;
        RECT 182.100 104.250 182.850 106.050 ;
        RECT 189.150 105.600 207.000 106.800 ;
        RECT 189.150 105.000 190.950 105.600 ;
        RECT 200.100 105.000 201.900 105.600 ;
        RECT 190.050 104.100 190.950 105.000 ;
        RECT 206.100 104.850 207.000 105.600 ;
        RECT 172.950 103.050 175.050 103.200 ;
        RECT 169.950 101.100 175.050 103.050 ;
        RECT 67.800 96.000 69.600 96.600 ;
        RECT 62.400 94.800 69.600 96.000 ;
        RECT 62.400 93.600 63.600 94.800 ;
        RECT 70.950 93.600 72.300 99.900 ;
        RECT 80.100 98.100 81.900 98.850 ;
        RECT 79.950 94.950 82.050 97.050 ;
        RECT 12.600 81.600 14.400 93.600 ;
        RECT 30.600 81.600 32.400 93.600 ;
        RECT 43.800 81.600 45.600 93.600 ;
        RECT 46.800 92.700 54.600 93.600 ;
        RECT 46.800 81.600 48.600 92.700 ;
        RECT 52.800 81.600 54.600 92.700 ;
        RECT 62.400 81.600 64.200 93.600 ;
        RECT 69.900 92.100 72.300 93.600 ;
        RECT 69.900 81.600 71.700 92.100 ;
        RECT 83.400 87.600 84.600 99.900 ;
        RECT 86.100 98.100 87.900 98.850 ;
        RECT 95.100 98.100 96.900 98.850 ;
        RECT 85.950 94.950 88.050 97.050 ;
        RECT 94.950 94.950 97.050 97.050 ;
        RECT 98.400 87.600 99.600 99.900 ;
        RECT 101.100 98.100 102.900 98.850 ;
        RECT 110.100 98.100 111.900 98.850 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 109.950 94.950 112.050 97.050 ;
        RECT 113.400 87.600 114.600 99.900 ;
        RECT 116.100 98.100 117.900 98.850 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 115.950 94.950 118.050 97.050 ;
        RECT 134.850 96.900 135.900 101.100 ;
        RECT 169.950 100.950 174.450 101.100 ;
        RECT 136.950 97.950 139.050 100.050 ;
        RECT 151.950 99.450 154.050 100.050 ;
        RECT 156.000 99.450 160.050 100.050 ;
        RECT 151.950 98.550 160.050 99.450 ;
        RECT 151.950 97.950 154.050 98.550 ;
        RECT 156.000 97.950 160.050 98.550 ;
        RECT 167.100 98.100 168.900 98.850 ;
        RECT 134.850 93.600 136.050 96.900 ;
        RECT 83.400 81.600 85.200 87.600 ;
        RECT 98.400 81.600 100.200 87.600 ;
        RECT 113.400 81.600 115.200 87.600 ;
        RECT 134.700 81.600 136.500 93.600 ;
        RECT 152.400 87.600 153.600 96.900 ;
        RECT 166.950 94.950 169.050 97.050 ;
        RECT 170.400 87.600 171.600 99.900 ;
        RECT 173.100 98.100 174.900 98.850 ;
        RECT 172.950 94.950 175.050 97.050 ;
        RECT 152.400 81.600 154.200 87.600 ;
        RECT 169.800 81.600 171.600 87.600 ;
        RECT 176.550 93.600 177.750 103.950 ;
        RECT 206.100 103.050 207.900 104.850 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 178.950 95.400 180.750 97.200 ;
        RECT 179.850 94.200 184.050 95.400 ;
        RECT 190.050 94.200 190.950 99.900 ;
        RECT 196.950 97.950 199.050 103.050 ;
        RECT 203.100 100.800 204.900 101.400 ;
        RECT 200.100 99.600 204.900 100.800 ;
        RECT 198.750 95.700 200.550 96.000 ;
        RECT 208.950 95.700 209.850 110.400 ;
        RECT 215.400 108.600 217.200 116.400 ;
        RECT 222.900 112.200 224.700 116.400 ;
        RECT 222.900 110.400 224.850 112.200 ;
        RECT 221.100 108.600 222.900 109.500 ;
        RECT 215.400 107.700 222.900 108.600 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 215.100 99.150 216.900 99.900 ;
        RECT 198.750 95.100 209.850 95.700 ;
        RECT 176.550 81.600 178.350 93.600 ;
        RECT 181.950 93.300 184.050 94.200 ;
        RECT 184.950 93.300 190.950 94.200 ;
        RECT 192.150 94.500 209.850 95.100 ;
        RECT 192.150 94.200 200.550 94.500 ;
        RECT 184.950 92.400 185.850 93.300 ;
        RECT 183.150 90.600 185.850 92.400 ;
        RECT 186.750 92.100 188.550 92.400 ;
        RECT 192.150 92.100 193.050 94.200 ;
        RECT 208.950 93.600 209.850 94.500 ;
        RECT 186.750 91.200 193.050 92.100 ;
        RECT 193.950 92.700 195.750 93.300 ;
        RECT 193.950 91.500 201.450 92.700 ;
        RECT 186.750 90.600 188.550 91.200 ;
        RECT 200.250 90.600 201.450 91.500 ;
        RECT 181.950 87.600 185.850 89.700 ;
        RECT 190.950 89.550 192.750 90.300 ;
        RECT 195.750 89.550 197.550 90.300 ;
        RECT 190.950 88.500 197.550 89.550 ;
        RECT 200.250 88.500 205.050 90.600 ;
        RECT 184.050 81.600 185.850 87.600 ;
        RECT 191.850 81.600 193.650 88.500 ;
        RECT 200.250 87.600 201.450 88.500 ;
        RECT 199.650 81.600 201.450 87.600 ;
        RECT 208.050 81.600 209.850 93.600 ;
        RECT 218.400 87.600 219.450 107.700 ;
        RECT 223.950 107.100 224.850 110.400 ;
        RECT 233.400 111.300 235.200 116.400 ;
        RECT 239.400 111.300 241.200 116.400 ;
        RECT 233.400 109.950 241.200 111.300 ;
        RECT 242.400 110.400 244.200 116.400 ;
        RECT 242.400 108.300 243.600 110.400 ;
        RECT 256.200 109.200 258.000 116.400 ;
        RECT 268.500 110.400 270.300 116.400 ;
        RECT 274.800 113.400 276.600 116.400 ;
        RECT 239.850 107.250 243.600 108.300 ;
        RECT 254.400 108.300 258.000 109.200 ;
        RECT 239.850 107.100 241.050 107.250 ;
        RECT 223.950 103.950 229.050 106.050 ;
        RECT 232.950 103.950 235.050 106.050 ;
        RECT 238.950 105.450 241.050 106.050 ;
        RECT 243.000 105.450 247.050 106.050 ;
        RECT 238.950 104.550 247.050 105.450 ;
        RECT 238.950 103.950 241.050 104.550 ;
        RECT 243.000 103.950 247.050 104.550 ;
        RECT 254.400 104.100 255.600 108.300 ;
        RECT 268.800 107.100 270.000 110.400 ;
        RECT 274.800 109.500 276.000 113.400 ;
        RECT 288.300 112.200 290.100 116.400 ;
        RECT 270.900 108.600 276.000 109.500 ;
        RECT 288.150 110.400 290.100 112.200 ;
        RECT 270.900 107.700 272.850 108.600 ;
        RECT 271.950 107.100 272.850 107.700 ;
        RECT 288.150 107.100 289.050 110.400 ;
        RECT 290.100 108.600 291.900 109.500 ;
        RECT 295.800 108.600 297.600 116.400 ;
        RECT 305.400 113.400 307.200 116.400 ;
        RECT 305.400 110.100 306.600 113.400 ;
        RECT 320.400 111.300 322.200 116.400 ;
        RECT 326.400 111.300 328.200 116.400 ;
        RECT 320.400 109.950 328.200 111.300 ;
        RECT 329.400 110.400 331.200 116.400 ;
        RECT 343.500 110.400 345.300 116.400 ;
        RECT 349.800 113.400 351.600 116.400 ;
        RECT 290.100 107.700 297.600 108.600 ;
        RECT 304.950 108.450 307.050 109.050 ;
        RECT 313.950 108.450 316.050 109.050 ;
        RECT 259.950 105.450 262.050 106.050 ;
        RECT 268.950 105.450 271.050 106.050 ;
        RECT 259.950 104.550 271.050 105.450 ;
        RECT 259.950 103.950 262.050 104.550 ;
        RECT 268.950 103.950 271.050 104.550 ;
        RECT 221.100 101.100 222.900 101.850 ;
        RECT 220.950 97.950 223.050 100.050 ;
        RECT 225.000 93.600 226.050 102.900 ;
        RECT 233.100 102.150 234.900 102.900 ;
        RECT 236.100 101.100 237.900 101.850 ;
        RECT 238.950 101.100 240.150 102.900 ;
        RECT 247.950 102.450 252.000 103.050 ;
        RECT 253.950 102.450 256.050 103.050 ;
        RECT 272.100 102.900 272.850 107.100 ;
        RECT 286.950 103.950 289.050 106.050 ;
        RECT 242.100 101.100 243.900 101.850 ;
        RECT 247.950 101.550 256.050 102.450 ;
        RECT 235.950 97.950 238.050 100.050 ;
        RECT 239.100 96.900 240.150 101.100 ;
        RECT 247.950 100.950 252.000 101.550 ;
        RECT 253.950 100.950 256.050 101.550 ;
        RECT 241.950 97.950 244.050 100.050 ;
        RECT 251.100 98.100 252.900 98.850 ;
        RECT 238.950 93.600 240.150 96.900 ;
        RECT 250.950 94.950 253.050 97.050 ;
        RECT 218.400 81.600 220.200 87.600 ;
        RECT 225.000 81.600 226.800 93.600 ;
        RECT 238.500 81.600 240.300 93.600 ;
        RECT 241.950 90.450 244.050 91.050 ;
        RECT 251.550 90.450 252.450 94.950 ;
        RECT 241.950 89.550 252.450 90.450 ;
        RECT 241.950 88.950 244.050 89.550 ;
        RECT 254.400 87.600 255.600 99.900 ;
        RECT 257.100 98.100 258.900 98.850 ;
        RECT 256.950 94.950 259.050 97.050 ;
        RECT 268.800 93.600 270.000 102.900 ;
        RECT 271.950 96.300 272.850 102.900 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 275.100 99.150 276.900 99.900 ;
        RECT 270.900 95.400 272.850 96.300 ;
        RECT 270.900 94.500 276.600 95.400 ;
        RECT 254.400 81.600 256.200 87.600 ;
        RECT 268.500 81.600 270.300 93.600 ;
        RECT 275.400 87.600 276.600 94.500 ;
        RECT 286.950 93.600 288.000 102.900 ;
        RECT 290.100 101.100 291.900 101.850 ;
        RECT 289.950 97.950 292.050 100.050 ;
        RECT 274.800 81.600 276.600 87.600 ;
        RECT 286.200 81.600 288.000 93.600 ;
        RECT 293.550 87.600 294.600 107.700 ;
        RECT 304.950 107.550 316.050 108.450 ;
        RECT 329.400 108.300 330.600 110.400 ;
        RECT 304.950 106.950 307.050 107.550 ;
        RECT 313.950 106.950 316.050 107.550 ;
        RECT 326.850 107.250 330.600 108.300 ;
        RECT 326.850 107.100 328.050 107.250 ;
        RECT 343.800 107.100 345.000 110.400 ;
        RECT 349.800 109.500 351.000 113.400 ;
        RECT 359.400 111.300 361.200 116.400 ;
        RECT 365.400 111.300 367.200 116.400 ;
        RECT 359.400 109.950 367.200 111.300 ;
        RECT 368.400 110.400 370.200 116.400 ;
        RECT 375.150 110.400 376.950 116.400 ;
        RECT 382.950 114.300 384.750 116.400 ;
        RECT 381.000 113.400 384.750 114.300 ;
        RECT 390.750 113.400 392.550 116.400 ;
        RECT 398.550 113.400 400.350 116.400 ;
        RECT 381.000 112.500 382.050 113.400 ;
        RECT 379.950 110.400 382.050 112.500 ;
        RECT 390.750 111.600 391.800 113.400 ;
        RECT 345.900 108.600 351.000 109.500 ;
        RECT 345.900 107.700 347.850 108.600 ;
        RECT 368.400 108.300 369.600 110.400 ;
        RECT 346.950 107.100 347.850 107.700 ;
        RECT 365.850 107.250 369.600 108.300 ;
        RECT 365.850 107.100 367.050 107.250 ;
        RECT 305.700 104.100 307.050 105.900 ;
        RECT 295.950 100.950 298.050 103.050 ;
        RECT 296.100 99.150 297.900 99.900 ;
        RECT 301.950 97.950 304.050 100.050 ;
        RECT 305.700 99.900 306.900 104.100 ;
        RECT 319.950 103.950 322.050 106.050 ;
        RECT 325.950 105.450 328.050 106.050 ;
        RECT 334.950 105.450 337.050 106.050 ;
        RECT 325.950 104.550 337.050 105.450 ;
        RECT 325.950 103.950 328.050 104.550 ;
        RECT 334.950 103.950 337.050 104.550 ;
        RECT 343.950 103.950 346.050 106.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 347.100 102.900 347.850 107.100 ;
        RECT 358.950 103.950 361.050 106.050 ;
        RECT 364.950 103.950 367.050 106.050 ;
        RECT 320.100 102.150 321.900 102.900 ;
        RECT 323.100 101.100 324.900 101.850 ;
        RECT 325.950 101.100 327.150 102.900 ;
        RECT 329.100 101.100 330.900 101.850 ;
        RECT 302.100 96.150 303.900 96.900 ;
        RECT 305.700 94.650 307.050 99.900 ;
        RECT 308.100 99.150 309.900 99.900 ;
        RECT 322.950 97.950 325.050 100.050 ;
        RECT 326.100 96.900 327.150 101.100 ;
        RECT 328.950 97.950 331.050 100.050 ;
        RECT 305.700 93.600 308.400 94.650 ;
        RECT 325.950 93.600 327.150 96.900 ;
        RECT 343.800 93.600 345.000 102.900 ;
        RECT 346.950 96.300 347.850 102.900 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 359.100 102.150 360.900 102.900 ;
        RECT 362.100 101.100 363.900 101.850 ;
        RECT 364.950 101.100 366.150 102.900 ;
        RECT 368.100 101.100 369.900 101.850 ;
        RECT 350.100 99.150 351.900 99.900 ;
        RECT 361.950 97.950 364.050 100.050 ;
        RECT 365.100 96.900 366.150 101.100 ;
        RECT 367.950 97.950 370.050 100.050 ;
        RECT 345.900 95.400 347.850 96.300 ;
        RECT 345.900 94.500 351.600 95.400 ;
        RECT 292.800 81.600 294.600 87.600 ;
        RECT 306.600 81.600 308.400 93.600 ;
        RECT 325.500 81.600 327.300 93.600 ;
        RECT 343.500 81.600 345.300 93.600 ;
        RECT 350.400 87.600 351.600 94.500 ;
        RECT 364.950 93.600 366.150 96.900 ;
        RECT 375.150 95.700 376.050 110.400 ;
        RECT 383.550 109.800 385.350 111.600 ;
        RECT 386.850 110.550 391.800 111.600 ;
        RECT 399.300 112.500 400.350 113.400 ;
        RECT 399.300 111.300 403.050 112.500 ;
        RECT 386.850 109.800 388.650 110.550 ;
        RECT 400.950 110.400 403.050 111.300 ;
        RECT 406.650 110.400 408.450 116.400 ;
        RECT 383.850 106.800 384.900 109.800 ;
        RECT 378.000 105.600 395.850 106.800 ;
        RECT 407.250 106.050 408.450 110.400 ;
        RECT 418.200 109.200 420.000 116.400 ;
        RECT 378.000 104.850 378.900 105.600 ;
        RECT 383.100 105.000 384.900 105.600 ;
        RECT 394.050 105.000 395.850 105.600 ;
        RECT 377.100 103.050 378.900 104.850 ;
        RECT 394.050 104.100 394.950 105.000 ;
        RECT 402.150 104.250 402.900 106.050 ;
        RECT 403.950 103.950 406.050 106.050 ;
        RECT 407.100 103.950 408.450 106.050 ;
        RECT 416.400 108.300 420.000 109.200 ;
        RECT 426.150 110.400 427.950 116.400 ;
        RECT 433.950 114.300 435.750 116.400 ;
        RECT 432.000 113.400 435.750 114.300 ;
        RECT 441.750 113.400 443.550 116.400 ;
        RECT 449.550 113.400 451.350 116.400 ;
        RECT 432.000 112.500 433.050 113.400 ;
        RECT 430.950 110.400 433.050 112.500 ;
        RECT 441.750 111.600 442.800 113.400 ;
        RECT 416.400 104.100 417.600 108.300 ;
        RECT 380.100 100.800 381.900 101.400 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 380.100 99.600 384.900 100.800 ;
        RECT 385.950 97.950 388.050 100.050 ;
        RECT 384.450 95.700 386.250 96.000 ;
        RECT 375.150 95.100 386.250 95.700 ;
        RECT 375.150 94.500 392.850 95.100 ;
        RECT 375.150 93.600 376.050 94.500 ;
        RECT 384.450 94.200 392.850 94.500 ;
        RECT 349.800 81.600 351.600 87.600 ;
        RECT 364.500 81.600 366.300 93.600 ;
        RECT 375.150 81.600 376.950 93.600 ;
        RECT 389.250 92.700 391.050 93.300 ;
        RECT 383.550 91.500 391.050 92.700 ;
        RECT 391.950 92.100 392.850 94.200 ;
        RECT 394.050 94.200 394.950 99.900 ;
        RECT 404.250 95.400 406.050 97.200 ;
        RECT 400.950 94.200 405.150 95.400 ;
        RECT 394.050 93.300 400.050 94.200 ;
        RECT 400.950 93.300 403.050 94.200 ;
        RECT 407.250 93.600 408.450 103.950 ;
        RECT 412.950 103.050 415.050 103.200 ;
        RECT 412.950 101.100 418.050 103.050 ;
        RECT 413.550 100.950 418.050 101.100 ;
        RECT 413.100 98.100 414.900 98.850 ;
        RECT 412.950 94.950 415.050 97.050 ;
        RECT 399.150 92.400 400.050 93.300 ;
        RECT 396.450 92.100 398.250 92.400 ;
        RECT 383.550 90.600 384.750 91.500 ;
        RECT 391.950 91.200 398.250 92.100 ;
        RECT 396.450 90.600 398.250 91.200 ;
        RECT 399.150 90.600 401.850 92.400 ;
        RECT 379.950 88.500 384.750 90.600 ;
        RECT 387.450 89.550 389.250 90.300 ;
        RECT 392.250 89.550 394.050 90.300 ;
        RECT 387.450 88.500 394.050 89.550 ;
        RECT 383.550 87.600 384.750 88.500 ;
        RECT 383.550 81.600 385.350 87.600 ;
        RECT 391.350 81.600 393.150 88.500 ;
        RECT 399.150 87.600 403.050 89.700 ;
        RECT 399.150 81.600 400.950 87.600 ;
        RECT 406.650 81.600 408.450 93.600 ;
        RECT 416.400 87.600 417.600 99.900 ;
        RECT 419.100 98.100 420.900 98.850 ;
        RECT 418.950 94.950 421.050 97.050 ;
        RECT 426.150 95.700 427.050 110.400 ;
        RECT 434.550 109.800 436.350 111.600 ;
        RECT 437.850 110.550 442.800 111.600 ;
        RECT 450.300 112.500 451.350 113.400 ;
        RECT 450.300 111.300 454.050 112.500 ;
        RECT 437.850 109.800 439.650 110.550 ;
        RECT 451.950 110.400 454.050 111.300 ;
        RECT 457.650 110.400 459.450 116.400 ;
        RECT 472.800 113.400 474.600 116.400 ;
        RECT 434.850 106.800 435.900 109.800 ;
        RECT 429.000 105.600 446.850 106.800 ;
        RECT 458.250 106.050 459.450 110.400 ;
        RECT 473.400 110.100 474.600 113.400 ;
        RECT 484.800 110.400 486.600 116.400 ;
        RECT 472.950 106.950 478.050 109.050 ;
        RECT 485.400 108.300 486.600 110.400 ;
        RECT 487.800 111.300 489.600 116.400 ;
        RECT 493.800 111.300 495.600 116.400 ;
        RECT 487.800 109.950 495.600 111.300 ;
        RECT 485.400 107.250 489.150 108.300 ;
        RECT 487.950 107.100 489.150 107.250 ;
        RECT 506.100 108.000 507.900 116.400 ;
        RECT 515.550 110.400 517.350 116.400 ;
        RECT 523.650 113.400 525.450 116.400 ;
        RECT 531.450 113.400 533.250 116.400 ;
        RECT 539.250 114.300 541.050 116.400 ;
        RECT 539.250 113.400 543.000 114.300 ;
        RECT 523.650 112.500 524.700 113.400 ;
        RECT 520.950 111.300 524.700 112.500 ;
        RECT 532.200 111.600 533.250 113.400 ;
        RECT 541.950 112.500 543.000 113.400 ;
        RECT 520.950 110.400 523.050 111.300 ;
        RECT 532.200 110.550 537.150 111.600 ;
        RECT 506.100 106.350 510.300 108.000 ;
        RECT 429.000 104.850 429.900 105.600 ;
        RECT 434.100 105.000 435.900 105.600 ;
        RECT 445.050 105.000 446.850 105.600 ;
        RECT 428.100 103.050 429.900 104.850 ;
        RECT 445.050 104.100 445.950 105.000 ;
        RECT 453.150 104.250 453.900 106.050 ;
        RECT 431.100 100.800 432.900 101.400 ;
        RECT 442.950 100.950 445.050 103.050 ;
        RECT 454.950 100.950 457.050 106.050 ;
        RECT 458.100 103.950 459.450 106.050 ;
        RECT 472.950 104.100 474.300 105.900 ;
        RECT 431.100 99.600 435.900 100.800 ;
        RECT 436.950 97.950 439.050 100.050 ;
        RECT 435.450 95.700 437.250 96.000 ;
        RECT 426.150 95.100 437.250 95.700 ;
        RECT 426.150 94.500 443.850 95.100 ;
        RECT 426.150 93.600 427.050 94.500 ;
        RECT 435.450 94.200 443.850 94.500 ;
        RECT 416.400 81.600 418.200 87.600 ;
        RECT 426.150 81.600 427.950 93.600 ;
        RECT 440.250 92.700 442.050 93.300 ;
        RECT 434.550 91.500 442.050 92.700 ;
        RECT 442.950 92.100 443.850 94.200 ;
        RECT 445.050 94.200 445.950 99.900 ;
        RECT 455.250 95.400 457.050 97.200 ;
        RECT 451.950 94.200 456.150 95.400 ;
        RECT 445.050 93.300 451.050 94.200 ;
        RECT 451.950 93.300 454.050 94.200 ;
        RECT 458.250 93.600 459.450 103.950 ;
        RECT 466.950 100.950 472.050 103.050 ;
        RECT 473.100 99.900 474.300 104.100 ;
        RECT 487.950 103.950 490.050 106.050 ;
        RECT 493.950 103.950 496.050 106.050 ;
        RECT 506.100 104.100 507.900 104.850 ;
        RECT 485.100 101.100 486.900 101.850 ;
        RECT 488.850 101.100 490.050 102.900 ;
        RECT 494.100 102.150 495.900 102.900 ;
        RECT 491.100 101.100 492.900 101.850 ;
        RECT 470.100 99.150 471.900 99.900 ;
        RECT 472.950 94.650 474.300 99.900 ;
        RECT 475.950 97.950 478.050 100.050 ;
        RECT 484.950 97.950 487.050 100.050 ;
        RECT 488.850 96.900 489.900 101.100 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 490.950 97.950 493.050 100.050 ;
        RECT 496.950 99.450 501.000 100.050 ;
        RECT 502.950 99.450 505.050 100.050 ;
        RECT 496.950 98.550 505.050 99.450 ;
        RECT 496.950 97.950 501.000 98.550 ;
        RECT 502.950 97.950 505.050 98.550 ;
        RECT 509.400 98.100 510.300 106.350 ;
        RECT 515.550 106.050 516.750 110.400 ;
        RECT 535.350 109.800 537.150 110.550 ;
        RECT 538.650 109.800 540.450 111.600 ;
        RECT 541.950 110.400 544.050 112.500 ;
        RECT 547.050 110.400 548.850 116.400 ;
        RECT 539.100 106.800 540.150 109.800 ;
        RECT 515.550 103.950 516.900 106.050 ;
        RECT 517.950 103.950 520.050 106.050 ;
        RECT 521.100 104.250 521.850 106.050 ;
        RECT 528.150 105.600 546.000 106.800 ;
        RECT 528.150 105.000 529.950 105.600 ;
        RECT 539.100 105.000 540.900 105.600 ;
        RECT 529.050 104.100 529.950 105.000 ;
        RECT 545.100 104.850 546.000 105.600 ;
        RECT 476.100 96.150 477.900 96.900 ;
        RECT 450.150 92.400 451.050 93.300 ;
        RECT 447.450 92.100 449.250 92.400 ;
        RECT 434.550 90.600 435.750 91.500 ;
        RECT 442.950 91.200 449.250 92.100 ;
        RECT 447.450 90.600 449.250 91.200 ;
        RECT 450.150 90.600 452.850 92.400 ;
        RECT 430.950 88.500 435.750 90.600 ;
        RECT 438.450 89.550 440.250 90.300 ;
        RECT 443.250 89.550 445.050 90.300 ;
        RECT 438.450 88.500 445.050 89.550 ;
        RECT 434.550 87.600 435.750 88.500 ;
        RECT 434.550 81.600 436.350 87.600 ;
        RECT 442.350 81.600 444.150 88.500 ;
        RECT 450.150 87.600 454.050 89.700 ;
        RECT 450.150 81.600 451.950 87.600 ;
        RECT 457.650 81.600 459.450 93.600 ;
        RECT 471.600 93.600 474.300 94.650 ;
        RECT 488.850 93.600 490.050 96.900 ;
        RECT 503.100 96.150 504.900 96.900 ;
        RECT 500.100 95.100 501.900 95.850 ;
        RECT 508.950 94.950 514.050 97.050 ;
        RECT 471.600 81.600 473.400 93.600 ;
        RECT 488.700 81.600 490.500 93.600 ;
        RECT 499.950 91.950 505.050 94.050 ;
        RECT 509.400 88.800 510.300 93.900 ;
        RECT 503.700 87.900 510.300 88.800 ;
        RECT 503.700 87.600 505.200 87.900 ;
        RECT 503.400 81.600 505.200 87.600 ;
        RECT 509.400 87.600 510.300 87.900 ;
        RECT 515.550 93.600 516.750 103.950 ;
        RECT 545.100 103.050 546.900 104.850 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 542.100 100.800 543.900 101.400 ;
        RECT 517.950 95.400 519.750 97.200 ;
        RECT 518.850 94.200 523.050 95.400 ;
        RECT 529.050 94.200 529.950 99.900 ;
        RECT 532.950 97.950 538.050 100.050 ;
        RECT 539.100 99.600 543.900 100.800 ;
        RECT 537.750 95.700 539.550 96.000 ;
        RECT 547.950 95.700 548.850 110.400 ;
        RECT 562.200 109.200 564.000 116.400 ;
        RECT 580.200 110.400 582.000 116.400 ;
        RECT 560.400 108.300 564.000 109.200 ;
        RECT 560.400 104.100 561.600 108.300 ;
        RECT 580.950 107.100 582.000 110.400 ;
        RECT 596.400 111.300 598.200 116.400 ;
        RECT 602.400 111.300 604.200 116.400 ;
        RECT 596.400 109.950 604.200 111.300 ;
        RECT 605.400 110.400 607.200 116.400 ;
        RECT 605.400 108.300 606.600 110.400 ;
        RECT 622.200 109.200 624.000 116.400 ;
        RECT 635.400 111.300 637.200 116.400 ;
        RECT 641.400 111.300 643.200 116.400 ;
        RECT 635.400 109.950 643.200 111.300 ;
        RECT 644.400 110.400 646.200 116.400 ;
        RECT 653.400 113.400 655.200 116.400 ;
        RECT 602.850 107.250 606.600 108.300 ;
        RECT 620.400 108.300 624.000 109.200 ;
        RECT 644.400 108.300 645.600 110.400 ;
        RECT 654.000 109.500 655.200 113.400 ;
        RECT 659.700 110.400 661.500 116.400 ;
        RECT 665.550 110.400 667.350 116.400 ;
        RECT 673.650 113.400 675.450 116.400 ;
        RECT 681.450 113.400 683.250 116.400 ;
        RECT 689.250 114.300 691.050 116.400 ;
        RECT 689.250 113.400 693.000 114.300 ;
        RECT 673.650 112.500 674.700 113.400 ;
        RECT 670.950 111.300 674.700 112.500 ;
        RECT 682.200 111.600 683.250 113.400 ;
        RECT 691.950 112.500 693.000 113.400 ;
        RECT 670.950 110.400 673.050 111.300 ;
        RECT 682.200 110.550 687.150 111.600 ;
        RECT 654.000 108.600 659.100 109.500 ;
        RECT 602.850 107.100 604.050 107.250 ;
        RECT 565.950 105.450 570.000 106.050 ;
        RECT 565.950 105.000 570.450 105.450 ;
        RECT 565.950 103.950 571.050 105.000 ;
        RECT 571.950 103.950 577.050 106.050 ;
        RECT 580.950 103.950 583.050 106.050 ;
        RECT 586.950 103.950 589.050 106.050 ;
        RECT 595.950 103.950 598.050 106.050 ;
        RECT 601.950 105.450 604.050 106.050 ;
        RECT 613.950 105.450 616.050 106.050 ;
        RECT 601.950 104.550 616.050 105.450 ;
        RECT 601.950 103.950 604.050 104.550 ;
        RECT 613.950 103.950 616.050 104.550 ;
        RECT 620.400 104.100 621.600 108.300 ;
        RECT 641.850 107.250 645.600 108.300 ;
        RECT 657.150 107.700 659.100 108.600 ;
        RECT 641.850 107.100 643.050 107.250 ;
        RECT 657.150 107.100 658.050 107.700 ;
        RECT 660.000 107.100 661.200 110.400 ;
        RECT 634.950 103.950 637.050 106.200 ;
        RECT 640.950 103.950 643.050 106.050 ;
        RECT 559.950 100.950 565.050 103.050 ;
        RECT 568.950 100.950 571.050 103.950 ;
        RECT 575.250 102.150 577.050 102.900 ;
        RECT 578.250 101.100 580.050 101.850 ;
        RECT 582.150 101.100 583.050 102.900 ;
        RECT 587.100 102.150 588.900 102.900 ;
        RECT 596.100 102.150 597.900 102.900 ;
        RECT 583.950 101.100 585.750 101.850 ;
        RECT 599.100 101.100 600.900 101.850 ;
        RECT 601.950 101.100 603.150 102.900 ;
        RECT 610.950 102.450 613.050 103.050 ;
        RECT 619.950 102.450 622.050 103.050 ;
        RECT 605.100 101.100 606.900 101.850 ;
        RECT 610.950 101.550 622.050 102.450 ;
        RECT 635.100 102.150 636.900 102.900 ;
        RECT 557.100 98.100 558.900 98.850 ;
        RECT 537.750 95.100 548.850 95.700 ;
        RECT 509.400 81.600 511.200 87.600 ;
        RECT 515.550 81.600 517.350 93.600 ;
        RECT 520.950 93.300 523.050 94.200 ;
        RECT 523.950 93.300 529.950 94.200 ;
        RECT 531.150 94.500 548.850 95.100 ;
        RECT 550.950 96.450 555.000 97.050 ;
        RECT 556.950 96.450 559.050 97.050 ;
        RECT 550.950 95.550 559.050 96.450 ;
        RECT 550.950 94.950 555.000 95.550 ;
        RECT 556.950 94.950 559.050 95.550 ;
        RECT 531.150 94.200 539.550 94.500 ;
        RECT 523.950 92.400 524.850 93.300 ;
        RECT 522.150 90.600 524.850 92.400 ;
        RECT 525.750 92.100 527.550 92.400 ;
        RECT 531.150 92.100 532.050 94.200 ;
        RECT 547.950 93.600 548.850 94.500 ;
        RECT 525.750 91.200 532.050 92.100 ;
        RECT 532.950 92.700 534.750 93.300 ;
        RECT 532.950 91.500 540.450 92.700 ;
        RECT 525.750 90.600 527.550 91.200 ;
        RECT 539.250 90.600 540.450 91.500 ;
        RECT 520.950 87.600 524.850 89.700 ;
        RECT 529.950 89.550 531.750 90.300 ;
        RECT 534.750 89.550 536.550 90.300 ;
        RECT 529.950 88.500 536.550 89.550 ;
        RECT 539.250 88.500 544.050 90.600 ;
        RECT 523.050 81.600 524.850 87.600 ;
        RECT 530.850 81.600 532.650 88.500 ;
        RECT 539.250 87.600 540.450 88.500 ;
        RECT 538.650 81.600 540.450 87.600 ;
        RECT 547.050 81.600 548.850 93.600 ;
        RECT 560.400 87.600 561.600 99.900 ;
        RECT 563.100 98.100 564.900 98.850 ;
        RECT 577.950 97.950 580.050 100.050 ;
        RECT 562.950 94.950 565.050 97.050 ;
        RECT 582.150 96.900 582.900 101.100 ;
        RECT 583.950 97.950 586.050 100.050 ;
        RECT 598.950 97.950 601.050 100.050 ;
        RECT 602.100 96.900 603.150 101.100 ;
        RECT 610.950 100.950 613.050 101.550 ;
        RECT 619.950 100.950 622.050 101.550 ;
        RECT 638.100 101.100 639.900 101.850 ;
        RECT 640.950 101.100 642.150 102.900 ;
        RECT 644.100 101.100 645.900 101.850 ;
        RECT 604.950 97.950 607.050 100.050 ;
        RECT 617.100 98.100 618.900 98.850 ;
        RECT 612.000 96.900 615.000 97.050 ;
        RECT 582.150 95.400 583.050 96.900 ;
        RECT 582.150 94.500 586.200 95.400 ;
        RECT 575.400 92.400 583.200 93.300 ;
        RECT 560.400 81.600 562.200 87.600 ;
        RECT 575.400 81.600 577.200 92.400 ;
        RECT 581.400 82.500 583.200 92.400 ;
        RECT 584.400 83.400 586.200 94.500 ;
        RECT 601.950 93.600 603.150 96.900 ;
        RECT 610.950 96.450 615.000 96.900 ;
        RECT 616.950 96.450 619.050 97.050 ;
        RECT 610.950 95.550 619.050 96.450 ;
        RECT 610.950 94.950 615.000 95.550 ;
        RECT 616.950 94.950 619.050 95.550 ;
        RECT 610.950 94.800 613.050 94.950 ;
        RECT 587.400 82.500 589.200 93.600 ;
        RECT 581.400 81.600 589.200 82.500 ;
        RECT 601.500 81.600 603.300 93.600 ;
        RECT 620.400 87.600 621.600 99.900 ;
        RECT 623.100 98.100 624.900 98.850 ;
        RECT 637.950 97.950 640.050 100.050 ;
        RECT 622.950 94.950 625.050 97.050 ;
        RECT 641.100 96.900 642.150 101.100 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 657.150 102.900 657.900 107.100 ;
        RECT 665.550 106.050 666.750 110.400 ;
        RECT 685.350 109.800 687.150 110.550 ;
        RECT 688.650 109.800 690.450 111.600 ;
        RECT 691.950 110.400 694.050 112.500 ;
        RECT 697.050 110.400 698.850 116.400 ;
        RECT 709.200 110.400 711.000 116.400 ;
        RECT 735.000 112.050 736.800 116.400 ;
        RECT 749.400 113.400 751.200 116.400 ;
        RECT 689.100 106.800 690.150 109.800 ;
        RECT 658.950 103.950 664.050 106.050 ;
        RECT 665.550 103.950 666.900 106.050 ;
        RECT 667.950 103.950 670.050 106.050 ;
        RECT 671.100 104.250 671.850 106.050 ;
        RECT 678.150 105.600 696.000 106.800 ;
        RECT 678.150 105.000 679.950 105.600 ;
        RECT 689.100 105.000 690.900 105.600 ;
        RECT 679.050 104.100 679.950 105.000 ;
        RECT 695.100 104.850 696.000 105.600 ;
        RECT 643.950 97.950 646.050 100.050 ;
        RECT 653.100 99.150 654.900 99.900 ;
        RECT 640.950 93.600 642.150 96.900 ;
        RECT 657.150 96.300 658.050 102.900 ;
        RECT 657.150 95.400 659.100 96.300 ;
        RECT 653.400 94.500 659.100 95.400 ;
        RECT 620.400 81.600 622.200 87.600 ;
        RECT 640.500 81.600 642.300 93.600 ;
        RECT 653.400 87.600 654.600 94.500 ;
        RECT 660.000 93.600 661.200 102.900 ;
        RECT 665.550 93.600 666.750 103.950 ;
        RECT 695.100 103.050 696.900 104.850 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 692.100 100.800 693.900 101.400 ;
        RECT 667.950 95.400 669.750 97.200 ;
        RECT 668.850 94.200 673.050 95.400 ;
        RECT 679.050 94.200 679.950 99.900 ;
        RECT 685.950 97.950 688.050 100.050 ;
        RECT 689.100 99.600 693.900 100.800 ;
        RECT 687.750 95.700 689.550 96.000 ;
        RECT 697.950 95.700 698.850 110.400 ;
        RECT 709.950 107.100 711.000 110.400 ;
        RECT 731.400 110.400 736.800 112.050 ;
        RECT 731.400 107.100 732.300 110.400 ;
        RECT 750.300 109.200 751.200 113.400 ;
        RECT 755.400 110.400 757.200 116.400 ;
        RECT 761.550 110.400 763.350 116.400 ;
        RECT 769.650 113.400 771.450 116.400 ;
        RECT 777.450 113.400 779.250 116.400 ;
        RECT 785.250 114.300 787.050 116.400 ;
        RECT 785.250 113.400 789.000 114.300 ;
        RECT 769.650 112.500 770.700 113.400 ;
        RECT 766.950 111.300 770.700 112.500 ;
        RECT 778.200 111.600 779.250 113.400 ;
        RECT 787.950 112.500 789.000 113.400 ;
        RECT 766.950 110.400 769.050 111.300 ;
        RECT 778.200 110.550 783.150 111.600 ;
        RECT 750.300 108.300 753.750 109.200 ;
        RECT 751.950 107.400 753.750 108.300 ;
        RECT 703.950 103.950 706.050 106.050 ;
        RECT 709.950 103.950 712.050 106.050 ;
        RECT 715.950 103.950 718.050 106.050 ;
        RECT 721.950 105.450 724.050 106.050 ;
        RECT 730.950 105.450 733.050 106.050 ;
        RECT 721.950 104.550 733.050 105.450 ;
        RECT 721.950 103.950 724.050 104.550 ;
        RECT 730.950 103.950 733.050 104.550 ;
        RECT 736.950 103.950 739.050 106.050 ;
        RECT 748.950 103.950 751.050 106.050 ;
        RECT 704.250 102.150 706.050 102.900 ;
        RECT 707.250 101.100 709.050 101.850 ;
        RECT 711.150 101.100 712.050 102.900 ;
        RECT 716.100 102.150 717.900 102.900 ;
        RECT 712.950 101.100 714.750 101.850 ;
        RECT 706.950 97.950 709.050 100.050 ;
        RECT 687.750 95.100 698.850 95.700 ;
        RECT 653.400 81.600 655.200 87.600 ;
        RECT 659.700 81.600 661.500 93.600 ;
        RECT 665.550 81.600 667.350 93.600 ;
        RECT 670.950 93.300 673.050 94.200 ;
        RECT 673.950 93.300 679.950 94.200 ;
        RECT 681.150 94.500 698.850 95.100 ;
        RECT 711.150 96.900 711.900 101.100 ;
        RECT 712.950 97.950 715.050 100.050 ;
        RECT 711.150 95.400 712.050 96.900 ;
        RECT 711.150 94.500 715.200 95.400 ;
        RECT 681.150 94.200 689.550 94.500 ;
        RECT 673.950 92.400 674.850 93.300 ;
        RECT 672.150 90.600 674.850 92.400 ;
        RECT 675.750 92.100 677.550 92.400 ;
        RECT 681.150 92.100 682.050 94.200 ;
        RECT 697.950 93.600 698.850 94.500 ;
        RECT 675.750 91.200 682.050 92.100 ;
        RECT 682.950 92.700 684.750 93.300 ;
        RECT 682.950 91.500 690.450 92.700 ;
        RECT 675.750 90.600 677.550 91.200 ;
        RECT 689.250 90.600 690.450 91.500 ;
        RECT 670.950 87.600 674.850 89.700 ;
        RECT 679.950 89.550 681.750 90.300 ;
        RECT 684.750 89.550 686.550 90.300 ;
        RECT 679.950 88.500 686.550 89.550 ;
        RECT 689.250 88.500 694.050 90.600 ;
        RECT 673.050 81.600 674.850 87.600 ;
        RECT 680.850 81.600 682.650 88.500 ;
        RECT 689.250 87.600 690.450 88.500 ;
        RECT 688.650 81.600 690.450 87.600 ;
        RECT 697.050 81.600 698.850 93.600 ;
        RECT 704.400 92.400 712.200 93.300 ;
        RECT 704.400 81.600 706.200 92.400 ;
        RECT 710.400 82.500 712.200 92.400 ;
        RECT 713.400 83.400 715.200 94.500 ;
        RECT 731.400 93.600 732.300 102.900 ;
        RECT 737.100 102.150 738.900 102.900 ;
        RECT 749.100 102.150 750.900 102.900 ;
        RECT 734.100 101.100 735.900 101.850 ;
        RECT 740.100 101.100 741.900 101.850 ;
        RECT 746.100 101.100 747.900 101.850 ;
        RECT 733.950 97.950 736.050 100.050 ;
        RECT 739.950 99.450 742.050 100.050 ;
        RECT 745.950 99.450 748.050 100.050 ;
        RECT 739.950 98.550 748.050 99.450 ;
        RECT 739.950 97.950 742.050 98.550 ;
        RECT 745.950 97.950 748.050 98.550 ;
        RECT 752.700 96.600 753.600 107.400 ;
        RECT 756.000 104.100 757.050 110.400 ;
        RECT 761.550 106.050 762.750 110.400 ;
        RECT 781.350 109.800 783.150 110.550 ;
        RECT 784.650 109.800 786.450 111.600 ;
        RECT 787.950 110.400 790.050 112.500 ;
        RECT 793.050 110.400 794.850 116.400 ;
        RECT 785.100 106.800 786.150 109.800 ;
        RECT 761.550 103.950 762.900 106.050 ;
        RECT 763.950 103.950 766.050 106.050 ;
        RECT 767.100 104.250 767.850 106.050 ;
        RECT 774.150 105.600 792.000 106.800 ;
        RECT 774.150 105.000 775.950 105.600 ;
        RECT 785.100 105.000 786.900 105.600 ;
        RECT 775.050 104.100 775.950 105.000 ;
        RECT 791.100 104.850 792.000 105.600 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 751.800 96.000 753.600 96.600 ;
        RECT 746.400 94.800 753.600 96.000 ;
        RECT 746.400 93.600 747.600 94.800 ;
        RECT 754.950 93.600 756.300 99.900 ;
        RECT 716.400 82.500 718.200 93.600 ;
        RECT 710.400 81.600 718.200 82.500 ;
        RECT 730.800 81.600 732.600 93.600 ;
        RECT 733.800 92.700 741.600 93.600 ;
        RECT 733.800 81.600 735.600 92.700 ;
        RECT 739.800 81.600 741.600 92.700 ;
        RECT 746.400 81.600 748.200 93.600 ;
        RECT 753.900 92.100 756.300 93.600 ;
        RECT 761.550 93.600 762.750 103.950 ;
        RECT 791.100 103.050 792.900 104.850 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 763.950 95.400 765.750 97.200 ;
        RECT 764.850 94.200 769.050 95.400 ;
        RECT 775.050 94.200 775.950 99.900 ;
        RECT 781.950 97.950 784.050 103.050 ;
        RECT 788.100 100.800 789.900 101.400 ;
        RECT 785.100 99.600 789.900 100.800 ;
        RECT 783.750 95.700 785.550 96.000 ;
        RECT 793.950 95.700 794.850 110.400 ;
        RECT 803.400 111.300 805.200 116.400 ;
        RECT 809.400 111.300 811.200 116.400 ;
        RECT 803.400 109.950 811.200 111.300 ;
        RECT 812.400 110.400 814.200 116.400 ;
        RECT 812.400 108.300 813.600 110.400 ;
        RECT 809.850 107.250 813.600 108.300 ;
        RECT 809.850 107.100 811.050 107.250 ;
        RECT 802.950 103.950 805.050 106.050 ;
        RECT 808.950 103.950 811.050 106.050 ;
        RECT 803.100 102.150 804.900 102.900 ;
        RECT 806.100 101.100 807.900 101.850 ;
        RECT 808.950 101.100 810.150 102.900 ;
        RECT 812.100 101.100 813.900 101.850 ;
        RECT 805.950 97.800 808.050 100.050 ;
        RECT 809.100 96.900 810.150 101.100 ;
        RECT 811.950 97.950 814.050 100.050 ;
        RECT 783.750 95.100 794.850 95.700 ;
        RECT 753.900 81.600 755.700 92.100 ;
        RECT 761.550 81.600 763.350 93.600 ;
        RECT 766.950 93.300 769.050 94.200 ;
        RECT 769.950 93.300 775.950 94.200 ;
        RECT 777.150 94.500 794.850 95.100 ;
        RECT 777.150 94.200 785.550 94.500 ;
        RECT 769.950 92.400 770.850 93.300 ;
        RECT 768.150 90.600 770.850 92.400 ;
        RECT 771.750 92.100 773.550 92.400 ;
        RECT 777.150 92.100 778.050 94.200 ;
        RECT 793.950 93.600 794.850 94.500 ;
        RECT 808.950 93.600 810.150 96.900 ;
        RECT 771.750 91.200 778.050 92.100 ;
        RECT 778.950 92.700 780.750 93.300 ;
        RECT 778.950 91.500 786.450 92.700 ;
        RECT 771.750 90.600 773.550 91.200 ;
        RECT 785.250 90.600 786.450 91.500 ;
        RECT 766.950 87.600 770.850 89.700 ;
        RECT 775.950 89.550 777.750 90.300 ;
        RECT 780.750 89.550 782.550 90.300 ;
        RECT 775.950 88.500 782.550 89.550 ;
        RECT 785.250 88.500 790.050 90.600 ;
        RECT 769.050 81.600 770.850 87.600 ;
        RECT 776.850 81.600 778.650 88.500 ;
        RECT 785.250 87.600 786.450 88.500 ;
        RECT 784.650 81.600 786.450 87.600 ;
        RECT 793.050 81.600 794.850 93.600 ;
        RECT 808.500 81.600 810.300 93.600 ;
        RECT 3.150 65.400 4.950 77.400 ;
        RECT 11.550 71.400 13.350 77.400 ;
        RECT 11.550 70.500 12.750 71.400 ;
        RECT 19.350 70.500 21.150 77.400 ;
        RECT 27.150 71.400 28.950 77.400 ;
        RECT 7.950 68.400 12.750 70.500 ;
        RECT 15.450 69.450 22.050 70.500 ;
        RECT 15.450 68.700 17.250 69.450 ;
        RECT 20.250 68.700 22.050 69.450 ;
        RECT 27.150 69.300 31.050 71.400 ;
        RECT 11.550 67.500 12.750 68.400 ;
        RECT 24.450 67.800 26.250 68.400 ;
        RECT 11.550 66.300 19.050 67.500 ;
        RECT 17.250 65.700 19.050 66.300 ;
        RECT 19.950 66.900 26.250 67.800 ;
        RECT 3.150 64.500 4.050 65.400 ;
        RECT 19.950 64.800 20.850 66.900 ;
        RECT 24.450 66.600 26.250 66.900 ;
        RECT 27.150 66.600 29.850 68.400 ;
        RECT 27.150 65.700 28.050 66.600 ;
        RECT 12.450 64.500 20.850 64.800 ;
        RECT 3.150 63.900 20.850 64.500 ;
        RECT 22.050 64.800 28.050 65.700 ;
        RECT 28.950 64.800 31.050 65.700 ;
        RECT 34.650 65.400 36.450 77.400 ;
        RECT 3.150 63.300 14.250 63.900 ;
        RECT 3.150 48.600 4.050 63.300 ;
        RECT 12.450 63.000 14.250 63.300 ;
        RECT 8.100 58.200 12.900 59.400 ;
        RECT 13.950 58.950 16.050 61.050 ;
        RECT 22.050 59.100 22.950 64.800 ;
        RECT 28.950 63.600 33.150 64.800 ;
        RECT 32.250 61.800 34.050 63.600 ;
        RECT 8.100 57.600 9.900 58.200 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 5.100 54.150 6.900 55.950 ;
        RECT 35.250 55.050 36.450 65.400 ;
        RECT 6.000 53.400 6.900 54.150 ;
        RECT 22.050 54.000 22.950 54.900 ;
        RECT 11.100 53.400 12.900 54.000 ;
        RECT 22.050 53.400 23.850 54.000 ;
        RECT 6.000 52.200 23.850 53.400 ;
        RECT 30.150 52.950 30.900 54.750 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 35.100 52.950 36.450 55.050 ;
        RECT 11.850 49.200 12.900 52.200 ;
        RECT 3.150 42.600 4.950 48.600 ;
        RECT 7.950 46.500 10.050 48.600 ;
        RECT 11.550 47.400 13.350 49.200 ;
        RECT 14.850 48.450 16.650 49.200 ;
        RECT 35.250 48.600 36.450 52.950 ;
        RECT 14.850 47.400 19.800 48.450 ;
        RECT 28.950 47.700 31.050 48.600 ;
        RECT 9.000 45.600 10.050 46.500 ;
        RECT 18.750 45.600 19.800 47.400 ;
        RECT 27.300 46.500 31.050 47.700 ;
        RECT 27.300 45.600 28.350 46.500 ;
        RECT 9.000 44.700 12.750 45.600 ;
        RECT 10.950 42.600 12.750 44.700 ;
        RECT 18.750 42.600 20.550 45.600 ;
        RECT 26.550 42.600 28.350 45.600 ;
        RECT 34.650 42.600 36.450 48.600 ;
        RECT 38.550 65.400 40.350 77.400 ;
        RECT 46.050 71.400 47.850 77.400 ;
        RECT 43.950 69.300 47.850 71.400 ;
        RECT 53.850 70.500 55.650 77.400 ;
        RECT 61.650 71.400 63.450 77.400 ;
        RECT 62.250 70.500 63.450 71.400 ;
        RECT 52.950 69.450 59.550 70.500 ;
        RECT 52.950 68.700 54.750 69.450 ;
        RECT 57.750 68.700 59.550 69.450 ;
        RECT 62.250 68.400 67.050 70.500 ;
        RECT 45.150 66.600 47.850 68.400 ;
        RECT 48.750 67.800 50.550 68.400 ;
        RECT 48.750 66.900 55.050 67.800 ;
        RECT 62.250 67.500 63.450 68.400 ;
        RECT 48.750 66.600 50.550 66.900 ;
        RECT 46.950 65.700 47.850 66.600 ;
        RECT 38.550 55.050 39.750 65.400 ;
        RECT 43.950 64.800 46.050 65.700 ;
        RECT 46.950 64.800 52.950 65.700 ;
        RECT 41.850 63.600 46.050 64.800 ;
        RECT 40.950 61.800 42.750 63.600 ;
        RECT 52.050 59.100 52.950 64.800 ;
        RECT 54.150 64.800 55.050 66.900 ;
        RECT 55.950 66.300 63.450 67.500 ;
        RECT 55.950 65.700 57.750 66.300 ;
        RECT 70.050 65.400 71.850 77.400 ;
        RECT 85.500 65.400 87.300 77.400 ;
        RECT 96.150 65.400 97.950 77.400 ;
        RECT 104.550 71.400 106.350 77.400 ;
        RECT 104.550 70.500 105.750 71.400 ;
        RECT 112.350 70.500 114.150 77.400 ;
        RECT 120.150 71.400 121.950 77.400 ;
        RECT 100.950 68.400 105.750 70.500 ;
        RECT 108.450 69.450 115.050 70.500 ;
        RECT 108.450 68.700 110.250 69.450 ;
        RECT 113.250 68.700 115.050 69.450 ;
        RECT 120.150 69.300 124.050 71.400 ;
        RECT 104.550 67.500 105.750 68.400 ;
        RECT 117.450 67.800 119.250 68.400 ;
        RECT 104.550 66.300 112.050 67.500 ;
        RECT 110.250 65.700 112.050 66.300 ;
        RECT 112.950 66.900 119.250 67.800 ;
        RECT 54.150 64.500 62.550 64.800 ;
        RECT 70.950 64.500 71.850 65.400 ;
        RECT 54.150 63.900 71.850 64.500 ;
        RECT 60.750 63.300 71.850 63.900 ;
        RECT 60.750 63.000 62.550 63.300 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 58.950 55.950 61.050 61.050 ;
        RECT 62.100 58.200 66.900 59.400 ;
        RECT 65.100 57.600 66.900 58.200 ;
        RECT 38.550 52.950 39.900 55.050 ;
        RECT 40.950 52.950 43.050 55.050 ;
        RECT 44.100 52.950 44.850 54.750 ;
        RECT 52.050 54.000 52.950 54.900 ;
        RECT 68.100 54.150 69.900 55.950 ;
        RECT 51.150 53.400 52.950 54.000 ;
        RECT 62.100 53.400 63.900 54.000 ;
        RECT 68.100 53.400 69.000 54.150 ;
        RECT 38.550 48.600 39.750 52.950 ;
        RECT 51.150 52.200 69.000 53.400 ;
        RECT 62.100 49.200 63.150 52.200 ;
        RECT 38.550 42.600 40.350 48.600 ;
        RECT 43.950 47.700 46.050 48.600 ;
        RECT 58.350 48.450 60.150 49.200 ;
        RECT 43.950 46.500 47.700 47.700 ;
        RECT 46.650 45.600 47.700 46.500 ;
        RECT 55.200 47.400 60.150 48.450 ;
        RECT 61.650 47.400 63.450 49.200 ;
        RECT 70.950 48.600 71.850 63.300 ;
        RECT 85.950 62.100 87.150 65.400 ;
        RECT 82.950 58.950 85.050 61.050 ;
        RECT 86.100 57.900 87.150 62.100 ;
        RECT 96.150 64.500 97.050 65.400 ;
        RECT 112.950 64.800 113.850 66.900 ;
        RECT 117.450 66.600 119.250 66.900 ;
        RECT 120.150 66.600 122.850 68.400 ;
        RECT 120.150 65.700 121.050 66.600 ;
        RECT 105.450 64.500 113.850 64.800 ;
        RECT 96.150 63.900 113.850 64.500 ;
        RECT 115.050 64.800 121.050 65.700 ;
        RECT 121.950 64.800 124.050 65.700 ;
        RECT 127.650 65.400 129.450 77.400 ;
        RECT 96.150 63.300 107.250 63.900 ;
        RECT 88.950 58.950 91.050 61.050 ;
        RECT 83.100 57.150 84.900 57.900 ;
        RECT 80.100 56.100 81.900 56.850 ;
        RECT 85.950 56.100 87.150 57.900 ;
        RECT 89.100 57.150 90.900 57.900 ;
        RECT 79.950 52.950 82.050 55.050 ;
        RECT 85.950 52.950 88.050 55.050 ;
        RECT 86.850 51.750 88.050 51.900 ;
        RECT 86.850 50.700 90.600 51.750 ;
        RECT 55.200 45.600 56.250 47.400 ;
        RECT 64.950 46.500 67.050 48.600 ;
        RECT 64.950 45.600 66.000 46.500 ;
        RECT 46.650 42.600 48.450 45.600 ;
        RECT 54.450 42.600 56.250 45.600 ;
        RECT 62.250 44.700 66.000 45.600 ;
        RECT 62.250 42.600 64.050 44.700 ;
        RECT 70.050 42.600 71.850 48.600 ;
        RECT 80.400 47.700 88.200 49.050 ;
        RECT 80.400 42.600 82.200 47.700 ;
        RECT 86.400 42.600 88.200 47.700 ;
        RECT 89.400 48.600 90.600 50.700 ;
        RECT 96.150 48.600 97.050 63.300 ;
        RECT 105.450 63.000 107.250 63.300 ;
        RECT 101.100 58.200 105.900 59.400 ;
        RECT 106.950 58.950 109.050 61.050 ;
        RECT 115.050 59.100 115.950 64.800 ;
        RECT 121.950 63.600 126.150 64.800 ;
        RECT 125.250 61.800 127.050 63.600 ;
        RECT 101.100 57.600 102.900 58.200 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 98.100 54.150 99.900 55.950 ;
        RECT 128.250 55.050 129.450 65.400 ;
        RECT 140.400 71.400 142.200 77.400 ;
        RECT 130.950 63.450 135.000 64.050 ;
        RECT 136.950 63.450 139.050 64.050 ;
        RECT 130.950 62.550 139.050 63.450 ;
        RECT 130.950 61.950 135.000 62.550 ;
        RECT 136.950 61.950 139.050 62.550 ;
        RECT 137.100 60.150 138.900 60.900 ;
        RECT 140.400 59.100 141.600 71.400 ;
        RECT 157.500 65.400 159.300 77.400 ;
        RECT 168.150 65.400 169.950 77.400 ;
        RECT 176.550 71.400 178.350 77.400 ;
        RECT 176.550 70.500 177.750 71.400 ;
        RECT 184.350 70.500 186.150 77.400 ;
        RECT 192.150 71.400 193.950 77.400 ;
        RECT 172.950 68.400 177.750 70.500 ;
        RECT 180.450 69.450 187.050 70.500 ;
        RECT 180.450 68.700 182.250 69.450 ;
        RECT 185.250 68.700 187.050 69.450 ;
        RECT 192.150 69.300 196.050 71.400 ;
        RECT 176.550 67.500 177.750 68.400 ;
        RECT 189.450 67.800 191.250 68.400 ;
        RECT 176.550 66.300 184.050 67.500 ;
        RECT 182.250 65.700 184.050 66.300 ;
        RECT 184.950 66.900 191.250 67.800 ;
        RECT 142.950 61.950 145.050 64.050 ;
        RECT 157.950 62.100 159.150 65.400 ;
        RECT 143.100 60.150 144.900 60.900 ;
        RECT 154.950 58.950 157.050 61.050 ;
        RECT 136.950 55.950 142.050 58.050 ;
        RECT 158.100 57.900 159.150 62.100 ;
        RECT 168.150 64.500 169.050 65.400 ;
        RECT 184.950 64.800 185.850 66.900 ;
        RECT 189.450 66.600 191.250 66.900 ;
        RECT 192.150 66.600 194.850 68.400 ;
        RECT 192.150 65.700 193.050 66.600 ;
        RECT 177.450 64.500 185.850 64.800 ;
        RECT 168.150 63.900 185.850 64.500 ;
        RECT 187.050 64.800 193.050 65.700 ;
        RECT 193.950 64.800 196.050 65.700 ;
        RECT 199.650 65.400 201.450 77.400 ;
        RECT 168.150 63.300 179.250 63.900 ;
        RECT 160.950 58.950 163.050 61.050 ;
        RECT 155.100 57.150 156.900 57.900 ;
        RECT 152.100 56.100 153.900 56.850 ;
        RECT 157.950 56.100 159.150 57.900 ;
        RECT 161.100 57.150 162.900 57.900 ;
        RECT 99.000 53.400 99.900 54.150 ;
        RECT 115.050 54.000 115.950 54.900 ;
        RECT 104.100 53.400 105.900 54.000 ;
        RECT 115.050 53.400 116.850 54.000 ;
        RECT 99.000 52.200 116.850 53.400 ;
        RECT 123.150 52.950 123.900 54.750 ;
        RECT 124.950 52.950 127.050 55.050 ;
        RECT 128.100 52.950 129.450 55.050 ;
        RECT 104.850 49.200 105.900 52.200 ;
        RECT 89.400 42.600 91.200 48.600 ;
        RECT 96.150 42.600 97.950 48.600 ;
        RECT 100.950 46.500 103.050 48.600 ;
        RECT 104.550 47.400 106.350 49.200 ;
        RECT 107.850 48.450 109.650 49.200 ;
        RECT 128.250 48.600 129.450 52.950 ;
        RECT 140.400 50.700 141.600 54.900 ;
        RECT 151.950 52.950 154.050 55.050 ;
        RECT 157.950 54.450 160.050 55.050 ;
        RECT 162.000 54.450 166.050 55.050 ;
        RECT 157.950 53.550 166.050 54.450 ;
        RECT 157.950 52.950 160.050 53.550 ;
        RECT 162.000 52.950 166.050 53.550 ;
        RECT 158.850 51.750 160.050 51.900 ;
        RECT 158.850 50.700 162.600 51.750 ;
        RECT 140.400 49.800 144.000 50.700 ;
        RECT 107.850 47.400 112.800 48.450 ;
        RECT 121.950 47.700 124.050 48.600 ;
        RECT 102.000 45.600 103.050 46.500 ;
        RECT 111.750 45.600 112.800 47.400 ;
        RECT 120.300 46.500 124.050 47.700 ;
        RECT 120.300 45.600 121.350 46.500 ;
        RECT 102.000 44.700 105.750 45.600 ;
        RECT 103.950 42.600 105.750 44.700 ;
        RECT 111.750 42.600 113.550 45.600 ;
        RECT 119.550 42.600 121.350 45.600 ;
        RECT 127.650 42.600 129.450 48.600 ;
        RECT 142.200 42.600 144.000 49.800 ;
        RECT 152.400 47.700 160.200 49.050 ;
        RECT 152.400 42.600 154.200 47.700 ;
        RECT 158.400 42.600 160.200 47.700 ;
        RECT 161.400 48.600 162.600 50.700 ;
        RECT 168.150 48.600 169.050 63.300 ;
        RECT 177.450 63.000 179.250 63.300 ;
        RECT 173.100 58.200 177.900 59.400 ;
        RECT 178.950 58.950 181.050 61.050 ;
        RECT 187.050 59.100 187.950 64.800 ;
        RECT 193.950 63.600 198.150 64.800 ;
        RECT 197.250 61.800 199.050 63.600 ;
        RECT 173.100 57.600 174.900 58.200 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 170.100 54.150 171.900 55.950 ;
        RECT 200.250 55.050 201.450 65.400 ;
        RECT 212.400 71.400 214.200 77.400 ;
        RECT 205.950 61.950 211.050 64.050 ;
        RECT 209.100 60.150 210.900 60.900 ;
        RECT 212.400 59.100 213.600 71.400 ;
        RECT 222.150 65.400 223.950 77.400 ;
        RECT 230.550 71.400 232.350 77.400 ;
        RECT 230.550 70.500 231.750 71.400 ;
        RECT 238.350 70.500 240.150 77.400 ;
        RECT 246.150 71.400 247.950 77.400 ;
        RECT 226.950 68.400 231.750 70.500 ;
        RECT 234.450 69.450 241.050 70.500 ;
        RECT 234.450 68.700 236.250 69.450 ;
        RECT 239.250 68.700 241.050 69.450 ;
        RECT 246.150 69.300 250.050 71.400 ;
        RECT 230.550 67.500 231.750 68.400 ;
        RECT 243.450 67.800 245.250 68.400 ;
        RECT 230.550 66.300 238.050 67.500 ;
        RECT 236.250 65.700 238.050 66.300 ;
        RECT 238.950 66.900 245.250 67.800 ;
        RECT 222.150 64.500 223.050 65.400 ;
        RECT 238.950 64.800 239.850 66.900 ;
        RECT 243.450 66.600 245.250 66.900 ;
        RECT 246.150 66.600 248.850 68.400 ;
        RECT 246.150 65.700 247.050 66.600 ;
        RECT 231.450 64.500 239.850 64.800 ;
        RECT 214.950 61.950 217.050 64.050 ;
        RECT 222.150 63.900 239.850 64.500 ;
        RECT 241.050 64.800 247.050 65.700 ;
        RECT 247.950 64.800 250.050 65.700 ;
        RECT 253.650 65.400 255.450 77.400 ;
        RECT 222.150 63.300 233.250 63.900 ;
        RECT 215.100 60.150 216.900 60.900 ;
        RECT 202.950 57.450 205.050 58.050 ;
        RECT 211.950 57.450 214.050 58.050 ;
        RECT 202.950 56.550 214.050 57.450 ;
        RECT 202.950 55.950 205.050 56.550 ;
        RECT 211.950 55.950 214.050 56.550 ;
        RECT 171.000 53.400 171.900 54.150 ;
        RECT 187.050 54.000 187.950 54.900 ;
        RECT 176.100 53.400 177.900 54.000 ;
        RECT 187.050 53.400 188.850 54.000 ;
        RECT 171.000 52.200 188.850 53.400 ;
        RECT 195.150 52.950 195.900 54.750 ;
        RECT 196.950 52.950 199.050 55.050 ;
        RECT 200.100 52.950 201.450 55.050 ;
        RECT 176.850 49.200 177.900 52.200 ;
        RECT 161.400 42.600 163.200 48.600 ;
        RECT 168.150 42.600 169.950 48.600 ;
        RECT 172.950 46.500 175.050 48.600 ;
        RECT 176.550 47.400 178.350 49.200 ;
        RECT 179.850 48.450 181.650 49.200 ;
        RECT 200.250 48.600 201.450 52.950 ;
        RECT 212.400 50.700 213.600 54.900 ;
        RECT 212.400 49.800 216.000 50.700 ;
        RECT 179.850 47.400 184.800 48.450 ;
        RECT 193.950 47.700 196.050 48.600 ;
        RECT 174.000 45.600 175.050 46.500 ;
        RECT 183.750 45.600 184.800 47.400 ;
        RECT 192.300 46.500 196.050 47.700 ;
        RECT 192.300 45.600 193.350 46.500 ;
        RECT 174.000 44.700 177.750 45.600 ;
        RECT 175.950 42.600 177.750 44.700 ;
        RECT 183.750 42.600 185.550 45.600 ;
        RECT 191.550 42.600 193.350 45.600 ;
        RECT 199.650 42.600 201.450 48.600 ;
        RECT 214.200 42.600 216.000 49.800 ;
        RECT 222.150 48.600 223.050 63.300 ;
        RECT 231.450 63.000 233.250 63.300 ;
        RECT 227.100 58.200 231.900 59.400 ;
        RECT 232.950 58.950 235.050 61.050 ;
        RECT 241.050 59.100 241.950 64.800 ;
        RECT 247.950 63.600 252.150 64.800 ;
        RECT 251.250 61.800 253.050 63.600 ;
        RECT 227.100 57.600 228.900 58.200 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 224.100 54.150 225.900 55.950 ;
        RECT 254.250 55.050 255.450 65.400 ;
        RECT 263.400 71.400 265.200 77.400 ;
        RECT 256.950 61.950 262.050 64.050 ;
        RECT 260.100 60.150 261.900 60.900 ;
        RECT 263.400 59.100 264.600 71.400 ;
        RECT 281.700 65.400 283.500 77.400 ;
        RECT 299.400 71.400 301.200 77.400 ;
        RECT 265.950 61.950 268.050 64.050 ;
        RECT 281.850 62.100 283.050 65.400 ;
        RECT 289.950 63.450 294.000 64.050 ;
        RECT 295.950 63.450 298.050 64.050 ;
        RECT 289.950 62.550 298.050 63.450 ;
        RECT 266.100 60.150 267.900 60.900 ;
        RECT 277.950 58.950 280.050 61.050 ;
        RECT 259.950 55.950 265.050 58.050 ;
        RECT 281.850 57.900 282.900 62.100 ;
        RECT 289.950 61.950 294.000 62.550 ;
        RECT 295.950 61.950 298.050 62.550 ;
        RECT 283.950 58.950 286.050 61.050 ;
        RECT 296.100 60.150 297.900 60.900 ;
        RECT 299.400 59.100 300.600 71.400 ;
        RECT 311.400 66.600 313.200 77.400 ;
        RECT 317.400 76.500 325.200 77.400 ;
        RECT 317.400 66.600 319.200 76.500 ;
        RECT 311.400 65.700 319.200 66.600 ;
        RECT 320.400 64.500 322.200 75.600 ;
        RECT 323.400 65.400 325.200 76.500 ;
        RECT 341.700 65.400 343.500 77.400 ;
        RECT 355.800 71.400 357.600 77.400 ;
        RECT 301.950 61.950 304.050 64.050 ;
        RECT 318.150 63.600 322.200 64.500 ;
        RECT 318.150 62.100 319.050 63.600 ;
        RECT 341.850 62.100 343.050 65.400 ;
        RECT 356.400 62.100 357.600 71.400 ;
        RECT 363.150 65.400 364.950 77.400 ;
        RECT 371.550 71.400 373.350 77.400 ;
        RECT 371.550 70.500 372.750 71.400 ;
        RECT 379.350 70.500 381.150 77.400 ;
        RECT 387.150 71.400 388.950 77.400 ;
        RECT 367.950 68.400 372.750 70.500 ;
        RECT 375.450 69.450 382.050 70.500 ;
        RECT 375.450 68.700 377.250 69.450 ;
        RECT 380.250 68.700 382.050 69.450 ;
        RECT 387.150 69.300 391.050 71.400 ;
        RECT 371.550 67.500 372.750 68.400 ;
        RECT 384.450 67.800 386.250 68.400 ;
        RECT 371.550 66.300 379.050 67.500 ;
        RECT 377.250 65.700 379.050 66.300 ;
        RECT 379.950 66.900 386.250 67.800 ;
        RECT 363.150 64.500 364.050 65.400 ;
        RECT 379.950 64.800 380.850 66.900 ;
        RECT 384.450 66.600 386.250 66.900 ;
        RECT 387.150 66.600 389.850 68.400 ;
        RECT 387.150 65.700 388.050 66.600 ;
        RECT 372.450 64.500 380.850 64.800 ;
        RECT 363.150 63.900 380.850 64.500 ;
        RECT 382.050 64.800 388.050 65.700 ;
        RECT 388.950 64.800 391.050 65.700 ;
        RECT 394.650 65.400 396.450 77.400 ;
        RECT 403.800 76.500 411.600 77.400 ;
        RECT 403.800 65.400 405.600 76.500 ;
        RECT 363.150 63.300 374.250 63.900 ;
        RECT 302.100 60.150 303.900 60.900 ;
        RECT 313.950 58.950 316.050 61.050 ;
        RECT 278.100 57.150 279.900 57.900 ;
        RECT 281.850 56.100 283.050 57.900 ;
        RECT 284.100 57.150 285.900 57.900 ;
        RECT 292.950 57.450 297.000 58.050 ;
        RECT 298.950 57.450 301.050 58.050 ;
        RECT 318.150 57.900 318.900 62.100 ;
        RECT 319.950 58.950 322.050 61.050 ;
        RECT 337.950 58.950 340.050 61.050 ;
        RECT 341.850 57.900 342.900 62.100 ;
        RECT 343.950 58.950 346.050 61.050 ;
        RECT 349.950 60.450 354.000 61.050 ;
        RECT 355.950 60.450 358.050 61.050 ;
        RECT 349.950 59.550 358.050 60.450 ;
        RECT 349.950 58.950 354.000 59.550 ;
        RECT 355.950 58.950 358.050 59.550 ;
        RECT 287.100 56.100 288.900 56.850 ;
        RECT 292.950 56.550 301.050 57.450 ;
        RECT 314.250 57.150 316.050 57.900 ;
        RECT 292.950 55.950 297.000 56.550 ;
        RECT 298.950 55.950 301.050 56.550 ;
        RECT 311.250 56.100 313.050 56.850 ;
        RECT 318.150 56.100 319.050 57.900 ;
        RECT 319.950 57.150 321.750 57.900 ;
        RECT 338.100 57.150 339.900 57.900 ;
        RECT 323.100 56.100 324.900 56.850 ;
        RECT 341.850 56.100 343.050 57.900 ;
        RECT 344.100 57.150 345.900 57.900 ;
        RECT 347.100 56.100 348.900 56.850 ;
        RECT 225.000 53.400 225.900 54.150 ;
        RECT 241.050 54.000 241.950 54.900 ;
        RECT 230.100 53.400 231.900 54.000 ;
        RECT 241.050 53.400 242.850 54.000 ;
        RECT 225.000 52.200 242.850 53.400 ;
        RECT 249.150 52.950 249.900 54.750 ;
        RECT 250.950 52.950 253.050 55.050 ;
        RECT 254.100 52.950 255.450 55.050 ;
        RECT 230.850 49.200 231.900 52.200 ;
        RECT 222.150 42.600 223.950 48.600 ;
        RECT 226.950 46.500 229.050 48.600 ;
        RECT 230.550 47.400 232.350 49.200 ;
        RECT 233.850 48.450 235.650 49.200 ;
        RECT 254.250 48.600 255.450 52.950 ;
        RECT 263.400 50.700 264.600 54.900 ;
        RECT 268.950 54.450 271.050 55.050 ;
        RECT 280.950 54.450 283.050 55.050 ;
        RECT 268.950 53.550 283.050 54.450 ;
        RECT 268.950 52.950 271.050 53.550 ;
        RECT 280.950 52.950 283.050 53.550 ;
        RECT 286.950 52.950 289.050 55.050 ;
        RECT 280.950 51.750 282.150 51.900 ;
        RECT 278.400 50.700 282.150 51.750 ;
        RECT 299.400 50.700 300.600 54.900 ;
        RECT 310.950 52.950 313.050 55.050 ;
        RECT 316.950 52.950 319.050 55.050 ;
        RECT 322.950 52.950 325.050 55.050 ;
        RECT 340.950 52.950 343.050 55.050 ;
        RECT 346.950 52.950 349.050 55.050 ;
        RECT 263.400 49.800 267.000 50.700 ;
        RECT 233.850 47.400 238.800 48.450 ;
        RECT 247.950 47.700 250.050 48.600 ;
        RECT 228.000 45.600 229.050 46.500 ;
        RECT 237.750 45.600 238.800 47.400 ;
        RECT 246.300 46.500 250.050 47.700 ;
        RECT 246.300 45.600 247.350 46.500 ;
        RECT 228.000 44.700 231.750 45.600 ;
        RECT 229.950 42.600 231.750 44.700 ;
        RECT 237.750 42.600 239.550 45.600 ;
        RECT 245.550 42.600 247.350 45.600 ;
        RECT 253.650 42.600 255.450 48.600 ;
        RECT 265.200 42.600 267.000 49.800 ;
        RECT 278.400 48.600 279.600 50.700 ;
        RECT 299.400 49.800 303.000 50.700 ;
        RECT 277.800 42.600 279.600 48.600 ;
        RECT 280.800 47.700 288.600 49.050 ;
        RECT 280.800 42.600 282.600 47.700 ;
        RECT 286.800 42.600 288.600 47.700 ;
        RECT 301.200 42.600 303.000 49.800 ;
        RECT 316.950 48.600 318.000 51.900 ;
        RECT 340.950 51.750 342.150 51.900 ;
        RECT 338.400 50.700 342.150 51.750 ;
        RECT 338.400 48.600 339.600 50.700 ;
        RECT 316.200 42.600 318.000 48.600 ;
        RECT 337.800 42.600 339.600 48.600 ;
        RECT 340.800 47.700 348.600 49.050 ;
        RECT 340.800 42.600 342.600 47.700 ;
        RECT 346.800 42.600 348.600 47.700 ;
        RECT 356.400 45.600 357.600 57.900 ;
        RECT 359.100 56.100 360.900 56.850 ;
        RECT 358.950 52.950 361.050 55.050 ;
        RECT 355.800 42.600 357.600 45.600 ;
        RECT 363.150 48.600 364.050 63.300 ;
        RECT 372.450 63.000 374.250 63.300 ;
        RECT 368.100 58.200 372.900 59.400 ;
        RECT 373.950 58.950 376.050 61.050 ;
        RECT 382.050 59.100 382.950 64.800 ;
        RECT 388.950 63.600 393.150 64.800 ;
        RECT 392.250 61.800 394.050 63.600 ;
        RECT 368.100 57.600 369.900 58.200 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 365.100 54.150 366.900 55.950 ;
        RECT 395.250 55.050 396.450 65.400 ;
        RECT 406.800 64.500 408.600 75.600 ;
        RECT 409.800 66.600 411.600 76.500 ;
        RECT 415.800 66.600 417.600 77.400 ;
        RECT 409.800 65.700 417.600 66.600 ;
        RECT 427.500 65.400 429.300 77.400 ;
        RECT 433.800 71.400 435.600 77.400 ;
        RECT 406.800 63.600 410.850 64.500 ;
        RECT 409.950 62.100 410.850 63.600 ;
        RECT 406.950 58.950 409.050 61.050 ;
        RECT 410.100 57.900 410.850 62.100 ;
        RECT 412.950 58.950 415.050 61.050 ;
        RECT 407.250 57.150 409.050 57.900 ;
        RECT 404.100 56.100 405.900 56.850 ;
        RECT 409.950 56.100 410.850 57.900 ;
        RECT 412.950 57.150 414.750 57.900 ;
        RECT 415.950 56.100 417.750 56.850 ;
        RECT 366.000 53.400 366.900 54.150 ;
        RECT 382.050 54.000 382.950 54.900 ;
        RECT 371.100 53.400 372.900 54.000 ;
        RECT 382.050 53.400 383.850 54.000 ;
        RECT 366.000 52.200 383.850 53.400 ;
        RECT 390.150 52.950 390.900 54.750 ;
        RECT 391.950 52.950 394.050 55.050 ;
        RECT 395.100 52.950 396.450 55.050 ;
        RECT 403.950 52.950 406.050 55.050 ;
        RECT 371.850 49.200 372.900 52.200 ;
        RECT 363.150 42.600 364.950 48.600 ;
        RECT 367.950 46.500 370.050 48.600 ;
        RECT 371.550 47.400 373.350 49.200 ;
        RECT 374.850 48.450 376.650 49.200 ;
        RECT 395.250 48.600 396.450 52.950 ;
        RECT 409.950 52.800 412.050 55.050 ;
        RECT 415.950 52.950 418.050 55.050 ;
        RECT 421.950 54.450 424.050 58.050 ;
        RECT 427.800 56.100 429.000 65.400 ;
        RECT 434.400 64.500 435.600 71.400 ;
        RECT 447.600 65.400 449.400 77.400 ;
        RECT 429.900 63.600 435.600 64.500 ;
        RECT 446.700 64.350 449.400 65.400 ;
        RECT 464.400 71.400 466.200 77.400 ;
        RECT 429.900 62.700 431.850 63.600 ;
        RECT 430.950 56.100 431.850 62.700 ;
        RECT 443.100 62.100 444.900 62.850 ;
        RECT 434.100 59.100 435.900 59.850 ;
        RECT 442.950 58.950 445.050 61.050 ;
        RECT 446.700 59.100 448.050 64.350 ;
        RECT 464.400 62.100 465.600 71.400 ;
        RECT 481.500 65.400 483.300 77.400 ;
        RECT 503.700 65.400 505.500 77.400 ;
        RECT 520.800 71.400 522.600 77.400 ;
        RECT 481.950 62.100 483.150 65.400 ;
        RECT 449.100 59.100 450.900 59.850 ;
        RECT 427.950 54.450 430.050 55.050 ;
        RECT 421.950 54.000 430.050 54.450 ;
        RECT 422.550 53.550 430.050 54.000 ;
        RECT 427.950 52.950 430.050 53.550 ;
        RECT 431.100 51.900 431.850 56.100 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 446.700 54.900 447.900 59.100 ;
        RECT 463.950 58.950 466.050 61.050 ;
        RECT 478.950 58.950 481.050 61.050 ;
        RECT 448.950 55.950 451.050 58.050 ;
        RECT 482.100 57.900 483.150 62.100 ;
        RECT 503.850 62.100 505.050 65.400 ;
        RECT 521.400 62.100 522.600 71.400 ;
        RECT 528.150 65.400 529.950 77.400 ;
        RECT 536.550 71.400 538.350 77.400 ;
        RECT 536.550 70.500 537.750 71.400 ;
        RECT 544.350 70.500 546.150 77.400 ;
        RECT 552.150 71.400 553.950 77.400 ;
        RECT 532.950 68.400 537.750 70.500 ;
        RECT 540.450 69.450 547.050 70.500 ;
        RECT 540.450 68.700 542.250 69.450 ;
        RECT 545.250 68.700 547.050 69.450 ;
        RECT 552.150 69.300 556.050 71.400 ;
        RECT 536.550 67.500 537.750 68.400 ;
        RECT 549.450 67.800 551.250 68.400 ;
        RECT 536.550 66.300 544.050 67.500 ;
        RECT 542.250 65.700 544.050 66.300 ;
        RECT 544.950 66.900 551.250 67.800 ;
        RECT 528.150 64.500 529.050 65.400 ;
        RECT 544.950 64.800 545.850 66.900 ;
        RECT 549.450 66.600 551.250 66.900 ;
        RECT 552.150 66.600 554.850 68.400 ;
        RECT 552.150 65.700 553.050 66.600 ;
        RECT 537.450 64.500 545.850 64.800 ;
        RECT 528.150 63.900 545.850 64.500 ;
        RECT 547.050 64.800 553.050 65.700 ;
        RECT 553.950 64.800 556.050 65.700 ;
        RECT 559.650 65.400 561.450 77.400 ;
        RECT 528.150 63.300 539.250 63.900 ;
        RECT 484.950 58.950 487.050 61.050 ;
        RECT 499.950 58.950 502.050 61.050 ;
        RECT 503.850 57.900 504.900 62.100 ;
        RECT 505.950 58.950 508.050 61.050 ;
        RECT 520.950 58.950 523.050 61.050 ;
        RECT 461.100 56.100 462.900 56.850 ;
        RECT 446.700 53.100 448.050 54.900 ;
        RECT 460.950 52.950 463.050 55.050 ;
        RECT 374.850 47.400 379.800 48.450 ;
        RECT 388.950 47.700 391.050 48.600 ;
        RECT 369.000 45.600 370.050 46.500 ;
        RECT 378.750 45.600 379.800 47.400 ;
        RECT 387.300 46.500 391.050 47.700 ;
        RECT 387.300 45.600 388.350 46.500 ;
        RECT 369.000 44.700 372.750 45.600 ;
        RECT 370.950 42.600 372.750 44.700 ;
        RECT 378.750 42.600 380.550 45.600 ;
        RECT 386.550 42.600 388.350 45.600 ;
        RECT 394.650 42.600 396.450 48.600 ;
        RECT 411.000 48.600 412.050 51.900 ;
        RECT 427.800 48.600 429.000 51.900 ;
        RECT 430.950 51.300 431.850 51.900 ;
        RECT 429.900 50.400 431.850 51.300 ;
        RECT 429.900 49.500 435.000 50.400 ;
        RECT 445.950 49.950 448.050 52.050 ;
        RECT 411.000 42.600 412.800 48.600 ;
        RECT 427.500 42.600 429.300 48.600 ;
        RECT 433.800 45.600 435.000 49.500 ;
        RECT 446.400 45.600 447.600 48.900 ;
        RECT 464.400 45.600 465.600 57.900 ;
        RECT 479.100 57.150 480.900 57.900 ;
        RECT 476.100 56.100 477.900 56.850 ;
        RECT 481.950 56.100 483.150 57.900 ;
        RECT 485.100 57.150 486.900 57.900 ;
        RECT 500.100 57.150 501.900 57.900 ;
        RECT 503.850 56.100 505.050 57.900 ;
        RECT 506.100 57.150 507.900 57.900 ;
        RECT 509.100 56.100 510.900 56.850 ;
        RECT 475.950 52.950 478.050 55.050 ;
        RECT 481.950 52.950 484.050 55.050 ;
        RECT 487.950 54.450 490.050 55.050 ;
        RECT 502.950 54.450 505.050 55.050 ;
        RECT 487.950 53.550 505.050 54.450 ;
        RECT 487.950 52.950 490.050 53.550 ;
        RECT 502.950 52.950 505.050 53.550 ;
        RECT 508.950 52.950 511.050 55.200 ;
        RECT 482.850 51.750 484.050 51.900 ;
        RECT 502.950 51.750 504.150 51.900 ;
        RECT 482.850 50.700 486.600 51.750 ;
        RECT 476.400 47.700 484.200 49.050 ;
        RECT 433.800 42.600 435.600 45.600 ;
        RECT 446.400 42.600 448.200 45.600 ;
        RECT 464.400 42.600 466.200 45.600 ;
        RECT 476.400 42.600 478.200 47.700 ;
        RECT 482.400 42.600 484.200 47.700 ;
        RECT 485.400 48.600 486.600 50.700 ;
        RECT 500.400 50.700 504.150 51.750 ;
        RECT 500.400 48.600 501.600 50.700 ;
        RECT 485.400 42.600 487.200 48.600 ;
        RECT 499.800 42.600 501.600 48.600 ;
        RECT 502.800 47.700 510.600 49.050 ;
        RECT 502.800 42.600 504.600 47.700 ;
        RECT 508.800 42.600 510.600 47.700 ;
        RECT 521.400 45.600 522.600 57.900 ;
        RECT 524.100 56.100 525.900 56.850 ;
        RECT 523.950 52.950 526.050 55.050 ;
        RECT 520.800 42.600 522.600 45.600 ;
        RECT 528.150 48.600 529.050 63.300 ;
        RECT 537.450 63.000 539.250 63.300 ;
        RECT 533.100 58.200 537.900 59.400 ;
        RECT 538.950 58.950 541.050 61.050 ;
        RECT 547.050 59.100 547.950 64.800 ;
        RECT 553.950 63.600 558.150 64.800 ;
        RECT 557.250 61.800 559.050 63.600 ;
        RECT 533.100 57.600 534.900 58.200 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 530.100 54.150 531.900 55.950 ;
        RECT 560.250 55.050 561.450 65.400 ;
        RECT 572.400 71.400 574.200 77.400 ;
        RECT 572.400 62.100 573.600 71.400 ;
        RECT 579.150 65.400 580.950 77.400 ;
        RECT 587.550 71.400 589.350 77.400 ;
        RECT 587.550 70.500 588.750 71.400 ;
        RECT 595.350 70.500 597.150 77.400 ;
        RECT 603.150 71.400 604.950 77.400 ;
        RECT 583.950 68.400 588.750 70.500 ;
        RECT 591.450 69.450 598.050 70.500 ;
        RECT 591.450 68.700 593.250 69.450 ;
        RECT 596.250 68.700 598.050 69.450 ;
        RECT 603.150 69.300 607.050 71.400 ;
        RECT 587.550 67.500 588.750 68.400 ;
        RECT 600.450 67.800 602.250 68.400 ;
        RECT 587.550 66.300 595.050 67.500 ;
        RECT 593.250 65.700 595.050 66.300 ;
        RECT 595.950 66.900 602.250 67.800 ;
        RECT 579.150 64.500 580.050 65.400 ;
        RECT 595.950 64.800 596.850 66.900 ;
        RECT 600.450 66.600 602.250 66.900 ;
        RECT 603.150 66.600 605.850 68.400 ;
        RECT 603.150 65.700 604.050 66.600 ;
        RECT 588.450 64.500 596.850 64.800 ;
        RECT 579.150 63.900 596.850 64.500 ;
        RECT 598.050 64.800 604.050 65.700 ;
        RECT 604.950 64.800 607.050 65.700 ;
        RECT 610.650 65.400 612.450 77.400 ;
        RECT 626.700 65.400 628.500 77.400 ;
        RECT 643.800 65.400 645.600 77.400 ;
        RECT 579.150 63.300 590.250 63.900 ;
        RECT 571.950 58.950 574.050 61.050 ;
        RECT 569.100 56.100 570.900 56.850 ;
        RECT 531.000 53.400 531.900 54.150 ;
        RECT 547.050 54.000 547.950 54.900 ;
        RECT 536.100 53.400 537.900 54.000 ;
        RECT 547.050 53.400 548.850 54.000 ;
        RECT 531.000 52.200 548.850 53.400 ;
        RECT 555.150 52.950 555.900 54.750 ;
        RECT 556.950 52.950 559.050 55.050 ;
        RECT 560.100 52.950 561.450 55.050 ;
        RECT 568.950 52.950 571.050 55.050 ;
        RECT 536.850 49.200 537.900 52.200 ;
        RECT 528.150 42.600 529.950 48.600 ;
        RECT 532.950 46.500 535.050 48.600 ;
        RECT 536.550 47.400 538.350 49.200 ;
        RECT 539.850 48.450 541.650 49.200 ;
        RECT 560.250 48.600 561.450 52.950 ;
        RECT 539.850 47.400 544.800 48.450 ;
        RECT 553.950 47.700 556.050 48.600 ;
        RECT 534.000 45.600 535.050 46.500 ;
        RECT 543.750 45.600 544.800 47.400 ;
        RECT 552.300 46.500 556.050 47.700 ;
        RECT 552.300 45.600 553.350 46.500 ;
        RECT 534.000 44.700 537.750 45.600 ;
        RECT 535.950 42.600 537.750 44.700 ;
        RECT 543.750 42.600 545.550 45.600 ;
        RECT 551.550 42.600 553.350 45.600 ;
        RECT 559.650 42.600 561.450 48.600 ;
        RECT 572.400 45.600 573.600 57.900 ;
        RECT 579.150 48.600 580.050 63.300 ;
        RECT 588.450 63.000 590.250 63.300 ;
        RECT 584.100 58.200 588.900 59.400 ;
        RECT 589.950 58.950 592.050 61.050 ;
        RECT 598.050 59.100 598.950 64.800 ;
        RECT 604.950 63.600 609.150 64.800 ;
        RECT 608.250 61.800 610.050 63.600 ;
        RECT 584.100 57.600 585.900 58.200 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 581.100 54.150 582.900 55.950 ;
        RECT 611.250 55.050 612.450 65.400 ;
        RECT 626.850 62.100 628.050 65.400 ;
        RECT 644.400 64.500 645.600 65.400 ;
        RECT 649.800 64.500 651.600 77.400 ;
        RECT 644.400 63.600 651.600 64.500 ;
        RECT 662.400 71.400 664.200 77.400 ;
        RECT 662.400 64.500 663.600 71.400 ;
        RECT 668.700 65.400 670.500 77.400 ;
        RECT 685.800 71.400 687.600 77.400 ;
        RECT 662.400 63.600 668.100 64.500 ;
        RECT 622.950 58.950 625.050 61.050 ;
        RECT 626.850 57.900 627.900 62.100 ;
        RECT 628.950 58.800 631.050 61.050 ;
        RECT 623.100 57.150 624.900 57.900 ;
        RECT 626.850 56.100 628.050 57.900 ;
        RECT 629.100 57.150 630.900 57.900 ;
        RECT 632.100 56.100 633.900 56.850 ;
        RECT 644.400 56.100 645.600 63.600 ;
        RECT 666.150 62.700 668.100 63.600 ;
        RECT 650.100 59.100 651.900 59.850 ;
        RECT 662.100 59.100 663.900 59.850 ;
        RECT 649.950 55.950 652.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 666.150 56.100 667.050 62.700 ;
        RECT 669.000 56.100 670.200 65.400 ;
        RECT 682.950 61.950 685.050 64.050 ;
        RECT 683.100 60.150 684.900 60.900 ;
        RECT 686.400 59.100 687.600 71.400 ;
        RECT 701.400 71.400 703.200 77.400 ;
        RECT 688.950 61.950 691.050 64.050 ;
        RECT 701.400 62.100 702.600 71.400 ;
        RECT 719.700 65.400 721.500 77.400 ;
        RECT 734.400 71.400 736.200 77.400 ;
        RECT 719.850 62.100 721.050 65.400 ;
        RECT 689.100 60.150 690.900 60.900 ;
        RECT 697.950 58.950 703.050 61.050 ;
        RECT 715.950 58.950 718.050 61.050 ;
        RECT 582.000 53.400 582.900 54.150 ;
        RECT 598.050 54.000 598.950 54.900 ;
        RECT 587.100 53.400 588.900 54.000 ;
        RECT 598.050 53.400 599.850 54.000 ;
        RECT 582.000 52.200 599.850 53.400 ;
        RECT 606.150 52.950 606.900 54.750 ;
        RECT 607.950 52.950 610.050 55.050 ;
        RECT 611.100 52.950 612.450 55.050 ;
        RECT 619.950 54.450 624.000 55.050 ;
        RECT 625.950 54.450 628.050 55.050 ;
        RECT 619.950 53.550 628.050 54.450 ;
        RECT 619.950 52.950 624.000 53.550 ;
        RECT 625.950 52.950 628.050 53.550 ;
        RECT 631.950 52.950 634.050 55.050 ;
        RECT 643.950 52.950 646.050 55.050 ;
        RECT 587.850 49.200 588.900 52.200 ;
        RECT 572.400 42.600 574.200 45.600 ;
        RECT 579.150 42.600 580.950 48.600 ;
        RECT 583.950 46.500 586.050 48.600 ;
        RECT 587.550 47.400 589.350 49.200 ;
        RECT 590.850 48.450 592.650 49.200 ;
        RECT 611.250 48.600 612.450 52.950 ;
        RECT 666.150 51.900 666.900 56.100 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 719.850 57.900 720.900 62.100 ;
        RECT 730.950 61.950 733.050 64.050 ;
        RECT 721.950 58.950 724.050 61.050 ;
        RECT 731.100 60.150 732.900 60.900 ;
        RECT 734.400 59.100 735.600 71.400 ;
        RECT 754.500 65.400 756.300 77.400 ;
        RECT 776.700 65.400 778.500 77.400 ;
        RECT 791.400 71.400 793.200 77.400 ;
        RECT 806.400 71.400 808.200 77.400 ;
        RECT 815.400 71.400 817.200 77.400 ;
        RECT 736.950 61.950 739.050 64.050 ;
        RECT 754.950 62.100 756.150 65.400 ;
        RECT 737.100 60.150 738.900 60.900 ;
        RECT 751.950 58.950 754.050 61.050 ;
        RECT 698.100 56.100 699.900 56.850 ;
        RECT 667.950 52.950 670.050 55.050 ;
        RECT 625.950 51.750 627.150 51.900 ;
        RECT 623.400 50.700 627.150 51.750 ;
        RECT 644.400 50.700 645.600 51.900 ;
        RECT 666.150 51.300 667.050 51.900 ;
        RECT 623.400 48.600 624.600 50.700 ;
        RECT 644.400 49.500 651.600 50.700 ;
        RECT 666.150 50.400 668.100 51.300 ;
        RECT 590.850 47.400 595.800 48.450 ;
        RECT 604.950 47.700 607.050 48.600 ;
        RECT 585.000 45.600 586.050 46.500 ;
        RECT 594.750 45.600 595.800 47.400 ;
        RECT 603.300 46.500 607.050 47.700 ;
        RECT 603.300 45.600 604.350 46.500 ;
        RECT 585.000 44.700 588.750 45.600 ;
        RECT 586.950 42.600 588.750 44.700 ;
        RECT 594.750 42.600 596.550 45.600 ;
        RECT 602.550 42.600 604.350 45.600 ;
        RECT 610.650 42.600 612.450 48.600 ;
        RECT 622.800 42.600 624.600 48.600 ;
        RECT 625.800 47.700 633.600 49.050 ;
        RECT 644.400 48.600 645.600 49.500 ;
        RECT 650.400 48.600 651.600 49.500 ;
        RECT 625.800 42.600 627.600 47.700 ;
        RECT 631.800 42.600 633.600 47.700 ;
        RECT 643.800 42.600 645.600 48.600 ;
        RECT 649.800 42.600 651.600 48.600 ;
        RECT 663.000 49.500 668.100 50.400 ;
        RECT 663.000 45.600 664.200 49.500 ;
        RECT 669.000 48.600 670.200 51.900 ;
        RECT 686.400 50.700 687.600 54.900 ;
        RECT 684.000 49.800 687.600 50.700 ;
        RECT 662.400 42.600 664.200 45.600 ;
        RECT 668.700 42.600 670.500 48.600 ;
        RECT 684.000 42.600 685.800 49.800 ;
        RECT 701.400 45.600 702.600 57.900 ;
        RECT 716.100 57.150 717.900 57.900 ;
        RECT 719.850 56.100 721.050 57.900 ;
        RECT 722.100 57.150 723.900 57.900 ;
        RECT 725.100 56.100 726.900 56.850 ;
        RECT 730.950 55.950 736.050 58.050 ;
        RECT 755.100 57.900 756.150 62.100 ;
        RECT 776.850 62.100 778.050 65.400 ;
        RECT 791.400 62.100 792.600 71.400 ;
        RECT 806.400 62.100 807.600 71.400 ;
        RECT 815.400 64.500 816.600 71.400 ;
        RECT 821.700 65.400 823.500 77.400 ;
        RECT 815.400 63.600 821.100 64.500 ;
        RECT 819.150 62.700 821.100 63.600 ;
        RECT 757.950 60.450 760.050 61.050 ;
        RECT 762.000 60.450 766.050 61.050 ;
        RECT 757.950 59.550 766.050 60.450 ;
        RECT 757.950 58.950 760.050 59.550 ;
        RECT 762.000 58.950 766.050 59.550 ;
        RECT 772.950 58.950 775.050 61.050 ;
        RECT 776.850 57.900 777.900 62.100 ;
        RECT 778.950 58.950 781.050 61.050 ;
        RECT 790.950 58.950 793.050 61.050 ;
        RECT 805.950 58.950 808.050 61.050 ;
        RECT 815.100 59.100 816.900 59.850 ;
        RECT 752.100 57.150 753.900 57.900 ;
        RECT 749.100 56.100 750.900 56.850 ;
        RECT 754.950 56.100 756.150 57.900 ;
        RECT 758.100 57.150 759.900 57.900 ;
        RECT 773.100 57.150 774.900 57.900 ;
        RECT 776.850 56.100 778.050 57.900 ;
        RECT 779.100 57.150 780.900 57.900 ;
        RECT 782.100 56.100 783.900 56.850 ;
        RECT 788.100 56.100 789.900 56.850 ;
        RECT 709.950 54.450 712.050 55.050 ;
        RECT 718.950 54.450 721.050 55.050 ;
        RECT 709.950 53.550 721.050 54.450 ;
        RECT 709.950 52.950 712.050 53.550 ;
        RECT 718.950 52.950 721.050 53.550 ;
        RECT 724.950 52.950 727.050 55.050 ;
        RECT 718.950 51.750 720.150 51.900 ;
        RECT 716.400 50.700 720.150 51.750 ;
        RECT 734.400 50.700 735.600 54.900 ;
        RECT 748.950 52.950 751.050 55.050 ;
        RECT 754.950 52.950 757.050 55.050 ;
        RECT 775.950 52.950 778.050 55.050 ;
        RECT 781.950 52.950 784.050 55.050 ;
        RECT 787.950 52.950 790.050 55.050 ;
        RECT 755.850 51.750 757.050 51.900 ;
        RECT 775.950 51.750 777.150 51.900 ;
        RECT 755.850 50.700 759.600 51.750 ;
        RECT 716.400 48.600 717.600 50.700 ;
        RECT 734.400 49.800 738.000 50.700 ;
        RECT 701.400 42.600 703.200 45.600 ;
        RECT 715.800 42.600 717.600 48.600 ;
        RECT 718.800 47.700 726.600 49.050 ;
        RECT 718.800 42.600 720.600 47.700 ;
        RECT 724.800 42.600 726.600 47.700 ;
        RECT 736.200 42.600 738.000 49.800 ;
        RECT 749.400 47.700 757.200 49.050 ;
        RECT 739.950 45.450 742.050 46.050 ;
        RECT 745.950 45.450 748.050 46.200 ;
        RECT 739.950 44.550 748.050 45.450 ;
        RECT 739.950 43.950 742.050 44.550 ;
        RECT 745.950 44.100 748.050 44.550 ;
        RECT 749.400 42.600 751.200 47.700 ;
        RECT 755.400 42.600 757.200 47.700 ;
        RECT 758.400 48.600 759.600 50.700 ;
        RECT 773.400 50.700 777.150 51.750 ;
        RECT 773.400 48.600 774.600 50.700 ;
        RECT 758.400 42.600 760.200 48.600 ;
        RECT 772.800 42.600 774.600 48.600 ;
        RECT 775.800 47.700 783.600 49.050 ;
        RECT 775.800 42.600 777.600 47.700 ;
        RECT 781.800 42.600 783.600 47.700 ;
        RECT 791.400 45.600 792.600 57.900 ;
        RECT 803.100 56.100 804.900 56.850 ;
        RECT 802.950 52.950 805.050 55.050 ;
        RECT 806.400 45.600 807.600 57.900 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 819.150 56.100 820.050 62.700 ;
        RECT 822.000 56.100 823.200 65.400 ;
        RECT 819.150 51.900 819.900 56.100 ;
        RECT 819.150 51.300 820.050 51.900 ;
        RECT 819.150 50.400 821.100 51.300 ;
        RECT 816.000 49.500 821.100 50.400 ;
        RECT 816.000 45.600 817.200 49.500 ;
        RECT 822.000 48.600 823.200 51.900 ;
        RECT 791.400 42.600 793.200 45.600 ;
        RECT 806.400 42.600 808.200 45.600 ;
        RECT 815.400 42.600 817.200 45.600 ;
        RECT 821.700 42.600 823.500 48.600 ;
        RECT 7.800 35.400 9.600 38.400 ;
        RECT 25.800 35.400 27.600 38.400 ;
        RECT 40.800 35.400 42.600 38.400 ;
        RECT 55.800 35.400 57.600 38.400 ;
        RECT 8.400 23.100 9.600 35.400 ;
        RECT 26.400 32.100 27.600 35.400 ;
        RECT 25.950 30.450 28.050 31.050 ;
        RECT 37.950 30.450 40.050 31.050 ;
        RECT 25.950 29.550 40.050 30.450 ;
        RECT 25.950 28.950 28.050 29.550 ;
        RECT 37.950 28.950 40.050 29.550 ;
        RECT 10.950 25.950 13.050 28.050 ;
        RECT 25.950 26.100 27.300 27.900 ;
        RECT 11.100 24.150 12.900 24.900 ;
        RECT 16.950 24.450 21.000 25.050 ;
        RECT 22.950 24.450 25.050 25.050 ;
        RECT 16.950 23.550 25.050 24.450 ;
        RECT 16.950 22.950 21.000 23.550 ;
        RECT 22.950 22.950 25.050 23.550 ;
        RECT 7.950 19.950 10.050 22.050 ;
        RECT 26.100 21.900 27.300 26.100 ;
        RECT 23.100 21.150 24.900 21.900 ;
        RECT 8.400 9.600 9.600 18.900 ;
        RECT 25.950 16.650 27.300 21.900 ;
        RECT 28.950 21.450 31.050 22.050 ;
        RECT 34.950 21.450 37.050 25.050 ;
        RECT 41.400 23.100 42.600 35.400 ;
        RECT 56.400 32.100 57.600 35.400 ;
        RECT 68.400 33.300 70.200 38.400 ;
        RECT 74.400 33.300 76.200 38.400 ;
        RECT 68.400 31.950 76.200 33.300 ;
        RECT 77.400 32.400 79.200 38.400 ;
        RECT 92.400 35.400 94.200 38.400 ;
        RECT 106.800 35.400 108.600 38.400 ;
        RECT 55.950 28.950 61.050 31.050 ;
        RECT 77.400 30.300 78.600 32.400 ;
        RECT 74.850 29.250 78.600 30.300 ;
        RECT 74.850 29.100 76.050 29.250 ;
        RECT 43.950 25.950 46.050 28.050 ;
        RECT 55.950 26.100 57.300 27.900 ;
        RECT 44.100 24.150 45.900 24.900 ;
        RECT 49.950 22.950 55.050 25.050 ;
        RECT 28.950 21.000 37.050 21.450 ;
        RECT 28.950 20.550 36.450 21.000 ;
        RECT 28.950 19.950 31.050 20.550 ;
        RECT 40.950 19.950 43.050 22.050 ;
        RECT 56.100 21.900 57.300 26.100 ;
        RECT 67.950 25.950 70.050 28.050 ;
        RECT 73.950 27.450 76.050 28.050 ;
        RECT 82.950 27.450 85.050 28.050 ;
        RECT 73.950 26.550 85.050 27.450 ;
        RECT 73.950 25.950 76.050 26.550 ;
        RECT 82.950 25.950 85.050 26.550 ;
        RECT 88.950 25.950 91.050 28.050 ;
        RECT 68.100 24.150 69.900 24.900 ;
        RECT 71.100 23.100 72.900 23.850 ;
        RECT 73.950 23.100 75.150 24.900 ;
        RECT 89.100 24.150 90.900 24.900 ;
        RECT 77.100 23.100 78.900 23.850 ;
        RECT 92.400 23.100 93.600 35.400 ;
        RECT 107.400 23.100 108.600 35.400 ;
        RECT 116.400 33.300 118.200 38.400 ;
        RECT 122.400 33.300 124.200 38.400 ;
        RECT 116.400 31.950 124.200 33.300 ;
        RECT 125.400 32.400 127.200 38.400 ;
        RECT 137.400 35.400 139.200 38.400 ;
        RECT 125.400 30.300 126.600 32.400 ;
        RECT 122.850 29.250 126.600 30.300 ;
        RECT 122.850 29.100 124.050 29.250 ;
        RECT 109.950 25.950 112.050 28.050 ;
        RECT 115.950 25.950 118.050 28.050 ;
        RECT 121.950 27.450 124.050 28.050 ;
        RECT 126.000 27.450 130.050 28.050 ;
        RECT 121.950 26.550 130.050 27.450 ;
        RECT 121.950 25.950 124.050 26.550 ;
        RECT 126.000 25.950 130.050 26.550 ;
        RECT 133.950 25.950 136.050 28.050 ;
        RECT 110.100 24.150 111.900 24.900 ;
        RECT 116.100 24.150 117.900 24.900 ;
        RECT 119.100 23.100 120.900 23.850 ;
        RECT 121.950 23.100 123.150 24.900 ;
        RECT 134.100 24.150 135.900 24.900 ;
        RECT 125.100 23.100 126.900 23.850 ;
        RECT 137.400 23.100 138.600 35.400 ;
        RECT 152.100 30.000 153.900 38.400 ;
        RECT 171.000 31.200 172.800 38.400 ;
        RECT 187.200 31.200 189.000 38.400 ;
        RECT 200.400 33.300 202.200 38.400 ;
        RECT 206.400 33.300 208.200 38.400 ;
        RECT 200.400 31.950 208.200 33.300 ;
        RECT 209.400 32.400 211.200 38.400 ;
        RECT 216.150 32.400 217.950 38.400 ;
        RECT 223.950 36.300 225.750 38.400 ;
        RECT 222.000 35.400 225.750 36.300 ;
        RECT 231.750 35.400 233.550 38.400 ;
        RECT 239.550 35.400 241.350 38.400 ;
        RECT 222.000 34.500 223.050 35.400 ;
        RECT 220.950 32.400 223.050 34.500 ;
        RECT 231.750 33.600 232.800 35.400 ;
        RECT 171.000 30.300 174.600 31.200 ;
        RECT 152.100 28.350 156.300 30.000 ;
        RECT 152.100 26.100 153.900 26.850 ;
        RECT 53.100 21.150 54.900 21.900 ;
        RECT 29.100 18.150 30.900 18.900 ;
        RECT 7.800 3.600 9.600 9.600 ;
        RECT 24.600 15.600 27.300 16.650 ;
        RECT 24.600 3.600 26.400 15.600 ;
        RECT 41.400 9.600 42.600 18.900 ;
        RECT 55.950 16.650 57.300 21.900 ;
        RECT 58.950 19.950 64.050 22.050 ;
        RECT 70.950 19.950 73.050 22.050 ;
        RECT 74.100 18.900 75.150 23.100 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 91.950 21.450 94.050 22.050 ;
        RECT 100.950 21.450 103.050 22.050 ;
        RECT 91.950 20.550 103.050 21.450 ;
        RECT 91.950 19.950 94.050 20.550 ;
        RECT 100.950 19.950 103.050 20.550 ;
        RECT 106.950 21.450 109.050 22.050 ;
        RECT 111.000 21.450 115.050 22.050 ;
        RECT 106.950 20.550 115.050 21.450 ;
        RECT 106.950 19.950 109.050 20.550 ;
        RECT 111.000 19.950 115.050 20.550 ;
        RECT 118.950 19.950 121.050 22.050 ;
        RECT 122.100 18.900 123.150 23.100 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 136.950 21.450 139.050 22.050 ;
        RECT 141.000 21.450 145.050 22.050 ;
        RECT 136.950 20.550 145.050 21.450 ;
        RECT 136.950 19.950 139.050 20.550 ;
        RECT 141.000 19.950 145.050 20.550 ;
        RECT 148.950 19.950 151.050 22.050 ;
        RECT 155.400 20.100 156.300 28.350 ;
        RECT 173.400 26.100 174.600 30.300 ;
        RECT 185.400 30.300 189.000 31.200 ;
        RECT 209.400 30.300 210.600 32.400 ;
        RECT 185.400 26.100 186.600 30.300 ;
        RECT 206.850 29.250 210.600 30.300 ;
        RECT 206.850 29.100 208.050 29.250 ;
        RECT 199.950 25.950 202.050 28.050 ;
        RECT 205.950 27.450 208.050 28.050 ;
        RECT 210.000 27.450 214.050 28.050 ;
        RECT 205.950 26.550 214.050 27.450 ;
        RECT 205.950 25.950 208.050 26.550 ;
        RECT 210.000 25.950 214.050 26.550 ;
        RECT 172.950 24.450 175.050 25.050 ;
        RECT 177.000 24.450 181.050 25.050 ;
        RECT 172.950 23.550 181.050 24.450 ;
        RECT 172.950 22.950 175.050 23.550 ;
        RECT 177.000 22.950 181.050 23.550 ;
        RECT 184.950 22.950 190.050 25.050 ;
        RECT 200.100 24.150 201.900 24.900 ;
        RECT 203.100 23.100 204.900 23.850 ;
        RECT 205.950 23.100 207.150 24.900 ;
        RECT 209.100 23.100 210.900 23.850 ;
        RECT 170.100 20.100 171.900 20.850 ;
        RECT 59.100 18.150 60.900 18.900 ;
        RECT 40.800 3.600 42.600 9.600 ;
        RECT 54.600 15.600 57.300 16.650 ;
        RECT 73.950 15.600 75.150 18.900 ;
        RECT 54.600 3.600 56.400 15.600 ;
        RECT 73.500 3.600 75.300 15.600 ;
        RECT 92.400 9.600 93.600 18.900 ;
        RECT 107.400 9.600 108.600 18.900 ;
        RECT 121.950 15.600 123.150 18.900 ;
        RECT 92.400 3.600 94.200 9.600 ;
        RECT 106.800 3.600 108.600 9.600 ;
        RECT 121.500 3.600 123.300 15.600 ;
        RECT 137.400 9.600 138.600 18.900 ;
        RECT 149.100 18.150 150.900 18.900 ;
        RECT 154.950 18.450 157.050 19.050 ;
        RECT 159.000 18.450 163.050 19.050 ;
        RECT 146.100 17.100 147.900 17.850 ;
        RECT 154.950 17.550 163.050 18.450 ;
        RECT 154.950 16.950 157.050 17.550 ;
        RECT 159.000 16.950 163.050 17.550 ;
        RECT 169.950 16.950 172.050 19.050 ;
        RECT 145.950 13.950 148.050 16.050 ;
        RECT 155.400 10.800 156.300 15.900 ;
        RECT 149.700 9.900 156.300 10.800 ;
        RECT 149.700 9.600 151.200 9.900 ;
        RECT 137.400 3.600 139.200 9.600 ;
        RECT 149.400 3.600 151.200 9.600 ;
        RECT 155.400 9.600 156.300 9.900 ;
        RECT 173.400 9.600 174.600 21.900 ;
        RECT 176.100 20.100 177.900 20.850 ;
        RECT 182.100 20.100 183.900 20.850 ;
        RECT 175.950 16.950 178.050 19.050 ;
        RECT 181.950 16.950 184.050 19.050 ;
        RECT 155.400 3.600 157.200 9.600 ;
        RECT 172.800 3.600 174.600 9.600 ;
        RECT 185.400 9.600 186.600 21.900 ;
        RECT 188.100 20.100 189.900 20.850 ;
        RECT 202.950 19.950 205.050 22.050 ;
        RECT 187.950 16.950 190.050 19.050 ;
        RECT 206.100 18.900 207.150 23.100 ;
        RECT 208.950 19.950 211.050 22.050 ;
        RECT 205.950 15.600 207.150 18.900 ;
        RECT 216.150 17.700 217.050 32.400 ;
        RECT 224.550 31.800 226.350 33.600 ;
        RECT 227.850 32.550 232.800 33.600 ;
        RECT 240.300 34.500 241.350 35.400 ;
        RECT 240.300 33.300 244.050 34.500 ;
        RECT 227.850 31.800 229.650 32.550 ;
        RECT 241.950 32.400 244.050 33.300 ;
        RECT 247.650 32.400 249.450 38.400 ;
        RECT 224.850 28.800 225.900 31.800 ;
        RECT 219.000 27.600 236.850 28.800 ;
        RECT 248.250 28.050 249.450 32.400 ;
        RECT 219.000 26.850 219.900 27.600 ;
        RECT 224.100 27.000 225.900 27.600 ;
        RECT 235.050 27.000 236.850 27.600 ;
        RECT 218.100 25.050 219.900 26.850 ;
        RECT 235.050 26.100 235.950 27.000 ;
        RECT 243.150 26.250 243.900 28.050 ;
        RECT 244.950 25.950 247.050 28.050 ;
        RECT 248.100 25.950 249.450 28.050 ;
        RECT 221.100 22.800 222.900 23.400 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 221.100 21.600 225.900 22.800 ;
        RECT 226.950 19.950 229.050 22.050 ;
        RECT 225.450 17.700 227.250 18.000 ;
        RECT 216.150 17.100 227.250 17.700 ;
        RECT 216.150 16.500 233.850 17.100 ;
        RECT 216.150 15.600 217.050 16.500 ;
        RECT 225.450 16.200 233.850 16.500 ;
        RECT 185.400 3.600 187.200 9.600 ;
        RECT 205.500 3.600 207.300 15.600 ;
        RECT 216.150 3.600 217.950 15.600 ;
        RECT 230.250 14.700 232.050 15.300 ;
        RECT 224.550 13.500 232.050 14.700 ;
        RECT 232.950 14.100 233.850 16.200 ;
        RECT 235.050 16.200 235.950 21.900 ;
        RECT 245.250 17.400 247.050 19.200 ;
        RECT 241.950 16.200 246.150 17.400 ;
        RECT 235.050 15.300 241.050 16.200 ;
        RECT 241.950 15.300 244.050 16.200 ;
        RECT 248.250 15.600 249.450 25.950 ;
        RECT 240.150 14.400 241.050 15.300 ;
        RECT 237.450 14.100 239.250 14.400 ;
        RECT 224.550 12.600 225.750 13.500 ;
        RECT 232.950 13.200 239.250 14.100 ;
        RECT 237.450 12.600 239.250 13.200 ;
        RECT 240.150 12.600 242.850 14.400 ;
        RECT 220.950 10.500 225.750 12.600 ;
        RECT 228.450 11.550 230.250 12.300 ;
        RECT 233.250 11.550 235.050 12.300 ;
        RECT 228.450 10.500 235.050 11.550 ;
        RECT 224.550 9.600 225.750 10.500 ;
        RECT 224.550 3.600 226.350 9.600 ;
        RECT 232.350 3.600 234.150 10.500 ;
        RECT 240.150 9.600 244.050 11.700 ;
        RECT 240.150 3.600 241.950 9.600 ;
        RECT 247.650 3.600 249.450 15.600 ;
        RECT 252.150 32.400 253.950 38.400 ;
        RECT 259.950 36.300 261.750 38.400 ;
        RECT 258.000 35.400 261.750 36.300 ;
        RECT 267.750 35.400 269.550 38.400 ;
        RECT 275.550 35.400 277.350 38.400 ;
        RECT 258.000 34.500 259.050 35.400 ;
        RECT 256.950 32.400 259.050 34.500 ;
        RECT 267.750 33.600 268.800 35.400 ;
        RECT 252.150 17.700 253.050 32.400 ;
        RECT 260.550 31.800 262.350 33.600 ;
        RECT 263.850 32.550 268.800 33.600 ;
        RECT 276.300 34.500 277.350 35.400 ;
        RECT 276.300 33.300 280.050 34.500 ;
        RECT 263.850 31.800 265.650 32.550 ;
        RECT 277.950 32.400 280.050 33.300 ;
        RECT 283.650 32.400 285.450 38.400 ;
        RECT 260.850 28.800 261.900 31.800 ;
        RECT 255.000 27.600 272.850 28.800 ;
        RECT 284.250 28.050 285.450 32.400 ;
        RECT 300.000 32.400 301.800 38.400 ;
        RECT 319.800 35.400 321.600 38.400 ;
        RECT 300.000 29.100 301.050 32.400 ;
        RECT 320.400 32.100 321.600 35.400 ;
        RECT 326.550 32.400 328.350 38.400 ;
        RECT 334.650 35.400 336.450 38.400 ;
        RECT 342.450 35.400 344.250 38.400 ;
        RECT 350.250 36.300 352.050 38.400 ;
        RECT 350.250 35.400 354.000 36.300 ;
        RECT 334.650 34.500 335.700 35.400 ;
        RECT 331.950 33.300 335.700 34.500 ;
        RECT 343.200 33.600 344.250 35.400 ;
        RECT 352.950 34.500 354.000 35.400 ;
        RECT 331.950 32.400 334.050 33.300 ;
        RECT 343.200 32.550 348.150 33.600 ;
        RECT 313.950 30.450 318.000 31.050 ;
        RECT 319.950 30.450 322.050 31.050 ;
        RECT 313.950 29.550 322.050 30.450 ;
        RECT 313.950 28.950 318.000 29.550 ;
        RECT 319.950 28.950 322.050 29.550 ;
        RECT 326.550 28.050 327.750 32.400 ;
        RECT 346.350 31.800 348.150 32.550 ;
        RECT 349.650 31.800 351.450 33.600 ;
        RECT 352.950 32.400 355.050 34.500 ;
        RECT 358.050 32.400 359.850 38.400 ;
        RECT 372.000 34.050 373.800 38.400 ;
        RECT 350.100 28.800 351.150 31.800 ;
        RECT 255.000 26.850 255.900 27.600 ;
        RECT 260.100 27.000 261.900 27.600 ;
        RECT 271.050 27.000 272.850 27.600 ;
        RECT 254.100 25.050 255.900 26.850 ;
        RECT 271.050 26.100 271.950 27.000 ;
        RECT 279.150 26.250 279.900 28.050 ;
        RECT 280.950 25.950 283.050 28.050 ;
        RECT 284.100 25.950 285.450 28.050 ;
        RECT 292.950 25.950 295.050 28.050 ;
        RECT 298.950 25.950 301.050 28.050 ;
        RECT 304.950 25.950 307.050 28.050 ;
        RECT 319.950 26.100 321.300 27.900 ;
        RECT 257.100 22.800 258.900 23.400 ;
        RECT 268.950 22.950 271.050 25.050 ;
        RECT 257.100 21.600 261.900 22.800 ;
        RECT 262.950 19.950 265.050 22.050 ;
        RECT 261.450 17.700 263.250 18.000 ;
        RECT 252.150 17.100 263.250 17.700 ;
        RECT 252.150 16.500 269.850 17.100 ;
        RECT 252.150 15.600 253.050 16.500 ;
        RECT 261.450 16.200 269.850 16.500 ;
        RECT 252.150 3.600 253.950 15.600 ;
        RECT 266.250 14.700 268.050 15.300 ;
        RECT 260.550 13.500 268.050 14.700 ;
        RECT 268.950 14.100 269.850 16.200 ;
        RECT 271.050 16.200 271.950 21.900 ;
        RECT 281.250 17.400 283.050 19.200 ;
        RECT 277.950 16.200 282.150 17.400 ;
        RECT 271.050 15.300 277.050 16.200 ;
        RECT 277.950 15.300 280.050 16.200 ;
        RECT 284.250 15.600 285.450 25.950 ;
        RECT 293.100 24.150 294.900 24.900 ;
        RECT 296.250 23.100 298.050 23.850 ;
        RECT 298.950 23.100 299.850 24.900 ;
        RECT 304.950 24.150 306.750 24.900 ;
        RECT 301.950 23.100 303.750 23.850 ;
        RECT 295.950 19.950 298.050 22.050 ;
        RECT 299.100 18.900 299.850 23.100 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 301.950 19.950 304.050 22.050 ;
        RECT 320.100 21.900 321.300 26.100 ;
        RECT 326.550 25.950 327.900 28.050 ;
        RECT 328.950 25.950 331.050 28.050 ;
        RECT 332.100 26.250 332.850 28.050 ;
        RECT 339.150 27.600 357.000 28.800 ;
        RECT 339.150 27.000 340.950 27.600 ;
        RECT 350.100 27.000 351.900 27.600 ;
        RECT 340.050 26.100 340.950 27.000 ;
        RECT 356.100 26.850 357.000 27.600 ;
        RECT 317.100 21.150 318.900 21.900 ;
        RECT 298.950 17.400 299.850 18.900 ;
        RECT 295.800 16.500 299.850 17.400 ;
        RECT 319.950 16.650 321.300 21.900 ;
        RECT 322.950 19.950 325.050 22.050 ;
        RECT 323.100 18.150 324.900 18.900 ;
        RECT 276.150 14.400 277.050 15.300 ;
        RECT 273.450 14.100 275.250 14.400 ;
        RECT 260.550 12.600 261.750 13.500 ;
        RECT 268.950 13.200 275.250 14.100 ;
        RECT 273.450 12.600 275.250 13.200 ;
        RECT 276.150 12.600 278.850 14.400 ;
        RECT 256.950 10.500 261.750 12.600 ;
        RECT 264.450 11.550 266.250 12.300 ;
        RECT 269.250 11.550 271.050 12.300 ;
        RECT 264.450 10.500 271.050 11.550 ;
        RECT 260.550 9.600 261.750 10.500 ;
        RECT 260.550 3.600 262.350 9.600 ;
        RECT 268.350 3.600 270.150 10.500 ;
        RECT 276.150 9.600 280.050 11.700 ;
        RECT 276.150 3.600 277.950 9.600 ;
        RECT 283.650 3.600 285.450 15.600 ;
        RECT 292.800 4.500 294.600 15.600 ;
        RECT 295.800 5.400 297.600 16.500 ;
        RECT 318.600 15.600 321.300 16.650 ;
        RECT 326.550 15.600 327.750 25.950 ;
        RECT 356.100 25.050 357.900 26.850 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 353.100 22.800 354.900 23.400 ;
        RECT 328.950 17.400 330.750 19.200 ;
        RECT 329.850 16.200 334.050 17.400 ;
        RECT 340.050 16.200 340.950 21.900 ;
        RECT 346.950 19.950 349.050 22.050 ;
        RECT 350.100 21.600 354.900 22.800 ;
        RECT 348.750 17.700 350.550 18.000 ;
        RECT 358.950 17.700 359.850 32.400 ;
        RECT 368.400 32.400 373.800 34.050 ;
        RECT 381.150 32.400 382.950 38.400 ;
        RECT 388.950 36.300 390.750 38.400 ;
        RECT 387.000 35.400 390.750 36.300 ;
        RECT 396.750 35.400 398.550 38.400 ;
        RECT 404.550 35.400 406.350 38.400 ;
        RECT 387.000 34.500 388.050 35.400 ;
        RECT 385.950 32.400 388.050 34.500 ;
        RECT 396.750 33.600 397.800 35.400 ;
        RECT 368.400 29.100 369.300 32.400 ;
        RECT 361.950 27.450 366.000 28.050 ;
        RECT 367.950 27.450 370.050 28.050 ;
        RECT 361.950 26.550 370.050 27.450 ;
        RECT 361.950 25.950 366.000 26.550 ;
        RECT 367.950 25.950 370.050 26.550 ;
        RECT 373.950 25.950 376.050 28.050 ;
        RECT 348.750 17.100 359.850 17.700 ;
        RECT 298.800 14.400 306.600 15.300 ;
        RECT 298.800 4.500 300.600 14.400 ;
        RECT 292.800 3.600 300.600 4.500 ;
        RECT 304.800 3.600 306.600 14.400 ;
        RECT 318.600 3.600 320.400 15.600 ;
        RECT 326.550 3.600 328.350 15.600 ;
        RECT 331.950 15.300 334.050 16.200 ;
        RECT 334.950 15.300 340.950 16.200 ;
        RECT 342.150 16.500 359.850 17.100 ;
        RECT 342.150 16.200 350.550 16.500 ;
        RECT 334.950 14.400 335.850 15.300 ;
        RECT 333.150 12.600 335.850 14.400 ;
        RECT 336.750 14.100 338.550 14.400 ;
        RECT 342.150 14.100 343.050 16.200 ;
        RECT 358.950 15.600 359.850 16.500 ;
        RECT 368.400 15.600 369.300 24.900 ;
        RECT 374.100 24.150 375.900 24.900 ;
        RECT 371.100 23.100 372.900 23.850 ;
        RECT 377.100 23.100 378.900 23.850 ;
        RECT 370.950 19.950 373.050 22.050 ;
        RECT 376.950 19.950 379.050 22.050 ;
        RECT 381.150 17.700 382.050 32.400 ;
        RECT 389.550 31.800 391.350 33.600 ;
        RECT 392.850 32.550 397.800 33.600 ;
        RECT 405.300 34.500 406.350 35.400 ;
        RECT 405.300 33.300 409.050 34.500 ;
        RECT 392.850 31.800 394.650 32.550 ;
        RECT 406.950 32.400 409.050 33.300 ;
        RECT 412.650 32.400 414.450 38.400 ;
        RECT 424.500 32.400 426.300 38.400 ;
        RECT 430.800 35.400 432.600 38.400 ;
        RECT 389.850 28.800 390.900 31.800 ;
        RECT 384.000 27.600 401.850 28.800 ;
        RECT 413.250 28.050 414.450 32.400 ;
        RECT 424.800 29.100 426.000 32.400 ;
        RECT 430.800 31.500 432.000 35.400 ;
        RECT 442.800 32.400 444.600 38.400 ;
        RECT 426.900 30.600 432.000 31.500 ;
        RECT 426.900 29.700 428.850 30.600 ;
        RECT 427.950 29.100 428.850 29.700 ;
        RECT 443.400 30.300 444.600 32.400 ;
        RECT 445.800 33.300 447.600 38.400 ;
        RECT 451.800 33.300 453.600 38.400 ;
        RECT 445.800 31.950 453.600 33.300 ;
        RECT 460.500 32.400 462.300 38.400 ;
        RECT 466.800 35.400 468.600 38.400 ;
        RECT 443.400 29.250 447.150 30.300 ;
        RECT 445.950 29.100 447.150 29.250 ;
        RECT 460.800 29.100 462.000 32.400 ;
        RECT 466.800 31.500 468.000 35.400 ;
        RECT 478.800 32.400 480.600 38.400 ;
        RECT 462.900 30.600 468.000 31.500 ;
        RECT 462.900 29.700 464.850 30.600 ;
        RECT 463.950 29.100 464.850 29.700 ;
        RECT 479.400 30.300 480.600 32.400 ;
        RECT 481.800 33.300 483.600 38.400 ;
        RECT 487.800 33.300 489.600 38.400 ;
        RECT 497.400 35.400 499.200 38.400 ;
        RECT 481.800 31.950 489.600 33.300 ;
        RECT 498.000 31.500 499.200 35.400 ;
        RECT 503.700 32.400 505.500 38.400 ;
        RECT 512.400 35.400 514.200 38.400 ;
        RECT 498.000 30.600 503.100 31.500 ;
        RECT 479.400 29.250 483.150 30.300 ;
        RECT 481.950 29.100 483.150 29.250 ;
        RECT 501.150 29.700 503.100 30.600 ;
        RECT 501.150 29.100 502.050 29.700 ;
        RECT 504.000 29.100 505.200 32.400 ;
        RECT 513.000 31.500 514.200 35.400 ;
        RECT 518.700 32.400 520.500 38.400 ;
        RECT 529.800 35.400 531.600 38.400 ;
        RECT 513.000 30.600 518.100 31.500 ;
        RECT 516.150 29.700 518.100 30.600 ;
        RECT 516.150 29.100 517.050 29.700 ;
        RECT 519.000 29.100 520.200 32.400 ;
        RECT 384.000 26.850 384.900 27.600 ;
        RECT 389.100 27.000 390.900 27.600 ;
        RECT 400.050 27.000 401.850 27.600 ;
        RECT 383.100 25.050 384.900 26.850 ;
        RECT 400.050 26.100 400.950 27.000 ;
        RECT 408.150 26.250 408.900 28.050 ;
        RECT 409.950 25.950 412.050 28.050 ;
        RECT 413.100 25.950 414.450 28.050 ;
        RECT 386.100 22.800 387.900 23.400 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 386.100 21.600 390.900 22.800 ;
        RECT 391.950 19.950 394.050 22.050 ;
        RECT 390.450 17.700 392.250 18.000 ;
        RECT 381.150 17.100 392.250 17.700 ;
        RECT 381.150 16.500 398.850 17.100 ;
        RECT 381.150 15.600 382.050 16.500 ;
        RECT 390.450 16.200 398.850 16.500 ;
        RECT 336.750 13.200 343.050 14.100 ;
        RECT 343.950 14.700 345.750 15.300 ;
        RECT 343.950 13.500 351.450 14.700 ;
        RECT 336.750 12.600 338.550 13.200 ;
        RECT 350.250 12.600 351.450 13.500 ;
        RECT 331.950 9.600 335.850 11.700 ;
        RECT 340.950 11.550 342.750 12.300 ;
        RECT 345.750 11.550 347.550 12.300 ;
        RECT 340.950 10.500 347.550 11.550 ;
        RECT 350.250 10.500 355.050 12.600 ;
        RECT 334.050 3.600 335.850 9.600 ;
        RECT 341.850 3.600 343.650 10.500 ;
        RECT 350.250 9.600 351.450 10.500 ;
        RECT 349.650 3.600 351.450 9.600 ;
        RECT 358.050 3.600 359.850 15.600 ;
        RECT 367.800 3.600 369.600 15.600 ;
        RECT 370.800 14.700 378.600 15.600 ;
        RECT 370.800 3.600 372.600 14.700 ;
        RECT 376.800 3.600 378.600 14.700 ;
        RECT 381.150 3.600 382.950 15.600 ;
        RECT 395.250 14.700 397.050 15.300 ;
        RECT 389.550 13.500 397.050 14.700 ;
        RECT 397.950 14.100 398.850 16.200 ;
        RECT 400.050 16.200 400.950 21.900 ;
        RECT 410.250 17.400 412.050 19.200 ;
        RECT 406.950 16.200 411.150 17.400 ;
        RECT 400.050 15.300 406.050 16.200 ;
        RECT 406.950 15.300 409.050 16.200 ;
        RECT 413.250 15.600 414.450 25.950 ;
        RECT 428.100 24.900 428.850 29.100 ;
        RECT 445.950 25.950 448.050 28.050 ;
        RECT 451.950 25.950 454.050 28.050 ;
        RECT 424.800 15.600 426.000 24.900 ;
        RECT 427.950 18.300 428.850 24.900 ;
        RECT 430.950 24.450 433.050 25.050 ;
        RECT 435.000 24.450 439.050 25.050 ;
        RECT 464.100 24.900 464.850 29.100 ;
        RECT 481.950 25.950 484.050 28.050 ;
        RECT 487.950 25.950 490.050 28.050 ;
        RECT 430.950 23.550 439.050 24.450 ;
        RECT 430.950 22.950 433.050 23.550 ;
        RECT 435.000 22.950 439.050 23.550 ;
        RECT 443.100 23.100 444.900 23.850 ;
        RECT 446.850 23.100 448.050 24.900 ;
        RECT 452.100 24.150 453.900 24.900 ;
        RECT 449.100 23.100 450.900 23.850 ;
        RECT 431.100 21.150 432.900 21.900 ;
        RECT 442.950 19.950 445.050 22.050 ;
        RECT 426.900 17.400 428.850 18.300 ;
        RECT 446.850 18.900 447.900 23.100 ;
        RECT 448.950 19.950 451.050 22.050 ;
        RECT 426.900 16.500 432.600 17.400 ;
        RECT 405.150 14.400 406.050 15.300 ;
        RECT 402.450 14.100 404.250 14.400 ;
        RECT 389.550 12.600 390.750 13.500 ;
        RECT 397.950 13.200 404.250 14.100 ;
        RECT 402.450 12.600 404.250 13.200 ;
        RECT 405.150 12.600 407.850 14.400 ;
        RECT 385.950 10.500 390.750 12.600 ;
        RECT 393.450 11.550 395.250 12.300 ;
        RECT 398.250 11.550 400.050 12.300 ;
        RECT 393.450 10.500 400.050 11.550 ;
        RECT 389.550 9.600 390.750 10.500 ;
        RECT 389.550 3.600 391.350 9.600 ;
        RECT 397.350 3.600 399.150 10.500 ;
        RECT 405.150 9.600 409.050 11.700 ;
        RECT 405.150 3.600 406.950 9.600 ;
        RECT 412.650 3.600 414.450 15.600 ;
        RECT 424.500 3.600 426.300 15.600 ;
        RECT 431.400 9.600 432.600 16.500 ;
        RECT 446.850 15.600 448.050 18.900 ;
        RECT 460.800 15.600 462.000 24.900 ;
        RECT 463.950 18.300 464.850 24.900 ;
        RECT 466.950 24.450 469.050 25.050 ;
        RECT 471.000 24.450 475.050 25.050 ;
        RECT 466.950 23.550 475.050 24.450 ;
        RECT 466.950 22.950 469.050 23.550 ;
        RECT 471.000 22.950 475.050 23.550 ;
        RECT 479.100 23.100 480.900 23.850 ;
        RECT 482.850 23.100 484.050 24.900 ;
        RECT 488.100 24.150 489.900 24.900 ;
        RECT 485.100 23.100 486.900 23.850 ;
        RECT 467.100 21.150 468.900 21.900 ;
        RECT 478.950 19.950 481.050 22.050 ;
        RECT 462.900 17.400 464.850 18.300 ;
        RECT 482.850 18.900 483.900 23.100 ;
        RECT 493.950 22.950 499.050 25.050 ;
        RECT 501.150 24.900 501.900 29.100 ;
        RECT 484.950 19.950 487.050 22.050 ;
        RECT 497.100 21.150 498.900 21.900 ;
        RECT 462.900 16.500 468.600 17.400 ;
        RECT 430.800 3.600 432.600 9.600 ;
        RECT 446.700 3.600 448.500 15.600 ;
        RECT 460.500 3.600 462.300 15.600 ;
        RECT 467.400 9.600 468.600 16.500 ;
        RECT 482.850 15.600 484.050 18.900 ;
        RECT 501.150 18.300 502.050 24.900 ;
        RECT 501.150 17.400 503.100 18.300 ;
        RECT 497.400 16.500 503.100 17.400 ;
        RECT 466.800 3.600 468.600 9.600 ;
        RECT 482.700 3.600 484.500 15.600 ;
        RECT 497.400 9.600 498.600 16.500 ;
        RECT 504.000 15.600 505.200 24.900 ;
        RECT 508.950 22.950 514.050 25.050 ;
        RECT 516.150 24.900 516.900 29.100 ;
        RECT 512.100 21.150 513.900 21.900 ;
        RECT 516.150 18.300 517.050 24.900 ;
        RECT 516.150 17.400 518.100 18.300 ;
        RECT 512.400 16.500 518.100 17.400 ;
        RECT 497.400 3.600 499.200 9.600 ;
        RECT 503.700 3.600 505.500 15.600 ;
        RECT 512.400 9.600 513.600 16.500 ;
        RECT 519.000 15.600 520.200 24.900 ;
        RECT 530.400 23.100 531.600 35.400 ;
        RECT 542.400 35.400 544.200 38.400 ;
        RECT 542.400 32.100 543.600 35.400 ;
        RECT 559.800 32.400 561.600 38.400 ;
        RECT 538.950 31.050 541.050 31.200 ;
        RECT 538.950 29.100 544.050 31.050 ;
        RECT 560.400 30.300 561.600 32.400 ;
        RECT 562.800 33.300 564.600 38.400 ;
        RECT 568.800 33.300 570.600 38.400 ;
        RECT 562.800 31.950 570.600 33.300 ;
        RECT 580.200 31.200 582.000 38.400 ;
        RECT 578.400 30.300 582.000 31.200 ;
        RECT 587.550 32.400 589.350 38.400 ;
        RECT 595.650 35.400 597.450 38.400 ;
        RECT 603.450 35.400 605.250 38.400 ;
        RECT 611.250 36.300 613.050 38.400 ;
        RECT 611.250 35.400 615.000 36.300 ;
        RECT 595.650 34.500 596.700 35.400 ;
        RECT 592.950 33.300 596.700 34.500 ;
        RECT 604.200 33.600 605.250 35.400 ;
        RECT 613.950 34.500 615.000 35.400 ;
        RECT 592.950 32.400 595.050 33.300 ;
        RECT 604.200 32.550 609.150 33.600 ;
        RECT 560.400 29.250 564.150 30.300 ;
        RECT 562.950 29.100 564.150 29.250 ;
        RECT 539.550 28.950 544.050 29.100 ;
        RECT 542.700 26.100 544.050 27.900 ;
        RECT 550.950 27.450 553.050 28.050 ;
        RECT 562.950 27.450 565.050 28.050 ;
        RECT 550.950 26.550 565.050 27.450 ;
        RECT 533.100 24.150 534.900 24.900 ;
        RECT 529.950 19.950 532.050 22.050 ;
        RECT 538.950 19.950 541.050 22.050 ;
        RECT 542.700 21.900 543.900 26.100 ;
        RECT 550.950 25.950 553.050 26.550 ;
        RECT 562.950 25.950 565.050 26.550 ;
        RECT 568.950 25.950 571.050 28.050 ;
        RECT 578.400 26.100 579.600 30.300 ;
        RECT 587.550 28.050 588.750 32.400 ;
        RECT 607.350 31.800 609.150 32.550 ;
        RECT 610.650 31.800 612.450 33.600 ;
        RECT 613.950 32.400 616.050 34.500 ;
        RECT 619.050 32.400 620.850 38.400 ;
        RECT 611.100 28.800 612.150 31.800 ;
        RECT 587.550 25.950 588.900 28.050 ;
        RECT 589.950 25.950 592.050 28.050 ;
        RECT 593.100 26.250 593.850 28.050 ;
        RECT 600.150 27.600 618.000 28.800 ;
        RECT 600.150 27.000 601.950 27.600 ;
        RECT 611.100 27.000 612.900 27.600 ;
        RECT 601.050 26.100 601.950 27.000 ;
        RECT 617.100 26.850 618.000 27.600 ;
        RECT 544.950 22.950 547.050 25.050 ;
        RECT 560.100 23.100 561.900 23.850 ;
        RECT 563.850 23.100 565.050 24.900 ;
        RECT 569.100 24.150 570.900 24.900 ;
        RECT 566.100 23.100 567.900 23.850 ;
        RECT 512.400 3.600 514.200 9.600 ;
        RECT 518.700 3.600 520.500 15.600 ;
        RECT 530.400 9.600 531.600 18.900 ;
        RECT 539.100 18.150 540.900 18.900 ;
        RECT 542.700 16.650 544.050 21.900 ;
        RECT 545.100 21.150 546.900 21.900 ;
        RECT 559.950 19.950 562.050 22.050 ;
        RECT 563.850 18.900 564.900 23.100 ;
        RECT 574.950 22.950 580.050 25.050 ;
        RECT 565.950 19.950 568.050 22.050 ;
        RECT 575.100 20.100 576.900 20.850 ;
        RECT 542.700 15.600 545.400 16.650 ;
        RECT 563.850 15.600 565.050 18.900 ;
        RECT 574.950 16.950 577.050 19.050 ;
        RECT 529.800 3.600 531.600 9.600 ;
        RECT 543.600 3.600 545.400 15.600 ;
        RECT 563.700 3.600 565.500 15.600 ;
        RECT 578.400 9.600 579.600 21.900 ;
        RECT 581.100 20.100 582.900 20.850 ;
        RECT 580.950 16.950 583.050 19.050 ;
        RECT 587.550 15.600 588.750 25.950 ;
        RECT 617.100 25.050 618.900 26.850 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 614.100 22.800 615.900 23.400 ;
        RECT 589.950 17.400 591.750 19.200 ;
        RECT 590.850 16.200 595.050 17.400 ;
        RECT 601.050 16.200 601.950 21.900 ;
        RECT 607.950 19.950 610.050 22.050 ;
        RECT 611.100 21.600 615.900 22.800 ;
        RECT 609.750 17.700 611.550 18.000 ;
        RECT 619.950 17.700 620.850 32.400 ;
        RECT 634.200 31.200 636.000 38.400 ;
        RECT 632.400 30.300 636.000 31.200 ;
        RECT 651.000 31.200 652.800 38.400 ;
        RECT 659.550 32.400 661.350 38.400 ;
        RECT 667.650 35.400 669.450 38.400 ;
        RECT 675.450 35.400 677.250 38.400 ;
        RECT 683.250 36.300 685.050 38.400 ;
        RECT 683.250 35.400 687.000 36.300 ;
        RECT 667.650 34.500 668.700 35.400 ;
        RECT 664.950 33.300 668.700 34.500 ;
        RECT 676.200 33.600 677.250 35.400 ;
        RECT 685.950 34.500 687.000 35.400 ;
        RECT 664.950 32.400 667.050 33.300 ;
        RECT 676.200 32.550 681.150 33.600 ;
        RECT 651.000 30.300 654.600 31.200 ;
        RECT 632.400 26.100 633.600 30.300 ;
        RECT 653.400 26.100 654.600 30.300 ;
        RECT 659.550 28.050 660.750 32.400 ;
        RECT 679.350 31.800 681.150 32.550 ;
        RECT 682.650 31.800 684.450 33.600 ;
        RECT 685.950 32.400 688.050 34.500 ;
        RECT 691.050 32.400 692.850 38.400 ;
        RECT 700.800 32.400 702.600 38.400 ;
        RECT 683.100 28.800 684.150 31.800 ;
        RECT 659.550 25.950 660.900 28.050 ;
        RECT 661.950 25.950 664.050 28.050 ;
        RECT 665.100 26.250 665.850 28.050 ;
        RECT 672.150 27.600 690.000 28.800 ;
        RECT 672.150 27.000 673.950 27.600 ;
        RECT 683.100 27.000 684.900 27.600 ;
        RECT 673.050 26.100 673.950 27.000 ;
        RECT 689.100 26.850 690.000 27.600 ;
        RECT 622.950 24.450 625.050 25.050 ;
        RECT 631.950 24.450 634.050 25.050 ;
        RECT 622.950 23.550 634.050 24.450 ;
        RECT 622.950 22.950 625.050 23.550 ;
        RECT 631.950 22.950 634.050 23.550 ;
        RECT 646.950 24.450 651.000 25.050 ;
        RECT 652.950 24.450 655.050 25.050 ;
        RECT 646.950 23.550 655.050 24.450 ;
        RECT 646.950 22.950 651.000 23.550 ;
        RECT 652.950 22.950 655.050 23.550 ;
        RECT 629.100 20.100 630.900 20.850 ;
        RECT 609.750 17.100 620.850 17.700 ;
        RECT 578.400 3.600 580.200 9.600 ;
        RECT 587.550 3.600 589.350 15.600 ;
        RECT 592.950 15.300 595.050 16.200 ;
        RECT 595.950 15.300 601.950 16.200 ;
        RECT 603.150 16.500 620.850 17.100 ;
        RECT 625.950 16.950 631.050 19.050 ;
        RECT 603.150 16.200 611.550 16.500 ;
        RECT 595.950 14.400 596.850 15.300 ;
        RECT 594.150 12.600 596.850 14.400 ;
        RECT 597.750 14.100 599.550 14.400 ;
        RECT 603.150 14.100 604.050 16.200 ;
        RECT 619.950 15.600 620.850 16.500 ;
        RECT 597.750 13.200 604.050 14.100 ;
        RECT 604.950 14.700 606.750 15.300 ;
        RECT 604.950 13.500 612.450 14.700 ;
        RECT 597.750 12.600 599.550 13.200 ;
        RECT 611.250 12.600 612.450 13.500 ;
        RECT 592.950 9.600 596.850 11.700 ;
        RECT 601.950 11.550 603.750 12.300 ;
        RECT 606.750 11.550 608.550 12.300 ;
        RECT 601.950 10.500 608.550 11.550 ;
        RECT 611.250 10.500 616.050 12.600 ;
        RECT 595.050 3.600 596.850 9.600 ;
        RECT 602.850 3.600 604.650 10.500 ;
        RECT 611.250 9.600 612.450 10.500 ;
        RECT 610.650 3.600 612.450 9.600 ;
        RECT 619.050 3.600 620.850 15.600 ;
        RECT 632.400 9.600 633.600 21.900 ;
        RECT 635.100 20.100 636.900 20.850 ;
        RECT 650.100 20.100 651.900 20.850 ;
        RECT 634.950 16.950 637.050 19.050 ;
        RECT 649.950 16.950 652.050 19.050 ;
        RECT 653.400 9.600 654.600 21.900 ;
        RECT 656.100 20.100 657.900 20.850 ;
        RECT 655.950 16.950 658.050 19.050 ;
        RECT 632.400 3.600 634.200 9.600 ;
        RECT 652.800 3.600 654.600 9.600 ;
        RECT 659.550 15.600 660.750 25.950 ;
        RECT 689.100 25.050 690.900 26.850 ;
        RECT 673.950 22.950 676.050 25.050 ;
        RECT 686.100 22.800 687.900 23.400 ;
        RECT 661.950 17.400 663.750 19.200 ;
        RECT 662.850 16.200 667.050 17.400 ;
        RECT 673.050 16.200 673.950 21.900 ;
        RECT 679.950 19.950 682.050 22.050 ;
        RECT 683.100 21.600 687.900 22.800 ;
        RECT 681.750 17.700 683.550 18.000 ;
        RECT 691.950 17.700 692.850 32.400 ;
        RECT 701.400 30.300 702.600 32.400 ;
        RECT 703.800 33.300 705.600 38.400 ;
        RECT 709.800 33.300 711.600 38.400 ;
        RECT 724.800 35.400 726.600 38.400 ;
        RECT 703.800 31.950 711.600 33.300 ;
        RECT 725.400 32.100 726.600 35.400 ;
        RECT 718.950 30.450 723.000 31.050 ;
        RECT 724.950 30.450 727.050 31.050 ;
        RECT 701.400 29.250 705.150 30.300 ;
        RECT 703.950 29.100 705.150 29.250 ;
        RECT 718.950 29.550 727.050 30.450 ;
        RECT 740.100 30.000 741.900 38.400 ;
        RECT 718.950 28.950 723.000 29.550 ;
        RECT 724.950 28.950 727.050 29.550 ;
        RECT 737.700 28.350 741.900 30.000 ;
        RECT 749.550 32.400 751.350 38.400 ;
        RECT 757.650 35.400 759.450 38.400 ;
        RECT 765.450 35.400 767.250 38.400 ;
        RECT 773.250 36.300 775.050 38.400 ;
        RECT 773.250 35.400 777.000 36.300 ;
        RECT 757.650 34.500 758.700 35.400 ;
        RECT 754.950 33.300 758.700 34.500 ;
        RECT 766.200 33.600 767.250 35.400 ;
        RECT 775.950 34.500 777.000 35.400 ;
        RECT 754.950 32.400 757.050 33.300 ;
        RECT 766.200 32.550 771.150 33.600 ;
        RECT 694.950 27.450 697.050 28.050 ;
        RECT 703.950 27.450 706.050 28.050 ;
        RECT 694.950 26.550 706.050 27.450 ;
        RECT 694.950 25.950 697.050 26.550 ;
        RECT 703.950 25.950 706.050 26.550 ;
        RECT 709.950 25.950 712.050 28.050 ;
        RECT 724.950 26.100 726.300 27.900 ;
        RECT 701.100 23.100 702.900 23.850 ;
        RECT 704.850 23.100 706.050 24.900 ;
        RECT 710.100 24.150 711.900 24.900 ;
        RECT 707.100 23.100 708.900 23.850 ;
        RECT 700.950 19.950 703.050 22.050 ;
        RECT 681.750 17.100 692.850 17.700 ;
        RECT 659.550 3.600 661.350 15.600 ;
        RECT 664.950 15.300 667.050 16.200 ;
        RECT 667.950 15.300 673.950 16.200 ;
        RECT 675.150 16.500 692.850 17.100 ;
        RECT 675.150 16.200 683.550 16.500 ;
        RECT 667.950 14.400 668.850 15.300 ;
        RECT 666.150 12.600 668.850 14.400 ;
        RECT 669.750 14.100 671.550 14.400 ;
        RECT 675.150 14.100 676.050 16.200 ;
        RECT 691.950 15.600 692.850 16.500 ;
        RECT 704.850 18.900 705.900 23.100 ;
        RECT 721.950 22.950 724.050 25.050 ;
        RECT 706.950 19.950 709.050 22.050 ;
        RECT 725.100 21.900 726.300 26.100 ;
        RECT 722.100 21.150 723.900 21.900 ;
        RECT 704.850 15.600 706.050 18.900 ;
        RECT 724.950 16.650 726.300 21.900 ;
        RECT 727.950 19.950 733.050 22.050 ;
        RECT 737.700 20.100 738.600 28.350 ;
        RECT 749.550 28.050 750.750 32.400 ;
        RECT 769.350 31.800 771.150 32.550 ;
        RECT 772.650 31.800 774.450 33.600 ;
        RECT 775.950 32.400 778.050 34.500 ;
        RECT 781.050 32.400 782.850 38.400 ;
        RECT 788.400 35.400 790.200 38.400 ;
        RECT 773.100 28.800 774.150 31.800 ;
        RECT 740.100 26.100 741.900 26.850 ;
        RECT 749.550 25.950 750.900 28.050 ;
        RECT 751.950 25.950 754.050 28.050 ;
        RECT 755.100 26.250 755.850 28.050 ;
        RECT 762.150 27.600 780.000 28.800 ;
        RECT 762.150 27.000 763.950 27.600 ;
        RECT 773.100 27.000 774.900 27.600 ;
        RECT 763.050 26.100 763.950 27.000 ;
        RECT 779.100 26.850 780.000 27.600 ;
        RECT 739.950 22.950 742.050 25.050 ;
        RECT 742.950 19.950 748.050 22.050 ;
        RECT 728.100 18.150 729.900 18.900 ;
        RECT 736.950 16.950 739.050 19.050 ;
        RECT 743.100 18.150 744.900 18.900 ;
        RECT 746.100 17.100 747.900 17.850 ;
        RECT 723.600 15.600 726.300 16.650 ;
        RECT 669.750 13.200 676.050 14.100 ;
        RECT 676.950 14.700 678.750 15.300 ;
        RECT 676.950 13.500 684.450 14.700 ;
        RECT 669.750 12.600 671.550 13.200 ;
        RECT 683.250 12.600 684.450 13.500 ;
        RECT 664.950 9.600 668.850 11.700 ;
        RECT 673.950 11.550 675.750 12.300 ;
        RECT 678.750 11.550 680.550 12.300 ;
        RECT 673.950 10.500 680.550 11.550 ;
        RECT 683.250 10.500 688.050 12.600 ;
        RECT 667.050 3.600 668.850 9.600 ;
        RECT 674.850 3.600 676.650 10.500 ;
        RECT 683.250 9.600 684.450 10.500 ;
        RECT 682.650 3.600 684.450 9.600 ;
        RECT 691.050 3.600 692.850 15.600 ;
        RECT 704.700 3.600 706.500 15.600 ;
        RECT 723.600 3.600 725.400 15.600 ;
        RECT 737.700 10.800 738.600 15.900 ;
        RECT 745.950 13.950 748.050 16.050 ;
        RECT 749.550 15.600 750.750 25.950 ;
        RECT 779.100 25.050 780.900 26.850 ;
        RECT 763.950 22.950 766.050 25.050 ;
        RECT 751.950 17.400 753.750 19.200 ;
        RECT 752.850 16.200 757.050 17.400 ;
        RECT 763.050 16.200 763.950 21.900 ;
        RECT 769.950 19.950 772.050 25.050 ;
        RECT 776.100 22.800 777.900 23.400 ;
        RECT 773.100 21.600 777.900 22.800 ;
        RECT 771.750 17.700 773.550 18.000 ;
        RECT 781.950 17.700 782.850 32.400 ;
        RECT 789.000 31.500 790.200 35.400 ;
        RECT 794.700 32.400 796.500 38.400 ;
        RECT 789.000 30.600 794.100 31.500 ;
        RECT 792.150 29.700 794.100 30.600 ;
        RECT 792.150 29.100 793.050 29.700 ;
        RECT 795.000 29.100 796.200 32.400 ;
        RECT 811.200 31.200 813.000 38.400 ;
        RECT 809.400 30.300 813.000 31.200 ;
        RECT 787.950 22.950 790.050 28.050 ;
        RECT 792.150 24.900 792.900 29.100 ;
        RECT 809.400 26.100 810.600 30.300 ;
        RECT 788.100 21.150 789.900 21.900 ;
        RECT 771.750 17.100 782.850 17.700 ;
        RECT 792.150 18.300 793.050 24.900 ;
        RECT 792.150 17.400 794.100 18.300 ;
        RECT 737.700 9.900 744.300 10.800 ;
        RECT 737.700 9.600 738.600 9.900 ;
        RECT 736.800 3.600 738.600 9.600 ;
        RECT 742.800 9.600 744.300 9.900 ;
        RECT 742.800 3.600 744.600 9.600 ;
        RECT 749.550 3.600 751.350 15.600 ;
        RECT 754.950 15.300 757.050 16.200 ;
        RECT 757.950 15.300 763.950 16.200 ;
        RECT 765.150 16.500 782.850 17.100 ;
        RECT 765.150 16.200 773.550 16.500 ;
        RECT 757.950 14.400 758.850 15.300 ;
        RECT 756.150 12.600 758.850 14.400 ;
        RECT 759.750 14.100 761.550 14.400 ;
        RECT 765.150 14.100 766.050 16.200 ;
        RECT 781.950 15.600 782.850 16.500 ;
        RECT 759.750 13.200 766.050 14.100 ;
        RECT 766.950 14.700 768.750 15.300 ;
        RECT 766.950 13.500 774.450 14.700 ;
        RECT 759.750 12.600 761.550 13.200 ;
        RECT 773.250 12.600 774.450 13.500 ;
        RECT 754.950 9.600 758.850 11.700 ;
        RECT 763.950 11.550 765.750 12.300 ;
        RECT 768.750 11.550 770.550 12.300 ;
        RECT 763.950 10.500 770.550 11.550 ;
        RECT 773.250 10.500 778.050 12.600 ;
        RECT 757.050 3.600 758.850 9.600 ;
        RECT 764.850 3.600 766.650 10.500 ;
        RECT 773.250 9.600 774.450 10.500 ;
        RECT 772.650 3.600 774.450 9.600 ;
        RECT 781.050 3.600 782.850 15.600 ;
        RECT 788.400 16.500 794.100 17.400 ;
        RECT 788.400 9.600 789.600 16.500 ;
        RECT 795.000 15.600 796.200 24.900 ;
        RECT 808.950 24.450 811.050 25.050 ;
        RECT 826.950 24.450 829.050 25.050 ;
        RECT 808.950 23.550 829.050 24.450 ;
        RECT 808.950 22.950 811.050 23.550 ;
        RECT 826.950 22.950 829.050 23.550 ;
        RECT 806.100 20.100 807.900 20.850 ;
        RECT 805.950 16.950 808.050 19.050 ;
        RECT 788.400 3.600 790.200 9.600 ;
        RECT 794.700 3.600 796.500 15.600 ;
        RECT 809.400 9.600 810.600 21.900 ;
        RECT 812.100 20.100 813.900 20.850 ;
        RECT 811.950 16.950 814.050 19.050 ;
        RECT 809.400 3.600 811.200 9.600 ;
      LAYER metal2 ;
        RECT 331.950 817.950 334.050 820.050 ;
        RECT 382.950 819.450 385.050 820.050 ;
        RECT 388.950 819.450 391.050 820.050 ;
        RECT 382.950 818.400 391.050 819.450 ;
        RECT 382.950 817.950 385.050 818.400 ;
        RECT 388.950 817.950 391.050 818.400 ;
        RECT 433.950 817.950 436.050 820.050 ;
        RECT 472.950 817.950 475.050 820.050 ;
        RECT 514.950 819.450 517.050 820.050 ;
        RECT 520.950 819.450 523.050 820.050 ;
        RECT 514.950 818.400 523.050 819.450 ;
        RECT 514.950 817.950 517.050 818.400 ;
        RECT 520.950 817.950 523.050 818.400 ;
        RECT 58.950 814.950 61.050 817.050 ;
        RECT 160.950 814.950 163.050 817.050 ;
        RECT 13.950 811.950 16.050 814.050 ;
        RECT 37.950 811.950 40.050 814.050 ;
        RECT 14.400 808.050 15.450 811.950 ;
        RECT 4.950 805.950 7.050 808.050 ;
        RECT 13.950 805.950 16.050 808.050 ;
        RECT 16.950 805.950 19.050 808.050 ;
        RECT 5.400 772.050 6.450 805.950 ;
        RECT 17.400 802.050 18.450 805.950 ;
        RECT 28.950 802.950 31.050 808.050 ;
        RECT 10.950 799.950 16.050 802.050 ;
        RECT 16.950 799.950 19.050 802.050 ;
        RECT 31.950 799.950 37.050 802.050 ;
        RECT 25.950 796.950 28.050 799.050 ;
        RECT 26.400 793.050 27.450 796.950 ;
        RECT 38.400 796.050 39.450 811.950 ;
        RECT 59.400 808.050 60.450 814.950 ;
        RECT 94.950 808.950 97.050 811.050 ;
        RECT 49.950 805.950 52.050 808.050 ;
        RECT 58.950 805.950 61.050 808.050 ;
        RECT 76.950 805.950 79.050 808.050 ;
        RECT 43.950 799.950 49.050 802.050 ;
        RECT 34.950 793.950 40.050 796.050 ;
        RECT 25.950 790.950 28.050 793.050 ;
        RECT 50.400 784.050 51.450 805.950 ;
        RECT 52.950 799.950 58.050 802.050 ;
        RECT 59.400 796.050 60.450 805.950 ;
        RECT 70.950 802.950 73.050 805.050 ;
        RECT 61.950 796.950 64.050 802.050 ;
        RECT 58.950 793.950 61.050 796.050 ;
        RECT 49.950 781.950 52.050 784.050 ;
        RECT 61.950 781.950 64.050 784.050 ;
        RECT 43.950 772.950 46.050 775.050 ;
        RECT 4.950 769.950 7.050 772.050 ;
        RECT 13.950 769.950 16.050 772.050 ;
        RECT 7.950 760.950 10.050 766.050 ;
        RECT 14.400 763.050 15.450 769.950 ;
        RECT 44.400 763.050 45.450 772.950 ;
        RECT 58.950 769.950 61.050 772.050 ;
        RECT 49.950 763.950 52.050 766.050 ;
        RECT 13.950 760.950 16.050 763.050 ;
        RECT 28.950 760.950 31.050 763.050 ;
        RECT 34.950 760.950 40.050 763.050 ;
        RECT 43.950 760.950 46.050 763.050 ;
        RECT 10.950 754.950 13.050 757.050 ;
        RECT 16.950 754.950 19.050 760.050 ;
        RECT 11.400 729.450 12.450 754.950 ;
        RECT 22.950 751.950 25.050 754.050 ;
        RECT 16.950 730.050 19.050 730.200 ;
        RECT 19.950 730.050 22.050 730.200 ;
        RECT 13.950 729.450 16.050 730.050 ;
        RECT 11.400 728.400 16.050 729.450 ;
        RECT 13.950 724.950 16.050 728.400 ;
        RECT 16.950 728.100 22.050 730.050 ;
        RECT 18.000 727.950 21.000 728.100 ;
        RECT 16.950 721.950 19.050 726.900 ;
        RECT 10.950 718.950 13.050 721.050 ;
        RECT 11.400 688.050 12.450 718.950 ;
        RECT 23.400 718.050 24.450 751.950 ;
        RECT 29.400 730.050 30.450 760.950 ;
        RECT 31.950 754.950 37.050 757.050 ;
        RECT 43.800 754.950 45.900 757.050 ;
        RECT 28.950 727.950 31.050 730.050 ;
        RECT 34.950 727.950 37.050 730.050 ;
        RECT 25.950 721.950 28.050 727.050 ;
        RECT 35.400 724.050 36.450 727.950 ;
        RECT 44.400 727.050 45.450 754.950 ;
        RECT 46.950 751.950 49.050 757.050 ;
        RECT 50.400 739.050 51.450 763.950 ;
        RECT 59.400 757.050 60.450 769.950 ;
        RECT 62.400 763.050 63.450 781.950 ;
        RECT 71.400 772.050 72.450 802.950 ;
        RECT 77.400 802.050 78.450 805.950 ;
        RECT 88.950 802.950 91.050 805.050 ;
        RECT 76.950 799.950 79.050 802.050 ;
        RECT 89.400 799.050 90.450 802.950 ;
        RECT 95.400 799.050 96.450 808.950 ;
        RECT 112.950 805.050 115.050 808.050 ;
        RECT 130.950 805.950 133.050 808.050 ;
        RECT 136.950 805.950 139.050 808.050 ;
        RECT 112.950 802.950 118.050 805.050 ;
        RECT 100.950 799.950 103.050 802.050 ;
        RECT 103.950 799.950 106.050 802.050 ;
        RECT 121.950 799.950 124.050 805.050 ;
        RECT 79.950 796.950 82.050 799.050 ;
        RECT 85.950 797.400 90.450 799.050 ;
        RECT 85.950 796.950 90.000 797.400 ;
        RECT 94.950 796.950 97.050 799.050 ;
        RECT 80.400 790.050 81.450 796.950 ;
        RECT 97.950 790.950 100.050 793.050 ;
        RECT 79.950 787.950 82.050 790.050 ;
        RECT 73.950 781.950 76.050 784.050 ;
        RECT 70.950 769.950 73.050 772.050 ;
        RECT 74.400 769.050 75.450 781.950 ;
        RECT 91.950 772.950 94.050 775.050 ;
        RECT 92.400 769.050 93.450 772.950 ;
        RECT 73.950 766.950 76.050 769.050 ;
        RECT 92.400 766.950 97.050 769.050 ;
        RECT 82.950 765.450 87.000 766.050 ;
        RECT 82.950 763.950 87.450 765.450 ;
        RECT 61.950 760.950 64.050 763.050 ;
        RECT 67.950 760.950 70.050 763.050 ;
        RECT 73.950 760.950 79.050 763.050 ;
        RECT 58.950 754.950 61.050 757.050 ;
        RECT 61.950 754.950 67.050 757.050 ;
        RECT 68.400 751.050 69.450 760.950 ;
        RECT 86.400 760.050 87.450 763.950 ;
        RECT 79.950 754.950 82.050 760.050 ;
        RECT 85.950 757.950 88.050 760.050 ;
        RECT 67.950 748.950 70.050 751.050 ;
        RECT 49.950 736.950 52.050 739.050 ;
        RECT 76.950 736.950 79.050 739.050 ;
        RECT 46.950 727.950 49.050 730.050 ;
        RECT 43.950 724.950 46.050 727.050 ;
        RECT 34.950 721.950 37.050 724.050 ;
        RECT 19.950 715.950 25.050 718.050 ;
        RECT 26.400 703.050 27.450 721.950 ;
        RECT 47.400 712.050 48.450 727.950 ;
        RECT 77.400 727.050 78.450 736.950 ;
        RECT 82.950 727.950 85.050 730.050 ;
        RECT 52.950 724.950 58.050 727.050 ;
        RECT 76.950 724.950 79.050 727.050 ;
        RECT 58.950 721.950 64.050 724.050 ;
        RECT 52.950 718.950 55.050 721.050 ;
        RECT 67.950 718.950 70.050 724.050 ;
        RECT 77.400 720.450 78.450 724.950 ;
        RECT 83.400 724.050 84.450 727.950 ;
        RECT 86.400 724.050 87.450 757.950 ;
        RECT 92.400 741.450 93.450 766.950 ;
        RECT 98.400 763.200 99.450 790.950 ;
        RECT 101.400 778.050 102.450 799.950 ;
        RECT 100.950 775.950 103.050 778.050 ;
        RECT 104.400 771.450 105.450 799.950 ;
        RECT 109.950 796.950 112.050 799.050 ;
        RECT 115.950 796.950 118.050 799.050 ;
        RECT 110.400 790.050 111.450 796.950 ;
        RECT 109.950 787.950 112.050 790.050 ;
        RECT 110.400 772.050 111.450 787.950 ;
        RECT 116.400 780.450 117.450 796.950 ;
        RECT 131.400 787.050 132.450 805.950 ;
        RECT 133.950 799.950 136.050 805.050 ;
        RECT 130.950 784.950 133.050 787.050 ;
        RECT 137.400 784.050 138.450 805.950 ;
        RECT 139.950 799.950 142.050 802.050 ;
        RECT 151.950 799.950 154.050 805.050 ;
        RECT 136.950 781.950 139.050 784.050 ;
        RECT 118.950 780.450 121.050 781.050 ;
        RECT 116.400 779.400 121.050 780.450 ;
        RECT 118.950 778.950 121.050 779.400 ;
        RECT 104.400 771.000 108.450 771.450 ;
        RECT 104.400 770.400 109.050 771.000 ;
        RECT 106.950 766.950 109.050 770.400 ;
        RECT 109.950 769.950 112.050 772.050 ;
        RECT 119.400 766.050 120.450 778.950 ;
        RECT 124.950 769.950 127.050 772.050 ;
        RECT 103.950 763.950 106.050 766.050 ;
        RECT 112.950 763.950 118.050 766.050 ;
        RECT 118.950 763.950 121.050 766.050 ;
        RECT 97.950 763.050 100.050 763.200 ;
        RECT 96.000 762.600 100.050 763.050 ;
        RECT 89.400 740.400 93.450 741.450 ;
        RECT 95.400 761.100 100.050 762.600 ;
        RECT 95.400 760.950 99.000 761.100 ;
        RECT 89.400 727.050 90.450 740.400 ;
        RECT 95.400 733.050 96.450 760.950 ;
        RECT 100.950 760.050 103.050 760.200 ;
        RECT 99.000 759.900 103.050 760.050 ;
        RECT 97.950 758.100 103.050 759.900 ;
        RECT 97.950 757.950 102.000 758.100 ;
        RECT 97.950 757.800 100.050 757.950 ;
        RECT 100.950 754.800 103.050 756.900 ;
        RECT 101.400 735.450 102.450 754.800 ;
        RECT 104.400 754.050 105.450 763.950 ;
        RECT 106.950 757.950 109.050 760.050 ;
        RECT 103.950 751.950 106.050 754.050 ;
        RECT 107.400 751.050 108.450 757.950 ;
        RECT 112.950 751.950 115.050 754.050 ;
        RECT 125.400 753.450 126.450 769.950 ;
        RECT 137.400 769.050 138.450 781.950 ;
        RECT 130.950 766.950 133.050 769.050 ;
        RECT 136.950 766.950 139.050 769.050 ;
        RECT 127.950 763.950 130.050 766.050 ;
        RECT 128.400 757.050 129.450 763.950 ;
        RECT 131.400 760.050 132.450 766.950 ;
        RECT 130.950 757.950 133.050 760.050 ;
        RECT 127.950 754.950 130.050 757.050 ;
        RECT 125.400 752.400 129.450 753.450 ;
        RECT 106.950 748.950 109.050 751.050 ;
        RECT 101.400 734.400 105.450 735.450 ;
        RECT 94.950 730.950 97.050 733.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 79.950 722.400 84.450 724.050 ;
        RECT 79.950 721.950 84.000 722.400 ;
        RECT 85.950 721.950 88.050 724.050 ;
        RECT 97.950 721.950 100.050 727.050 ;
        RECT 77.400 719.400 81.450 720.450 ;
        RECT 46.950 709.950 49.050 712.050 ;
        RECT 25.950 700.950 28.050 703.050 ;
        RECT 31.950 691.950 34.050 694.050 ;
        RECT 10.950 685.950 13.050 688.050 ;
        RECT 16.950 687.450 21.000 688.050 ;
        RECT 22.950 687.450 25.050 691.050 ;
        RECT 32.400 688.050 33.450 691.950 ;
        RECT 53.400 688.050 54.450 718.950 ;
        RECT 61.950 715.950 64.050 718.050 ;
        RECT 62.400 709.050 63.450 715.950 ;
        RECT 61.950 706.950 64.050 709.050 ;
        RECT 76.950 697.950 79.050 700.050 ;
        RECT 70.950 691.950 73.050 694.050 ;
        RECT 16.950 686.400 25.050 687.450 ;
        RECT 16.950 685.950 21.000 686.400 ;
        RECT 22.950 685.950 25.050 686.400 ;
        RECT 31.950 685.950 34.050 688.050 ;
        RECT 11.400 682.050 12.450 685.950 ;
        RECT 28.950 685.050 31.050 685.200 ;
        RECT 25.950 683.100 31.050 685.050 ;
        RECT 25.950 682.950 30.000 683.100 ;
        RECT 34.950 682.950 37.050 685.050 ;
        RECT 37.950 682.950 40.050 688.050 ;
        RECT 52.950 685.950 55.050 688.050 ;
        RECT 71.400 685.050 72.450 691.950 ;
        RECT 46.950 682.950 49.050 685.050 ;
        RECT 64.950 682.950 67.050 685.050 ;
        RECT 70.950 682.950 73.050 685.050 ;
        RECT 10.950 679.950 13.050 682.050 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 25.950 679.950 28.050 682.950 ;
        RECT 14.400 657.450 15.450 679.950 ;
        RECT 28.950 679.800 31.050 681.900 ;
        RECT 29.400 676.050 30.450 679.800 ;
        RECT 35.400 679.050 36.450 682.950 ;
        RECT 34.950 676.950 37.050 679.050 ;
        RECT 28.950 673.950 31.050 676.050 ;
        RECT 11.400 656.400 15.450 657.450 ;
        RECT 11.400 643.050 12.450 656.400 ;
        RECT 13.950 652.950 16.050 655.050 ;
        RECT 14.400 649.050 15.450 652.950 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 19.950 646.950 22.050 649.050 ;
        RECT 20.400 643.050 21.450 646.950 ;
        RECT 7.950 640.950 10.050 643.050 ;
        RECT 10.950 640.950 13.050 643.050 ;
        RECT 16.950 640.950 21.450 643.050 ;
        RECT 22.950 640.950 25.050 643.050 ;
        RECT 8.400 610.050 9.450 640.950 ;
        RECT 7.950 607.950 10.050 610.050 ;
        RECT 13.950 607.950 19.050 610.050 ;
        RECT 16.950 601.950 19.050 604.050 ;
        RECT 7.950 598.950 10.050 601.050 ;
        RECT 8.400 574.050 9.450 598.950 ;
        RECT 17.400 595.050 18.450 601.950 ;
        RECT 20.400 601.050 21.450 640.950 ;
        RECT 19.950 598.950 22.050 601.050 ;
        RECT 23.400 598.050 24.450 640.950 ;
        RECT 29.400 613.050 30.450 673.950 ;
        RECT 31.950 643.950 34.050 649.050 ;
        RECT 35.400 646.050 36.450 676.950 ;
        RECT 34.950 643.950 37.050 646.050 ;
        RECT 38.400 640.050 39.450 682.950 ;
        RECT 47.400 676.050 48.450 682.950 ;
        RECT 65.400 679.050 66.450 682.950 ;
        RECT 49.950 676.950 54.900 679.050 ;
        RECT 55.950 676.950 58.050 679.050 ;
        RECT 64.950 676.950 67.050 679.050 ;
        RECT 46.950 673.950 49.050 676.050 ;
        RECT 56.400 658.050 57.450 676.950 ;
        RECT 71.400 658.200 72.450 682.950 ;
        RECT 77.400 679.050 78.450 697.950 ;
        RECT 80.400 679.050 81.450 719.400 ;
        RECT 86.400 718.050 87.450 721.950 ;
        RECT 82.950 716.400 87.450 718.050 ;
        RECT 82.950 715.950 87.000 716.400 ;
        RECT 104.400 697.050 105.450 734.400 ;
        RECT 109.950 727.950 112.050 730.050 ;
        RECT 110.400 724.050 111.450 727.950 ;
        RECT 113.400 724.050 114.450 751.950 ;
        RECT 115.950 739.950 118.050 742.050 ;
        RECT 116.400 730.050 117.450 739.950 ;
        RECT 121.950 736.950 124.050 739.050 ;
        RECT 122.400 730.050 123.450 736.950 ;
        RECT 128.400 730.050 129.450 752.400 ;
        RECT 140.400 748.050 141.450 799.950 ;
        RECT 148.950 793.950 151.050 799.050 ;
        RECT 154.950 796.950 160.050 799.050 ;
        RECT 149.400 766.200 150.450 793.950 ;
        RECT 161.400 772.050 162.450 814.950 ;
        RECT 166.950 802.950 169.050 808.050 ;
        RECT 184.950 805.950 187.050 808.050 ;
        RECT 226.950 805.950 229.050 808.050 ;
        RECT 241.950 805.950 247.050 808.050 ;
        RECT 259.950 805.950 262.050 808.050 ;
        RECT 265.950 807.450 270.000 808.050 ;
        RECT 265.950 805.950 270.450 807.450 ;
        RECT 280.950 805.950 283.050 808.050 ;
        RECT 286.950 805.950 289.050 808.050 ;
        RECT 307.950 805.950 310.050 811.050 ;
        RECT 319.950 808.950 322.050 811.050 ;
        RECT 316.950 808.050 319.050 808.200 ;
        RECT 313.950 806.100 319.050 808.050 ;
        RECT 313.950 805.950 318.000 806.100 ;
        RECT 163.950 796.950 166.050 799.050 ;
        RECT 160.950 769.950 163.050 772.050 ;
        RECT 142.950 763.950 145.050 766.050 ;
        RECT 148.950 764.100 151.050 766.200 ;
        RECT 139.950 745.950 142.050 748.050 ;
        RECT 136.950 736.950 139.050 739.050 ;
        RECT 133.950 730.950 136.050 733.050 ;
        RECT 115.950 727.950 118.050 730.050 ;
        RECT 121.950 727.950 124.050 730.050 ;
        RECT 127.950 727.950 130.050 730.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 109.950 721.950 112.050 724.050 ;
        RECT 112.950 721.950 115.050 724.050 ;
        RECT 118.950 721.950 124.050 724.050 ;
        RECT 113.400 718.050 114.450 721.950 ;
        RECT 112.950 715.950 115.050 718.050 ;
        RECT 115.950 712.950 118.050 715.050 ;
        RECT 103.950 694.950 106.050 697.050 ;
        RECT 88.950 688.950 91.050 691.050 ;
        RECT 106.950 688.950 109.050 691.050 ;
        RECT 89.400 685.050 90.450 688.950 ;
        RECT 88.950 682.950 91.050 685.050 ;
        RECT 94.950 682.950 100.050 685.050 ;
        RECT 100.950 682.950 103.050 688.050 ;
        RECT 76.800 676.950 78.900 679.050 ;
        RECT 79.950 676.950 82.050 679.050 ;
        RECT 91.950 676.950 97.050 679.050 ;
        RECT 46.950 655.950 49.050 658.050 ;
        RECT 55.950 655.950 58.050 658.050 ;
        RECT 64.950 655.950 67.050 658.050 ;
        RECT 70.950 656.100 73.050 658.200 ;
        RECT 47.400 640.050 48.450 655.950 ;
        RECT 52.950 652.950 55.050 655.050 ;
        RECT 53.400 649.200 54.450 652.950 ;
        RECT 65.400 652.050 66.450 655.950 ;
        RECT 64.950 649.950 67.050 652.050 ;
        RECT 70.950 649.950 73.050 654.900 ;
        RECT 94.950 649.950 97.050 652.050 ;
        RECT 52.950 647.100 55.050 649.200 ;
        RECT 65.400 646.050 66.450 649.950 ;
        RECT 49.950 645.900 54.000 646.050 ;
        RECT 49.950 643.950 55.050 645.900 ;
        RECT 64.800 643.950 66.900 646.050 ;
        RECT 68.100 643.950 73.050 646.050 ;
        RECT 76.950 643.950 79.050 646.050 ;
        RECT 82.950 643.950 88.050 646.050 ;
        RECT 52.950 643.800 55.050 643.950 ;
        RECT 55.950 640.950 58.050 643.050 ;
        RECT 37.950 637.950 40.050 640.050 ;
        RECT 46.950 637.950 49.050 640.050 ;
        RECT 49.950 637.950 52.050 640.050 ;
        RECT 28.950 610.950 31.050 613.050 ;
        RECT 25.950 604.950 28.050 610.050 ;
        RECT 34.950 607.950 37.050 613.050 ;
        RECT 40.950 610.950 43.050 613.050 ;
        RECT 46.950 610.950 49.050 613.050 ;
        RECT 31.950 604.950 34.050 607.050 ;
        RECT 27.000 603.450 31.050 604.050 ;
        RECT 26.400 601.950 31.050 603.450 ;
        RECT 22.950 595.950 25.050 598.050 ;
        RECT 26.400 595.050 27.450 601.950 ;
        RECT 32.400 598.050 33.450 604.950 ;
        RECT 31.950 595.950 34.050 598.050 ;
        RECT 16.950 592.950 19.050 595.050 ;
        RECT 25.950 592.950 28.050 595.050 ;
        RECT 10.950 574.950 13.050 577.050 ;
        RECT 7.950 571.950 10.050 574.050 ;
        RECT 11.400 568.050 12.450 574.950 ;
        RECT 13.950 571.950 19.050 574.050 ;
        RECT 25.950 571.950 28.050 574.050 ;
        RECT 34.950 572.100 37.050 577.050 ;
        RECT 10.950 565.950 13.050 568.050 ;
        RECT 16.950 565.950 22.050 568.050 ;
        RECT 11.400 550.050 12.450 565.950 ;
        RECT 10.950 547.950 13.050 550.050 ;
        RECT 13.950 532.950 16.050 535.050 ;
        RECT 14.400 529.050 15.450 532.950 ;
        RECT 20.400 529.050 21.450 565.950 ;
        RECT 22.950 562.950 25.050 568.050 ;
        RECT 26.400 535.050 27.450 571.950 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 29.400 559.050 30.450 568.950 ;
        RECT 34.950 568.800 37.050 570.900 ;
        RECT 31.950 562.950 34.050 568.050 ;
        RECT 35.400 562.050 36.450 568.800 ;
        RECT 34.950 559.950 37.050 562.050 ;
        RECT 28.950 556.950 31.050 559.050 ;
        RECT 41.400 555.450 42.450 610.950 ;
        RECT 47.400 607.050 48.450 610.950 ;
        RECT 46.950 604.950 49.050 607.050 ;
        RECT 50.400 601.050 51.450 637.950 ;
        RECT 52.950 607.950 55.050 610.050 ;
        RECT 49.950 598.950 52.050 601.050 ;
        RECT 50.400 580.050 51.450 598.950 ;
        RECT 49.950 577.950 52.050 580.050 ;
        RECT 53.400 574.050 54.450 607.950 ;
        RECT 49.950 572.400 54.450 574.050 ;
        RECT 49.950 571.950 54.000 572.400 ;
        RECT 49.950 568.950 52.050 571.950 ;
        RECT 46.950 565.950 49.050 568.050 ;
        RECT 47.400 559.050 48.450 565.950 ;
        RECT 52.950 562.950 55.050 568.050 ;
        RECT 46.950 556.950 49.050 559.050 ;
        RECT 41.400 554.400 45.450 555.450 ;
        RECT 31.950 535.050 34.050 535.200 ;
        RECT 25.950 532.950 28.050 535.050 ;
        RECT 28.950 533.100 34.050 535.050 ;
        RECT 28.950 532.950 33.000 533.100 ;
        RECT 13.950 526.950 16.050 529.050 ;
        RECT 19.950 526.050 22.050 529.050 ;
        RECT 31.950 527.100 34.050 531.900 ;
        RECT 37.950 529.950 40.050 532.050 ;
        RECT 16.800 525.000 18.900 526.050 ;
        RECT 19.950 525.000 22.200 526.050 ;
        RECT 33.000 525.900 37.050 526.050 ;
        RECT 16.800 523.950 19.050 525.000 ;
        RECT 20.100 523.950 22.200 525.000 ;
        RECT 31.950 523.950 37.050 525.900 ;
        RECT 4.950 520.950 7.050 523.050 ;
        RECT 16.950 520.950 19.050 523.950 ;
        RECT 31.950 523.800 34.050 523.950 ;
        RECT 5.400 496.050 6.450 520.950 ;
        RECT 4.950 493.950 7.050 496.050 ;
        RECT 22.950 493.950 25.050 496.050 ;
        RECT 31.950 493.950 34.050 496.050 ;
        RECT 7.950 490.050 10.050 490.200 ;
        RECT 10.950 490.050 13.050 490.200 ;
        RECT 7.950 488.100 13.050 490.050 ;
        RECT 9.000 487.950 12.000 488.100 ;
        RECT 7.950 484.800 10.050 486.900 ;
        RECT 13.950 484.950 16.050 490.050 ;
        RECT 19.950 487.950 22.050 493.050 ;
        RECT 1.950 466.950 4.050 469.050 ;
        RECT 2.400 454.200 3.450 466.950 ;
        RECT 1.950 452.100 4.050 454.200 ;
        RECT 4.950 451.950 7.050 454.050 ;
        RECT 1.950 448.800 4.050 450.900 ;
        RECT 2.400 436.050 3.450 448.800 ;
        RECT 1.950 433.950 4.050 436.050 ;
        RECT 5.400 418.050 6.450 451.950 ;
        RECT 8.400 451.200 9.450 484.800 ;
        RECT 23.400 469.050 24.450 493.950 ;
        RECT 32.400 484.050 33.450 493.950 ;
        RECT 38.400 484.050 39.450 529.950 ;
        RECT 44.400 523.050 45.450 554.400 ;
        RECT 47.400 541.050 48.450 556.950 ;
        RECT 56.400 547.050 57.450 640.950 ;
        RECT 70.950 625.950 73.050 628.050 ;
        RECT 64.950 616.950 67.050 619.050 ;
        RECT 58.950 604.950 61.050 607.050 ;
        RECT 55.950 544.950 58.050 547.050 ;
        RECT 46.950 538.950 49.050 541.050 ;
        RECT 55.950 538.950 58.050 541.050 ;
        RECT 46.950 532.950 49.050 535.050 ;
        RECT 47.400 529.050 48.450 532.950 ;
        RECT 46.950 526.950 49.050 529.050 ;
        RECT 49.800 523.950 51.900 526.050 ;
        RECT 53.100 525.000 55.200 526.050 ;
        RECT 52.950 523.950 55.200 525.000 ;
        RECT 43.950 520.950 46.050 523.050 ;
        RECT 50.400 516.450 51.450 523.950 ;
        RECT 52.950 520.950 55.050 523.950 ;
        RECT 56.400 520.050 57.450 538.950 ;
        RECT 55.950 517.950 58.050 520.050 ;
        RECT 50.400 515.400 54.450 516.450 ;
        RECT 43.950 499.950 46.050 502.050 ;
        RECT 44.400 493.050 45.450 499.950 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 53.400 490.050 54.450 515.400 ;
        RECT 59.400 510.450 60.450 604.950 ;
        RECT 65.400 604.050 66.450 616.950 ;
        RECT 71.400 613.050 72.450 625.950 ;
        RECT 77.400 613.050 78.450 643.950 ;
        RECT 95.400 640.050 96.450 649.950 ;
        RECT 94.950 637.950 97.050 640.050 ;
        RECT 91.950 631.950 94.050 634.050 ;
        RECT 79.950 613.950 82.050 616.050 ;
        RECT 70.950 610.950 73.050 613.050 ;
        RECT 76.950 610.950 79.050 613.050 ;
        RECT 67.950 604.950 73.050 607.050 ;
        RECT 64.950 601.950 67.050 604.050 ;
        RECT 70.950 598.950 73.050 601.050 ;
        RECT 61.950 577.950 64.050 580.050 ;
        RECT 62.400 571.050 63.450 577.950 ;
        RECT 62.400 569.400 67.050 571.050 ;
        RECT 63.000 568.950 67.050 569.400 ;
        RECT 71.400 565.050 72.450 598.950 ;
        RECT 80.400 577.200 81.450 613.950 ;
        RECT 82.950 610.950 85.050 613.050 ;
        RECT 83.400 607.050 84.450 610.950 ;
        RECT 82.950 604.950 85.050 607.050 ;
        RECT 88.950 604.950 91.050 607.050 ;
        RECT 89.400 601.050 90.450 604.950 ;
        RECT 92.400 601.050 93.450 631.950 ;
        RECT 98.400 607.050 99.450 682.950 ;
        RECT 100.950 676.950 103.050 679.050 ;
        RECT 103.950 676.950 106.050 679.050 ;
        RECT 101.400 646.050 102.450 676.950 ;
        RECT 104.400 664.050 105.450 676.950 ;
        RECT 107.400 673.050 108.450 688.950 ;
        RECT 106.950 670.950 109.050 673.050 ;
        RECT 103.950 661.950 106.050 664.050 ;
        RECT 100.950 643.950 103.050 646.050 ;
        RECT 101.400 613.050 102.450 643.950 ;
        RECT 104.400 634.050 105.450 661.950 ;
        RECT 106.950 649.950 109.050 652.050 ;
        RECT 107.400 646.050 108.450 649.950 ;
        RECT 106.950 643.950 109.050 646.050 ;
        RECT 103.950 631.950 106.050 634.050 ;
        RECT 107.400 628.050 108.450 643.950 ;
        RECT 112.950 640.950 115.050 643.050 ;
        RECT 106.950 625.950 109.050 628.050 ;
        RECT 113.400 619.050 114.450 640.950 ;
        RECT 112.950 616.950 115.050 619.050 ;
        RECT 109.950 613.950 112.050 616.050 ;
        RECT 100.950 610.950 103.050 613.050 ;
        RECT 110.400 610.050 111.450 613.950 ;
        RECT 109.950 607.950 112.050 610.050 ;
        RECT 97.950 604.950 100.050 607.050 ;
        RECT 100.950 604.950 106.050 607.050 ;
        RECT 113.400 604.050 114.450 616.950 ;
        RECT 116.400 610.050 117.450 712.950 ;
        RECT 118.950 700.950 121.050 703.050 ;
        RECT 119.400 679.050 120.450 700.950 ;
        RECT 121.950 682.950 124.050 688.050 ;
        RECT 118.950 676.950 121.050 679.050 ;
        RECT 125.400 652.050 126.450 724.950 ;
        RECT 128.400 715.050 129.450 727.950 ;
        RECT 134.400 724.050 135.450 730.950 ;
        RECT 133.950 721.950 136.050 724.050 ;
        RECT 133.950 715.950 136.050 718.050 ;
        RECT 127.950 712.950 130.050 715.050 ;
        RECT 134.400 712.050 135.450 715.950 ;
        RECT 133.950 709.950 136.050 712.050 ;
        RECT 137.400 709.050 138.450 736.950 ;
        RECT 143.400 733.050 144.450 763.950 ;
        RECT 148.950 757.950 151.050 762.900 ;
        RECT 154.950 760.950 157.050 766.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 145.950 754.950 148.050 757.050 ;
        RECT 151.950 754.950 154.050 757.050 ;
        RECT 157.950 754.950 160.050 757.050 ;
        RECT 142.950 730.950 145.050 733.050 ;
        RECT 146.400 727.200 147.450 754.950 ;
        RECT 152.400 748.050 153.450 754.950 ;
        RECT 158.400 748.050 159.450 754.950 ;
        RECT 151.950 745.950 154.050 748.050 ;
        RECT 157.950 745.950 160.050 748.050 ;
        RECT 161.400 733.050 162.450 757.950 ;
        RECT 164.400 757.050 165.450 796.950 ;
        RECT 167.400 796.050 168.450 802.950 ;
        RECT 166.950 793.950 169.050 796.050 ;
        RECT 185.400 781.050 186.450 805.950 ;
        RECT 187.950 799.950 190.050 805.050 ;
        RECT 193.950 800.100 196.050 805.050 ;
        RECT 208.950 802.950 211.050 805.050 ;
        RECT 193.950 796.800 196.050 798.900 ;
        RECT 184.950 778.950 187.050 781.050 ;
        RECT 175.950 766.950 178.050 769.050 ;
        RECT 187.950 766.950 190.050 769.050 ;
        RECT 176.400 763.050 177.450 766.950 ;
        RECT 166.950 760.950 169.050 763.050 ;
        RECT 175.950 760.950 178.050 763.050 ;
        RECT 181.950 760.950 187.050 763.050 ;
        RECT 163.950 754.950 166.050 757.050 ;
        RECT 167.400 739.050 168.450 760.950 ;
        RECT 172.950 754.950 175.050 757.050 ;
        RECT 178.950 754.950 184.050 757.050 ;
        RECT 166.950 736.950 169.050 739.050 ;
        RECT 151.950 727.950 154.050 733.050 ;
        RECT 160.950 730.950 163.050 733.050 ;
        RECT 163.950 727.950 166.050 730.050 ;
        RECT 139.950 724.950 142.050 727.050 ;
        RECT 145.950 725.100 148.050 727.200 ;
        RECT 136.950 706.950 139.050 709.050 ;
        RECT 127.950 685.950 130.050 688.050 ;
        RECT 128.400 682.050 129.450 685.950 ;
        RECT 133.950 682.950 136.050 688.050 ;
        RECT 137.400 682.050 138.450 706.950 ;
        RECT 140.400 703.050 141.450 724.950 ;
        RECT 145.950 721.800 148.050 723.900 ;
        RECT 139.950 700.950 142.050 703.050 ;
        RECT 142.950 694.950 145.050 697.050 ;
        RECT 139.950 685.950 142.050 691.050 ;
        RECT 127.950 679.950 130.050 682.050 ;
        RECT 136.950 679.950 139.050 682.050 ;
        RECT 128.400 655.200 129.450 679.950 ;
        RECT 136.950 670.950 139.050 673.050 ;
        RECT 130.950 661.950 133.050 664.050 ;
        RECT 127.950 653.100 130.050 655.200 ;
        RECT 131.400 652.050 132.450 661.950 ;
        RECT 137.400 655.050 138.450 670.950 ;
        RECT 143.400 670.050 144.450 694.950 ;
        RECT 142.950 667.950 145.050 670.050 ;
        RECT 146.400 658.050 147.450 721.800 ;
        RECT 152.400 690.450 153.450 727.950 ;
        RECT 164.400 709.050 165.450 727.950 ;
        RECT 173.400 724.050 174.450 754.950 ;
        RECT 188.400 751.050 189.450 766.950 ;
        RECT 194.400 763.050 195.450 796.800 ;
        RECT 209.400 778.050 210.450 802.950 ;
        RECT 227.400 802.050 228.450 805.950 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 211.950 799.950 217.050 802.050 ;
        RECT 223.950 799.950 226.050 802.050 ;
        RECT 226.950 799.950 229.050 802.050 ;
        RECT 224.400 796.050 225.450 799.950 ;
        RECT 229.950 796.950 232.050 802.050 ;
        RECT 247.950 799.950 250.050 802.050 ;
        RECT 214.950 793.950 220.050 796.050 ;
        RECT 223.950 793.950 226.050 796.050 ;
        RECT 230.400 787.050 231.450 796.950 ;
        RECT 244.950 793.950 247.050 799.050 ;
        RECT 248.400 787.050 249.450 799.950 ;
        RECT 251.400 796.050 252.450 802.950 ;
        RECT 260.400 802.050 261.450 805.950 ;
        RECT 259.950 799.950 262.050 802.050 ;
        RECT 262.950 796.950 265.050 802.050 ;
        RECT 250.950 793.950 253.050 796.050 ;
        RECT 211.950 784.950 214.050 787.050 ;
        RECT 229.950 784.950 232.050 787.050 ;
        RECT 247.950 784.950 250.050 787.050 ;
        RECT 208.950 775.950 211.050 778.050 ;
        RECT 205.950 763.950 208.050 766.050 ;
        RECT 190.950 761.400 195.450 763.050 ;
        RECT 190.950 760.950 195.000 761.400 ;
        RECT 191.400 757.050 192.450 760.950 ;
        RECT 193.950 757.950 199.050 760.050 ;
        RECT 190.950 754.950 193.050 757.050 ;
        RECT 199.950 754.950 202.050 760.050 ;
        RECT 187.950 748.950 190.050 751.050 ;
        RECT 178.950 745.950 181.050 748.050 ;
        RECT 169.950 721.950 172.050 724.050 ;
        RECT 173.400 722.400 178.050 724.050 ;
        RECT 174.000 721.950 178.050 722.400 ;
        RECT 170.400 718.050 171.450 721.950 ;
        RECT 169.950 715.950 172.050 718.050 ;
        RECT 163.950 706.950 166.050 709.050 ;
        RECT 179.400 706.050 180.450 745.950 ;
        RECT 193.950 739.950 196.050 742.050 ;
        RECT 184.950 733.950 187.050 736.050 ;
        RECT 185.400 730.050 186.450 733.950 ;
        RECT 184.950 727.950 187.050 730.050 ;
        RECT 181.950 724.950 184.050 727.050 ;
        RECT 190.950 724.950 193.050 730.050 ;
        RECT 178.950 703.950 181.050 706.050 ;
        RECT 175.950 700.950 178.050 703.050 ;
        RECT 160.950 697.950 163.050 700.050 ;
        RECT 149.400 689.400 153.450 690.450 ;
        RECT 149.400 664.050 150.450 689.400 ;
        RECT 151.950 685.950 154.050 688.050 ;
        RECT 152.400 676.050 153.450 685.950 ;
        RECT 161.400 685.200 162.450 697.950 ;
        RECT 163.950 688.950 166.050 691.050 ;
        RECT 160.950 683.100 163.050 685.200 ;
        RECT 157.950 681.900 162.000 682.050 ;
        RECT 157.950 679.950 163.050 681.900 ;
        RECT 160.950 679.800 163.050 679.950 ;
        RECT 151.950 673.950 154.050 676.050 ;
        RECT 151.950 667.950 154.050 670.050 ;
        RECT 148.950 661.950 151.050 664.050 ;
        RECT 152.400 661.050 153.450 667.950 ;
        RECT 164.400 667.050 165.450 688.950 ;
        RECT 169.950 685.950 172.050 688.050 ;
        RECT 170.400 682.050 171.450 685.950 ;
        RECT 169.950 679.950 172.050 682.050 ;
        RECT 163.950 664.950 166.050 667.050 ;
        RECT 169.950 661.950 172.050 664.050 ;
        RECT 151.950 658.950 154.050 661.050 ;
        RECT 163.950 658.950 166.050 661.050 ;
        RECT 145.950 655.950 148.050 658.050 ;
        RECT 136.950 652.950 139.050 655.050 ;
        RECT 121.950 650.400 126.450 652.050 ;
        RECT 129.000 651.900 132.450 652.050 ;
        RECT 121.950 649.950 126.000 650.400 ;
        RECT 127.950 650.250 132.450 651.900 ;
        RECT 127.950 649.950 132.000 650.250 ;
        RECT 133.950 649.950 136.050 652.050 ;
        RECT 127.950 649.800 130.050 649.950 ;
        RECT 118.950 640.950 121.050 646.050 ;
        RECT 124.950 643.950 130.050 646.050 ;
        RECT 134.400 625.050 135.450 649.950 ;
        RECT 133.950 622.950 136.050 625.050 ;
        RECT 115.950 607.950 118.050 610.050 ;
        RECT 121.950 607.950 124.050 610.050 ;
        RECT 127.950 607.950 130.050 613.050 ;
        RECT 106.950 601.950 112.050 604.050 ;
        RECT 112.950 601.950 118.050 604.050 ;
        RECT 88.950 598.950 91.050 601.050 ;
        RECT 91.950 598.950 94.050 601.050 ;
        RECT 92.400 592.050 93.450 598.950 ;
        RECT 91.950 589.950 94.050 592.050 ;
        RECT 88.950 580.950 91.050 583.050 ;
        RECT 103.950 580.950 106.050 583.050 ;
        RECT 79.950 575.100 82.050 577.200 ;
        RECT 79.950 571.800 82.050 573.900 ;
        RECT 85.950 571.950 88.050 577.050 ;
        RECT 61.950 562.950 64.050 565.050 ;
        RECT 67.950 562.950 70.050 565.050 ;
        RECT 70.950 562.950 73.050 565.050 ;
        RECT 62.400 529.050 63.450 562.950 ;
        RECT 64.950 553.950 67.050 556.050 ;
        RECT 65.400 529.050 66.450 553.950 ;
        RECT 68.400 553.050 69.450 562.950 ;
        RECT 67.950 550.950 70.050 553.050 ;
        RECT 70.950 547.950 73.050 550.050 ;
        RECT 67.950 544.950 70.050 547.050 ;
        RECT 61.950 526.950 64.050 529.050 ;
        RECT 64.950 524.100 67.050 529.050 ;
        RECT 64.950 520.800 67.050 522.900 ;
        RECT 59.400 509.400 63.450 510.450 ;
        RECT 40.950 489.450 45.000 490.050 ;
        RECT 40.950 487.950 45.450 489.450 ;
        RECT 52.950 487.950 55.050 490.050 ;
        RECT 31.950 481.950 34.050 484.050 ;
        RECT 37.950 481.950 40.050 484.050 ;
        RECT 22.950 466.950 25.050 469.050 ;
        RECT 40.950 463.950 43.050 466.050 ;
        RECT 10.950 460.950 13.050 463.050 ;
        RECT 22.950 460.950 25.050 463.050 ;
        RECT 7.950 449.100 10.050 451.200 ;
        RECT 11.400 448.050 12.450 460.950 ;
        RECT 16.950 454.950 19.050 457.050 ;
        RECT 13.950 448.950 16.050 454.050 ;
        RECT 7.950 445.800 10.050 447.900 ;
        RECT 10.950 445.950 13.050 448.050 ;
        RECT 4.950 415.950 7.050 418.050 ;
        RECT 1.950 364.950 4.050 367.050 ;
        RECT 2.400 217.050 3.450 364.950 ;
        RECT 8.400 343.050 9.450 445.800 ;
        RECT 17.400 442.050 18.450 454.950 ;
        RECT 23.400 451.050 24.450 460.950 ;
        RECT 37.950 454.950 40.050 457.050 ;
        RECT 22.950 448.950 25.050 451.050 ;
        RECT 28.950 450.450 33.000 451.050 ;
        RECT 28.950 448.950 33.450 450.450 ;
        RECT 25.950 442.950 28.050 448.050 ;
        RECT 32.400 442.050 33.450 448.950 ;
        RECT 34.950 442.950 37.050 448.050 ;
        RECT 16.950 439.950 19.050 442.050 ;
        RECT 31.950 439.950 34.050 442.050 ;
        RECT 19.950 433.950 22.050 436.050 ;
        RECT 20.400 418.050 21.450 433.950 ;
        RECT 28.950 427.950 31.050 430.050 ;
        RECT 29.400 418.050 30.450 427.950 ;
        RECT 10.950 415.950 16.050 418.050 ;
        RECT 19.950 415.950 22.050 418.050 ;
        RECT 28.950 415.950 31.050 418.050 ;
        RECT 38.400 415.050 39.450 454.950 ;
        RECT 16.950 409.950 22.050 412.050 ;
        RECT 22.950 409.950 28.050 412.050 ;
        RECT 31.950 409.950 34.050 415.050 ;
        RECT 37.950 412.950 40.050 415.050 ;
        RECT 41.400 411.450 42.450 463.950 ;
        RECT 44.400 445.050 45.450 487.950 ;
        RECT 46.950 484.950 49.050 487.050 ;
        RECT 47.400 481.050 48.450 484.950 ;
        RECT 46.950 478.950 49.050 481.050 ;
        RECT 53.400 457.050 54.450 487.950 ;
        RECT 58.950 478.950 61.050 481.050 ;
        RECT 55.950 469.950 58.050 472.050 ;
        RECT 52.950 454.950 55.050 457.050 ;
        RECT 46.950 448.950 49.050 451.050 ;
        RECT 43.950 442.950 46.050 445.050 ;
        RECT 43.950 427.950 46.050 430.050 ;
        RECT 44.400 415.050 45.450 427.950 ;
        RECT 47.400 418.050 48.450 448.950 ;
        RECT 52.950 445.950 55.050 451.050 ;
        RECT 56.400 445.050 57.450 469.950 ;
        RECT 55.950 442.950 58.050 445.050 ;
        RECT 59.400 418.050 60.450 478.950 ;
        RECT 62.400 421.200 63.450 509.400 ;
        RECT 65.400 502.050 66.450 520.800 ;
        RECT 64.950 499.950 67.050 502.050 ;
        RECT 64.950 493.950 67.050 496.050 ;
        RECT 65.400 472.050 66.450 493.950 ;
        RECT 64.950 469.950 67.050 472.050 ;
        RECT 68.400 466.050 69.450 544.950 ;
        RECT 71.400 529.050 72.450 547.950 ;
        RECT 80.400 529.050 81.450 571.800 ;
        RECT 89.400 568.050 90.450 580.950 ;
        RECT 97.950 571.950 100.050 574.050 ;
        RECT 98.400 568.200 99.450 571.950 ;
        RECT 104.400 571.050 105.450 580.950 ;
        RECT 122.400 574.050 123.450 607.950 ;
        RECT 137.400 607.050 138.450 652.950 ;
        RECT 146.400 649.200 147.450 655.950 ;
        RECT 139.950 646.950 145.050 649.050 ;
        RECT 145.950 647.100 148.050 649.200 ;
        RECT 151.950 646.200 154.050 649.050 ;
        RECT 147.000 645.900 150.000 646.050 ;
        RECT 145.950 645.300 150.000 645.900 ;
        RECT 145.950 643.950 150.450 645.300 ;
        RECT 151.800 645.000 154.050 646.200 ;
        RECT 164.400 646.050 165.450 658.950 ;
        RECT 151.800 644.100 153.900 645.000 ;
        RECT 163.950 643.950 166.050 646.050 ;
        RECT 145.950 643.800 148.050 643.950 ;
        RECT 145.950 640.800 148.050 642.900 ;
        RECT 146.400 607.050 147.450 640.800 ;
        RECT 137.400 606.000 142.050 607.050 ;
        RECT 136.950 604.950 142.050 606.000 ;
        RECT 145.950 604.950 148.050 607.050 ;
        RECT 136.950 602.100 139.050 604.950 ;
        RECT 136.950 595.950 139.050 600.900 ;
        RECT 142.950 598.950 145.050 601.050 ;
        RECT 137.400 592.050 138.450 595.950 ;
        RECT 136.950 589.950 139.050 592.050 ;
        RECT 143.400 583.050 144.450 598.950 ;
        RECT 142.950 580.950 145.050 583.050 ;
        RECT 127.950 574.950 130.050 577.050 ;
        RECT 142.950 574.950 145.050 577.050 ;
        RECT 115.950 571.950 118.050 574.050 ;
        RECT 121.950 571.950 124.050 574.050 ;
        RECT 103.950 568.950 106.050 571.050 ;
        RECT 82.950 565.950 85.050 568.050 ;
        RECT 88.950 565.950 91.050 568.050 ;
        RECT 97.950 566.100 100.050 568.200 ;
        RECT 106.950 565.950 112.050 568.050 ;
        RECT 83.400 562.050 84.450 565.950 ;
        RECT 97.950 562.800 100.050 564.900 ;
        RECT 82.950 559.950 85.050 562.050 ;
        RECT 70.950 526.950 73.050 529.050 ;
        RECT 80.400 528.450 85.050 529.050 ;
        RECT 77.400 527.400 85.050 528.450 ;
        RECT 77.400 523.050 78.450 527.400 ;
        RECT 81.000 526.950 85.050 527.400 ;
        RECT 88.950 526.950 91.050 532.050 ;
        RECT 98.400 529.050 99.450 562.800 ;
        RECT 100.950 559.950 103.050 562.050 ;
        RECT 106.950 559.950 112.050 562.050 ;
        RECT 97.950 526.950 100.050 529.050 ;
        RECT 73.950 521.400 78.450 523.050 ;
        RECT 73.950 520.950 78.000 521.400 ;
        RECT 79.950 520.950 82.050 525.900 ;
        RECT 101.400 523.050 102.450 559.950 ;
        RECT 109.950 544.950 112.050 547.050 ;
        RECT 110.400 529.050 111.450 544.950 ;
        RECT 116.400 532.200 117.450 571.950 ;
        RECT 128.400 571.050 129.450 574.950 ;
        RECT 127.950 568.950 130.050 571.050 ;
        RECT 121.950 565.950 127.050 568.050 ;
        RECT 143.400 565.050 144.450 574.950 ;
        RECT 145.950 571.950 148.050 574.050 ;
        RECT 146.400 568.050 147.450 571.950 ;
        RECT 149.400 571.050 150.450 643.950 ;
        RECT 170.400 643.050 171.450 661.950 ;
        RECT 176.400 661.050 177.450 700.950 ;
        RECT 178.950 688.950 181.050 691.050 ;
        RECT 179.400 682.050 180.450 688.950 ;
        RECT 182.400 685.050 183.450 724.950 ;
        RECT 194.400 724.050 195.450 739.950 ;
        RECT 206.400 736.200 207.450 763.950 ;
        RECT 212.400 763.050 213.450 784.950 ;
        RECT 251.400 778.050 252.450 793.950 ;
        RECT 229.950 775.950 232.050 778.050 ;
        RECT 250.950 775.950 253.050 778.050 ;
        RECT 211.950 760.950 214.050 763.050 ;
        RECT 217.950 760.950 220.050 766.050 ;
        RECT 230.400 763.200 231.450 775.950 ;
        RECT 232.950 769.950 235.050 772.050 ;
        RECT 229.950 761.100 232.050 763.200 ;
        RECT 220.950 754.950 223.050 757.050 ;
        RECT 229.950 754.950 232.050 759.900 ;
        RECT 221.400 745.050 222.450 754.950 ;
        RECT 220.950 742.950 223.050 745.050 ;
        RECT 226.950 739.950 229.050 742.050 ;
        RECT 196.950 733.950 199.050 736.050 ;
        RECT 205.950 734.100 208.050 736.200 ;
        RECT 217.950 733.950 220.050 736.050 ;
        RECT 223.950 733.950 226.050 736.050 ;
        RECT 197.400 724.050 198.450 733.950 ;
        RECT 218.400 730.050 219.450 733.950 ;
        RECT 199.950 727.950 202.050 730.050 ;
        RECT 184.950 721.950 190.050 724.050 ;
        RECT 193.950 721.950 196.050 724.050 ;
        RECT 196.950 721.950 199.050 724.050 ;
        RECT 200.400 718.050 201.450 727.950 ;
        RECT 208.950 725.100 211.050 730.050 ;
        RECT 217.950 727.950 220.050 730.050 ;
        RECT 208.950 721.800 211.050 723.900 ;
        RECT 211.950 721.950 217.050 724.050 ;
        RECT 202.950 718.950 205.050 721.050 ;
        RECT 199.950 715.950 202.050 718.050 ;
        RECT 184.950 694.950 187.050 697.050 ;
        RECT 185.400 691.050 186.450 694.950 ;
        RECT 196.950 691.950 199.050 694.050 ;
        RECT 184.950 688.950 187.050 691.050 ;
        RECT 190.950 688.950 193.050 691.050 ;
        RECT 191.400 685.050 192.450 688.950 ;
        RECT 197.400 685.050 198.450 691.950 ;
        RECT 203.400 691.050 204.450 718.950 ;
        RECT 209.400 715.050 210.450 721.800 ;
        RECT 218.400 718.050 219.450 727.950 ;
        RECT 224.400 724.050 225.450 733.950 ;
        RECT 227.400 727.050 228.450 739.950 ;
        RECT 226.950 724.950 229.050 727.050 ;
        RECT 223.950 721.950 226.050 724.050 ;
        RECT 229.950 718.950 232.050 721.050 ;
        RECT 218.400 716.400 223.050 718.050 ;
        RECT 219.000 715.950 223.050 716.400 ;
        RECT 208.950 712.950 211.050 715.050 ;
        RECT 223.950 706.950 226.050 709.050 ;
        RECT 211.950 694.950 214.050 697.050 ;
        RECT 202.950 688.950 205.050 691.050 ;
        RECT 178.950 679.950 181.050 682.050 ;
        RECT 181.950 679.950 184.050 685.050 ;
        RECT 190.950 682.950 193.050 685.050 ;
        RECT 196.950 682.950 199.050 685.050 ;
        RECT 193.950 676.950 196.050 682.050 ;
        RECT 202.950 676.950 205.050 679.050 ;
        RECT 175.950 658.950 178.050 661.050 ;
        RECT 172.950 655.950 175.050 658.050 ;
        RECT 173.400 649.050 174.450 655.950 ;
        RECT 172.950 646.950 175.050 649.050 ;
        RECT 176.400 643.050 177.450 658.950 ;
        RECT 203.400 655.200 204.450 676.950 ;
        RECT 212.400 658.200 213.450 694.950 ;
        RECT 220.950 688.950 223.050 691.050 ;
        RECT 214.950 682.950 220.050 685.050 ;
        RECT 221.400 679.050 222.450 688.950 ;
        RECT 224.400 685.050 225.450 706.950 ;
        RECT 230.400 691.200 231.450 718.950 ;
        RECT 233.400 697.050 234.450 769.950 ;
        RECT 263.400 769.050 264.450 796.950 ;
        RECT 259.950 767.400 264.450 769.050 ;
        RECT 259.950 766.950 264.000 767.400 ;
        RECT 241.950 763.950 244.050 766.050 ;
        RECT 235.950 760.950 241.050 763.050 ;
        RECT 238.950 754.950 241.050 757.050 ;
        RECT 239.400 745.050 240.450 754.950 ;
        RECT 238.950 742.950 241.050 745.050 ;
        RECT 242.400 736.050 243.450 763.950 ;
        RECT 244.950 760.950 247.050 763.050 ;
        RECT 256.950 760.950 259.050 766.050 ;
        RECT 245.400 748.050 246.450 760.950 ;
        RECT 250.950 757.950 256.050 760.050 ;
        RECT 254.400 751.200 255.450 757.950 ;
        RECT 269.400 757.050 270.450 805.950 ;
        RECT 271.950 799.950 277.050 802.050 ;
        RECT 272.400 757.050 273.450 799.950 ;
        RECT 281.400 799.050 282.450 805.950 ;
        RECT 287.400 802.050 288.450 805.950 ;
        RECT 316.950 802.800 319.050 804.900 ;
        RECT 286.950 799.950 289.050 802.050 ;
        RECT 292.950 799.950 295.050 802.050 ;
        RECT 280.950 796.950 283.050 799.050 ;
        RECT 274.950 763.050 277.050 766.050 ;
        RECT 293.400 763.050 294.450 799.950 ;
        RECT 304.950 796.950 307.050 802.050 ;
        RECT 310.950 799.950 313.050 802.050 ;
        RECT 301.950 790.950 304.050 793.050 ;
        RECT 274.950 760.950 280.050 763.050 ;
        RECT 280.950 760.950 283.050 763.050 ;
        RECT 286.950 760.950 292.050 763.050 ;
        RECT 293.400 761.400 298.050 763.050 ;
        RECT 294.000 760.950 298.050 761.400 ;
        RECT 265.950 754.950 268.050 757.050 ;
        RECT 268.800 754.950 270.900 757.050 ;
        RECT 272.100 754.950 274.200 757.050 ;
        RECT 274.950 754.950 280.050 757.050 ;
        RECT 253.950 749.100 256.050 751.200 ;
        RECT 244.950 745.950 247.050 748.050 ;
        RECT 253.950 745.800 256.050 747.900 ;
        RECT 244.950 739.950 247.050 742.050 ;
        RECT 235.950 733.950 238.050 736.050 ;
        RECT 241.950 733.950 244.050 736.050 ;
        RECT 236.400 724.050 237.450 733.950 ;
        RECT 238.950 727.950 244.050 730.050 ;
        RECT 245.400 724.050 246.450 739.950 ;
        RECT 250.950 727.950 253.050 730.050 ;
        RECT 251.400 724.050 252.450 727.950 ;
        RECT 236.400 722.400 241.050 724.050 ;
        RECT 237.000 721.950 241.050 722.400 ;
        RECT 244.950 721.950 247.050 724.050 ;
        RECT 250.950 721.950 253.050 724.050 ;
        RECT 254.400 709.050 255.450 745.800 ;
        RECT 258.000 729.450 262.050 730.050 ;
        RECT 257.400 727.950 262.050 729.450 ;
        RECT 253.950 706.950 256.050 709.050 ;
        RECT 232.950 694.950 235.050 697.050 ;
        RECT 257.400 694.050 258.450 727.950 ;
        RECT 266.400 727.050 267.450 754.950 ;
        RECT 281.400 751.050 282.450 760.950 ;
        RECT 302.400 757.050 303.450 790.950 ;
        RECT 311.400 790.050 312.450 799.950 ;
        RECT 310.950 787.950 313.050 790.050 ;
        RECT 317.400 775.050 318.450 802.800 ;
        RECT 316.950 772.950 319.050 775.050 ;
        RECT 320.400 771.450 321.450 808.950 ;
        RECT 332.400 808.050 333.450 817.950 ;
        RECT 385.950 814.950 388.050 817.050 ;
        RECT 415.950 814.950 418.050 817.050 ;
        RECT 352.950 808.050 355.050 808.200 ;
        RECT 322.950 803.100 325.050 808.050 ;
        RECT 331.950 805.950 334.050 808.050 ;
        RECT 340.950 805.950 343.050 808.050 ;
        RECT 349.950 806.100 355.050 808.050 ;
        RECT 349.950 805.950 354.000 806.100 ;
        RECT 322.950 799.800 325.050 801.900 ;
        RECT 328.950 799.950 331.050 802.050 ;
        RECT 323.400 793.050 324.450 799.800 ;
        RECT 322.950 790.950 325.050 793.050 ;
        RECT 329.400 790.050 330.450 799.950 ;
        RECT 328.950 787.950 331.050 790.050 ;
        RECT 325.950 784.950 328.050 787.050 ;
        RECT 326.400 772.050 327.450 784.950 ;
        RECT 341.400 784.050 342.450 805.950 ;
        RECT 346.950 796.950 349.050 802.050 ;
        RECT 352.950 799.950 355.050 804.900 ;
        RECT 364.950 803.100 367.050 808.050 ;
        RECT 379.950 805.950 382.050 808.050 ;
        RECT 361.950 801.900 366.000 802.050 ;
        RECT 361.950 799.950 367.050 801.900 ;
        RECT 349.950 790.950 352.050 793.050 ;
        RECT 340.950 781.950 343.050 784.050 ;
        RECT 317.400 770.400 321.450 771.450 ;
        RECT 317.400 766.050 318.450 770.400 ;
        RECT 325.950 769.950 328.050 772.050 ;
        RECT 319.950 768.450 324.000 769.050 ;
        RECT 337.950 768.450 342.000 769.050 ;
        RECT 319.950 766.950 324.450 768.450 ;
        RECT 337.950 766.950 342.450 768.450 ;
        RECT 304.950 763.950 307.050 766.050 ;
        RECT 292.950 754.950 295.050 757.050 ;
        RECT 301.950 754.950 304.050 757.050 ;
        RECT 293.400 751.050 294.450 754.950 ;
        RECT 280.950 748.950 283.050 751.050 ;
        RECT 292.950 748.950 295.050 751.050 ;
        RECT 305.400 742.050 306.450 763.950 ;
        RECT 310.950 760.950 313.050 763.050 ;
        RECT 316.950 761.100 319.050 766.050 ;
        RECT 311.400 750.450 312.450 760.950 ;
        RECT 313.950 759.900 318.000 760.050 ;
        RECT 313.950 757.950 319.050 759.900 ;
        RECT 316.950 757.800 319.050 757.950 ;
        RECT 311.400 749.400 315.450 750.450 ;
        RECT 298.950 739.950 301.050 742.050 ;
        RECT 304.950 739.950 307.050 742.050 ;
        RECT 295.950 733.950 298.050 736.050 ;
        RECT 277.800 727.950 279.900 730.050 ;
        RECT 280.950 727.950 283.050 730.050 ;
        RECT 289.950 727.950 295.050 730.050 ;
        RECT 265.950 724.950 268.050 727.050 ;
        RECT 271.950 724.950 274.050 727.050 ;
        RECT 259.950 721.950 265.050 724.050 ;
        RECT 268.950 721.950 271.050 724.050 ;
        RECT 256.950 691.950 259.050 694.050 ;
        RECT 229.950 689.100 232.050 691.200 ;
        RECT 238.950 688.950 241.050 691.050 ;
        RECT 229.950 685.800 232.050 687.900 ;
        RECT 223.950 679.950 226.050 685.050 ;
        RECT 214.950 676.950 217.050 679.050 ;
        RECT 220.950 676.950 223.050 679.050 ;
        RECT 211.950 656.100 214.050 658.200 ;
        RECT 202.950 653.100 205.050 655.200 ;
        RECT 211.950 652.800 214.050 654.900 ;
        RECT 184.950 649.950 187.050 652.050 ;
        RECT 181.950 646.950 184.050 649.050 ;
        RECT 182.400 643.050 183.450 646.950 ;
        RECT 160.950 640.950 163.050 643.050 ;
        RECT 169.950 640.950 172.050 643.050 ;
        RECT 175.950 640.950 178.050 643.050 ;
        RECT 181.950 640.950 184.050 643.050 ;
        RECT 154.950 625.950 157.050 628.050 ;
        RECT 155.400 601.050 156.450 625.950 ;
        RECT 161.400 622.050 162.450 640.950 ;
        RECT 160.950 619.950 163.050 622.050 ;
        RECT 157.950 613.950 160.050 616.050 ;
        RECT 158.400 607.050 159.450 613.950 ;
        RECT 170.400 607.050 171.450 640.950 ;
        RECT 176.400 628.050 177.450 640.950 ;
        RECT 175.950 625.950 178.050 628.050 ;
        RECT 178.950 619.950 181.050 622.050 ;
        RECT 157.950 604.950 160.050 607.050 ;
        RECT 163.950 604.950 169.050 607.050 ;
        RECT 169.950 604.950 172.050 607.050 ;
        RECT 154.950 598.950 157.050 601.050 ;
        RECT 158.400 597.450 159.450 604.950 ;
        RECT 175.950 601.950 178.050 604.050 ;
        RECT 155.400 596.400 159.450 597.450 ;
        RECT 155.400 574.050 156.450 596.400 ;
        RECT 160.950 595.950 163.050 601.050 ;
        RECT 166.950 598.950 169.050 601.050 ;
        RECT 167.400 592.050 168.450 598.950 ;
        RECT 169.950 592.950 172.050 595.050 ;
        RECT 166.950 589.950 169.050 592.050 ;
        RECT 167.400 577.050 168.450 589.950 ;
        RECT 166.950 574.950 169.050 577.050 ;
        RECT 154.950 571.950 157.050 574.050 ;
        RECT 170.400 573.450 171.450 592.950 ;
        RECT 167.400 572.400 171.450 573.450 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 145.950 565.950 148.050 568.050 ;
        RECT 136.950 559.950 139.050 565.050 ;
        RECT 142.950 562.950 145.050 565.050 ;
        RECT 139.950 544.950 142.050 547.050 ;
        RECT 133.950 535.950 136.050 538.050 ;
        RECT 115.950 530.100 118.050 532.200 ;
        RECT 103.950 526.950 106.050 529.050 ;
        RECT 109.950 526.950 112.050 529.050 ;
        RECT 82.950 520.950 88.050 523.050 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 70.950 517.950 73.050 520.050 ;
        RECT 71.400 496.050 72.450 517.950 ;
        RECT 76.950 514.950 79.050 517.050 ;
        RECT 70.950 493.950 73.050 496.050 ;
        RECT 77.400 490.050 78.450 514.950 ;
        RECT 104.400 502.050 105.450 526.950 ;
        RECT 115.950 526.800 118.050 528.900 ;
        RECT 106.950 523.950 109.050 526.050 ;
        RECT 107.400 517.050 108.450 523.950 ;
        RECT 116.400 523.050 117.450 526.800 ;
        RECT 121.950 523.950 124.050 529.050 ;
        RECT 127.950 528.450 132.000 529.050 ;
        RECT 127.950 526.950 132.450 528.450 ;
        RECT 112.950 520.950 115.050 523.050 ;
        RECT 116.400 521.400 121.050 523.050 ;
        RECT 117.000 520.950 121.050 521.400 ;
        RECT 124.950 520.950 127.050 523.050 ;
        RECT 106.950 514.950 109.050 517.050 ;
        RECT 113.400 511.050 114.450 520.950 ;
        RECT 112.950 508.950 115.050 511.050 ;
        RECT 97.950 499.950 100.050 502.050 ;
        RECT 103.950 499.950 106.050 502.050 ;
        RECT 79.950 493.950 85.050 496.050 ;
        RECT 98.400 493.050 99.450 499.950 ;
        RECT 109.950 493.950 112.050 496.050 ;
        RECT 115.950 493.950 118.050 496.050 ;
        RECT 118.950 493.950 124.050 496.050 ;
        RECT 97.950 490.950 100.050 493.050 ;
        RECT 76.950 487.950 79.050 490.050 ;
        RECT 82.950 484.950 85.050 490.050 ;
        RECT 100.950 487.950 103.050 490.050 ;
        RECT 94.950 484.950 97.050 487.050 ;
        RECT 73.950 469.950 76.050 472.050 ;
        RECT 64.800 463.950 66.900 466.050 ;
        RECT 68.100 463.950 70.200 466.050 ;
        RECT 65.400 454.050 66.450 463.950 ;
        RECT 74.400 457.050 75.450 469.950 ;
        RECT 82.950 463.950 85.050 466.050 ;
        RECT 73.950 454.950 76.050 457.050 ;
        RECT 64.950 451.950 67.050 454.050 ;
        RECT 70.950 448.950 76.050 451.050 ;
        RECT 79.950 448.950 82.050 454.050 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 65.400 442.050 66.450 445.950 ;
        RECT 67.950 442.950 70.050 448.050 ;
        RECT 73.950 442.950 76.050 445.050 ;
        RECT 64.950 439.950 67.050 442.050 ;
        RECT 70.950 439.950 73.050 442.050 ;
        RECT 67.950 436.950 70.050 439.050 ;
        RECT 61.950 419.100 64.050 421.200 ;
        RECT 68.400 418.050 69.450 436.950 ;
        RECT 46.950 415.950 49.050 418.050 ;
        RECT 58.950 415.950 61.050 418.050 ;
        RECT 43.950 412.950 46.050 415.050 ;
        RECT 47.400 412.050 48.450 415.950 ;
        RECT 61.950 415.800 64.050 417.900 ;
        RECT 67.950 415.950 70.050 418.050 ;
        RECT 38.400 410.400 42.450 411.450 ;
        RECT 32.400 406.050 33.450 409.950 ;
        RECT 31.950 403.950 34.050 406.050 ;
        RECT 34.950 379.950 37.050 382.050 ;
        RECT 13.950 370.950 16.050 376.050 ;
        RECT 25.950 373.950 28.050 376.050 ;
        RECT 19.950 370.950 25.050 373.050 ;
        RECT 16.950 364.950 22.050 367.050 ;
        RECT 7.950 340.950 10.050 343.050 ;
        RECT 26.400 340.050 27.450 373.950 ;
        RECT 35.400 370.050 36.450 379.950 ;
        RECT 38.400 373.050 39.450 410.400 ;
        RECT 46.950 409.950 49.050 412.050 ;
        RECT 40.950 406.950 43.050 409.050 ;
        RECT 41.400 382.200 42.450 406.950 ;
        RECT 46.950 403.950 52.050 406.050 ;
        RECT 62.400 384.450 63.450 415.800 ;
        RECT 64.950 409.950 67.050 412.050 ;
        RECT 65.400 391.050 66.450 409.950 ;
        RECT 71.400 409.050 72.450 439.950 ;
        RECT 74.400 436.050 75.450 442.950 ;
        RECT 83.400 442.050 84.450 463.950 ;
        RECT 91.950 460.950 94.050 463.050 ;
        RECT 92.400 451.050 93.450 460.950 ;
        RECT 95.400 457.050 96.450 484.950 ;
        RECT 101.400 484.050 102.450 487.950 ;
        RECT 100.950 481.950 103.050 484.050 ;
        RECT 103.950 481.950 106.050 487.050 ;
        RECT 110.400 484.050 111.450 493.950 ;
        RECT 109.950 481.950 112.050 484.050 ;
        RECT 100.950 463.950 103.050 466.050 ;
        RECT 94.950 451.950 97.050 457.050 ;
        RECT 88.950 445.950 91.050 451.050 ;
        RECT 91.950 448.950 94.050 451.050 ;
        RECT 94.950 442.950 97.050 445.050 ;
        RECT 82.950 439.950 85.050 442.050 ;
        RECT 73.950 433.950 76.050 436.050 ;
        RECT 95.400 430.050 96.450 442.950 ;
        RECT 94.950 427.950 97.050 430.050 ;
        RECT 76.950 415.950 79.050 421.050 ;
        RECT 77.400 409.050 78.450 415.950 ;
        RECT 101.400 415.050 102.450 463.950 ;
        RECT 106.950 447.450 109.050 451.050 ;
        RECT 112.950 448.950 115.050 454.050 ;
        RECT 106.950 447.000 111.450 447.450 ;
        RECT 107.400 446.400 111.450 447.000 ;
        RECT 110.400 418.050 111.450 446.400 ;
        RECT 116.400 445.050 117.450 493.950 ;
        RECT 125.400 492.450 126.450 520.950 ;
        RECT 131.400 511.050 132.450 526.950 ;
        RECT 130.950 508.950 133.050 511.050 ;
        RECT 127.950 499.950 130.050 502.050 ;
        RECT 122.400 491.400 126.450 492.450 ;
        RECT 118.950 484.950 121.050 490.050 ;
        RECT 122.400 463.050 123.450 491.400 ;
        RECT 128.400 490.050 129.450 499.950 ;
        RECT 130.950 491.100 133.050 496.050 ;
        RECT 124.950 488.400 129.450 490.050 ;
        RECT 124.950 487.950 129.000 488.400 ;
        RECT 130.950 487.800 133.050 489.900 ;
        RECT 131.400 484.050 132.450 487.800 ;
        RECT 130.950 481.950 133.050 484.050 ;
        RECT 134.400 481.050 135.450 535.950 ;
        RECT 140.400 493.200 141.450 544.950 ;
        RECT 149.400 538.050 150.450 568.950 ;
        RECT 167.400 547.050 168.450 572.400 ;
        RECT 176.400 571.200 177.450 601.950 ;
        RECT 179.400 601.050 180.450 619.950 ;
        RECT 181.950 604.950 184.050 610.050 ;
        RECT 185.400 604.200 186.450 649.950 ;
        RECT 202.950 649.800 205.050 651.900 ;
        RECT 190.950 643.950 193.050 646.050 ;
        RECT 187.950 613.950 190.050 616.050 ;
        RECT 188.400 607.050 189.450 613.950 ;
        RECT 187.950 604.950 190.050 607.050 ;
        RECT 184.950 602.100 187.050 604.200 ;
        RECT 191.400 604.050 192.450 643.950 ;
        RECT 203.400 628.050 204.450 649.800 ;
        RECT 212.400 646.050 213.450 652.800 ;
        RECT 215.400 652.050 216.450 676.950 ;
        RECT 230.400 670.050 231.450 685.800 ;
        RECT 239.400 685.050 240.450 688.950 ;
        RECT 241.950 685.950 244.050 691.050 ;
        RECT 247.950 685.950 250.050 688.050 ;
        RECT 238.950 682.950 241.050 685.050 ;
        RECT 232.950 679.950 238.050 682.050 ;
        RECT 248.400 679.050 249.450 685.950 ;
        RECT 257.400 685.050 258.450 691.950 ;
        RECT 265.950 690.450 268.050 691.050 ;
        RECT 269.400 690.450 270.450 721.950 ;
        RECT 272.400 715.050 273.450 724.950 ;
        RECT 278.400 724.050 279.450 727.950 ;
        RECT 277.950 721.950 280.050 724.050 ;
        RECT 271.950 712.950 274.050 715.050 ;
        RECT 271.950 703.950 274.050 709.050 ;
        RECT 277.950 706.950 280.050 709.050 ;
        RECT 274.950 697.950 277.050 700.050 ;
        RECT 271.950 694.950 274.050 697.050 ;
        RECT 265.950 689.400 270.450 690.450 ;
        RECT 265.950 688.950 268.050 689.400 ;
        RECT 266.400 685.050 267.450 688.950 ;
        RECT 272.400 685.050 273.450 694.950 ;
        RECT 275.400 685.050 276.450 697.950 ;
        RECT 278.400 691.050 279.450 706.950 ;
        RECT 277.950 688.950 280.050 691.050 ;
        RECT 281.400 685.050 282.450 727.950 ;
        RECT 296.400 724.050 297.450 733.950 ;
        RECT 283.950 721.950 289.050 724.050 ;
        RECT 292.950 722.400 297.450 724.050 ;
        RECT 292.950 721.950 297.000 722.400 ;
        RECT 287.400 718.050 288.450 721.950 ;
        RECT 299.400 720.450 300.450 739.950 ;
        RECT 307.950 733.950 310.050 736.050 ;
        RECT 304.950 727.950 307.050 730.050 ;
        RECT 305.400 724.050 306.450 727.950 ;
        RECT 308.400 727.050 309.450 733.950 ;
        RECT 314.400 730.050 315.450 749.400 ;
        RECT 313.950 727.950 316.050 730.050 ;
        RECT 307.950 724.950 310.050 727.050 ;
        RECT 304.950 721.950 307.050 724.050 ;
        RECT 296.400 719.400 300.450 720.450 ;
        RECT 286.950 717.450 289.050 718.050 ;
        RECT 286.950 716.400 291.450 717.450 ;
        RECT 286.950 715.950 289.050 716.400 ;
        RECT 256.950 682.950 259.050 685.050 ;
        RECT 265.950 682.950 268.050 685.050 ;
        RECT 271.950 682.950 274.050 685.050 ;
        RECT 274.950 682.950 277.050 685.050 ;
        RECT 280.950 682.950 283.050 685.050 ;
        RECT 283.950 682.950 289.050 685.050 ;
        RECT 241.950 676.950 244.050 679.050 ;
        RECT 248.400 676.950 253.050 679.050 ;
        RECT 256.950 676.950 259.050 679.050 ;
        RECT 262.950 676.950 265.050 679.050 ;
        RECT 229.950 667.950 232.050 670.050 ;
        RECT 217.950 661.950 220.050 664.050 ;
        RECT 214.950 649.950 217.050 652.050 ;
        RECT 205.950 643.950 208.050 646.050 ;
        RECT 211.950 643.950 214.050 646.050 ;
        RECT 206.400 640.050 207.450 643.950 ;
        RECT 205.950 637.950 208.050 640.050 ;
        RECT 202.950 625.950 205.050 628.050 ;
        RECT 202.950 619.950 205.050 622.050 ;
        RECT 199.950 616.950 202.050 619.050 ;
        RECT 193.950 610.950 196.050 613.050 ;
        RECT 178.950 598.950 181.050 601.050 ;
        RECT 184.950 598.800 187.050 600.900 ;
        RECT 190.950 598.950 193.050 604.050 ;
        RECT 185.400 595.050 186.450 598.800 ;
        RECT 191.400 597.450 192.450 598.950 ;
        RECT 188.400 596.400 192.450 597.450 ;
        RECT 184.950 592.950 187.050 595.050 ;
        RECT 188.400 592.050 189.450 596.400 ;
        RECT 187.950 589.950 190.050 592.050 ;
        RECT 194.400 586.050 195.450 610.950 ;
        RECT 200.400 607.050 201.450 616.950 ;
        RECT 203.400 613.050 204.450 619.950 ;
        RECT 218.400 616.200 219.450 661.950 ;
        RECT 229.950 655.950 232.050 658.050 ;
        RECT 230.400 652.050 231.450 655.950 ;
        RECT 229.950 649.950 232.050 652.050 ;
        RECT 235.950 651.450 240.000 652.050 ;
        RECT 235.950 649.950 240.450 651.450 ;
        RECT 226.950 640.950 229.050 646.050 ;
        RECT 232.950 643.950 235.050 646.050 ;
        RECT 233.400 634.050 234.450 643.950 ;
        RECT 232.950 631.950 235.050 634.050 ;
        RECT 239.400 628.050 240.450 649.950 ;
        RECT 242.400 646.050 243.450 676.950 ;
        RECT 248.400 652.050 249.450 676.950 ;
        RECT 257.400 661.050 258.450 676.950 ;
        RECT 259.950 673.950 262.050 676.050 ;
        RECT 256.950 658.950 259.050 661.050 ;
        RECT 247.950 649.950 250.050 652.050 ;
        RECT 256.950 649.950 259.050 652.050 ;
        RECT 241.950 643.950 244.050 646.050 ;
        RECT 250.950 643.950 256.050 646.050 ;
        RECT 244.950 640.950 247.050 643.050 ;
        RECT 232.950 625.950 235.050 628.050 ;
        RECT 238.950 625.950 241.050 628.050 ;
        RECT 211.950 613.950 214.050 616.050 ;
        RECT 217.950 614.100 220.050 616.200 ;
        RECT 223.950 613.950 226.050 616.050 ;
        RECT 202.950 610.950 205.050 613.050 ;
        RECT 199.950 604.950 202.050 607.050 ;
        RECT 196.950 592.950 199.050 595.050 ;
        RECT 178.950 583.950 181.050 586.050 ;
        RECT 193.950 583.950 196.050 586.050 ;
        RECT 169.950 568.950 172.050 571.050 ;
        RECT 175.950 569.100 178.050 571.200 ;
        RECT 170.400 562.050 171.450 568.950 ;
        RECT 169.950 559.950 172.050 562.050 ;
        RECT 166.950 544.950 169.050 547.050 ;
        RECT 166.950 538.950 169.050 541.050 ;
        RECT 148.950 535.950 151.050 538.050 ;
        RECT 154.950 535.950 157.050 538.050 ;
        RECT 142.950 529.950 145.050 535.050 ;
        RECT 148.950 529.950 151.050 532.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 143.400 502.050 144.450 523.950 ;
        RECT 145.950 505.950 148.050 508.050 ;
        RECT 142.950 499.950 145.050 502.050 ;
        RECT 146.400 496.050 147.450 505.950 ;
        RECT 149.400 505.050 150.450 529.950 ;
        RECT 151.950 526.950 154.050 529.050 ;
        RECT 148.950 502.950 151.050 505.050 ;
        RECT 152.400 499.050 153.450 526.950 ;
        RECT 151.950 496.950 154.050 499.050 ;
        RECT 145.950 493.950 148.050 496.050 ;
        RECT 139.950 491.100 142.050 493.200 ;
        RECT 155.400 493.050 156.450 535.950 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 157.950 520.950 160.050 523.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 139.950 484.950 142.050 489.900 ;
        RECT 133.950 478.950 136.050 481.050 ;
        RECT 121.950 460.950 124.050 463.050 ;
        RECT 151.950 460.950 154.050 463.050 ;
        RECT 127.950 448.950 130.050 454.050 ;
        RECT 133.950 445.950 136.050 451.050 ;
        RECT 139.950 448.950 142.050 451.050 ;
        RECT 115.950 442.950 118.050 445.050 ;
        RECT 121.950 442.950 127.050 445.050 ;
        RECT 130.950 442.950 133.050 445.050 ;
        RECT 131.400 436.050 132.450 442.950 ;
        RECT 130.950 433.950 133.050 436.050 ;
        RECT 118.950 421.950 121.050 424.050 ;
        RECT 106.950 415.950 109.050 418.050 ;
        RECT 109.950 415.950 112.050 418.050 ;
        RECT 82.950 412.950 85.050 415.050 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 70.950 403.950 73.050 409.050 ;
        RECT 77.400 407.400 82.050 409.050 ;
        RECT 78.000 406.950 82.050 407.400 ;
        RECT 83.400 394.050 84.450 412.950 ;
        RECT 107.400 412.050 108.450 415.950 ;
        RECT 119.400 412.050 120.450 421.950 ;
        RECT 140.400 421.200 141.450 448.950 ;
        RECT 152.400 445.050 153.450 460.950 ;
        RECT 158.400 454.050 159.450 520.950 ;
        RECT 164.400 520.050 165.450 526.950 ;
        RECT 167.400 523.050 168.450 538.950 ;
        RECT 170.400 538.050 171.450 559.950 ;
        RECT 179.400 541.050 180.450 583.950 ;
        RECT 184.950 580.950 187.050 583.050 ;
        RECT 181.950 568.950 184.050 571.050 ;
        RECT 178.950 538.950 181.050 541.050 ;
        RECT 169.950 535.950 172.050 538.050 ;
        RECT 182.400 535.050 183.450 568.950 ;
        RECT 185.400 562.050 186.450 580.950 ;
        RECT 187.950 571.950 190.050 574.050 ;
        RECT 188.400 565.050 189.450 571.950 ;
        RECT 197.400 571.050 198.450 592.950 ;
        RECT 200.400 583.050 201.450 604.950 ;
        RECT 205.950 601.950 208.050 604.050 ;
        RECT 202.950 598.950 205.050 601.050 ;
        RECT 199.950 580.950 202.050 583.050 ;
        RECT 203.400 574.050 204.450 598.950 ;
        RECT 206.400 598.050 207.450 601.950 ;
        RECT 205.950 595.950 208.050 598.050 ;
        RECT 208.950 580.950 211.050 583.050 ;
        RECT 202.950 571.950 205.050 574.050 ;
        RECT 205.950 571.950 208.050 574.050 ;
        RECT 196.950 568.950 199.050 571.050 ;
        RECT 188.400 563.400 193.050 565.050 ;
        RECT 189.000 562.950 193.050 563.400 ;
        RECT 196.950 562.950 199.050 565.050 ;
        RECT 184.950 559.950 187.050 562.050 ;
        RECT 191.400 559.050 192.450 562.950 ;
        RECT 190.950 556.950 193.050 559.050 ;
        RECT 197.400 556.050 198.450 562.950 ;
        RECT 199.950 559.950 202.050 562.050 ;
        RECT 184.950 553.950 187.050 556.050 ;
        RECT 196.950 553.950 199.050 556.050 ;
        RECT 181.950 532.950 184.050 535.050 ;
        RECT 169.950 528.450 174.000 529.050 ;
        RECT 169.950 526.950 174.450 528.450 ;
        RECT 178.950 526.950 184.050 529.050 ;
        RECT 173.400 523.050 174.450 526.950 ;
        RECT 166.950 520.950 169.050 523.050 ;
        RECT 172.950 520.950 175.050 523.050 ;
        RECT 163.950 517.950 166.050 520.050 ;
        RECT 164.400 508.050 165.450 517.950 ;
        RECT 163.950 505.950 166.050 508.050 ;
        RECT 185.400 502.050 186.450 553.950 ;
        RECT 194.100 547.950 196.200 550.050 ;
        RECT 187.950 538.950 190.050 541.050 ;
        RECT 188.400 529.050 189.450 538.950 ;
        RECT 187.950 526.950 190.050 529.050 ;
        RECT 184.950 499.950 187.050 502.050 ;
        RECT 160.950 490.950 166.050 493.050 ;
        RECT 169.950 487.950 172.050 493.050 ;
        RECT 175.950 490.950 178.050 496.050 ;
        RECT 160.950 463.950 163.050 466.050 ;
        RECT 157.950 451.950 160.050 454.050 ;
        RECT 161.400 451.050 162.450 463.950 ;
        RECT 166.950 460.950 169.050 463.050 ;
        RECT 167.400 451.050 168.450 460.950 ;
        RECT 170.400 454.050 171.450 487.950 ;
        RECT 178.950 484.950 181.050 487.050 ;
        RECT 184.950 484.950 187.050 490.050 ;
        RECT 179.400 481.050 180.450 484.950 ;
        RECT 178.950 478.950 181.050 481.050 ;
        RECT 169.950 451.950 172.050 454.050 ;
        RECT 160.950 448.950 163.050 451.050 ;
        RECT 166.950 448.950 169.050 451.050 ;
        RECT 175.950 448.950 178.050 451.050 ;
        RECT 151.950 442.950 154.050 445.050 ;
        RECT 157.950 442.950 160.050 448.050 ;
        RECT 148.950 439.950 151.050 442.050 ;
        RECT 121.950 415.950 124.050 421.050 ;
        RECT 139.950 419.100 142.050 421.200 ;
        RECT 103.950 410.400 108.450 412.050 ;
        RECT 103.950 409.950 108.000 410.400 ;
        RECT 118.950 409.950 121.050 412.050 ;
        RECT 124.950 409.950 127.050 415.050 ;
        RECT 130.950 409.950 133.050 415.050 ;
        RECT 139.950 412.950 142.050 417.900 ;
        RECT 145.950 415.950 148.050 418.050 ;
        RECT 85.950 403.950 88.050 409.050 ;
        RECT 94.950 406.950 97.050 409.050 ;
        RECT 73.950 391.950 76.050 394.050 ;
        RECT 82.950 391.950 85.050 394.050 ;
        RECT 64.950 388.950 67.050 391.050 ;
        RECT 59.400 383.400 63.450 384.450 ;
        RECT 40.950 380.100 43.050 382.200 ;
        RECT 40.950 373.950 43.050 378.900 ;
        RECT 37.950 370.950 40.050 373.050 ;
        RECT 41.400 370.050 42.450 373.950 ;
        RECT 55.950 370.950 58.050 373.050 ;
        RECT 34.950 364.950 37.050 370.050 ;
        RECT 40.950 367.950 43.050 370.050 ;
        RECT 49.950 367.950 55.050 370.050 ;
        RECT 56.400 367.050 57.450 370.950 ;
        RECT 55.950 364.950 58.050 367.050 ;
        RECT 43.950 361.950 46.050 364.050 ;
        RECT 37.950 355.950 40.050 358.050 ;
        RECT 38.400 340.050 39.450 355.950 ;
        RECT 44.400 342.450 45.450 361.950 ;
        RECT 59.400 355.050 60.450 383.400 ;
        RECT 70.950 376.950 73.050 379.050 ;
        RECT 61.950 367.950 64.050 373.050 ;
        RECT 71.400 367.050 72.450 376.950 ;
        RECT 67.950 365.400 72.450 367.050 ;
        RECT 67.950 364.950 72.000 365.400 ;
        RECT 74.400 361.050 75.450 391.950 ;
        RECT 79.950 388.950 82.050 391.050 ;
        RECT 76.950 364.950 79.050 370.050 ;
        RECT 73.950 358.950 76.050 361.050 ;
        RECT 49.950 352.950 52.050 355.050 ;
        RECT 58.950 352.950 61.050 355.050 ;
        RECT 41.400 341.400 45.450 342.450 ;
        RECT 26.400 337.950 31.050 340.050 ;
        RECT 37.950 337.950 40.050 340.050 ;
        RECT 4.950 334.950 7.050 337.050 ;
        RECT 5.400 310.050 6.450 334.950 ;
        RECT 7.950 328.950 10.050 334.050 ;
        RECT 26.400 331.050 27.450 337.950 ;
        RECT 41.400 337.050 42.450 341.400 ;
        RECT 43.950 337.950 46.050 340.050 ;
        RECT 46.950 337.950 49.050 343.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 44.400 334.050 45.450 337.950 ;
        RECT 50.400 334.050 51.450 352.950 ;
        RECT 58.950 340.950 61.050 343.050 ;
        RECT 59.400 334.050 60.450 340.950 ;
        RECT 61.950 334.950 64.050 340.050 ;
        RECT 80.400 334.050 81.450 388.950 ;
        RECT 88.950 385.950 91.050 388.050 ;
        RECT 82.950 379.950 85.050 382.050 ;
        RECT 83.400 373.050 84.450 379.950 ;
        RECT 89.400 373.050 90.450 385.950 ;
        RECT 95.400 373.050 96.450 406.950 ;
        RECT 106.950 403.950 109.050 409.050 ;
        RECT 125.400 406.050 126.450 409.950 ;
        RECT 124.950 403.950 127.050 406.050 ;
        RECT 139.950 391.950 142.050 394.050 ;
        RECT 121.950 388.950 124.050 391.050 ;
        RECT 103.950 385.950 106.050 388.050 ;
        RECT 97.950 373.950 100.050 379.050 ;
        RECT 82.950 370.950 85.050 373.050 ;
        RECT 88.950 370.950 91.050 373.050 ;
        RECT 94.950 370.950 97.050 373.050 ;
        RECT 95.400 367.050 96.450 370.950 ;
        RECT 104.400 370.050 105.450 385.950 ;
        RECT 109.950 379.050 112.050 382.050 ;
        RECT 112.950 379.050 115.050 379.200 ;
        RECT 109.950 377.100 115.050 379.050 ;
        RECT 109.950 376.950 114.000 377.100 ;
        RECT 118.950 376.950 121.050 379.050 ;
        RECT 106.950 370.950 109.050 376.050 ;
        RECT 112.950 373.800 115.050 375.900 ;
        RECT 103.950 367.950 106.050 370.050 ;
        RECT 85.950 364.950 91.050 367.050 ;
        RECT 94.950 364.950 97.050 367.050 ;
        RECT 82.950 358.950 85.050 361.050 ;
        RECT 83.400 340.200 84.450 358.950 ;
        RECT 97.950 352.950 100.050 355.050 ;
        RECT 82.950 338.100 85.050 340.200 ;
        RECT 84.000 336.900 88.050 337.050 ;
        RECT 82.950 334.950 88.050 336.900 ;
        RECT 82.950 334.800 85.050 334.950 ;
        RECT 37.950 333.450 40.050 334.050 ;
        RECT 43.950 333.450 46.050 334.050 ;
        RECT 37.950 332.400 46.050 333.450 ;
        RECT 37.950 331.950 40.050 332.400 ;
        RECT 43.950 331.950 46.050 332.400 ;
        RECT 49.950 331.950 52.050 334.050 ;
        RECT 58.950 331.950 61.050 334.050 ;
        RECT 13.950 328.950 16.050 331.050 ;
        RECT 25.950 328.950 28.050 331.050 ;
        RECT 40.950 328.950 43.050 331.050 ;
        RECT 14.400 325.050 15.450 328.950 ;
        RECT 13.950 322.950 16.050 325.050 ;
        RECT 37.950 322.950 40.050 325.050 ;
        RECT 4.950 307.950 7.050 310.050 ;
        RECT 13.950 307.950 16.050 310.050 ;
        RECT 34.950 307.950 37.050 310.050 ;
        RECT 7.950 302.400 10.050 304.500 ;
        RECT 4.950 298.950 7.050 301.050 ;
        RECT 5.400 286.050 6.450 298.950 ;
        RECT 4.950 283.950 7.050 286.050 ;
        RECT 8.700 282.600 9.900 302.400 ;
        RECT 14.400 301.050 15.450 307.950 ;
        RECT 28.950 303.300 31.050 305.400 ;
        RECT 13.950 298.950 16.050 301.050 ;
        RECT 28.950 299.700 30.150 303.300 ;
        RECT 28.950 297.600 31.050 299.700 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 13.950 283.950 16.050 286.050 ;
        RECT 7.950 280.500 10.050 282.600 ;
        RECT 14.400 274.050 15.450 283.950 ;
        RECT 20.400 283.050 21.450 289.950 ;
        RECT 19.950 280.950 22.050 283.050 ;
        RECT 28.950 282.600 30.150 297.600 ;
        RECT 35.400 289.050 36.450 307.950 ;
        RECT 31.950 287.400 36.450 289.050 ;
        RECT 38.400 298.050 39.450 322.950 ;
        RECT 41.400 301.200 42.450 328.950 ;
        RECT 50.400 328.050 51.450 331.950 ;
        RECT 64.950 328.950 67.050 334.050 ;
        RECT 79.950 328.950 82.050 334.050 ;
        RECT 91.950 331.950 94.050 337.050 ;
        RECT 49.950 325.950 52.050 328.050 ;
        RECT 55.950 325.950 61.050 328.050 ;
        RECT 73.950 322.950 76.050 328.050 ;
        RECT 88.950 319.950 91.050 322.050 ;
        RECT 46.950 304.950 49.050 307.050 ;
        RECT 40.950 299.100 43.050 301.200 ;
        RECT 47.400 298.050 48.450 304.950 ;
        RECT 58.950 303.300 61.050 305.400 ;
        RECT 52.950 298.950 55.050 301.050 ;
        RECT 59.850 299.700 61.050 303.300 ;
        RECT 79.950 302.400 82.050 304.500 ;
        RECT 38.400 297.900 42.000 298.050 ;
        RECT 38.400 295.950 43.050 297.900 ;
        RECT 46.950 295.950 49.050 298.050 ;
        RECT 31.950 286.950 36.000 287.400 ;
        RECT 13.950 271.950 16.050 274.050 ;
        RECT 7.950 266.400 10.050 268.500 ;
        RECT 4.950 262.950 7.050 265.050 ;
        RECT 5.400 250.050 6.450 262.950 ;
        RECT 4.950 247.950 7.050 250.050 ;
        RECT 8.700 246.600 9.900 266.400 ;
        RECT 13.950 265.950 16.050 268.050 ;
        RECT 14.400 259.050 15.450 265.950 ;
        RECT 20.400 259.050 21.450 280.950 ;
        RECT 28.950 280.500 31.050 282.600 ;
        RECT 38.400 274.050 39.450 295.950 ;
        RECT 40.950 295.800 43.050 295.950 ;
        RECT 53.400 295.050 54.450 298.950 ;
        RECT 58.950 297.600 61.050 299.700 ;
        RECT 43.950 292.950 46.050 295.050 ;
        RECT 52.950 292.950 55.050 295.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 22.950 271.950 25.050 274.050 ;
        RECT 37.950 271.950 40.050 274.050 ;
        RECT 13.950 256.950 16.050 259.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 13.950 247.950 16.050 250.050 ;
        RECT 7.950 244.500 10.050 246.600 ;
        RECT 14.400 217.050 15.450 247.950 ;
        RECT 23.400 217.050 24.450 271.950 ;
        RECT 28.950 266.400 31.050 268.500 ;
        RECT 28.950 251.400 30.150 266.400 ;
        RECT 41.400 264.450 42.450 289.950 ;
        RECT 38.400 263.400 42.450 264.450 ;
        RECT 31.950 259.950 37.050 262.050 ;
        RECT 38.400 256.200 39.450 263.400 ;
        RECT 44.400 262.050 45.450 292.950 ;
        RECT 49.950 286.950 52.050 289.050 ;
        RECT 52.950 286.950 58.050 289.050 ;
        RECT 46.950 265.950 49.050 268.050 ;
        RECT 47.400 262.050 48.450 265.950 ;
        RECT 40.950 259.950 43.050 262.050 ;
        RECT 43.800 259.950 45.900 262.050 ;
        RECT 46.950 259.950 49.050 262.050 ;
        RECT 37.950 254.100 40.050 256.200 ;
        RECT 28.950 249.300 31.050 251.400 ;
        RECT 37.950 250.800 40.050 252.900 ;
        RECT 28.950 245.700 30.150 249.300 ;
        RECT 34.950 247.950 37.050 250.050 ;
        RECT 28.950 243.600 31.050 245.700 ;
        RECT 1.950 214.950 4.050 217.050 ;
        RECT 10.950 214.950 13.050 217.050 ;
        RECT 13.950 214.950 16.050 217.050 ;
        RECT 19.950 215.400 24.450 217.050 ;
        RECT 19.950 214.950 24.000 215.400 ;
        RECT 11.400 211.050 12.450 214.950 ;
        RECT 35.400 214.050 36.450 247.950 ;
        RECT 38.400 220.050 39.450 250.800 ;
        RECT 37.950 217.950 40.050 220.050 ;
        RECT 41.400 217.050 42.450 259.950 ;
        RECT 43.950 253.950 49.050 256.050 ;
        RECT 50.400 250.050 51.450 286.950 ;
        RECT 59.850 282.600 61.050 297.600 ;
        RECT 67.950 289.950 70.050 292.050 ;
        RECT 73.950 289.950 76.050 295.050 ;
        RECT 68.400 283.050 69.450 289.950 ;
        RECT 58.950 280.500 61.050 282.600 ;
        RECT 67.950 280.950 70.050 283.050 ;
        RECT 80.100 282.600 81.300 302.400 ;
        RECT 55.950 271.950 58.050 274.050 ;
        RECT 56.400 262.050 57.450 271.950 ;
        RECT 68.400 265.050 69.450 280.950 ;
        RECT 79.950 280.500 82.050 282.600 ;
        RECT 82.950 274.950 85.050 277.050 ;
        RECT 67.950 262.950 70.050 265.050 ;
        RECT 55.950 259.950 58.050 262.050 ;
        RECT 61.950 259.950 67.050 262.050 ;
        RECT 79.950 259.950 82.050 262.050 ;
        RECT 52.950 253.950 58.050 256.050 ;
        RECT 67.950 253.950 70.050 256.050 ;
        RECT 49.950 247.950 52.050 250.050 ;
        RECT 68.400 223.050 69.450 253.950 ;
        RECT 80.400 250.050 81.450 259.950 ;
        RECT 83.400 256.050 84.450 274.950 ;
        RECT 82.950 253.950 85.050 256.050 ;
        RECT 79.950 247.950 82.050 250.050 ;
        RECT 67.950 220.950 70.050 223.050 ;
        RECT 73.950 220.950 76.050 223.050 ;
        RECT 49.950 217.950 55.050 220.050 ;
        RECT 58.950 217.950 61.050 220.050 ;
        RECT 40.950 214.950 43.050 217.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 1.950 208.950 4.050 211.050 ;
        RECT 10.950 208.950 13.050 211.050 ;
        RECT 13.950 208.950 19.050 211.050 ;
        RECT 22.950 208.950 28.050 211.050 ;
        RECT 46.950 208.950 49.050 211.050 ;
        RECT 2.400 61.050 3.450 208.950 ;
        RECT 34.950 190.950 37.050 193.050 ;
        RECT 19.950 188.400 22.050 190.500 ;
        RECT 10.950 181.950 19.050 184.050 ;
        RECT 7.950 175.950 10.050 178.050 ;
        RECT 8.400 154.050 9.450 175.950 ;
        RECT 7.950 151.950 10.050 154.050 ;
        RECT 7.950 146.400 10.050 148.500 ;
        RECT 8.700 126.600 9.900 146.400 ;
        RECT 7.950 124.500 10.050 126.600 ;
        RECT 14.400 120.450 15.450 181.950 ;
        RECT 20.850 173.400 22.050 188.400 ;
        RECT 35.400 181.050 36.450 190.950 ;
        RECT 40.950 188.400 43.050 190.500 ;
        RECT 28.950 178.950 31.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 19.950 171.300 22.050 173.400 ;
        RECT 20.850 167.700 22.050 171.300 ;
        RECT 19.950 165.600 22.050 167.700 ;
        RECT 29.400 157.050 30.450 178.950 ;
        RECT 41.100 168.600 42.300 188.400 ;
        RECT 43.950 181.950 46.050 184.050 ;
        RECT 44.400 178.050 45.450 181.950 ;
        RECT 43.950 175.950 46.050 178.050 ;
        RECT 40.950 166.500 43.050 168.600 ;
        RECT 19.950 154.950 22.050 157.050 ;
        RECT 28.950 154.950 31.050 157.050 ;
        RECT 16.950 133.950 19.050 139.050 ;
        RECT 20.400 136.050 21.450 154.950 ;
        RECT 37.950 151.950 40.050 154.050 ;
        RECT 28.950 147.300 31.050 149.400 ;
        RECT 28.950 143.700 30.150 147.300 ;
        RECT 28.950 141.600 31.050 143.700 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 16.950 121.950 19.050 124.050 ;
        RECT 11.400 119.400 15.450 120.450 ;
        RECT 11.400 103.050 12.450 119.400 ;
        RECT 13.950 112.950 16.050 115.050 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 7.950 68.400 10.050 70.500 ;
        RECT 4.950 64.950 7.050 67.050 ;
        RECT 1.950 58.950 4.050 61.050 ;
        RECT 5.400 55.050 6.450 64.950 ;
        RECT 4.950 52.950 7.050 55.050 ;
        RECT 8.700 48.600 9.900 68.400 ;
        RECT 14.400 67.050 15.450 112.950 ;
        RECT 17.400 103.050 18.450 121.950 ;
        RECT 16.950 100.950 19.050 103.050 ;
        RECT 13.950 64.950 16.050 67.050 ;
        RECT 13.950 58.950 19.050 61.050 ;
        RECT 20.400 58.050 21.450 133.950 ;
        RECT 28.950 126.600 30.150 141.600 ;
        RECT 38.400 136.050 39.450 151.950 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 31.950 132.450 36.000 133.050 ;
        RECT 31.950 130.950 36.450 132.450 ;
        RECT 28.950 124.500 31.050 126.600 ;
        RECT 35.400 124.050 36.450 130.950 ;
        RECT 37.950 127.950 40.050 130.050 ;
        RECT 34.950 121.950 37.050 124.050 ;
        RECT 38.400 112.200 39.450 127.950 ;
        RECT 47.400 118.050 48.450 208.950 ;
        RECT 49.950 205.950 52.050 208.050 ;
        RECT 50.400 151.050 51.450 205.950 ;
        RECT 53.400 175.050 54.450 211.950 ;
        RECT 55.950 181.950 58.050 187.050 ;
        RECT 59.400 181.050 60.450 217.950 ;
        RECT 74.400 217.050 75.450 220.950 ;
        RECT 83.400 217.200 84.450 253.950 ;
        RECT 89.400 223.050 90.450 319.950 ;
        RECT 98.400 307.050 99.450 352.950 ;
        RECT 100.950 349.950 103.050 352.050 ;
        RECT 101.400 310.050 102.450 349.950 ;
        RECT 113.400 343.050 114.450 373.800 ;
        RECT 119.400 367.050 120.450 376.950 ;
        RECT 118.950 364.950 121.050 367.050 ;
        RECT 103.950 340.950 106.050 343.050 ;
        RECT 112.950 340.950 115.050 343.050 ;
        RECT 100.950 307.950 103.050 310.050 ;
        RECT 97.950 304.950 100.050 307.050 ;
        RECT 104.400 295.050 105.450 340.950 ;
        RECT 109.950 334.950 115.050 337.050 ;
        RECT 115.950 334.950 121.050 337.050 ;
        RECT 122.400 334.050 123.450 388.950 ;
        RECT 130.950 373.950 136.050 376.050 ;
        RECT 140.400 373.050 141.450 391.950 ;
        RECT 146.400 388.050 147.450 415.950 ;
        RECT 149.400 415.050 150.450 439.950 ;
        RECT 152.400 418.050 153.450 442.950 ;
        RECT 169.950 439.950 172.050 445.050 ;
        RECT 176.400 436.050 177.450 448.950 ;
        RECT 179.400 445.200 180.450 478.950 ;
        RECT 188.400 478.050 189.450 526.950 ;
        RECT 194.400 523.050 195.450 547.950 ;
        RECT 196.950 544.950 199.050 547.050 ;
        RECT 197.400 538.200 198.450 544.950 ;
        RECT 196.950 536.100 199.050 538.200 ;
        RECT 196.950 532.800 199.050 534.900 ;
        RECT 192.000 522.900 195.450 523.050 ;
        RECT 190.950 521.250 195.450 522.900 ;
        RECT 190.950 520.950 195.000 521.250 ;
        RECT 190.950 520.800 193.050 520.950 ;
        RECT 197.400 496.050 198.450 532.800 ;
        RECT 200.400 532.050 201.450 559.950 ;
        RECT 206.400 550.050 207.450 571.950 ;
        RECT 209.400 568.050 210.450 580.950 ;
        RECT 212.400 571.050 213.450 613.950 ;
        RECT 214.950 612.900 219.000 613.050 ;
        RECT 214.950 610.950 220.050 612.900 ;
        RECT 217.950 610.800 220.050 610.950 ;
        RECT 224.400 610.050 225.450 613.950 ;
        RECT 226.950 610.950 229.050 613.050 ;
        RECT 233.400 612.450 234.450 625.950 ;
        RECT 245.400 616.050 246.450 640.950 ;
        RECT 253.950 622.950 256.050 625.050 ;
        RECT 244.950 613.950 247.050 616.050 ;
        RECT 233.400 611.400 237.450 612.450 ;
        RECT 223.950 607.950 226.050 610.050 ;
        RECT 220.950 607.050 223.050 607.200 ;
        RECT 217.950 605.100 223.050 607.050 ;
        RECT 217.950 604.950 222.000 605.100 ;
        RECT 219.000 603.900 222.000 604.050 ;
        RECT 219.000 603.300 223.050 603.900 ;
        RECT 218.400 601.950 223.050 603.300 ;
        RECT 218.400 595.050 219.450 601.950 ;
        RECT 220.950 601.800 223.050 601.950 ;
        RECT 220.950 595.950 223.050 598.050 ;
        RECT 217.950 592.950 220.050 595.050 ;
        RECT 221.400 592.050 222.450 595.950 ;
        RECT 220.950 589.950 223.050 592.050 ;
        RECT 227.400 577.050 228.450 610.950 ;
        RECT 232.950 604.950 235.050 610.050 ;
        RECT 226.950 574.950 229.050 577.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 220.950 568.950 223.050 571.050 ;
        RECT 208.950 565.950 211.050 568.050 ;
        RECT 214.950 565.950 220.050 568.050 ;
        RECT 205.950 547.950 208.050 550.050 ;
        RECT 199.950 529.950 202.050 532.050 ;
        RECT 200.400 511.050 201.450 529.950 ;
        RECT 218.400 529.050 219.450 565.950 ;
        RECT 221.400 538.050 222.450 568.950 ;
        RECT 223.950 565.950 226.050 571.050 ;
        RECT 236.400 568.050 237.450 611.400 ;
        RECT 247.950 610.950 250.050 613.050 ;
        RECT 238.950 607.950 241.050 610.050 ;
        RECT 235.950 565.950 238.050 568.050 ;
        RECT 226.950 559.950 229.050 565.050 ;
        RECT 235.950 559.950 238.050 562.050 ;
        RECT 236.400 556.050 237.450 559.950 ;
        RECT 235.950 553.950 238.050 556.050 ;
        RECT 220.950 535.950 223.050 538.050 ;
        RECT 235.950 535.950 238.050 538.050 ;
        RECT 218.400 527.400 223.050 529.050 ;
        RECT 219.000 526.950 223.050 527.400 ;
        RECT 226.950 526.950 232.050 529.050 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 202.950 523.950 205.050 526.050 ;
        RECT 203.400 520.050 204.450 523.950 ;
        RECT 217.950 520.950 220.050 523.050 ;
        RECT 223.950 520.950 226.050 523.050 ;
        RECT 229.950 520.950 232.050 523.050 ;
        RECT 202.950 517.950 205.050 520.050 ;
        RECT 199.950 508.950 202.050 511.050 ;
        RECT 208.950 508.950 211.050 511.050 ;
        RECT 199.950 502.950 202.050 505.050 ;
        RECT 196.950 493.950 199.050 496.050 ;
        RECT 197.400 490.050 198.450 493.950 ;
        RECT 200.400 493.050 201.450 502.950 ;
        RECT 205.950 496.950 208.050 499.050 ;
        RECT 199.950 490.950 205.050 493.050 ;
        RECT 206.400 490.050 207.450 496.950 ;
        RECT 196.950 487.950 199.050 490.050 ;
        RECT 205.950 489.450 208.050 490.050 ;
        RECT 203.400 488.400 208.050 489.450 ;
        RECT 190.950 484.950 193.050 487.050 ;
        RECT 187.950 475.950 190.050 478.050 ;
        RECT 191.400 466.050 192.450 484.950 ;
        RECT 203.400 466.050 204.450 488.400 ;
        RECT 205.950 487.950 208.050 488.400 ;
        RECT 209.400 484.050 210.450 508.950 ;
        RECT 218.400 493.050 219.450 520.950 ;
        RECT 224.400 502.050 225.450 520.950 ;
        RECT 223.950 499.950 226.050 502.050 ;
        RECT 230.400 499.050 231.450 520.950 ;
        RECT 233.400 517.050 234.450 526.950 ;
        RECT 232.950 514.950 235.050 517.050 ;
        RECT 236.400 508.050 237.450 535.950 ;
        RECT 239.400 529.050 240.450 607.950 ;
        RECT 248.400 601.050 249.450 610.950 ;
        RECT 254.400 610.050 255.450 622.950 ;
        RECT 257.400 612.450 258.450 649.950 ;
        RECT 260.400 615.450 261.450 673.950 ;
        RECT 263.400 670.050 264.450 676.950 ;
        RECT 268.950 673.950 271.050 679.050 ;
        RECT 274.950 676.950 280.050 679.050 ;
        RECT 280.950 673.950 283.050 676.050 ;
        RECT 262.950 667.950 265.050 670.050 ;
        RECT 281.400 664.050 282.450 673.950 ;
        RECT 280.950 661.950 283.050 664.050 ;
        RECT 290.400 655.050 291.450 716.400 ;
        RECT 296.400 694.050 297.450 719.400 ;
        RECT 316.950 718.950 319.050 721.050 ;
        RECT 298.950 715.950 304.050 718.050 ;
        RECT 313.950 697.950 316.050 700.050 ;
        RECT 304.950 694.950 307.050 697.050 ;
        RECT 295.950 691.950 298.050 694.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 293.400 676.050 294.450 679.950 ;
        RECT 296.400 679.050 297.450 691.950 ;
        RECT 301.950 688.950 304.050 694.050 ;
        RECT 305.400 685.050 306.450 694.950 ;
        RECT 310.950 685.950 313.050 688.050 ;
        RECT 304.950 682.950 307.050 685.050 ;
        RECT 306.000 681.450 310.050 682.050 ;
        RECT 305.400 679.950 310.050 681.450 ;
        RECT 295.950 676.950 298.050 679.050 ;
        RECT 292.950 673.950 295.050 676.050 ;
        RECT 295.950 655.950 298.050 658.050 ;
        RECT 289.950 652.950 292.050 655.050 ;
        RECT 286.950 649.950 289.050 652.050 ;
        RECT 292.950 649.950 295.050 652.050 ;
        RECT 277.950 644.100 280.050 649.050 ;
        RECT 280.950 643.950 286.050 646.050 ;
        RECT 277.950 640.800 280.050 642.900 ;
        RECT 268.950 628.950 271.050 631.050 ;
        RECT 260.400 614.400 264.450 615.450 ;
        RECT 257.400 611.400 261.450 612.450 ;
        RECT 260.400 610.050 261.450 611.400 ;
        RECT 254.400 608.400 259.050 610.050 ;
        RECT 255.000 607.950 259.050 608.400 ;
        RECT 259.950 607.950 262.050 610.050 ;
        RECT 250.950 604.950 253.050 607.050 ;
        RECT 241.950 598.950 244.050 601.050 ;
        RECT 247.950 598.950 250.050 601.050 ;
        RECT 242.400 595.050 243.450 598.950 ;
        RECT 241.950 592.950 244.050 595.050 ;
        RECT 251.400 574.050 252.450 604.950 ;
        RECT 253.950 601.950 259.050 604.050 ;
        RECT 260.400 601.050 261.450 607.950 ;
        RECT 259.950 598.950 262.050 601.050 ;
        RECT 263.400 577.050 264.450 614.400 ;
        RECT 269.400 610.200 270.450 628.950 ;
        RECT 278.400 619.050 279.450 640.800 ;
        RECT 287.400 640.050 288.450 649.950 ;
        RECT 289.950 643.950 292.050 646.050 ;
        RECT 286.950 637.950 289.050 640.050 ;
        RECT 277.950 616.950 280.050 619.050 ;
        RECT 283.950 616.950 286.050 619.050 ;
        RECT 268.950 608.100 271.050 610.200 ;
        RECT 268.950 604.800 271.050 606.900 ;
        RECT 262.950 574.950 265.050 577.050 ;
        RECT 250.950 571.950 253.050 574.050 ;
        RECT 256.950 573.450 261.000 574.050 ;
        RECT 256.950 571.950 261.450 573.450 ;
        RECT 265.950 571.950 268.050 574.050 ;
        RECT 247.950 565.950 250.050 568.050 ;
        RECT 253.950 565.950 256.050 568.050 ;
        RECT 248.400 559.050 249.450 565.950 ;
        RECT 247.950 556.950 250.050 559.050 ;
        RECT 254.400 553.050 255.450 565.950 ;
        RECT 253.950 550.950 256.050 553.050 ;
        RECT 254.400 529.050 255.450 550.950 ;
        RECT 260.400 541.050 261.450 571.950 ;
        RECT 262.950 562.800 265.050 564.900 ;
        RECT 259.950 538.950 262.050 541.050 ;
        RECT 238.950 526.950 241.050 529.050 ;
        RECT 253.950 526.950 256.050 529.050 ;
        RECT 259.950 526.950 262.050 532.050 ;
        RECT 250.950 520.950 253.050 523.050 ;
        RECT 256.950 520.950 259.050 523.050 ;
        RECT 235.950 505.950 238.050 508.050 ;
        RECT 232.950 502.950 235.050 505.050 ;
        RECT 229.950 496.950 232.050 499.050 ;
        RECT 233.400 496.050 234.450 502.950 ;
        RECT 217.950 490.950 220.050 493.050 ;
        RECT 226.950 490.950 229.050 493.050 ;
        RECT 232.950 490.950 235.050 496.050 ;
        RECT 238.950 493.950 241.050 496.050 ;
        RECT 208.950 481.950 211.050 484.050 ;
        RECT 217.950 483.450 220.050 487.050 ;
        RECT 215.400 482.400 220.050 483.450 ;
        RECT 209.400 478.050 210.450 481.950 ;
        RECT 205.800 475.950 207.900 478.050 ;
        RECT 209.100 477.450 211.200 478.050 ;
        RECT 209.100 476.400 213.450 477.450 ;
        RECT 209.100 475.950 211.200 476.400 ;
        RECT 190.950 463.950 193.050 466.050 ;
        RECT 202.950 463.950 205.050 466.050 ;
        RECT 193.950 457.950 196.050 460.050 ;
        RECT 194.400 454.050 195.450 457.950 ;
        RECT 181.950 451.950 184.050 454.050 ;
        RECT 184.950 451.950 187.050 454.050 ;
        RECT 193.950 451.950 196.050 454.050 ;
        RECT 182.400 448.050 183.450 451.950 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 178.950 443.100 181.050 445.200 ;
        RECT 178.950 439.800 181.050 441.900 ;
        RECT 166.950 433.950 169.050 436.050 ;
        RECT 175.950 433.950 178.050 436.050 ;
        RECT 154.950 421.950 157.050 424.050 ;
        RECT 151.950 415.950 154.050 418.050 ;
        RECT 148.950 409.950 151.050 415.050 ;
        RECT 155.400 412.050 156.450 421.950 ;
        RECT 157.950 415.950 160.050 421.050 ;
        RECT 167.400 415.050 168.450 433.950 ;
        RECT 179.400 424.050 180.450 439.800 ;
        RECT 178.950 421.950 181.050 424.050 ;
        RECT 169.950 418.950 172.050 421.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 154.950 409.950 157.050 412.050 ;
        RECT 145.950 385.950 148.050 388.050 ;
        RECT 160.950 379.950 163.050 382.050 ;
        RECT 142.950 376.950 145.050 379.050 ;
        RECT 127.950 367.950 130.050 373.050 ;
        RECT 139.950 370.950 142.050 373.050 ;
        RECT 143.400 370.050 144.450 376.950 ;
        RECT 133.950 367.950 139.050 370.050 ;
        RECT 142.950 367.950 145.050 370.050 ;
        RECT 151.950 367.950 154.050 370.050 ;
        RECT 152.400 352.050 153.450 367.950 ;
        RECT 161.400 367.050 162.450 379.950 ;
        RECT 170.400 379.050 171.450 418.950 ;
        RECT 172.950 409.950 175.050 415.050 ;
        RECT 178.950 412.950 184.050 415.050 ;
        RECT 185.400 411.450 186.450 451.950 ;
        RECT 187.950 448.950 190.050 451.050 ;
        RECT 179.400 411.000 186.450 411.450 ;
        RECT 178.950 410.400 186.450 411.000 ;
        RECT 178.950 406.950 181.050 410.400 ;
        RECT 188.400 409.050 189.450 448.950 ;
        RECT 190.950 445.950 193.050 448.050 ;
        RECT 191.400 442.050 192.450 445.950 ;
        RECT 202.950 444.450 205.050 448.050 ;
        RECT 200.400 444.000 205.050 444.450 ;
        RECT 200.400 443.400 204.450 444.000 ;
        RECT 190.950 439.950 193.050 442.050 ;
        RECT 200.400 436.050 201.450 443.400 ;
        RECT 206.400 441.450 207.450 475.950 ;
        RECT 212.400 454.050 213.450 476.400 ;
        RECT 215.400 460.050 216.450 482.400 ;
        RECT 217.950 482.100 220.050 482.400 ;
        RECT 227.400 481.050 228.450 490.950 ;
        RECT 239.400 490.050 240.450 493.950 ;
        RECT 244.950 490.950 247.050 493.050 ;
        RECT 238.950 487.950 241.050 490.050 ;
        RECT 217.950 478.800 220.050 480.900 ;
        RECT 226.950 478.950 229.050 481.050 ;
        RECT 218.400 472.050 219.450 478.800 ;
        RECT 229.950 475.950 232.050 478.050 ;
        RECT 217.950 469.950 220.050 472.050 ;
        RECT 217.950 463.950 220.050 466.050 ;
        RECT 214.950 457.950 217.050 460.050 ;
        RECT 218.400 457.050 219.450 463.950 ;
        RECT 220.950 460.950 223.050 463.050 ;
        RECT 211.950 451.950 214.050 454.050 ;
        RECT 217.950 451.950 220.050 457.050 ;
        RECT 211.950 442.950 214.050 445.050 ;
        RECT 203.400 440.400 207.450 441.450 ;
        RECT 199.950 433.950 202.050 436.050 ;
        RECT 190.950 415.950 193.050 418.050 ;
        RECT 184.950 407.400 189.450 409.050 ;
        RECT 184.950 406.950 189.000 407.400 ;
        RECT 179.400 379.050 180.450 406.950 ;
        RECT 191.400 394.050 192.450 415.950 ;
        RECT 200.400 412.050 201.450 433.950 ;
        RECT 203.400 412.050 204.450 440.400 ;
        RECT 205.950 436.950 208.050 439.050 ;
        RECT 206.400 415.200 207.450 436.950 ;
        RECT 212.400 436.050 213.450 442.950 ;
        RECT 211.950 433.950 214.050 436.050 ;
        RECT 218.400 432.450 219.450 451.950 ;
        RECT 221.400 448.050 222.450 460.950 ;
        RECT 220.950 445.950 223.050 448.050 ;
        RECT 230.400 445.050 231.450 475.950 ;
        RECT 239.400 463.050 240.450 487.950 ;
        RECT 245.400 486.450 246.450 490.950 ;
        RECT 251.400 490.050 252.450 520.950 ;
        RECT 257.400 517.050 258.450 520.950 ;
        RECT 259.950 517.950 262.050 520.050 ;
        RECT 256.950 514.950 259.050 517.050 ;
        RECT 260.400 496.050 261.450 517.950 ;
        RECT 253.950 490.950 256.050 496.050 ;
        RECT 259.950 493.950 262.050 496.050 ;
        RECT 250.950 487.950 253.050 490.050 ;
        RECT 254.400 487.050 255.450 490.950 ;
        RECT 256.950 487.950 259.050 490.050 ;
        RECT 245.400 485.400 249.450 486.450 ;
        RECT 244.950 478.950 247.050 481.050 ;
        RECT 232.950 460.950 235.050 463.050 ;
        RECT 238.950 460.950 241.050 463.050 ;
        RECT 233.400 451.050 234.450 460.950 ;
        RECT 238.950 454.950 241.050 457.050 ;
        RECT 239.400 451.050 240.450 454.950 ;
        RECT 232.950 448.950 235.050 451.050 ;
        RECT 238.950 448.950 241.050 451.050 ;
        RECT 229.950 442.950 232.050 445.050 ;
        RECT 235.950 442.950 238.050 448.050 ;
        RECT 241.950 442.950 244.050 445.050 ;
        RECT 242.400 436.050 243.450 442.950 ;
        RECT 241.950 433.950 244.050 436.050 ;
        RECT 215.400 431.400 219.450 432.450 ;
        RECT 208.950 415.950 211.050 421.050 ;
        RECT 205.950 413.100 208.050 415.200 ;
        RECT 199.950 409.950 202.050 412.050 ;
        RECT 203.400 411.900 207.000 412.050 ;
        RECT 203.400 410.250 208.050 411.900 ;
        RECT 204.000 409.950 208.050 410.250 ;
        RECT 211.950 409.950 214.050 412.050 ;
        RECT 205.950 409.800 208.050 409.950 ;
        RECT 190.950 391.950 193.050 394.050 ;
        RECT 199.950 391.950 202.050 394.050 ;
        RECT 169.950 376.950 172.050 379.050 ;
        RECT 179.400 377.400 184.050 379.050 ;
        RECT 180.000 376.950 184.050 377.400 ;
        RECT 166.950 373.950 169.050 376.050 ;
        RECT 160.950 364.950 163.050 367.050 ;
        RECT 151.950 349.950 154.050 352.050 ;
        RECT 130.950 337.950 133.050 340.050 ;
        RECT 145.950 337.950 151.050 340.050 ;
        RECT 154.950 337.950 160.050 340.050 ;
        RECT 121.950 331.950 124.050 334.050 ;
        RECT 115.950 328.950 118.050 331.050 ;
        RECT 116.400 295.050 117.450 328.950 ;
        RECT 124.950 325.950 127.050 328.050 ;
        RECT 125.400 295.050 126.450 325.950 ;
        RECT 131.400 295.050 132.450 337.950 ;
        RECT 133.950 334.950 136.050 337.050 ;
        RECT 134.400 328.050 135.450 334.950 ;
        RECT 136.950 328.950 139.050 334.050 ;
        RECT 142.950 328.950 148.050 331.050 ;
        RECT 151.950 328.950 154.050 337.050 ;
        RECT 157.950 328.950 160.050 334.050 ;
        RECT 133.950 325.950 136.050 328.050 ;
        RECT 161.400 322.050 162.450 364.950 ;
        RECT 163.950 337.950 166.050 340.050 ;
        RECT 160.950 319.950 163.050 322.050 ;
        RECT 164.400 318.450 165.450 337.950 ;
        RECT 167.400 334.050 168.450 373.950 ;
        RECT 178.950 370.950 181.050 376.050 ;
        RECT 200.400 373.050 201.450 391.950 ;
        RECT 202.950 388.950 205.050 391.050 ;
        RECT 203.400 385.050 204.450 388.950 ;
        RECT 202.950 382.950 205.050 385.050 ;
        RECT 174.000 369.450 178.050 370.050 ;
        RECT 173.400 367.950 178.050 369.450 ;
        RECT 193.950 367.950 196.050 373.050 ;
        RECT 199.950 370.950 202.050 373.050 ;
        RECT 173.400 340.050 174.450 367.950 ;
        RECT 203.400 367.050 204.450 382.950 ;
        RECT 212.400 375.450 213.450 409.950 ;
        RECT 215.400 376.050 216.450 431.400 ;
        RECT 217.950 427.950 220.050 430.050 ;
        RECT 218.400 415.050 219.450 427.950 ;
        RECT 223.950 421.950 226.050 424.050 ;
        RECT 232.950 421.950 235.050 424.050 ;
        RECT 220.950 418.950 223.050 421.050 ;
        RECT 221.400 415.050 222.450 418.950 ;
        RECT 224.400 415.050 225.450 421.950 ;
        RECT 233.400 418.050 234.450 421.950 ;
        RECT 245.400 421.200 246.450 478.950 ;
        RECT 248.400 445.050 249.450 485.400 ;
        RECT 253.950 484.950 256.050 487.050 ;
        RECT 257.400 481.050 258.450 487.950 ;
        RECT 256.950 478.950 259.050 481.050 ;
        RECT 250.950 448.950 253.050 451.050 ;
        RECT 247.950 442.950 250.050 445.050 ;
        RECT 244.950 419.100 247.050 421.200 ;
        RECT 247.950 418.050 250.050 418.200 ;
        RECT 251.400 418.050 252.450 448.950 ;
        RECT 260.400 445.050 261.450 493.950 ;
        RECT 263.400 448.050 264.450 562.800 ;
        RECT 266.400 553.050 267.450 571.950 ;
        RECT 265.950 550.950 268.050 553.050 ;
        RECT 265.950 544.950 268.050 547.050 ;
        RECT 266.400 523.050 267.450 544.950 ;
        RECT 269.400 535.050 270.450 604.800 ;
        RECT 271.950 598.950 274.050 604.050 ;
        RECT 277.950 598.950 280.050 604.050 ;
        RECT 271.950 589.950 274.050 592.050 ;
        RECT 272.400 580.050 273.450 589.950 ;
        RECT 277.950 586.950 280.050 589.050 ;
        RECT 278.400 583.050 279.450 586.950 ;
        RECT 284.400 586.050 285.450 616.950 ;
        RECT 290.400 610.200 291.450 643.950 ;
        RECT 293.400 637.050 294.450 649.950 ;
        RECT 292.950 634.950 295.050 637.050 ;
        RECT 296.400 612.450 297.450 655.950 ;
        RECT 301.950 649.950 304.050 655.050 ;
        RECT 305.400 646.050 306.450 679.950 ;
        RECT 307.950 661.950 310.050 664.050 ;
        RECT 304.950 643.950 307.050 646.050 ;
        RECT 308.400 639.450 309.450 661.950 ;
        RECT 311.400 643.050 312.450 685.950 ;
        RECT 314.400 649.050 315.450 697.950 ;
        RECT 317.400 658.050 318.450 718.950 ;
        RECT 323.400 715.050 324.450 766.950 ;
        RECT 325.950 763.950 328.050 766.050 ;
        RECT 326.400 736.050 327.450 763.950 ;
        RECT 334.950 761.100 337.050 766.050 ;
        RECT 331.950 759.900 336.000 760.050 ;
        RECT 331.950 757.950 337.050 759.900 ;
        RECT 334.950 757.800 337.050 757.950 ;
        RECT 337.950 754.950 340.050 757.050 ;
        RECT 338.400 745.050 339.450 754.950 ;
        RECT 341.400 748.050 342.450 766.950 ;
        RECT 343.950 763.950 346.050 766.050 ;
        RECT 344.400 760.050 345.450 763.950 ;
        RECT 350.400 760.050 351.450 790.950 ;
        RECT 353.400 769.050 354.450 799.950 ;
        RECT 364.950 799.800 367.050 799.950 ;
        RECT 358.950 793.950 361.050 799.050 ;
        RECT 370.800 796.950 372.900 799.050 ;
        RECT 373.950 796.950 376.050 802.050 ;
        RECT 367.950 790.950 370.050 793.050 ;
        RECT 352.950 766.950 355.050 769.050 ;
        RECT 358.950 766.950 364.050 769.050 ;
        RECT 368.400 763.050 369.450 790.950 ;
        RECT 371.400 766.050 372.450 796.950 ;
        RECT 380.400 793.050 381.450 805.950 ;
        RECT 386.400 805.050 387.450 814.950 ;
        RECT 397.950 805.950 400.050 808.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 388.950 799.950 391.050 805.050 ;
        RECT 379.950 790.950 382.050 793.050 ;
        RECT 389.400 778.050 390.450 799.950 ;
        RECT 391.950 793.950 394.050 799.050 ;
        RECT 398.400 790.050 399.450 805.950 ;
        RECT 409.950 802.950 412.050 808.050 ;
        RECT 416.400 802.050 417.450 814.950 ;
        RECT 427.950 808.950 430.050 811.050 ;
        RECT 418.950 805.950 421.050 808.050 ;
        RECT 406.950 799.950 409.050 802.050 ;
        RECT 412.950 800.400 417.450 802.050 ;
        RECT 412.950 799.950 417.000 800.400 ;
        RECT 407.400 796.050 408.450 799.950 ;
        RECT 419.400 799.050 420.450 805.950 ;
        RECT 428.400 805.050 429.450 808.950 ;
        RECT 434.400 808.050 435.450 817.950 ;
        RECT 433.950 805.950 436.050 808.050 ;
        RECT 427.950 802.950 430.050 805.050 ;
        RECT 448.950 802.950 451.050 808.050 ;
        RECT 454.950 805.950 457.050 808.050 ;
        RECT 463.950 805.950 466.050 811.050 ;
        RECT 473.400 808.050 474.450 817.950 ;
        RECT 517.950 814.950 520.050 817.050 ;
        RECT 719.400 816.000 726.450 816.450 ;
        RECT 718.950 815.400 726.450 816.000 ;
        RECT 472.950 805.950 475.050 808.050 ;
        RECT 429.000 801.450 433.050 802.050 ;
        RECT 428.400 799.950 433.050 801.450 ;
        RECT 445.950 799.950 448.050 802.050 ;
        RECT 418.950 796.950 421.050 799.050 ;
        RECT 406.950 793.950 409.050 796.050 ;
        RECT 424.950 793.950 427.050 796.050 ;
        RECT 425.400 790.050 426.450 793.950 ;
        RECT 428.400 793.050 429.450 799.950 ;
        RECT 433.950 793.950 436.050 799.050 ;
        RECT 446.400 793.050 447.450 799.950 ;
        RECT 449.400 796.050 450.450 802.950 ;
        RECT 455.400 802.050 456.450 805.950 ;
        RECT 478.950 802.950 481.050 808.050 ;
        RECT 484.950 805.950 487.050 811.050 ;
        RECT 502.950 805.950 505.050 811.050 ;
        RECT 511.950 805.950 514.050 811.050 ;
        RECT 518.400 808.050 519.450 814.950 ;
        RECT 718.950 814.050 721.050 815.400 ;
        RECT 535.950 811.950 538.050 814.050 ;
        RECT 550.950 811.950 553.050 814.050 ;
        RECT 586.950 811.950 589.050 814.050 ;
        RECT 703.950 811.950 706.050 814.050 ;
        RECT 718.800 813.000 721.050 814.050 ;
        RECT 722.100 813.000 724.200 814.050 ;
        RECT 718.800 811.950 720.900 813.000 ;
        RECT 721.950 811.950 724.200 813.000 ;
        RECT 517.950 805.950 520.050 808.050 ;
        RECT 536.400 802.050 537.450 811.950 ;
        RECT 551.400 808.050 552.450 811.950 ;
        RECT 551.400 806.400 556.050 808.050 ;
        RECT 552.000 805.950 556.050 806.400 ;
        RECT 565.950 805.950 568.050 808.050 ;
        RECT 570.000 807.450 574.050 808.050 ;
        RECT 569.400 805.950 574.050 807.450 ;
        RECT 538.950 802.950 541.050 805.050 ;
        RECT 541.950 802.950 544.050 805.050 ;
        RECT 451.950 800.400 456.450 802.050 ;
        RECT 451.950 799.950 456.000 800.400 ;
        RECT 460.950 799.950 463.050 802.050 ;
        RECT 466.950 799.950 472.050 802.050 ;
        RECT 472.950 799.950 478.050 802.050 ;
        RECT 493.950 799.950 496.050 802.050 ;
        RECT 499.950 799.950 502.050 802.050 ;
        RECT 511.950 799.950 517.050 802.050 ;
        RECT 520.950 799.950 523.050 802.050 ;
        RECT 535.950 799.950 538.050 802.050 ;
        RECT 448.950 793.950 451.050 796.050 ;
        RECT 461.400 793.050 462.450 799.950 ;
        RECT 427.950 790.950 430.050 793.050 ;
        RECT 445.950 790.950 448.050 793.050 ;
        RECT 460.950 790.950 463.050 793.050 ;
        RECT 487.950 790.950 490.050 793.050 ;
        RECT 397.950 787.950 400.050 790.050 ;
        RECT 424.950 787.950 427.050 790.050 ;
        RECT 394.950 781.950 397.050 784.050 ;
        RECT 376.950 775.950 379.050 778.050 ;
        RECT 388.950 775.950 391.050 778.050 ;
        RECT 373.950 772.950 376.050 775.050 ;
        RECT 370.950 763.950 373.050 766.050 ;
        RECT 355.950 760.950 361.050 763.050 ;
        RECT 364.950 760.950 367.050 763.050 ;
        RECT 367.950 760.950 370.050 763.050 ;
        RECT 343.950 757.950 346.050 760.050 ;
        RECT 350.400 758.400 355.050 760.050 ;
        RECT 351.000 757.950 355.050 758.400 ;
        RECT 346.950 756.450 351.000 757.050 ;
        RECT 346.950 756.000 351.450 756.450 ;
        RECT 346.950 754.950 352.050 756.000 ;
        RECT 343.950 751.950 346.050 754.050 ;
        RECT 349.950 751.950 352.050 754.950 ;
        RECT 340.950 745.950 343.050 748.050 ;
        RECT 337.950 742.950 340.050 745.050 ;
        RECT 325.950 733.950 328.050 736.050 ;
        RECT 344.400 727.050 345.450 751.950 ;
        RECT 365.400 748.050 366.450 760.950 ;
        RECT 374.400 760.050 375.450 772.950 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 370.950 757.050 373.050 757.200 ;
        RECT 370.950 756.600 375.000 757.050 ;
        RECT 370.950 755.100 375.450 756.600 ;
        RECT 372.000 754.950 375.450 755.100 ;
        RECT 370.950 748.950 373.050 753.900 ;
        RECT 364.950 745.950 367.050 748.050 ;
        RECT 367.950 733.950 370.050 736.050 ;
        RECT 358.950 727.950 361.050 730.050 ;
        RECT 328.950 723.450 333.000 724.050 ;
        RECT 328.950 721.950 333.450 723.450 ;
        RECT 334.950 721.950 337.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 349.950 724.950 352.050 727.050 ;
        RECT 332.400 721.050 333.450 721.950 ;
        RECT 350.400 721.050 351.450 724.950 ;
        RECT 359.400 721.050 360.450 727.950 ;
        RECT 368.400 727.050 369.450 733.950 ;
        RECT 367.950 724.950 370.050 727.050 ;
        RECT 370.950 721.950 373.050 727.050 ;
        RECT 331.950 718.950 334.050 721.050 ;
        RECT 340.950 718.950 346.050 721.050 ;
        RECT 349.950 718.950 352.050 721.050 ;
        RECT 358.950 718.950 361.050 721.050 ;
        RECT 322.950 712.950 325.050 715.050 ;
        RECT 322.950 682.950 325.050 688.050 ;
        RECT 328.950 685.950 331.050 688.050 ;
        RECT 329.400 664.050 330.450 685.950 ;
        RECT 332.400 685.050 333.450 718.950 ;
        RECT 334.950 715.950 337.050 718.050 ;
        RECT 331.950 682.950 334.050 685.050 ;
        RECT 319.950 661.950 322.050 664.050 ;
        RECT 328.950 661.950 331.050 664.050 ;
        RECT 316.950 655.950 319.050 658.050 ;
        RECT 320.400 649.200 321.450 661.950 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 319.950 647.100 322.050 649.200 ;
        RECT 316.950 645.900 321.000 646.050 ;
        RECT 316.950 643.950 322.050 645.900 ;
        RECT 328.950 643.950 331.050 649.050 ;
        RECT 319.950 643.800 322.050 643.950 ;
        RECT 332.400 643.050 333.450 682.950 ;
        RECT 335.400 682.200 336.450 715.950 ;
        RECT 346.950 697.950 349.050 700.050 ;
        RECT 347.400 691.050 348.450 697.950 ;
        RECT 343.950 688.950 346.050 691.050 ;
        RECT 346.950 688.950 349.050 691.050 ;
        RECT 334.950 680.100 337.050 682.200 ;
        RECT 334.950 676.800 337.050 678.900 ;
        RECT 335.400 651.450 336.450 676.800 ;
        RECT 344.400 673.050 345.450 688.950 ;
        RECT 346.950 679.950 349.050 685.050 ;
        RECT 350.400 679.050 351.450 718.950 ;
        RECT 374.400 718.050 375.450 754.950 ;
        RECT 370.950 715.950 376.050 718.050 ;
        RECT 352.950 706.950 355.050 709.050 ;
        RECT 358.950 706.950 361.050 709.050 ;
        RECT 353.400 679.050 354.450 706.950 ;
        RECT 359.400 685.050 360.450 706.950 ;
        RECT 364.950 688.950 367.050 691.050 ;
        RECT 365.400 685.050 366.450 688.950 ;
        RECT 377.400 688.050 378.450 775.950 ;
        RECT 391.950 772.950 394.050 775.050 ;
        RECT 382.950 763.950 385.050 766.050 ;
        RECT 383.400 724.050 384.450 763.950 ;
        RECT 385.950 763.050 388.050 763.200 ;
        RECT 388.950 763.050 391.050 763.200 ;
        RECT 392.400 763.050 393.450 772.950 ;
        RECT 385.950 761.100 391.050 763.050 ;
        RECT 387.000 760.950 390.000 761.100 ;
        RECT 385.950 757.800 388.050 759.900 ;
        RECT 391.950 757.950 394.050 763.050 ;
        RECT 386.400 736.050 387.450 757.800 ;
        RECT 388.950 751.950 391.050 757.050 ;
        RECT 385.950 733.950 388.050 736.050 ;
        RECT 386.400 727.050 387.450 733.950 ;
        RECT 395.400 732.450 396.450 781.950 ;
        RECT 397.950 769.950 400.050 772.050 ;
        RECT 398.400 766.050 399.450 769.950 ;
        RECT 409.950 766.950 415.050 769.050 ;
        RECT 421.950 766.950 424.050 769.050 ;
        RECT 397.950 763.950 400.050 766.050 ;
        RECT 406.950 760.950 415.050 763.050 ;
        RECT 400.950 757.950 406.050 760.050 ;
        RECT 415.950 754.950 418.050 757.050 ;
        RECT 418.950 754.950 421.050 757.050 ;
        RECT 403.950 745.950 406.050 748.050 ;
        RECT 392.400 732.000 396.450 732.450 ;
        RECT 391.950 731.400 396.450 732.000 ;
        RECT 391.950 727.950 394.050 731.400 ;
        RECT 404.400 730.050 405.450 745.950 ;
        RECT 416.400 742.050 417.450 754.950 ;
        RECT 415.950 739.950 418.050 742.050 ;
        RECT 394.950 727.950 397.050 730.050 ;
        RECT 403.950 727.950 406.050 730.050 ;
        RECT 388.950 727.050 391.050 727.200 ;
        RECT 386.400 725.550 391.050 727.050 ;
        RECT 387.000 725.100 391.050 725.550 ;
        RECT 387.000 724.950 390.000 725.100 ;
        RECT 382.950 721.950 385.050 724.050 ;
        RECT 390.000 723.900 394.050 724.050 ;
        RECT 388.950 721.950 394.050 723.900 ;
        RECT 388.950 721.800 391.050 721.950 ;
        RECT 379.950 718.950 382.050 721.050 ;
        RECT 380.400 697.050 381.450 718.950 ;
        RECT 395.400 718.050 396.450 727.950 ;
        RECT 406.950 721.950 409.050 727.050 ;
        RECT 409.950 721.950 415.050 724.050 ;
        RECT 394.950 715.950 397.050 718.050 ;
        RECT 400.950 709.950 403.050 712.050 ;
        RECT 385.950 706.950 388.050 709.050 ;
        RECT 379.950 694.950 382.050 697.050 ;
        RECT 386.400 691.050 387.450 706.950 ;
        RECT 388.950 691.950 391.050 694.050 ;
        RECT 385.950 688.950 388.050 691.050 ;
        RECT 376.950 685.950 379.050 688.050 ;
        RECT 382.950 685.050 385.050 685.200 ;
        RECT 385.950 685.050 388.050 685.200 ;
        RECT 389.400 685.050 390.450 691.950 ;
        RECT 401.400 685.050 402.450 709.950 ;
        RECT 416.400 709.050 417.450 739.950 ;
        RECT 419.400 730.050 420.450 754.950 ;
        RECT 422.400 754.050 423.450 766.950 ;
        RECT 421.950 751.950 424.050 754.050 ;
        RECT 418.950 727.950 421.050 730.050 ;
        RECT 415.950 706.950 418.050 709.050 ;
        RECT 418.950 697.950 421.050 700.050 ;
        RECT 403.950 691.950 409.050 694.050 ;
        RECT 412.950 691.950 418.050 694.050 ;
        RECT 409.950 688.950 412.050 691.050 ;
        RECT 355.950 682.950 361.050 685.050 ;
        RECT 364.950 679.950 367.050 685.050 ;
        RECT 370.950 682.950 373.050 685.050 ;
        RECT 382.950 683.100 388.050 685.050 ;
        RECT 384.000 682.950 387.000 683.100 ;
        RECT 388.950 682.950 391.050 685.050 ;
        RECT 394.950 682.950 400.050 685.050 ;
        RECT 401.400 683.400 406.050 685.050 ;
        RECT 402.000 682.950 406.050 683.400 ;
        RECT 349.950 676.950 352.050 679.050 ;
        RECT 352.950 676.950 355.050 679.050 ;
        RECT 361.950 678.450 364.050 679.050 ;
        RECT 371.400 678.450 372.450 682.950 ;
        RECT 379.950 681.900 384.000 682.050 ;
        RECT 379.950 679.950 385.050 681.900 ;
        RECT 382.950 679.800 385.050 679.950 ;
        RECT 410.400 679.050 411.450 688.950 ;
        RECT 419.400 685.050 420.450 697.950 ;
        RECT 422.400 688.050 423.450 751.950 ;
        RECT 425.400 727.050 426.450 787.950 ;
        RECT 428.400 730.050 429.450 790.950 ;
        RECT 448.950 778.950 451.050 781.050 ;
        RECT 449.400 766.050 450.450 778.950 ;
        RECT 484.950 775.950 487.050 778.050 ;
        RECT 475.950 772.950 478.050 775.050 ;
        RECT 463.950 769.950 466.050 772.050 ;
        RECT 433.950 760.950 439.050 763.050 ;
        RECT 442.950 760.950 445.050 766.050 ;
        RECT 448.950 763.950 451.050 766.050 ;
        RECT 433.950 754.050 436.050 757.050 ;
        RECT 439.950 754.950 442.050 760.050 ;
        RECT 449.400 757.050 450.450 763.950 ;
        RECT 457.950 761.100 460.050 766.050 ;
        RECT 464.400 760.050 465.450 769.950 ;
        RECT 466.950 763.950 469.050 766.050 ;
        RECT 457.950 757.800 460.050 759.900 ;
        RECT 463.950 757.950 466.050 760.050 ;
        RECT 467.400 759.450 468.450 763.950 ;
        RECT 476.400 763.050 477.450 772.950 ;
        RECT 485.400 766.050 486.450 775.950 ;
        RECT 484.950 763.950 487.050 766.050 ;
        RECT 469.950 762.450 474.000 763.050 ;
        RECT 469.950 760.950 474.450 762.450 ;
        RECT 475.950 760.950 478.050 763.050 ;
        RECT 488.400 762.450 489.450 790.950 ;
        RECT 490.950 781.950 493.050 784.050 ;
        RECT 485.400 761.400 489.450 762.450 ;
        RECT 467.400 758.400 471.450 759.450 ;
        RECT 445.950 755.400 450.450 757.050 ;
        RECT 445.950 754.950 450.000 755.400 ;
        RECT 458.400 754.050 459.450 757.800 ;
        RECT 466.950 754.950 469.050 757.050 ;
        RECT 433.800 753.000 436.050 754.050 ;
        RECT 433.800 751.950 435.900 753.000 ;
        RECT 437.100 751.950 439.200 754.050 ;
        RECT 451.950 751.950 454.050 754.050 ;
        RECT 457.950 751.950 460.050 754.050 ;
        RECT 437.400 742.050 438.450 751.950 ;
        RECT 436.950 739.950 439.050 742.050 ;
        RECT 452.400 741.450 453.450 751.950 ;
        RECT 467.400 742.050 468.450 754.950 ;
        RECT 457.950 741.450 460.050 742.050 ;
        RECT 452.400 740.400 460.050 741.450 ;
        RECT 457.950 739.950 460.050 740.400 ;
        RECT 466.950 739.950 469.050 742.050 ;
        RECT 451.950 736.950 454.050 739.050 ;
        RECT 427.950 727.950 430.050 730.050 ;
        RECT 433.950 727.950 436.050 733.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 424.950 718.950 427.050 721.050 ;
        RECT 430.950 718.950 433.050 724.050 ;
        RECT 439.950 721.950 445.050 724.050 ;
        RECT 449.400 721.050 450.450 724.950 ;
        RECT 452.400 724.050 453.450 736.950 ;
        RECT 466.950 733.950 469.050 736.050 ;
        RECT 467.400 730.050 468.450 733.950 ;
        RECT 470.400 733.050 471.450 758.400 ;
        RECT 473.400 736.050 474.450 760.950 ;
        RECT 476.400 754.050 477.450 760.950 ;
        RECT 485.400 757.050 486.450 761.400 ;
        RECT 491.400 760.050 492.450 781.950 ;
        RECT 494.400 772.050 495.450 799.950 ;
        RECT 496.950 784.950 499.050 787.050 ;
        RECT 493.950 769.950 496.050 772.050 ;
        RECT 494.400 763.050 495.450 769.950 ;
        RECT 497.400 769.050 498.450 784.950 ;
        RECT 496.950 766.950 499.050 769.050 ;
        RECT 493.950 760.950 496.050 763.050 ;
        RECT 490.950 757.950 493.050 760.050 ;
        RECT 500.400 757.050 501.450 799.950 ;
        RECT 521.400 793.050 522.450 799.950 ;
        RECT 520.950 790.950 523.050 793.050 ;
        RECT 532.950 790.950 535.050 796.050 ;
        RECT 533.400 778.050 534.450 790.950 ;
        RECT 536.400 787.050 537.450 799.950 ;
        RECT 539.400 796.050 540.450 802.950 ;
        RECT 542.400 799.050 543.450 802.950 ;
        RECT 566.400 802.050 567.450 805.950 ;
        RECT 550.950 799.950 553.050 802.050 ;
        RECT 556.950 799.950 559.050 802.050 ;
        RECT 565.950 799.950 568.050 802.050 ;
        RECT 541.950 796.950 547.050 799.050 ;
        RECT 551.400 796.050 552.450 799.950 ;
        RECT 538.950 793.950 541.050 796.050 ;
        RECT 550.950 793.950 553.050 796.050 ;
        RECT 535.950 784.950 538.050 787.050 ;
        RECT 539.400 784.050 540.450 793.950 ;
        RECT 538.950 781.950 541.050 784.050 ;
        RECT 532.950 775.950 535.050 778.050 ;
        RECT 508.950 766.950 511.050 769.050 ;
        RECT 523.950 766.950 529.050 769.050 ;
        RECT 509.400 763.050 510.450 766.950 ;
        RECT 539.400 766.050 540.450 781.950 ;
        RECT 557.400 778.050 558.450 799.950 ;
        RECT 569.400 790.050 570.450 805.950 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 571.950 799.950 577.050 802.050 ;
        RECT 568.950 787.950 571.050 790.050 ;
        RECT 565.950 781.950 568.050 784.050 ;
        RECT 561.000 780.450 565.050 781.050 ;
        RECT 560.400 778.950 565.050 780.450 ;
        RECT 556.950 775.950 559.050 778.050 ;
        RECT 544.950 772.950 547.050 775.050 ;
        RECT 538.950 763.950 541.050 766.050 ;
        RECT 508.950 760.950 511.050 763.050 ;
        RECT 514.950 760.950 520.050 763.050 ;
        RECT 526.950 760.950 529.050 763.050 ;
        RECT 484.950 754.950 487.050 757.050 ;
        RECT 499.950 754.950 502.050 757.050 ;
        RECT 475.950 751.950 478.050 754.050 ;
        RECT 493.950 751.950 496.050 754.050 ;
        RECT 511.950 751.950 514.050 757.050 ;
        RECT 475.950 742.950 478.050 745.050 ;
        RECT 472.950 733.950 475.050 736.050 ;
        RECT 469.950 730.950 472.050 733.050 ;
        RECT 476.400 730.050 477.450 742.950 ;
        RECT 460.950 725.100 463.050 730.050 ;
        RECT 466.950 727.950 469.050 730.050 ;
        RECT 472.950 727.950 475.050 730.050 ;
        RECT 475.950 727.950 478.050 730.050 ;
        RECT 487.950 727.950 493.050 730.050 ;
        RECT 451.950 721.950 454.050 724.050 ;
        RECT 462.000 723.900 466.050 724.050 ;
        RECT 460.950 723.450 466.050 723.900 ;
        RECT 458.400 722.400 466.050 723.450 ;
        RECT 448.950 718.950 451.050 721.050 ;
        RECT 425.400 691.050 426.450 718.950 ;
        RECT 431.400 711.450 432.450 718.950 ;
        RECT 431.400 710.400 435.450 711.450 ;
        RECT 424.950 688.950 427.050 691.050 ;
        RECT 421.950 685.950 424.050 688.050 ;
        RECT 430.950 685.950 433.050 688.050 ;
        RECT 415.950 682.950 421.050 685.050 ;
        RECT 361.950 677.400 372.450 678.450 ;
        RECT 361.950 676.950 364.050 677.400 ;
        RECT 391.950 676.950 397.050 679.050 ;
        RECT 409.950 676.950 412.050 679.050 ;
        RECT 412.950 676.950 418.050 679.050 ;
        RECT 367.950 673.950 370.050 676.050 ;
        RECT 343.950 670.950 346.050 673.050 ;
        RECT 364.950 661.950 367.050 664.050 ;
        RECT 340.950 652.050 343.050 652.200 ;
        RECT 343.950 652.050 346.050 652.200 ;
        RECT 365.400 652.050 366.450 661.950 ;
        RECT 368.400 658.050 369.450 673.950 ;
        RECT 370.950 664.950 373.050 667.050 ;
        RECT 367.950 655.950 370.050 658.050 ;
        RECT 335.400 650.400 339.450 651.450 ;
        RECT 310.950 640.950 313.050 643.050 ;
        RECT 325.950 640.950 328.050 643.050 ;
        RECT 331.950 640.950 334.050 643.050 ;
        RECT 308.400 638.400 312.450 639.450 ;
        RECT 301.950 634.950 304.050 637.050 ;
        RECT 293.400 611.400 297.450 612.450 ;
        RECT 289.950 608.100 292.050 610.200 ;
        RECT 293.400 607.050 294.450 611.400 ;
        RECT 289.950 601.950 292.050 606.900 ;
        RECT 292.950 604.950 295.050 607.050 ;
        RECT 295.950 604.950 298.050 610.050 ;
        RECT 296.400 589.050 297.450 604.950 ;
        RECT 298.950 595.950 301.050 601.050 ;
        RECT 295.950 586.950 298.050 589.050 ;
        RECT 284.400 584.400 289.050 586.050 ;
        RECT 285.000 583.950 289.050 584.400 ;
        RECT 298.950 583.950 301.050 586.050 ;
        RECT 277.950 580.950 280.050 583.050 ;
        RECT 289.950 580.950 292.050 583.050 ;
        RECT 271.950 577.950 274.050 580.050 ;
        RECT 278.400 574.050 279.450 580.950 ;
        RECT 290.400 574.050 291.450 580.950 ;
        RECT 295.950 577.950 298.050 580.050 ;
        RECT 292.950 574.950 295.050 577.050 ;
        RECT 277.950 571.950 280.050 574.050 ;
        RECT 283.950 571.950 286.050 574.050 ;
        RECT 289.950 571.950 292.050 574.050 ;
        RECT 277.950 565.950 280.050 568.050 ;
        RECT 268.950 532.950 271.050 535.050 ;
        RECT 278.400 529.050 279.450 565.950 ;
        RECT 271.950 525.450 274.050 529.050 ;
        RECT 277.950 526.950 280.050 529.050 ;
        RECT 269.400 525.000 274.050 525.450 ;
        RECT 269.400 524.400 273.450 525.000 ;
        RECT 265.950 520.950 268.050 523.050 ;
        RECT 265.950 505.950 268.050 508.050 ;
        RECT 266.400 454.200 267.450 505.950 ;
        RECT 269.400 505.050 270.450 524.400 ;
        RECT 284.400 523.050 285.450 571.950 ;
        RECT 293.400 570.450 294.450 574.950 ;
        RECT 290.400 569.400 294.450 570.450 ;
        RECT 290.400 532.050 291.450 569.400 ;
        RECT 296.400 568.050 297.450 577.950 ;
        RECT 299.400 576.450 300.450 583.950 ;
        RECT 302.400 583.050 303.450 634.950 ;
        RECT 311.400 613.200 312.450 638.400 ;
        RECT 313.950 634.950 316.050 640.050 ;
        RECT 319.950 634.950 322.050 637.050 ;
        RECT 320.400 631.050 321.450 634.950 ;
        RECT 319.800 628.950 321.900 631.050 ;
        RECT 323.100 628.950 325.200 631.050 ;
        RECT 310.950 611.100 313.050 613.200 ;
        RECT 310.950 607.800 313.050 609.900 ;
        RECT 304.950 598.950 307.050 604.050 ;
        RECT 301.950 580.950 304.050 583.050 ;
        RECT 299.400 575.400 303.450 576.450 ;
        RECT 298.950 571.950 301.050 574.050 ;
        RECT 292.950 565.950 295.050 568.050 ;
        RECT 295.950 565.950 298.050 568.050 ;
        RECT 293.400 547.050 294.450 565.950 ;
        RECT 299.400 562.050 300.450 571.950 ;
        RECT 302.400 571.050 303.450 575.400 ;
        RECT 305.400 574.050 306.450 598.950 ;
        RECT 311.400 586.050 312.450 607.800 ;
        RECT 320.400 604.050 321.450 628.950 ;
        RECT 323.400 610.050 324.450 628.950 ;
        RECT 326.400 616.050 327.450 640.950 ;
        RECT 325.950 613.950 328.050 616.050 ;
        RECT 338.400 610.050 339.450 650.400 ;
        RECT 340.950 650.100 346.050 652.050 ;
        RECT 342.000 649.950 345.000 650.100 ;
        RECT 340.800 646.800 342.900 648.900 ;
        RECT 344.100 646.800 346.200 648.900 ;
        RECT 352.950 646.950 355.050 652.050 ;
        RECT 364.950 649.950 367.050 652.050 ;
        RECT 341.400 625.050 342.450 646.800 ;
        RECT 344.400 631.050 345.450 646.800 ;
        RECT 346.950 634.950 349.050 640.050 ;
        RECT 343.950 628.950 346.050 631.050 ;
        RECT 340.950 622.950 343.050 625.050 ;
        RECT 340.950 613.950 343.050 616.050 ;
        RECT 322.950 607.950 325.050 610.050 ;
        RECT 325.950 607.950 328.050 610.050 ;
        RECT 331.950 607.950 334.050 610.050 ;
        RECT 337.950 607.950 340.050 610.050 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 320.400 600.450 321.450 601.950 ;
        RECT 317.400 599.400 321.450 600.450 ;
        RECT 313.950 595.950 316.050 598.050 ;
        RECT 310.950 583.950 313.050 586.050 ;
        RECT 304.950 571.950 307.050 574.050 ;
        RECT 301.950 568.950 304.050 571.050 ;
        RECT 298.950 559.950 301.050 562.050 ;
        RECT 292.950 544.950 295.050 547.050 ;
        RECT 298.950 538.950 301.050 541.050 ;
        RECT 289.950 529.950 292.050 532.050 ;
        RECT 295.950 530.100 298.050 535.050 ;
        RECT 280.950 520.950 285.450 523.050 ;
        RECT 271.950 511.950 274.050 514.050 ;
        RECT 268.950 502.950 271.050 505.050 ;
        RECT 272.400 496.050 273.450 511.950 ;
        RECT 284.400 502.050 285.450 520.950 ;
        RECT 290.400 510.450 291.450 529.950 ;
        RECT 295.950 523.950 298.050 528.900 ;
        RECT 290.400 509.400 294.450 510.450 ;
        RECT 286.950 505.950 289.050 508.050 ;
        RECT 283.950 499.950 286.050 502.050 ;
        RECT 268.950 493.950 271.050 496.050 ;
        RECT 271.950 493.950 274.050 496.050 ;
        RECT 269.400 490.050 270.450 493.950 ;
        RECT 268.950 487.950 271.050 490.050 ;
        RECT 272.400 478.050 273.450 493.950 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 284.400 487.050 285.450 490.950 ;
        RECT 287.400 490.050 288.450 505.950 ;
        RECT 286.950 487.950 289.050 490.050 ;
        RECT 274.950 484.950 277.050 487.050 ;
        RECT 280.950 484.950 283.050 487.050 ;
        RECT 283.950 484.950 286.050 487.050 ;
        RECT 271.950 475.950 274.050 478.050 ;
        RECT 265.950 452.100 268.050 454.200 ;
        RECT 265.950 448.800 268.050 450.900 ;
        RECT 268.950 448.950 274.050 451.050 ;
        RECT 262.950 445.950 265.050 448.050 ;
        RECT 256.950 439.950 259.050 445.050 ;
        RECT 259.950 442.950 262.050 445.050 ;
        RECT 257.400 430.200 258.450 439.950 ;
        RECT 263.400 436.050 264.450 445.950 ;
        RECT 262.950 433.950 265.050 436.050 ;
        RECT 256.950 428.100 259.050 430.200 ;
        RECT 266.400 427.050 267.450 448.800 ;
        RECT 275.400 445.050 276.450 484.950 ;
        RECT 281.400 478.050 282.450 484.950 ;
        RECT 289.950 480.450 292.050 484.050 ;
        RECT 287.400 480.000 292.050 480.450 ;
        RECT 287.400 479.400 291.450 480.000 ;
        RECT 280.950 475.950 283.050 478.050 ;
        RECT 268.950 442.950 271.050 445.050 ;
        RECT 274.800 442.950 276.900 445.050 ;
        RECT 277.950 442.950 280.050 445.050 ;
        RECT 256.950 424.800 259.050 426.900 ;
        RECT 265.950 424.950 268.050 427.050 ;
        RECT 232.950 415.950 235.050 418.050 ;
        RECT 246.000 417.900 250.050 418.050 ;
        RECT 244.950 416.100 250.050 417.900 ;
        RECT 244.950 415.950 249.000 416.100 ;
        RECT 250.950 415.950 253.050 418.050 ;
        RECT 244.950 415.800 247.050 415.950 ;
        RECT 217.800 414.000 219.900 415.050 ;
        RECT 217.800 412.950 220.050 414.000 ;
        RECT 221.100 412.950 223.200 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 217.950 409.950 220.050 412.950 ;
        RECT 241.950 406.950 244.050 412.050 ;
        RECT 242.400 394.050 243.450 406.950 ;
        RECT 241.950 391.950 244.050 394.050 ;
        RECT 245.400 385.050 246.450 415.800 ;
        RECT 247.950 409.950 250.050 414.900 ;
        RECT 257.400 412.050 258.450 424.800 ;
        RECT 269.400 424.050 270.450 442.950 ;
        RECT 268.950 421.950 271.050 424.050 ;
        RECT 259.950 418.950 262.050 421.050 ;
        RECT 274.950 418.950 277.050 421.050 ;
        RECT 253.950 410.400 258.450 412.050 ;
        RECT 253.950 409.950 258.000 410.400 ;
        RECT 260.400 409.050 261.450 418.950 ;
        RECT 262.950 415.950 268.050 418.050 ;
        RECT 268.950 414.450 271.050 418.050 ;
        RECT 266.400 414.000 271.050 414.450 ;
        RECT 266.400 413.400 270.450 414.000 ;
        RECT 259.950 406.950 262.050 409.050 ;
        RECT 244.950 382.950 247.050 385.050 ;
        RECT 266.400 376.050 267.450 413.400 ;
        RECT 275.400 412.050 276.450 418.950 ;
        RECT 278.400 418.050 279.450 442.950 ;
        RECT 287.400 442.050 288.450 479.400 ;
        RECT 289.950 448.950 292.050 454.050 ;
        RECT 293.400 451.050 294.450 509.400 ;
        RECT 299.400 496.050 300.450 538.950 ;
        RECT 302.400 538.200 303.450 568.950 ;
        RECT 314.400 550.200 315.450 595.950 ;
        RECT 317.400 571.050 318.450 599.400 ;
        RECT 322.950 571.950 325.050 574.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 313.950 548.100 316.050 550.200 ;
        RECT 313.950 544.800 316.050 546.900 ;
        RECT 307.950 538.950 310.050 541.050 ;
        RECT 301.950 536.100 304.050 538.200 ;
        RECT 301.950 529.950 304.050 534.900 ;
        RECT 308.400 532.050 309.450 538.950 ;
        RECT 307.950 529.950 310.050 532.050 ;
        RECT 307.950 523.950 310.050 526.050 ;
        RECT 298.950 493.950 301.050 496.050 ;
        RECT 304.950 487.950 307.050 493.050 ;
        RECT 298.950 484.950 301.050 487.050 ;
        RECT 299.400 481.050 300.450 484.950 ;
        RECT 298.950 478.950 301.050 481.050 ;
        RECT 308.400 460.050 309.450 523.950 ;
        RECT 314.400 505.050 315.450 544.800 ;
        RECT 317.400 535.050 318.450 568.950 ;
        RECT 323.400 568.050 324.450 571.950 ;
        RECT 326.400 568.050 327.450 607.950 ;
        RECT 328.950 601.950 331.050 604.050 ;
        RECT 329.400 574.050 330.450 601.950 ;
        RECT 332.400 592.050 333.450 607.950 ;
        RECT 334.950 601.950 337.050 607.050 ;
        RECT 331.950 589.950 334.050 592.050 ;
        RECT 337.950 586.950 340.050 589.050 ;
        RECT 334.950 580.950 337.050 583.050 ;
        RECT 335.400 574.050 336.450 580.950 ;
        RECT 328.950 571.950 331.050 574.050 ;
        RECT 334.950 571.950 337.050 574.050 ;
        RECT 338.400 568.050 339.450 586.950 ;
        RECT 323.400 566.400 328.050 568.050 ;
        RECT 324.000 565.950 328.050 566.400 ;
        RECT 337.950 565.950 340.050 568.050 ;
        RECT 341.400 541.050 342.450 613.950 ;
        RECT 353.400 613.050 354.450 646.950 ;
        RECT 355.950 631.950 358.050 634.050 ;
        RECT 352.950 610.950 355.050 613.050 ;
        RECT 349.950 604.950 352.050 607.050 ;
        RECT 343.950 601.950 349.050 604.050 ;
        RECT 350.400 601.050 351.450 604.950 ;
        RECT 349.950 598.950 352.050 601.050 ;
        RECT 356.400 576.450 357.450 631.950 ;
        RECT 365.400 628.050 366.450 649.950 ;
        RECT 368.400 646.050 369.450 655.950 ;
        RECT 367.950 643.950 370.050 646.050 ;
        RECT 371.400 634.050 372.450 664.950 ;
        RECT 392.400 664.050 393.450 676.950 ;
        RECT 391.950 661.950 394.050 664.050 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 388.950 646.950 391.050 652.050 ;
        RECT 394.950 649.950 400.050 652.050 ;
        RECT 406.950 649.950 409.050 652.050 ;
        RECT 383.400 643.050 384.450 646.950 ;
        RECT 400.950 643.950 403.050 646.050 ;
        RECT 403.950 643.950 406.050 649.050 ;
        RECT 382.950 640.950 385.050 643.050 ;
        RECT 370.950 631.950 373.050 634.050 ;
        RECT 364.950 625.950 367.050 628.050 ;
        RECT 373.950 625.950 376.050 628.050 ;
        RECT 361.950 607.950 364.050 610.050 ;
        RECT 358.950 601.950 361.050 604.050 ;
        RECT 359.400 595.050 360.450 601.950 ;
        RECT 358.950 592.950 361.050 595.050 ;
        RECT 362.400 577.050 363.450 607.950 ;
        RECT 374.400 604.050 375.450 625.950 ;
        RECT 376.950 604.950 382.050 607.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 385.950 601.950 388.050 607.050 ;
        RECT 388.950 604.950 391.050 607.050 ;
        RECT 368.400 577.050 369.450 601.950 ;
        RECT 376.950 598.950 379.050 601.050 ;
        RECT 379.950 598.950 385.050 601.050 ;
        RECT 370.950 592.950 373.050 595.050 ;
        RECT 371.400 583.050 372.450 592.950 ;
        RECT 370.950 580.950 373.050 583.050 ;
        RECT 353.400 575.400 357.450 576.450 ;
        RECT 343.950 568.950 346.050 571.050 ;
        RECT 346.950 568.950 349.050 571.050 ;
        RECT 344.400 565.050 345.450 568.950 ;
        RECT 347.400 565.050 348.450 568.950 ;
        RECT 353.400 568.200 354.450 575.400 ;
        RECT 361.950 574.950 364.050 577.050 ;
        RECT 367.950 574.950 370.050 577.050 ;
        RECT 364.950 573.450 367.050 574.050 ;
        RECT 356.400 572.400 367.050 573.450 ;
        RECT 352.950 566.100 355.050 568.200 ;
        RECT 343.950 562.950 346.050 565.050 ;
        RECT 346.950 562.950 349.050 565.050 ;
        RECT 352.950 559.950 355.050 564.900 ;
        RECT 350.100 556.950 352.200 559.050 ;
        RECT 319.950 538.950 322.050 541.050 ;
        RECT 340.950 538.950 343.050 541.050 ;
        RECT 316.950 532.950 319.050 535.050 ;
        RECT 320.400 532.050 321.450 538.950 ;
        RECT 322.950 532.950 325.050 535.050 ;
        RECT 319.950 529.950 322.050 532.050 ;
        RECT 323.400 514.050 324.450 532.950 ;
        RECT 325.950 529.950 331.050 532.050 ;
        RECT 339.000 528.450 343.050 529.050 ;
        RECT 338.400 526.950 343.050 528.450 ;
        RECT 346.950 526.950 349.050 529.050 ;
        RECT 325.950 523.950 328.050 526.050 ;
        RECT 322.950 513.450 325.050 514.050 ;
        RECT 320.400 512.400 325.050 513.450 ;
        RECT 313.950 502.950 316.050 505.050 ;
        RECT 310.950 493.950 313.050 496.050 ;
        RECT 313.950 493.950 316.050 496.050 ;
        RECT 311.400 490.050 312.450 493.950 ;
        RECT 310.950 487.950 313.050 490.050 ;
        RECT 314.400 481.050 315.450 493.950 ;
        RECT 320.400 492.450 321.450 512.400 ;
        RECT 322.950 511.950 325.050 512.400 ;
        RECT 317.400 491.400 321.450 492.450 ;
        RECT 313.950 478.950 316.050 481.050 ;
        RECT 301.950 457.950 304.050 460.050 ;
        RECT 307.950 457.950 310.050 460.050 ;
        RECT 292.950 448.950 295.050 451.050 ;
        RECT 295.950 448.950 298.050 454.050 ;
        RECT 293.400 445.050 294.450 448.950 ;
        RECT 302.400 448.050 303.450 457.950 ;
        RECT 304.950 454.950 307.050 457.050 ;
        RECT 301.950 447.450 304.050 448.050 ;
        RECT 299.400 446.400 304.050 447.450 ;
        RECT 292.950 442.950 295.050 445.050 ;
        RECT 286.950 439.950 289.050 442.050 ;
        RECT 299.400 424.050 300.450 446.400 ;
        RECT 301.950 445.950 304.050 446.400 ;
        RECT 305.400 445.050 306.450 454.950 ;
        RECT 307.950 448.950 310.050 451.050 ;
        RECT 304.950 442.950 307.050 445.050 ;
        RECT 308.400 442.050 309.450 448.950 ;
        RECT 310.950 445.950 313.050 448.050 ;
        RECT 307.950 439.950 310.050 442.050 ;
        RECT 311.400 436.050 312.450 445.950 ;
        RECT 317.400 442.050 318.450 491.400 ;
        RECT 319.950 487.950 325.050 490.050 ;
        RECT 326.400 463.050 327.450 523.950 ;
        RECT 328.950 505.950 331.050 508.050 ;
        RECT 329.400 496.050 330.450 505.950 ;
        RECT 328.950 493.950 331.050 496.050 ;
        RECT 338.400 493.050 339.450 526.950 ;
        RECT 340.950 520.950 346.050 523.050 ;
        RECT 347.400 519.450 348.450 526.950 ;
        RECT 350.400 523.050 351.450 556.950 ;
        RECT 352.950 535.950 355.050 538.050 ;
        RECT 349.950 520.950 352.050 523.050 ;
        RECT 344.400 518.400 348.450 519.450 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 337.950 486.450 343.050 487.050 ;
        RECT 344.400 486.450 345.450 518.400 ;
        RECT 353.400 511.050 354.450 535.950 ;
        RECT 352.950 508.950 355.050 511.050 ;
        RECT 349.950 500.400 352.050 502.500 ;
        RECT 346.950 493.950 349.050 499.050 ;
        RECT 337.950 485.400 345.450 486.450 ;
        RECT 350.850 485.400 352.050 500.400 ;
        RECT 337.950 484.950 343.050 485.400 ;
        RECT 349.950 483.300 352.050 485.400 ;
        RECT 350.850 479.700 352.050 483.300 ;
        RECT 349.950 477.600 352.050 479.700 ;
        RECT 352.950 469.950 355.050 472.050 ;
        RECT 328.950 466.950 331.050 469.050 ;
        RECT 325.950 460.950 328.050 463.050 ;
        RECT 326.400 454.200 327.450 460.950 ;
        RECT 319.950 448.950 322.050 454.050 ;
        RECT 325.950 452.100 328.050 454.200 ;
        RECT 322.950 451.050 325.050 451.200 ;
        RECT 322.950 450.900 327.000 451.050 ;
        RECT 322.950 449.100 328.050 450.900 ;
        RECT 324.000 448.950 328.050 449.100 ;
        RECT 325.950 448.800 328.050 448.950 ;
        RECT 322.950 442.950 325.050 447.900 ;
        RECT 329.400 445.050 330.450 466.950 ;
        RECT 343.950 459.300 346.050 461.400 ;
        RECT 344.850 455.700 346.050 459.300 ;
        RECT 331.950 448.950 334.050 454.050 ;
        RECT 343.950 453.600 346.050 455.700 ;
        RECT 328.950 442.950 331.050 445.050 ;
        RECT 316.950 439.950 319.050 442.050 ;
        RECT 340.950 439.950 343.050 445.050 ;
        RECT 344.850 438.600 346.050 453.600 ;
        RECT 353.400 448.050 354.450 469.950 ;
        RECT 356.400 466.050 357.450 572.400 ;
        RECT 364.950 571.950 367.050 572.400 ;
        RECT 370.950 571.950 373.050 574.050 ;
        RECT 358.950 568.950 361.050 571.050 ;
        RECT 359.400 517.050 360.450 568.950 ;
        RECT 361.950 562.950 364.050 568.050 ;
        RECT 367.950 565.950 370.050 571.050 ;
        RECT 368.400 559.050 369.450 565.950 ;
        RECT 371.400 562.050 372.450 571.950 ;
        RECT 370.950 559.950 373.050 562.050 ;
        RECT 367.950 556.950 370.050 559.050 ;
        RECT 364.950 529.950 370.050 532.050 ;
        RECT 371.400 531.450 372.450 559.950 ;
        RECT 377.400 550.050 378.450 598.950 ;
        RECT 386.400 592.050 387.450 601.950 ;
        RECT 385.950 589.950 388.050 592.050 ;
        RECT 382.950 583.950 385.050 586.050 ;
        RECT 383.400 574.050 384.450 583.950 ;
        RECT 382.950 571.950 385.050 574.050 ;
        RECT 383.400 568.050 384.450 571.950 ;
        RECT 382.950 565.950 385.050 568.050 ;
        RECT 389.400 556.050 390.450 604.950 ;
        RECT 391.950 598.950 394.050 604.050 ;
        RECT 394.950 595.950 397.050 598.050 ;
        RECT 395.400 571.050 396.450 595.950 ;
        RECT 401.400 592.050 402.450 643.950 ;
        RECT 407.400 640.050 408.450 649.950 ;
        RECT 412.950 646.950 415.050 649.050 ;
        RECT 409.950 640.950 412.050 646.050 ;
        RECT 406.950 637.950 409.050 640.050 ;
        RECT 409.950 595.950 412.050 601.050 ;
        RECT 397.800 589.950 399.900 592.050 ;
        RECT 401.100 589.950 403.200 592.050 ;
        RECT 398.400 571.200 399.450 589.950 ;
        RECT 413.400 586.050 414.450 646.950 ;
        RECT 415.950 628.950 418.050 631.050 ;
        RECT 416.400 625.050 417.450 628.950 ;
        RECT 415.950 622.950 418.050 625.050 ;
        RECT 419.400 622.050 420.450 682.950 ;
        RECT 424.950 679.950 427.050 685.050 ;
        RECT 431.400 679.050 432.450 685.950 ;
        RECT 430.950 676.950 433.050 679.050 ;
        RECT 434.400 675.450 435.450 710.400 ;
        RECT 451.950 694.950 454.050 697.050 ;
        RECT 436.950 691.950 439.050 694.050 ;
        RECT 437.400 688.050 438.450 691.950 ;
        RECT 452.400 691.050 453.450 694.950 ;
        RECT 451.950 688.950 454.050 691.050 ;
        RECT 436.950 685.950 439.050 688.050 ;
        RECT 445.950 683.100 448.050 688.050 ;
        RECT 436.950 679.950 439.050 682.050 ;
        RECT 442.950 681.900 447.000 682.050 ;
        RECT 442.950 679.950 448.050 681.900 ;
        RECT 431.400 674.400 435.450 675.450 ;
        RECT 424.950 670.950 427.050 673.050 ;
        RECT 421.950 655.950 424.050 658.050 ;
        RECT 418.950 619.950 421.050 622.050 ;
        RECT 418.950 607.050 421.050 610.050 ;
        RECT 415.950 604.950 421.050 607.050 ;
        RECT 422.400 604.200 423.450 655.950 ;
        RECT 425.400 643.050 426.450 670.950 ;
        RECT 431.400 646.050 432.450 674.400 ;
        RECT 437.400 673.050 438.450 679.950 ;
        RECT 445.950 679.800 448.050 679.950 ;
        RECT 436.950 670.950 439.050 673.050 ;
        RECT 452.400 658.050 453.450 688.950 ;
        RECT 458.400 688.050 459.450 722.400 ;
        RECT 460.950 721.950 466.050 722.400 ;
        RECT 460.950 721.800 463.050 721.950 ;
        RECT 469.950 718.950 472.050 724.050 ;
        RECT 463.950 703.950 466.050 706.050 ;
        RECT 464.400 688.050 465.450 703.950 ;
        RECT 473.400 697.050 474.450 727.950 ;
        RECT 481.950 726.450 486.000 727.050 ;
        RECT 481.950 724.950 486.450 726.450 ;
        RECT 485.400 706.050 486.450 724.950 ;
        RECT 487.950 718.950 490.050 724.050 ;
        RECT 484.950 703.950 487.050 706.050 ;
        RECT 488.400 702.450 489.450 718.950 ;
        RECT 494.400 703.050 495.450 751.950 ;
        RECT 523.950 739.950 526.050 742.050 ;
        RECT 527.400 741.450 528.450 760.950 ;
        RECT 529.950 759.450 534.000 760.050 ;
        RECT 529.950 757.950 534.450 759.450 ;
        RECT 529.950 754.950 532.050 757.950 ;
        RECT 527.400 740.400 531.450 741.450 ;
        RECT 524.400 730.050 525.450 739.950 ;
        RECT 526.950 736.950 529.050 739.050 ;
        RECT 527.400 730.050 528.450 736.950 ;
        RECT 502.950 727.950 505.050 730.050 ;
        RECT 523.950 727.950 526.050 730.050 ;
        RECT 526.950 727.950 529.050 730.050 ;
        RECT 503.400 724.050 504.450 727.950 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 517.950 724.950 523.050 727.050 ;
        RECT 502.950 721.950 505.050 724.050 ;
        RECT 496.950 712.950 499.050 715.050 ;
        RECT 485.400 701.400 489.450 702.450 ;
        RECT 472.950 694.950 475.050 697.050 ;
        RECT 457.950 685.950 460.050 688.050 ;
        RECT 463.950 685.950 466.050 688.050 ;
        RECT 481.950 685.050 484.050 688.050 ;
        RECT 485.400 685.200 486.450 701.400 ;
        RECT 493.950 700.950 496.050 703.050 ;
        RECT 487.950 697.950 490.050 700.050 ;
        RECT 484.950 685.050 487.050 685.200 ;
        RECT 488.400 685.050 489.450 697.950 ;
        RECT 481.950 684.000 487.050 685.050 ;
        RECT 482.400 683.100 487.050 684.000 ;
        RECT 482.400 682.950 486.000 683.100 ;
        RECT 487.950 682.950 490.050 685.050 ;
        RECT 454.950 676.950 457.050 682.050 ;
        RECT 482.400 679.050 483.450 682.950 ;
        RECT 488.400 679.050 489.450 682.950 ;
        RECT 497.400 679.050 498.450 712.950 ;
        RECT 503.400 709.050 504.450 721.950 ;
        RECT 505.950 718.950 508.050 724.050 ;
        RECT 506.400 715.050 507.450 718.950 ;
        RECT 505.950 712.950 508.050 715.050 ;
        RECT 502.950 706.950 505.050 709.050 ;
        RECT 512.400 706.050 513.450 724.950 ;
        RECT 523.950 718.950 526.050 724.050 ;
        RECT 511.950 703.950 514.050 706.050 ;
        RECT 512.400 700.050 513.450 703.950 ;
        RECT 511.950 697.950 514.050 700.050 ;
        RECT 517.950 685.050 520.050 688.050 ;
        RECT 527.400 687.450 528.450 727.950 ;
        RECT 524.400 687.000 528.450 687.450 ;
        RECT 514.950 682.950 520.050 685.050 ;
        RECT 523.950 686.400 528.450 687.000 ;
        RECT 523.950 682.950 526.050 686.400 ;
        RECT 520.950 679.950 523.050 682.050 ;
        RECT 481.950 676.950 484.050 679.050 ;
        RECT 487.950 676.950 490.050 679.050 ;
        RECT 496.950 676.950 499.050 679.050 ;
        RECT 511.950 676.950 514.050 679.050 ;
        RECT 490.950 664.950 493.050 667.050 ;
        RECT 460.950 658.950 463.050 661.050 ;
        RECT 451.950 655.950 454.050 658.050 ;
        RECT 452.400 652.050 453.450 655.950 ;
        RECT 451.950 649.950 454.050 652.050 ;
        RECT 461.400 649.050 462.450 658.950 ;
        RECT 463.950 652.050 466.050 652.200 ;
        RECT 463.950 650.100 469.050 652.050 ;
        RECT 465.000 649.950 469.050 650.100 ;
        RECT 472.950 649.950 475.050 655.050 ;
        RECT 433.950 646.950 436.050 649.050 ;
        RECT 424.950 640.950 427.050 643.050 ;
        RECT 430.950 640.950 433.050 646.050 ;
        RECT 434.400 640.050 435.450 646.950 ;
        RECT 436.950 643.950 439.050 649.050 ;
        RECT 460.950 646.950 463.050 649.050 ;
        RECT 463.950 646.800 466.050 648.900 ;
        RECT 478.950 647.100 481.050 652.050 ;
        RECT 445.950 640.050 448.050 643.050 ;
        RECT 451.950 640.950 454.050 646.050 ;
        RECT 433.950 637.950 436.050 640.050 ;
        RECT 439.950 637.950 442.050 640.050 ;
        RECT 445.800 639.000 448.050 640.050 ;
        RECT 445.800 637.950 447.900 639.000 ;
        RECT 449.100 637.950 451.200 640.050 ;
        RECT 430.950 607.950 433.050 610.050 ;
        RECT 427.950 607.050 430.050 607.200 ;
        RECT 424.950 605.100 430.050 607.050 ;
        RECT 424.950 604.950 429.000 605.100 ;
        RECT 421.950 602.100 424.050 604.200 ;
        RECT 427.950 601.800 430.050 603.900 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 416.400 595.050 417.450 598.950 ;
        RECT 421.950 598.800 424.050 600.900 ;
        RECT 415.950 592.950 418.050 595.050 ;
        RECT 422.400 592.050 423.450 598.800 ;
        RECT 421.950 589.950 424.050 592.050 ;
        RECT 400.950 583.950 403.050 586.050 ;
        RECT 412.950 583.950 415.050 586.050 ;
        RECT 401.400 574.050 402.450 583.950 ;
        RECT 400.950 571.950 403.050 574.050 ;
        RECT 415.950 571.950 418.050 574.050 ;
        RECT 391.950 569.400 396.450 571.050 ;
        RECT 391.950 568.950 396.000 569.400 ;
        RECT 397.950 569.100 400.050 571.200 ;
        RECT 388.950 553.950 391.050 556.050 ;
        RECT 376.950 547.950 379.050 550.050 ;
        RECT 373.950 531.450 376.050 532.050 ;
        RECT 371.400 530.400 376.050 531.450 ;
        RECT 373.950 529.950 376.050 530.400 ;
        RECT 370.950 523.950 373.050 528.900 ;
        RECT 374.400 523.050 375.450 529.950 ;
        RECT 377.400 529.050 378.450 547.950 ;
        RECT 377.400 527.400 382.050 529.050 ;
        RECT 378.000 526.950 382.050 527.400 ;
        RECT 382.950 526.950 388.050 529.050 ;
        RECT 373.950 520.950 376.050 523.050 ;
        RECT 376.950 520.950 379.050 523.050 ;
        RECT 382.950 520.950 385.050 523.050 ;
        RECT 377.400 517.050 378.450 520.950 ;
        RECT 358.950 514.950 361.050 517.050 ;
        RECT 376.950 514.950 379.050 517.050 ;
        RECT 361.950 505.950 364.050 508.050 ;
        RECT 358.950 502.950 361.050 505.050 ;
        RECT 359.400 496.200 360.450 502.950 ;
        RECT 358.950 494.100 361.050 496.200 ;
        RECT 358.950 490.800 361.050 492.900 ;
        RECT 359.400 472.050 360.450 490.800 ;
        RECT 358.950 469.950 361.050 472.050 ;
        RECT 355.950 463.950 358.050 466.050 ;
        RECT 362.400 465.450 363.450 505.950 ;
        RECT 370.950 500.400 373.050 502.500 ;
        RECT 364.950 487.950 367.050 493.050 ;
        RECT 371.100 480.600 372.300 500.400 ;
        RECT 383.400 498.450 384.450 520.950 ;
        RECT 385.950 514.950 388.050 517.050 ;
        RECT 380.400 497.400 384.450 498.450 ;
        RECT 370.950 478.500 373.050 480.600 ;
        RECT 359.400 464.400 363.450 465.450 ;
        RECT 359.400 451.050 360.450 464.400 ;
        RECT 370.950 463.950 373.050 466.050 ;
        RECT 364.950 458.400 367.050 460.500 ;
        RECT 358.950 448.950 361.050 451.050 ;
        RECT 352.950 445.950 355.050 448.050 ;
        RECT 343.950 436.500 346.050 438.600 ;
        RECT 310.950 433.950 313.050 436.050 ;
        RECT 283.950 418.950 286.050 424.050 ;
        RECT 286.950 421.950 289.050 424.050 ;
        RECT 298.950 421.950 301.050 424.050 ;
        RECT 340.950 422.400 343.050 424.500 ;
        RECT 277.950 415.950 280.050 418.050 ;
        RECT 287.400 412.050 288.450 421.950 ;
        RECT 292.950 412.950 295.050 418.050 ;
        RECT 301.950 415.950 304.050 418.050 ;
        RECT 319.950 415.950 322.050 421.050 ;
        RECT 268.950 409.950 271.050 412.050 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 286.950 409.950 289.050 412.050 ;
        RECT 209.400 374.400 213.450 375.450 ;
        RECT 205.950 370.950 208.050 373.050 ;
        RECT 196.950 361.950 199.050 367.050 ;
        RECT 202.950 364.950 205.050 367.050 ;
        RECT 206.400 364.050 207.450 370.950 ;
        RECT 209.400 367.050 210.450 374.400 ;
        RECT 214.950 373.950 217.050 376.050 ;
        RECT 211.950 372.450 214.050 373.050 ;
        RECT 217.950 372.450 220.050 373.050 ;
        RECT 211.950 371.400 220.050 372.450 ;
        RECT 211.950 370.950 214.050 371.400 ;
        RECT 217.950 370.950 220.050 371.400 ;
        RECT 223.950 367.950 226.050 373.050 ;
        RECT 235.950 370.950 238.050 376.050 ;
        RECT 265.950 373.950 268.050 376.050 ;
        RECT 241.950 367.950 244.050 373.050 ;
        RECT 269.400 370.050 270.450 409.950 ;
        RECT 298.950 406.950 301.050 412.050 ;
        RECT 302.400 406.050 303.450 415.950 ;
        RECT 307.950 409.950 313.050 412.050 ;
        RECT 316.950 409.950 319.050 415.050 ;
        RECT 292.950 403.950 295.050 406.050 ;
        RECT 301.950 403.950 304.050 406.050 ;
        RECT 322.950 403.950 325.050 409.050 ;
        RECT 293.400 382.050 294.450 403.950 ;
        RECT 341.700 402.600 342.900 422.400 ;
        RECT 346.950 415.950 349.050 418.050 ;
        RECT 347.400 412.050 348.450 415.950 ;
        RECT 353.400 415.050 354.450 445.950 ;
        RECT 355.950 442.950 358.050 445.050 ;
        RECT 356.400 421.050 357.450 442.950 ;
        RECT 365.100 438.600 366.300 458.400 ;
        RECT 364.950 436.500 367.050 438.600 ;
        RECT 361.950 422.400 364.050 424.500 ;
        RECT 355.950 418.950 358.050 421.050 ;
        RECT 346.950 409.950 349.050 412.050 ;
        RECT 352.950 409.950 355.050 415.050 ;
        RECT 361.950 407.400 363.150 422.400 ;
        RECT 364.950 415.950 367.050 421.050 ;
        RECT 361.950 405.300 364.050 407.400 ;
        RECT 340.950 400.500 343.050 402.600 ;
        RECT 361.950 401.700 363.150 405.300 ;
        RECT 361.950 399.600 364.050 401.700 ;
        RECT 367.950 394.950 370.050 397.050 ;
        RECT 292.950 379.950 295.050 382.050 ;
        RECT 301.950 381.300 304.050 383.400 ;
        RECT 293.400 373.050 294.450 379.950 ;
        RECT 302.850 377.700 304.050 381.300 ;
        RECT 322.950 380.400 325.050 382.500 ;
        RECT 301.950 375.600 304.050 377.700 ;
        RECT 292.950 370.950 295.050 373.050 ;
        RECT 250.950 367.950 253.050 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 286.950 367.950 289.050 370.050 ;
        RECT 208.950 364.950 211.050 367.050 ;
        RECT 211.950 364.950 217.050 367.050 ;
        RECT 220.950 364.950 223.050 367.050 ;
        RECT 225.000 366.450 229.050 367.050 ;
        RECT 224.400 364.950 229.050 366.450 ;
        RECT 232.950 364.950 235.050 367.050 ;
        RECT 244.950 364.950 247.050 367.050 ;
        RECT 205.950 361.950 208.050 364.050 ;
        RECT 187.950 355.950 190.050 358.050 ;
        RECT 178.950 343.950 181.050 346.050 ;
        RECT 179.400 340.050 180.450 343.950 ;
        RECT 188.400 340.050 189.450 355.950 ;
        RECT 214.950 349.950 217.050 352.050 ;
        RECT 208.950 344.400 211.050 346.500 ;
        RECT 172.950 334.950 175.050 340.050 ;
        RECT 178.950 337.950 181.050 340.050 ;
        RECT 187.950 337.950 190.050 340.050 ;
        RECT 193.950 337.950 196.050 340.050 ;
        RECT 199.950 339.450 204.000 340.050 ;
        RECT 199.950 337.950 204.450 339.450 ;
        RECT 166.950 331.950 169.050 334.050 ;
        RECT 161.400 317.400 165.450 318.450 ;
        RECT 145.950 303.300 148.050 305.400 ;
        RECT 146.850 299.700 148.050 303.300 ;
        RECT 145.950 297.600 148.050 299.700 ;
        RECT 136.950 295.050 139.050 295.200 ;
        RECT 94.950 292.950 100.050 295.050 ;
        RECT 103.950 292.950 106.050 295.050 ;
        RECT 115.950 292.950 118.050 295.050 ;
        RECT 121.950 292.950 127.050 295.050 ;
        RECT 130.950 292.950 133.050 295.050 ;
        RECT 133.950 293.100 139.050 295.050 ;
        RECT 133.950 292.950 138.000 293.100 ;
        RECT 139.950 292.950 142.050 295.050 ;
        RECT 94.950 286.950 97.050 289.050 ;
        RECT 95.400 277.050 96.450 286.950 ;
        RECT 94.950 274.950 97.050 277.050 ;
        RECT 98.400 274.050 99.450 292.950 ;
        RECT 100.950 286.950 103.050 292.050 ;
        RECT 106.950 286.950 109.050 289.050 ;
        RECT 97.950 271.950 100.050 274.050 ;
        RECT 107.400 271.050 108.450 286.950 ;
        RECT 100.950 268.950 103.050 271.050 ;
        RECT 106.950 268.950 109.050 271.050 ;
        RECT 94.950 266.400 97.050 268.500 ;
        RECT 95.700 246.600 96.900 266.400 ;
        RECT 101.400 256.050 102.450 268.950 ;
        RECT 115.950 266.400 118.050 268.500 ;
        RECT 122.400 268.050 123.450 292.950 ;
        RECT 124.950 286.950 127.050 289.050 ;
        RECT 136.950 286.950 139.050 291.900 ;
        RECT 109.950 262.950 112.050 265.050 ;
        RECT 110.400 259.050 111.450 262.950 ;
        RECT 106.950 256.950 112.050 259.050 ;
        RECT 100.950 253.950 103.050 256.050 ;
        RECT 115.950 251.400 117.150 266.400 ;
        RECT 121.950 265.950 124.050 268.050 ;
        RECT 118.950 259.950 121.050 265.050 ;
        RECT 115.950 249.300 118.050 251.400 ;
        RECT 94.950 244.500 97.050 246.600 ;
        RECT 115.950 245.700 117.150 249.300 ;
        RECT 115.950 243.600 118.050 245.700 ;
        RECT 115.950 232.950 118.050 235.050 ;
        RECT 88.950 220.950 91.050 223.050 ;
        RECT 109.950 220.950 112.050 223.050 ;
        RECT 67.950 211.950 70.050 217.050 ;
        RECT 73.950 214.950 76.050 217.050 ;
        RECT 82.950 215.100 85.050 217.200 ;
        RECT 89.400 217.050 90.450 220.950 ;
        RECT 110.400 217.050 111.450 220.950 ;
        RECT 88.950 214.950 91.050 217.050 ;
        RECT 68.400 196.050 69.450 211.950 ;
        RECT 67.950 193.950 70.050 196.050 ;
        RECT 61.950 190.950 64.050 193.050 ;
        RECT 62.400 184.050 63.450 190.950 ;
        RECT 70.950 187.950 73.050 190.050 ;
        RECT 61.950 181.950 64.050 184.050 ;
        RECT 58.950 175.950 61.050 181.050 ;
        RECT 52.950 172.950 55.050 175.050 ;
        RECT 64.950 172.950 67.050 178.050 ;
        RECT 49.950 148.950 52.050 151.050 ;
        RECT 64.950 145.950 67.050 148.050 ;
        RECT 52.950 136.950 61.050 139.050 ;
        RECT 65.400 133.050 66.450 145.950 ;
        RECT 71.400 142.200 72.450 187.950 ;
        RECT 74.400 184.200 75.450 214.950 ;
        RECT 82.950 211.800 85.050 213.900 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 103.950 212.100 106.050 217.050 ;
        RECT 109.950 214.950 112.050 217.050 ;
        RECT 79.950 205.950 82.050 208.050 ;
        RECT 73.950 182.100 76.050 184.200 ;
        RECT 80.400 181.050 81.450 205.950 ;
        RECT 83.400 187.050 84.450 211.800 ;
        RECT 95.400 208.050 96.450 211.950 ;
        RECT 116.400 211.050 117.450 232.950 ;
        RECT 122.400 211.050 123.450 265.950 ;
        RECT 125.400 256.050 126.450 286.950 ;
        RECT 127.950 259.950 133.050 262.050 ;
        RECT 124.950 253.950 127.050 256.050 ;
        RECT 128.400 250.050 129.450 259.950 ;
        RECT 130.950 253.950 136.050 256.050 ;
        RECT 127.950 247.950 130.050 250.050 ;
        RECT 131.400 229.050 132.450 253.950 ;
        RECT 133.950 247.950 136.050 250.050 ;
        RECT 130.950 226.950 133.050 229.050 ;
        RECT 127.950 220.950 130.050 223.050 ;
        RECT 128.400 214.050 129.450 220.950 ;
        RECT 134.400 214.050 135.450 247.950 ;
        RECT 140.400 241.050 141.450 292.950 ;
        RECT 142.950 286.950 145.050 292.050 ;
        RECT 146.850 282.600 148.050 297.600 ;
        RECT 161.400 295.050 162.450 317.400 ;
        RECT 179.400 309.450 180.450 337.950 ;
        RECT 190.950 331.950 193.050 334.050 ;
        RECT 191.400 328.050 192.450 331.950 ;
        RECT 190.950 325.950 193.050 328.050 ;
        RECT 194.400 324.450 195.450 337.950 ;
        RECT 196.950 328.950 199.050 334.050 ;
        RECT 176.400 308.400 180.450 309.450 ;
        RECT 191.400 323.400 195.450 324.450 ;
        RECT 166.950 302.400 169.050 304.500 ;
        RECT 160.950 292.950 163.050 295.050 ;
        RECT 151.950 289.950 157.050 292.050 ;
        RECT 145.950 280.500 148.050 282.600 ;
        RECT 145.950 266.400 148.050 268.500 ;
        RECT 146.700 246.600 147.900 266.400 ;
        RECT 151.950 262.950 154.050 265.050 ;
        RECT 152.400 259.050 153.450 262.950 ;
        RECT 155.400 259.050 156.450 289.950 ;
        RECT 167.100 282.600 168.300 302.400 ;
        RECT 166.950 280.500 169.050 282.600 ;
        RECT 166.950 266.400 169.050 268.500 ;
        RECT 151.950 256.950 154.050 259.050 ;
        RECT 154.950 256.950 160.050 259.050 ;
        RECT 166.950 251.400 168.150 266.400 ;
        RECT 169.950 256.950 172.050 262.050 ;
        RECT 166.950 249.300 169.050 251.400 ;
        RECT 145.950 244.500 148.050 246.600 ;
        RECT 166.950 245.700 168.150 249.300 ;
        RECT 166.950 243.600 169.050 245.700 ;
        RECT 139.950 238.950 142.050 241.050 ;
        RECT 145.950 238.950 148.050 241.050 ;
        RECT 127.950 211.950 130.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 142.950 211.950 145.050 214.050 ;
        RECT 100.950 208.950 103.050 211.050 ;
        RECT 105.000 210.900 109.050 211.050 ;
        RECT 103.950 208.950 109.050 210.900 ;
        RECT 115.950 208.950 118.050 211.050 ;
        RECT 121.950 208.950 124.050 211.050 ;
        RECT 94.950 205.950 97.050 208.050 ;
        RECT 101.400 196.050 102.450 208.950 ;
        RECT 103.950 208.800 106.050 208.950 ;
        RECT 136.950 205.950 139.050 211.050 ;
        RECT 88.950 193.950 91.050 196.050 ;
        RECT 100.950 193.950 103.050 196.050 ;
        RECT 130.950 193.950 133.050 196.050 ;
        RECT 82.950 184.950 85.050 187.050 ;
        RECT 73.950 178.800 76.050 180.900 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 70.950 140.100 73.050 142.200 ;
        RECT 74.400 139.050 75.450 178.800 ;
        RECT 76.950 169.950 79.050 178.050 ;
        RECT 83.400 175.050 84.450 184.950 ;
        RECT 85.950 178.950 88.050 184.050 ;
        RECT 89.400 178.050 90.450 193.950 ;
        RECT 100.950 187.950 103.050 190.050 ;
        RECT 115.950 188.400 118.050 190.500 ;
        RECT 101.400 184.050 102.450 187.950 ;
        RECT 91.950 181.950 97.050 184.050 ;
        RECT 100.950 181.950 103.050 184.050 ;
        RECT 112.950 181.950 115.050 187.050 ;
        RECT 88.950 175.950 91.050 178.050 ;
        RECT 91.950 175.950 94.050 178.050 ;
        RECT 94.950 175.950 100.050 178.050 ;
        RECT 103.950 175.950 106.050 178.050 ;
        RECT 82.950 172.950 85.050 175.050 ;
        RECT 77.400 148.050 78.450 169.950 ;
        RECT 76.950 145.950 79.050 148.050 ;
        RECT 88.950 142.950 91.050 145.050 ;
        RECT 85.950 139.950 88.050 142.050 ;
        RECT 69.000 138.900 72.000 139.050 ;
        RECT 67.950 136.950 73.050 138.900 ;
        RECT 74.400 137.400 79.050 139.050 ;
        RECT 75.000 136.950 79.050 137.400 ;
        RECT 67.950 136.800 70.050 136.950 ;
        RECT 70.950 136.800 73.050 136.950 ;
        RECT 55.950 130.950 58.050 133.050 ;
        RECT 65.400 131.400 70.050 133.050 ;
        RECT 66.000 130.950 70.050 131.400 ;
        RECT 56.400 124.050 57.450 130.950 ;
        RECT 55.950 121.950 58.050 124.050 ;
        RECT 46.950 115.950 49.050 118.050 ;
        RECT 31.950 109.950 34.050 112.050 ;
        RECT 37.950 110.100 40.050 112.200 ;
        RECT 22.950 106.950 25.050 109.050 ;
        RECT 23.400 100.050 24.450 106.950 ;
        RECT 32.400 103.050 33.450 109.950 ;
        RECT 37.950 103.950 40.050 108.900 ;
        RECT 40.950 103.950 43.050 106.050 ;
        RECT 46.950 103.950 52.050 106.050 ;
        RECT 61.950 103.950 67.050 106.050 ;
        RECT 23.400 98.400 28.050 100.050 ;
        RECT 24.000 97.950 28.050 98.400 ;
        RECT 31.950 97.950 34.050 103.050 ;
        RECT 41.400 76.050 42.450 103.950 ;
        RECT 43.950 97.950 49.050 100.050 ;
        RECT 52.950 97.950 58.050 100.050 ;
        RECT 61.950 97.950 67.050 100.050 ;
        RECT 68.400 85.050 69.450 130.950 ;
        RECT 73.950 127.950 76.050 133.050 ;
        RECT 79.950 103.950 82.050 106.050 ;
        RECT 76.950 100.950 79.050 103.050 ;
        RECT 77.400 94.050 78.450 100.950 ;
        RECT 80.400 97.050 81.450 103.950 ;
        RECT 86.400 100.050 87.450 139.950 ;
        RECT 89.400 130.050 90.450 142.950 ;
        RECT 92.400 136.050 93.450 175.950 ;
        RECT 104.400 160.050 105.450 175.950 ;
        RECT 116.850 173.400 118.050 188.400 ;
        RECT 124.950 178.950 130.050 181.050 ;
        RECT 131.400 178.050 132.450 193.950 ;
        RECT 136.950 188.400 139.050 190.500 ;
        RECT 143.400 190.050 144.450 211.950 ;
        RECT 130.950 175.950 133.050 178.050 ;
        RECT 115.950 171.300 118.050 173.400 ;
        RECT 116.850 167.700 118.050 171.300 ;
        RECT 137.100 168.600 138.300 188.400 ;
        RECT 142.950 187.950 145.050 190.050 ;
        RECT 115.950 165.600 118.050 167.700 ;
        RECT 136.950 166.500 139.050 168.600 ;
        RECT 103.950 157.950 106.050 160.050 ;
        RECT 121.950 157.950 124.050 160.050 ;
        RECT 97.950 148.950 100.050 151.050 ;
        RECT 109.950 148.950 112.050 151.050 ;
        RECT 98.400 139.050 99.450 148.950 ;
        RECT 110.400 139.050 111.450 148.950 ;
        RECT 97.950 136.950 100.050 139.050 ;
        RECT 109.950 136.950 112.050 139.050 ;
        RECT 115.950 136.950 118.050 139.050 ;
        RECT 91.950 130.950 94.050 136.050 ;
        RECT 116.400 133.050 117.450 136.950 ;
        RECT 122.400 136.050 123.450 157.950 ;
        RECT 142.950 147.450 145.050 148.050 ;
        RECT 146.400 147.450 147.450 238.950 ;
        RECT 172.950 226.950 175.050 229.050 ;
        RECT 157.950 220.950 160.050 223.050 ;
        RECT 148.950 214.950 151.050 217.050 ;
        RECT 149.400 211.050 150.450 214.950 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 148.950 208.950 151.050 211.050 ;
        RECT 155.400 208.050 156.450 211.950 ;
        RECT 154.950 205.950 157.050 208.050 ;
        RECT 151.950 181.950 154.050 187.050 ;
        RECT 152.400 172.050 153.450 181.950 ;
        RECT 158.400 181.050 159.450 220.950 ;
        RECT 173.400 217.050 174.450 226.950 ;
        RECT 176.400 223.050 177.450 308.400 ;
        RECT 181.950 302.400 184.050 304.500 ;
        RECT 182.700 282.600 183.900 302.400 ;
        RECT 191.400 295.050 192.450 323.400 ;
        RECT 203.400 322.050 204.450 337.950 ;
        RECT 209.700 324.600 210.900 344.400 ;
        RECT 215.400 334.050 216.450 349.950 ;
        RECT 221.400 339.450 222.450 364.950 ;
        RECT 218.400 338.400 222.450 339.450 ;
        RECT 214.950 331.950 217.050 334.050 ;
        RECT 208.950 322.500 211.050 324.600 ;
        RECT 202.950 319.950 205.050 322.050 ;
        RECT 193.950 313.950 196.050 316.050 ;
        RECT 190.950 292.950 193.050 295.050 ;
        RECT 194.400 292.050 195.450 313.950 ;
        RECT 218.400 310.050 219.450 338.400 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 221.400 328.050 222.450 334.950 ;
        RECT 220.950 325.950 223.050 328.050 ;
        RECT 221.400 316.050 222.450 325.950 ;
        RECT 220.950 313.950 223.050 316.050 ;
        RECT 217.950 307.950 220.050 310.050 ;
        RECT 202.950 303.300 205.050 305.400 ;
        RECT 202.950 299.700 204.150 303.300 ;
        RECT 217.950 302.400 220.050 304.500 ;
        RECT 202.950 297.600 205.050 299.700 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 202.950 282.600 204.150 297.600 ;
        RECT 205.950 288.450 210.000 289.050 ;
        RECT 205.950 286.950 210.450 288.450 ;
        RECT 209.400 283.050 210.450 286.950 ;
        RECT 181.950 280.500 184.050 282.600 ;
        RECT 202.950 280.500 205.050 282.600 ;
        RECT 208.950 280.950 211.050 283.050 ;
        RECT 218.700 282.600 219.900 302.400 ;
        RECT 224.400 298.200 225.450 364.950 ;
        RECT 233.400 352.050 234.450 364.950 ;
        RECT 232.950 349.950 235.050 352.050 ;
        RECT 229.950 344.400 232.050 346.500 ;
        RECT 229.950 329.400 231.150 344.400 ;
        RECT 232.950 337.950 238.050 340.050 ;
        RECT 238.950 337.950 244.050 340.050 ;
        RECT 229.950 327.300 232.050 329.400 ;
        RECT 229.950 323.700 231.150 327.300 ;
        RECT 229.950 321.600 232.050 323.700 ;
        RECT 229.950 313.950 232.050 316.050 ;
        RECT 226.950 307.950 229.050 310.050 ;
        RECT 223.950 296.100 226.050 298.200 ;
        RECT 227.400 295.050 228.450 307.950 ;
        RECT 225.000 294.900 228.450 295.050 ;
        RECT 223.950 293.250 228.450 294.900 ;
        RECT 223.950 292.950 228.000 293.250 ;
        RECT 223.950 292.800 226.050 292.950 ;
        RECT 230.400 292.050 231.450 313.950 ;
        RECT 242.400 310.050 243.450 337.950 ;
        RECT 245.400 337.050 246.450 364.950 ;
        RECT 244.950 331.950 247.050 337.050 ;
        RECT 251.400 328.050 252.450 367.950 ;
        RECT 287.400 361.050 288.450 367.950 ;
        RECT 292.950 361.950 295.050 367.050 ;
        RECT 297.000 366.450 301.050 367.050 ;
        RECT 296.400 364.950 301.050 366.450 ;
        RECT 296.400 361.050 297.450 364.950 ;
        RECT 286.950 358.950 289.050 361.050 ;
        RECT 295.950 358.950 298.050 361.050 ;
        RECT 302.850 360.600 304.050 375.600 ;
        RECT 310.950 373.950 313.050 376.050 ;
        RECT 311.400 370.050 312.450 373.950 ;
        RECT 316.950 370.950 319.050 373.050 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 287.400 355.050 288.450 358.950 ;
        RECT 301.950 358.500 304.050 360.600 ;
        RECT 286.950 352.950 289.050 355.050 ;
        RECT 311.400 352.050 312.450 367.950 ;
        RECT 317.400 364.050 318.450 370.950 ;
        RECT 316.950 361.950 319.050 364.050 ;
        RECT 323.100 360.600 324.300 380.400 ;
        RECT 343.950 370.950 346.050 373.050 ;
        RECT 349.950 370.950 355.050 373.050 ;
        RECT 344.400 367.050 345.450 370.950 ;
        RECT 331.950 361.950 334.050 367.050 ;
        RECT 343.950 364.950 346.050 367.050 ;
        RECT 346.950 361.950 349.050 367.050 ;
        RECT 322.950 358.500 325.050 360.600 ;
        RECT 298.950 349.950 301.050 352.050 ;
        RECT 310.950 349.950 313.050 352.050 ;
        RECT 325.950 349.950 328.050 352.050 ;
        RECT 289.950 344.400 292.050 346.500 ;
        RECT 265.950 340.950 268.050 343.050 ;
        RECT 256.950 334.950 262.050 337.050 ;
        RECT 250.950 325.950 253.050 328.050 ;
        RECT 253.950 319.950 256.050 322.050 ;
        RECT 241.950 307.950 244.050 310.050 ;
        RECT 238.950 303.300 241.050 305.400 ;
        RECT 238.950 299.700 240.150 303.300 ;
        RECT 238.950 297.600 241.050 299.700 ;
        RECT 223.950 289.800 226.050 291.900 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 217.950 280.500 220.050 282.600 ;
        RECT 178.950 265.950 181.050 268.050 ;
        RECT 179.400 262.050 180.450 265.950 ;
        RECT 178.950 259.950 181.050 262.050 ;
        RECT 184.950 259.950 187.050 265.050 ;
        RECT 205.950 261.450 210.000 262.050 ;
        RECT 205.950 259.950 210.450 261.450 ;
        RECT 205.950 256.950 208.050 259.950 ;
        RECT 181.950 253.950 187.050 256.050 ;
        RECT 187.950 253.950 190.050 256.050 ;
        RECT 202.950 255.450 207.000 256.050 ;
        RECT 202.950 253.950 207.450 255.450 ;
        RECT 188.400 247.050 189.450 253.950 ;
        RECT 206.400 250.050 207.450 253.950 ;
        RECT 209.400 253.050 210.450 259.950 ;
        RECT 224.400 259.050 225.450 289.800 ;
        RECT 238.950 282.600 240.150 297.600 ;
        RECT 254.400 295.050 255.450 319.950 ;
        RECT 253.950 292.950 259.050 295.050 ;
        RECT 259.950 289.950 262.050 295.050 ;
        RECT 241.950 288.450 246.000 289.050 ;
        RECT 241.950 286.950 246.450 288.450 ;
        RECT 250.950 286.950 256.050 289.050 ;
        RECT 238.950 280.500 241.050 282.600 ;
        RECT 229.950 268.950 232.050 271.050 ;
        RECT 220.950 256.950 226.050 259.050 ;
        RECT 211.950 253.950 214.050 256.050 ;
        RECT 226.950 253.950 229.050 259.050 ;
        RECT 208.950 250.950 211.050 253.050 ;
        RECT 212.400 250.050 213.450 253.950 ;
        RECT 205.950 247.950 208.050 250.050 ;
        RECT 211.950 247.950 214.050 250.050 ;
        RECT 187.950 244.950 190.050 247.050 ;
        RECT 230.400 223.050 231.450 268.950 ;
        RECT 232.950 262.950 235.050 268.050 ;
        RECT 235.950 262.950 238.050 265.050 ;
        RECT 175.950 220.950 178.050 223.050 ;
        RECT 205.950 217.950 208.050 220.050 ;
        RECT 211.950 217.950 214.050 223.050 ;
        RECT 229.950 220.950 232.050 223.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 172.950 211.950 175.050 217.050 ;
        RECT 181.950 214.950 187.050 217.050 ;
        RECT 190.950 214.950 196.050 217.050 ;
        RECT 196.950 211.950 199.050 217.050 ;
        RECT 202.950 214.950 205.050 217.050 ;
        RECT 163.950 205.950 166.050 211.050 ;
        RECT 167.400 199.050 168.450 211.950 ;
        RECT 203.400 211.050 204.450 214.950 ;
        RECT 206.400 211.050 207.450 217.950 ;
        RECT 220.950 214.950 226.050 217.050 ;
        RECT 229.950 214.950 235.050 217.050 ;
        RECT 223.950 211.950 226.050 214.950 ;
        RECT 236.400 214.050 237.450 262.950 ;
        RECT 245.400 262.050 246.450 286.950 ;
        RECT 251.400 283.050 252.450 286.950 ;
        RECT 256.950 283.950 259.050 286.050 ;
        RECT 250.950 280.950 253.050 283.050 ;
        RECT 257.400 271.050 258.450 283.950 ;
        RECT 266.400 277.050 267.450 340.950 ;
        RECT 280.950 337.950 283.050 340.050 ;
        RECT 283.950 337.950 289.050 340.050 ;
        RECT 271.950 331.950 274.050 337.050 ;
        RECT 274.950 331.950 280.050 334.050 ;
        RECT 281.400 301.050 282.450 337.950 ;
        RECT 290.850 329.400 292.050 344.400 ;
        RECT 299.400 337.050 300.450 349.950 ;
        RECT 310.950 344.400 313.050 346.500 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 304.950 334.950 307.050 340.050 ;
        RECT 289.950 327.300 292.050 329.400 ;
        RECT 290.850 323.700 292.050 327.300 ;
        RECT 289.950 321.600 292.050 323.700 ;
        RECT 283.950 307.950 286.050 310.050 ;
        RECT 280.950 298.950 283.050 301.050 ;
        RECT 274.950 292.950 280.050 295.050 ;
        RECT 284.400 292.050 285.450 307.950 ;
        RECT 289.950 298.950 292.050 301.050 ;
        RECT 290.400 295.050 291.450 298.950 ;
        RECT 299.400 298.050 300.450 334.950 ;
        RECT 304.950 328.950 307.050 331.050 ;
        RECT 298.950 295.950 301.050 298.050 ;
        RECT 289.950 292.950 292.050 295.050 ;
        RECT 283.950 289.950 286.050 292.050 ;
        RECT 295.950 286.950 298.050 292.050 ;
        RECT 292.950 283.950 295.050 286.050 ;
        RECT 265.950 274.950 268.050 277.050 ;
        RECT 256.950 268.950 259.050 271.050 ;
        RECT 280.950 265.950 283.050 268.050 ;
        RECT 259.950 262.950 262.050 265.050 ;
        RECT 265.950 262.950 271.050 265.050 ;
        RECT 244.950 256.950 247.050 262.050 ;
        RECT 250.950 256.950 256.050 259.050 ;
        RECT 260.400 256.050 261.450 262.950 ;
        RECT 281.400 262.050 282.450 265.950 ;
        RECT 286.950 262.950 289.050 265.050 ;
        RECT 268.950 256.950 274.050 259.050 ;
        RECT 280.950 256.950 283.050 262.050 ;
        RECT 241.950 250.950 244.050 256.050 ;
        RECT 260.400 254.400 265.050 256.050 ;
        RECT 261.000 253.950 265.050 254.400 ;
        RECT 283.950 253.950 286.050 256.050 ;
        RECT 250.950 250.950 253.050 253.050 ;
        RECT 241.950 235.950 244.050 238.050 ;
        RECT 242.400 217.050 243.450 235.950 ;
        RECT 241.950 214.950 244.050 217.050 ;
        RECT 235.950 211.950 238.050 214.050 ;
        RECT 181.950 208.950 184.050 211.050 ;
        RECT 202.950 208.950 205.050 211.050 ;
        RECT 205.950 208.950 208.050 211.050 ;
        RECT 214.950 208.950 217.050 211.050 ;
        RECT 220.950 208.950 223.050 211.050 ;
        RECT 226.950 208.950 229.050 211.050 ;
        RECT 169.950 205.950 175.050 208.050 ;
        RECT 182.400 199.050 183.450 208.950 ;
        RECT 166.950 196.950 169.050 199.050 ;
        RECT 181.950 196.950 184.050 199.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 167.400 178.050 168.450 196.950 ;
        RECT 193.950 190.950 196.050 193.050 ;
        RECT 169.950 187.950 172.050 190.050 ;
        RECT 178.950 188.400 181.050 190.500 ;
        RECT 170.400 184.050 171.450 187.950 ;
        RECT 169.950 181.950 172.050 184.050 ;
        RECT 172.950 181.950 178.050 184.050 ;
        RECT 166.950 175.950 169.050 178.050 ;
        RECT 179.850 173.400 181.050 188.400 ;
        RECT 194.400 181.050 195.450 190.950 ;
        RECT 199.950 188.400 202.050 190.500 ;
        RECT 215.400 190.050 216.450 208.950 ;
        RECT 221.400 205.050 222.450 208.950 ;
        RECT 220.950 202.950 223.050 205.050 ;
        RECT 227.400 202.050 228.450 208.950 ;
        RECT 232.950 202.950 235.050 205.050 ;
        RECT 226.950 199.950 229.050 202.050 ;
        RECT 217.950 196.950 220.050 199.050 ;
        RECT 187.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 151.950 169.950 154.050 172.050 ;
        RECT 178.950 171.300 181.050 173.400 ;
        RECT 179.850 167.700 181.050 171.300 ;
        RECT 184.950 169.950 187.050 172.050 ;
        RECT 178.950 165.600 181.050 167.700 ;
        RECT 142.950 146.400 147.450 147.450 ;
        RECT 142.950 145.950 145.050 146.400 ;
        RECT 157.950 145.950 160.050 148.050 ;
        RECT 127.950 139.950 130.050 145.050 ;
        RECT 133.950 139.950 136.050 142.050 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 103.950 130.950 109.050 133.050 ;
        RECT 112.950 130.950 115.050 133.050 ;
        RECT 115.950 130.950 118.050 133.050 ;
        RECT 88.950 127.950 91.050 130.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 103.950 100.950 109.050 103.050 ;
        RECT 79.950 94.950 82.050 97.050 ;
        RECT 85.950 94.950 88.050 100.050 ;
        RECT 92.400 97.050 93.450 100.950 ;
        RECT 113.400 97.050 114.450 130.950 ;
        RECT 122.400 100.050 123.450 133.950 ;
        RECT 134.400 130.050 135.450 139.950 ;
        RECT 143.400 136.050 144.450 145.950 ;
        RECT 158.400 142.050 159.450 145.950 ;
        RECT 151.950 136.950 154.050 142.050 ;
        RECT 157.950 139.950 160.050 142.050 ;
        RECT 160.950 139.950 166.050 142.050 ;
        RECT 175.950 136.950 178.050 142.050 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 160.950 133.950 163.050 136.050 ;
        RECT 157.950 130.950 160.050 133.050 ;
        RECT 133.950 127.950 136.050 130.050 ;
        RECT 145.950 127.950 148.050 130.050 ;
        RECT 146.400 108.450 147.450 127.950 ;
        RECT 151.950 121.950 154.050 124.050 ;
        RECT 146.400 108.000 150.450 108.450 ;
        RECT 146.400 107.400 151.050 108.000 ;
        RECT 130.950 103.950 136.050 106.050 ;
        RECT 139.950 103.950 142.050 106.050 ;
        RECT 148.950 103.950 151.050 107.400 ;
        RECT 124.950 100.950 127.050 103.050 ;
        RECT 92.400 95.400 97.050 97.050 ;
        RECT 93.000 94.950 97.050 95.400 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 100.950 91.950 103.050 97.050 ;
        RECT 106.950 94.950 109.050 97.050 ;
        RECT 109.950 95.400 114.450 97.050 ;
        RECT 109.950 94.950 114.000 95.400 ;
        RECT 115.950 94.950 118.050 100.050 ;
        RECT 121.950 97.950 124.050 100.050 ;
        RECT 67.950 82.950 70.050 85.050 ;
        RECT 79.950 82.950 82.050 85.050 ;
        RECT 80.400 79.050 81.450 82.950 ;
        RECT 79.950 76.950 82.050 79.050 ;
        RECT 40.950 73.950 43.050 76.050 ;
        RECT 76.950 73.950 79.050 76.050 ;
        RECT 28.950 69.300 31.050 71.400 ;
        RECT 43.950 69.300 46.050 71.400 ;
        RECT 28.950 65.700 30.150 69.300 ;
        RECT 44.850 65.700 46.050 69.300 ;
        RECT 64.950 68.400 67.050 70.500 ;
        RECT 28.950 63.600 31.050 65.700 ;
        RECT 43.950 63.600 46.050 65.700 ;
        RECT 13.950 52.950 16.050 55.050 ;
        RECT 19.950 52.950 22.050 58.050 ;
        RECT 7.950 46.500 10.050 48.600 ;
        RECT 14.400 46.050 15.450 52.950 ;
        RECT 16.950 49.950 19.050 52.050 ;
        RECT 13.950 43.950 16.050 46.050 ;
        RECT 17.400 28.050 18.450 49.950 ;
        RECT 28.950 48.600 30.150 63.600 ;
        RECT 31.950 49.950 34.050 55.050 ;
        RECT 39.000 54.450 43.050 55.050 ;
        RECT 38.400 52.950 43.050 54.450 ;
        RECT 28.950 46.500 31.050 48.600 ;
        RECT 19.950 43.950 22.050 46.050 ;
        RECT 20.400 31.050 21.450 43.950 ;
        RECT 38.400 43.050 39.450 52.950 ;
        RECT 44.850 48.600 46.050 63.600 ;
        RECT 49.950 55.950 55.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 59.400 52.050 60.450 55.950 ;
        RECT 58.950 49.950 61.050 52.050 ;
        RECT 65.100 48.600 66.300 68.400 ;
        RECT 43.950 46.500 46.050 48.600 ;
        RECT 64.950 46.500 67.050 48.600 ;
        RECT 37.950 40.950 40.050 43.050 ;
        RECT 43.950 40.950 46.050 43.050 ;
        RECT 61.950 40.950 64.050 43.050 ;
        RECT 19.950 28.950 22.050 31.050 ;
        RECT 10.950 25.950 16.050 28.050 ;
        RECT 16.950 22.950 19.050 28.050 ;
        RECT 20.400 22.050 21.450 28.950 ;
        RECT 37.950 25.950 40.050 31.050 ;
        RECT 44.400 28.050 45.450 40.950 ;
        RECT 49.950 28.950 52.050 31.050 ;
        RECT 58.950 28.950 61.050 31.050 ;
        RECT 43.950 25.950 46.050 28.050 ;
        RECT 7.950 19.950 13.050 22.050 ;
        RECT 19.950 19.950 22.050 22.050 ;
        RECT 34.950 19.950 37.050 25.050 ;
        RECT 44.400 22.050 45.450 25.950 ;
        RECT 50.400 25.050 51.450 28.950 ;
        RECT 49.950 22.950 52.050 25.050 ;
        RECT 40.950 16.950 43.050 22.050 ;
        RECT 43.950 19.950 46.050 22.050 ;
        RECT 59.400 13.050 60.450 28.950 ;
        RECT 62.400 22.050 63.450 40.950 ;
        RECT 77.400 31.050 78.450 73.950 ;
        RECT 80.400 55.050 81.450 76.950 ;
        RECT 100.950 68.400 103.050 70.500 ;
        RECT 82.950 58.950 85.050 61.050 ;
        RECT 88.950 58.950 91.050 61.050 ;
        RECT 79.950 52.950 82.050 55.050 ;
        RECT 83.400 43.050 84.450 58.950 ;
        RECT 85.950 49.950 88.050 55.050 ;
        RECT 82.950 40.950 85.050 43.050 ;
        RECT 89.400 40.050 90.450 58.950 ;
        RECT 101.700 48.600 102.900 68.400 ;
        RECT 107.400 61.050 108.450 94.950 ;
        RECT 125.400 82.050 126.450 100.950 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 136.950 97.950 139.050 103.050 ;
        RECT 131.400 94.050 132.450 97.950 ;
        RECT 130.950 91.950 133.050 94.050 ;
        RECT 136.950 91.950 139.050 94.050 ;
        RECT 140.400 93.450 141.450 103.950 ;
        RECT 142.950 100.950 145.050 103.050 ;
        RECT 143.400 97.050 144.450 100.950 ;
        RECT 152.400 99.450 153.450 121.950 ;
        RECT 158.400 103.050 159.450 130.950 ;
        RECT 149.400 98.400 153.450 99.450 ;
        RECT 142.950 94.950 145.050 97.050 ;
        RECT 140.400 92.400 144.450 93.450 ;
        RECT 124.950 79.950 127.050 82.050 ;
        RECT 112.950 67.950 115.050 70.050 ;
        RECT 121.950 69.300 124.050 71.400 ;
        RECT 106.950 58.950 109.050 61.050 ;
        RECT 113.400 58.050 114.450 67.950 ;
        RECT 121.950 65.700 123.150 69.300 ;
        RECT 121.950 63.600 124.050 65.700 ;
        RECT 112.950 55.950 115.050 58.050 ;
        RECT 121.950 48.600 123.150 63.600 ;
        RECT 130.950 61.950 133.050 64.050 ;
        RECT 131.400 55.050 132.450 61.950 ;
        RECT 137.400 58.050 138.450 91.950 ;
        RECT 143.400 64.050 144.450 92.400 ;
        RECT 142.950 61.950 145.050 64.050 ;
        RECT 136.950 55.950 139.050 58.050 ;
        RECT 124.950 52.950 130.050 55.050 ;
        RECT 130.950 52.950 133.050 55.050 ;
        RECT 143.400 52.050 144.450 61.950 ;
        RECT 149.400 60.450 150.450 98.400 ;
        RECT 157.950 97.950 160.050 103.050 ;
        RECT 161.400 97.050 162.450 133.950 ;
        RECT 185.400 133.050 186.450 169.950 ;
        RECT 188.400 135.450 189.450 178.950 ;
        RECT 200.100 168.600 201.300 188.400 ;
        RECT 214.950 187.950 217.050 190.050 ;
        RECT 211.950 181.950 214.050 187.050 ;
        RECT 218.400 186.450 219.450 196.950 ;
        RECT 220.950 190.950 223.050 193.050 ;
        RECT 215.400 185.400 219.450 186.450 ;
        RECT 215.400 178.050 216.450 185.400 ;
        RECT 221.400 184.050 222.450 190.950 ;
        RECT 217.950 182.400 222.450 184.050 ;
        RECT 217.950 181.950 222.000 182.400 ;
        RECT 233.400 181.050 234.450 202.950 ;
        RECT 226.950 178.950 232.050 181.050 ;
        RECT 232.950 178.950 235.050 181.050 ;
        RECT 214.950 175.950 217.050 178.050 ;
        RECT 220.950 175.950 223.050 178.050 ;
        RECT 221.400 169.050 222.450 175.950 ;
        RECT 199.950 166.500 202.050 168.600 ;
        RECT 220.950 166.950 223.050 169.050 ;
        RECT 190.950 136.950 193.050 142.050 ;
        RECT 188.400 134.400 192.450 135.450 ;
        RECT 178.950 130.950 181.050 133.050 ;
        RECT 185.400 131.400 190.050 133.050 ;
        RECT 186.000 130.950 190.050 131.400 ;
        RECT 179.400 123.450 180.450 130.950 ;
        RECT 176.400 122.400 180.450 123.450 ;
        RECT 172.950 109.950 175.050 112.050 ;
        RECT 173.400 103.200 174.450 109.950 ;
        RECT 176.400 109.050 177.450 122.400 ;
        RECT 181.950 110.400 184.050 112.500 ;
        RECT 176.400 107.400 181.050 109.050 ;
        RECT 177.000 106.950 181.050 107.400 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 172.950 101.100 175.050 103.200 ;
        RECT 167.400 97.050 168.450 100.950 ;
        RECT 160.950 94.950 163.050 97.050 ;
        RECT 166.950 94.950 169.050 97.050 ;
        RECT 172.950 94.950 175.050 99.900 ;
        RECT 182.850 95.400 184.050 110.400 ;
        RECT 191.400 103.050 192.450 134.400 ;
        RECT 196.950 133.950 199.050 139.050 ;
        RECT 211.950 136.950 214.050 142.050 ;
        RECT 233.400 139.050 234.450 178.950 ;
        RECT 217.950 136.950 223.050 139.050 ;
        RECT 223.950 136.950 226.050 139.050 ;
        RECT 232.950 136.950 235.050 139.050 ;
        RECT 193.950 132.450 198.000 133.050 ;
        RECT 193.950 130.950 198.450 132.450 ;
        RECT 214.950 130.950 217.050 133.050 ;
        RECT 197.400 103.050 198.450 130.950 ;
        RECT 202.950 110.400 205.050 112.500 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 181.950 93.300 184.050 95.400 ;
        RECT 182.850 89.700 184.050 93.300 ;
        RECT 181.950 87.600 184.050 89.700 ;
        RECT 154.950 79.950 157.050 82.050 ;
        RECT 155.400 61.050 156.450 79.950 ;
        RECT 166.950 76.950 169.050 79.050 ;
        RECT 163.950 61.050 166.050 61.200 ;
        RECT 146.400 59.400 150.450 60.450 ;
        RECT 142.950 49.950 145.050 52.050 ;
        RECT 100.950 46.500 103.050 48.600 ;
        RECT 121.950 46.500 124.050 48.600 ;
        RECT 146.400 46.050 147.450 59.400 ;
        RECT 154.950 58.950 157.050 61.050 ;
        RECT 160.950 59.100 166.050 61.050 ;
        RECT 160.950 58.950 165.000 59.100 ;
        RECT 151.950 49.950 154.050 55.050 ;
        RECT 163.950 52.950 166.050 57.900 ;
        RECT 127.950 43.950 130.050 46.050 ;
        RECT 145.950 43.950 148.050 46.050 ;
        RECT 88.950 37.950 91.050 40.050 ;
        RECT 76.950 28.950 79.050 31.050 ;
        RECT 118.950 28.950 121.050 31.050 ;
        RECT 64.950 25.950 70.050 28.050 ;
        RECT 61.950 16.950 64.050 22.050 ;
        RECT 70.950 19.950 73.050 25.050 ;
        RECT 77.400 22.050 78.450 28.950 ;
        RECT 82.950 25.950 85.050 28.050 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 71.400 13.050 72.450 19.950 ;
        RECT 83.400 13.050 84.450 25.950 ;
        RECT 88.950 22.950 91.050 28.050 ;
        RECT 106.950 25.950 112.050 28.050 ;
        RECT 112.950 25.950 118.050 28.050 ;
        RECT 119.400 22.050 120.450 28.950 ;
        RECT 128.400 28.050 129.450 43.950 ;
        RECT 127.950 25.950 130.050 28.050 ;
        RECT 133.950 25.950 136.050 31.050 ;
        RECT 100.950 16.950 103.050 22.050 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 118.950 19.950 121.050 22.050 ;
        RECT 113.400 16.050 114.450 19.950 ;
        RECT 124.950 16.950 127.050 22.050 ;
        RECT 142.950 19.950 145.050 25.050 ;
        RECT 151.950 22.950 157.050 25.050 ;
        RECT 167.400 22.200 168.450 76.950 ;
        RECT 191.400 76.050 192.450 100.950 ;
        RECT 203.100 90.600 204.300 110.400 ;
        RECT 215.400 109.050 216.450 130.950 ;
        RECT 214.950 106.950 217.050 109.050 ;
        RECT 218.400 103.050 219.450 136.950 ;
        RECT 224.400 133.050 225.450 136.950 ;
        RECT 236.400 133.050 237.450 211.950 ;
        RECT 242.400 201.450 243.450 214.950 ;
        RECT 242.400 200.400 246.450 201.450 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 242.400 142.050 243.450 160.950 ;
        RECT 245.400 145.050 246.450 200.400 ;
        RECT 244.950 142.950 247.050 145.050 ;
        RECT 251.400 142.050 252.450 250.950 ;
        RECT 255.000 222.450 259.050 223.050 ;
        RECT 254.400 220.950 259.050 222.450 ;
        RECT 254.400 202.050 255.450 220.950 ;
        RECT 263.400 220.200 264.450 253.950 ;
        RECT 284.400 244.050 285.450 253.950 ;
        RECT 283.950 241.950 286.050 244.050 ;
        RECT 287.400 238.050 288.450 262.950 ;
        RECT 293.400 262.050 294.450 283.950 ;
        RECT 298.950 274.950 301.050 277.050 ;
        RECT 292.950 259.950 295.050 262.050 ;
        RECT 293.400 256.050 294.450 259.950 ;
        RECT 299.400 259.050 300.450 274.950 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 292.950 253.950 295.050 256.050 ;
        RECT 305.400 253.050 306.450 328.950 ;
        RECT 311.100 324.600 312.300 344.400 ;
        RECT 326.400 334.050 327.450 349.950 ;
        RECT 349.950 346.950 352.050 349.050 ;
        RECT 328.950 337.950 334.050 340.050 ;
        RECT 337.950 337.950 343.050 340.050 ;
        RECT 343.950 337.950 346.050 343.050 ;
        RECT 350.400 340.050 351.450 346.950 ;
        RECT 349.950 337.950 352.050 340.050 ;
        RECT 326.400 332.400 331.050 334.050 ;
        RECT 327.000 331.950 331.050 332.400 ;
        RECT 334.950 331.950 337.050 337.050 ;
        RECT 344.400 331.050 345.450 337.950 ;
        RECT 343.950 328.950 346.050 331.050 ;
        RECT 310.950 322.500 313.050 324.600 ;
        RECT 353.400 313.050 354.450 370.950 ;
        RECT 361.950 349.950 364.050 352.050 ;
        RECT 355.950 343.950 358.050 346.050 ;
        RECT 356.400 337.050 357.450 343.950 ;
        RECT 362.400 337.050 363.450 349.950 ;
        RECT 368.400 346.050 369.450 394.950 ;
        RECT 367.950 343.950 370.050 346.050 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 361.950 334.950 364.050 337.050 ;
        RECT 367.950 334.950 370.050 337.050 ;
        RECT 371.400 336.450 372.450 463.950 ;
        RECT 380.400 451.050 381.450 497.400 ;
        RECT 386.400 496.050 387.450 514.950 ;
        RECT 392.400 505.050 393.450 568.950 ;
        RECT 399.000 567.900 403.050 568.050 ;
        RECT 397.950 565.950 403.050 567.900 ;
        RECT 406.950 565.950 409.050 571.050 ;
        RECT 397.950 565.800 400.050 565.950 ;
        RECT 416.400 565.050 417.450 571.950 ;
        RECT 424.950 568.950 427.050 574.050 ;
        RECT 428.400 567.450 429.450 601.800 ;
        RECT 431.400 589.050 432.450 607.950 ;
        RECT 434.400 604.050 435.450 637.950 ;
        RECT 440.400 615.450 441.450 637.950 ;
        RECT 440.400 614.400 444.450 615.450 ;
        RECT 439.950 607.950 442.050 610.050 ;
        RECT 440.400 604.050 441.450 607.950 ;
        RECT 433.950 601.950 436.050 604.050 ;
        RECT 439.950 601.950 442.050 604.050 ;
        RECT 443.400 601.050 444.450 614.400 ;
        RECT 449.400 601.050 450.450 637.950 ;
        RECT 464.400 631.050 465.450 646.800 ;
        RECT 491.400 646.050 492.450 664.950 ;
        RECT 497.400 652.050 498.450 676.950 ;
        RECT 512.400 661.050 513.450 676.950 ;
        RECT 517.950 670.950 520.050 673.050 ;
        RECT 499.950 660.450 504.000 661.050 ;
        RECT 499.950 660.000 504.450 660.450 ;
        RECT 499.950 658.950 505.050 660.000 ;
        RECT 511.950 658.950 514.050 661.050 ;
        RECT 502.950 655.950 505.050 658.950 ;
        RECT 493.950 650.400 498.450 652.050 ;
        RECT 493.950 649.950 498.000 650.400 ;
        RECT 499.950 649.950 502.050 655.050 ;
        RECT 514.950 649.950 517.050 655.050 ;
        RECT 490.950 643.950 493.050 646.050 ;
        RECT 508.950 643.950 511.050 649.050 ;
        RECT 518.400 648.450 519.450 670.950 ;
        RECT 521.400 652.050 522.450 679.950 ;
        RECT 530.400 679.050 531.450 740.400 ;
        RECT 533.400 682.050 534.450 757.950 ;
        RECT 545.400 754.050 546.450 772.950 ;
        RECT 547.950 763.950 550.050 766.050 ;
        RECT 552.000 765.450 556.050 766.050 ;
        RECT 551.400 763.950 556.050 765.450 ;
        RECT 544.950 751.950 547.050 754.050 ;
        RECT 548.400 739.200 549.450 763.950 ;
        RECT 551.400 742.050 552.450 763.950 ;
        RECT 556.950 754.950 559.050 760.050 ;
        RECT 556.950 747.450 559.050 751.050 ;
        RECT 554.400 747.000 559.050 747.450 ;
        RECT 554.400 746.400 558.450 747.000 ;
        RECT 550.950 739.950 553.050 742.050 ;
        RECT 547.950 737.100 550.050 739.200 ;
        RECT 554.400 736.050 555.450 746.400 ;
        RECT 560.400 745.050 561.450 778.950 ;
        RECT 566.400 775.050 567.450 781.950 ;
        RECT 565.950 772.950 568.050 775.050 ;
        RECT 568.950 769.950 571.050 772.050 ;
        RECT 562.950 760.050 565.050 766.050 ;
        RECT 569.400 763.050 570.450 769.950 ;
        RECT 571.950 766.950 574.050 769.050 ;
        RECT 568.950 760.950 571.050 763.050 ;
        RECT 562.800 759.000 565.050 760.050 ;
        RECT 566.100 759.000 568.200 760.050 ;
        RECT 562.800 757.950 564.900 759.000 ;
        RECT 565.950 757.950 568.200 759.000 ;
        RECT 565.950 754.950 568.050 757.950 ;
        RECT 572.400 757.050 573.450 766.950 ;
        RECT 578.400 759.450 579.450 802.950 ;
        RECT 580.950 796.950 583.050 802.050 ;
        RECT 587.400 799.050 588.450 811.950 ;
        RECT 592.950 805.950 595.050 808.050 ;
        RECT 601.950 805.950 604.050 808.050 ;
        RECT 613.950 805.950 619.050 808.050 ;
        RECT 622.950 805.950 625.050 811.050 ;
        RECT 704.400 808.050 705.450 811.950 ;
        RECT 721.950 808.950 724.050 811.950 ;
        RECT 725.400 810.450 726.450 815.400 ;
        RECT 745.950 814.950 748.050 817.050 ;
        RECT 739.950 811.950 742.050 814.050 ;
        RECT 725.400 809.400 735.450 810.450 ;
        RECT 734.400 808.050 735.450 809.400 ;
        RECT 740.400 808.050 741.450 811.950 ;
        RECT 586.950 796.950 589.050 799.050 ;
        RECT 593.400 793.050 594.450 805.950 ;
        RECT 598.950 802.950 601.050 805.050 ;
        RECT 592.950 790.950 595.050 793.050 ;
        RECT 592.950 781.950 595.050 784.050 ;
        RECT 583.950 775.950 586.050 778.050 ;
        RECT 580.950 769.950 583.050 772.050 ;
        RECT 575.400 758.400 579.450 759.450 ;
        RECT 571.950 754.950 574.050 757.050 ;
        RECT 568.950 751.950 571.050 754.050 ;
        RECT 559.950 742.950 562.050 745.050 ;
        RECT 547.950 733.800 550.050 735.900 ;
        RECT 553.950 733.950 556.050 736.050 ;
        RECT 548.400 730.050 549.450 733.800 ;
        RECT 569.400 730.050 570.450 751.950 ;
        RECT 575.400 732.450 576.450 758.400 ;
        RECT 577.950 754.950 580.050 757.050 ;
        RECT 578.400 751.050 579.450 754.950 ;
        RECT 577.950 750.450 580.050 751.050 ;
        RECT 581.400 750.450 582.450 769.950 ;
        RECT 584.400 766.050 585.450 775.950 ;
        RECT 583.950 763.950 586.050 766.050 ;
        RECT 593.400 763.050 594.450 781.950 ;
        RECT 599.400 778.050 600.450 802.950 ;
        RECT 602.400 802.050 603.450 805.950 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 643.950 802.950 646.050 808.050 ;
        RECT 652.950 805.950 655.050 808.050 ;
        RECT 685.950 805.950 691.050 808.050 ;
        RECT 703.950 805.950 706.050 808.050 ;
        RECT 601.950 799.950 604.050 802.050 ;
        RECT 613.950 799.950 616.050 802.050 ;
        RECT 602.400 784.050 603.450 799.950 ;
        RECT 604.950 793.950 607.050 799.050 ;
        RECT 601.950 781.950 604.050 784.050 ;
        RECT 598.950 775.950 601.050 778.050 ;
        RECT 595.950 769.950 598.050 772.050 ;
        RECT 596.400 763.050 597.450 769.950 ;
        RECT 601.950 763.050 604.050 763.200 ;
        RECT 605.400 763.050 606.450 793.950 ;
        RECT 610.950 781.950 613.050 784.050 ;
        RECT 586.950 757.950 589.050 763.050 ;
        RECT 592.950 760.950 595.050 763.050 ;
        RECT 595.950 760.950 598.050 763.050 ;
        RECT 598.950 761.100 604.050 763.050 ;
        RECT 598.950 760.950 603.000 761.100 ;
        RECT 604.950 760.950 607.050 763.050 ;
        RECT 589.950 754.950 592.050 757.050 ;
        RECT 595.950 754.950 598.050 757.050 ;
        RECT 601.950 754.950 604.050 759.900 ;
        RECT 611.400 757.050 612.450 781.950 ;
        RECT 614.400 778.050 615.450 799.950 ;
        RECT 619.950 796.950 622.050 802.050 ;
        RECT 625.950 796.950 628.050 799.050 ;
        RECT 626.400 781.050 627.450 796.950 ;
        RECT 625.950 778.950 628.050 781.050 ;
        RECT 613.950 775.950 616.050 778.050 ;
        RECT 629.400 769.200 630.450 802.950 ;
        RECT 631.950 796.950 637.050 799.050 ;
        RECT 653.400 796.050 654.450 805.950 ;
        RECT 679.950 800.100 682.050 805.050 ;
        RECT 685.950 799.950 688.050 802.050 ;
        RECT 691.950 799.950 694.050 802.050 ;
        RECT 709.950 799.950 712.050 808.050 ;
        RECT 730.950 805.950 733.050 808.050 ;
        RECT 734.400 806.400 739.050 808.050 ;
        RECT 735.000 805.950 739.050 806.400 ;
        RECT 739.950 805.950 742.050 808.050 ;
        RECT 724.950 802.950 727.050 805.050 ;
        RECT 673.950 796.950 676.050 799.050 ;
        RECT 652.950 793.950 655.050 796.050 ;
        RECT 640.950 772.950 643.050 775.050 ;
        RECT 616.950 766.950 619.050 769.050 ;
        RECT 628.950 767.100 631.050 769.200 ;
        RECT 617.400 757.050 618.450 766.950 ;
        RECT 628.950 763.800 631.050 765.900 ;
        RECT 634.950 763.950 637.050 766.050 ;
        RECT 610.950 754.950 613.050 757.050 ;
        RECT 616.950 754.950 619.050 757.050 ;
        RECT 577.950 749.400 582.450 750.450 ;
        RECT 577.950 748.950 580.050 749.400 ;
        RECT 590.400 745.050 591.450 754.950 ;
        RECT 596.400 745.050 597.450 754.950 ;
        RECT 601.950 748.950 604.050 751.050 ;
        RECT 577.950 742.950 580.050 745.050 ;
        RECT 589.950 742.950 592.050 745.050 ;
        RECT 595.950 742.950 598.050 745.050 ;
        RECT 572.400 731.400 576.450 732.450 ;
        RECT 541.950 726.450 544.050 730.050 ;
        RECT 547.950 727.950 550.050 730.050 ;
        RECT 553.950 727.950 556.050 730.050 ;
        RECT 568.950 727.950 571.050 730.050 ;
        RECT 539.400 725.400 544.050 726.450 ;
        RECT 535.950 721.950 538.050 724.050 ;
        RECT 536.400 718.050 537.450 721.950 ;
        RECT 535.950 715.950 538.050 718.050 ;
        RECT 535.950 703.950 538.050 706.050 ;
        RECT 536.400 682.050 537.450 703.950 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 535.950 679.950 538.050 682.050 ;
        RECT 539.400 679.050 540.450 725.400 ;
        RECT 541.950 724.950 544.050 725.400 ;
        RECT 544.950 718.950 547.050 724.050 ;
        RECT 550.950 718.950 553.050 724.050 ;
        RECT 550.950 706.950 553.050 709.050 ;
        RECT 551.400 703.050 552.450 706.950 ;
        RECT 550.950 700.950 553.050 703.050 ;
        RECT 554.400 700.050 555.450 727.950 ;
        RECT 559.950 724.950 565.050 727.050 ;
        RECT 572.400 724.050 573.450 731.400 ;
        RECT 574.950 727.950 577.050 730.050 ;
        RECT 568.950 722.400 573.450 724.050 ;
        RECT 568.950 721.950 573.000 722.400 ;
        RECT 568.950 720.450 571.050 721.950 ;
        RECT 566.400 719.400 571.050 720.450 ;
        RECT 553.950 697.950 556.050 700.050 ;
        RECT 559.950 697.950 562.050 700.050 ;
        RECT 541.950 688.950 544.050 691.050 ;
        RECT 542.400 685.200 543.450 688.950 ;
        RECT 541.950 683.100 544.050 685.200 ;
        RECT 541.950 679.800 544.050 681.900 ;
        RECT 529.950 676.950 532.050 679.050 ;
        RECT 538.950 676.950 541.050 679.050 ;
        RECT 532.950 673.950 535.050 676.050 ;
        RECT 533.400 667.050 534.450 673.950 ;
        RECT 539.400 673.050 540.450 676.950 ;
        RECT 542.400 676.050 543.450 679.800 ;
        RECT 554.400 679.050 555.450 697.950 ;
        RECT 560.400 688.050 561.450 697.950 ;
        RECT 566.400 691.050 567.450 719.400 ;
        RECT 568.950 718.950 571.050 719.400 ;
        RECT 575.400 700.050 576.450 727.950 ;
        RECT 578.400 718.050 579.450 742.950 ;
        RECT 583.950 739.950 586.050 742.050 ;
        RECT 584.400 730.050 585.450 739.950 ;
        RECT 602.400 730.050 603.450 748.950 ;
        RECT 629.400 745.050 630.450 763.800 ;
        RECT 635.400 751.050 636.450 763.950 ;
        RECT 641.400 760.050 642.450 772.950 ;
        RECT 643.950 763.950 646.050 769.050 ;
        RECT 649.950 763.950 652.050 766.050 ;
        RECT 640.950 757.950 643.050 760.050 ;
        RECT 634.950 748.950 637.050 751.050 ;
        RECT 628.950 742.950 631.050 745.050 ;
        RECT 643.950 742.950 646.050 745.050 ;
        RECT 634.950 736.950 637.050 739.050 ;
        RECT 583.950 727.950 586.050 730.050 ;
        RECT 595.950 724.950 598.050 730.050 ;
        RECT 601.950 727.950 604.050 730.050 ;
        RECT 607.950 727.950 610.050 733.050 ;
        RECT 635.400 730.200 636.450 736.950 ;
        RECT 634.950 728.100 637.050 730.200 ;
        RECT 644.400 727.050 645.450 742.950 ;
        RECT 619.950 724.950 622.050 727.050 ;
        RECT 604.950 721.950 607.050 724.050 ;
        RECT 610.950 721.950 613.050 724.050 ;
        RECT 583.950 718.950 586.050 721.050 ;
        RECT 589.950 718.950 592.050 721.050 ;
        RECT 577.950 715.950 580.050 718.050 ;
        RECT 580.950 712.950 583.050 715.050 ;
        RECT 574.950 697.950 577.050 700.050 ;
        RECT 559.950 685.950 562.050 688.050 ;
        RECT 565.950 685.950 568.050 691.050 ;
        RECT 541.950 673.950 544.050 676.050 ;
        RECT 544.950 675.450 547.050 679.050 ;
        RECT 550.950 677.400 555.450 679.050 ;
        RECT 550.950 676.950 555.000 677.400 ;
        RECT 544.950 675.000 549.450 675.450 ;
        RECT 545.400 674.400 549.450 675.000 ;
        RECT 538.950 670.950 541.050 673.050 ;
        RECT 544.950 670.950 547.050 673.050 ;
        RECT 532.950 664.950 535.050 667.050 ;
        RECT 538.950 664.950 541.050 667.050 ;
        RECT 529.950 658.950 532.050 661.050 ;
        RECT 520.950 649.950 523.050 652.050 ;
        RECT 526.950 649.950 529.050 652.050 ;
        RECT 515.400 647.400 519.450 648.450 ;
        RECT 454.950 628.950 457.050 631.050 ;
        RECT 463.950 628.950 466.050 631.050 ;
        RECT 451.950 604.950 454.050 610.050 ;
        RECT 455.400 603.450 456.450 628.950 ;
        RECT 491.400 622.050 492.450 643.950 ;
        RECT 499.800 628.950 501.900 631.050 ;
        RECT 490.950 619.950 493.050 622.050 ;
        RECT 478.950 610.950 481.050 613.050 ;
        RECT 457.950 604.950 460.050 610.050 ;
        RECT 466.950 607.950 469.050 610.050 ;
        RECT 452.400 602.400 456.450 603.450 ;
        RECT 442.950 598.950 445.050 601.050 ;
        RECT 448.950 598.950 451.050 601.050 ;
        RECT 449.400 595.050 450.450 598.950 ;
        RECT 448.950 592.950 451.050 595.050 ;
        RECT 430.950 586.950 433.050 589.050 ;
        RECT 445.950 586.950 448.050 589.050 ;
        RECT 442.950 580.950 445.050 583.050 ;
        RECT 436.950 574.950 439.050 577.050 ;
        RECT 430.950 571.950 433.050 574.050 ;
        RECT 425.400 567.000 429.450 567.450 ;
        RECT 424.950 566.400 429.450 567.000 ;
        RECT 415.950 562.950 418.050 565.050 ;
        RECT 424.950 559.950 427.050 566.400 ;
        RECT 397.950 536.400 400.050 538.500 ;
        RECT 418.950 537.300 421.050 539.400 ;
        RECT 398.700 516.600 399.900 536.400 ;
        RECT 409.950 532.950 412.050 535.050 ;
        RECT 418.950 533.700 420.150 537.300 ;
        RECT 410.400 526.050 411.450 532.950 ;
        RECT 418.950 531.600 421.050 533.700 ;
        RECT 403.950 520.950 406.050 526.050 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 397.950 514.500 400.050 516.600 ;
        RECT 391.950 502.950 394.050 505.050 ;
        RECT 388.950 499.950 391.050 502.050 ;
        RECT 384.000 495.450 388.050 496.050 ;
        RECT 383.400 493.950 388.050 495.450 ;
        RECT 383.400 481.050 384.450 493.950 ;
        RECT 389.400 490.050 390.450 499.950 ;
        RECT 391.950 490.950 394.050 496.050 ;
        RECT 388.950 487.950 391.050 490.050 ;
        RECT 394.950 487.950 400.050 490.050 ;
        RECT 400.950 487.950 403.050 493.050 ;
        RECT 382.950 478.950 385.050 481.050 ;
        RECT 379.950 448.950 382.050 451.050 ;
        RECT 376.950 445.950 379.050 448.050 ;
        RECT 373.950 442.950 376.050 445.050 ;
        RECT 374.400 415.050 375.450 442.950 ;
        RECT 377.400 442.050 378.450 445.950 ;
        RECT 383.400 445.050 384.450 478.950 ;
        RECT 403.950 475.950 406.050 478.050 ;
        RECT 404.400 466.050 405.450 475.950 ;
        RECT 403.950 463.950 406.050 466.050 ;
        RECT 394.950 458.400 397.050 460.500 ;
        RECT 382.950 442.950 385.050 445.050 ;
        RECT 376.950 439.950 379.050 442.050 ;
        RECT 395.700 438.600 396.900 458.400 ;
        RECT 400.950 448.950 403.050 454.050 ;
        RECT 410.400 448.050 411.450 523.950 ;
        RECT 418.950 516.600 420.150 531.600 ;
        RECT 425.400 523.050 426.450 559.950 ;
        RECT 431.400 550.050 432.450 571.950 ;
        RECT 437.400 571.050 438.450 574.950 ;
        RECT 443.400 571.050 444.450 580.950 ;
        RECT 446.400 574.050 447.450 586.950 ;
        RECT 445.950 571.950 448.050 574.050 ;
        RECT 436.950 565.950 439.050 571.050 ;
        RECT 442.950 565.950 445.050 571.050 ;
        RECT 431.400 548.400 436.050 550.050 ;
        RECT 432.000 547.950 436.050 548.400 ;
        RECT 439.950 526.950 442.050 532.050 ;
        RECT 421.950 521.400 426.450 523.050 ;
        RECT 421.950 520.950 426.000 521.400 ;
        RECT 418.950 514.500 421.050 516.600 ;
        RECT 421.950 508.950 424.050 511.050 ;
        RECT 422.400 487.050 423.450 508.950 ;
        RECT 430.950 490.950 436.050 493.050 ;
        RECT 412.950 481.950 415.050 487.050 ;
        RECT 421.950 484.950 424.050 487.050 ;
        RECT 415.950 459.300 418.050 461.400 ;
        RECT 415.950 455.700 417.150 459.300 ;
        RECT 415.950 453.600 418.050 455.700 ;
        RECT 406.950 442.950 409.050 448.050 ;
        RECT 409.950 445.950 412.050 448.050 ;
        RECT 415.950 438.600 417.150 453.600 ;
        RECT 422.400 445.050 423.450 484.950 ;
        RECT 427.950 481.950 430.050 487.050 ;
        RECT 440.400 486.450 441.450 526.950 ;
        RECT 448.950 487.950 451.050 493.050 ;
        RECT 442.950 486.450 445.050 487.050 ;
        RECT 440.400 485.400 445.050 486.450 ;
        RECT 442.950 484.950 445.050 485.400 ;
        RECT 436.950 481.800 439.050 483.900 ;
        RECT 424.950 457.950 427.050 460.050 ;
        RECT 418.950 443.400 423.450 445.050 ;
        RECT 418.950 442.950 423.000 443.400 ;
        RECT 394.950 436.500 397.050 438.600 ;
        RECT 415.950 436.500 418.050 438.600 ;
        RECT 382.950 433.950 385.050 436.050 ;
        RECT 383.400 421.050 384.450 433.950 ;
        RECT 382.950 418.950 385.050 421.050 ;
        RECT 373.950 409.950 376.050 415.050 ;
        RECT 412.950 406.950 415.050 409.050 ;
        RECT 413.400 403.050 414.450 406.950 ;
        RECT 425.400 403.050 426.450 457.950 ;
        RECT 429.000 447.450 433.050 448.050 ;
        RECT 428.400 445.950 433.050 447.450 ;
        RECT 428.400 442.050 429.450 445.950 ;
        RECT 437.400 445.050 438.450 481.800 ;
        RECT 443.400 460.050 444.450 484.950 ;
        RECT 452.400 475.050 453.450 602.400 ;
        RECT 454.950 595.950 457.050 601.050 ;
        RECT 460.950 599.100 463.050 604.050 ;
        RECT 460.950 595.800 463.050 597.900 ;
        RECT 457.950 586.950 460.050 589.050 ;
        RECT 458.400 574.050 459.450 586.950 ;
        RECT 457.950 571.950 460.050 574.050 ;
        RECT 458.400 531.450 459.450 571.950 ;
        RECT 461.400 568.050 462.450 595.800 ;
        RECT 467.400 595.050 468.450 607.950 ;
        RECT 479.400 598.050 480.450 610.950 ;
        RECT 500.400 610.050 501.450 628.950 ;
        RECT 499.950 607.950 502.050 610.050 ;
        RECT 481.950 598.950 484.050 604.050 ;
        RECT 487.950 601.950 490.050 604.050 ;
        RECT 478.950 595.950 481.050 598.050 ;
        RECT 488.400 595.050 489.450 601.950 ;
        RECT 500.400 601.050 501.450 607.950 ;
        RECT 515.400 607.200 516.450 647.400 ;
        RECT 527.400 646.050 528.450 649.950 ;
        RECT 517.950 643.950 520.050 646.050 ;
        RECT 518.400 637.050 519.450 643.950 ;
        RECT 523.950 640.950 526.050 646.050 ;
        RECT 526.950 643.950 529.050 646.050 ;
        RECT 527.400 640.050 528.450 643.950 ;
        RECT 526.950 637.950 529.050 640.050 ;
        RECT 517.950 634.950 520.050 637.050 ;
        RECT 523.950 619.950 526.050 622.050 ;
        RECT 517.950 613.950 520.050 616.050 ;
        RECT 502.950 603.450 505.050 604.050 ;
        RECT 508.950 603.450 511.050 607.050 ;
        RECT 514.950 605.100 517.050 607.200 ;
        RECT 502.950 603.000 511.050 603.450 ;
        RECT 502.950 602.400 510.450 603.000 ;
        RECT 502.950 601.950 505.050 602.400 ;
        RECT 514.950 601.800 517.050 603.900 ;
        RECT 499.950 598.950 502.050 601.050 ;
        RECT 505.950 598.950 508.050 601.050 ;
        RECT 502.950 595.950 505.050 598.050 ;
        RECT 466.950 592.950 469.050 595.050 ;
        RECT 487.950 592.950 490.050 595.050 ;
        RECT 472.950 589.950 475.050 592.050 ;
        RECT 490.950 589.950 493.050 592.050 ;
        RECT 473.400 583.050 474.450 589.950 ;
        RECT 475.950 583.950 478.050 586.050 ;
        RECT 472.950 580.950 475.050 583.050 ;
        RECT 476.400 574.050 477.450 583.950 ;
        RECT 481.950 580.950 484.050 583.050 ;
        RECT 475.950 571.950 478.050 574.050 ;
        RECT 482.400 571.050 483.450 580.950 ;
        RECT 484.950 571.950 490.050 574.050 ;
        RECT 481.950 568.950 484.050 571.050 ;
        RECT 460.950 565.950 463.050 568.050 ;
        RECT 463.950 565.950 466.050 568.050 ;
        RECT 458.400 530.400 462.450 531.450 ;
        RECT 454.950 529.050 457.050 529.200 ;
        RECT 454.950 527.100 460.050 529.050 ;
        RECT 456.000 526.950 460.050 527.100 ;
        RECT 454.950 520.950 457.050 525.900 ;
        RECT 461.400 523.050 462.450 530.400 ;
        RECT 464.400 523.050 465.450 565.950 ;
        RECT 478.950 559.950 481.050 565.050 ;
        RECT 479.400 553.050 480.450 559.950 ;
        RECT 478.950 550.950 481.050 553.050 ;
        RECT 485.400 549.450 486.450 571.950 ;
        RECT 491.400 568.050 492.450 589.950 ;
        RECT 503.400 586.050 504.450 595.950 ;
        RECT 502.950 583.950 505.050 586.050 ;
        RECT 506.400 574.050 507.450 598.950 ;
        RECT 515.400 598.050 516.450 601.800 ;
        RECT 508.950 595.950 511.050 598.050 ;
        RECT 514.950 595.950 517.050 598.050 ;
        RECT 509.400 586.050 510.450 595.950 ;
        RECT 518.400 589.050 519.450 613.950 ;
        RECT 524.400 607.050 525.450 619.950 ;
        RECT 530.400 616.050 531.450 658.950 ;
        RECT 532.950 643.950 538.050 646.050 ;
        RECT 532.950 634.950 535.050 637.050 ;
        RECT 533.400 622.050 534.450 634.950 ;
        RECT 535.950 622.950 538.050 625.050 ;
        RECT 532.950 619.950 535.050 622.050 ;
        RECT 529.950 613.950 532.050 616.050 ;
        RECT 536.400 607.050 537.450 622.950 ;
        RECT 539.400 607.200 540.450 664.950 ;
        RECT 541.950 646.950 544.050 649.050 ;
        RECT 542.400 643.050 543.450 646.950 ;
        RECT 545.400 646.050 546.450 670.950 ;
        RECT 548.400 667.050 549.450 674.400 ;
        RECT 553.950 667.950 556.050 670.050 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 554.400 661.050 555.450 667.950 ;
        RECT 553.950 658.950 556.050 661.050 ;
        RECT 547.950 652.950 550.050 655.050 ;
        RECT 548.400 646.050 549.450 652.950 ;
        RECT 550.950 649.950 556.050 652.050 ;
        RECT 560.400 648.450 561.450 685.950 ;
        RECT 571.950 676.950 574.050 682.050 ;
        RECT 581.400 679.050 582.450 712.950 ;
        RECT 584.400 688.050 585.450 718.950 ;
        RECT 590.400 706.050 591.450 718.950 ;
        RECT 605.400 715.050 606.450 721.950 ;
        RECT 604.950 712.950 607.050 715.050 ;
        RECT 589.950 703.950 592.050 706.050 ;
        RECT 586.950 688.950 589.050 691.050 ;
        RECT 598.950 688.950 601.050 691.050 ;
        RECT 583.950 685.950 586.050 688.050 ;
        RECT 587.400 685.050 588.450 688.950 ;
        RECT 599.400 685.050 600.450 688.950 ;
        RECT 611.400 685.050 612.450 721.950 ;
        RECT 620.400 706.050 621.450 724.950 ;
        RECT 634.950 724.800 637.050 726.900 ;
        RECT 643.950 724.950 646.050 727.050 ;
        RECT 625.950 718.950 628.050 724.050 ;
        RECT 635.400 715.050 636.450 724.800 ;
        RECT 640.950 721.950 643.050 724.050 ;
        RECT 634.950 712.950 637.050 715.050 ;
        RECT 619.950 703.950 622.050 706.050 ;
        RECT 634.950 700.950 637.050 703.050 ;
        RECT 622.950 697.950 625.050 700.050 ;
        RECT 586.950 682.950 589.050 685.050 ;
        RECT 592.950 682.950 595.050 685.050 ;
        RECT 598.950 682.950 601.050 685.050 ;
        RECT 604.950 682.950 607.050 685.050 ;
        RECT 610.950 682.950 613.050 685.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 580.950 676.950 583.050 679.050 ;
        RECT 565.950 676.050 568.050 676.200 ;
        RECT 568.950 676.050 571.050 676.200 ;
        RECT 565.950 674.100 571.050 676.050 ;
        RECT 567.000 673.950 570.000 674.100 ;
        RECT 574.950 673.950 577.050 676.050 ;
        RECT 568.950 670.800 571.050 672.900 ;
        RECT 569.400 658.050 570.450 670.800 ;
        RECT 571.950 658.950 574.050 661.050 ;
        RECT 568.950 655.950 571.050 658.050 ;
        RECT 572.400 652.050 573.450 658.950 ;
        RECT 575.400 658.050 576.450 673.950 ;
        RECT 581.400 667.050 582.450 676.950 ;
        RECT 580.950 664.950 583.050 667.050 ;
        RECT 574.950 655.950 577.050 658.050 ;
        RECT 568.950 649.950 571.050 652.050 ;
        RECT 571.950 649.950 574.050 652.050 ;
        RECT 560.400 647.400 564.450 648.450 ;
        RECT 544.950 643.950 547.050 646.050 ;
        RECT 548.400 644.400 553.050 646.050 ;
        RECT 549.000 643.950 553.050 644.400 ;
        RECT 556.950 643.950 559.050 646.050 ;
        RECT 541.950 640.950 544.050 643.050 ;
        RECT 550.950 640.950 553.050 643.950 ;
        RECT 542.400 637.050 543.450 640.950 ;
        RECT 553.950 637.950 556.050 640.050 ;
        RECT 541.950 634.950 544.050 637.050 ;
        RECT 545.400 636.000 552.450 636.450 ;
        RECT 544.950 635.400 552.450 636.000 ;
        RECT 544.950 631.950 547.050 635.400 ;
        RECT 551.400 616.050 552.450 635.400 ;
        RECT 550.950 613.950 553.050 616.050 ;
        RECT 554.400 613.050 555.450 637.950 ;
        RECT 557.400 622.050 558.450 643.950 ;
        RECT 563.400 642.450 564.450 647.400 ;
        RECT 560.400 642.000 564.450 642.450 ;
        RECT 559.950 641.400 564.450 642.000 ;
        RECT 569.400 642.450 570.450 649.950 ;
        RECT 577.950 646.950 583.050 649.050 ;
        RECT 569.400 642.000 573.450 642.450 ;
        RECT 569.400 641.400 574.050 642.000 ;
        RECT 559.950 637.950 562.050 641.400 ;
        RECT 571.950 637.950 574.050 641.400 ;
        RECT 574.950 640.950 577.050 646.050 ;
        RECT 584.400 643.050 585.450 679.950 ;
        RECT 593.400 679.050 594.450 682.950 ;
        RECT 586.950 676.950 592.050 679.050 ;
        RECT 592.950 676.950 595.050 679.050 ;
        RECT 586.950 655.950 589.050 658.050 ;
        RECT 583.950 640.950 586.050 643.050 ;
        RECT 587.400 640.050 588.450 655.950 ;
        RECT 593.400 649.050 594.450 676.950 ;
        RECT 598.950 667.950 601.050 670.050 ;
        RECT 592.950 646.950 595.050 649.050 ;
        RECT 599.400 646.050 600.450 667.950 ;
        RECT 605.400 658.050 606.450 682.950 ;
        RECT 623.400 679.050 624.450 697.950 ;
        RECT 631.950 685.050 634.050 685.200 ;
        RECT 625.950 682.950 628.050 685.050 ;
        RECT 630.000 684.600 634.050 685.050 ;
        RECT 629.400 683.100 634.050 684.600 ;
        RECT 629.400 682.950 633.000 683.100 ;
        RECT 626.400 679.200 627.450 682.950 ;
        RECT 610.950 676.950 613.050 679.050 ;
        RECT 613.950 676.950 619.050 679.050 ;
        RECT 622.950 676.950 625.050 679.050 ;
        RECT 625.950 677.100 628.050 679.200 ;
        RECT 611.400 673.050 612.450 676.950 ;
        RECT 607.800 670.950 609.900 673.050 ;
        RECT 611.100 670.950 613.200 673.050 ;
        RECT 608.400 667.050 609.450 670.950 ;
        RECT 607.950 664.950 610.050 667.050 ;
        RECT 604.950 655.950 607.050 658.050 ;
        RECT 616.950 655.950 619.050 658.050 ;
        RECT 607.950 649.950 610.050 652.050 ;
        RECT 601.950 646.950 604.050 649.050 ;
        RECT 589.950 640.950 592.050 646.050 ;
        RECT 598.950 643.950 601.050 646.050 ;
        RECT 586.950 637.950 589.050 640.050 ;
        RECT 574.950 634.950 577.050 637.050 ;
        RECT 556.950 619.950 559.050 622.050 ;
        RECT 553.950 607.950 556.050 613.050 ;
        RECT 520.950 604.950 523.050 607.050 ;
        RECT 523.950 604.950 526.050 607.050 ;
        RECT 529.950 604.950 532.050 607.050 ;
        RECT 532.950 605.400 537.450 607.050 ;
        RECT 532.950 604.950 537.000 605.400 ;
        RECT 538.950 605.100 541.050 607.200 ;
        RECT 557.400 607.050 558.450 619.950 ;
        RECT 562.950 610.950 565.050 616.050 ;
        RECT 517.950 586.950 520.050 589.050 ;
        RECT 508.950 583.950 511.050 586.050 ;
        RECT 505.950 571.950 508.050 574.050 ;
        RECT 513.000 573.900 516.000 574.050 ;
        RECT 511.950 571.950 517.050 573.900 ;
        RECT 511.950 571.800 514.050 571.950 ;
        RECT 514.950 571.800 517.050 571.950 ;
        RECT 490.950 565.950 493.050 568.050 ;
        RECT 496.950 565.950 502.050 568.050 ;
        RECT 514.950 567.450 517.050 568.050 ;
        RECT 521.400 567.450 522.450 604.950 ;
        RECT 530.400 601.050 531.450 604.950 ;
        RECT 538.950 601.800 541.050 603.900 ;
        RECT 544.950 601.950 547.050 607.050 ;
        RECT 556.950 604.950 559.050 607.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 523.950 598.950 526.050 601.050 ;
        RECT 529.950 598.950 532.050 601.050 ;
        RECT 524.400 574.050 525.450 598.950 ;
        RECT 532.950 595.950 535.050 598.050 ;
        RECT 533.400 583.050 534.450 595.950 ;
        RECT 539.400 586.050 540.450 601.800 ;
        RECT 538.950 583.950 541.050 586.050 ;
        RECT 544.950 583.950 547.050 586.050 ;
        RECT 532.950 580.950 535.050 583.050 ;
        RECT 533.400 574.050 534.450 580.950 ;
        RECT 545.400 574.050 546.450 583.950 ;
        RECT 560.400 583.050 561.450 601.950 ;
        RECT 559.950 580.950 562.050 583.050 ;
        RECT 565.950 577.950 568.050 580.050 ;
        RECT 523.950 571.950 526.050 574.050 ;
        RECT 526.950 571.950 529.050 574.050 ;
        RECT 532.950 571.950 535.050 574.050 ;
        RECT 544.950 571.950 547.050 574.050 ;
        RECT 553.950 571.950 556.050 574.050 ;
        RECT 562.950 571.950 565.050 577.050 ;
        RECT 527.400 568.050 528.450 571.950 ;
        RECT 538.950 568.050 541.050 568.200 ;
        RECT 514.950 566.400 522.450 567.450 ;
        RECT 514.950 565.950 517.050 566.400 ;
        RECT 508.950 562.950 511.050 565.050 ;
        RECT 509.400 559.050 510.450 562.950 ;
        RECT 508.950 556.950 511.050 559.050 ;
        RECT 479.400 548.400 486.450 549.450 ;
        RECT 469.950 536.400 472.050 538.500 ;
        RECT 460.950 520.950 463.050 523.050 ;
        RECT 464.400 521.400 469.050 523.050 ;
        RECT 465.000 520.950 469.050 521.400 ;
        RECT 461.400 514.050 462.450 520.950 ;
        RECT 463.950 514.950 466.050 517.050 ;
        RECT 470.700 516.600 471.900 536.400 ;
        RECT 475.950 523.950 478.050 529.050 ;
        RECT 460.950 511.950 463.050 514.050 ;
        RECT 454.950 502.950 457.050 505.050 ;
        RECT 455.400 487.050 456.450 502.950 ;
        RECT 464.400 493.050 465.450 514.950 ;
        RECT 469.950 514.500 472.050 516.600 ;
        RECT 472.950 508.950 475.050 511.050 ;
        RECT 473.400 496.050 474.450 508.950 ;
        RECT 479.400 502.050 480.450 548.400 ;
        RECT 490.950 537.300 493.050 539.400 ;
        RECT 499.950 538.950 502.050 541.050 ;
        RECT 481.950 532.950 484.050 535.050 ;
        RECT 490.950 533.700 492.150 537.300 ;
        RECT 482.400 526.050 483.450 532.950 ;
        RECT 490.950 531.600 493.050 533.700 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 490.950 516.600 492.150 531.600 ;
        RECT 493.950 520.950 496.050 526.050 ;
        RECT 500.400 523.050 501.450 538.950 ;
        RECT 505.950 536.400 508.050 538.500 ;
        RECT 502.950 532.950 505.050 535.050 ;
        RECT 503.400 526.050 504.450 532.950 ;
        RECT 502.950 523.950 505.050 526.050 ;
        RECT 499.950 520.950 502.050 523.050 ;
        RECT 506.700 516.600 507.900 536.400 ;
        RECT 511.950 523.950 514.050 526.050 ;
        RECT 514.950 523.950 520.050 526.050 ;
        RECT 490.950 514.500 493.050 516.600 ;
        RECT 505.950 514.500 508.050 516.600 ;
        RECT 499.950 511.950 502.050 514.050 ;
        RECT 478.950 499.950 481.050 502.050 ;
        RECT 500.400 501.450 501.450 511.950 ;
        RECT 512.400 508.050 513.450 523.950 ;
        RECT 521.400 523.050 522.450 566.400 ;
        RECT 523.950 565.950 526.050 568.050 ;
        RECT 526.950 565.950 529.050 568.050 ;
        RECT 524.400 550.050 525.450 565.950 ;
        RECT 529.950 562.950 532.050 568.050 ;
        RECT 538.950 566.100 544.050 568.050 ;
        RECT 540.000 565.950 544.050 566.100 ;
        RECT 538.950 562.800 541.050 564.900 ;
        RECT 523.950 547.950 526.050 550.050 ;
        RECT 526.950 537.300 529.050 539.400 ;
        RECT 526.950 533.700 528.150 537.300 ;
        RECT 526.950 531.600 529.050 533.700 ;
        RECT 520.950 520.950 523.050 523.050 ;
        RECT 517.950 514.950 520.050 517.050 ;
        RECT 526.950 516.600 528.150 531.600 ;
        RECT 532.950 526.950 535.050 529.050 ;
        RECT 529.950 520.950 532.050 526.050 ;
        RECT 511.950 505.950 514.050 508.050 ;
        RECT 514.950 502.950 517.050 505.050 ;
        RECT 497.400 500.400 501.450 501.450 ;
        RECT 479.400 496.050 480.450 499.950 ;
        RECT 472.950 493.950 475.050 496.050 ;
        RECT 478.950 493.950 481.050 496.050 ;
        RECT 493.950 493.950 496.050 496.050 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 466.950 487.950 472.050 490.050 ;
        RECT 454.950 484.950 457.050 487.050 ;
        RECT 460.950 484.950 463.050 487.050 ;
        RECT 475.950 484.950 478.050 490.050 ;
        RECT 490.950 487.950 493.050 493.050 ;
        RECT 494.400 486.450 495.450 493.950 ;
        RECT 497.400 490.050 498.450 500.400 ;
        RECT 515.400 496.050 516.450 502.950 ;
        RECT 499.950 493.950 505.050 496.050 ;
        RECT 508.950 493.950 511.050 496.050 ;
        RECT 514.950 493.950 517.050 496.050 ;
        RECT 496.950 487.950 499.050 490.050 ;
        RECT 494.400 485.400 498.450 486.450 ;
        RECT 461.400 481.050 462.450 484.950 ;
        RECT 460.950 478.950 463.050 481.050 ;
        RECT 493.950 478.950 496.050 481.050 ;
        RECT 451.950 472.950 454.050 475.050 ;
        RECT 475.950 472.950 478.050 475.050 ;
        RECT 442.950 457.950 445.050 460.050 ;
        RECT 448.950 458.400 451.050 460.500 ;
        RECT 469.950 459.300 472.050 461.400 ;
        RECT 439.950 448.950 442.050 451.050 ;
        RECT 436.950 442.950 439.050 445.050 ;
        RECT 427.950 439.950 430.050 442.050 ;
        RECT 406.950 400.950 409.050 403.050 ;
        RECT 412.950 400.950 415.050 403.050 ;
        RECT 424.950 400.950 427.050 403.050 ;
        RECT 391.950 380.400 394.050 382.500 ;
        RECT 379.950 373.950 382.050 376.050 ;
        RECT 380.400 370.050 381.450 373.950 ;
        RECT 379.950 367.950 385.050 370.050 ;
        RECT 383.400 352.050 384.450 367.950 ;
        RECT 385.950 364.950 388.050 367.050 ;
        RECT 382.950 349.950 385.050 352.050 ;
        RECT 379.950 344.400 382.050 346.500 ;
        RECT 371.400 335.400 375.450 336.450 ;
        RECT 368.400 331.050 369.450 334.950 ;
        RECT 358.950 328.950 364.050 331.050 ;
        RECT 367.950 328.950 370.050 331.050 ;
        RECT 352.950 310.950 355.050 313.050 ;
        RECT 368.400 310.050 369.450 328.950 ;
        RECT 374.400 325.050 375.450 335.400 ;
        RECT 376.950 334.950 379.050 340.050 ;
        RECT 380.850 329.400 382.050 344.400 ;
        RECT 379.950 327.300 382.050 329.400 ;
        RECT 373.950 322.950 376.050 325.050 ;
        RECT 380.850 323.700 382.050 327.300 ;
        RECT 379.950 321.600 382.050 323.700 ;
        RECT 367.950 307.950 370.050 310.050 ;
        RECT 331.950 303.300 334.050 305.400 ;
        RECT 332.850 299.700 334.050 303.300 ;
        RECT 352.950 302.400 355.050 304.500 ;
        RECT 331.950 297.600 334.050 299.700 ;
        RECT 313.950 292.950 316.050 295.050 ;
        RECT 316.950 292.950 322.050 295.050 ;
        RECT 314.400 289.050 315.450 292.950 ;
        RECT 313.950 286.950 316.050 289.050 ;
        RECT 319.950 286.950 325.050 289.050 ;
        RECT 325.950 286.950 331.050 289.050 ;
        RECT 307.950 283.950 310.050 286.050 ;
        RECT 304.950 250.950 307.050 253.050 ;
        RECT 289.950 241.950 292.050 244.050 ;
        RECT 286.950 235.950 289.050 238.050 ;
        RECT 283.950 226.950 286.050 229.050 ;
        RECT 262.950 218.100 265.050 220.200 ;
        RECT 268.950 217.950 271.050 220.050 ;
        RECT 271.950 217.950 274.050 220.050 ;
        RECT 258.000 216.450 262.050 217.050 ;
        RECT 257.400 214.950 262.050 216.450 ;
        RECT 257.400 211.050 258.450 214.950 ;
        RECT 262.950 211.950 265.050 216.900 ;
        RECT 256.950 208.950 259.050 211.050 ;
        RECT 253.950 199.950 256.050 202.050 ;
        RECT 263.400 172.050 264.450 211.950 ;
        RECT 269.400 184.050 270.450 217.950 ;
        RECT 272.400 196.050 273.450 217.950 ;
        RECT 284.400 217.200 285.450 226.950 ;
        RECT 286.950 220.950 289.050 223.050 ;
        RECT 274.950 214.950 280.050 217.050 ;
        RECT 283.950 215.100 286.050 217.200 ;
        RECT 283.950 211.800 286.050 213.900 ;
        RECT 277.950 208.950 283.050 211.050 ;
        RECT 271.950 193.950 274.050 196.050 ;
        RECT 268.950 181.950 271.050 184.050 ;
        RECT 271.950 175.950 274.050 181.050 ;
        RECT 284.400 178.050 285.450 211.800 ;
        RECT 287.400 181.200 288.450 220.950 ;
        RECT 290.400 214.200 291.450 241.950 ;
        RECT 292.950 214.950 295.050 217.050 ;
        RECT 298.950 214.950 304.050 217.050 ;
        RECT 289.950 212.100 292.050 214.200 ;
        RECT 293.400 211.050 294.450 214.950 ;
        RECT 295.950 211.950 298.050 214.050 ;
        RECT 308.400 213.450 309.450 283.950 ;
        RECT 332.850 282.600 334.050 297.600 ;
        RECT 340.950 295.950 343.050 298.050 ;
        RECT 341.400 292.050 342.450 295.950 ;
        RECT 340.950 289.950 343.050 292.050 ;
        RECT 331.950 280.500 334.050 282.600 ;
        RECT 328.950 274.950 331.050 277.050 ;
        RECT 310.950 259.950 313.050 265.050 ;
        RECT 329.400 262.200 330.450 274.950 ;
        RECT 341.400 265.050 342.450 289.950 ;
        RECT 346.950 286.950 349.050 292.050 ;
        RECT 353.100 282.600 354.300 302.400 ;
        RECT 376.950 301.950 379.050 304.050 ;
        RECT 377.400 295.050 378.450 301.950 ;
        RECT 367.950 292.950 373.050 295.050 ;
        RECT 376.950 292.950 379.050 295.050 ;
        RECT 367.950 288.450 372.000 289.050 ;
        RECT 367.950 286.950 372.450 288.450 ;
        RECT 373.950 286.950 379.050 289.050 ;
        RECT 352.950 280.500 355.050 282.600 ;
        RECT 371.400 277.050 372.450 286.950 ;
        RECT 355.950 274.950 358.050 277.050 ;
        RECT 370.950 274.950 373.050 277.050 ;
        RECT 340.950 262.950 343.050 265.050 ;
        RECT 322.950 257.100 325.050 262.050 ;
        RECT 328.950 260.100 331.050 262.200 ;
        RECT 328.950 256.800 331.050 258.900 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 313.950 253.950 316.050 256.050 ;
        RECT 319.950 255.900 324.000 256.050 ;
        RECT 319.950 253.950 325.050 255.900 ;
        RECT 314.400 244.050 315.450 253.950 ;
        RECT 322.950 253.800 325.050 253.950 ;
        RECT 325.950 250.950 328.050 256.050 ;
        RECT 313.950 241.950 316.050 244.050 ;
        RECT 329.400 229.050 330.450 256.800 ;
        RECT 338.400 247.050 339.450 256.950 ;
        RECT 340.950 250.950 346.050 253.050 ;
        RECT 349.950 250.950 352.050 253.050 ;
        RECT 337.950 244.950 340.050 247.050 ;
        RECT 328.950 226.950 331.050 229.050 ;
        RECT 316.950 224.400 319.050 226.500 ;
        RECT 337.950 225.300 340.050 227.400 ;
        RECT 305.400 212.400 309.450 213.450 ;
        RECT 291.000 210.900 294.450 211.050 ;
        RECT 289.950 209.400 294.450 210.900 ;
        RECT 289.950 208.950 294.000 209.400 ;
        RECT 289.950 208.800 292.050 208.950 ;
        RECT 289.950 199.950 292.050 202.050 ;
        RECT 290.400 184.050 291.450 199.950 ;
        RECT 296.400 196.050 297.450 211.950 ;
        RECT 305.400 205.050 306.450 212.400 ;
        RECT 307.950 208.950 310.050 211.050 ;
        RECT 304.950 202.950 307.050 205.050 ;
        RECT 295.950 193.950 298.050 196.050 ;
        RECT 295.950 184.950 298.050 187.050 ;
        RECT 289.950 181.950 292.050 184.050 ;
        RECT 286.950 179.100 289.050 181.200 ;
        RECT 296.400 178.050 297.450 184.950 ;
        RECT 301.950 178.950 304.050 184.050 ;
        RECT 277.950 175.950 283.050 178.050 ;
        RECT 283.950 175.950 286.050 178.050 ;
        RECT 286.950 175.800 289.050 177.900 ;
        RECT 295.950 175.950 298.050 178.050 ;
        RECT 262.950 169.950 265.050 172.050 ;
        RECT 280.950 151.950 283.050 154.050 ;
        RECT 241.950 139.950 244.050 142.050 ;
        RECT 247.950 140.400 252.450 142.050 ;
        RECT 247.950 139.950 252.000 140.400 ;
        RECT 256.950 139.950 259.050 145.050 ;
        RECT 281.400 142.050 282.450 151.950 ;
        RECT 262.950 136.950 265.050 142.050 ;
        RECT 273.000 141.450 277.050 142.050 ;
        RECT 272.400 139.950 277.050 141.450 ;
        RECT 280.950 139.950 283.050 142.050 ;
        RECT 272.400 136.050 273.450 139.950 ;
        RECT 287.400 139.050 288.450 175.800 ;
        RECT 296.400 151.050 297.450 175.950 ;
        RECT 302.400 160.050 303.450 178.950 ;
        RECT 305.400 178.050 306.450 202.950 ;
        RECT 308.400 199.050 309.450 208.950 ;
        RECT 317.700 204.600 318.900 224.400 ;
        RECT 337.950 221.700 339.150 225.300 ;
        RECT 337.950 219.600 340.050 221.700 ;
        RECT 322.950 214.950 328.050 217.050 ;
        RECT 328.950 211.950 331.050 214.050 ;
        RECT 316.950 202.500 319.050 204.600 ;
        RECT 325.950 202.950 328.050 205.050 ;
        RECT 307.950 196.950 310.050 199.050 ;
        RECT 307.950 181.950 310.050 187.050 ;
        RECT 326.400 184.050 327.450 202.950 ;
        RECT 325.950 181.950 328.050 184.050 ;
        RECT 329.400 181.200 330.450 211.950 ;
        RECT 337.950 204.600 339.150 219.600 ;
        RECT 340.950 205.950 343.050 211.050 ;
        RECT 350.400 208.050 351.450 250.950 ;
        RECT 356.400 223.200 357.450 274.950 ;
        RECT 386.400 274.050 387.450 364.950 ;
        RECT 392.700 360.600 393.900 380.400 ;
        RECT 397.950 370.950 400.050 373.050 ;
        RECT 398.400 361.050 399.450 370.950 ;
        RECT 400.950 367.950 406.050 370.050 ;
        RECT 391.950 358.500 394.050 360.600 ;
        RECT 397.950 358.950 400.050 361.050 ;
        RECT 388.950 349.950 391.050 352.050 ;
        RECT 389.400 337.050 390.450 349.950 ;
        RECT 400.950 344.400 403.050 346.500 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 389.400 331.050 390.450 334.950 ;
        RECT 394.950 331.950 397.050 334.050 ;
        RECT 388.950 328.950 391.050 331.050 ;
        RECT 395.400 319.050 396.450 331.950 ;
        RECT 401.100 324.600 402.300 344.400 ;
        RECT 400.950 322.500 403.050 324.600 ;
        RECT 394.950 316.950 397.050 319.050 ;
        RECT 403.950 316.950 406.050 319.050 ;
        RECT 388.950 310.950 391.050 313.050 ;
        RECT 389.400 289.050 390.450 310.950 ;
        RECT 397.950 307.950 400.050 310.050 ;
        RECT 398.400 298.050 399.450 307.950 ;
        RECT 397.950 295.950 400.050 298.050 ;
        RECT 391.950 294.450 396.000 295.050 ;
        RECT 391.950 292.950 396.450 294.450 ;
        RECT 400.950 292.950 403.050 295.050 ;
        RECT 388.950 286.950 391.050 289.050 ;
        RECT 385.950 271.950 388.050 274.050 ;
        RECT 367.950 268.950 370.050 271.050 ;
        RECT 361.950 266.400 364.050 268.500 ;
        RECT 358.950 259.950 361.050 262.050 ;
        RECT 359.400 256.050 360.450 259.950 ;
        RECT 358.950 253.950 361.050 256.050 ;
        RECT 362.850 251.400 364.050 266.400 ;
        RECT 361.950 249.300 364.050 251.400 ;
        RECT 362.850 245.700 364.050 249.300 ;
        RECT 361.950 243.600 364.050 245.700 ;
        RECT 368.400 238.050 369.450 268.950 ;
        RECT 382.950 266.400 385.050 268.500 ;
        RECT 370.950 262.950 373.050 265.050 ;
        RECT 371.400 259.050 372.450 262.950 ;
        RECT 370.950 256.950 373.050 259.050 ;
        RECT 376.950 253.950 379.050 259.050 ;
        RECT 370.950 250.950 373.050 253.050 ;
        RECT 367.950 235.950 370.050 238.050 ;
        RECT 358.950 226.950 361.050 229.050 ;
        RECT 355.950 221.100 358.050 223.200 ;
        RECT 359.400 220.050 360.450 226.950 ;
        RECT 357.000 219.900 360.450 220.050 ;
        RECT 355.950 218.250 360.450 219.900 ;
        RECT 355.950 217.950 360.000 218.250 ;
        RECT 361.950 217.950 364.050 223.050 ;
        RECT 355.950 217.800 358.050 217.950 ;
        RECT 352.950 211.950 355.050 214.050 ;
        RECT 349.950 205.950 352.050 208.050 ;
        RECT 337.950 202.500 340.050 204.600 ;
        RECT 337.950 184.050 340.050 184.200 ;
        RECT 340.950 184.050 343.050 184.200 ;
        RECT 337.950 182.100 343.050 184.050 ;
        RECT 339.000 181.950 342.000 182.100 ;
        RECT 346.950 181.950 349.050 184.050 ;
        RECT 313.950 178.950 319.050 181.050 ;
        RECT 328.950 179.100 331.050 181.200 ;
        RECT 304.950 175.950 307.050 178.050 ;
        RECT 307.950 175.950 313.050 178.050 ;
        RECT 316.950 177.450 319.050 178.950 ;
        RECT 340.950 178.050 343.050 180.900 ;
        RECT 327.000 177.900 330.000 178.050 ;
        RECT 316.950 176.400 321.450 177.450 ;
        RECT 316.950 175.950 319.050 176.400 ;
        RECT 301.950 157.950 304.050 160.050 ;
        RECT 301.950 151.950 304.050 154.050 ;
        RECT 289.950 148.950 292.050 151.050 ;
        RECT 295.950 148.950 298.050 151.050 ;
        RECT 286.950 136.950 289.050 139.050 ;
        RECT 238.950 133.950 244.050 136.050 ;
        RECT 271.950 133.950 274.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 220.950 131.400 225.450 133.050 ;
        RECT 220.950 130.950 225.000 131.400 ;
        RECT 235.950 130.950 238.050 133.050 ;
        RECT 214.950 101.400 219.450 103.050 ;
        RECT 214.950 100.950 219.000 101.400 ;
        RECT 221.400 100.050 222.450 130.950 ;
        RECT 226.950 103.950 229.050 106.050 ;
        RECT 232.950 103.950 235.050 109.050 ;
        RECT 241.950 103.950 247.050 106.050 ;
        RECT 259.950 103.950 262.050 106.050 ;
        RECT 262.950 103.950 265.050 106.050 ;
        RECT 227.400 100.050 228.450 103.950 ;
        RECT 220.950 97.950 223.050 100.050 ;
        RECT 226.950 97.950 229.050 100.050 ;
        RECT 232.950 97.950 238.050 100.050 ;
        RECT 241.950 97.950 247.050 100.050 ;
        RECT 247.950 97.950 250.050 103.050 ;
        RECT 260.400 97.050 261.450 103.950 ;
        RECT 256.950 95.400 261.450 97.050 ;
        RECT 256.950 94.950 261.000 95.400 ;
        RECT 202.950 88.500 205.050 90.600 ;
        RECT 241.950 88.950 244.050 91.050 ;
        RECT 205.950 82.950 208.050 85.050 ;
        RECT 184.950 73.950 187.050 76.050 ;
        RECT 190.950 73.950 193.050 76.050 ;
        RECT 172.950 68.400 175.050 70.500 ;
        RECT 185.400 70.050 186.450 73.950 ;
        RECT 173.700 48.600 174.900 68.400 ;
        RECT 184.950 67.950 187.050 70.050 ;
        RECT 193.950 69.300 196.050 71.400 ;
        RECT 178.950 55.950 181.050 61.050 ;
        RECT 185.400 58.050 186.450 67.950 ;
        RECT 193.950 65.700 195.150 69.300 ;
        RECT 199.950 67.950 202.050 70.050 ;
        RECT 193.950 63.600 196.050 65.700 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 193.950 48.600 195.150 63.600 ;
        RECT 196.950 52.950 199.050 58.050 ;
        RECT 200.400 52.050 201.450 67.950 ;
        RECT 206.400 64.050 207.450 82.950 ;
        RECT 232.950 73.950 235.050 76.050 ;
        RECT 214.950 67.950 217.050 70.050 ;
        RECT 226.950 68.400 229.050 70.500 ;
        RECT 215.400 64.050 216.450 67.950 ;
        RECT 205.950 61.950 208.050 64.050 ;
        RECT 214.950 61.950 217.050 64.050 ;
        RECT 202.950 55.950 205.050 61.050 ;
        RECT 206.400 55.050 207.450 61.950 ;
        RECT 205.950 52.950 208.050 55.050 ;
        RECT 199.950 49.950 202.050 52.050 ;
        RECT 172.950 46.500 175.050 48.600 ;
        RECT 193.950 46.500 196.050 48.600 ;
        RECT 187.950 37.950 190.050 40.050 ;
        RECT 188.400 25.050 189.450 37.950 ;
        RECT 200.400 28.050 201.450 49.950 ;
        RECT 227.700 48.600 228.900 68.400 ;
        RECT 233.400 61.050 234.450 73.950 ;
        RECT 242.400 61.050 243.450 88.950 ;
        RECT 247.950 69.300 250.050 71.400 ;
        RECT 257.400 70.050 258.450 94.950 ;
        RECT 263.400 76.050 264.450 103.950 ;
        RECT 274.950 100.950 277.050 103.050 ;
        RECT 275.400 85.050 276.450 100.950 ;
        RECT 268.950 82.950 271.050 85.050 ;
        RECT 274.950 82.950 277.050 85.050 ;
        RECT 269.400 79.050 270.450 82.950 ;
        RECT 268.950 76.950 271.050 79.050 ;
        RECT 262.950 73.950 265.050 76.050 ;
        RECT 247.950 65.700 249.150 69.300 ;
        RECT 256.950 67.950 259.050 70.050 ;
        RECT 278.400 67.050 279.450 133.950 ;
        RECT 286.950 112.950 289.050 115.050 ;
        RECT 287.400 106.050 288.450 112.950 ;
        RECT 286.950 103.950 289.050 106.050 ;
        RECT 290.400 100.050 291.450 148.950 ;
        RECT 295.950 142.950 298.050 145.050 ;
        RECT 292.950 133.950 295.050 139.050 ;
        RECT 296.400 133.050 297.450 142.950 ;
        RECT 298.950 139.950 301.050 142.050 ;
        RECT 295.950 130.950 298.050 133.050 ;
        RECT 295.950 100.950 298.050 106.050 ;
        RECT 299.400 100.050 300.450 139.950 ;
        RECT 302.400 136.050 303.450 151.950 ;
        RECT 320.400 139.050 321.450 176.400 ;
        RECT 325.950 175.950 331.050 177.900 ;
        RECT 334.950 175.950 340.050 178.050 ;
        RECT 340.800 177.000 343.050 178.050 ;
        RECT 340.800 175.950 342.900 177.000 ;
        RECT 344.100 175.950 346.200 178.050 ;
        RECT 325.950 175.800 328.050 175.950 ;
        RECT 328.950 175.800 331.050 175.950 ;
        RECT 337.950 169.950 340.050 172.050 ;
        RECT 331.950 157.950 334.050 160.050 ;
        RECT 332.400 142.050 333.450 157.950 ;
        RECT 338.400 142.050 339.450 169.950 ;
        RECT 344.400 163.050 345.450 175.950 ;
        RECT 347.400 172.050 348.450 181.950 ;
        RECT 346.950 169.950 349.050 172.050 ;
        RECT 353.400 169.050 354.450 211.950 ;
        RECT 368.400 211.050 369.450 235.950 ;
        RECT 371.400 229.050 372.450 250.950 ;
        RECT 383.100 246.600 384.300 266.400 ;
        RECT 395.400 256.050 396.450 292.950 ;
        RECT 401.400 289.050 402.450 292.950 ;
        RECT 404.400 289.050 405.450 316.950 ;
        RECT 400.800 286.950 402.900 289.050 ;
        RECT 403.950 286.950 406.050 289.050 ;
        RECT 407.400 265.050 408.450 400.950 ;
        RECT 412.950 381.300 415.050 383.400 ;
        RECT 412.950 377.700 414.150 381.300 ;
        RECT 412.950 375.600 415.050 377.700 ;
        RECT 412.950 360.600 414.150 375.600 ;
        RECT 424.950 373.950 427.050 376.050 ;
        RECT 415.950 370.950 418.050 373.050 ;
        RECT 416.400 367.050 417.450 370.950 ;
        RECT 415.950 364.950 418.050 367.050 ;
        RECT 421.950 364.950 424.050 367.050 ;
        RECT 422.400 361.050 423.450 364.950 ;
        RECT 425.400 361.050 426.450 373.950 ;
        RECT 428.400 369.450 429.450 439.950 ;
        RECT 430.950 415.950 433.050 421.050 ;
        RECT 440.400 420.450 441.450 448.950 ;
        RECT 449.700 438.600 450.900 458.400 ;
        RECT 469.950 455.700 471.150 459.300 ;
        RECT 469.950 453.600 472.050 455.700 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 448.950 436.500 451.050 438.600 ;
        RECT 455.400 421.200 456.450 445.950 ;
        RECT 460.950 442.950 463.050 448.050 ;
        RECT 461.400 424.050 462.450 442.950 ;
        RECT 469.950 438.600 471.150 453.600 ;
        RECT 476.400 445.050 477.450 472.950 ;
        RECT 484.950 457.950 487.050 460.050 ;
        RECT 485.400 448.050 486.450 457.950 ;
        RECT 494.400 454.050 495.450 478.950 ;
        RECT 497.400 472.050 498.450 485.400 ;
        RECT 502.950 478.950 505.050 481.050 ;
        RECT 496.950 469.950 499.050 472.050 ;
        RECT 499.950 463.950 502.050 466.050 ;
        RECT 500.400 457.050 501.450 463.950 ;
        RECT 503.400 463.050 504.450 478.950 ;
        RECT 509.400 478.050 510.450 493.950 ;
        RECT 518.400 490.050 519.450 514.950 ;
        RECT 526.950 514.500 529.050 516.600 ;
        RECT 533.400 505.050 534.450 526.950 ;
        RECT 539.400 526.050 540.450 562.800 ;
        RECT 554.400 559.050 555.450 571.950 ;
        RECT 566.400 568.050 567.450 577.950 ;
        RECT 569.400 574.050 570.450 601.950 ;
        RECT 575.400 601.050 576.450 634.950 ;
        RECT 580.950 625.950 583.050 628.050 ;
        RECT 577.950 619.950 580.050 622.050 ;
        RECT 578.400 610.050 579.450 619.950 ;
        RECT 577.950 607.950 580.050 610.050 ;
        RECT 574.950 598.950 577.050 601.050 ;
        RECT 575.400 580.050 576.450 598.950 ;
        RECT 574.950 577.950 577.050 580.050 ;
        RECT 581.400 577.200 582.450 625.950 ;
        RECT 602.400 622.050 603.450 646.950 ;
        RECT 608.400 646.050 609.450 649.950 ;
        RECT 613.950 646.950 616.050 652.050 ;
        RECT 617.400 646.050 618.450 655.950 ;
        RECT 623.400 654.450 624.450 676.950 ;
        RECT 625.950 673.800 628.050 675.900 ;
        RECT 626.400 661.050 627.450 673.800 ;
        RECT 629.400 661.050 630.450 682.950 ;
        RECT 631.950 676.950 634.050 681.900 ;
        RECT 635.400 667.050 636.450 700.950 ;
        RECT 641.400 673.050 642.450 721.950 ;
        RECT 644.400 721.050 645.450 724.950 ;
        RECT 650.400 724.050 651.450 763.950 ;
        RECT 653.400 760.050 654.450 793.950 ;
        RECT 674.400 790.050 675.450 796.950 ;
        RECT 679.950 793.950 682.050 798.900 ;
        RECT 686.400 790.050 687.450 799.950 ;
        RECT 673.950 787.950 676.050 790.050 ;
        RECT 685.950 787.950 688.050 790.050 ;
        RECT 674.400 775.050 675.450 787.950 ;
        RECT 685.950 775.950 688.050 778.050 ;
        RECT 673.950 772.950 676.050 775.050 ;
        RECT 664.950 766.950 667.050 769.050 ;
        RECT 658.950 760.950 661.050 766.050 ;
        RECT 652.950 757.950 655.050 760.050 ;
        RECT 659.400 751.050 660.450 760.950 ;
        RECT 665.400 760.050 666.450 766.950 ;
        RECT 673.950 760.950 676.050 766.050 ;
        RECT 679.950 763.950 682.050 769.050 ;
        RECT 664.950 757.950 667.050 760.050 ;
        RECT 682.950 757.950 685.050 763.050 ;
        RECT 673.950 751.950 676.050 757.050 ;
        RECT 658.950 748.950 661.050 751.050 ;
        RECT 686.400 739.050 687.450 775.950 ;
        RECT 688.950 763.950 691.050 766.050 ;
        RECT 676.950 736.950 679.050 739.050 ;
        RECT 685.950 736.950 688.050 739.050 ;
        RECT 658.950 727.950 661.050 733.050 ;
        RECT 667.950 724.950 670.050 727.050 ;
        RECT 646.950 721.950 652.050 724.050 ;
        RECT 643.950 718.950 646.050 721.050 ;
        RECT 658.950 718.950 661.050 724.050 ;
        RECT 664.950 718.950 667.050 724.050 ;
        RECT 652.950 709.950 655.050 712.050 ;
        RECT 653.400 691.050 654.450 709.950 ;
        RECT 652.950 688.950 655.050 691.050 ;
        RECT 658.950 688.950 661.050 691.050 ;
        RECT 643.950 685.950 646.050 688.050 ;
        RECT 640.950 670.950 643.050 673.050 ;
        RECT 634.950 664.950 637.050 667.050 ;
        RECT 644.400 661.050 645.450 685.950 ;
        RECT 649.950 682.950 655.050 685.050 ;
        RECT 646.950 676.950 649.050 682.050 ;
        RECT 659.400 679.050 660.450 688.950 ;
        RECT 661.950 682.950 664.050 685.050 ;
        RECT 658.950 676.950 661.050 679.050 ;
        RECT 662.400 678.450 663.450 682.950 ;
        RECT 668.400 682.050 669.450 724.950 ;
        RECT 677.400 724.050 678.450 736.950 ;
        RECT 689.400 730.050 690.450 763.950 ;
        RECT 692.400 754.050 693.450 799.950 ;
        RECT 715.950 796.950 718.050 802.050 ;
        RECT 718.950 796.950 724.050 799.050 ;
        RECT 716.400 778.050 717.450 796.950 ;
        RECT 715.950 775.950 718.050 778.050 ;
        RECT 725.400 772.200 726.450 802.950 ;
        RECT 731.400 799.050 732.450 805.950 ;
        RECT 737.400 802.050 738.450 805.950 ;
        RECT 740.400 802.050 741.450 805.950 ;
        RECT 746.400 805.050 747.450 814.950 ;
        RECT 814.950 813.450 817.050 814.050 ;
        RECT 800.400 812.400 817.050 813.450 ;
        RECT 787.950 810.450 790.050 811.050 ;
        RECT 779.400 810.000 790.050 810.450 ;
        RECT 778.950 809.400 790.050 810.000 ;
        RECT 748.950 805.950 751.050 808.050 ;
        RECT 757.950 805.950 760.050 808.050 ;
        RECT 760.950 805.950 763.050 808.050 ;
        RECT 778.950 805.950 781.050 809.400 ;
        RECT 787.950 808.950 790.050 809.400 ;
        RECT 736.950 799.950 739.050 802.050 ;
        RECT 739.950 799.950 742.050 802.050 ;
        RECT 745.950 799.950 748.050 805.050 ;
        RECT 727.950 797.400 732.450 799.050 ;
        RECT 727.950 796.950 732.000 797.400 ;
        RECT 724.950 770.100 727.050 772.200 ;
        RECT 724.950 766.800 727.050 768.900 ;
        RECT 694.950 757.950 697.050 763.050 ;
        RECT 700.950 760.950 703.050 763.050 ;
        RECT 712.950 760.950 715.050 766.050 ;
        RECT 718.950 760.950 721.050 763.050 ;
        RECT 701.400 757.050 702.450 760.950 ;
        RECT 697.950 754.950 700.050 757.050 ;
        RECT 700.950 754.950 703.050 757.050 ;
        RECT 691.950 751.950 694.050 754.050 ;
        RECT 691.950 733.950 694.050 736.050 ;
        RECT 682.950 727.950 685.050 730.050 ;
        RECT 683.400 724.050 684.450 727.950 ;
        RECT 685.950 724.950 688.050 730.050 ;
        RECT 688.950 727.950 691.050 730.050 ;
        RECT 676.950 721.950 679.050 724.050 ;
        RECT 682.950 721.950 685.050 724.050 ;
        RECT 673.950 709.950 676.050 712.050 ;
        RECT 670.950 685.950 673.050 688.050 ;
        RECT 671.400 682.050 672.450 685.950 ;
        RECT 664.950 679.950 669.450 682.050 ;
        RECT 670.950 679.950 673.050 682.050 ;
        RECT 662.400 677.400 666.450 678.450 ;
        RECT 625.800 658.950 627.900 661.050 ;
        RECT 629.100 658.950 631.200 661.050 ;
        RECT 634.950 658.950 637.050 661.050 ;
        RECT 643.950 658.950 646.050 661.050 ;
        RECT 620.400 653.400 624.450 654.450 ;
        RECT 607.950 643.950 610.050 646.050 ;
        RECT 610.950 643.950 613.050 646.050 ;
        RECT 616.950 645.450 619.050 646.050 ;
        RECT 614.400 644.400 619.050 645.450 ;
        RECT 611.400 640.050 612.450 643.950 ;
        RECT 610.950 637.950 613.050 640.050 ;
        RECT 601.950 619.950 604.050 622.050 ;
        RECT 607.950 613.950 610.050 616.050 ;
        RECT 601.950 607.950 604.050 613.050 ;
        RECT 608.400 604.050 609.450 613.950 ;
        RECT 614.400 610.050 615.450 644.400 ;
        RECT 616.950 643.950 619.050 644.400 ;
        RECT 620.400 639.450 621.450 653.400 ;
        RECT 622.950 649.950 628.050 652.050 ;
        RECT 635.400 649.050 636.450 658.950 ;
        RECT 665.400 652.050 666.450 677.400 ;
        RECT 668.400 664.050 669.450 679.950 ;
        RECT 667.950 661.950 670.050 664.050 ;
        RECT 674.400 658.050 675.450 709.950 ;
        RECT 678.000 690.450 682.050 691.050 ;
        RECT 677.400 688.950 682.050 690.450 ;
        RECT 677.400 676.050 678.450 688.950 ;
        RECT 692.400 688.050 693.450 733.950 ;
        RECT 694.950 727.950 697.050 730.050 ;
        RECT 695.400 706.050 696.450 727.950 ;
        RECT 698.400 712.050 699.450 754.950 ;
        RECT 703.950 751.950 706.050 757.050 ;
        RECT 706.950 754.950 712.050 757.050 ;
        RECT 704.400 733.050 705.450 751.950 ;
        RECT 712.950 745.950 715.050 748.050 ;
        RECT 703.950 730.950 706.050 733.050 ;
        RECT 704.400 715.050 705.450 730.950 ;
        RECT 713.400 724.050 714.450 745.950 ;
        RECT 719.400 733.050 720.450 760.950 ;
        RECT 718.950 730.950 721.050 733.050 ;
        RECT 715.950 727.950 718.050 730.050 ;
        RECT 721.950 727.950 724.050 730.050 ;
        RECT 706.950 721.950 709.050 724.050 ;
        RECT 712.950 721.950 715.050 724.050 ;
        RECT 703.950 712.950 706.050 715.050 ;
        RECT 697.950 709.950 700.050 712.050 ;
        RECT 694.950 703.950 697.050 706.050 ;
        RECT 707.400 694.050 708.450 721.950 ;
        RECT 716.400 703.050 717.450 727.950 ;
        RECT 722.400 718.050 723.450 727.950 ;
        RECT 725.400 724.050 726.450 766.800 ;
        RECT 749.400 766.050 750.450 805.950 ;
        RECT 758.400 802.050 759.450 805.950 ;
        RECT 761.400 802.050 762.450 805.950 ;
        RECT 784.950 802.950 787.050 808.050 ;
        RECT 800.400 805.050 801.450 812.400 ;
        RECT 814.950 811.950 817.050 812.400 ;
        RECT 823.950 811.950 826.050 814.050 ;
        RECT 802.950 808.950 805.050 811.050 ;
        RECT 811.950 808.950 814.050 811.050 ;
        RECT 803.400 805.200 804.450 808.950 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 802.950 803.100 805.050 805.200 ;
        RECT 805.950 802.050 808.050 805.050 ;
        RECT 757.950 799.950 760.050 802.050 ;
        RECT 760.950 799.950 763.050 802.050 ;
        RECT 766.950 799.950 769.050 802.050 ;
        RECT 781.950 801.450 786.000 802.050 ;
        RECT 781.950 799.950 786.450 801.450 ;
        RECT 754.950 796.950 757.050 799.050 ;
        RECT 730.950 760.950 733.050 766.050 ;
        RECT 748.950 765.450 751.050 766.050 ;
        RECT 746.400 764.400 751.050 765.450 ;
        RECT 736.950 760.950 739.050 763.050 ;
        RECT 727.950 754.950 730.050 760.050 ;
        RECT 733.950 754.950 736.050 757.050 ;
        RECT 734.400 742.050 735.450 754.950 ;
        RECT 733.950 739.950 736.050 742.050 ;
        RECT 724.950 721.950 727.050 724.050 ;
        RECT 721.950 715.950 724.050 718.050 ;
        RECT 722.400 709.050 723.450 715.950 ;
        RECT 721.950 706.950 724.050 709.050 ;
        RECT 733.950 703.950 736.050 706.050 ;
        RECT 715.950 700.950 718.050 703.050 ;
        RECT 706.950 691.950 709.050 694.050 ;
        RECT 691.950 685.950 694.050 688.050 ;
        RECT 700.950 686.100 703.050 691.050 ;
        RECT 718.950 688.950 721.050 691.050 ;
        RECT 709.950 685.950 712.050 688.050 ;
        RECT 712.950 685.950 715.050 688.050 ;
        RECT 682.950 685.050 685.050 685.200 ;
        RECT 703.950 685.050 706.050 685.200 ;
        RECT 681.000 684.600 685.050 685.050 ;
        RECT 702.000 684.900 706.050 685.050 ;
        RECT 680.400 683.100 685.050 684.600 ;
        RECT 700.950 683.100 706.050 684.900 ;
        RECT 680.400 682.950 684.000 683.100 ;
        RECT 700.950 682.950 705.000 683.100 ;
        RECT 676.950 673.950 679.050 676.050 ;
        RECT 673.950 655.950 676.050 658.050 ;
        RECT 680.400 652.050 681.450 682.950 ;
        RECT 700.950 682.800 703.050 682.950 ;
        RECT 684.000 681.900 688.050 682.050 ;
        RECT 705.000 681.900 709.050 682.050 ;
        RECT 682.950 679.950 688.050 681.900 ;
        RECT 703.950 679.950 709.050 681.900 ;
        RECT 682.950 679.800 685.050 679.950 ;
        RECT 703.950 679.800 706.050 679.950 ;
        RECT 697.950 661.950 700.050 664.050 ;
        RECT 682.950 655.950 685.050 658.050 ;
        RECT 658.950 649.950 661.050 652.050 ;
        RECT 664.950 649.950 667.050 652.050 ;
        RECT 670.950 649.950 676.050 652.050 ;
        RECT 679.950 649.950 682.050 652.050 ;
        RECT 634.950 646.950 637.050 649.050 ;
        RECT 631.950 643.950 634.050 646.050 ;
        RECT 628.950 640.950 631.050 643.050 ;
        RECT 620.400 638.400 624.450 639.450 ;
        RECT 623.400 625.050 624.450 638.400 ;
        RECT 622.950 622.950 625.050 625.050 ;
        RECT 623.400 610.050 624.450 622.950 ;
        RECT 629.400 613.050 630.450 640.950 ;
        RECT 628.950 610.950 631.050 613.050 ;
        RECT 613.950 607.950 616.050 610.050 ;
        RECT 619.950 608.400 624.450 610.050 ;
        RECT 619.950 607.950 624.000 608.400 ;
        RECT 625.950 607.950 628.050 610.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 607.950 601.950 610.050 604.050 ;
        RECT 583.950 598.950 586.050 601.050 ;
        RECT 580.950 575.100 583.050 577.200 ;
        RECT 568.950 571.950 571.050 574.050 ;
        RECT 574.950 571.950 577.050 574.050 ;
        RECT 565.950 565.950 568.050 568.050 ;
        RECT 571.950 565.950 574.050 571.050 ;
        RECT 566.400 559.050 567.450 565.950 ;
        RECT 575.400 562.050 576.450 571.950 ;
        RECT 580.950 571.800 583.050 573.900 ;
        RECT 581.400 562.050 582.450 571.800 ;
        RECT 584.400 568.050 585.450 598.950 ;
        RECT 586.950 595.950 589.050 598.050 ;
        RECT 587.400 574.050 588.450 595.950 ;
        RECT 595.950 580.950 598.050 583.050 ;
        RECT 596.400 574.050 597.450 580.950 ;
        RECT 602.400 574.050 603.450 601.950 ;
        RECT 626.400 598.050 627.450 607.950 ;
        RECT 629.400 601.050 630.450 610.950 ;
        RECT 632.400 610.050 633.450 643.950 ;
        RECT 637.950 640.950 643.050 643.050 ;
        RECT 646.950 640.950 649.050 643.050 ;
        RECT 640.950 628.950 643.050 631.050 ;
        RECT 641.400 610.050 642.450 628.950 ;
        RECT 631.950 604.950 634.050 610.050 ;
        RECT 640.950 607.950 643.050 610.050 ;
        RECT 647.400 607.050 648.450 640.950 ;
        RECT 634.950 601.950 637.050 607.050 ;
        RECT 643.950 604.950 649.050 607.050 ;
        RECT 652.950 604.950 655.050 610.050 ;
        RECT 628.950 598.950 631.050 601.050 ;
        RECT 610.950 595.950 613.050 598.050 ;
        RECT 625.950 595.950 628.050 598.050 ;
        RECT 586.950 571.950 589.050 574.050 ;
        RECT 589.950 571.950 592.050 574.050 ;
        RECT 595.950 571.950 598.050 574.050 ;
        RECT 602.400 572.400 607.050 574.050 ;
        RECT 603.000 571.950 607.050 572.400 ;
        RECT 590.400 568.050 591.450 571.950 ;
        RECT 584.400 566.400 589.050 568.050 ;
        RECT 585.000 565.950 589.050 566.400 ;
        RECT 589.950 565.950 592.050 568.050 ;
        RECT 592.950 562.950 595.050 568.050 ;
        RECT 598.950 565.950 604.050 568.050 ;
        RECT 568.950 559.950 571.050 562.050 ;
        RECT 574.950 559.950 577.050 562.050 ;
        RECT 580.950 559.950 583.050 562.050 ;
        RECT 553.950 556.950 556.050 559.050 ;
        RECT 559.950 556.950 562.050 559.050 ;
        RECT 565.950 556.950 568.050 559.050 ;
        RECT 556.950 550.950 559.050 553.050 ;
        RECT 547.950 535.950 550.050 538.050 ;
        RECT 548.400 532.050 549.450 535.950 ;
        RECT 548.400 530.400 553.050 532.050 ;
        RECT 549.000 529.950 553.050 530.400 ;
        RECT 557.400 526.200 558.450 550.950 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 556.950 524.100 559.050 526.200 ;
        RECT 539.400 505.050 540.450 523.950 ;
        RECT 556.950 520.800 559.050 522.900 ;
        RECT 557.400 517.050 558.450 520.800 ;
        RECT 556.950 514.950 559.050 517.050 ;
        RECT 547.950 511.950 550.050 514.050 ;
        RECT 532.950 502.950 535.050 505.050 ;
        RECT 538.950 502.950 541.050 505.050 ;
        RECT 526.950 499.950 529.050 502.050 ;
        RECT 527.400 490.050 528.450 499.950 ;
        RECT 538.950 496.950 541.050 499.050 ;
        RECT 532.950 490.950 538.050 493.050 ;
        RECT 511.950 487.950 517.050 490.050 ;
        RECT 517.950 487.950 520.050 490.050 ;
        RECT 526.950 487.950 529.050 490.050 ;
        RECT 539.400 487.050 540.450 496.950 ;
        RECT 544.950 493.950 547.050 496.050 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 538.950 484.950 541.050 487.050 ;
        RECT 508.950 475.950 511.050 478.050 ;
        RECT 505.950 463.950 508.050 466.050 ;
        RECT 523.950 463.950 526.050 466.050 ;
        RECT 502.950 460.950 505.050 463.050 ;
        RECT 499.950 454.950 502.050 457.050 ;
        RECT 487.950 451.950 490.050 454.050 ;
        RECT 493.950 451.950 496.050 454.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 472.950 442.950 478.050 445.050 ;
        RECT 469.950 436.500 472.050 438.600 ;
        RECT 488.400 436.050 489.450 451.950 ;
        RECT 494.400 448.050 495.450 451.950 ;
        RECT 506.400 451.050 507.450 463.950 ;
        RECT 511.950 457.950 514.050 460.050 ;
        RECT 512.400 451.050 513.450 457.950 ;
        RECT 505.950 448.950 508.050 451.050 ;
        RECT 511.950 448.950 514.050 451.050 ;
        RECT 520.950 448.950 523.050 451.050 ;
        RECT 493.950 445.950 496.050 448.050 ;
        RECT 502.950 442.950 505.050 448.050 ;
        RECT 521.400 445.050 522.450 448.950 ;
        RECT 524.400 445.050 525.450 463.950 ;
        RECT 535.950 458.400 538.050 460.500 ;
        RECT 508.950 442.950 511.050 445.050 ;
        RECT 520.950 442.950 523.050 445.050 ;
        RECT 523.950 442.950 526.050 445.050 ;
        RECT 487.950 433.950 490.050 436.050 ;
        RECT 509.400 433.050 510.450 442.950 ;
        RECT 536.700 438.600 537.900 458.400 ;
        RECT 542.400 457.050 543.450 487.950 ;
        RECT 545.400 481.050 546.450 493.950 ;
        RECT 548.400 490.050 549.450 511.950 ;
        RECT 553.950 493.950 556.050 496.050 ;
        RECT 547.950 487.950 550.050 490.050 ;
        RECT 554.400 484.050 555.450 493.950 ;
        RECT 560.400 490.050 561.450 556.950 ;
        RECT 566.400 538.200 567.450 556.950 ;
        RECT 565.950 536.100 568.050 538.200 ;
        RECT 565.950 532.800 568.050 534.900 ;
        RECT 566.400 529.050 567.450 532.800 ;
        RECT 565.950 526.950 568.050 529.050 ;
        RECT 569.400 523.050 570.450 559.950 ;
        RECT 611.400 553.050 612.450 595.950 ;
        RECT 629.400 594.450 630.450 598.950 ;
        RECT 626.400 593.400 630.450 594.450 ;
        RECT 619.950 580.950 622.050 583.050 ;
        RECT 620.400 574.050 621.450 580.950 ;
        RECT 619.950 571.950 622.050 574.050 ;
        RECT 613.950 568.950 619.050 571.050 ;
        RECT 626.400 568.050 627.450 593.400 ;
        RECT 635.400 589.050 636.450 601.950 ;
        RECT 659.400 601.050 660.450 649.950 ;
        RECT 665.400 631.050 666.450 649.950 ;
        RECT 683.400 646.050 684.450 655.950 ;
        RECT 688.950 649.950 694.050 652.050 ;
        RECT 698.400 646.050 699.450 661.950 ;
        RECT 710.400 646.050 711.450 685.950 ;
        RECT 713.400 679.050 714.450 685.950 ;
        RECT 712.950 676.950 715.050 679.050 ;
        RECT 719.400 673.050 720.450 688.950 ;
        RECT 721.950 682.950 724.050 685.050 ;
        RECT 718.950 670.950 721.050 673.050 ;
        RECT 719.400 652.050 720.450 670.950 ;
        RECT 722.400 661.050 723.450 682.950 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 721.950 658.950 724.050 661.050 ;
        RECT 712.950 646.950 715.050 652.050 ;
        RECT 718.950 649.950 721.050 652.050 ;
        RECT 725.400 649.200 726.450 679.950 ;
        RECT 730.950 658.950 733.050 661.050 ;
        RECT 724.950 647.100 727.050 649.200 ;
        RECT 731.400 646.050 732.450 658.950 ;
        RECT 734.400 654.450 735.450 703.950 ;
        RECT 737.400 700.050 738.450 760.950 ;
        RECT 739.950 754.950 745.050 757.050 ;
        RECT 746.400 744.450 747.450 764.400 ;
        RECT 748.950 763.950 751.050 764.400 ;
        RECT 755.400 763.050 756.450 796.950 ;
        RECT 767.400 793.050 768.450 799.950 ;
        RECT 778.950 793.950 781.050 796.050 ;
        RECT 766.950 790.950 769.050 793.050 ;
        RECT 763.950 772.950 766.050 775.050 ;
        RECT 760.950 766.950 763.050 769.050 ;
        RECT 761.400 763.050 762.450 766.950 ;
        RECT 754.950 760.950 757.050 763.050 ;
        RECT 760.950 760.950 763.050 763.050 ;
        RECT 748.950 754.950 754.050 757.050 ;
        RECT 757.950 754.950 760.050 757.050 ;
        RECT 743.400 743.400 747.450 744.450 ;
        RECT 743.400 727.050 744.450 743.400 ;
        RECT 745.950 739.950 748.050 742.050 ;
        RECT 746.400 730.050 747.450 739.950 ;
        RECT 745.950 727.950 748.050 730.050 ;
        RECT 742.950 724.950 745.050 727.050 ;
        RECT 746.400 724.050 747.450 727.950 ;
        RECT 758.400 726.450 759.450 754.950 ;
        RECT 764.400 727.050 765.450 772.950 ;
        RECT 767.400 769.050 768.450 790.950 ;
        RECT 766.950 766.950 769.050 769.050 ;
        RECT 775.950 763.950 778.050 766.050 ;
        RECT 776.400 751.050 777.450 763.950 ;
        RECT 779.400 763.200 780.450 793.950 ;
        RECT 785.400 772.200 786.450 799.950 ;
        RECT 793.950 796.950 796.050 802.050 ;
        RECT 804.000 801.900 808.050 802.050 ;
        RECT 802.950 799.950 808.050 801.900 ;
        RECT 812.400 802.050 813.450 808.950 ;
        RECT 824.400 808.050 825.450 811.950 ;
        RECT 817.950 802.950 820.050 808.050 ;
        RECT 823.950 805.950 826.050 808.050 ;
        RECT 812.400 800.400 817.050 802.050 ;
        RECT 813.000 799.950 817.050 800.400 ;
        RECT 802.950 799.800 805.050 799.950 ;
        RECT 799.950 796.950 802.050 799.050 ;
        RECT 800.400 775.050 801.450 796.950 ;
        RECT 808.950 793.950 811.050 799.050 ;
        RECT 820.950 796.950 823.050 802.050 ;
        RECT 799.950 772.950 802.050 775.050 ;
        RECT 784.950 770.100 787.050 772.200 ;
        RECT 793.950 769.950 796.050 772.050 ;
        RECT 783.000 768.900 786.000 769.050 ;
        RECT 781.950 766.950 787.050 768.900 ;
        RECT 781.950 766.800 784.050 766.950 ;
        RECT 784.950 766.800 787.050 766.950 ;
        RECT 778.950 763.050 781.050 763.200 ;
        RECT 794.400 763.050 795.450 769.950 ;
        RECT 799.950 766.950 802.050 769.050 ;
        RECT 800.400 763.050 801.450 766.950 ;
        RECT 778.950 761.100 784.050 763.050 ;
        RECT 780.000 760.950 784.050 761.100 ;
        RECT 778.950 754.950 781.050 759.900 ;
        RECT 793.950 757.950 796.050 763.050 ;
        RECT 796.950 760.950 799.050 763.050 ;
        RECT 799.950 760.950 802.050 763.050 ;
        RECT 805.950 760.950 808.050 763.050 ;
        RECT 797.400 757.050 798.450 760.950 ;
        RECT 806.400 757.050 807.450 760.950 ;
        RECT 809.400 757.050 810.450 793.950 ;
        RECT 814.950 760.950 820.050 763.050 ;
        RECT 823.950 762.450 828.000 763.050 ;
        RECT 823.950 760.950 828.450 762.450 ;
        RECT 796.950 754.950 799.050 757.050 ;
        RECT 805.800 754.950 807.900 757.050 ;
        RECT 808.950 754.950 811.050 757.050 ;
        RECT 814.950 754.950 817.050 757.050 ;
        RECT 820.950 754.950 823.050 757.050 ;
        RECT 775.950 748.950 778.050 751.050 ;
        RECT 776.400 730.050 777.450 748.950 ;
        RECT 815.400 745.050 816.450 754.950 ;
        RECT 814.950 742.950 817.050 745.050 ;
        RECT 799.950 733.950 802.050 736.050 ;
        RECT 775.950 727.950 778.050 730.050 ;
        RECT 755.400 725.400 759.450 726.450 ;
        RECT 739.950 718.950 742.050 724.050 ;
        RECT 745.950 721.950 748.050 724.050 ;
        RECT 736.950 697.950 739.050 700.050 ;
        RECT 740.400 688.050 741.450 718.950 ;
        RECT 736.950 684.450 739.050 688.050 ;
        RECT 739.950 685.950 742.050 688.050 ;
        RECT 746.400 685.050 747.450 721.950 ;
        RECT 748.950 715.950 751.050 718.050 ;
        RECT 749.400 700.050 750.450 715.950 ;
        RECT 748.950 697.950 751.050 700.050 ;
        RECT 751.950 685.950 754.050 688.050 ;
        RECT 742.950 684.450 745.050 685.050 ;
        RECT 736.950 684.000 745.050 684.450 ;
        RECT 737.400 683.400 745.050 684.000 ;
        RECT 746.400 683.400 751.050 685.050 ;
        RECT 742.950 682.950 745.050 683.400 ;
        RECT 747.000 682.950 751.050 683.400 ;
        RECT 752.400 679.050 753.450 685.950 ;
        RECT 736.950 676.950 742.050 679.050 ;
        RECT 745.950 676.950 751.050 679.050 ;
        RECT 751.950 676.950 754.050 679.050 ;
        RECT 755.400 675.450 756.450 725.400 ;
        RECT 763.950 724.950 766.050 727.050 ;
        RECT 757.950 721.950 763.050 724.050 ;
        RECT 766.950 718.950 769.050 721.050 ;
        RECT 757.950 715.950 763.050 718.050 ;
        RECT 762.000 681.450 766.050 682.050 ;
        RECT 761.400 681.000 766.050 681.450 ;
        RECT 760.950 679.950 766.050 681.000 ;
        RECT 760.950 676.950 763.050 679.950 ;
        RECT 767.400 679.050 768.450 718.950 ;
        RECT 776.400 718.050 777.450 727.950 ;
        RECT 784.950 724.950 790.050 727.050 ;
        RECT 790.950 724.950 796.050 727.050 ;
        RECT 778.950 721.950 784.050 724.050 ;
        RECT 800.400 721.050 801.450 733.950 ;
        RECT 821.400 727.200 822.450 754.950 ;
        RECT 827.400 751.050 828.450 760.950 ;
        RECT 826.950 748.950 829.050 751.050 ;
        RECT 823.950 733.950 826.050 736.050 ;
        RECT 820.950 727.050 823.050 727.200 ;
        RECT 817.950 725.100 823.050 727.050 ;
        RECT 817.950 724.950 822.000 725.100 ;
        RECT 824.400 724.050 825.450 733.950 ;
        RECT 826.950 724.950 829.050 727.050 ;
        RECT 822.000 723.900 825.450 724.050 ;
        RECT 820.950 722.250 825.450 723.900 ;
        RECT 820.950 721.950 825.000 722.250 ;
        RECT 820.950 721.800 823.050 721.950 ;
        RECT 790.950 718.950 793.050 721.050 ;
        RECT 799.950 718.950 802.050 721.050 ;
        RECT 776.400 716.400 781.050 718.050 ;
        RECT 777.000 715.950 781.050 716.400 ;
        RECT 791.400 688.050 792.450 718.950 ;
        RECT 805.950 715.950 808.050 721.050 ;
        RECT 811.950 718.950 814.050 721.050 ;
        RECT 821.400 720.450 822.450 721.800 ;
        RECT 818.400 719.400 822.450 720.450 ;
        RECT 812.400 688.050 813.450 718.950 ;
        RECT 814.950 715.950 817.050 718.050 ;
        RECT 787.800 687.000 789.900 688.050 ;
        RECT 787.800 685.950 790.050 687.000 ;
        RECT 791.100 685.950 793.200 688.050 ;
        RECT 799.950 685.950 805.050 688.050 ;
        RECT 808.950 686.400 813.450 688.050 ;
        RECT 808.950 685.950 813.000 686.400 ;
        RECT 769.950 682.950 775.050 685.050 ;
        RECT 781.950 679.950 784.050 685.050 ;
        RECT 787.950 682.950 790.050 685.950 ;
        RECT 808.950 682.950 811.050 685.950 ;
        RECT 815.400 685.050 816.450 715.950 ;
        RECT 814.950 682.950 817.050 685.050 ;
        RECT 793.950 679.950 796.050 682.050 ;
        RECT 766.950 676.950 769.050 679.050 ;
        RECT 775.950 676.950 781.050 679.050 ;
        RECT 784.950 676.950 787.050 679.050 ;
        RECT 755.400 674.400 759.450 675.450 ;
        RECT 754.950 670.950 757.050 673.050 ;
        RECT 734.400 653.400 738.450 654.450 ;
        RECT 733.950 646.950 736.050 652.050 ;
        RECT 670.950 640.950 673.050 646.050 ;
        RECT 676.950 640.950 679.050 646.050 ;
        RECT 682.950 643.950 685.050 646.050 ;
        RECT 694.950 640.950 697.050 646.050 ;
        RECT 698.400 644.400 703.050 646.050 ;
        RECT 699.000 643.950 703.050 644.400 ;
        RECT 709.950 643.950 712.050 646.050 ;
        RECT 724.950 643.800 727.050 645.900 ;
        RECT 730.950 643.950 733.050 646.050 ;
        RECT 725.400 640.050 726.450 643.800 ;
        RECT 725.400 638.400 730.050 640.050 ;
        RECT 726.000 637.950 730.050 638.400 ;
        RECT 664.950 628.950 667.050 631.050 ;
        RECT 670.950 628.950 673.050 631.050 ;
        RECT 667.950 613.950 670.050 616.050 ;
        RECT 668.400 607.050 669.450 613.950 ;
        RECT 671.400 607.050 672.450 628.950 ;
        RECT 703.950 625.950 706.050 628.050 ;
        RECT 679.950 622.950 682.050 625.050 ;
        RECT 667.950 604.950 670.050 607.050 ;
        RECT 670.950 604.950 673.050 607.050 ;
        RECT 673.950 606.450 678.000 607.050 ;
        RECT 673.950 604.950 678.450 606.450 ;
        RECT 671.400 601.050 672.450 604.950 ;
        RECT 646.950 598.950 652.050 601.050 ;
        RECT 658.950 598.950 661.050 601.050 ;
        RECT 670.950 598.950 673.050 601.050 ;
        RECT 664.950 595.950 667.050 598.050 ;
        RECT 634.950 586.950 637.050 589.050 ;
        RECT 649.950 586.950 652.050 589.050 ;
        RECT 634.950 571.950 637.050 574.050 ;
        RECT 622.950 562.950 625.050 568.050 ;
        RECT 625.950 565.950 628.050 568.050 ;
        RECT 628.950 565.950 631.050 571.050 ;
        RECT 635.400 567.450 636.450 571.950 ;
        RECT 650.400 571.050 651.450 586.950 ;
        RECT 665.400 574.050 666.450 595.950 ;
        RECT 677.400 589.050 678.450 604.950 ;
        RECT 676.950 586.950 679.050 589.050 ;
        RECT 652.950 571.950 658.050 574.050 ;
        RECT 664.950 571.950 667.050 574.050 ;
        RECT 643.950 568.950 646.050 571.050 ;
        RECT 649.950 568.950 652.050 571.050 ;
        RECT 670.950 568.950 673.050 571.050 ;
        RECT 635.400 566.400 639.450 567.450 ;
        RECT 610.950 550.950 613.050 553.050 ;
        RECT 574.950 547.950 577.050 550.050 ;
        RECT 604.950 547.950 607.050 550.050 ;
        RECT 571.950 535.950 574.050 538.050 ;
        RECT 568.950 520.950 571.050 523.050 ;
        RECT 572.400 493.050 573.450 535.950 ;
        RECT 575.400 535.050 576.450 547.950 ;
        RECT 589.950 544.950 592.050 547.050 ;
        RECT 583.950 541.950 586.050 544.050 ;
        RECT 574.950 532.950 577.050 535.050 ;
        RECT 574.950 526.950 577.050 529.050 ;
        RECT 577.950 526.950 580.050 529.050 ;
        RECT 575.400 523.050 576.450 526.950 ;
        RECT 574.950 520.950 577.050 523.050 ;
        RECT 578.400 502.050 579.450 526.950 ;
        RECT 580.950 520.950 583.050 526.050 ;
        RECT 580.950 504.450 583.050 505.050 ;
        RECT 584.400 504.450 585.450 541.950 ;
        RECT 586.950 538.950 589.050 541.050 ;
        RECT 587.400 532.050 588.450 538.950 ;
        RECT 590.400 535.050 591.450 544.950 ;
        RECT 589.950 532.950 592.050 535.050 ;
        RECT 586.950 529.950 589.050 532.050 ;
        RECT 592.950 526.950 595.050 532.050 ;
        RECT 598.950 529.950 601.050 532.050 ;
        RECT 586.950 523.950 592.050 526.050 ;
        RECT 599.400 520.050 600.450 529.950 ;
        RECT 605.400 522.450 606.450 547.950 ;
        RECT 607.950 529.950 610.050 532.050 ;
        RECT 602.400 521.400 606.450 522.450 ;
        RECT 586.950 517.950 589.050 520.050 ;
        RECT 598.950 517.950 601.050 520.050 ;
        RECT 580.950 503.400 585.450 504.450 ;
        RECT 580.950 502.950 583.050 503.400 ;
        RECT 577.950 499.950 580.050 502.050 ;
        RECT 581.400 496.050 582.450 502.950 ;
        RECT 577.950 494.400 582.450 496.050 ;
        RECT 577.950 493.950 582.000 494.400 ;
        RECT 565.950 490.950 571.050 493.050 ;
        RECT 571.950 490.950 574.050 493.050 ;
        RECT 587.400 490.050 588.450 517.950 ;
        RECT 602.400 514.050 603.450 521.400 ;
        RECT 604.950 517.950 607.050 520.050 ;
        RECT 601.950 511.950 604.050 514.050 ;
        RECT 605.400 499.050 606.450 517.950 ;
        RECT 608.400 517.050 609.450 529.950 ;
        RECT 619.950 528.450 622.050 529.050 ;
        RECT 623.400 528.450 624.450 562.950 ;
        RECT 626.400 541.050 627.450 565.950 ;
        RECT 634.950 559.950 637.050 565.050 ;
        RECT 628.950 556.950 631.050 559.050 ;
        RECT 625.950 538.950 628.050 541.050 ;
        RECT 629.400 529.050 630.450 556.950 ;
        RECT 638.400 538.050 639.450 566.400 ;
        RECT 644.400 565.050 645.450 568.950 ;
        RECT 658.950 565.950 661.050 568.050 ;
        RECT 643.950 562.950 646.050 565.050 ;
        RECT 640.950 550.950 643.050 553.050 ;
        RECT 637.950 535.950 640.050 538.050 ;
        RECT 619.950 527.400 624.450 528.450 ;
        RECT 619.950 523.950 622.050 527.400 ;
        RECT 628.950 526.950 631.050 529.050 ;
        RECT 634.950 526.950 637.050 532.050 ;
        RECT 625.950 520.950 628.050 523.050 ;
        RECT 637.950 520.950 640.050 526.050 ;
        RECT 607.950 514.950 610.050 517.050 ;
        RECT 626.400 511.050 627.450 520.950 ;
        RECT 625.950 508.950 628.050 511.050 ;
        RECT 625.950 502.950 628.050 505.050 ;
        RECT 604.950 496.950 607.050 499.050 ;
        RECT 559.950 487.950 562.050 490.050 ;
        RECT 586.950 487.950 589.050 490.050 ;
        RECT 553.950 481.950 556.050 484.050 ;
        RECT 544.950 478.950 547.050 481.050 ;
        RECT 560.400 466.050 561.450 487.950 ;
        RECT 605.400 487.050 606.450 496.950 ;
        RECT 626.400 496.050 627.450 502.950 ;
        RECT 607.950 490.950 610.050 496.050 ;
        RECT 616.950 493.950 619.050 496.050 ;
        RECT 625.950 493.950 628.050 496.050 ;
        RECT 617.400 487.050 618.450 493.950 ;
        RECT 619.950 487.950 622.050 493.050 ;
        RECT 626.400 490.050 627.450 493.950 ;
        RECT 625.950 487.950 628.050 490.050 ;
        RECT 628.950 487.950 631.050 493.050 ;
        RECT 641.400 492.450 642.450 550.950 ;
        RECT 659.400 544.050 660.450 565.950 ;
        RECT 664.950 562.950 667.050 568.050 ;
        RECT 664.950 556.950 667.050 559.050 ;
        RECT 658.950 541.950 661.050 544.050 ;
        RECT 659.400 532.050 660.450 541.950 ;
        RECT 658.950 529.950 661.050 532.050 ;
        RECT 646.950 523.950 649.050 526.050 ;
        RECT 652.950 523.950 655.050 529.050 ;
        RECT 665.400 526.050 666.450 556.950 ;
        RECT 671.400 547.050 672.450 568.950 ;
        RECT 680.400 553.050 681.450 622.950 ;
        RECT 688.950 610.950 691.050 616.050 ;
        RECT 688.950 607.050 691.050 607.200 ;
        RECT 688.950 605.100 694.050 607.050 ;
        RECT 690.000 604.950 694.050 605.100 ;
        RECT 688.950 598.950 691.050 603.900 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 695.400 589.050 696.450 601.950 ;
        RECT 694.950 586.950 697.050 589.050 ;
        RECT 691.950 562.950 694.050 565.050 ;
        RECT 697.950 562.950 700.050 565.050 ;
        RECT 692.400 559.050 693.450 562.950 ;
        RECT 691.800 556.950 693.900 559.050 ;
        RECT 695.100 556.950 697.200 559.050 ;
        RECT 679.950 550.950 682.050 553.050 ;
        RECT 670.950 544.950 673.050 547.050 ;
        RECT 670.950 535.950 673.050 538.050 ;
        RECT 682.950 535.950 685.050 538.050 ;
        RECT 671.400 532.050 672.450 535.950 ;
        RECT 670.950 529.950 673.050 532.050 ;
        RECT 673.950 529.950 676.050 532.050 ;
        RECT 676.950 529.950 679.050 532.050 ;
        RECT 647.400 505.050 648.450 523.950 ;
        RECT 658.950 520.950 661.050 526.050 ;
        RECT 664.950 523.950 667.050 526.050 ;
        RECT 646.950 502.950 649.050 505.050 ;
        RECT 641.400 491.400 645.450 492.450 ;
        RECT 640.950 490.050 643.050 490.200 ;
        RECT 637.950 488.100 643.050 490.050 ;
        RECT 637.950 487.950 642.000 488.100 ;
        RECT 592.950 484.950 598.050 487.050 ;
        RECT 601.950 485.400 606.450 487.050 ;
        RECT 601.950 484.950 606.000 485.400 ;
        RECT 616.950 484.950 619.050 487.050 ;
        RECT 622.950 481.950 625.050 487.050 ;
        RECT 640.950 484.800 643.050 486.900 ;
        RECT 559.950 463.950 562.050 466.050 ;
        RECT 580.950 463.950 583.050 466.050 ;
        RECT 556.950 459.300 559.050 461.400 ;
        RECT 541.950 454.950 544.050 457.050 ;
        RECT 556.950 455.700 558.150 459.300 ;
        RECT 556.950 453.600 559.050 455.700 ;
        RECT 541.950 448.950 544.050 451.050 ;
        RECT 542.400 439.050 543.450 448.950 ;
        RECT 547.950 445.950 550.050 448.050 ;
        RECT 535.950 436.500 538.050 438.600 ;
        RECT 541.950 436.950 544.050 439.050 ;
        RECT 508.950 430.950 511.050 433.050 ;
        RECT 460.950 421.950 463.050 424.050 ;
        RECT 499.950 422.400 502.050 424.500 ;
        RECT 437.400 420.000 441.450 420.450 ;
        RECT 436.950 419.400 441.450 420.000 ;
        RECT 436.950 415.950 439.050 419.400 ;
        RECT 454.950 419.100 457.050 421.200 ;
        RECT 454.950 415.800 457.050 417.900 ;
        RECT 433.950 409.950 436.050 412.050 ;
        RECT 455.400 411.450 456.450 415.800 ;
        RECT 452.400 411.000 456.450 411.450 ;
        RECT 451.950 410.400 456.450 411.000 ;
        RECT 434.400 403.050 435.450 409.950 ;
        RECT 445.950 406.950 448.050 409.050 ;
        RECT 451.950 406.950 454.050 410.400 ;
        RECT 457.950 409.950 460.050 415.050 ;
        RECT 469.950 412.950 472.050 415.050 ;
        RECT 484.950 412.950 487.050 418.050 ;
        RECT 490.950 415.950 493.050 418.050 ;
        RECT 433.950 400.950 436.050 403.050 ;
        RECT 446.400 399.450 447.450 406.950 ;
        RECT 452.400 400.050 453.450 406.950 ;
        RECT 443.400 398.400 447.450 399.450 ;
        RECT 430.950 370.950 433.050 376.050 ;
        RECT 443.400 373.050 444.450 398.400 ;
        RECT 451.950 397.950 454.050 400.050 ;
        RECT 470.400 397.050 471.450 412.950 ;
        RECT 478.950 409.950 484.050 412.050 ;
        RECT 487.950 406.950 490.050 412.050 ;
        RECT 491.400 400.050 492.450 415.950 ;
        RECT 500.700 402.600 501.900 422.400 ;
        RECT 511.950 421.950 514.050 424.050 ;
        RECT 520.950 422.400 523.050 424.500 ;
        RECT 512.400 415.050 513.450 421.950 ;
        RECT 505.950 409.950 508.050 415.050 ;
        RECT 511.950 412.950 514.050 415.050 ;
        RECT 520.950 407.400 522.150 422.400 ;
        RECT 548.400 421.050 549.450 445.950 ;
        RECT 556.950 438.600 558.150 453.600 ;
        RECT 581.400 451.050 582.450 463.950 ;
        RECT 641.400 457.050 642.450 484.800 ;
        RECT 640.950 454.950 643.050 457.050 ;
        RECT 574.950 448.950 577.050 451.050 ;
        RECT 580.950 448.950 583.050 451.050 ;
        RECT 628.950 448.950 634.050 451.050 ;
        RECT 637.950 448.950 640.050 454.050 ;
        RECT 559.950 442.950 565.050 445.050 ;
        RECT 571.950 442.950 574.050 445.050 ;
        RECT 556.950 436.500 559.050 438.600 ;
        RECT 547.950 418.950 550.050 421.050 ;
        RECT 562.950 418.950 565.050 421.050 ;
        RECT 523.950 412.950 526.050 418.050 ;
        RECT 541.950 412.950 544.050 418.050 ;
        RECT 553.950 412.950 559.050 415.050 ;
        RECT 520.950 405.300 523.050 407.400 ;
        RECT 538.950 406.950 541.050 412.050 ;
        RECT 544.950 406.950 547.050 412.050 ;
        RECT 499.950 400.500 502.050 402.600 ;
        RECT 520.950 401.700 522.150 405.300 ;
        RECT 490.950 397.950 493.050 400.050 ;
        RECT 511.950 397.950 514.050 400.050 ;
        RECT 520.950 399.600 523.050 401.700 ;
        RECT 469.950 394.950 472.050 397.050 ;
        RECT 470.400 385.050 471.450 394.950 ;
        RECT 469.950 382.950 472.050 385.050 ;
        RECT 481.950 380.400 484.050 382.500 ;
        RECT 502.950 381.300 505.050 383.400 ;
        RECT 436.950 370.950 439.050 373.050 ;
        RECT 442.950 370.950 445.050 373.050 ;
        RECT 460.950 370.950 463.050 373.050 ;
        RECT 466.950 370.950 469.050 373.050 ;
        RECT 472.950 370.950 475.050 373.050 ;
        RECT 428.400 368.400 432.450 369.450 ;
        RECT 412.950 358.500 415.050 360.600 ;
        RECT 421.800 358.950 423.900 361.050 ;
        RECT 425.100 358.950 427.200 361.050 ;
        RECT 415.950 344.400 418.050 346.500 ;
        RECT 416.700 324.600 417.900 344.400 ;
        RECT 421.950 340.950 424.050 343.050 ;
        RECT 422.400 334.050 423.450 340.950 ;
        RECT 431.400 340.050 432.450 368.400 ;
        RECT 433.950 364.950 436.050 370.050 ;
        RECT 437.400 367.050 438.450 370.950 ;
        RECT 451.950 367.950 457.050 370.050 ;
        RECT 436.950 364.950 439.050 367.050 ;
        RECT 461.400 364.050 462.450 370.950 ;
        RECT 463.950 364.950 466.050 370.050 ;
        RECT 442.950 358.950 445.050 364.050 ;
        RECT 460.950 361.950 463.050 364.050 ;
        RECT 461.400 355.050 462.450 361.950 ;
        RECT 460.950 352.950 463.050 355.050 ;
        RECT 436.950 344.400 439.050 346.500 ;
        RECT 430.950 337.950 433.050 340.050 ;
        RECT 427.950 334.950 430.050 337.050 ;
        RECT 421.950 331.950 424.050 334.050 ;
        RECT 428.400 331.050 429.450 334.950 ;
        RECT 427.950 328.950 430.050 331.050 ;
        RECT 415.950 322.500 418.050 324.600 ;
        RECT 428.400 316.050 429.450 328.950 ;
        RECT 431.400 319.050 432.450 337.950 ;
        RECT 436.950 329.400 438.150 344.400 ;
        RECT 454.950 343.950 457.050 346.050 ;
        RECT 439.950 339.450 444.000 340.050 ;
        RECT 439.950 337.950 444.450 339.450 ;
        RECT 445.950 337.950 448.050 343.050 ;
        RECT 443.400 331.050 444.450 337.950 ;
        RECT 455.400 334.050 456.450 343.950 ;
        RECT 457.950 334.950 460.050 340.050 ;
        RECT 464.400 337.050 465.450 364.950 ;
        RECT 467.400 352.050 468.450 370.950 ;
        RECT 473.400 367.050 474.450 370.950 ;
        RECT 472.950 364.950 475.050 367.050 ;
        RECT 482.700 360.600 483.900 380.400 ;
        RECT 493.950 376.950 496.050 379.050 ;
        RECT 502.950 377.700 504.150 381.300 ;
        RECT 487.950 370.950 493.050 373.050 ;
        RECT 494.400 370.050 495.450 376.950 ;
        RECT 502.950 375.600 505.050 377.700 ;
        RECT 493.950 367.950 496.050 370.050 ;
        RECT 496.950 364.950 499.050 367.050 ;
        RECT 481.950 358.500 484.050 360.600 ;
        RECT 484.950 352.950 487.050 355.050 ;
        RECT 466.950 349.950 469.050 352.050 ;
        RECT 478.950 349.950 481.050 352.050 ;
        RECT 466.950 340.950 469.050 346.050 ;
        RECT 479.400 343.050 480.450 349.950 ;
        RECT 478.950 340.950 481.050 343.050 ;
        RECT 463.950 334.950 466.050 337.050 ;
        RECT 475.950 334.950 481.050 337.050 ;
        RECT 454.950 331.950 457.050 334.050 ;
        RECT 460.950 331.950 463.050 334.050 ;
        RECT 436.950 327.300 439.050 329.400 ;
        RECT 442.950 328.950 445.050 331.050 ;
        RECT 436.950 323.700 438.150 327.300 ;
        RECT 436.950 321.600 439.050 323.700 ;
        RECT 448.950 322.950 451.050 325.050 ;
        RECT 430.950 316.950 433.050 319.050 ;
        RECT 436.950 316.950 439.050 319.050 ;
        RECT 427.950 313.950 430.050 316.050 ;
        RECT 424.950 301.950 427.050 304.050 ;
        RECT 415.950 295.950 418.050 298.050 ;
        RECT 409.950 292.950 415.050 295.050 ;
        RECT 416.400 277.050 417.450 295.950 ;
        RECT 418.950 292.950 421.050 295.050 ;
        RECT 425.400 294.450 426.450 301.950 ;
        RECT 427.950 295.950 430.050 301.050 ;
        RECT 433.950 295.950 436.050 298.050 ;
        RECT 425.400 294.000 429.450 294.450 ;
        RECT 425.400 293.400 430.050 294.000 ;
        RECT 419.400 283.050 420.450 292.950 ;
        RECT 427.950 289.950 430.050 293.400 ;
        RECT 421.950 286.950 427.050 289.050 ;
        RECT 430.950 286.950 433.050 289.050 ;
        RECT 418.950 280.950 421.050 283.050 ;
        RECT 424.950 280.950 427.050 283.050 ;
        RECT 415.950 274.950 418.050 277.050 ;
        RECT 406.950 262.950 409.050 265.050 ;
        RECT 403.950 259.950 406.050 262.050 ;
        RECT 409.950 259.950 412.050 262.050 ;
        RECT 391.950 250.950 394.050 256.050 ;
        RECT 394.950 253.950 397.050 256.050 ;
        RECT 404.400 253.050 405.450 259.950 ;
        RECT 406.950 253.950 409.050 256.050 ;
        RECT 403.950 250.950 406.050 253.050 ;
        RECT 382.950 244.500 385.050 246.600 ;
        RECT 407.400 235.050 408.450 253.950 ;
        RECT 410.400 238.050 411.450 259.950 ;
        RECT 415.950 256.950 418.050 262.050 ;
        RECT 425.400 256.050 426.450 280.950 ;
        RECT 427.950 268.950 430.050 271.050 ;
        RECT 428.400 262.050 429.450 268.950 ;
        RECT 427.950 259.950 430.050 262.050 ;
        RECT 427.950 256.050 430.050 256.200 ;
        RECT 418.950 250.950 421.050 256.050 ;
        RECT 424.950 254.100 430.050 256.050 ;
        RECT 424.950 253.950 429.000 254.100 ;
        RECT 421.950 238.950 424.050 241.050 ;
        RECT 409.950 235.950 412.050 238.050 ;
        RECT 406.950 232.950 409.050 235.050 ;
        RECT 370.950 226.950 373.050 229.050 ;
        RECT 370.950 220.950 373.050 223.050 ;
        RECT 371.400 217.050 372.450 220.950 ;
        RECT 370.950 214.950 373.050 217.050 ;
        RECT 373.950 214.950 376.050 217.050 ;
        RECT 376.950 216.450 381.000 217.050 ;
        RECT 376.950 214.950 381.450 216.450 ;
        RECT 385.950 214.950 388.050 217.050 ;
        RECT 397.950 214.950 400.050 217.050 ;
        RECT 374.400 211.050 375.450 214.950 ;
        RECT 380.400 211.050 381.450 214.950 ;
        RECT 367.950 208.950 370.050 211.050 ;
        RECT 373.950 208.950 376.050 211.050 ;
        RECT 379.950 208.950 382.050 211.050 ;
        RECT 361.950 188.400 364.050 190.500 ;
        RECT 368.400 190.050 369.450 208.950 ;
        RECT 386.400 208.050 387.450 214.950 ;
        RECT 398.400 211.050 399.450 214.950 ;
        RECT 407.400 211.050 408.450 232.950 ;
        RECT 415.950 214.950 421.050 217.050 ;
        RECT 422.400 214.050 423.450 238.950 ;
        RECT 425.400 223.050 426.450 253.950 ;
        RECT 427.950 250.800 430.050 252.900 ;
        RECT 428.400 238.050 429.450 250.800 ;
        RECT 431.400 247.050 432.450 286.950 ;
        RECT 434.400 286.050 435.450 295.950 ;
        RECT 433.950 283.950 436.050 286.050 ;
        RECT 437.400 279.450 438.450 316.950 ;
        RECT 439.950 310.950 442.050 313.050 ;
        RECT 440.400 289.050 441.450 310.950 ;
        RECT 442.950 292.950 448.050 295.050 ;
        RECT 440.400 287.400 445.050 289.050 ;
        RECT 441.000 286.950 445.050 287.400 ;
        RECT 434.400 278.400 438.450 279.450 ;
        RECT 430.950 244.950 433.050 247.050 ;
        RECT 434.400 241.050 435.450 278.400 ;
        RECT 436.950 262.950 439.050 268.050 ;
        RECT 443.400 267.450 444.450 286.950 ;
        RECT 443.400 266.400 447.450 267.450 ;
        RECT 442.950 262.950 445.050 265.050 ;
        RECT 436.950 253.950 442.050 256.050 ;
        RECT 433.950 238.950 436.050 241.050 ;
        RECT 427.800 235.950 429.900 238.050 ;
        RECT 431.100 235.950 433.200 238.050 ;
        RECT 424.950 220.950 427.050 223.050 ;
        RECT 421.950 211.950 424.050 214.050 ;
        RECT 397.950 208.950 400.050 211.050 ;
        RECT 400.950 208.950 403.050 211.050 ;
        RECT 406.950 208.950 409.050 211.050 ;
        RECT 409.950 208.950 415.050 211.050 ;
        RECT 385.950 205.950 388.050 208.050 ;
        RECT 388.950 190.950 391.050 193.050 ;
        RECT 355.950 181.950 358.050 184.050 ;
        RECT 358.950 181.950 361.050 184.050 ;
        RECT 352.950 166.950 355.050 169.050 ;
        RECT 343.950 160.950 346.050 163.050 ;
        RECT 356.400 142.050 357.450 181.950 ;
        RECT 359.400 178.050 360.450 181.950 ;
        RECT 358.950 175.950 361.050 178.050 ;
        RECT 362.850 173.400 364.050 188.400 ;
        RECT 367.950 187.950 370.050 190.050 ;
        RECT 382.950 188.400 385.050 190.500 ;
        RECT 376.950 181.950 379.050 184.050 ;
        RECT 370.950 178.950 376.050 181.050 ;
        RECT 377.400 178.050 378.450 181.950 ;
        RECT 376.950 175.950 379.050 178.050 ;
        RECT 361.950 171.300 364.050 173.400 ;
        RECT 362.850 167.700 364.050 171.300 ;
        RECT 383.100 168.600 384.300 188.400 ;
        RECT 361.950 165.600 364.050 167.700 ;
        RECT 382.950 166.500 385.050 168.600 ;
        RECT 389.400 148.050 390.450 190.950 ;
        RECT 391.950 175.950 394.050 181.050 ;
        RECT 401.400 178.050 402.450 208.950 ;
        RECT 422.400 193.050 423.450 211.950 ;
        RECT 428.400 211.050 429.450 235.950 ;
        RECT 427.950 208.950 430.050 211.050 ;
        RECT 421.950 190.950 424.050 193.050 ;
        RECT 409.950 184.950 412.050 187.050 ;
        RECT 403.950 181.950 409.050 184.050 ;
        RECT 400.950 175.950 403.050 178.050 ;
        RECT 403.950 175.950 409.050 178.050 ;
        RECT 410.400 172.050 411.450 184.950 ;
        RECT 421.950 181.950 427.050 184.050 ;
        RECT 412.950 178.950 415.050 181.050 ;
        RECT 409.950 169.950 412.050 172.050 ;
        RECT 394.950 148.950 397.050 151.050 ;
        RECT 388.950 145.950 391.050 148.050 ;
        RECT 395.400 145.050 396.450 148.950 ;
        RECT 403.950 146.400 406.050 148.500 ;
        RECT 394.950 142.950 397.050 145.050 ;
        RECT 331.950 139.950 334.050 142.050 ;
        RECT 337.950 139.950 340.050 142.050 ;
        RECT 348.000 141.450 352.050 142.050 ;
        RECT 347.400 139.950 352.050 141.450 ;
        RECT 355.950 139.950 358.050 142.050 ;
        RECT 388.950 139.950 391.050 142.050 ;
        RECT 397.950 139.950 400.050 142.050 ;
        RECT 319.950 136.950 322.050 139.050 ;
        RECT 325.950 136.950 328.050 139.050 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 307.950 130.950 310.050 133.050 ;
        RECT 322.950 130.950 325.050 136.050 ;
        RECT 308.400 103.050 309.450 130.950 ;
        RECT 326.400 124.050 327.450 136.950 ;
        RECT 332.400 136.050 333.450 139.950 ;
        RECT 331.950 133.950 334.050 136.050 ;
        RECT 338.400 124.050 339.450 139.950 ;
        RECT 347.400 136.050 348.450 139.950 ;
        RECT 367.950 139.050 370.050 139.200 ;
        RECT 346.950 133.950 349.050 136.050 ;
        RECT 361.950 133.950 364.050 139.050 ;
        RECT 367.950 137.100 373.050 139.050 ;
        RECT 369.000 136.950 373.050 137.100 ;
        RECT 376.950 136.950 382.050 139.050 ;
        RECT 367.950 130.950 370.050 135.900 ;
        RECT 382.950 133.950 385.050 139.050 ;
        RECT 389.400 136.050 390.450 139.950 ;
        RECT 388.950 133.950 391.050 136.050 ;
        RECT 325.950 121.950 328.050 124.050 ;
        RECT 337.950 121.950 340.050 124.050 ;
        RECT 322.950 112.950 325.050 115.050 ;
        RECT 313.950 103.950 316.050 109.050 ;
        RECT 316.950 103.950 322.050 106.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 323.400 100.050 324.450 112.950 ;
        RECT 337.950 109.950 340.050 112.050 ;
        RECT 334.950 103.950 337.050 106.050 ;
        RECT 289.950 94.950 292.050 100.050 ;
        RECT 298.950 97.950 301.050 100.050 ;
        RECT 301.950 94.950 304.050 100.050 ;
        RECT 322.950 97.950 325.050 100.050 ;
        RECT 328.950 97.950 331.050 103.050 ;
        RECT 319.950 88.950 322.050 91.050 ;
        RECT 286.950 70.950 289.050 73.050 ;
        RECT 301.950 70.950 304.050 73.050 ;
        RECT 247.950 63.600 250.050 65.700 ;
        RECT 277.950 64.950 280.050 67.050 ;
        RECT 283.950 64.950 286.050 67.050 ;
        RECT 232.950 58.950 235.050 61.050 ;
        RECT 241.950 58.950 244.050 61.050 ;
        RECT 238.950 55.950 241.050 58.050 ;
        RECT 239.400 52.050 240.450 55.950 ;
        RECT 232.950 49.950 235.050 52.050 ;
        RECT 238.950 49.950 241.050 52.050 ;
        RECT 226.950 46.500 229.050 48.600 ;
        RECT 208.950 43.950 211.050 46.050 ;
        RECT 199.950 25.950 202.050 28.050 ;
        RECT 178.950 24.450 181.050 25.050 ;
        RECT 184.950 24.450 187.050 25.050 ;
        RECT 178.950 23.400 187.050 24.450 ;
        RECT 178.950 22.950 181.050 23.400 ;
        RECT 184.950 22.950 187.050 23.400 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 148.950 16.950 151.050 22.050 ;
        RECT 166.950 20.100 169.050 22.200 ;
        RECT 160.950 16.950 166.050 19.050 ;
        RECT 168.000 18.900 172.050 19.050 ;
        RECT 166.950 16.950 172.050 18.900 ;
        RECT 175.950 16.950 178.050 19.050 ;
        RECT 181.950 16.950 184.050 22.050 ;
        RECT 202.950 19.950 205.050 25.050 ;
        RECT 209.400 22.050 210.450 43.950 ;
        RECT 220.950 32.400 223.050 34.500 ;
        RECT 211.950 22.950 214.050 28.050 ;
        RECT 208.950 19.950 211.050 22.050 ;
        RECT 166.950 16.800 169.050 16.950 ;
        RECT 112.950 13.950 115.050 16.050 ;
        RECT 142.950 13.950 148.050 16.050 ;
        RECT 176.400 13.050 177.450 16.950 ;
        RECT 187.950 13.950 190.050 19.050 ;
        RECT 58.950 10.950 61.050 13.050 ;
        RECT 70.950 10.950 73.050 13.050 ;
        RECT 82.950 10.950 85.050 13.050 ;
        RECT 175.950 10.950 178.050 13.050 ;
        RECT 221.700 12.600 222.900 32.400 ;
        RECT 233.400 25.050 234.450 49.950 ;
        RECT 247.950 48.600 249.150 63.600 ;
        RECT 253.950 61.950 256.050 64.050 ;
        RECT 256.950 61.950 259.050 64.050 ;
        RECT 250.950 58.950 253.050 61.050 ;
        RECT 251.400 55.050 252.450 58.950 ;
        RECT 254.400 58.050 255.450 61.950 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 250.950 52.950 253.050 55.050 ;
        RECT 247.950 46.500 250.050 48.600 ;
        RECT 257.400 40.050 258.450 61.950 ;
        RECT 265.950 58.950 268.050 64.050 ;
        RECT 284.400 61.050 285.450 64.950 ;
        RECT 287.400 64.050 288.450 70.950 ;
        RECT 302.400 64.050 303.450 70.950 ;
        RECT 286.950 61.950 289.050 64.050 ;
        RECT 289.950 61.950 292.050 64.050 ;
        RECT 301.950 61.950 304.050 64.050 ;
        RECT 274.950 58.950 280.050 61.050 ;
        RECT 283.950 58.950 286.050 61.050 ;
        RECT 259.950 55.950 262.050 58.050 ;
        RECT 260.400 46.050 261.450 55.950 ;
        RECT 287.400 55.050 288.450 61.950 ;
        RECT 268.950 52.950 271.050 55.050 ;
        RECT 286.950 52.950 289.050 55.050 ;
        RECT 259.950 43.950 262.050 46.050 ;
        RECT 247.950 37.950 250.050 40.050 ;
        RECT 256.950 37.950 259.050 40.050 ;
        RECT 241.950 32.400 244.050 34.500 ;
        RECT 226.950 19.950 229.050 25.050 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 241.950 17.400 243.150 32.400 ;
        RECT 248.400 28.050 249.450 37.950 ;
        RECT 269.400 37.050 270.450 52.950 ;
        RECT 262.950 34.950 265.050 37.050 ;
        RECT 268.950 34.950 271.050 37.050 ;
        RECT 256.950 32.400 259.050 34.500 ;
        RECT 244.950 25.950 249.450 28.050 ;
        RECT 248.400 19.050 249.450 25.950 ;
        RECT 241.950 15.300 244.050 17.400 ;
        RECT 247.950 16.950 250.050 19.050 ;
        RECT 220.950 10.500 223.050 12.600 ;
        RECT 241.950 11.700 243.150 15.300 ;
        RECT 257.700 12.600 258.900 32.400 ;
        RECT 263.400 22.050 264.450 34.950 ;
        RECT 277.950 32.400 280.050 34.500 ;
        RECT 268.950 22.950 274.050 25.050 ;
        RECT 262.950 19.950 265.050 22.050 ;
        RECT 277.950 17.400 279.150 32.400 ;
        RECT 290.400 28.050 291.450 61.950 ;
        RECT 320.400 61.050 321.450 88.950 ;
        RECT 329.400 61.050 330.450 97.950 ;
        RECT 335.400 61.050 336.450 103.950 ;
        RECT 338.400 100.050 339.450 109.950 ;
        RECT 368.400 106.050 369.450 130.950 ;
        RECT 385.950 127.950 388.050 133.050 ;
        RECT 391.950 121.950 394.050 124.050 ;
        RECT 379.950 110.400 382.050 112.500 ;
        RECT 370.950 106.950 373.050 109.050 ;
        RECT 340.950 103.950 346.050 106.050 ;
        RECT 355.950 103.950 361.050 106.050 ;
        RECT 364.950 103.950 367.050 106.050 ;
        RECT 367.950 103.950 370.050 106.050 ;
        RECT 337.950 97.950 340.050 100.050 ;
        RECT 341.400 73.050 342.450 103.950 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 350.400 88.050 351.450 100.950 ;
        RECT 365.400 100.050 366.450 103.950 ;
        RECT 371.400 100.050 372.450 106.950 ;
        RECT 358.950 97.950 364.050 100.050 ;
        RECT 364.950 97.950 367.050 100.050 ;
        RECT 367.950 98.400 372.450 100.050 ;
        RECT 367.950 97.950 372.000 98.400 ;
        RECT 380.700 90.600 381.900 110.400 ;
        RECT 392.400 103.050 393.450 121.950 ;
        RECT 398.400 118.050 399.450 139.950 ;
        RECT 404.700 126.600 405.900 146.400 ;
        RECT 413.400 141.450 414.450 178.950 ;
        RECT 428.400 178.050 429.450 208.950 ;
        RECT 431.400 184.200 432.450 235.950 ;
        RECT 443.400 231.450 444.450 262.950 ;
        RECT 446.400 238.050 447.450 266.400 ;
        RECT 449.400 250.050 450.450 322.950 ;
        RECT 457.950 319.950 460.050 322.050 ;
        RECT 451.950 301.950 454.050 304.050 ;
        RECT 452.400 295.200 453.450 301.950 ;
        RECT 451.950 293.100 454.050 295.200 ;
        RECT 451.950 287.100 454.050 291.900 ;
        RECT 458.400 288.450 459.450 319.950 ;
        RECT 461.400 313.050 462.450 331.950 ;
        RECT 469.950 328.950 472.050 334.050 ;
        RECT 485.400 322.050 486.450 352.950 ;
        RECT 497.400 346.050 498.450 364.950 ;
        RECT 502.950 360.600 504.150 375.600 ;
        RECT 505.950 361.950 508.050 367.050 ;
        RECT 502.950 358.500 505.050 360.600 ;
        RECT 496.950 343.950 499.050 346.050 ;
        RECT 497.400 337.050 498.450 343.950 ;
        RECT 512.400 340.050 513.450 397.950 ;
        RECT 517.950 380.400 520.050 382.500 ;
        RECT 538.950 381.300 541.050 383.400 ;
        RECT 518.700 360.600 519.900 380.400 ;
        RECT 529.950 376.950 532.050 379.050 ;
        RECT 538.950 377.700 540.150 381.300 ;
        RECT 530.400 370.050 531.450 376.950 ;
        RECT 538.950 375.600 541.050 377.700 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 529.950 367.950 532.050 370.050 ;
        RECT 517.950 358.500 520.050 360.600 ;
        RECT 524.400 343.050 525.450 367.950 ;
        RECT 538.950 360.600 540.150 375.600 ;
        RECT 547.950 370.950 550.050 373.050 ;
        RECT 548.400 367.050 549.450 370.950 ;
        RECT 541.950 364.950 547.050 367.050 ;
        RECT 547.950 364.950 550.050 367.050 ;
        RECT 556.950 364.950 559.050 370.050 ;
        RECT 538.950 358.500 541.050 360.600 ;
        RECT 523.950 340.950 526.050 343.050 ;
        RECT 511.950 337.950 514.050 340.050 ;
        RECT 529.950 337.950 532.050 343.050 ;
        RECT 548.400 340.050 549.450 364.950 ;
        RECT 550.950 361.950 553.050 364.050 ;
        RECT 532.950 337.950 538.050 340.050 ;
        RECT 547.950 337.950 550.050 340.050 ;
        RECT 490.950 334.950 493.050 337.050 ;
        RECT 496.950 334.950 499.050 337.050 ;
        RECT 484.950 319.950 487.050 322.050 ;
        RECT 472.950 313.950 475.050 316.050 ;
        RECT 460.950 310.950 463.050 313.050 ;
        RECT 463.950 303.300 466.050 305.400 ;
        RECT 464.850 299.700 466.050 303.300 ;
        RECT 469.950 301.950 472.050 304.050 ;
        RECT 463.950 297.600 466.050 299.700 ;
        RECT 455.400 287.400 459.450 288.450 ;
        RECT 451.950 283.800 454.050 285.900 ;
        RECT 452.400 256.050 453.450 283.800 ;
        RECT 455.400 271.050 456.450 287.400 ;
        RECT 460.950 283.950 463.050 289.050 ;
        RECT 464.850 282.600 466.050 297.600 ;
        RECT 463.950 280.500 466.050 282.600 ;
        RECT 470.400 280.050 471.450 301.950 ;
        RECT 473.400 292.050 474.450 313.950 ;
        RECT 484.950 302.400 487.050 304.500 ;
        RECT 472.950 289.950 475.050 292.050 ;
        RECT 478.950 289.950 481.050 295.050 ;
        RECT 473.400 280.050 474.450 289.950 ;
        RECT 478.950 280.950 481.050 283.050 ;
        RECT 485.100 282.600 486.300 302.400 ;
        RECT 491.400 283.050 492.450 334.950 ;
        RECT 512.400 331.050 513.450 337.950 ;
        RECT 520.950 331.950 523.050 337.050 ;
        RECT 523.950 331.950 529.050 334.050 ;
        RECT 505.950 328.950 511.050 331.050 ;
        RECT 512.400 329.400 517.050 331.050 ;
        RECT 513.000 328.950 517.050 329.400 ;
        RECT 532.950 328.950 535.050 334.050 ;
        RECT 544.950 328.950 547.050 334.050 ;
        RECT 547.950 325.950 550.050 328.050 ;
        RECT 541.950 310.950 544.050 313.050 ;
        RECT 496.950 295.950 499.050 298.050 ;
        RECT 502.950 295.950 508.050 298.050 ;
        RECT 493.950 289.950 496.050 292.050 ;
        RECT 457.950 277.950 460.050 280.050 ;
        RECT 469.800 277.950 471.900 280.050 ;
        RECT 473.100 277.950 475.200 280.050 ;
        RECT 454.950 268.950 457.050 271.050 ;
        RECT 458.400 262.050 459.450 277.950 ;
        RECT 469.950 262.950 475.050 265.050 ;
        RECT 457.950 259.950 460.050 262.050 ;
        RECT 463.950 257.100 466.050 262.050 ;
        RECT 451.950 253.950 454.050 256.050 ;
        RECT 460.950 255.900 465.000 256.050 ;
        RECT 460.950 253.950 466.050 255.900 ;
        RECT 448.950 247.950 451.050 250.050 ;
        RECT 445.950 235.950 448.050 238.050 ;
        RECT 461.400 235.050 462.450 253.950 ;
        RECT 463.950 253.800 466.050 253.950 ;
        RECT 469.950 250.950 472.050 259.050 ;
        RECT 475.950 253.950 478.050 259.050 ;
        RECT 472.950 247.950 475.050 250.050 ;
        RECT 460.950 232.950 463.050 235.050 ;
        RECT 443.400 230.400 447.450 231.450 ;
        RECT 439.950 224.400 442.050 226.500 ;
        RECT 433.950 214.950 436.050 217.050 ;
        RECT 434.400 198.450 435.450 214.950 ;
        RECT 440.700 204.600 441.900 224.400 ;
        RECT 439.950 202.500 442.050 204.600 ;
        RECT 434.400 197.400 438.450 198.450 ;
        RECT 430.950 182.100 433.050 184.200 ;
        RECT 433.950 181.050 436.050 181.200 ;
        RECT 432.000 180.900 436.050 181.050 ;
        RECT 430.950 179.100 436.050 180.900 ;
        RECT 430.950 178.950 435.000 179.100 ;
        RECT 430.950 178.800 433.050 178.950 ;
        RECT 418.950 175.950 421.050 178.050 ;
        RECT 424.950 176.400 429.450 178.050 ;
        RECT 424.950 175.950 429.000 176.400 ;
        RECT 419.400 172.050 420.450 175.950 ;
        RECT 433.950 175.800 436.050 177.900 ;
        RECT 418.950 169.950 421.050 172.050 ;
        RECT 430.950 157.950 433.050 160.050 ;
        RECT 431.400 151.050 432.450 157.950 ;
        RECT 424.950 147.300 427.050 149.400 ;
        RECT 430.950 148.950 433.050 151.050 ;
        RECT 424.950 143.700 426.150 147.300 ;
        RECT 424.950 141.600 427.050 143.700 ;
        RECT 413.400 140.400 417.450 141.450 ;
        RECT 409.950 139.050 412.050 139.200 ;
        RECT 409.950 138.600 414.000 139.050 ;
        RECT 409.950 137.100 414.450 138.600 ;
        RECT 411.000 136.950 414.450 137.100 ;
        RECT 409.950 133.800 412.050 135.900 ;
        RECT 403.950 124.500 406.050 126.600 ;
        RECT 397.950 115.950 400.050 118.050 ;
        RECT 406.950 115.950 409.050 118.050 ;
        RECT 400.950 110.400 403.050 112.500 ;
        RECT 385.950 97.950 388.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 379.950 88.500 382.050 90.600 ;
        RECT 349.950 85.950 352.050 88.050 ;
        RECT 392.400 76.050 393.450 100.950 ;
        RECT 400.950 95.400 402.150 110.400 ;
        RECT 403.950 103.950 406.050 106.050 ;
        RECT 404.400 100.050 405.450 103.950 ;
        RECT 403.950 97.950 406.050 100.050 ;
        RECT 400.950 93.300 403.050 95.400 ;
        RECT 400.950 89.700 402.150 93.300 ;
        RECT 400.950 87.600 403.050 89.700 ;
        RECT 379.950 73.950 382.050 76.050 ;
        RECT 391.950 73.950 394.050 76.050 ;
        RECT 397.950 73.950 400.050 76.050 ;
        RECT 340.950 70.950 343.050 73.050 ;
        RECT 367.950 68.400 370.050 70.500 ;
        RECT 292.950 55.950 295.050 61.050 ;
        RECT 313.950 55.950 316.050 61.050 ;
        RECT 319.950 58.950 322.050 61.050 ;
        RECT 328.950 58.950 331.050 61.050 ;
        RECT 335.400 59.400 340.050 61.050 ;
        RECT 336.000 58.950 340.050 59.400 ;
        RECT 343.950 58.950 346.050 64.050 ;
        RECT 349.950 58.950 352.050 61.050 ;
        RECT 355.950 58.950 358.050 61.050 ;
        RECT 310.950 52.950 313.050 55.050 ;
        RECT 316.950 52.950 319.050 55.050 ;
        RECT 322.950 52.950 325.050 58.050 ;
        RECT 350.400 55.050 351.450 58.950 ;
        RECT 356.400 55.050 357.450 58.950 ;
        RECT 337.950 52.950 343.050 55.050 ;
        RECT 346.950 53.400 351.450 55.050 ;
        RECT 346.950 52.950 351.000 53.400 ;
        RECT 355.800 52.950 357.900 55.050 ;
        RECT 292.950 43.950 295.050 46.050 ;
        RECT 293.400 28.050 294.450 43.950 ;
        RECT 311.400 34.050 312.450 52.950 ;
        RECT 317.400 37.050 318.450 52.950 ;
        RECT 323.400 46.050 324.450 52.950 ;
        RECT 343.950 49.950 346.050 52.050 ;
        RECT 358.950 49.950 361.050 55.050 ;
        RECT 322.950 43.950 325.050 46.050 ;
        RECT 316.950 34.950 319.050 37.050 ;
        RECT 304.950 31.950 307.050 34.050 ;
        RECT 310.950 31.950 313.050 34.050 ;
        RECT 322.950 31.950 325.050 34.050 ;
        RECT 331.950 32.400 334.050 34.500 ;
        RECT 305.400 28.050 306.450 31.950 ;
        RECT 313.950 28.950 316.050 31.050 ;
        RECT 280.950 25.950 286.050 28.050 ;
        RECT 289.950 25.950 292.050 28.050 ;
        RECT 292.950 25.950 295.050 28.050 ;
        RECT 298.950 25.950 301.050 28.050 ;
        RECT 304.950 25.950 307.050 28.050 ;
        RECT 290.400 22.050 291.450 25.950 ;
        RECT 289.950 19.950 292.050 22.050 ;
        RECT 292.950 19.950 298.050 22.050 ;
        RECT 277.950 15.300 280.050 17.400 ;
        RECT 241.950 9.600 244.050 11.700 ;
        RECT 256.950 10.500 259.050 12.600 ;
        RECT 277.950 11.700 279.150 15.300 ;
        RECT 277.950 9.600 280.050 11.700 ;
        RECT 299.400 10.050 300.450 25.950 ;
        RECT 314.400 22.050 315.450 28.950 ;
        RECT 316.950 22.950 319.050 28.050 ;
        RECT 301.950 16.950 304.050 22.050 ;
        RECT 313.950 19.950 316.050 22.050 ;
        RECT 317.400 16.050 318.450 22.950 ;
        RECT 323.400 22.050 324.450 31.950 ;
        RECT 325.950 25.950 331.050 28.050 ;
        RECT 322.950 19.950 325.050 22.050 ;
        RECT 332.850 17.400 334.050 32.400 ;
        RECT 344.400 25.050 345.450 49.950 ;
        RECT 368.700 48.600 369.900 68.400 ;
        RECT 373.950 58.950 376.050 64.050 ;
        RECT 380.400 58.050 381.450 73.950 ;
        RECT 388.950 69.300 391.050 71.400 ;
        RECT 388.950 65.700 390.150 69.300 ;
        RECT 388.950 63.600 391.050 65.700 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 388.950 48.600 390.150 63.600 ;
        RECT 394.950 61.950 397.050 64.050 ;
        RECT 395.400 55.050 396.450 61.950 ;
        RECT 391.950 52.950 397.050 55.050 ;
        RECT 367.950 46.500 370.050 48.600 ;
        RECT 388.950 46.500 391.050 48.600 ;
        RECT 373.950 40.950 376.050 43.050 ;
        RECT 367.950 34.950 370.050 37.050 ;
        RECT 352.950 32.400 355.050 34.500 ;
        RECT 340.950 22.950 346.050 25.050 ;
        RECT 337.950 19.950 340.050 22.050 ;
        RECT 316.950 13.950 319.050 16.050 ;
        RECT 331.950 15.300 334.050 17.400 ;
        RECT 332.850 11.700 334.050 15.300 ;
        RECT 338.400 13.050 339.450 19.950 ;
        RECT 346.950 16.950 349.050 22.050 ;
        RECT 298.950 7.950 301.050 10.050 ;
        RECT 331.950 9.600 334.050 11.700 ;
        RECT 337.950 10.950 340.050 13.050 ;
        RECT 353.100 12.600 354.300 32.400 ;
        RECT 361.950 25.950 364.050 28.050 ;
        RECT 362.400 22.050 363.450 25.950 ;
        RECT 361.950 19.950 364.050 22.050 ;
        RECT 364.950 13.950 367.050 16.050 ;
        RECT 352.950 10.500 355.050 12.600 ;
        RECT 365.400 10.050 366.450 13.950 ;
        RECT 364.950 7.950 367.050 10.050 ;
        RECT 368.400 7.050 369.450 34.950 ;
        RECT 374.400 28.050 375.450 40.950 ;
        RECT 379.950 31.950 382.050 34.050 ;
        RECT 385.950 32.400 388.050 34.500 ;
        RECT 373.950 25.950 376.050 28.050 ;
        RECT 380.400 22.050 381.450 31.950 ;
        RECT 370.950 19.950 373.050 22.050 ;
        RECT 376.950 19.950 382.050 22.050 ;
        RECT 371.400 13.050 372.450 19.950 ;
        RECT 370.950 10.950 373.050 13.050 ;
        RECT 386.700 12.600 387.900 32.400 ;
        RECT 391.950 28.950 394.050 31.050 ;
        RECT 392.400 22.050 393.450 28.950 ;
        RECT 398.400 25.050 399.450 73.950 ;
        RECT 407.400 70.050 408.450 115.950 ;
        RECT 406.950 67.950 409.050 70.050 ;
        RECT 406.950 58.950 409.050 64.050 ;
        RECT 410.400 58.200 411.450 133.800 ;
        RECT 413.400 130.050 414.450 136.950 ;
        RECT 416.400 136.050 417.450 140.400 ;
        RECT 415.950 133.950 418.050 136.050 ;
        RECT 412.950 127.950 415.050 130.050 ;
        RECT 416.400 124.050 417.450 133.950 ;
        RECT 424.950 126.600 426.150 141.600 ;
        RECT 431.400 133.050 432.450 148.950 ;
        RECT 434.400 133.200 435.450 175.800 ;
        RECT 437.400 139.050 438.450 197.400 ;
        RECT 446.400 148.050 447.450 230.400 ;
        RECT 448.950 223.950 451.050 226.050 ;
        RECT 460.950 225.300 463.050 227.400 ;
        RECT 449.400 217.050 450.450 223.950 ;
        RECT 460.950 221.700 462.150 225.300 ;
        RECT 460.950 219.600 463.050 221.700 ;
        RECT 448.950 214.950 451.050 217.050 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 452.400 205.050 453.450 211.950 ;
        RECT 451.950 202.950 454.050 205.050 ;
        RECT 460.950 204.600 462.150 219.600 ;
        RECT 466.950 217.950 469.050 220.050 ;
        RECT 467.400 211.050 468.450 217.950 ;
        RECT 463.950 209.400 468.450 211.050 ;
        RECT 463.950 208.950 468.000 209.400 ;
        RECT 460.950 202.500 463.050 204.600 ;
        RECT 451.950 187.950 454.050 190.050 ;
        RECT 448.950 157.950 451.050 160.050 ;
        RECT 445.950 145.950 448.050 148.050 ;
        RECT 436.950 136.950 439.050 139.050 ;
        RECT 442.950 136.950 445.050 142.050 ;
        RECT 449.400 139.050 450.450 157.950 ;
        RECT 452.400 157.050 453.450 187.950 ;
        RECT 473.400 166.050 474.450 247.950 ;
        RECT 479.400 216.450 480.450 280.950 ;
        RECT 484.950 280.500 487.050 282.600 ;
        RECT 490.950 280.950 493.050 283.050 ;
        RECT 494.400 264.450 495.450 289.950 ;
        RECT 497.400 277.050 498.450 295.950 ;
        RECT 496.950 274.950 499.050 277.050 ;
        RECT 497.400 267.450 498.450 274.950 ;
        RECT 499.950 267.450 502.050 268.050 ;
        RECT 497.400 266.400 502.050 267.450 ;
        RECT 499.950 265.950 502.050 266.400 ;
        RECT 491.400 263.400 495.450 264.450 ;
        RECT 491.400 256.050 492.450 263.400 ;
        RECT 500.400 262.200 501.450 265.950 ;
        RECT 493.950 259.950 496.050 262.050 ;
        RECT 499.950 260.100 502.050 262.200 ;
        RECT 506.400 262.050 507.450 295.950 ;
        RECT 523.950 292.950 526.050 298.050 ;
        RECT 529.950 294.450 534.000 295.050 ;
        RECT 529.950 292.950 534.450 294.450 ;
        RECT 535.950 292.950 541.050 295.050 ;
        RECT 517.950 286.950 520.050 292.050 ;
        RECT 526.950 289.950 529.050 292.050 ;
        RECT 533.400 291.450 534.450 292.950 ;
        RECT 542.400 292.050 543.450 310.950 ;
        RECT 548.400 292.050 549.450 325.950 ;
        RECT 551.400 310.050 552.450 361.950 ;
        RECT 556.950 344.400 559.050 346.500 ;
        RECT 557.700 324.600 558.900 344.400 ;
        RECT 563.400 343.050 564.450 418.950 ;
        RECT 572.400 415.050 573.450 442.950 ;
        RECT 571.950 409.950 574.050 415.050 ;
        RECT 575.400 400.050 576.450 448.950 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 577.950 442.950 580.050 445.050 ;
        RECT 586.950 442.950 589.050 445.050 ;
        RECT 578.400 439.050 579.450 442.950 ;
        RECT 577.950 436.950 580.050 439.050 ;
        RECT 577.950 415.950 580.050 421.050 ;
        RECT 587.400 418.050 588.450 442.950 ;
        RECT 598.950 422.400 601.050 424.500 ;
        RECT 614.400 424.050 615.450 445.950 ;
        RECT 589.950 418.950 592.050 421.050 ;
        RECT 586.950 412.950 589.050 418.050 ;
        RECT 577.950 409.950 583.050 412.050 ;
        RECT 574.950 397.950 577.050 400.050 ;
        RECT 583.950 381.300 586.050 383.400 ;
        RECT 568.950 376.950 571.050 379.050 ;
        RECT 584.850 377.700 586.050 381.300 ;
        RECT 562.950 340.950 565.050 343.050 ;
        RECT 569.400 337.050 570.450 376.950 ;
        RECT 583.950 375.600 586.050 377.700 ;
        RECT 571.950 370.950 574.050 373.050 ;
        RECT 572.400 349.050 573.450 370.950 ;
        RECT 574.950 361.950 577.050 367.050 ;
        RECT 577.950 364.950 583.050 367.050 ;
        RECT 584.850 360.600 586.050 375.600 ;
        RECT 590.400 364.050 591.450 418.950 ;
        RECT 599.700 402.600 600.900 422.400 ;
        RECT 613.950 421.950 616.050 424.050 ;
        RECT 619.950 422.400 622.050 424.500 ;
        RECT 614.400 415.050 615.450 421.950 ;
        RECT 610.950 413.400 615.450 415.050 ;
        RECT 610.950 412.950 615.000 413.400 ;
        RECT 607.950 409.950 610.050 412.050 ;
        RECT 598.950 400.500 601.050 402.600 ;
        RECT 608.400 397.050 609.450 409.950 ;
        RECT 607.950 394.950 610.050 397.050 ;
        RECT 604.950 380.400 607.050 382.500 ;
        RECT 592.950 376.950 595.050 379.050 ;
        RECT 593.400 370.050 594.450 376.950 ;
        RECT 598.950 370.950 601.050 373.050 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 589.950 361.950 592.050 364.050 ;
        RECT 583.950 358.500 586.050 360.600 ;
        RECT 599.400 358.050 600.450 370.950 ;
        RECT 605.100 360.600 606.300 380.400 ;
        RECT 611.400 379.050 612.450 412.950 ;
        RECT 619.950 407.400 621.150 422.400 ;
        RECT 622.950 412.950 625.050 418.050 ;
        RECT 619.950 405.300 622.050 407.400 ;
        RECT 619.950 401.700 621.150 405.300 ;
        RECT 619.950 399.600 622.050 401.700 ;
        RECT 622.950 394.950 625.050 397.050 ;
        RECT 610.950 376.950 613.050 379.050 ;
        RECT 619.950 370.950 622.050 373.050 ;
        RECT 610.950 361.950 613.050 364.050 ;
        RECT 604.950 358.500 607.050 360.600 ;
        RECT 598.950 355.950 601.050 358.050 ;
        RECT 571.950 346.950 574.050 349.050 ;
        RECT 598.950 346.950 601.050 349.050 ;
        RECT 577.950 344.400 580.050 346.500 ;
        RECT 568.950 334.950 571.050 337.050 ;
        RECT 562.950 331.950 565.050 334.050 ;
        RECT 556.950 322.500 559.050 324.600 ;
        RECT 550.950 307.950 553.050 310.050 ;
        RECT 553.950 298.950 556.050 301.050 ;
        RECT 533.400 290.400 537.450 291.450 ;
        RECT 518.400 283.050 519.450 286.950 ;
        RECT 527.400 286.050 528.450 289.950 ;
        RECT 529.950 286.950 535.050 289.050 ;
        RECT 526.950 283.950 529.050 286.050 ;
        RECT 517.950 280.950 520.050 283.050 ;
        RECT 532.950 277.950 535.050 280.050 ;
        RECT 523.950 266.400 526.050 268.500 ;
        RECT 505.950 259.950 508.050 262.050 ;
        RECT 508.950 259.950 511.050 262.050 ;
        RECT 490.950 253.950 493.050 256.050 ;
        RECT 481.950 250.950 484.050 253.050 ;
        RECT 482.400 217.050 483.450 250.950 ;
        RECT 490.950 232.950 493.050 235.050 ;
        RECT 484.950 217.950 490.050 220.050 ;
        RECT 476.400 215.400 480.450 216.450 ;
        RECT 472.950 163.950 475.050 166.050 ;
        RECT 451.950 154.950 454.050 157.050 ;
        RECT 472.950 151.950 475.050 154.050 ;
        RECT 451.950 145.950 454.050 148.050 ;
        RECT 448.950 136.950 451.050 139.050 ;
        RECT 452.400 136.050 453.450 145.950 ;
        RECT 454.950 136.950 457.050 139.050 ;
        RECT 427.950 131.400 432.450 133.050 ;
        RECT 427.950 130.950 432.000 131.400 ;
        RECT 433.950 131.100 436.050 133.200 ;
        RECT 436.950 130.950 442.050 133.050 ;
        RECT 445.950 130.950 451.050 133.050 ;
        RECT 451.950 130.950 454.050 136.050 ;
        RECT 435.000 129.900 438.000 130.050 ;
        RECT 433.950 129.300 438.000 129.900 ;
        RECT 433.950 127.950 438.450 129.300 ;
        RECT 433.950 127.800 436.050 127.950 ;
        RECT 424.950 124.500 427.050 126.600 ;
        RECT 415.950 121.950 418.050 124.050 ;
        RECT 424.950 118.950 427.050 121.050 ;
        RECT 418.950 109.950 421.050 112.050 ;
        RECT 412.950 106.950 415.050 109.050 ;
        RECT 413.400 103.200 414.450 106.950 ;
        RECT 412.950 101.100 415.050 103.200 ;
        RECT 412.950 94.950 415.050 99.900 ;
        RECT 419.400 97.050 420.450 109.950 ;
        RECT 425.400 100.050 426.450 118.950 ;
        RECT 430.950 110.400 433.050 112.500 ;
        RECT 424.950 97.950 427.050 100.050 ;
        RECT 418.950 94.950 421.050 97.050 ;
        RECT 431.700 90.600 432.900 110.400 ;
        RECT 437.400 100.050 438.450 127.950 ;
        RECT 455.400 121.050 456.450 136.950 ;
        RECT 463.950 133.950 466.050 136.050 ;
        RECT 454.950 118.950 457.050 121.050 ;
        RECT 460.950 118.950 463.050 121.050 ;
        RECT 451.950 110.400 454.050 112.500 ;
        RECT 442.950 100.950 445.050 106.050 ;
        RECT 436.950 99.450 441.000 100.050 ;
        RECT 436.950 97.950 441.450 99.450 ;
        RECT 430.950 88.500 433.050 90.600 ;
        RECT 412.950 76.950 415.050 79.050 ;
        RECT 413.400 61.050 414.450 76.950 ;
        RECT 433.950 67.950 436.050 70.050 ;
        RECT 412.950 58.950 415.050 61.050 ;
        RECT 424.950 58.950 427.050 61.050 ;
        RECT 403.950 52.950 406.050 58.050 ;
        RECT 409.950 56.100 412.050 58.200 ;
        RECT 409.950 52.800 412.050 54.900 ;
        RECT 415.950 52.950 421.050 55.050 ;
        RECT 421.950 52.950 424.050 58.050 ;
        RECT 410.400 49.050 411.450 52.800 ;
        RECT 409.950 46.950 412.050 49.050 ;
        RECT 406.950 32.400 409.050 34.500 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 391.950 19.950 394.050 22.050 ;
        RECT 406.950 17.400 408.150 32.400 ;
        RECT 416.400 31.050 417.450 52.950 ;
        RECT 425.400 51.450 426.450 58.950 ;
        RECT 434.400 58.050 435.450 67.950 ;
        RECT 440.400 61.050 441.450 97.950 ;
        RECT 451.950 95.400 453.150 110.400 ;
        RECT 461.400 103.050 462.450 118.950 ;
        RECT 454.950 99.450 457.050 103.050 ;
        RECT 460.950 100.950 463.050 103.050 ;
        RECT 454.950 99.000 459.450 99.450 ;
        RECT 455.400 98.400 459.450 99.000 ;
        RECT 451.950 93.300 454.050 95.400 ;
        RECT 451.950 89.700 453.150 93.300 ;
        RECT 451.950 87.600 454.050 89.700 ;
        RECT 458.400 76.050 459.450 98.400 ;
        RECT 464.400 88.050 465.450 133.950 ;
        RECT 473.400 133.050 474.450 151.950 ;
        RECT 472.950 130.950 475.050 133.050 ;
        RECT 473.400 112.050 474.450 130.950 ;
        RECT 472.950 109.950 475.050 112.050 ;
        RECT 476.400 109.050 477.450 215.400 ;
        RECT 481.950 214.950 484.050 217.050 ;
        RECT 481.950 208.950 487.050 211.050 ;
        RECT 487.950 208.950 490.050 214.050 ;
        RECT 491.400 142.050 492.450 232.950 ;
        RECT 494.400 226.050 495.450 259.950 ;
        RECT 499.950 256.800 502.050 258.900 ;
        RECT 493.950 223.950 496.050 226.050 ;
        RECT 500.400 220.050 501.450 256.800 ;
        RECT 493.950 219.450 498.000 220.050 ;
        RECT 493.950 217.950 498.450 219.450 ;
        RECT 497.400 214.050 498.450 217.950 ;
        RECT 499.950 214.950 502.050 220.050 ;
        RECT 509.400 217.200 510.450 259.950 ;
        RECT 514.950 256.950 517.050 262.050 ;
        RECT 520.950 259.950 523.050 265.050 ;
        RECT 517.950 253.950 520.050 256.050 ;
        RECT 508.950 215.100 511.050 217.200 ;
        RECT 496.950 211.950 499.050 214.050 ;
        RECT 510.000 213.900 514.050 214.050 ;
        RECT 508.950 211.950 514.050 213.900 ;
        RECT 493.950 202.950 496.050 205.050 ;
        RECT 494.400 181.050 495.450 202.950 ;
        RECT 493.950 178.950 496.050 181.050 ;
        RECT 490.950 139.950 493.050 142.050 ;
        RECT 481.950 136.950 484.050 139.050 ;
        RECT 487.950 136.950 490.050 139.050 ;
        RECT 482.400 133.050 483.450 136.950 ;
        RECT 481.950 130.950 484.050 133.050 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 485.400 126.450 486.450 130.950 ;
        RECT 482.400 125.400 486.450 126.450 ;
        RECT 475.950 106.950 478.050 109.050 ;
        RECT 466.950 100.950 469.050 103.050 ;
        RECT 463.950 85.950 466.050 88.050 ;
        RECT 457.950 73.950 460.050 76.050 ;
        RECT 460.950 67.950 463.050 70.050 ;
        RECT 440.400 58.950 445.050 61.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 419.400 51.000 426.450 51.450 ;
        RECT 418.950 50.400 426.450 51.000 ;
        RECT 418.950 46.950 421.050 50.400 ;
        RECT 440.400 46.050 441.450 58.950 ;
        RECT 448.950 53.100 451.050 58.050 ;
        RECT 461.400 55.050 462.450 67.950 ;
        RECT 467.400 61.050 468.450 100.950 ;
        RECT 475.950 97.950 481.050 100.050 ;
        RECT 482.400 97.050 483.450 125.400 ;
        RECT 488.400 106.050 489.450 136.950 ;
        RECT 494.400 136.050 495.450 178.950 ;
        RECT 497.400 160.050 498.450 211.950 ;
        RECT 508.950 211.800 511.050 211.950 ;
        RECT 518.400 208.050 519.450 253.950 ;
        RECT 524.850 251.400 526.050 266.400 ;
        RECT 533.400 259.050 534.450 277.950 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 523.950 249.300 526.050 251.400 ;
        RECT 524.850 245.700 526.050 249.300 ;
        RECT 536.400 247.050 537.450 290.400 ;
        RECT 541.950 289.950 544.050 292.050 ;
        RECT 547.950 291.450 550.050 292.050 ;
        RECT 547.950 290.400 552.450 291.450 ;
        RECT 547.950 289.950 550.050 290.400 ;
        RECT 538.950 286.950 541.050 289.050 ;
        RECT 539.400 256.050 540.450 286.950 ;
        RECT 544.950 266.400 547.050 268.500 ;
        RECT 538.950 253.950 541.050 256.050 ;
        RECT 523.950 243.600 526.050 245.700 ;
        RECT 535.950 244.950 538.050 247.050 ;
        RECT 545.100 246.600 546.300 266.400 ;
        RECT 536.400 229.050 537.450 244.950 ;
        RECT 544.950 244.500 547.050 246.600 ;
        RECT 551.400 238.050 552.450 290.400 ;
        RECT 554.400 289.050 555.450 298.950 ;
        RECT 563.400 289.050 564.450 331.950 ;
        RECT 577.950 329.400 579.150 344.400 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 580.950 334.950 583.050 340.050 ;
        RECT 577.950 327.300 580.050 329.400 ;
        RECT 586.950 328.950 589.050 334.050 ;
        RECT 577.950 323.700 579.150 327.300 ;
        RECT 577.950 321.600 580.050 323.700 ;
        RECT 583.950 322.950 586.050 325.050 ;
        RECT 584.400 301.050 585.450 322.950 ;
        RECT 593.400 304.050 594.450 340.950 ;
        RECT 599.400 337.050 600.450 346.950 ;
        RECT 604.950 340.950 607.050 343.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 598.950 307.950 601.050 310.050 ;
        RECT 592.950 301.950 595.050 304.050 ;
        RECT 583.950 298.950 586.050 301.050 ;
        RECT 571.950 295.050 574.050 298.050 ;
        RECT 586.950 295.950 592.050 298.050 ;
        RECT 599.400 295.050 600.450 307.950 ;
        RECT 605.400 298.050 606.450 340.950 ;
        RECT 604.950 295.950 607.050 298.050 ;
        RECT 565.950 292.950 568.050 295.050 ;
        RECT 570.000 294.450 574.050 295.050 ;
        RECT 569.400 292.950 574.050 294.450 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 553.950 286.950 556.050 289.050 ;
        RECT 562.950 286.950 565.050 289.050 ;
        RECT 554.400 268.050 555.450 286.950 ;
        RECT 566.400 286.050 567.450 292.950 ;
        RECT 565.950 283.950 568.050 286.050 ;
        RECT 553.950 265.950 556.050 268.050 ;
        RECT 565.950 262.950 568.050 268.050 ;
        RECT 562.950 256.950 565.050 259.050 ;
        RECT 553.950 253.950 559.050 256.050 ;
        RECT 563.400 253.050 564.450 256.950 ;
        RECT 562.950 250.950 565.050 253.050 ;
        RECT 556.950 244.950 559.050 247.050 ;
        RECT 550.950 235.950 553.050 238.050 ;
        RECT 535.950 226.950 538.050 229.050 ;
        RECT 557.400 217.050 558.450 244.950 ;
        RECT 520.950 214.950 526.050 217.050 ;
        RECT 529.950 214.950 532.050 217.050 ;
        RECT 535.950 214.950 538.050 217.050 ;
        RECT 556.950 214.950 559.050 217.050 ;
        RECT 526.950 208.950 529.050 211.050 ;
        RECT 517.950 205.950 520.050 208.050 ;
        RECT 523.950 187.950 526.050 190.050 ;
        RECT 524.400 184.050 525.450 187.950 ;
        RECT 527.400 187.050 528.450 208.950 ;
        RECT 530.400 199.050 531.450 214.950 ;
        RECT 536.400 211.050 537.450 214.950 ;
        RECT 557.400 211.050 558.450 214.950 ;
        RECT 562.950 211.950 568.050 214.050 ;
        RECT 532.950 209.400 537.450 211.050 ;
        RECT 532.950 208.950 537.000 209.400 ;
        RECT 547.950 208.950 553.050 211.050 ;
        RECT 556.950 208.950 559.050 211.050 ;
        RECT 553.950 205.950 556.050 208.050 ;
        RECT 529.950 196.950 532.050 199.050 ;
        RECT 554.400 193.050 555.450 205.950 ;
        RECT 529.950 190.950 532.050 193.050 ;
        RECT 553.950 190.950 556.050 193.050 ;
        RECT 526.950 184.950 529.050 187.050 ;
        RECT 514.950 181.950 517.050 184.050 ;
        RECT 523.950 181.950 526.050 184.050 ;
        RECT 515.400 175.050 516.450 181.950 ;
        RECT 517.950 175.950 520.050 181.050 ;
        RECT 530.400 178.050 531.450 190.950 ;
        RECT 541.950 188.400 544.050 190.500 ;
        RECT 532.950 181.950 535.050 187.050 ;
        RECT 535.950 181.950 541.050 184.050 ;
        RECT 520.950 175.950 526.050 178.050 ;
        RECT 529.950 175.950 532.050 178.050 ;
        RECT 505.950 172.950 508.050 175.050 ;
        RECT 514.950 172.950 517.050 175.050 ;
        RECT 542.850 173.400 544.050 188.400 ;
        RECT 556.950 187.950 559.050 190.050 ;
        RECT 562.950 188.400 565.050 190.500 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 496.950 157.950 499.050 160.050 ;
        RECT 506.400 154.050 507.450 172.950 ;
        RECT 505.950 151.950 508.050 154.050 ;
        RECT 499.950 147.300 502.050 149.400 ;
        RECT 500.850 143.700 502.050 147.300 ;
        RECT 499.950 141.600 502.050 143.700 ;
        RECT 496.950 136.950 499.050 139.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 497.400 133.050 498.450 136.950 ;
        RECT 490.950 132.450 495.000 133.050 ;
        RECT 490.950 132.000 495.450 132.450 ;
        RECT 490.950 130.950 496.050 132.000 ;
        RECT 496.950 130.950 499.050 133.050 ;
        RECT 493.950 127.950 496.050 130.950 ;
        RECT 500.850 126.600 502.050 141.600 ;
        RECT 511.950 136.950 514.050 142.050 ;
        RECT 505.950 133.950 511.050 136.050 ;
        RECT 499.950 124.500 502.050 126.600 ;
        RECT 509.400 121.050 510.450 133.950 ;
        RECT 508.950 118.950 511.050 121.050 ;
        RECT 515.400 112.050 516.450 172.950 ;
        RECT 541.950 171.300 544.050 173.400 ;
        RECT 542.850 167.700 544.050 171.300 ;
        RECT 526.950 163.950 529.050 166.050 ;
        RECT 541.950 165.600 544.050 167.700 ;
        RECT 520.950 146.400 523.050 148.500 ;
        RECT 521.100 126.600 522.300 146.400 ;
        RECT 527.400 145.050 528.450 163.950 ;
        RECT 551.400 154.050 552.450 178.950 ;
        RECT 557.400 178.050 558.450 187.950 ;
        RECT 556.950 175.950 559.050 178.050 ;
        RECT 563.100 168.600 564.300 188.400 ;
        RECT 569.400 187.050 570.450 292.950 ;
        RECT 605.400 292.050 606.450 295.950 ;
        RECT 611.400 295.050 612.450 361.950 ;
        RECT 620.400 337.200 621.450 370.950 ;
        RECT 623.400 367.050 624.450 394.950 ;
        RECT 625.950 370.950 628.050 376.050 ;
        RECT 629.400 367.050 630.450 448.950 ;
        RECT 644.400 447.450 645.450 491.400 ;
        RECT 649.950 490.950 652.050 496.050 ;
        RECT 655.950 493.950 658.050 499.050 ;
        RECT 665.400 493.050 666.450 523.950 ;
        RECT 674.400 496.050 675.450 529.950 ;
        RECT 677.400 526.050 678.450 529.950 ;
        RECT 683.400 529.050 684.450 535.950 ;
        RECT 682.950 526.950 685.050 529.050 ;
        RECT 676.950 523.950 679.050 526.050 ;
        RECT 685.950 520.950 688.050 526.050 ;
        RECT 679.950 511.950 682.050 514.050 ;
        RECT 667.950 493.950 670.050 496.050 ;
        RECT 673.950 493.950 676.050 496.050 ;
        RECT 655.950 487.950 661.050 490.050 ;
        RECT 664.950 487.950 667.050 493.050 ;
        RECT 668.400 460.050 669.450 493.950 ;
        RECT 680.400 493.050 681.450 511.950 ;
        RECT 695.400 508.050 696.450 556.950 ;
        RECT 698.400 526.200 699.450 562.950 ;
        RECT 697.950 524.100 700.050 526.200 ;
        RECT 704.400 523.050 705.450 625.950 ;
        RECT 706.950 616.950 709.050 619.050 ;
        RECT 707.400 610.050 708.450 616.950 ;
        RECT 706.950 607.950 709.050 610.050 ;
        RECT 707.400 595.050 708.450 607.950 ;
        RECT 715.950 601.950 718.050 607.050 ;
        RECT 721.950 604.950 727.050 607.050 ;
        RECT 733.950 604.950 736.050 607.050 ;
        RECT 734.400 601.050 735.450 604.950 ;
        RECT 709.950 598.950 712.050 601.050 ;
        RECT 718.950 598.950 721.050 601.050 ;
        RECT 706.950 592.950 709.050 595.050 ;
        RECT 710.400 574.050 711.450 598.950 ;
        RECT 719.400 595.050 720.450 598.950 ;
        RECT 733.950 595.950 736.050 601.050 ;
        RECT 718.950 592.950 721.050 595.050 ;
        RECT 712.950 574.950 715.050 580.050 ;
        RECT 737.400 576.450 738.450 653.400 ;
        RECT 739.950 652.950 742.050 655.050 ;
        RECT 740.400 583.050 741.450 652.950 ;
        RECT 742.950 649.950 745.050 652.050 ;
        RECT 743.400 613.050 744.450 649.950 ;
        RECT 755.400 649.050 756.450 670.950 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 745.800 640.950 747.900 643.050 ;
        RECT 748.950 640.950 751.050 643.050 ;
        RECT 746.400 637.050 747.450 640.950 ;
        RECT 745.950 634.950 748.050 637.050 ;
        RECT 742.950 610.950 745.050 613.050 ;
        RECT 749.400 607.050 750.450 640.950 ;
        RECT 755.400 625.050 756.450 646.950 ;
        RECT 758.400 646.050 759.450 674.400 ;
        RECT 757.950 643.950 760.050 646.050 ;
        RECT 767.400 643.050 768.450 676.950 ;
        RECT 785.400 655.050 786.450 676.950 ;
        RECT 775.950 649.950 778.050 655.050 ;
        RECT 784.950 652.950 787.050 655.050 ;
        RECT 778.950 646.950 781.050 652.050 ;
        RECT 781.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 760.950 637.950 763.050 643.050 ;
        RECT 766.950 640.950 769.050 643.050 ;
        RECT 769.950 640.950 772.050 646.050 ;
        RECT 772.950 640.950 778.050 643.050 ;
        RECT 763.950 637.950 766.050 640.050 ;
        RECT 754.950 622.950 757.050 625.050 ;
        RECT 751.950 619.950 754.050 622.050 ;
        RECT 760.950 619.950 763.050 622.050 ;
        RECT 752.400 607.050 753.450 619.950 ;
        RECT 757.950 610.950 760.050 613.050 ;
        RECT 742.950 604.950 745.050 607.050 ;
        RECT 748.950 604.950 751.050 607.050 ;
        RECT 751.950 604.950 754.050 607.050 ;
        RECT 739.950 580.950 742.050 583.050 ;
        RECT 716.400 575.400 723.450 576.450 ;
        RECT 737.400 575.400 741.450 576.450 ;
        RECT 709.950 571.950 712.050 574.050 ;
        RECT 716.400 573.450 717.450 575.400 ;
        RECT 713.400 572.400 717.450 573.450 ;
        RECT 713.400 571.050 714.450 572.400 ;
        RECT 718.950 571.950 721.050 574.050 ;
        RECT 706.950 565.950 709.050 571.050 ;
        RECT 712.950 565.950 715.050 571.050 ;
        RECT 719.400 568.050 720.450 571.950 ;
        RECT 722.400 571.050 723.450 575.400 ;
        RECT 736.950 571.950 739.050 574.050 ;
        RECT 722.400 569.400 727.050 571.050 ;
        RECT 723.000 568.950 727.050 569.400 ;
        RECT 737.400 568.050 738.450 571.950 ;
        RECT 718.950 565.950 721.050 568.050 ;
        RECT 727.950 565.950 733.050 568.050 ;
        RECT 736.950 565.950 739.050 568.050 ;
        RECT 724.950 547.950 727.050 550.050 ;
        RECT 725.400 541.050 726.450 547.950 ;
        RECT 736.950 544.950 739.050 547.050 ;
        RECT 724.950 538.950 727.050 541.050 ;
        RECT 715.950 529.050 718.050 529.200 ;
        RECT 709.950 526.950 712.050 529.050 ;
        RECT 715.950 528.600 720.000 529.050 ;
        RECT 715.950 527.100 720.450 528.600 ;
        RECT 717.000 526.950 720.450 527.100 ;
        RECT 697.950 520.800 700.050 522.900 ;
        RECT 703.950 520.950 706.050 523.050 ;
        RECT 698.400 514.050 699.450 520.800 ;
        RECT 710.400 520.050 711.450 526.950 ;
        RECT 715.950 523.050 718.050 525.900 ;
        RECT 712.950 522.000 718.050 523.050 ;
        RECT 712.950 520.950 717.450 522.000 ;
        RECT 709.950 517.950 712.050 520.050 ;
        RECT 697.950 511.950 700.050 514.050 ;
        RECT 712.950 508.950 715.050 511.050 ;
        RECT 694.950 505.950 697.050 508.050 ;
        RECT 709.950 505.950 712.050 508.050 ;
        RECT 691.950 499.950 694.050 502.050 ;
        RECT 703.950 499.950 706.050 502.050 ;
        RECT 685.950 493.950 688.050 496.050 ;
        RECT 679.950 490.950 682.050 493.050 ;
        RECT 670.950 489.450 673.050 490.200 ;
        RECT 676.950 489.450 679.050 490.050 ;
        RECT 670.950 488.400 679.050 489.450 ;
        RECT 670.950 488.100 673.050 488.400 ;
        RECT 676.950 487.950 679.050 488.400 ;
        RECT 670.950 484.800 673.050 486.900 ;
        RECT 682.950 484.950 685.050 490.050 ;
        RECT 667.950 457.950 670.050 460.050 ;
        RECT 671.400 454.050 672.450 484.800 ;
        RECT 686.400 472.050 687.450 493.950 ;
        RECT 688.950 484.950 691.050 487.050 ;
        RECT 685.950 469.950 688.050 472.050 ;
        RECT 689.400 466.050 690.450 484.950 ;
        RECT 692.400 481.050 693.450 499.950 ;
        RECT 697.950 490.950 700.050 496.050 ;
        RECT 700.950 490.050 703.050 490.200 ;
        RECT 704.400 490.050 705.450 499.950 ;
        RECT 706.950 493.950 709.050 496.050 ;
        RECT 700.950 488.550 705.450 490.050 ;
        RECT 700.950 488.100 705.000 488.550 ;
        RECT 702.000 487.950 705.000 488.100 ;
        RECT 707.400 487.050 708.450 493.950 ;
        RECT 700.950 481.950 703.050 486.900 ;
        RECT 706.950 484.950 709.050 487.050 ;
        RECT 703.950 481.950 706.050 484.050 ;
        RECT 691.950 478.950 694.050 481.050 ;
        RECT 694.950 469.950 697.050 472.050 ;
        RECT 688.950 463.950 691.050 466.050 ;
        RECT 679.950 457.950 682.050 460.050 ;
        RECT 680.400 454.050 681.450 457.950 ;
        RECT 695.400 457.050 696.450 469.950 ;
        RECT 649.950 448.950 652.050 451.050 ;
        RECT 661.950 449.100 664.050 454.050 ;
        RECT 667.950 453.000 672.450 454.050 ;
        RECT 667.950 451.950 673.050 453.000 ;
        RECT 679.950 451.950 682.050 454.050 ;
        RECT 685.950 451.950 688.050 457.050 ;
        RECT 694.950 454.950 697.050 457.050 ;
        RECT 670.950 448.950 673.050 451.950 ;
        RECT 691.950 448.950 697.050 451.050 ;
        RECT 644.400 446.400 648.450 447.450 ;
        RECT 634.950 442.950 637.050 445.050 ;
        RECT 640.950 442.950 646.050 445.050 ;
        RECT 635.400 418.200 636.450 442.950 ;
        RECT 647.400 427.050 648.450 446.400 ;
        RECT 646.950 424.950 649.050 427.050 ;
        RECT 650.400 421.050 651.450 448.950 ;
        RECT 661.950 445.800 664.050 447.900 ;
        RECT 655.950 439.950 658.050 445.050 ;
        RECT 662.400 442.050 663.450 445.800 ;
        RECT 688.950 442.950 691.050 448.050 ;
        RECT 694.950 442.950 700.050 445.050 ;
        RECT 661.950 439.950 664.050 442.050 ;
        RECT 658.950 424.950 661.050 427.050 ;
        RECT 637.950 418.950 640.050 421.050 ;
        RECT 649.950 418.950 652.050 421.050 ;
        RECT 634.950 416.100 637.050 418.200 ;
        RECT 634.950 412.800 637.050 414.900 ;
        RECT 635.400 370.050 636.450 412.800 ;
        RECT 638.400 412.050 639.450 418.950 ;
        RECT 640.950 415.950 643.050 418.050 ;
        RECT 646.950 417.450 651.000 418.050 ;
        RECT 646.950 415.950 651.450 417.450 ;
        RECT 641.400 412.050 642.450 415.950 ;
        RECT 650.400 412.050 651.450 415.950 ;
        RECT 637.950 409.950 640.050 412.050 ;
        RECT 640.950 409.950 643.050 412.050 ;
        RECT 643.950 409.950 646.050 412.050 ;
        RECT 649.950 411.450 652.050 412.050 ;
        RECT 649.950 410.400 654.450 411.450 ;
        RECT 649.950 409.950 652.050 410.400 ;
        RECT 644.400 400.050 645.450 409.950 ;
        RECT 643.950 397.950 646.050 400.050 ;
        RECT 646.950 382.950 649.050 385.050 ;
        RECT 637.950 373.050 640.050 376.050 ;
        RECT 637.950 370.950 646.050 373.050 ;
        RECT 622.950 364.950 625.050 367.050 ;
        RECT 628.950 364.950 631.050 367.050 ;
        RECT 634.950 364.950 637.050 370.050 ;
        RECT 613.950 334.950 616.050 337.050 ;
        RECT 619.950 335.100 622.050 337.200 ;
        RECT 614.400 331.050 615.450 334.950 ;
        RECT 629.400 334.050 630.450 364.950 ;
        RECT 631.950 343.950 634.050 346.050 ;
        RECT 613.950 328.950 616.050 331.050 ;
        RECT 619.950 328.950 622.050 333.900 ;
        RECT 628.950 331.950 631.050 334.050 ;
        RECT 632.400 331.050 633.450 343.950 ;
        RECT 647.400 337.050 648.450 382.950 ;
        RECT 653.400 370.050 654.450 410.400 ;
        RECT 659.400 391.050 660.450 424.950 ;
        RECT 670.950 422.400 673.050 424.500 ;
        RECT 661.950 415.950 664.050 421.050 ;
        RECT 664.950 415.950 670.050 418.050 ;
        RECT 658.950 388.950 661.050 391.050 ;
        RECT 665.400 379.050 666.450 415.950 ;
        RECT 671.850 407.400 673.050 422.400 ;
        RECT 679.950 421.950 682.050 424.050 ;
        RECT 691.950 422.400 694.050 424.500 ;
        RECT 680.400 415.050 681.450 421.950 ;
        RECT 679.950 412.950 682.050 415.050 ;
        RECT 670.950 405.300 673.050 407.400 ;
        RECT 671.850 401.700 673.050 405.300 ;
        RECT 670.950 399.600 673.050 401.700 ;
        RECT 664.950 376.950 667.050 379.050 ;
        RECT 670.950 376.950 673.050 379.050 ;
        RECT 671.400 370.050 672.450 376.950 ;
        RECT 680.400 376.200 681.450 412.950 ;
        RECT 682.950 409.950 688.050 412.050 ;
        RECT 692.100 402.600 693.300 422.400 ;
        RECT 700.950 415.950 703.050 418.050 ;
        RECT 691.950 400.500 694.050 402.600 ;
        RECT 682.950 397.950 685.050 400.050 ;
        RECT 679.950 374.100 682.050 376.200 ;
        RECT 683.400 373.050 684.450 397.950 ;
        RECT 691.950 391.950 694.050 394.050 ;
        RECT 688.950 385.950 691.050 388.050 ;
        RECT 689.400 373.050 690.450 385.950 ;
        RECT 673.950 370.950 676.050 373.050 ;
        RECT 681.000 372.900 685.050 373.050 ;
        RECT 679.950 370.950 685.050 372.900 ;
        RECT 688.950 370.950 691.050 373.050 ;
        RECT 652.950 367.950 655.050 370.050 ;
        RECT 664.950 364.950 667.050 370.050 ;
        RECT 670.950 367.950 673.050 370.050 ;
        RECT 655.950 361.950 658.050 364.050 ;
        RECT 652.950 343.950 655.050 346.050 ;
        RECT 640.950 331.950 643.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 631.950 328.950 634.050 331.050 ;
        RECT 634.950 328.950 640.050 331.050 ;
        RECT 614.400 325.050 615.450 328.950 ;
        RECT 647.400 328.050 648.450 334.950 ;
        RECT 646.950 325.950 649.050 328.050 ;
        RECT 613.950 322.950 616.050 325.050 ;
        RECT 622.950 301.950 625.050 304.050 ;
        RECT 637.950 301.950 640.050 304.050 ;
        RECT 610.950 292.950 613.050 295.050 ;
        RECT 613.950 292.950 619.050 295.050 ;
        RECT 619.950 292.950 622.050 295.050 ;
        RECT 574.950 289.050 577.050 292.050 ;
        RECT 580.950 289.950 583.050 292.050 ;
        RECT 604.950 289.950 607.050 292.050 ;
        RECT 573.000 288.450 577.050 289.050 ;
        RECT 572.400 286.950 577.050 288.450 ;
        RECT 572.400 253.050 573.450 286.950 ;
        RECT 581.400 286.050 582.450 289.950 ;
        RECT 580.950 283.950 583.050 286.050 ;
        RECT 613.950 283.950 616.050 289.050 ;
        RECT 595.950 271.950 598.050 274.050 ;
        RECT 574.950 268.950 577.050 271.050 ;
        RECT 575.400 265.050 576.450 268.950 ;
        RECT 577.950 265.950 580.050 268.050 ;
        RECT 574.950 262.950 577.050 265.050 ;
        RECT 575.400 256.050 576.450 262.950 ;
        RECT 578.400 262.050 579.450 265.950 ;
        RECT 596.400 262.050 597.450 271.950 ;
        RECT 601.950 265.950 604.050 268.050 ;
        RECT 602.400 262.050 603.450 265.950 ;
        RECT 577.950 259.950 580.050 262.050 ;
        RECT 589.950 259.950 592.050 262.050 ;
        RECT 595.950 259.950 598.050 262.050 ;
        RECT 601.950 259.950 604.050 262.050 ;
        RECT 607.950 259.950 610.050 265.050 ;
        RECT 620.400 262.050 621.450 292.950 ;
        RECT 623.400 292.050 624.450 301.950 ;
        RECT 638.400 298.050 639.450 301.950 ;
        RECT 649.950 298.950 652.050 301.050 ;
        RECT 630.000 294.450 634.050 295.050 ;
        RECT 629.400 292.950 634.050 294.450 ;
        RECT 637.950 292.950 640.050 298.050 ;
        RECT 646.950 295.950 649.050 298.050 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 623.400 268.050 624.450 289.950 ;
        RECT 625.950 283.950 628.050 286.050 ;
        RECT 629.400 285.450 630.450 292.950 ;
        RECT 631.950 286.950 637.050 289.050 ;
        RECT 629.400 284.400 633.450 285.450 ;
        RECT 622.950 265.950 625.050 268.050 ;
        RECT 626.400 262.050 627.450 283.950 ;
        RECT 619.950 259.950 622.050 262.050 ;
        RECT 625.950 259.950 628.050 262.050 ;
        RECT 574.950 253.950 577.050 256.050 ;
        RECT 577.950 253.950 583.050 256.050 ;
        RECT 571.950 250.950 574.050 253.050 ;
        RECT 571.950 241.950 574.050 244.050 ;
        RECT 572.400 217.050 573.450 241.950 ;
        RECT 574.950 217.950 577.050 220.050 ;
        RECT 571.950 211.950 574.050 217.050 ;
        RECT 575.400 211.050 576.450 217.950 ;
        RECT 574.950 208.950 577.050 211.050 ;
        RECT 575.400 199.050 576.450 208.950 ;
        RECT 574.950 196.950 577.050 199.050 ;
        RECT 590.400 198.450 591.450 259.950 ;
        RECT 604.950 250.950 607.050 256.050 ;
        RECT 607.950 253.950 613.050 256.050 ;
        RECT 616.950 253.950 619.050 256.050 ;
        RECT 601.950 235.950 604.050 238.050 ;
        RECT 607.950 235.950 610.050 238.050 ;
        RECT 598.950 226.950 601.050 229.050 ;
        RECT 590.400 197.400 594.450 198.450 ;
        RECT 589.950 193.950 592.050 196.050 ;
        RECT 568.950 184.950 571.050 187.050 ;
        RECT 590.400 184.050 591.450 193.950 ;
        RECT 571.950 181.950 574.050 184.050 ;
        RECT 589.950 181.950 592.050 184.050 ;
        RECT 562.950 166.500 565.050 168.600 ;
        RECT 562.950 160.950 565.050 163.050 ;
        RECT 544.950 151.950 547.050 154.050 ;
        RECT 550.950 151.950 553.050 154.050 ;
        RECT 556.950 151.950 559.050 154.050 ;
        RECT 526.950 142.950 529.050 145.050 ;
        RECT 545.400 142.050 546.450 151.950 ;
        RECT 550.950 147.300 553.050 149.400 ;
        RECT 551.850 143.700 553.050 147.300 ;
        RECT 544.950 139.950 547.050 142.050 ;
        RECT 550.950 141.600 553.050 143.700 ;
        RECT 526.950 136.950 529.050 139.050 ;
        RECT 532.950 136.950 535.050 139.050 ;
        RECT 520.950 124.500 523.050 126.600 ;
        RECT 490.950 109.950 493.050 112.050 ;
        RECT 514.950 109.950 517.050 112.050 ;
        RECT 520.950 110.400 523.050 112.500 ;
        RECT 487.950 103.950 490.050 106.050 ;
        RECT 491.400 100.050 492.450 109.950 ;
        RECT 511.950 106.950 514.050 109.050 ;
        RECT 493.950 105.450 498.000 106.050 ;
        RECT 493.950 103.950 498.450 105.450 ;
        RECT 497.400 100.050 498.450 103.950 ;
        RECT 505.950 100.950 508.050 103.050 ;
        RECT 484.950 97.950 487.050 100.050 ;
        RECT 490.950 97.950 493.050 100.050 ;
        RECT 496.950 97.950 499.050 100.050 ;
        RECT 502.950 97.950 505.050 100.050 ;
        RECT 481.950 94.950 484.050 97.050 ;
        RECT 485.400 91.050 486.450 97.950 ;
        RECT 493.950 94.950 496.050 97.050 ;
        RECT 484.950 88.950 487.050 91.050 ;
        RECT 478.950 82.950 481.050 85.050 ;
        RECT 479.400 61.050 480.450 82.950 ;
        RECT 463.950 58.950 468.450 61.050 ;
        RECT 478.950 58.950 481.050 61.050 ;
        RECT 484.950 58.950 490.050 61.050 ;
        RECT 467.400 55.050 468.450 58.950 ;
        RECT 445.950 51.900 450.000 52.050 ;
        RECT 445.950 49.950 451.050 51.900 ;
        RECT 460.950 49.950 463.050 55.050 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 472.950 52.950 478.050 55.050 ;
        RECT 481.950 52.950 484.050 55.050 ;
        RECT 487.950 52.950 490.050 55.050 ;
        RECT 448.950 49.800 451.050 49.950 ;
        RECT 421.950 43.950 424.050 46.050 ;
        RECT 439.950 43.950 442.050 46.050 ;
        RECT 415.950 28.950 418.050 31.050 ;
        RECT 422.400 28.050 423.450 43.950 ;
        RECT 409.950 22.950 412.050 28.050 ;
        RECT 421.950 25.950 424.050 28.050 ;
        RECT 436.950 22.950 439.050 28.050 ;
        RECT 442.950 25.950 448.050 28.050 ;
        RECT 451.950 25.950 454.050 31.050 ;
        RECT 467.400 28.050 468.450 52.950 ;
        RECT 482.400 40.050 483.450 52.950 ;
        RECT 481.950 37.950 484.050 40.050 ;
        RECT 488.400 36.450 489.450 52.950 ;
        RECT 494.400 52.050 495.450 94.950 ;
        RECT 497.400 64.050 498.450 97.950 ;
        RECT 503.400 94.050 504.450 97.950 ;
        RECT 502.950 91.950 505.050 94.050 ;
        RECT 506.400 91.050 507.450 100.950 ;
        RECT 512.400 97.050 513.450 106.950 ;
        RECT 517.950 100.950 520.050 106.050 ;
        RECT 511.950 94.950 514.050 97.050 ;
        RECT 521.850 95.400 523.050 110.400 ;
        RECT 527.400 106.050 528.450 136.950 ;
        RECT 529.950 127.950 532.050 133.050 ;
        RECT 529.950 118.950 532.050 121.050 ;
        RECT 526.950 103.950 529.050 106.050 ;
        RECT 530.400 103.050 531.450 118.950 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 520.950 93.300 523.050 95.400 ;
        RECT 499.950 88.950 502.050 91.050 ;
        RECT 505.800 88.950 507.900 91.050 ;
        RECT 509.100 88.950 511.200 91.050 ;
        RECT 521.850 89.700 523.050 93.300 ;
        RECT 500.400 70.050 501.450 88.950 ;
        RECT 499.950 67.950 502.050 70.050 ;
        RECT 496.950 61.950 499.050 64.050 ;
        RECT 500.400 61.050 501.450 67.950 ;
        RECT 509.400 61.050 510.450 88.950 ;
        RECT 520.950 87.600 523.050 89.700 ;
        RECT 530.400 76.050 531.450 100.950 ;
        RECT 533.400 100.050 534.450 136.950 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 539.400 127.050 540.450 133.950 ;
        RECT 546.000 132.450 550.050 133.050 ;
        RECT 545.400 130.950 550.050 132.450 ;
        RECT 538.950 124.950 541.050 127.050 ;
        RECT 545.400 121.050 546.450 130.950 ;
        RECT 551.850 126.600 553.050 141.600 ;
        RECT 557.400 136.050 558.450 151.950 ;
        RECT 556.950 133.950 562.050 136.050 ;
        RECT 550.950 124.500 553.050 126.600 ;
        RECT 544.950 118.950 547.050 121.050 ;
        RECT 550.950 118.950 553.050 121.050 ;
        RECT 541.950 110.400 544.050 112.500 ;
        RECT 532.950 97.950 535.050 100.050 ;
        RECT 535.950 97.950 538.050 100.050 ;
        RECT 536.400 79.050 537.450 97.950 ;
        RECT 542.100 90.600 543.300 110.400 ;
        RECT 551.400 97.050 552.450 118.950 ;
        RECT 556.950 109.950 559.050 112.050 ;
        RECT 550.950 94.950 553.050 97.050 ;
        RECT 551.400 91.050 552.450 94.950 ;
        RECT 557.400 94.050 558.450 109.950 ;
        RECT 559.950 106.950 562.050 109.050 ;
        RECT 560.400 103.050 561.450 106.950 ;
        RECT 563.400 103.050 564.450 160.950 ;
        RECT 572.400 153.450 573.450 181.950 ;
        RECT 579.000 177.450 583.050 178.050 ;
        RECT 578.400 175.950 583.050 177.450 ;
        RECT 586.950 175.950 592.050 178.050 ;
        RECT 578.400 163.050 579.450 175.950 ;
        RECT 580.950 166.950 583.050 169.050 ;
        RECT 577.950 160.950 580.050 163.050 ;
        RECT 566.400 152.400 573.450 153.450 ;
        RECT 566.400 139.050 567.450 152.400 ;
        RECT 571.950 146.400 574.050 148.500 ;
        RECT 565.950 136.950 568.050 139.050 ;
        RECT 572.100 126.600 573.300 146.400 ;
        RECT 577.950 139.950 580.050 142.050 ;
        RECT 571.950 124.500 574.050 126.600 ;
        RECT 565.950 103.950 568.050 109.050 ;
        RECT 571.950 103.950 574.050 106.050 ;
        RECT 559.950 100.950 562.050 103.050 ;
        RECT 562.950 100.950 565.050 103.050 ;
        RECT 568.950 100.950 571.050 103.050 ;
        RECT 562.950 94.950 568.050 97.050 ;
        RECT 556.950 91.950 559.050 94.050 ;
        RECT 541.950 88.500 544.050 90.600 ;
        RECT 550.950 88.950 553.050 91.050 ;
        RECT 535.950 76.950 538.050 79.050 ;
        RECT 523.950 73.950 526.050 76.050 ;
        RECT 529.950 73.950 532.050 76.050 ;
        RECT 544.950 73.950 547.050 76.050 ;
        RECT 499.950 58.950 502.050 61.050 ;
        RECT 505.950 59.400 510.450 61.050 ;
        RECT 505.950 58.950 510.000 59.400 ;
        RECT 520.950 58.950 523.050 64.050 ;
        RECT 508.950 53.100 511.050 58.050 ;
        RECT 521.400 55.050 522.450 58.950 ;
        RECT 524.400 55.050 525.450 73.950 ;
        RECT 532.950 68.400 535.050 70.500 ;
        RECT 520.950 52.950 523.050 55.050 ;
        RECT 523.950 52.950 526.050 55.050 ;
        RECT 493.950 49.950 496.050 52.050 ;
        RECT 508.950 49.800 511.050 51.900 ;
        RECT 493.950 37.950 496.050 40.050 ;
        RECT 485.400 35.400 489.450 36.450 ;
        RECT 466.950 25.950 469.050 28.050 ;
        RECT 472.950 22.950 475.050 28.050 ;
        RECT 478.950 25.950 484.050 28.050 ;
        RECT 485.400 22.050 486.450 35.400 ;
        RECT 487.950 31.950 490.050 34.050 ;
        RECT 488.400 28.050 489.450 31.950 ;
        RECT 487.950 25.950 490.050 28.050 ;
        RECT 494.400 25.050 495.450 37.950 ;
        RECT 509.400 25.050 510.450 49.800 ;
        RECT 524.400 45.450 525.450 52.950 ;
        RECT 533.700 48.600 534.900 68.400 ;
        RECT 538.950 58.950 541.050 64.050 ;
        RECT 545.400 58.050 546.450 73.950 ;
        RECT 553.950 69.300 556.050 71.400 ;
        RECT 553.950 65.700 555.150 69.300 ;
        RECT 553.950 63.600 556.050 65.700 ;
        RECT 569.400 64.050 570.450 100.950 ;
        RECT 544.950 55.950 547.050 58.050 ;
        RECT 553.950 48.600 555.150 63.600 ;
        RECT 568.950 61.950 571.050 64.050 ;
        RECT 572.400 61.050 573.450 103.950 ;
        RECT 578.400 100.050 579.450 139.950 ;
        RECT 581.400 121.050 582.450 166.950 ;
        RECT 589.950 136.950 592.050 142.050 ;
        RECT 593.400 141.450 594.450 197.400 ;
        RECT 595.950 196.950 598.050 199.050 ;
        RECT 596.400 187.050 597.450 196.950 ;
        RECT 595.950 184.950 598.050 187.050 ;
        RECT 596.400 165.450 597.450 184.950 ;
        RECT 599.400 169.050 600.450 226.950 ;
        RECT 602.400 202.050 603.450 235.950 ;
        RECT 604.950 232.950 607.050 235.050 ;
        RECT 601.950 199.950 604.050 202.050 ;
        RECT 605.400 190.050 606.450 232.950 ;
        RECT 604.950 187.950 607.050 190.050 ;
        RECT 601.950 181.950 604.050 184.050 ;
        RECT 604.950 181.950 607.050 184.050 ;
        RECT 602.400 178.050 603.450 181.950 ;
        RECT 605.400 178.050 606.450 181.950 ;
        RECT 601.950 175.950 604.050 178.050 ;
        RECT 604.950 175.950 607.050 178.050 ;
        RECT 598.950 166.950 601.050 169.050 ;
        RECT 596.400 164.400 600.450 165.450 ;
        RECT 593.400 141.000 597.450 141.450 ;
        RECT 593.400 140.400 598.050 141.000 ;
        RECT 595.950 136.950 598.050 140.400 ;
        RECT 583.950 130.950 586.050 133.050 ;
        RECT 592.950 130.950 598.050 133.050 ;
        RECT 580.950 118.950 583.050 121.050 ;
        RECT 584.400 112.050 585.450 130.950 ;
        RECT 595.950 118.950 598.050 121.050 ;
        RECT 583.950 109.950 586.050 112.050 ;
        RECT 580.950 103.950 586.050 106.050 ;
        RECT 586.950 103.950 589.050 109.050 ;
        RECT 596.400 106.050 597.450 118.950 ;
        RECT 595.950 103.950 598.050 106.050 ;
        RECT 577.950 94.950 580.050 100.050 ;
        RECT 583.950 97.950 586.050 100.050 ;
        RECT 584.400 94.050 585.450 97.950 ;
        RECT 583.950 91.950 586.050 94.050 ;
        RECT 596.400 82.050 597.450 103.950 ;
        RECT 599.400 103.050 600.450 164.400 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 602.400 109.050 603.450 133.950 ;
        RECT 608.400 112.050 609.450 235.950 ;
        RECT 617.400 226.050 618.450 253.950 ;
        RECT 619.950 250.950 622.050 253.050 ;
        RECT 610.950 223.950 613.050 226.050 ;
        RECT 616.950 223.950 619.050 226.050 ;
        RECT 611.400 181.050 612.450 223.950 ;
        RECT 613.950 211.950 619.050 214.050 ;
        RECT 616.950 205.950 619.050 208.050 ;
        RECT 617.400 184.050 618.450 205.950 ;
        RECT 616.950 181.950 619.050 184.050 ;
        RECT 610.950 175.950 613.050 181.050 ;
        RECT 620.400 180.450 621.450 250.950 ;
        RECT 632.400 244.050 633.450 284.400 ;
        RECT 635.400 280.050 636.450 286.950 ;
        RECT 634.950 277.950 637.050 280.050 ;
        RECT 635.400 247.050 636.450 277.950 ;
        RECT 640.950 268.950 643.050 271.050 ;
        RECT 641.400 262.050 642.450 268.950 ;
        RECT 637.950 259.950 640.050 262.050 ;
        RECT 640.950 259.950 643.050 262.050 ;
        RECT 638.400 256.050 639.450 259.950 ;
        RECT 637.950 253.950 640.050 256.050 ;
        RECT 634.950 244.950 637.050 247.050 ;
        RECT 631.950 241.950 634.050 244.050 ;
        RECT 632.400 229.050 633.450 241.950 ;
        RECT 631.950 226.950 634.050 229.050 ;
        RECT 625.950 224.400 628.050 226.500 ;
        RECT 622.950 220.950 625.050 223.050 ;
        RECT 623.400 208.050 624.450 220.950 ;
        RECT 622.950 205.950 625.050 208.050 ;
        RECT 626.700 204.600 627.900 224.400 ;
        RECT 638.400 223.050 639.450 253.950 ;
        RECT 643.950 250.950 646.050 256.050 ;
        RECT 644.400 235.050 645.450 250.950 ;
        RECT 647.400 238.050 648.450 295.950 ;
        RECT 650.400 294.450 651.450 298.950 ;
        RECT 653.400 298.050 654.450 343.950 ;
        RECT 656.400 307.050 657.450 361.950 ;
        RECT 674.400 340.050 675.450 370.950 ;
        RECT 679.950 370.800 682.050 370.950 ;
        RECT 692.400 367.050 693.450 391.950 ;
        RECT 701.400 388.050 702.450 415.950 ;
        RECT 704.400 415.050 705.450 481.950 ;
        RECT 710.400 454.050 711.450 505.950 ;
        RECT 713.400 496.050 714.450 508.950 ;
        RECT 712.950 493.950 715.050 496.050 ;
        RECT 716.400 492.450 717.450 520.950 ;
        RECT 719.400 520.050 720.450 526.950 ;
        RECT 725.400 526.050 726.450 538.950 ;
        RECT 737.400 529.050 738.450 544.950 ;
        RECT 740.400 535.050 741.450 575.400 ;
        RECT 743.400 541.050 744.450 604.950 ;
        RECT 748.950 598.950 751.050 601.050 ;
        RECT 754.950 598.950 757.050 604.050 ;
        RECT 749.400 592.050 750.450 598.950 ;
        RECT 748.950 589.950 751.050 592.050 ;
        RECT 751.950 580.950 754.050 583.050 ;
        RECT 752.400 574.050 753.450 580.950 ;
        RECT 751.950 571.950 754.050 574.050 ;
        RECT 748.950 565.950 751.050 568.050 ;
        RECT 745.950 550.950 748.050 553.050 ;
        RECT 742.950 538.950 745.050 541.050 ;
        RECT 739.950 532.950 742.050 535.050 ;
        RECT 746.400 529.050 747.450 550.950 ;
        RECT 749.400 547.050 750.450 565.950 ;
        RECT 748.950 544.950 751.050 547.050 ;
        RECT 752.400 544.050 753.450 571.950 ;
        RECT 751.950 541.950 754.050 544.050 ;
        RECT 758.400 538.050 759.450 610.950 ;
        RECT 761.400 607.050 762.450 619.950 ;
        RECT 760.950 604.950 763.050 607.050 ;
        RECT 764.400 574.050 765.450 637.950 ;
        RECT 766.950 616.950 769.050 619.050 ;
        RECT 767.400 601.050 768.450 616.950 ;
        RECT 766.950 598.950 769.050 601.050 ;
        RECT 772.950 598.950 775.050 604.050 ;
        RECT 775.950 577.950 778.050 580.050 ;
        RECT 766.950 574.950 769.050 577.050 ;
        RECT 760.950 572.400 765.450 574.050 ;
        RECT 760.950 571.950 765.000 572.400 ;
        RECT 767.400 553.050 768.450 574.950 ;
        RECT 776.400 568.050 777.450 577.950 ;
        RECT 782.400 576.450 783.450 646.950 ;
        RECT 788.400 625.050 789.450 646.950 ;
        RECT 794.400 646.050 795.450 679.950 ;
        RECT 805.950 658.950 808.050 661.050 ;
        RECT 796.950 646.950 799.050 652.050 ;
        RECT 790.950 644.400 795.450 646.050 ;
        RECT 790.950 643.950 795.000 644.400 ;
        RECT 806.400 643.050 807.450 658.950 ;
        RECT 815.400 646.050 816.450 682.950 ;
        RECT 818.400 679.050 819.450 719.400 ;
        RECT 820.950 715.950 826.050 718.050 ;
        RECT 827.400 697.050 828.450 724.950 ;
        RECT 820.950 694.950 823.050 697.050 ;
        RECT 826.950 694.950 829.050 697.050 ;
        RECT 821.400 685.050 822.450 694.950 ;
        RECT 829.950 691.950 832.050 694.050 ;
        RECT 820.950 682.950 823.050 685.050 ;
        RECT 817.950 676.950 820.050 679.050 ;
        RECT 823.950 676.950 826.050 682.050 ;
        RECT 820.950 646.950 826.050 649.050 ;
        RECT 826.950 646.950 829.050 649.050 ;
        RECT 814.950 643.950 817.050 646.050 ;
        RECT 799.950 640.950 802.050 643.050 ;
        RECT 800.400 637.050 801.450 640.950 ;
        RECT 805.950 637.950 808.050 643.050 ;
        RECT 817.950 640.950 820.050 646.050 ;
        RECT 823.950 640.950 826.050 643.050 ;
        RECT 811.950 637.950 817.050 640.050 ;
        RECT 799.950 634.950 802.050 637.050 ;
        RECT 796.950 625.950 799.050 628.050 ;
        RECT 787.950 622.950 790.050 625.050 ;
        RECT 790.950 616.950 793.050 619.050 ;
        RECT 787.950 610.950 790.050 613.050 ;
        RECT 784.950 601.950 787.050 607.050 ;
        RECT 788.400 598.050 789.450 610.950 ;
        RECT 791.400 607.200 792.450 616.950 ;
        RECT 797.400 610.050 798.450 625.950 ;
        RECT 811.950 622.950 814.050 625.050 ;
        RECT 790.950 605.100 793.050 607.200 ;
        RECT 796.950 604.950 799.050 610.050 ;
        RECT 802.950 607.950 805.050 610.050 ;
        RECT 792.000 603.900 796.050 604.050 ;
        RECT 790.950 601.950 796.050 603.900 ;
        RECT 790.950 601.800 793.050 601.950 ;
        RECT 787.950 595.950 790.050 598.050 ;
        RECT 787.950 589.950 790.050 592.050 ;
        RECT 782.400 575.400 786.450 576.450 ;
        RECT 781.950 568.950 784.050 574.050 ;
        RECT 769.950 565.950 772.050 568.050 ;
        RECT 775.950 565.950 778.050 568.050 ;
        RECT 766.950 550.950 769.050 553.050 ;
        RECT 763.950 541.950 766.050 544.050 ;
        RECT 751.950 535.950 754.050 538.050 ;
        RECT 757.950 535.950 760.050 538.050 ;
        RECT 748.950 532.950 751.050 535.050 ;
        RECT 730.950 526.950 733.050 529.050 ;
        RECT 737.400 527.400 742.050 529.050 ;
        RECT 738.000 526.950 742.050 527.400 ;
        RECT 745.950 526.950 748.050 529.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 731.400 523.050 732.450 526.950 ;
        RECT 727.800 520.950 729.900 523.050 ;
        RECT 731.100 520.950 733.200 523.050 ;
        RECT 736.950 520.950 742.050 523.050 ;
        RECT 718.950 517.950 721.050 520.050 ;
        RECT 718.950 511.950 721.050 514.050 ;
        RECT 719.400 496.050 720.450 511.950 ;
        RECT 728.400 496.050 729.450 520.950 ;
        RECT 742.950 517.950 745.050 523.050 ;
        RECT 749.400 499.050 750.450 532.950 ;
        RECT 752.400 523.050 753.450 535.950 ;
        RECT 764.400 529.050 765.450 541.950 ;
        RECT 757.950 523.950 760.050 529.050 ;
        RECT 763.950 526.950 766.050 529.050 ;
        RECT 751.950 520.950 754.050 523.050 ;
        RECT 754.950 522.450 757.050 523.050 ;
        RECT 754.950 521.400 762.450 522.450 ;
        RECT 754.950 520.950 757.050 521.400 ;
        RECT 757.950 517.950 760.050 520.050 ;
        RECT 758.400 514.050 759.450 517.950 ;
        RECT 761.400 517.050 762.450 521.400 ;
        RECT 760.950 514.950 763.050 517.050 ;
        RECT 757.950 511.950 760.050 514.050 ;
        RECT 764.400 511.050 765.450 526.950 ;
        RECT 770.400 526.050 771.450 565.950 ;
        RECT 785.400 559.050 786.450 575.400 ;
        RECT 784.950 556.950 787.050 559.050 ;
        RECT 775.950 529.950 778.050 535.050 ;
        RECT 781.950 529.950 787.050 532.050 ;
        RECT 769.950 523.950 772.050 526.050 ;
        RECT 772.950 523.950 775.050 526.050 ;
        RECT 766.950 520.950 769.050 523.050 ;
        RECT 763.950 508.950 766.050 511.050 ;
        RECT 767.400 502.050 768.450 520.950 ;
        RECT 769.950 517.950 772.050 520.050 ;
        RECT 770.400 514.050 771.450 517.950 ;
        RECT 769.950 511.950 772.050 514.050 ;
        RECT 754.950 499.950 757.050 502.050 ;
        RECT 766.950 499.950 769.050 502.050 ;
        RECT 733.950 496.950 736.050 499.050 ;
        RECT 748.950 496.950 751.050 499.050 ;
        RECT 718.950 493.950 721.050 496.050 ;
        RECT 727.950 493.950 730.050 496.050 ;
        RECT 713.400 491.400 717.450 492.450 ;
        RECT 713.400 469.050 714.450 491.400 ;
        RECT 715.950 487.950 718.050 490.050 ;
        RECT 716.400 484.050 717.450 487.950 ;
        RECT 719.400 487.050 720.450 493.950 ;
        RECT 721.950 487.950 727.050 490.050 ;
        RECT 727.950 487.950 733.050 490.050 ;
        RECT 718.950 484.950 721.050 487.050 ;
        RECT 715.950 481.950 718.050 484.050 ;
        RECT 712.950 466.950 715.050 469.050 ;
        RECT 718.950 460.950 721.050 463.050 ;
        RECT 715.950 457.950 718.050 460.050 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 709.950 445.950 712.050 448.050 ;
        RECT 710.400 418.050 711.450 445.950 ;
        RECT 716.400 445.050 717.450 457.950 ;
        RECT 719.400 454.050 720.450 460.950 ;
        RECT 730.950 454.950 733.050 457.050 ;
        RECT 718.950 451.950 721.050 454.050 ;
        RECT 715.950 442.950 718.050 445.050 ;
        RECT 719.400 418.050 720.450 451.950 ;
        RECT 731.400 451.050 732.450 454.950 ;
        RECT 724.950 445.950 727.050 451.050 ;
        RECT 730.950 448.950 733.050 451.050 ;
        RECT 730.950 439.950 733.050 442.050 ;
        RECT 724.950 427.950 727.050 430.050 ;
        RECT 709.950 415.950 712.050 418.050 ;
        RECT 718.950 415.950 721.050 418.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 709.950 409.950 712.050 412.050 ;
        RECT 715.950 409.950 721.050 412.050 ;
        RECT 706.950 406.950 709.050 409.050 ;
        RECT 700.950 385.950 703.050 388.050 ;
        RECT 694.950 373.950 697.050 376.050 ;
        RECT 679.950 364.950 682.050 367.050 ;
        RECT 685.950 364.950 688.050 367.050 ;
        RECT 691.950 364.950 694.050 367.050 ;
        RECT 676.950 358.950 679.050 361.050 ;
        RECT 658.950 337.950 664.050 340.050 ;
        RECT 667.950 334.950 670.050 340.050 ;
        RECT 670.950 337.950 676.050 340.050 ;
        RECT 661.950 331.950 667.050 334.050 ;
        RECT 670.950 331.950 673.050 334.050 ;
        RECT 671.400 313.050 672.450 331.950 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 655.950 304.950 658.050 307.050 ;
        RECT 677.400 301.050 678.450 358.950 ;
        RECT 680.400 352.050 681.450 364.950 ;
        RECT 686.400 358.050 687.450 364.950 ;
        RECT 685.950 355.950 688.050 358.050 ;
        RECT 679.950 349.950 682.050 352.050 ;
        RECT 682.950 344.400 685.050 346.500 ;
        RECT 683.700 324.600 684.900 344.400 ;
        RECT 695.400 337.050 696.450 373.950 ;
        RECT 707.400 373.050 708.450 406.950 ;
        RECT 710.400 400.050 711.450 409.950 ;
        RECT 721.950 406.950 724.050 412.050 ;
        RECT 709.950 397.950 712.050 400.050 ;
        RECT 706.950 370.950 709.050 373.050 ;
        RECT 712.950 370.950 715.050 376.050 ;
        RECT 721.950 373.050 724.050 376.050 ;
        RECT 725.400 373.050 726.450 427.950 ;
        RECT 731.400 412.050 732.450 439.950 ;
        RECT 734.400 429.450 735.450 496.950 ;
        RECT 736.950 493.950 739.050 496.050 ;
        RECT 737.400 453.450 738.450 493.950 ;
        RECT 739.950 490.950 742.050 496.050 ;
        RECT 751.950 493.950 754.050 496.050 ;
        RECT 745.950 490.950 748.050 493.050 ;
        RECT 746.400 481.050 747.450 490.950 ;
        RECT 748.950 489.450 751.050 493.050 ;
        RECT 752.400 489.450 753.450 493.950 ;
        RECT 755.400 490.050 756.450 499.950 ;
        RECT 773.400 496.050 774.450 523.950 ;
        RECT 766.950 493.950 772.050 496.050 ;
        RECT 772.950 493.950 775.050 496.050 ;
        RECT 776.400 490.050 777.450 529.950 ;
        RECT 778.950 523.950 781.050 526.050 ;
        RECT 748.950 488.400 753.450 489.450 ;
        RECT 748.950 484.950 751.050 488.400 ;
        RECT 754.950 484.950 757.050 490.050 ;
        RECT 766.950 487.950 772.050 490.050 ;
        RECT 775.950 487.950 778.050 490.050 ;
        RECT 776.400 484.050 777.450 487.950 ;
        RECT 775.950 481.950 778.050 484.050 ;
        RECT 745.950 478.950 748.050 481.050 ;
        RECT 779.400 469.050 780.450 523.950 ;
        RECT 788.400 508.050 789.450 589.950 ;
        RECT 799.950 586.950 802.050 589.050 ;
        RECT 790.950 574.950 793.050 577.050 ;
        RECT 791.400 571.200 792.450 574.950 ;
        RECT 790.950 569.100 793.050 571.200 ;
        RECT 796.950 568.950 799.050 574.050 ;
        RECT 792.000 567.900 795.000 568.050 ;
        RECT 790.950 565.950 796.050 567.900 ;
        RECT 790.950 565.800 793.050 565.950 ;
        RECT 793.950 565.800 796.050 565.950 ;
        RECT 800.400 532.050 801.450 586.950 ;
        RECT 803.400 574.050 804.450 607.950 ;
        RECT 812.400 604.050 813.450 622.950 ;
        RECT 817.950 610.950 820.050 613.050 ;
        RECT 814.950 604.950 817.050 610.050 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 818.400 595.050 819.450 610.950 ;
        RECT 817.950 592.950 820.050 595.050 ;
        RECT 824.400 589.050 825.450 640.950 ;
        RECT 823.950 586.950 826.050 589.050 ;
        RECT 808.950 577.950 811.050 580.050 ;
        RECT 802.950 571.950 805.050 574.050 ;
        RECT 803.400 535.050 804.450 571.950 ;
        RECT 809.400 568.050 810.450 577.950 ;
        RECT 817.950 574.950 820.050 577.050 ;
        RECT 808.950 565.950 811.050 568.050 ;
        RECT 814.950 565.950 817.050 571.050 ;
        RECT 802.950 532.950 808.050 535.050 ;
        RECT 790.950 529.950 793.050 532.050 ;
        RECT 799.950 529.950 802.050 532.050 ;
        RECT 791.400 517.050 792.450 529.950 ;
        RECT 800.400 529.050 801.450 529.950 ;
        RECT 800.400 527.400 805.050 529.050 ;
        RECT 801.000 526.950 805.050 527.400 ;
        RECT 818.400 526.050 819.450 574.950 ;
        RECT 823.950 571.950 826.050 574.050 ;
        RECT 824.400 535.050 825.450 571.950 ;
        RECT 823.950 532.950 826.050 535.050 ;
        RECT 796.950 523.950 802.050 526.050 ;
        RECT 817.950 523.950 820.050 526.050 ;
        RECT 790.950 514.950 793.050 517.050 ;
        RECT 787.950 505.950 790.050 508.050 ;
        RECT 784.950 496.950 787.050 499.050 ;
        RECT 781.950 493.950 784.050 496.050 ;
        RECT 782.400 487.200 783.450 493.950 ;
        RECT 781.950 485.100 784.050 487.200 ;
        RECT 781.950 481.800 784.050 483.900 ;
        RECT 748.950 466.950 751.050 469.050 ;
        RECT 766.950 466.950 769.050 469.050 ;
        RECT 778.950 466.950 781.050 469.050 ;
        RECT 737.400 452.400 741.450 453.450 ;
        RECT 736.950 445.950 739.050 451.050 ;
        RECT 734.400 428.400 738.450 429.450 ;
        RECT 733.950 424.950 736.050 427.050 ;
        RECT 734.400 418.050 735.450 424.950 ;
        RECT 733.950 415.950 736.050 418.050 ;
        RECT 730.950 409.950 733.050 412.050 ;
        RECT 730.950 388.950 733.050 391.050 ;
        RECT 727.950 385.950 730.050 388.050 ;
        RECT 721.950 371.400 726.450 373.050 ;
        RECT 721.950 370.950 726.000 371.400 ;
        RECT 703.950 364.950 706.050 367.050 ;
        RECT 704.400 352.050 705.450 364.950 ;
        RECT 707.400 364.050 708.450 370.950 ;
        RECT 712.950 367.050 715.050 367.200 ;
        RECT 709.950 365.100 715.050 367.050 ;
        RECT 709.950 364.950 714.000 365.100 ;
        RECT 724.950 364.950 727.050 370.050 ;
        RECT 706.950 361.950 709.050 364.050 ;
        RECT 712.950 361.800 715.050 363.900 ;
        RECT 709.950 352.950 712.050 355.050 ;
        RECT 703.950 349.950 706.050 352.050 ;
        RECT 703.950 344.400 706.050 346.500 ;
        RECT 688.950 331.950 691.050 337.050 ;
        RECT 694.950 334.950 697.050 337.050 ;
        RECT 703.950 329.400 705.150 344.400 ;
        RECT 706.950 334.950 709.050 340.050 ;
        RECT 703.950 327.300 706.050 329.400 ;
        RECT 682.950 322.500 685.050 324.600 ;
        RECT 703.950 323.700 705.150 327.300 ;
        RECT 697.950 319.950 700.050 322.050 ;
        RECT 703.950 321.600 706.050 323.700 ;
        RECT 676.950 298.950 679.050 301.050 ;
        RECT 688.950 298.950 691.050 301.050 ;
        RECT 652.950 295.950 655.050 298.050 ;
        RECT 655.950 294.450 658.050 295.050 ;
        RECT 650.400 293.400 658.050 294.450 ;
        RECT 650.400 241.050 651.450 293.400 ;
        RECT 655.950 292.950 658.050 293.400 ;
        RECT 661.950 292.950 664.050 295.050 ;
        RECT 676.950 292.950 679.050 295.050 ;
        RECT 652.950 289.050 655.050 292.050 ;
        RECT 662.400 289.050 663.450 292.950 ;
        RECT 652.800 288.000 655.050 289.050 ;
        RECT 652.800 286.950 654.900 288.000 ;
        RECT 655.950 286.950 658.050 289.050 ;
        RECT 661.950 286.950 664.050 289.050 ;
        RECT 652.950 253.950 655.050 259.050 ;
        RECT 649.950 238.950 652.050 241.050 ;
        RECT 646.950 235.950 649.050 238.050 ;
        RECT 643.950 232.950 646.050 235.050 ;
        RECT 646.950 225.300 649.050 227.400 ;
        RECT 637.950 220.950 640.050 223.050 ;
        RECT 646.950 221.700 648.150 225.300 ;
        RECT 646.950 219.600 649.050 221.700 ;
        RECT 631.950 214.950 634.050 217.050 ;
        RECT 632.400 211.050 633.450 214.950 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 631.950 208.950 634.050 211.050 ;
        RECT 625.950 202.500 628.050 204.600 ;
        RECT 634.950 199.950 637.050 202.050 ;
        RECT 622.950 193.950 625.050 196.050 ;
        RECT 623.400 184.050 624.450 193.950 ;
        RECT 631.950 190.950 634.050 193.050 ;
        RECT 622.950 181.950 625.050 184.050 ;
        RECT 620.400 179.400 624.450 180.450 ;
        RECT 616.950 175.950 622.050 178.050 ;
        RECT 610.950 145.950 613.050 148.050 ;
        RECT 611.400 133.050 612.450 145.950 ;
        RECT 619.950 142.950 622.050 145.050 ;
        RECT 613.950 136.950 619.050 139.050 ;
        RECT 610.950 130.950 616.050 133.050 ;
        RECT 620.400 121.050 621.450 142.950 ;
        RECT 623.400 139.050 624.450 179.400 ;
        RECT 625.950 175.950 631.050 178.050 ;
        RECT 622.950 136.950 625.050 139.050 ;
        RECT 619.950 118.950 622.050 121.050 ;
        RECT 607.950 109.950 610.050 112.050 ;
        RECT 601.950 106.950 604.050 109.050 ;
        RECT 613.950 105.450 618.000 106.050 ;
        RECT 613.950 103.950 618.450 105.450 ;
        RECT 598.950 94.950 601.050 103.050 ;
        RECT 604.950 97.950 610.050 100.050 ;
        RECT 610.950 98.100 613.050 103.050 ;
        RECT 610.950 94.800 613.050 96.900 ;
        RECT 577.950 79.950 580.050 82.050 ;
        RECT 595.950 79.950 598.050 82.050 ;
        RECT 571.950 58.950 574.050 61.050 ;
        RECT 556.950 49.950 559.050 55.050 ;
        RECT 565.950 52.950 571.050 55.050 ;
        RECT 532.950 46.500 535.050 48.600 ;
        RECT 553.950 46.500 556.050 48.600 ;
        RECT 524.400 44.400 528.450 45.450 ;
        RECT 527.400 25.050 528.450 44.400 ;
        RECT 529.950 40.950 532.050 43.050 ;
        RECT 493.950 22.950 496.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 526.950 22.950 529.050 25.050 ;
        RECT 530.400 22.050 531.450 40.950 ;
        RECT 538.950 29.100 541.050 34.050 ;
        RECT 559.950 31.950 562.050 34.050 ;
        RECT 550.950 25.950 553.050 28.050 ;
        RECT 442.950 19.950 445.050 22.050 ;
        RECT 406.950 15.300 409.050 17.400 ;
        RECT 443.400 16.050 444.450 19.950 ;
        RECT 448.950 16.950 451.050 22.050 ;
        RECT 478.950 19.950 481.050 22.050 ;
        RECT 484.950 19.950 487.050 22.050 ;
        RECT 529.950 19.950 532.050 22.050 ;
        RECT 538.950 19.950 541.050 25.050 ;
        RECT 544.950 22.950 550.050 25.050 ;
        RECT 385.950 10.500 388.050 12.600 ;
        RECT 406.950 11.700 408.150 15.300 ;
        RECT 442.950 13.950 445.050 16.050 ;
        RECT 406.950 9.600 409.050 11.700 ;
        RECT 479.400 7.050 480.450 19.950 ;
        RECT 551.400 19.050 552.450 25.950 ;
        RECT 560.400 22.050 561.450 31.950 ;
        RECT 572.400 28.050 573.450 58.950 ;
        RECT 578.400 43.050 579.450 79.950 ;
        RECT 611.400 73.050 612.450 94.800 ;
        RECT 583.950 68.400 586.050 70.500 ;
        RECT 604.950 69.300 607.050 71.400 ;
        RECT 610.950 70.950 613.050 73.050 ;
        RECT 584.700 48.600 585.900 68.400 ;
        RECT 604.950 65.700 606.150 69.300 ;
        RECT 589.950 58.950 592.050 64.050 ;
        RECT 604.950 63.600 607.050 65.700 ;
        RECT 592.950 55.950 598.050 58.050 ;
        RECT 604.950 48.600 606.150 63.600 ;
        RECT 611.400 55.050 612.450 70.950 ;
        RECT 617.400 64.050 618.450 103.950 ;
        RECT 619.950 94.950 625.050 97.050 ;
        RECT 629.400 64.200 630.450 175.950 ;
        RECT 632.400 160.050 633.450 190.950 ;
        RECT 635.400 181.050 636.450 199.950 ;
        RECT 634.950 178.950 637.050 181.050 ;
        RECT 631.950 157.950 634.050 160.050 ;
        RECT 638.400 154.050 639.450 211.950 ;
        RECT 646.950 204.600 648.150 219.600 ;
        RECT 656.400 217.050 657.450 286.950 ;
        RECT 664.950 283.950 667.050 289.050 ;
        RECT 670.950 286.950 676.050 289.050 ;
        RECT 667.950 277.950 670.050 280.050 ;
        RECT 664.950 262.950 667.050 265.050 ;
        RECT 658.950 256.950 661.050 262.050 ;
        RECT 665.400 253.050 666.450 262.950 ;
        RECT 668.400 259.050 669.450 277.950 ;
        RECT 677.400 274.050 678.450 292.950 ;
        RECT 679.950 289.950 685.050 292.050 ;
        RECT 685.950 280.950 688.050 286.050 ;
        RECT 676.950 273.450 679.050 274.050 ;
        RECT 674.400 272.400 679.050 273.450 ;
        RECT 667.950 256.950 670.050 259.050 ;
        RECT 674.400 256.050 675.450 272.400 ;
        RECT 676.950 271.950 679.050 272.400 ;
        RECT 682.950 256.950 685.050 262.050 ;
        RECT 673.950 253.950 676.050 256.050 ;
        RECT 679.950 253.950 682.050 256.050 ;
        RECT 664.950 250.950 667.050 253.050 ;
        RECT 661.950 238.950 664.050 241.050 ;
        RECT 676.950 238.950 679.050 241.050 ;
        RECT 662.400 217.050 663.450 238.950 ;
        RECT 677.400 229.050 678.450 238.950 ;
        RECT 676.950 226.950 679.050 229.050 ;
        RECT 655.950 214.950 658.050 217.050 ;
        RECT 661.950 214.950 664.050 217.050 ;
        RECT 667.950 214.950 673.050 217.050 ;
        RECT 655.950 208.950 658.050 211.050 ;
        RECT 664.950 208.950 670.050 211.050 ;
        RECT 649.950 207.450 654.000 208.050 ;
        RECT 649.950 205.950 654.450 207.450 ;
        RECT 646.950 202.500 649.050 204.600 ;
        RECT 643.950 187.950 646.050 190.050 ;
        RECT 640.950 181.950 643.050 184.050 ;
        RECT 641.400 178.050 642.450 181.950 ;
        RECT 640.950 175.950 643.050 178.050 ;
        RECT 637.950 151.950 640.050 154.050 ;
        RECT 644.400 148.050 645.450 187.950 ;
        RECT 653.400 184.050 654.450 205.950 ;
        RECT 649.950 182.400 654.450 184.050 ;
        RECT 649.950 181.950 654.000 182.400 ;
        RECT 656.400 178.050 657.450 208.950 ;
        RECT 680.400 187.050 681.450 253.950 ;
        RECT 683.400 253.050 684.450 256.950 ;
        RECT 689.400 256.050 690.450 298.950 ;
        RECT 691.950 289.950 697.050 292.050 ;
        RECT 698.400 283.050 699.450 319.950 ;
        RECT 706.950 310.950 709.050 313.050 ;
        RECT 707.400 295.050 708.450 310.950 ;
        RECT 700.950 292.950 703.050 295.050 ;
        RECT 706.950 292.950 709.050 295.050 ;
        RECT 697.950 280.950 700.050 283.050 ;
        RECT 701.400 280.050 702.450 292.950 ;
        RECT 700.950 277.950 703.050 280.050 ;
        RECT 701.400 274.050 702.450 277.950 ;
        RECT 700.950 271.950 703.050 274.050 ;
        RECT 706.950 259.050 709.050 262.050 ;
        RECT 710.400 259.200 711.450 352.950 ;
        RECT 713.400 328.050 714.450 361.800 ;
        RECT 715.950 337.950 718.050 340.050 ;
        RECT 712.950 325.950 715.050 328.050 ;
        RECT 716.400 319.050 717.450 337.950 ;
        RECT 718.950 331.950 721.050 334.050 ;
        RECT 715.950 316.950 718.050 319.050 ;
        RECT 719.400 313.050 720.450 331.950 ;
        RECT 718.950 310.950 721.050 313.050 ;
        RECT 715.950 304.950 718.050 307.050 ;
        RECT 712.950 295.950 715.050 298.050 ;
        RECT 713.400 292.050 714.450 295.950 ;
        RECT 712.950 289.950 715.050 292.050 ;
        RECT 716.400 289.200 717.450 304.950 ;
        RECT 715.950 287.100 718.050 289.200 ;
        RECT 719.400 289.050 720.450 310.950 ;
        RECT 728.400 301.050 729.450 385.950 ;
        RECT 731.400 367.050 732.450 388.950 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 730.950 364.950 733.050 367.050 ;
        RECT 730.950 349.950 733.050 352.050 ;
        RECT 731.400 334.050 732.450 349.950 ;
        RECT 734.400 340.050 735.450 367.950 ;
        RECT 737.400 346.050 738.450 428.400 ;
        RECT 740.400 388.050 741.450 452.400 ;
        RECT 749.400 451.050 750.450 466.950 ;
        RECT 767.400 451.050 768.450 466.950 ;
        RECT 778.950 460.950 781.050 463.050 ;
        RECT 748.950 445.950 751.050 451.050 ;
        RECT 754.950 447.450 757.050 451.050 ;
        RECT 757.950 448.950 763.050 451.050 ;
        RECT 766.950 448.950 769.050 451.050 ;
        RECT 772.950 448.950 775.050 451.050 ;
        RECT 754.950 447.000 759.450 447.450 ;
        RECT 755.400 446.400 760.050 447.000 ;
        RECT 742.950 439.950 745.050 442.050 ;
        RECT 743.400 394.050 744.450 439.950 ;
        RECT 749.400 427.050 750.450 445.950 ;
        RECT 757.950 442.950 760.050 446.400 ;
        RECT 773.400 445.050 774.450 448.950 ;
        RECT 779.400 445.050 780.450 460.950 ;
        RECT 782.400 451.050 783.450 481.800 ;
        RECT 785.400 475.050 786.450 496.950 ;
        RECT 797.400 496.050 798.450 523.950 ;
        RECT 814.950 520.950 817.050 523.050 ;
        RECT 805.950 511.950 808.050 514.050 ;
        RECT 796.950 493.950 799.050 496.050 ;
        RECT 787.950 484.950 790.050 490.050 ;
        RECT 797.400 489.450 798.450 493.950 ;
        RECT 806.400 493.050 807.450 511.950 ;
        RECT 815.400 499.050 816.450 520.950 ;
        RECT 823.950 505.950 826.050 508.050 ;
        RECT 814.950 496.950 817.050 499.050 ;
        RECT 817.950 493.950 823.050 496.050 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 794.400 489.000 798.450 489.450 ;
        RECT 793.950 488.400 798.450 489.000 ;
        RECT 808.950 489.450 811.050 490.050 ;
        RECT 814.950 489.450 817.050 490.050 ;
        RECT 808.950 488.400 817.050 489.450 ;
        RECT 793.950 484.950 796.050 488.400 ;
        RECT 808.950 487.950 811.050 488.400 ;
        RECT 814.950 487.950 817.050 488.400 ;
        RECT 802.950 484.950 805.050 487.050 ;
        RECT 784.950 472.950 787.050 475.050 ;
        RECT 795.000 456.450 799.050 457.050 ;
        RECT 794.400 454.950 799.050 456.450 ;
        RECT 781.950 448.950 784.050 451.050 ;
        RECT 763.950 442.950 769.050 445.050 ;
        RECT 769.950 442.950 772.050 445.050 ;
        RECT 772.950 442.950 775.050 445.050 ;
        RECT 779.400 443.400 784.050 445.050 ;
        RECT 780.000 442.950 784.050 443.400 ;
        RECT 770.400 430.050 771.450 442.950 ;
        RECT 769.950 427.950 772.050 430.050 ;
        RECT 748.950 424.950 751.050 427.050 ;
        RECT 766.950 422.400 769.050 424.500 ;
        RECT 787.950 422.400 790.050 424.500 ;
        RECT 745.950 415.950 748.050 421.050 ;
        RECT 751.950 412.950 754.050 418.050 ;
        RECT 757.950 417.450 762.000 418.050 ;
        RECT 757.950 415.950 762.450 417.450 ;
        RECT 745.950 409.950 751.050 412.050 ;
        RECT 754.950 406.950 757.050 412.050 ;
        RECT 761.400 406.050 762.450 415.950 ;
        RECT 760.950 403.950 763.050 406.050 ;
        RECT 767.700 402.600 768.900 422.400 ;
        RECT 772.950 409.950 775.050 415.050 ;
        RECT 778.950 412.950 781.050 415.050 ;
        RECT 766.950 400.500 769.050 402.600 ;
        RECT 742.950 391.950 745.050 394.050 ;
        RECT 739.950 385.950 742.050 388.050 ;
        RECT 772.950 385.950 775.050 388.050 ;
        RECT 742.950 380.400 745.050 382.500 ;
        RECT 763.950 381.300 766.050 383.400 ;
        RECT 743.700 360.600 744.900 380.400 ;
        RECT 754.950 376.950 757.050 379.050 ;
        RECT 763.950 377.700 765.150 381.300 ;
        RECT 755.400 370.050 756.450 376.950 ;
        RECT 763.950 375.600 766.050 377.700 ;
        RECT 748.950 364.950 751.050 370.050 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 742.950 358.500 745.050 360.600 ;
        RECT 755.400 352.050 756.450 367.950 ;
        RECT 763.950 360.600 765.150 375.600 ;
        RECT 766.950 366.450 771.000 367.050 ;
        RECT 766.950 364.950 771.450 366.450 ;
        RECT 770.400 361.050 771.450 364.950 ;
        RECT 763.950 358.500 766.050 360.600 ;
        RECT 769.950 358.950 772.050 361.050 ;
        RECT 773.400 355.050 774.450 385.950 ;
        RECT 779.400 379.050 780.450 412.950 ;
        RECT 787.950 407.400 789.150 422.400 ;
        RECT 790.950 415.950 793.050 421.050 ;
        RECT 781.950 403.950 784.050 406.050 ;
        RECT 787.950 405.300 790.050 407.400 ;
        RECT 778.950 376.950 781.050 379.050 ;
        RECT 782.400 370.050 783.450 403.950 ;
        RECT 787.950 401.700 789.150 405.300 ;
        RECT 787.950 399.600 790.050 401.700 ;
        RECT 794.400 400.050 795.450 454.950 ;
        RECT 796.950 448.950 802.050 451.050 ;
        RECT 803.400 448.050 804.450 484.950 ;
        RECT 808.950 481.950 814.050 484.050 ;
        RECT 808.950 475.950 811.050 478.050 ;
        RECT 805.950 451.950 808.050 454.050 ;
        RECT 802.950 445.950 805.050 448.050 ;
        RECT 796.950 421.950 799.050 424.050 ;
        RECT 793.950 397.950 796.050 400.050 ;
        RECT 784.950 388.950 787.050 391.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 772.950 352.950 775.050 355.050 ;
        RECT 754.950 349.950 757.050 352.050 ;
        RECT 766.950 349.950 769.050 352.050 ;
        RECT 736.950 343.950 739.050 346.050 ;
        RECT 754.950 344.400 757.050 346.500 ;
        RECT 733.950 337.950 736.050 340.050 ;
        RECT 739.950 334.950 742.050 340.050 ;
        RECT 745.950 339.450 750.000 340.050 ;
        RECT 745.950 337.950 750.450 339.450 ;
        RECT 730.950 331.950 733.050 334.050 ;
        RECT 733.950 331.950 739.050 334.050 ;
        RECT 742.950 331.950 745.050 334.050 ;
        RECT 743.400 328.050 744.450 331.950 ;
        RECT 742.950 325.950 745.050 328.050 ;
        RECT 727.950 298.950 730.050 301.050 ;
        RECT 739.950 298.950 742.050 301.050 ;
        RECT 724.950 292.950 727.050 298.050 ;
        RECT 730.950 294.450 735.000 295.050 ;
        RECT 730.950 292.950 735.450 294.450 ;
        RECT 734.400 289.050 735.450 292.950 ;
        RECT 719.400 287.400 724.050 289.050 ;
        RECT 720.000 286.950 724.050 287.400 ;
        RECT 727.950 286.950 730.050 289.050 ;
        RECT 733.950 286.950 736.050 289.050 ;
        RECT 715.950 283.800 718.050 285.900 ;
        RECT 716.400 265.050 717.450 283.800 ;
        RECT 724.950 268.950 727.050 271.050 ;
        RECT 715.950 262.950 718.050 265.050 ;
        RECT 712.950 259.950 715.050 262.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 706.800 258.000 709.050 259.050 ;
        RECT 706.800 256.950 708.900 258.000 ;
        RECT 710.100 257.100 712.200 259.200 ;
        RECT 688.950 253.950 691.050 256.050 ;
        RECT 683.400 251.400 688.050 253.050 ;
        RECT 684.000 250.950 688.050 251.400 ;
        RECT 691.950 250.950 697.050 253.050 ;
        RECT 695.400 247.050 696.450 250.950 ;
        RECT 694.950 244.950 697.050 247.050 ;
        RECT 698.400 229.050 699.450 256.950 ;
        RECT 703.950 253.950 706.050 256.050 ;
        RECT 700.950 247.950 703.050 250.050 ;
        RECT 688.950 226.950 691.050 229.050 ;
        RECT 697.950 226.950 700.050 229.050 ;
        RECT 682.950 217.950 685.050 220.050 ;
        RECT 683.400 214.050 684.450 217.950 ;
        RECT 689.400 217.050 690.450 226.950 ;
        RECT 701.400 226.050 702.450 247.950 ;
        RECT 704.400 241.050 705.450 253.950 ;
        RECT 709.950 250.950 712.050 255.900 ;
        RECT 713.400 250.050 714.450 259.950 ;
        RECT 715.950 256.950 718.050 259.050 ;
        RECT 718.950 256.950 721.050 259.050 ;
        RECT 712.950 247.950 715.050 250.050 ;
        RECT 703.950 238.950 706.050 241.050 ;
        RECT 700.950 223.950 703.050 226.050 ;
        RECT 691.950 220.950 694.050 223.050 ;
        RECT 688.950 214.950 691.050 217.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 664.950 181.950 667.050 187.050 ;
        RECT 679.950 184.950 682.050 187.050 ;
        RECT 673.950 181.950 676.050 184.050 ;
        RECT 688.950 181.950 691.050 187.050 ;
        RECT 652.950 176.400 657.450 178.050 ;
        RECT 652.950 175.950 657.000 176.400 ;
        RECT 667.950 175.950 673.050 178.050 ;
        RECT 643.950 145.950 646.050 148.050 ;
        RECT 653.400 142.050 654.450 175.950 ;
        RECT 674.400 166.050 675.450 181.950 ;
        RECT 676.950 175.950 682.050 178.050 ;
        RECT 685.950 175.950 688.050 181.050 ;
        RECT 673.950 163.950 676.050 166.050 ;
        RECT 686.400 163.050 687.450 175.950 ;
        RECT 692.400 175.050 693.450 220.950 ;
        RECT 697.950 214.050 700.050 217.050 ;
        RECT 703.950 214.950 706.050 217.050 ;
        RECT 706.950 214.950 712.050 217.050 ;
        RECT 696.000 213.450 700.050 214.050 ;
        RECT 695.400 211.950 700.050 213.450 ;
        RECT 695.400 208.050 696.450 211.950 ;
        RECT 704.400 208.050 705.450 214.950 ;
        RECT 694.800 205.950 696.900 208.050 ;
        RECT 697.950 205.950 700.050 208.050 ;
        RECT 703.950 205.950 706.050 208.050 ;
        RECT 712.950 205.950 715.050 211.050 ;
        RECT 694.950 181.950 697.050 184.050 ;
        RECT 695.400 178.050 696.450 181.950 ;
        RECT 698.400 181.200 699.450 205.950 ;
        RECT 703.950 199.950 706.050 202.050 ;
        RECT 704.400 184.050 705.450 199.950 ;
        RECT 709.950 184.950 712.050 187.050 ;
        RECT 697.950 179.100 700.050 181.200 ;
        RECT 703.950 178.950 706.050 184.050 ;
        RECT 710.400 178.050 711.450 184.950 ;
        RECT 716.400 183.450 717.450 256.950 ;
        RECT 719.400 211.050 720.450 256.950 ;
        RECT 725.400 253.050 726.450 268.950 ;
        RECT 728.400 256.050 729.450 286.950 ;
        RECT 740.400 265.050 741.450 298.950 ;
        RECT 743.400 286.050 744.450 325.950 ;
        RECT 745.950 301.950 748.050 304.050 ;
        RECT 746.400 295.050 747.450 301.950 ;
        RECT 749.400 298.050 750.450 337.950 ;
        RECT 755.700 324.600 756.900 344.400 ;
        RECT 767.400 337.050 768.450 349.950 ;
        RECT 785.400 349.050 786.450 388.950 ;
        RECT 790.950 379.950 793.050 382.050 ;
        RECT 791.400 373.050 792.450 379.950 ;
        RECT 797.400 375.450 798.450 421.950 ;
        RECT 799.950 415.950 805.050 418.050 ;
        RECT 800.400 376.200 801.450 415.950 ;
        RECT 802.950 409.950 805.050 412.050 ;
        RECT 803.400 406.050 804.450 409.950 ;
        RECT 802.950 403.950 805.050 406.050 ;
        RECT 806.400 402.450 807.450 451.950 ;
        RECT 803.400 401.400 807.450 402.450 ;
        RECT 803.400 391.050 804.450 401.400 ;
        RECT 805.950 397.950 808.050 400.050 ;
        RECT 802.950 388.950 805.050 391.050 ;
        RECT 802.950 379.950 805.050 382.050 ;
        RECT 794.400 374.400 798.450 375.450 ;
        RECT 790.950 370.950 793.050 373.050 ;
        RECT 790.950 361.950 793.050 364.050 ;
        RECT 784.950 346.950 787.050 349.050 ;
        RECT 775.950 344.400 778.050 346.500 ;
        RECT 760.950 331.950 763.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 754.950 322.500 757.050 324.600 ;
        RECT 757.950 316.950 760.050 319.050 ;
        RECT 748.950 295.950 751.050 298.050 ;
        RECT 758.400 295.050 759.450 316.950 ;
        RECT 763.950 301.950 766.050 304.050 ;
        RECT 745.950 292.950 748.050 295.050 ;
        RECT 751.950 289.950 754.050 295.050 ;
        RECT 757.950 292.950 760.050 295.050 ;
        RECT 758.400 289.050 759.450 292.950 ;
        RECT 754.950 287.400 759.450 289.050 ;
        RECT 754.950 286.950 759.000 287.400 ;
        RECT 742.950 283.950 745.050 286.050 ;
        RECT 751.950 283.950 754.050 286.050 ;
        RECT 739.950 262.950 742.050 265.050 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 727.950 253.950 730.050 256.050 ;
        RECT 734.400 253.050 735.450 256.950 ;
        RECT 724.950 250.950 727.050 253.050 ;
        RECT 730.950 251.400 735.450 253.050 ;
        RECT 730.950 250.950 735.000 251.400 ;
        RECT 742.950 250.950 745.050 256.050 ;
        RECT 748.950 250.950 751.050 253.050 ;
        RECT 749.400 247.050 750.450 250.950 ;
        RECT 748.950 244.950 751.050 247.050 ;
        RECT 752.400 241.050 753.450 283.950 ;
        RECT 760.950 277.950 763.050 280.050 ;
        RECT 757.950 265.950 760.050 268.050 ;
        RECT 754.950 262.950 757.050 265.050 ;
        RECT 730.950 238.950 733.050 241.050 ;
        RECT 751.950 238.950 754.050 241.050 ;
        RECT 731.400 223.050 732.450 238.950 ;
        RECT 745.950 225.300 748.050 227.400 ;
        RECT 730.950 217.950 733.050 223.050 ;
        RECT 746.850 221.700 748.050 225.300 ;
        RECT 736.950 217.950 739.050 220.050 ;
        RECT 739.950 217.950 742.050 220.050 ;
        RECT 745.950 219.600 748.050 221.700 ;
        RECT 755.400 220.050 756.450 262.950 ;
        RECT 758.400 220.050 759.450 265.950 ;
        RECT 761.400 265.050 762.450 277.950 ;
        RECT 764.400 268.050 765.450 301.950 ;
        RECT 770.400 292.050 771.450 334.950 ;
        RECT 775.950 329.400 777.150 344.400 ;
        RECT 784.950 340.950 787.050 343.050 ;
        RECT 778.950 334.950 781.050 340.050 ;
        RECT 775.950 327.300 778.050 329.400 ;
        RECT 775.950 323.700 777.150 327.300 ;
        RECT 775.950 321.600 778.050 323.700 ;
        RECT 775.950 293.100 778.050 298.050 ;
        RECT 769.950 289.950 775.050 292.050 ;
        RECT 775.950 286.950 778.050 291.900 ;
        RECT 785.400 291.450 786.450 340.950 ;
        RECT 791.400 337.050 792.450 361.950 ;
        RECT 794.400 339.450 795.450 374.400 ;
        RECT 799.950 374.100 802.050 376.200 ;
        RECT 803.400 373.050 804.450 379.950 ;
        RECT 796.950 370.950 799.050 373.050 ;
        RECT 801.000 372.900 804.450 373.050 ;
        RECT 799.950 371.250 804.450 372.900 ;
        RECT 799.950 370.950 804.000 371.250 ;
        RECT 797.400 346.050 798.450 370.950 ;
        RECT 799.950 370.800 802.050 370.950 ;
        RECT 806.400 367.050 807.450 397.950 ;
        RECT 809.400 394.050 810.450 475.950 ;
        RECT 811.950 460.950 814.050 463.050 ;
        RECT 808.950 391.950 811.050 394.050 ;
        RECT 812.400 388.050 813.450 460.950 ;
        RECT 817.950 442.950 820.050 445.050 ;
        RECT 818.400 436.050 819.450 442.950 ;
        RECT 817.950 433.950 820.050 436.050 ;
        RECT 824.400 424.050 825.450 505.950 ;
        RECT 827.400 478.050 828.450 646.950 ;
        RECT 830.400 574.050 831.450 691.950 ;
        RECT 829.950 571.950 832.050 574.050 ;
        RECT 829.950 532.950 832.050 535.050 ;
        RECT 826.950 475.950 829.050 478.050 ;
        RECT 830.400 463.050 831.450 532.950 ;
        RECT 829.950 460.950 832.050 463.050 ;
        RECT 823.950 421.950 826.050 424.050 ;
        RECT 826.950 412.950 829.050 415.050 ;
        RECT 817.950 406.950 820.050 409.050 ;
        RECT 814.950 403.950 817.050 406.050 ;
        RECT 811.950 385.950 814.050 388.050 ;
        RECT 811.950 379.950 814.050 382.050 ;
        RECT 812.400 373.050 813.450 379.950 ;
        RECT 815.400 376.050 816.450 403.950 ;
        RECT 818.400 400.050 819.450 406.950 ;
        RECT 823.950 403.950 826.050 409.050 ;
        RECT 817.950 397.950 820.050 400.050 ;
        RECT 827.400 396.450 828.450 412.950 ;
        RECT 824.400 395.400 828.450 396.450 ;
        RECT 824.400 379.050 825.450 395.400 ;
        RECT 826.950 391.950 829.050 394.050 ;
        RECT 817.950 376.950 820.050 379.050 ;
        RECT 823.950 376.950 826.050 379.050 ;
        RECT 814.950 373.950 817.050 376.050 ;
        RECT 818.400 373.050 819.450 376.950 ;
        RECT 820.950 373.950 823.050 376.050 ;
        RECT 811.950 370.950 814.050 373.050 ;
        RECT 817.950 370.950 820.050 373.050 ;
        RECT 802.950 364.950 805.050 367.050 ;
        RECT 806.400 365.400 811.050 367.050 ;
        RECT 807.000 364.950 811.050 365.400 ;
        RECT 814.950 364.950 817.050 370.050 ;
        RECT 803.400 361.050 804.450 364.950 ;
        RECT 802.950 358.950 805.050 361.050 ;
        RECT 799.950 346.950 802.050 349.050 ;
        RECT 796.950 343.950 799.050 346.050 ;
        RECT 794.400 338.400 798.450 339.450 ;
        RECT 787.950 331.950 790.050 337.050 ;
        RECT 791.400 334.950 796.050 337.050 ;
        RECT 785.400 290.400 789.450 291.450 ;
        RECT 784.950 286.950 787.050 289.050 ;
        RECT 769.950 283.950 772.050 286.050 ;
        RECT 763.950 265.950 766.050 268.050 ;
        RECT 760.950 262.950 763.050 265.050 ;
        RECT 763.950 256.950 766.050 262.050 ;
        RECT 770.400 256.050 771.450 283.950 ;
        RECT 781.950 268.950 784.050 271.050 ;
        RECT 775.950 259.950 778.050 262.050 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 769.950 253.950 772.050 256.050 ;
        RECT 766.950 224.400 769.050 226.500 ;
        RECT 721.950 211.950 724.050 214.050 ;
        RECT 733.950 211.950 736.050 217.050 ;
        RECT 718.950 208.950 721.050 211.050 ;
        RECT 713.400 182.400 717.450 183.450 ;
        RECT 695.400 177.900 699.000 178.050 ;
        RECT 695.400 176.250 700.050 177.900 ;
        RECT 696.000 175.950 700.050 176.250 ;
        RECT 709.950 175.950 712.050 178.050 ;
        RECT 697.950 175.800 700.050 175.950 ;
        RECT 691.950 172.950 694.050 175.050 ;
        RECT 697.950 172.800 700.050 174.900 ;
        RECT 685.950 160.950 688.050 163.050 ;
        RECT 694.950 154.950 697.050 157.050 ;
        RECT 658.950 147.300 661.050 149.400 ;
        RECT 659.850 143.700 661.050 147.300 ;
        RECT 679.950 146.400 682.050 148.500 ;
        RECT 634.950 139.950 637.050 142.050 ;
        RECT 637.950 139.950 643.050 142.050 ;
        RECT 646.950 139.950 652.050 142.050 ;
        RECT 652.950 139.950 655.050 142.050 ;
        RECT 658.950 141.600 661.050 143.700 ;
        RECT 635.400 106.200 636.450 139.950 ;
        RECT 643.950 133.950 646.050 136.050 ;
        RECT 634.950 106.050 637.050 106.200 ;
        RECT 633.000 105.600 637.050 106.050 ;
        RECT 632.400 104.100 637.050 105.600 ;
        RECT 632.400 103.950 636.000 104.100 ;
        RECT 640.950 103.950 643.050 106.050 ;
        RECT 632.400 79.050 633.450 103.950 ;
        RECT 634.950 100.050 637.050 102.900 ;
        RECT 634.950 99.000 640.050 100.050 ;
        RECT 635.400 98.400 640.050 99.000 ;
        RECT 636.000 97.950 640.050 98.400 ;
        RECT 641.400 85.050 642.450 103.950 ;
        RECT 644.400 100.050 645.450 133.950 ;
        RECT 652.950 130.950 658.050 133.050 ;
        RECT 653.400 127.050 654.450 130.950 ;
        RECT 652.950 124.950 655.050 127.050 ;
        RECT 659.850 126.600 661.050 141.600 ;
        RECT 673.950 136.950 676.050 142.050 ;
        RECT 667.950 133.950 670.050 136.050 ;
        RECT 658.950 124.500 661.050 126.600 ;
        RECT 664.950 120.450 667.050 124.050 ;
        RECT 662.400 120.000 667.050 120.450 ;
        RECT 662.400 119.400 666.450 120.000 ;
        RECT 662.400 106.050 663.450 119.400 ;
        RECT 668.400 118.050 669.450 133.950 ;
        RECT 680.100 126.600 681.300 146.400 ;
        RECT 688.950 139.950 691.050 142.050 ;
        RECT 689.400 133.050 690.450 139.950 ;
        RECT 691.950 136.950 694.050 139.050 ;
        RECT 695.400 138.450 696.450 154.950 ;
        RECT 698.400 142.050 699.450 172.800 ;
        RECT 713.400 145.050 714.450 182.400 ;
        RECT 722.400 181.050 723.450 211.950 ;
        RECT 737.400 211.050 738.450 217.950 ;
        RECT 736.950 208.950 739.050 211.050 ;
        RECT 737.400 193.050 738.450 208.950 ;
        RECT 736.950 190.950 739.050 193.050 ;
        RECT 727.950 184.950 730.050 187.050 ;
        RECT 715.950 175.950 718.050 181.050 ;
        RECT 721.950 178.950 724.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 715.950 163.950 718.050 166.050 ;
        RECT 703.950 142.950 706.050 145.050 ;
        RECT 712.950 142.950 715.050 145.050 ;
        RECT 697.950 141.450 702.000 142.050 ;
        RECT 697.950 139.950 702.450 141.450 ;
        RECT 695.400 137.400 699.450 138.450 ;
        RECT 688.950 130.950 691.050 133.050 ;
        RECT 692.400 130.050 693.450 136.950 ;
        RECT 691.950 127.950 694.050 130.050 ;
        RECT 679.950 124.500 682.050 126.600 ;
        RECT 667.950 115.950 670.050 118.050 ;
        RECT 679.950 115.950 682.050 118.050 ;
        RECT 664.950 108.450 667.050 112.050 ;
        RECT 670.950 110.400 673.050 112.500 ;
        RECT 664.950 108.000 669.450 108.450 ;
        RECT 665.400 107.400 670.050 108.000 ;
        RECT 661.950 103.950 664.050 106.050 ;
        RECT 667.950 103.950 670.050 107.400 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 643.950 97.950 646.050 100.050 ;
        RECT 653.400 88.050 654.450 100.950 ;
        RECT 671.850 95.400 673.050 110.400 ;
        RECT 680.400 106.050 681.450 115.950 ;
        RECT 691.950 110.400 694.050 112.500 ;
        RECT 679.950 100.950 682.050 106.050 ;
        RECT 670.950 93.300 673.050 95.400 ;
        RECT 671.850 89.700 673.050 93.300 ;
        RECT 652.950 85.950 655.050 88.050 ;
        RECT 670.950 87.600 673.050 89.700 ;
        RECT 640.950 82.950 643.050 85.050 ;
        RECT 631.950 76.950 634.050 79.050 ;
        RECT 616.950 61.950 619.050 64.050 ;
        RECT 628.950 62.100 631.050 64.200 ;
        RECT 649.950 61.950 652.050 64.050 ;
        RECT 622.950 58.950 625.050 61.050 ;
        RECT 607.950 53.400 612.450 55.050 ;
        RECT 607.950 52.950 612.000 53.400 ;
        RECT 619.950 52.950 622.050 55.050 ;
        RECT 583.950 46.500 586.050 48.600 ;
        RECT 604.950 46.500 607.050 48.600 ;
        RECT 577.950 40.950 580.050 43.050 ;
        RECT 620.400 37.050 621.450 52.950 ;
        RECT 607.950 34.950 610.050 37.050 ;
        RECT 619.950 34.950 622.050 37.050 ;
        RECT 574.950 31.950 577.050 34.050 ;
        RECT 592.950 32.400 595.050 34.500 ;
        RECT 565.950 25.950 571.050 28.050 ;
        RECT 571.950 25.950 574.050 28.050 ;
        RECT 559.950 19.950 562.050 22.050 ;
        RECT 565.950 19.950 568.050 22.050 ;
        RECT 550.950 16.950 553.050 19.050 ;
        RECT 566.400 16.050 567.450 19.950 ;
        RECT 569.400 19.050 570.450 25.950 ;
        RECT 575.400 25.050 576.450 31.950 ;
        RECT 574.950 22.950 577.050 25.050 ;
        RECT 577.950 24.450 580.050 25.050 ;
        RECT 577.950 24.000 588.450 24.450 ;
        RECT 577.950 23.400 589.050 24.000 ;
        RECT 577.950 22.950 580.050 23.400 ;
        RECT 568.950 16.950 571.050 19.050 ;
        RECT 571.950 16.950 577.050 19.050 ;
        RECT 580.950 16.950 583.050 22.050 ;
        RECT 586.950 19.950 589.050 23.400 ;
        RECT 589.950 22.950 592.050 28.050 ;
        RECT 593.850 17.400 595.050 32.400 ;
        RECT 601.950 22.950 604.050 28.050 ;
        RECT 608.400 22.050 609.450 34.950 ;
        RECT 613.950 32.400 616.050 34.500 ;
        RECT 607.950 19.950 610.050 22.050 ;
        RECT 565.950 13.950 568.050 16.050 ;
        RECT 592.950 15.300 595.050 17.400 ;
        RECT 593.850 11.700 595.050 15.300 ;
        RECT 614.100 12.600 615.300 32.400 ;
        RECT 623.400 25.050 624.450 58.950 ;
        RECT 628.950 55.950 631.050 60.900 ;
        RECT 643.950 58.950 646.050 61.050 ;
        RECT 644.400 55.050 645.450 58.950 ;
        RECT 650.400 58.050 651.450 61.950 ;
        RECT 653.400 61.050 654.450 85.950 ;
        RECT 680.400 70.050 681.450 100.950 ;
        RECT 685.950 97.950 688.050 103.050 ;
        RECT 692.100 90.600 693.300 110.400 ;
        RECT 691.950 88.500 694.050 90.600 ;
        RECT 682.950 70.950 685.050 73.050 ;
        RECT 673.950 67.950 676.050 70.050 ;
        RECT 679.950 67.950 682.050 70.050 ;
        RECT 652.950 58.950 655.050 61.050 ;
        RECT 649.950 55.950 652.050 58.050 ;
        RECT 661.950 55.950 664.050 61.050 ;
        RECT 631.950 49.950 634.050 55.050 ;
        RECT 643.950 52.950 646.050 55.050 ;
        RECT 649.950 49.950 652.050 52.050 ;
        RECT 667.950 49.950 670.050 55.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 646.950 22.950 649.050 25.050 ;
        RECT 626.400 19.050 627.450 22.950 ;
        RECT 625.950 13.950 628.050 19.050 ;
        RECT 631.950 16.950 637.050 19.050 ;
        RECT 647.400 13.050 648.450 22.950 ;
        RECT 650.400 19.050 651.450 49.950 ;
        RECT 664.950 32.400 667.050 34.500 ;
        RECT 655.950 22.950 658.050 25.050 ;
        RECT 661.950 22.950 664.050 28.050 ;
        RECT 656.400 19.050 657.450 22.950 ;
        RECT 649.950 16.950 652.050 19.050 ;
        RECT 655.950 16.950 658.050 19.050 ;
        RECT 665.850 17.400 667.050 32.400 ;
        RECT 674.400 28.050 675.450 67.950 ;
        RECT 683.400 64.050 684.450 70.950 ;
        RECT 682.950 61.950 685.050 64.050 ;
        RECT 688.950 61.950 691.050 67.050 ;
        RECT 698.400 61.050 699.450 137.400 ;
        RECT 701.400 124.050 702.450 139.950 ;
        RECT 700.950 121.950 703.050 124.050 ;
        RECT 704.400 106.050 705.450 142.950 ;
        RECT 706.950 134.100 709.050 139.050 ;
        RECT 709.950 136.950 715.050 139.050 ;
        RECT 706.950 127.950 709.050 132.900 ;
        RECT 716.400 112.050 717.450 163.950 ;
        RECT 718.950 142.950 721.050 145.050 ;
        RECT 719.400 139.050 720.450 142.950 ;
        RECT 725.400 139.050 726.450 178.950 ;
        RECT 728.400 145.050 729.450 184.950 ;
        RECT 733.950 178.950 736.050 184.050 ;
        RECT 740.400 180.450 741.450 217.950 ;
        RECT 742.950 205.950 745.050 211.050 ;
        RECT 746.850 204.600 748.050 219.600 ;
        RECT 754.800 217.950 756.900 220.050 ;
        RECT 758.100 217.950 760.200 220.050 ;
        RECT 751.950 211.950 757.050 214.050 ;
        RECT 760.950 211.950 763.050 217.050 ;
        RECT 745.950 202.500 748.050 204.600 ;
        RECT 751.950 187.950 754.050 190.050 ;
        RECT 752.400 184.050 753.450 187.950 ;
        RECT 755.400 184.050 756.450 211.950 ;
        RECT 767.100 204.600 768.300 224.400 ;
        RECT 766.950 202.500 769.050 204.600 ;
        RECT 773.400 202.050 774.450 256.950 ;
        RECT 772.950 199.950 775.050 202.050 ;
        RECT 763.950 196.950 766.050 199.050 ;
        RECT 751.950 181.950 754.050 184.050 ;
        RECT 754.950 181.950 757.050 184.050 ;
        RECT 759.000 183.450 763.050 184.050 ;
        RECT 758.400 181.950 763.050 183.450 ;
        RECT 737.400 179.400 741.450 180.450 ;
        RECT 737.400 169.050 738.450 179.400 ;
        RECT 742.950 175.950 745.050 178.050 ;
        RECT 754.950 175.950 757.050 178.050 ;
        RECT 736.950 166.950 739.050 169.050 ;
        RECT 736.950 160.950 739.050 163.050 ;
        RECT 727.950 142.950 730.050 145.050 ;
        RECT 737.400 139.050 738.450 160.950 ;
        RECT 743.400 145.050 744.450 175.950 ;
        RECT 742.950 142.950 745.050 145.050 ;
        RECT 718.950 136.950 721.050 139.050 ;
        RECT 724.950 136.950 727.050 139.050 ;
        RECT 729.000 138.450 733.050 139.050 ;
        RECT 728.400 136.950 733.050 138.450 ;
        RECT 736.950 136.950 739.050 139.050 ;
        RECT 721.950 130.950 727.050 133.050 ;
        RECT 724.950 115.950 727.050 118.050 ;
        RECT 715.950 109.950 718.050 112.050 ;
        RECT 703.950 103.950 706.050 106.050 ;
        RECT 709.950 100.950 712.050 106.050 ;
        RECT 715.950 101.100 718.050 106.050 ;
        RECT 721.950 103.950 724.050 106.050 ;
        RECT 722.400 100.050 723.450 103.950 ;
        RECT 706.950 94.950 709.050 100.050 ;
        RECT 712.950 99.900 717.000 100.050 ;
        RECT 712.950 97.950 718.050 99.900 ;
        RECT 721.950 97.950 724.050 100.050 ;
        RECT 715.950 97.800 718.050 97.950 ;
        RECT 697.950 58.950 700.050 61.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 686.400 46.050 687.450 55.950 ;
        RECT 707.400 52.050 708.450 94.950 ;
        RECT 725.400 79.050 726.450 115.950 ;
        RECT 724.950 76.950 727.050 79.050 ;
        RECT 724.950 70.950 727.050 73.050 ;
        RECT 715.950 58.950 718.050 64.050 ;
        RECT 721.950 58.950 724.050 64.050 ;
        RECT 725.400 55.050 726.450 70.950 ;
        RECT 728.400 67.050 729.450 136.950 ;
        RECT 743.400 133.050 744.450 142.950 ;
        RECT 755.400 139.050 756.450 175.950 ;
        RECT 758.400 157.050 759.450 181.950 ;
        RECT 764.400 178.050 765.450 196.950 ;
        RECT 776.400 190.050 777.450 259.950 ;
        RECT 782.400 256.050 783.450 268.950 ;
        RECT 785.400 262.050 786.450 286.950 ;
        RECT 788.400 264.450 789.450 290.400 ;
        RECT 791.400 271.050 792.450 334.950 ;
        RECT 797.400 313.050 798.450 338.400 ;
        RECT 796.950 310.950 799.050 313.050 ;
        RECT 800.400 304.050 801.450 346.950 ;
        RECT 803.400 334.050 804.450 358.950 ;
        RECT 811.950 343.950 814.050 346.050 ;
        RECT 805.950 340.950 808.050 343.050 ;
        RECT 806.400 337.050 807.450 340.950 ;
        RECT 812.400 337.050 813.450 343.950 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 821.400 334.050 822.450 373.950 ;
        RECT 802.950 331.950 805.050 334.050 ;
        RECT 808.950 331.950 811.050 334.050 ;
        RECT 820.950 331.950 823.050 334.050 ;
        RECT 802.950 310.950 805.050 313.050 ;
        RECT 799.950 301.950 802.050 304.050 ;
        RECT 796.950 294.450 799.050 298.050 ;
        RECT 799.950 295.950 802.050 298.050 ;
        RECT 794.400 293.400 799.050 294.450 ;
        RECT 790.950 268.950 793.050 271.050 ;
        RECT 788.400 263.400 792.450 264.450 ;
        RECT 785.400 261.000 790.050 262.050 ;
        RECT 784.950 259.950 790.050 261.000 ;
        RECT 784.950 257.100 787.050 259.950 ;
        RECT 791.400 256.050 792.450 263.400 ;
        RECT 782.400 255.900 786.000 256.050 ;
        RECT 782.400 254.250 787.050 255.900 ;
        RECT 783.000 253.950 787.050 254.250 ;
        RECT 790.950 253.950 793.050 256.050 ;
        RECT 784.950 253.800 787.050 253.950 ;
        RECT 791.400 220.200 792.450 253.950 ;
        RECT 778.950 215.100 781.050 220.050 ;
        RECT 781.950 217.950 787.050 220.050 ;
        RECT 790.950 218.100 793.050 220.200 ;
        RECT 790.950 214.800 793.050 216.900 ;
        RECT 780.000 213.900 784.050 214.050 ;
        RECT 778.950 211.950 784.050 213.900 ;
        RECT 778.950 211.800 781.050 211.950 ;
        RECT 787.950 208.950 790.050 211.050 ;
        RECT 769.950 187.950 772.050 190.050 ;
        RECT 775.950 187.950 778.050 190.050 ;
        RECT 763.950 172.950 766.050 178.050 ;
        RECT 757.950 154.950 760.050 157.050 ;
        RECT 766.950 148.950 769.050 151.050 ;
        RECT 745.950 136.950 751.050 139.050 ;
        RECT 754.950 136.950 757.050 139.050 ;
        RECT 767.400 136.200 768.450 148.950 ;
        RECT 770.400 139.050 771.450 187.950 ;
        RECT 772.950 184.950 775.050 187.050 ;
        RECT 773.400 142.050 774.450 184.950 ;
        RECT 778.950 178.950 781.050 184.050 ;
        RECT 778.950 172.950 784.050 175.050 ;
        RECT 788.400 174.450 789.450 208.950 ;
        RECT 791.400 187.050 792.450 214.800 ;
        RECT 794.400 199.050 795.450 293.400 ;
        RECT 796.950 292.950 799.050 293.400 ;
        RECT 800.400 274.050 801.450 295.950 ;
        RECT 803.400 277.050 804.450 310.950 ;
        RECT 809.400 301.050 810.450 331.950 ;
        RECT 805.950 298.950 808.050 301.050 ;
        RECT 806.400 292.200 807.450 298.950 ;
        RECT 808.950 295.950 811.050 301.050 ;
        RECT 817.950 298.950 820.050 301.050 ;
        RECT 818.400 295.050 819.450 298.950 ;
        RECT 811.950 292.950 817.050 295.050 ;
        RECT 818.400 293.400 823.050 295.050 ;
        RECT 819.000 292.950 823.050 293.400 ;
        RECT 805.950 290.100 808.050 292.200 ;
        RECT 805.950 286.800 808.050 288.900 ;
        RECT 808.950 286.950 814.050 289.050 ;
        RECT 817.950 286.950 820.050 289.050 ;
        RECT 806.400 283.050 807.450 286.800 ;
        RECT 805.950 280.950 808.050 283.050 ;
        RECT 802.950 274.950 805.050 277.050 ;
        RECT 799.950 271.950 802.050 274.050 ;
        RECT 799.950 266.400 802.050 268.500 ;
        RECT 796.950 259.950 799.050 265.050 ;
        RECT 800.850 251.400 802.050 266.400 ;
        RECT 799.950 249.300 802.050 251.400 ;
        RECT 800.850 245.700 802.050 249.300 ;
        RECT 799.950 243.600 802.050 245.700 ;
        RECT 796.950 217.950 799.050 220.050 ;
        RECT 797.400 211.050 798.450 217.950 ;
        RECT 806.400 217.050 807.450 280.950 ;
        RECT 811.950 274.950 814.050 277.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 805.950 214.950 808.050 217.050 ;
        RECT 796.950 208.950 799.050 211.050 ;
        RECT 793.950 196.950 796.050 199.050 ;
        RECT 796.950 188.400 799.050 190.500 ;
        RECT 790.950 184.950 793.050 187.050 ;
        RECT 788.400 173.400 792.450 174.450 ;
        RECT 787.950 169.950 790.050 172.050 ;
        RECT 775.950 160.950 778.050 163.050 ;
        RECT 772.950 139.950 775.050 142.050 ;
        RECT 776.400 139.050 777.450 160.950 ;
        RECT 788.400 154.050 789.450 169.950 ;
        RECT 787.950 151.950 790.050 154.050 ;
        RECT 784.950 150.450 789.000 151.050 ;
        RECT 784.950 148.950 789.450 150.450 ;
        RECT 784.950 142.950 787.050 145.050 ;
        RECT 788.400 144.450 789.450 148.950 ;
        RECT 791.400 148.050 792.450 173.400 ;
        RECT 797.700 168.600 798.900 188.400 ;
        RECT 809.400 184.050 810.450 256.950 ;
        RECT 812.400 211.200 813.450 274.950 ;
        RECT 818.400 273.450 819.450 286.950 ;
        RECT 815.400 272.400 819.450 273.450 ;
        RECT 815.400 256.050 816.450 272.400 ;
        RECT 820.950 266.400 823.050 268.500 ;
        RECT 814.950 253.950 817.050 256.050 ;
        RECT 821.100 246.600 822.300 266.400 ;
        RECT 820.950 244.500 823.050 246.600 ;
        RECT 811.950 209.100 814.050 211.200 ;
        RECT 817.950 188.400 820.050 190.500 ;
        RECT 802.950 175.950 805.050 181.050 ;
        RECT 808.950 178.950 811.050 184.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 796.950 166.500 799.050 168.600 ;
        RECT 805.950 166.950 808.050 169.050 ;
        RECT 790.950 145.950 793.050 148.050 ;
        RECT 796.950 145.950 799.050 148.050 ;
        RECT 788.400 144.000 795.450 144.450 ;
        RECT 788.400 143.400 796.050 144.000 ;
        RECT 785.400 139.050 786.450 142.950 ;
        RECT 790.950 139.950 793.050 142.050 ;
        RECT 793.950 139.950 796.050 143.400 ;
        RECT 769.950 136.950 772.050 139.050 ;
        RECT 775.950 136.950 778.050 139.050 ;
        RECT 784.950 136.950 787.050 139.050 ;
        RECT 766.950 134.100 769.050 136.200 ;
        RECT 791.400 136.050 792.450 139.950 ;
        RECT 730.950 130.950 736.050 133.050 ;
        RECT 739.950 131.400 744.450 133.050 ;
        RECT 739.950 130.950 744.000 131.400 ;
        RECT 748.950 130.950 751.050 133.050 ;
        RECT 739.950 118.950 742.050 121.050 ;
        RECT 736.950 103.950 739.050 109.050 ;
        RECT 733.950 94.950 736.050 100.050 ;
        RECT 740.400 85.050 741.450 118.950 ;
        RECT 745.950 109.950 748.050 112.050 ;
        RECT 746.400 100.050 747.450 109.950 ;
        RECT 749.400 109.050 750.450 130.950 ;
        RECT 751.950 127.950 754.050 133.050 ;
        RECT 757.950 130.950 760.050 133.050 ;
        RECT 748.950 103.950 751.050 109.050 ;
        RECT 751.950 100.950 757.050 103.050 ;
        RECT 745.950 97.950 748.050 100.050 ;
        RECT 739.950 82.950 742.050 85.050 ;
        RECT 745.950 76.950 748.050 79.050 ;
        RECT 730.950 67.950 733.050 70.050 ;
        RECT 742.950 67.950 745.050 70.050 ;
        RECT 727.950 64.950 730.050 67.050 ;
        RECT 731.400 64.050 732.450 67.950 ;
        RECT 730.950 61.950 733.050 64.050 ;
        RECT 736.950 61.950 739.050 64.050 ;
        RECT 737.400 58.050 738.450 61.950 ;
        RECT 727.950 55.950 733.050 58.050 ;
        RECT 736.950 55.950 739.050 58.050 ;
        RECT 709.950 52.950 712.050 55.050 ;
        RECT 724.950 52.950 727.050 55.050 ;
        RECT 706.950 49.950 709.050 52.050 ;
        RECT 685.950 43.950 688.050 46.050 ;
        RECT 685.950 32.400 688.050 34.500 ;
        RECT 710.400 33.450 711.450 52.950 ;
        RECT 739.950 43.950 742.050 46.050 ;
        RECT 707.400 32.400 711.450 33.450 ;
        RECT 673.950 22.950 676.050 28.050 ;
        RECT 679.950 19.950 682.050 25.050 ;
        RECT 664.950 15.300 667.050 17.400 ;
        RECT 592.950 9.600 595.050 11.700 ;
        RECT 613.950 10.500 616.050 12.600 ;
        RECT 646.950 10.950 649.050 13.050 ;
        RECT 665.850 11.700 667.050 15.300 ;
        RECT 686.100 12.600 687.300 32.400 ;
        RECT 694.950 25.950 697.050 28.050 ;
        RECT 695.400 22.050 696.450 25.950 ;
        RECT 707.400 22.050 708.450 32.400 ;
        RECT 709.950 25.950 712.050 31.050 ;
        RECT 715.950 28.950 721.050 31.050 ;
        RECT 740.400 25.050 741.450 43.950 ;
        RECT 743.400 37.050 744.450 67.950 ;
        RECT 746.400 46.200 747.450 76.950 ;
        RECT 748.950 70.950 751.050 73.050 ;
        RECT 749.400 55.050 750.450 70.950 ;
        RECT 758.400 64.050 759.450 130.950 ;
        RECT 766.950 130.800 769.050 132.900 ;
        RECT 778.950 130.950 781.050 136.050 ;
        RECT 790.950 130.950 793.050 136.050 ;
        RECT 797.400 133.050 798.450 145.950 ;
        RECT 799.950 139.950 802.050 142.050 ;
        RECT 796.950 130.950 799.050 133.050 ;
        RECT 767.400 118.050 768.450 130.800 ;
        RECT 784.950 127.950 790.050 130.050 ;
        RECT 775.950 118.950 778.050 121.050 ;
        RECT 766.950 115.950 769.050 118.050 ;
        RECT 766.950 110.400 769.050 112.500 ;
        RECT 762.000 105.450 766.050 106.050 ;
        RECT 761.400 103.950 766.050 105.450 ;
        RECT 751.950 58.950 754.050 64.050 ;
        RECT 757.950 61.950 760.050 64.050 ;
        RECT 748.950 52.950 751.050 55.050 ;
        RECT 754.950 52.950 757.050 58.050 ;
        RECT 761.400 55.050 762.450 103.950 ;
        RECT 767.850 95.400 769.050 110.400 ;
        RECT 776.400 106.050 777.450 118.950 ;
        RECT 787.950 110.400 790.050 112.500 ;
        RECT 781.950 106.950 784.050 109.050 ;
        RECT 775.950 100.950 778.050 106.050 ;
        RECT 782.400 103.050 783.450 106.950 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 766.950 93.300 769.050 95.400 ;
        RECT 767.850 89.700 769.050 93.300 ;
        RECT 788.100 90.600 789.300 110.400 ;
        RECT 800.400 106.050 801.450 139.950 ;
        RECT 802.950 130.950 805.050 133.050 ;
        RECT 803.400 127.050 804.450 130.950 ;
        RECT 802.950 124.950 805.050 127.050 ;
        RECT 800.400 103.950 805.050 106.050 ;
        RECT 793.950 100.950 796.050 103.050 ;
        RECT 766.950 87.600 769.050 89.700 ;
        RECT 787.950 88.500 790.050 90.600 ;
        RECT 781.950 64.950 784.050 67.050 ;
        RECT 763.950 58.950 769.050 61.050 ;
        RECT 772.950 58.950 775.050 61.050 ;
        RECT 775.950 58.950 781.050 61.050 ;
        RECT 760.950 52.950 763.050 55.050 ;
        RECT 769.950 49.950 772.050 52.050 ;
        RECT 745.950 44.100 748.050 46.200 ;
        RECT 745.950 40.800 748.050 42.900 ;
        RECT 742.950 34.950 745.050 37.050 ;
        RECT 746.400 25.050 747.450 40.800 ;
        RECT 754.950 32.400 757.050 34.500 ;
        RECT 721.950 22.950 727.050 25.050 ;
        RECT 739.950 22.950 742.050 25.050 ;
        RECT 694.950 19.950 697.050 22.050 ;
        RECT 700.950 19.950 703.050 22.050 ;
        RECT 706.950 19.950 709.050 22.050 ;
        RECT 730.950 19.950 733.050 22.050 ;
        RECT 745.950 19.950 748.050 25.050 ;
        RECT 751.950 22.950 754.050 28.050 ;
        RECT 701.400 13.050 702.450 19.950 ;
        RECT 731.400 16.050 732.450 19.950 ;
        RECT 736.950 16.950 739.050 19.050 ;
        RECT 755.850 17.400 757.050 32.400 ;
        RECT 763.950 22.950 766.050 28.050 ;
        RECT 770.400 25.050 771.450 49.950 ;
        RECT 773.400 46.050 774.450 58.950 ;
        RECT 782.400 55.050 783.450 64.950 ;
        RECT 787.950 58.950 793.050 61.050 ;
        RECT 775.950 49.950 778.050 55.050 ;
        RECT 781.950 52.950 784.050 55.050 ;
        RECT 787.950 52.950 790.050 55.050 ;
        RECT 772.950 43.950 775.050 46.050 ;
        RECT 788.400 43.050 789.450 52.950 ;
        RECT 787.950 40.950 790.050 43.050 ;
        RECT 781.950 34.950 784.050 37.050 ;
        RECT 787.950 34.950 790.050 37.050 ;
        RECT 775.950 32.400 778.050 34.500 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 730.950 13.950 733.050 16.050 ;
        RECT 737.400 13.050 738.450 16.950 ;
        RECT 742.950 13.950 748.050 16.050 ;
        RECT 754.950 15.300 757.050 17.400 ;
        RECT 664.950 9.600 667.050 11.700 ;
        RECT 685.950 10.500 688.050 12.600 ;
        RECT 700.950 10.950 703.050 13.050 ;
        RECT 736.950 10.950 739.050 13.050 ;
        RECT 755.850 11.700 757.050 15.300 ;
        RECT 776.100 12.600 777.300 32.400 ;
        RECT 778.950 28.950 781.050 31.050 ;
        RECT 779.400 16.050 780.450 28.950 ;
        RECT 778.950 13.950 781.050 16.050 ;
        RECT 782.400 13.050 783.450 34.950 ;
        RECT 788.400 28.050 789.450 34.950 ;
        RECT 787.950 25.950 790.050 28.050 ;
        RECT 794.400 25.050 795.450 100.950 ;
        RECT 796.950 73.950 799.050 76.050 ;
        RECT 793.950 22.950 796.050 25.050 ;
        RECT 797.400 19.050 798.450 73.950 ;
        RECT 800.400 67.050 801.450 103.950 ;
        RECT 806.400 103.200 807.450 166.950 ;
        RECT 809.400 121.050 810.450 178.950 ;
        RECT 812.400 154.050 813.450 178.950 ;
        RECT 817.950 173.400 819.150 188.400 ;
        RECT 820.950 178.950 823.050 184.050 ;
        RECT 817.950 171.300 820.050 173.400 ;
        RECT 817.950 167.700 819.150 171.300 ;
        RECT 817.950 165.600 820.050 167.700 ;
        RECT 811.950 151.950 814.050 154.050 ;
        RECT 820.950 151.950 823.050 154.050 ;
        RECT 821.400 142.050 822.450 151.950 ;
        RECT 811.950 139.950 817.050 142.050 ;
        RECT 820.950 139.950 823.050 142.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 808.950 118.950 811.050 121.050 ;
        RECT 808.950 103.950 811.050 109.050 ;
        RECT 805.950 101.100 808.050 103.200 ;
        RECT 812.400 100.050 813.450 133.950 ;
        RECT 817.950 130.950 820.050 133.050 ;
        RECT 805.950 97.800 808.050 99.900 ;
        RECT 811.950 97.950 814.050 100.050 ;
        RECT 806.400 73.050 807.450 97.800 ;
        RECT 808.950 82.950 811.050 85.050 ;
        RECT 805.950 70.950 808.050 73.050 ;
        RECT 799.950 64.950 802.050 67.050 ;
        RECT 806.400 61.050 807.450 70.950 ;
        RECT 805.950 58.950 808.050 61.050 ;
        RECT 802.950 52.950 805.050 55.050 ;
        RECT 803.400 31.050 804.450 52.950 ;
        RECT 809.400 37.050 810.450 82.950 ;
        RECT 818.400 79.050 819.450 130.950 ;
        RECT 817.950 76.950 820.050 79.050 ;
        RECT 814.950 64.950 817.050 67.050 ;
        RECT 815.400 58.050 816.450 64.950 ;
        RECT 814.950 55.950 817.050 58.050 ;
        RECT 808.950 34.950 811.050 37.050 ;
        RECT 802.950 28.950 805.050 31.050 ;
        RECT 827.400 25.050 828.450 391.950 ;
        RECT 811.950 22.950 814.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 812.400 19.050 813.450 22.950 ;
        RECT 796.950 16.950 799.050 19.050 ;
        RECT 802.950 16.950 808.050 19.050 ;
        RECT 811.950 16.950 814.050 19.050 ;
        RECT 754.950 9.600 757.050 11.700 ;
        RECT 775.950 10.500 778.050 12.600 ;
        RECT 781.950 10.950 784.050 13.050 ;
        RECT 367.950 4.950 370.050 7.050 ;
        RECT 478.950 4.950 481.050 7.050 ;
      LAYER metal3 ;
        RECT 331.950 819.600 334.050 820.050 ;
        RECT 382.950 819.600 385.050 820.050 ;
        RECT 331.950 818.400 385.050 819.600 ;
        RECT 331.950 817.950 334.050 818.400 ;
        RECT 382.950 817.950 385.050 818.400 ;
        RECT 388.950 819.600 391.050 820.050 ;
        RECT 433.950 819.600 436.050 820.050 ;
        RECT 388.950 818.400 436.050 819.600 ;
        RECT 388.950 817.950 391.050 818.400 ;
        RECT 433.950 817.950 436.050 818.400 ;
        RECT 472.950 819.600 475.050 820.050 ;
        RECT 514.950 819.600 517.050 820.050 ;
        RECT 472.950 818.400 517.050 819.600 ;
        RECT 472.950 817.950 475.050 818.400 ;
        RECT 514.950 817.950 517.050 818.400 ;
        RECT 520.950 819.600 523.050 820.050 ;
        RECT 520.950 818.400 651.600 819.600 ;
        RECT 520.950 817.950 523.050 818.400 ;
        RECT 58.950 816.600 61.050 817.050 ;
        RECT 160.950 816.600 163.050 817.050 ;
        RECT 58.950 815.400 163.050 816.600 ;
        RECT 58.950 814.950 61.050 815.400 ;
        RECT 160.950 814.950 163.050 815.400 ;
        RECT 385.950 816.600 388.050 817.050 ;
        RECT 415.950 816.600 418.050 817.050 ;
        RECT 517.950 816.600 520.050 817.050 ;
        RECT 385.950 815.400 520.050 816.600 ;
        RECT 650.400 816.600 651.600 818.400 ;
        RECT 745.950 816.600 748.050 817.050 ;
        RECT 650.400 815.400 748.050 816.600 ;
        RECT 385.950 814.950 388.050 815.400 ;
        RECT 415.950 814.950 418.050 815.400 ;
        RECT 517.950 814.950 520.050 815.400 ;
        RECT 745.950 814.950 748.050 815.400 ;
        RECT 13.950 813.600 16.050 814.050 ;
        RECT 37.950 813.600 40.050 814.050 ;
        RECT 13.950 812.400 40.050 813.600 ;
        RECT 13.950 811.950 16.050 812.400 ;
        RECT 37.950 811.950 40.050 812.400 ;
        RECT 535.950 813.600 538.050 814.050 ;
        RECT 550.950 813.600 553.050 814.050 ;
        RECT 586.950 813.600 589.050 814.050 ;
        RECT 535.950 812.400 589.050 813.600 ;
        RECT 535.950 811.950 538.050 812.400 ;
        RECT 550.950 811.950 553.050 812.400 ;
        RECT 586.950 811.950 589.050 812.400 ;
        RECT 703.950 813.600 706.050 814.050 ;
        RECT 718.800 813.600 720.900 814.050 ;
        RECT 703.950 812.400 720.900 813.600 ;
        RECT 703.950 811.950 706.050 812.400 ;
        RECT 718.800 811.950 720.900 812.400 ;
        RECT 722.100 813.600 724.200 814.050 ;
        RECT 739.950 813.600 742.050 814.050 ;
        RECT 722.100 812.400 742.050 813.600 ;
        RECT 722.100 811.950 724.200 812.400 ;
        RECT 739.950 811.950 742.050 812.400 ;
        RECT 814.950 813.600 817.050 814.050 ;
        RECT 823.950 813.600 826.050 814.050 ;
        RECT 814.950 812.400 826.050 813.600 ;
        RECT 814.950 811.950 817.050 812.400 ;
        RECT 823.950 811.950 826.050 812.400 ;
        RECT 307.950 810.600 310.050 811.050 ;
        RECT 319.950 810.600 322.050 811.050 ;
        RECT 307.950 809.400 322.050 810.600 ;
        RECT 307.950 808.950 310.050 809.400 ;
        RECT 319.950 808.950 322.050 809.400 ;
        RECT 427.950 810.600 430.050 811.050 ;
        RECT 463.950 810.600 466.050 811.050 ;
        RECT 484.950 810.600 487.050 811.050 ;
        RECT 427.950 809.400 487.050 810.600 ;
        RECT 427.950 808.950 430.050 809.400 ;
        RECT 463.950 808.950 466.050 809.400 ;
        RECT 484.950 808.950 487.050 809.400 ;
        RECT 502.950 810.600 505.050 811.050 ;
        RECT 511.950 810.600 514.050 811.050 ;
        RECT 622.950 810.600 625.050 811.050 ;
        RECT 502.950 809.400 625.050 810.600 ;
        RECT 502.950 808.950 505.050 809.400 ;
        RECT 511.950 808.950 514.050 809.400 ;
        RECT 622.950 808.950 625.050 809.400 ;
        RECT 787.950 810.600 790.050 811.050 ;
        RECT 802.950 810.600 805.050 811.050 ;
        RECT 811.950 810.600 814.050 811.050 ;
        RECT 787.950 809.400 814.050 810.600 ;
        RECT 787.950 808.950 790.050 809.400 ;
        RECT 802.950 808.950 805.050 809.400 ;
        RECT 811.950 808.950 814.050 809.400 ;
        RECT 16.950 807.600 19.050 808.050 ;
        RECT 28.950 807.600 31.050 808.050 ;
        RECT 112.950 807.600 115.050 808.050 ;
        RECT 16.950 806.400 115.050 807.600 ;
        RECT 16.950 805.950 19.050 806.400 ;
        RECT 28.950 805.950 31.050 806.400 ;
        RECT 112.950 805.950 115.050 806.400 ;
        RECT 244.950 807.600 247.050 808.050 ;
        RECT 259.950 807.600 262.050 808.050 ;
        RECT 244.950 806.400 262.050 807.600 ;
        RECT 244.950 805.950 247.050 806.400 ;
        RECT 259.950 805.950 262.050 806.400 ;
        RECT 316.950 807.600 319.050 808.200 ;
        RECT 331.950 807.600 334.050 808.050 ;
        RECT 316.950 806.400 334.050 807.600 ;
        RECT 316.950 806.100 319.050 806.400 ;
        RECT 331.950 805.950 334.050 806.400 ;
        RECT 352.950 807.600 355.050 808.200 ;
        RECT 364.950 807.600 367.050 808.050 ;
        RECT 379.950 807.600 382.050 808.050 ;
        RECT 418.950 807.600 421.050 808.050 ;
        RECT 352.950 806.400 421.050 807.600 ;
        RECT 352.950 806.100 355.050 806.400 ;
        RECT 364.950 805.950 367.050 806.400 ;
        RECT 379.950 805.950 382.050 806.400 ;
        RECT 418.950 805.950 421.050 806.400 ;
        RECT 601.950 807.600 604.050 808.050 ;
        RECT 613.950 807.600 616.050 808.050 ;
        RECT 601.950 806.400 616.050 807.600 ;
        RECT 601.950 805.950 604.050 806.400 ;
        RECT 613.950 805.950 616.050 806.400 ;
        RECT 652.950 807.600 655.050 808.050 ;
        RECT 685.950 807.600 688.050 808.050 ;
        RECT 652.950 806.400 688.050 807.600 ;
        RECT 652.950 805.950 655.050 806.400 ;
        RECT 685.950 805.950 688.050 806.400 ;
        RECT 709.950 807.600 712.050 808.050 ;
        RECT 730.950 807.600 733.050 808.050 ;
        RECT 709.950 806.400 733.050 807.600 ;
        RECT 709.950 805.950 712.050 806.400 ;
        RECT 730.950 805.950 733.050 806.400 ;
        RECT 739.950 807.600 742.050 808.050 ;
        RECT 760.950 807.600 763.050 808.050 ;
        RECT 739.950 806.400 763.050 807.600 ;
        RECT 739.950 805.950 742.050 806.400 ;
        RECT 760.950 805.950 763.050 806.400 ;
        RECT 88.950 804.600 91.050 805.050 ;
        RECT 115.950 804.600 118.050 805.050 ;
        RECT 121.950 804.600 124.050 805.050 ;
        RECT 88.950 803.400 111.600 804.600 ;
        RECT 88.950 802.950 91.050 803.400 ;
        RECT 13.950 801.600 16.050 802.050 ;
        RECT 34.950 801.600 37.050 802.050 ;
        RECT 43.950 801.600 46.050 802.050 ;
        RECT 55.950 801.600 58.050 802.050 ;
        RECT 13.950 800.400 58.050 801.600 ;
        RECT 13.950 799.950 16.050 800.400 ;
        RECT 34.950 799.950 37.050 800.400 ;
        RECT 43.950 799.950 46.050 800.400 ;
        RECT 55.950 799.950 58.050 800.400 ;
        RECT 76.950 801.600 79.050 802.050 ;
        RECT 100.950 801.600 103.050 802.050 ;
        RECT 76.950 800.400 103.050 801.600 ;
        RECT 76.950 799.950 79.050 800.400 ;
        RECT 100.950 799.950 103.050 800.400 ;
        RECT 61.950 798.600 64.050 799.050 ;
        RECT 94.950 798.600 97.050 799.050 ;
        RECT 61.950 797.400 97.050 798.600 ;
        RECT 110.400 798.600 111.600 803.400 ;
        RECT 115.950 803.400 124.050 804.600 ;
        RECT 115.950 802.950 118.050 803.400 ;
        RECT 121.950 802.950 124.050 803.400 ;
        RECT 133.950 801.600 136.050 805.050 ;
        RECT 166.950 804.600 169.050 805.050 ;
        RECT 187.950 804.600 190.050 805.050 ;
        RECT 166.950 803.400 190.050 804.600 ;
        RECT 166.950 802.950 169.050 803.400 ;
        RECT 187.950 802.950 190.050 803.400 ;
        RECT 316.950 804.600 319.050 804.900 ;
        RECT 322.950 804.600 325.050 805.200 ;
        RECT 316.950 803.400 325.050 804.600 ;
        RECT 316.950 802.800 319.050 803.400 ;
        RECT 322.950 803.100 325.050 803.400 ;
        RECT 139.950 801.600 142.050 802.050 ;
        RECT 151.950 801.600 154.050 802.050 ;
        RECT 193.950 801.600 196.050 802.200 ;
        RECT 133.950 801.000 142.050 801.600 ;
        RECT 134.400 800.400 142.050 801.000 ;
        RECT 139.950 799.950 142.050 800.400 ;
        RECT 146.400 800.400 154.050 801.600 ;
        RECT 146.400 798.600 147.600 800.400 ;
        RECT 151.950 799.950 154.050 800.400 ;
        RECT 164.400 800.400 196.050 801.600 ;
        RECT 164.400 799.050 165.600 800.400 ;
        RECT 193.950 800.100 196.050 800.400 ;
        RECT 214.950 801.600 217.050 802.050 ;
        RECT 226.950 801.600 229.050 802.050 ;
        RECT 247.950 801.600 250.050 802.050 ;
        RECT 214.950 800.400 250.050 801.600 ;
        RECT 214.950 799.950 217.050 800.400 ;
        RECT 226.950 799.950 229.050 800.400 ;
        RECT 247.950 799.950 250.050 800.400 ;
        RECT 262.950 801.600 265.050 802.050 ;
        RECT 271.950 801.600 274.050 802.050 ;
        RECT 286.950 801.600 289.050 802.050 ;
        RECT 262.950 800.400 289.050 801.600 ;
        RECT 352.950 801.600 355.050 804.900 ;
        RECT 388.950 804.600 391.050 805.050 ;
        RECT 409.950 804.600 412.050 805.050 ;
        RECT 388.950 803.400 412.050 804.600 ;
        RECT 388.950 802.950 391.050 803.400 ;
        RECT 409.950 802.950 412.050 803.400 ;
        RECT 448.950 804.600 451.050 805.050 ;
        RECT 478.950 804.600 481.050 805.050 ;
        RECT 541.950 804.600 544.050 805.050 ;
        RECT 448.950 803.400 544.050 804.600 ;
        RECT 448.950 802.950 451.050 803.400 ;
        RECT 478.950 802.950 481.050 803.400 ;
        RECT 541.950 802.950 544.050 803.400 ;
        RECT 577.950 804.600 580.050 805.050 ;
        RECT 643.950 804.600 646.050 805.050 ;
        RECT 577.950 803.400 646.050 804.600 ;
        RECT 577.950 802.950 580.050 803.400 ;
        RECT 643.950 802.950 646.050 803.400 ;
        RECT 745.950 804.600 748.050 805.050 ;
        RECT 784.950 804.600 787.050 808.050 ;
        RECT 799.950 804.600 802.050 805.050 ;
        RECT 745.950 804.000 787.050 804.600 ;
        RECT 745.950 803.400 786.600 804.000 ;
        RECT 788.400 803.400 802.050 804.600 ;
        RECT 745.950 802.950 748.050 803.400 ;
        RECT 364.950 801.600 367.050 801.900 ;
        RECT 373.950 801.600 376.050 802.050 ;
        RECT 352.950 801.000 376.050 801.600 ;
        RECT 353.400 800.400 376.050 801.000 ;
        RECT 262.950 799.950 265.050 800.400 ;
        RECT 271.950 799.950 274.050 800.400 ;
        RECT 286.950 799.950 289.050 800.400 ;
        RECT 364.950 799.800 367.050 800.400 ;
        RECT 373.950 799.950 376.050 800.400 ;
        RECT 469.950 799.950 475.050 802.050 ;
        RECT 499.950 801.600 502.050 802.050 ;
        RECT 511.950 801.600 514.050 802.050 ;
        RECT 499.950 800.400 514.050 801.600 ;
        RECT 499.950 799.950 502.050 800.400 ;
        RECT 511.950 799.950 514.050 800.400 ;
        RECT 565.950 801.600 568.050 802.050 ;
        RECT 571.950 801.600 574.050 802.050 ;
        RECT 565.950 800.400 574.050 801.600 ;
        RECT 565.950 799.950 568.050 800.400 ;
        RECT 571.950 799.950 574.050 800.400 ;
        RECT 679.950 801.600 682.050 802.200 ;
        RECT 709.950 801.600 712.050 802.050 ;
        RECT 679.950 800.400 712.050 801.600 ;
        RECT 679.950 800.100 682.050 800.400 ;
        RECT 709.950 799.950 712.050 800.400 ;
        RECT 736.950 801.600 739.050 802.050 ;
        RECT 757.950 801.600 760.050 802.050 ;
        RECT 788.400 801.600 789.600 803.400 ;
        RECT 799.950 802.950 802.050 803.400 ;
        RECT 805.950 804.600 808.050 805.050 ;
        RECT 817.950 804.600 820.050 805.050 ;
        RECT 805.950 803.400 820.050 804.600 ;
        RECT 805.950 802.950 808.050 803.400 ;
        RECT 817.950 802.950 820.050 803.400 ;
        RECT 736.950 800.400 760.050 801.600 ;
        RECT 736.950 799.950 739.050 800.400 ;
        RECT 757.950 799.950 760.050 800.400 ;
        RECT 761.400 800.400 789.600 801.600 ;
        RECT 793.950 801.600 796.050 802.050 ;
        RECT 802.950 801.600 805.050 801.900 ;
        RECT 793.950 800.400 805.050 801.600 ;
        RECT 110.400 797.400 147.600 798.600 ;
        RECT 157.950 798.600 160.050 799.050 ;
        RECT 163.950 798.600 166.050 799.050 ;
        RECT 157.950 797.400 166.050 798.600 ;
        RECT 61.950 796.950 64.050 797.400 ;
        RECT 94.950 796.950 97.050 797.400 ;
        RECT 157.950 796.950 160.050 797.400 ;
        RECT 163.950 796.950 166.050 797.400 ;
        RECT 229.950 798.600 232.050 799.050 ;
        RECT 244.950 798.600 247.050 799.050 ;
        RECT 229.950 797.400 247.050 798.600 ;
        RECT 229.950 796.950 232.050 797.400 ;
        RECT 244.950 796.950 247.050 797.400 ;
        RECT 280.950 798.600 283.050 799.050 ;
        RECT 304.950 798.600 307.050 799.050 ;
        RECT 346.950 798.600 349.050 799.050 ;
        RECT 358.950 798.600 361.050 799.050 ;
        RECT 280.950 797.400 361.050 798.600 ;
        RECT 280.950 796.950 283.050 797.400 ;
        RECT 304.950 796.950 307.050 797.400 ;
        RECT 346.950 796.950 349.050 797.400 ;
        RECT 358.950 796.950 361.050 797.400 ;
        RECT 391.950 798.600 394.050 799.050 ;
        RECT 391.950 797.400 408.600 798.600 ;
        RECT 391.950 796.950 394.050 797.400 ;
        RECT 407.400 796.050 408.600 797.400 ;
        RECT 37.950 795.600 40.050 796.050 ;
        RECT 58.950 795.600 61.050 796.050 ;
        RECT 37.950 794.400 61.050 795.600 ;
        RECT 37.950 793.950 40.050 794.400 ;
        RECT 58.950 793.950 61.050 794.400 ;
        RECT 148.950 795.600 151.050 796.050 ;
        RECT 166.950 795.600 169.050 796.050 ;
        RECT 148.950 794.400 169.050 795.600 ;
        RECT 148.950 793.950 151.050 794.400 ;
        RECT 166.950 793.950 169.050 794.400 ;
        RECT 217.950 795.600 220.050 796.050 ;
        RECT 223.950 795.600 226.050 796.050 ;
        RECT 250.950 795.600 253.050 796.050 ;
        RECT 217.950 794.400 253.050 795.600 ;
        RECT 217.950 793.950 220.050 794.400 ;
        RECT 223.950 793.950 226.050 794.400 ;
        RECT 250.950 793.950 253.050 794.400 ;
        RECT 406.950 795.600 409.050 796.050 ;
        RECT 424.950 795.600 427.050 796.050 ;
        RECT 406.950 794.400 427.050 795.600 ;
        RECT 433.950 795.600 436.050 799.050 ;
        RECT 541.950 798.600 544.050 799.050 ;
        RECT 580.950 798.600 583.050 799.050 ;
        RECT 541.950 797.400 583.050 798.600 ;
        RECT 541.950 796.950 544.050 797.400 ;
        RECT 580.950 796.950 583.050 797.400 ;
        RECT 604.950 798.600 607.050 799.050 ;
        RECT 619.950 798.600 622.050 799.050 ;
        RECT 604.950 797.400 622.050 798.600 ;
        RECT 604.950 796.950 607.050 797.400 ;
        RECT 619.950 796.950 622.050 797.400 ;
        RECT 625.950 798.600 628.050 799.050 ;
        RECT 631.950 798.600 634.050 799.050 ;
        RECT 625.950 797.400 634.050 798.600 ;
        RECT 625.950 796.950 628.050 797.400 ;
        RECT 631.950 796.950 634.050 797.400 ;
        RECT 715.950 796.950 721.050 799.050 ;
        RECT 754.950 798.600 757.050 799.050 ;
        RECT 761.400 798.600 762.600 800.400 ;
        RECT 793.950 799.950 796.050 800.400 ;
        RECT 802.950 799.800 805.050 800.400 ;
        RECT 754.950 797.400 762.600 798.600 ;
        RECT 808.950 798.600 811.050 799.050 ;
        RECT 820.950 798.600 823.050 799.050 ;
        RECT 808.950 797.400 823.050 798.600 ;
        RECT 754.950 796.950 757.050 797.400 ;
        RECT 808.950 796.950 811.050 797.400 ;
        RECT 820.950 796.950 823.050 797.400 ;
        RECT 448.950 795.600 451.050 796.050 ;
        RECT 433.950 795.000 451.050 795.600 ;
        RECT 434.400 794.400 451.050 795.000 ;
        RECT 406.950 793.950 409.050 794.400 ;
        RECT 424.950 793.950 427.050 794.400 ;
        RECT 448.950 793.950 451.050 794.400 ;
        RECT 538.950 795.600 541.050 796.050 ;
        RECT 550.950 795.600 553.050 796.050 ;
        RECT 538.950 794.400 553.050 795.600 ;
        RECT 538.950 793.950 541.050 794.400 ;
        RECT 550.950 793.950 553.050 794.400 ;
        RECT 652.950 795.600 655.050 796.050 ;
        RECT 679.950 795.600 682.050 796.050 ;
        RECT 652.950 794.400 682.050 795.600 ;
        RECT 652.950 793.950 655.050 794.400 ;
        RECT 679.950 793.950 682.050 794.400 ;
        RECT 25.950 792.600 28.050 793.050 ;
        RECT 97.950 792.600 100.050 793.050 ;
        RECT 25.950 791.400 100.050 792.600 ;
        RECT 25.950 790.950 28.050 791.400 ;
        RECT 97.950 790.950 100.050 791.400 ;
        RECT 301.950 792.600 304.050 793.050 ;
        RECT 322.950 792.600 325.050 793.050 ;
        RECT 349.950 792.600 352.050 793.050 ;
        RECT 301.950 791.400 352.050 792.600 ;
        RECT 301.950 790.950 304.050 791.400 ;
        RECT 322.950 790.950 325.050 791.400 ;
        RECT 349.950 790.950 352.050 791.400 ;
        RECT 367.950 792.600 370.050 793.050 ;
        RECT 379.950 792.600 382.050 793.050 ;
        RECT 367.950 791.400 382.050 792.600 ;
        RECT 367.950 790.950 370.050 791.400 ;
        RECT 379.950 790.950 382.050 791.400 ;
        RECT 427.950 792.600 430.050 793.050 ;
        RECT 445.950 792.600 448.050 793.050 ;
        RECT 460.950 792.600 463.050 793.050 ;
        RECT 427.950 791.400 463.050 792.600 ;
        RECT 427.950 790.950 430.050 791.400 ;
        RECT 445.950 790.950 448.050 791.400 ;
        RECT 460.950 790.950 463.050 791.400 ;
        RECT 487.950 792.600 490.050 793.050 ;
        RECT 520.950 792.600 523.050 793.050 ;
        RECT 532.950 792.600 535.050 793.050 ;
        RECT 487.950 791.400 535.050 792.600 ;
        RECT 487.950 790.950 490.050 791.400 ;
        RECT 520.950 790.950 523.050 791.400 ;
        RECT 532.950 790.950 535.050 791.400 ;
        RECT 592.950 792.600 595.050 793.050 ;
        RECT 766.950 792.600 769.050 793.050 ;
        RECT 592.950 791.400 769.050 792.600 ;
        RECT 592.950 790.950 595.050 791.400 ;
        RECT 766.950 790.950 769.050 791.400 ;
        RECT 79.950 789.600 82.050 790.050 ;
        RECT 109.950 789.600 112.050 790.050 ;
        RECT 79.950 788.400 112.050 789.600 ;
        RECT 79.950 787.950 82.050 788.400 ;
        RECT 109.950 787.950 112.050 788.400 ;
        RECT 310.950 789.600 313.050 790.050 ;
        RECT 328.950 789.600 331.050 790.050 ;
        RECT 397.950 789.600 400.050 790.050 ;
        RECT 310.950 788.400 400.050 789.600 ;
        RECT 310.950 787.950 313.050 788.400 ;
        RECT 328.950 787.950 331.050 788.400 ;
        RECT 397.950 787.950 400.050 788.400 ;
        RECT 424.950 789.600 427.050 790.050 ;
        RECT 568.950 789.600 571.050 790.050 ;
        RECT 424.950 788.400 571.050 789.600 ;
        RECT 424.950 787.950 427.050 788.400 ;
        RECT 568.950 787.950 571.050 788.400 ;
        RECT 673.950 789.600 676.050 790.050 ;
        RECT 685.950 789.600 688.050 790.050 ;
        RECT 673.950 788.400 688.050 789.600 ;
        RECT 673.950 787.950 676.050 788.400 ;
        RECT 685.950 787.950 688.050 788.400 ;
        RECT 130.950 786.600 133.050 787.050 ;
        RECT 211.950 786.600 214.050 787.050 ;
        RECT 229.950 786.600 232.050 787.050 ;
        RECT 130.950 785.400 232.050 786.600 ;
        RECT 130.950 784.950 133.050 785.400 ;
        RECT 211.950 784.950 214.050 785.400 ;
        RECT 229.950 784.950 232.050 785.400 ;
        RECT 247.950 786.600 250.050 787.050 ;
        RECT 325.950 786.600 328.050 787.050 ;
        RECT 247.950 785.400 328.050 786.600 ;
        RECT 247.950 784.950 250.050 785.400 ;
        RECT 325.950 784.950 328.050 785.400 ;
        RECT 496.950 786.600 499.050 787.050 ;
        RECT 535.950 786.600 538.050 787.050 ;
        RECT 496.950 785.400 538.050 786.600 ;
        RECT 496.950 784.950 499.050 785.400 ;
        RECT 535.950 784.950 538.050 785.400 ;
        RECT 49.950 783.600 52.050 784.050 ;
        RECT 61.950 783.600 64.050 784.050 ;
        RECT 73.950 783.600 76.050 784.050 ;
        RECT 136.950 783.600 139.050 784.050 ;
        RECT 49.950 782.400 139.050 783.600 ;
        RECT 49.950 781.950 52.050 782.400 ;
        RECT 61.950 781.950 64.050 782.400 ;
        RECT 73.950 781.950 76.050 782.400 ;
        RECT 136.950 781.950 139.050 782.400 ;
        RECT 340.950 783.600 343.050 784.050 ;
        RECT 394.950 783.600 397.050 784.050 ;
        RECT 340.950 782.400 397.050 783.600 ;
        RECT 340.950 781.950 343.050 782.400 ;
        RECT 394.950 781.950 397.050 782.400 ;
        RECT 490.950 783.600 493.050 784.050 ;
        RECT 538.950 783.600 541.050 784.050 ;
        RECT 490.950 782.400 541.050 783.600 ;
        RECT 490.950 781.950 493.050 782.400 ;
        RECT 538.950 781.950 541.050 782.400 ;
        RECT 565.950 783.600 568.050 784.050 ;
        RECT 592.950 783.600 595.050 784.050 ;
        RECT 565.950 782.400 595.050 783.600 ;
        RECT 565.950 781.950 568.050 782.400 ;
        RECT 592.950 781.950 595.050 782.400 ;
        RECT 601.950 783.600 604.050 784.050 ;
        RECT 610.950 783.600 613.050 784.050 ;
        RECT 601.950 782.400 613.050 783.600 ;
        RECT 601.950 781.950 604.050 782.400 ;
        RECT 610.950 781.950 613.050 782.400 ;
        RECT 118.950 780.600 121.050 781.050 ;
        RECT 184.950 780.600 187.050 781.050 ;
        RECT 448.950 780.600 451.050 781.050 ;
        RECT 118.950 779.400 451.050 780.600 ;
        RECT 118.950 778.950 121.050 779.400 ;
        RECT 184.950 778.950 187.050 779.400 ;
        RECT 448.950 778.950 451.050 779.400 ;
        RECT 562.950 780.600 565.050 781.050 ;
        RECT 625.950 780.600 628.050 781.050 ;
        RECT 562.950 779.400 628.050 780.600 ;
        RECT 562.950 778.950 565.050 779.400 ;
        RECT 625.950 778.950 628.050 779.400 ;
        RECT 100.950 777.600 103.050 778.050 ;
        RECT 208.950 777.600 211.050 778.050 ;
        RECT 229.950 777.600 232.050 778.050 ;
        RECT 100.950 776.400 232.050 777.600 ;
        RECT 100.950 775.950 103.050 776.400 ;
        RECT 208.950 775.950 211.050 776.400 ;
        RECT 229.950 775.950 232.050 776.400 ;
        RECT 250.950 777.600 253.050 778.050 ;
        RECT 376.950 777.600 379.050 778.050 ;
        RECT 250.950 776.400 379.050 777.600 ;
        RECT 250.950 775.950 253.050 776.400 ;
        RECT 376.950 775.950 379.050 776.400 ;
        RECT 388.950 777.600 391.050 778.050 ;
        RECT 484.950 777.600 487.050 778.050 ;
        RECT 388.950 776.400 487.050 777.600 ;
        RECT 388.950 775.950 391.050 776.400 ;
        RECT 484.950 775.950 487.050 776.400 ;
        RECT 532.950 777.600 535.050 778.050 ;
        RECT 556.950 777.600 559.050 778.050 ;
        RECT 532.950 776.400 559.050 777.600 ;
        RECT 532.950 775.950 535.050 776.400 ;
        RECT 556.950 775.950 559.050 776.400 ;
        RECT 583.950 777.600 586.050 778.050 ;
        RECT 598.950 777.600 601.050 778.050 ;
        RECT 613.950 777.600 616.050 778.050 ;
        RECT 583.950 776.400 616.050 777.600 ;
        RECT 583.950 775.950 586.050 776.400 ;
        RECT 598.950 775.950 601.050 776.400 ;
        RECT 613.950 775.950 616.050 776.400 ;
        RECT 685.950 777.600 688.050 778.050 ;
        RECT 715.950 777.600 718.050 778.050 ;
        RECT 685.950 776.400 718.050 777.600 ;
        RECT 685.950 775.950 688.050 776.400 ;
        RECT 715.950 775.950 718.050 776.400 ;
        RECT 43.950 774.600 46.050 775.050 ;
        RECT 91.950 774.600 94.050 775.050 ;
        RECT 43.950 773.400 94.050 774.600 ;
        RECT 43.950 772.950 46.050 773.400 ;
        RECT 91.950 772.950 94.050 773.400 ;
        RECT 316.950 774.600 319.050 775.050 ;
        RECT 373.950 774.600 376.050 775.050 ;
        RECT 316.950 773.400 376.050 774.600 ;
        RECT 316.950 772.950 319.050 773.400 ;
        RECT 373.950 772.950 376.050 773.400 ;
        RECT 391.950 774.600 394.050 775.050 ;
        RECT 475.950 774.600 478.050 775.050 ;
        RECT 391.950 773.400 478.050 774.600 ;
        RECT 391.950 772.950 394.050 773.400 ;
        RECT 475.950 772.950 478.050 773.400 ;
        RECT 544.950 774.600 547.050 775.050 ;
        RECT 565.950 774.600 568.050 775.050 ;
        RECT 544.950 773.400 568.050 774.600 ;
        RECT 544.950 772.950 547.050 773.400 ;
        RECT 565.950 772.950 568.050 773.400 ;
        RECT 640.950 774.600 643.050 775.050 ;
        RECT 673.950 774.600 676.050 775.050 ;
        RECT 640.950 773.400 676.050 774.600 ;
        RECT 640.950 772.950 643.050 773.400 ;
        RECT 673.950 772.950 676.050 773.400 ;
        RECT 763.950 774.600 766.050 775.050 ;
        RECT 799.950 774.600 802.050 775.050 ;
        RECT 763.950 773.400 802.050 774.600 ;
        RECT 763.950 772.950 766.050 773.400 ;
        RECT 799.950 772.950 802.050 773.400 ;
        RECT 4.950 771.600 7.050 772.050 ;
        RECT 13.950 771.600 16.050 772.050 ;
        RECT 4.950 770.400 16.050 771.600 ;
        RECT 4.950 769.950 7.050 770.400 ;
        RECT 13.950 769.950 16.050 770.400 ;
        RECT 58.950 771.600 61.050 772.050 ;
        RECT 70.950 771.600 73.050 772.050 ;
        RECT 58.950 770.400 73.050 771.600 ;
        RECT 58.950 769.950 61.050 770.400 ;
        RECT 70.950 769.950 73.050 770.400 ;
        RECT 109.950 771.600 112.050 772.050 ;
        RECT 124.950 771.600 127.050 772.050 ;
        RECT 109.950 770.400 127.050 771.600 ;
        RECT 109.950 769.950 112.050 770.400 ;
        RECT 124.950 769.950 127.050 770.400 ;
        RECT 160.950 771.600 163.050 772.050 ;
        RECT 232.950 771.600 235.050 772.050 ;
        RECT 160.950 770.400 235.050 771.600 ;
        RECT 160.950 769.950 163.050 770.400 ;
        RECT 232.950 769.950 235.050 770.400 ;
        RECT 325.950 771.600 328.050 772.050 ;
        RECT 397.950 771.600 400.050 772.050 ;
        RECT 325.950 770.400 400.050 771.600 ;
        RECT 325.950 769.950 328.050 770.400 ;
        RECT 397.950 769.950 400.050 770.400 ;
        RECT 463.950 771.600 466.050 772.050 ;
        RECT 493.950 771.600 496.050 772.050 ;
        RECT 463.950 770.400 496.050 771.600 ;
        RECT 463.950 769.950 466.050 770.400 ;
        RECT 493.950 769.950 496.050 770.400 ;
        RECT 568.950 771.600 571.050 772.050 ;
        RECT 580.950 771.600 583.050 772.050 ;
        RECT 568.950 770.400 583.050 771.600 ;
        RECT 568.950 769.950 571.050 770.400 ;
        RECT 580.950 769.950 583.050 770.400 ;
        RECT 595.950 771.600 598.050 772.050 ;
        RECT 724.950 771.600 727.050 772.200 ;
        RECT 784.950 771.600 787.050 772.200 ;
        RECT 793.950 771.600 796.050 772.050 ;
        RECT 595.950 770.400 642.600 771.600 ;
        RECT 595.950 769.950 598.050 770.400 ;
        RECT 106.950 768.600 109.050 769.050 ;
        RECT 130.950 768.600 133.050 769.050 ;
        RECT 136.950 768.600 139.050 769.050 ;
        RECT 106.950 767.400 114.600 768.600 ;
        RECT 106.950 766.950 109.050 767.400 ;
        RECT 113.400 766.050 114.600 767.400 ;
        RECT 130.950 767.400 139.050 768.600 ;
        RECT 130.950 766.950 133.050 767.400 ;
        RECT 136.950 766.950 139.050 767.400 ;
        RECT 175.950 768.600 178.050 769.050 ;
        RECT 187.950 768.600 190.050 769.050 ;
        RECT 175.950 767.400 190.050 768.600 ;
        RECT 175.950 766.950 178.050 767.400 ;
        RECT 187.950 766.950 190.050 767.400 ;
        RECT 352.950 768.600 355.050 769.050 ;
        RECT 361.950 768.600 364.050 769.050 ;
        RECT 352.950 767.400 364.050 768.600 ;
        RECT 352.950 766.950 355.050 767.400 ;
        RECT 361.950 766.950 364.050 767.400 ;
        RECT 412.950 768.600 415.050 769.050 ;
        RECT 421.950 768.600 424.050 769.050 ;
        RECT 412.950 767.400 424.050 768.600 ;
        RECT 412.950 766.950 415.050 767.400 ;
        RECT 421.950 766.950 424.050 767.400 ;
        RECT 508.950 768.600 511.050 769.050 ;
        RECT 526.950 768.600 529.050 769.050 ;
        RECT 571.950 768.600 574.050 769.050 ;
        RECT 616.950 768.600 619.050 769.050 ;
        RECT 628.950 768.600 631.050 769.200 ;
        RECT 508.950 767.400 631.050 768.600 ;
        RECT 641.400 769.050 642.600 770.400 ;
        RECT 724.950 770.400 796.050 771.600 ;
        RECT 724.950 770.100 727.050 770.400 ;
        RECT 784.950 770.100 787.050 770.400 ;
        RECT 793.950 769.950 796.050 770.400 ;
        RECT 641.400 768.600 646.050 769.050 ;
        RECT 664.950 768.600 667.050 769.050 ;
        RECT 679.950 768.600 682.050 769.050 ;
        RECT 641.400 767.400 682.050 768.600 ;
        RECT 508.950 766.950 511.050 767.400 ;
        RECT 526.950 766.950 529.050 767.400 ;
        RECT 571.950 766.950 574.050 767.400 ;
        RECT 616.950 766.950 619.050 767.400 ;
        RECT 628.950 767.100 631.050 767.400 ;
        RECT 642.000 766.950 646.050 767.400 ;
        RECT 664.950 766.950 667.050 767.400 ;
        RECT 679.950 766.950 682.050 767.400 ;
        RECT 724.950 768.600 727.050 768.900 ;
        RECT 760.950 768.600 763.050 769.050 ;
        RECT 724.950 767.400 763.050 768.600 ;
        RECT 724.950 766.800 727.050 767.400 ;
        RECT 760.950 766.950 763.050 767.400 ;
        RECT 766.950 768.600 769.050 769.050 ;
        RECT 781.950 768.600 784.050 768.900 ;
        RECT 799.950 768.600 802.050 769.050 ;
        RECT 766.950 767.400 802.050 768.600 ;
        RECT 766.950 766.950 769.050 767.400 ;
        RECT 781.950 766.800 784.050 767.400 ;
        RECT 799.950 766.950 802.050 767.400 ;
        RECT 7.950 765.600 10.050 766.050 ;
        RECT 49.950 765.600 52.050 766.050 ;
        RECT 7.950 764.400 52.050 765.600 ;
        RECT 113.400 765.600 118.050 766.050 ;
        RECT 142.950 765.600 145.050 766.050 ;
        RECT 113.400 764.400 145.050 765.600 ;
        RECT 7.950 763.950 10.050 764.400 ;
        RECT 49.950 763.950 52.050 764.400 ;
        RECT 114.000 763.950 118.050 764.400 ;
        RECT 142.950 763.950 145.050 764.400 ;
        RECT 148.950 765.600 151.050 766.200 ;
        RECT 154.950 765.600 157.050 766.050 ;
        RECT 148.950 764.400 157.050 765.600 ;
        RECT 148.950 764.100 151.050 764.400 ;
        RECT 154.950 763.950 157.050 764.400 ;
        RECT 13.950 762.600 16.050 763.050 ;
        RECT 34.950 762.600 37.050 763.050 ;
        RECT 13.950 761.400 37.050 762.600 ;
        RECT 13.950 760.950 16.050 761.400 ;
        RECT 34.950 760.950 37.050 761.400 ;
        RECT 67.950 762.600 70.050 763.050 ;
        RECT 73.950 762.600 76.050 763.050 ;
        RECT 67.950 761.400 76.050 762.600 ;
        RECT 67.950 760.950 70.050 761.400 ;
        RECT 73.950 760.950 76.050 761.400 ;
        RECT 184.950 762.600 187.050 763.050 ;
        RECT 217.950 762.600 220.050 766.050 ;
        RECT 256.950 765.600 259.050 766.050 ;
        RECT 274.950 765.600 277.050 766.050 ;
        RECT 256.950 764.400 277.050 765.600 ;
        RECT 256.950 763.950 259.050 764.400 ;
        RECT 274.950 763.950 277.050 764.400 ;
        RECT 316.950 765.600 319.050 766.050 ;
        RECT 334.950 765.600 337.050 766.050 ;
        RECT 316.950 764.400 337.050 765.600 ;
        RECT 316.950 763.950 319.050 764.400 ;
        RECT 334.950 763.950 337.050 764.400 ;
        RECT 370.950 765.600 373.050 766.050 ;
        RECT 382.950 765.600 385.050 766.050 ;
        RECT 370.950 764.400 385.050 765.600 ;
        RECT 370.950 763.950 373.050 764.400 ;
        RECT 382.950 763.950 385.050 764.400 ;
        RECT 238.950 762.600 241.050 763.050 ;
        RECT 244.950 762.600 247.050 763.050 ;
        RECT 184.950 761.400 195.600 762.600 ;
        RECT 217.950 762.000 247.050 762.600 ;
        RECT 218.400 761.400 247.050 762.000 ;
        RECT 184.950 760.950 187.050 761.400 ;
        RECT 16.950 756.600 19.050 760.050 ;
        RECT 85.950 759.600 88.050 760.050 ;
        RECT 97.950 759.600 100.050 759.900 ;
        RECT 85.950 758.400 100.050 759.600 ;
        RECT 85.950 757.950 88.050 758.400 ;
        RECT 97.950 757.800 100.050 758.400 ;
        RECT 148.950 759.600 151.050 760.050 ;
        RECT 160.950 759.600 163.050 760.050 ;
        RECT 148.950 758.400 163.050 759.600 ;
        RECT 194.400 759.600 195.600 761.400 ;
        RECT 238.950 760.950 241.050 761.400 ;
        RECT 244.950 760.950 247.050 761.400 ;
        RECT 277.950 762.600 280.050 763.050 ;
        RECT 286.950 762.600 289.050 763.050 ;
        RECT 310.950 762.600 313.050 763.050 ;
        RECT 277.950 761.400 313.050 762.600 ;
        RECT 277.950 760.950 280.050 761.400 ;
        RECT 286.950 760.950 289.050 761.400 ;
        RECT 310.950 760.950 313.050 761.400 ;
        RECT 358.950 762.600 361.050 763.050 ;
        RECT 367.950 762.600 370.050 763.050 ;
        RECT 358.950 761.400 370.050 762.600 ;
        RECT 358.950 760.950 361.050 761.400 ;
        RECT 367.950 760.950 370.050 761.400 ;
        RECT 388.950 762.600 391.050 763.200 ;
        RECT 409.950 762.600 415.050 763.050 ;
        RECT 433.950 762.600 436.050 763.050 ;
        RECT 388.950 761.400 436.050 762.600 ;
        RECT 442.950 762.600 445.050 766.050 ;
        RECT 466.950 765.600 469.050 766.050 ;
        RECT 458.400 765.000 469.050 765.600 ;
        RECT 457.950 764.400 469.050 765.000 ;
        RECT 457.950 762.600 460.050 764.400 ;
        RECT 466.950 763.950 469.050 764.400 ;
        RECT 562.950 765.600 565.050 766.050 ;
        RECT 583.950 765.600 586.050 766.050 ;
        RECT 562.950 764.400 586.050 765.600 ;
        RECT 562.950 763.950 565.050 764.400 ;
        RECT 583.950 763.950 586.050 764.400 ;
        RECT 658.950 765.600 661.050 766.050 ;
        RECT 688.950 765.600 691.050 766.050 ;
        RECT 712.950 765.600 715.050 766.050 ;
        RECT 658.950 765.000 675.600 765.600 ;
        RECT 658.950 764.400 676.050 765.000 ;
        RECT 658.950 763.950 661.050 764.400 ;
        RECT 601.950 763.050 604.050 763.200 ;
        RECT 442.950 762.000 460.050 762.600 ;
        RECT 443.400 761.400 460.050 762.000 ;
        RECT 388.950 761.100 391.050 761.400 ;
        RECT 409.950 760.950 415.050 761.400 ;
        RECT 433.950 760.950 436.050 761.400 ;
        RECT 457.950 761.100 460.050 761.400 ;
        RECT 517.950 762.600 520.050 763.050 ;
        RECT 526.950 762.600 529.050 763.050 ;
        RECT 595.950 762.600 598.050 763.050 ;
        RECT 517.950 761.400 529.050 762.600 ;
        RECT 517.950 760.950 520.050 761.400 ;
        RECT 526.950 760.950 529.050 761.400 ;
        RECT 584.400 761.400 598.050 762.600 ;
        RECT 196.950 759.600 202.050 760.050 ;
        RECT 194.400 758.400 202.050 759.600 ;
        RECT 148.950 757.950 151.050 758.400 ;
        RECT 160.950 757.950 163.050 758.400 ;
        RECT 196.950 757.950 202.050 758.400 ;
        RECT 229.950 759.600 232.050 759.900 ;
        RECT 250.950 759.600 253.050 760.050 ;
        RECT 229.950 758.400 253.050 759.600 ;
        RECT 229.950 757.800 232.050 758.400 ;
        RECT 250.950 757.950 253.050 758.400 ;
        RECT 316.950 759.600 319.050 759.900 ;
        RECT 334.950 759.600 337.050 759.900 ;
        RECT 343.950 759.600 346.050 760.050 ;
        RECT 316.950 758.400 346.050 759.600 ;
        RECT 316.950 757.800 319.050 758.400 ;
        RECT 334.950 757.800 337.050 758.400 ;
        RECT 343.950 757.950 346.050 758.400 ;
        RECT 373.950 759.600 376.050 760.050 ;
        RECT 385.950 759.600 388.050 759.900 ;
        RECT 373.950 758.400 388.050 759.600 ;
        RECT 373.950 757.950 376.050 758.400 ;
        RECT 385.950 757.800 388.050 758.400 ;
        RECT 391.950 759.600 394.050 760.050 ;
        RECT 400.950 759.600 403.050 760.050 ;
        RECT 391.950 758.400 403.050 759.600 ;
        RECT 391.950 757.950 394.050 758.400 ;
        RECT 400.950 757.950 403.050 758.400 ;
        RECT 439.950 759.600 442.050 760.050 ;
        RECT 463.950 759.600 466.050 760.050 ;
        RECT 439.950 758.400 466.050 759.600 ;
        RECT 439.950 757.950 442.050 758.400 ;
        RECT 463.950 757.950 466.050 758.400 ;
        RECT 556.950 759.600 559.050 760.050 ;
        RECT 562.800 759.600 564.900 760.050 ;
        RECT 556.950 758.400 564.900 759.600 ;
        RECT 556.950 757.950 559.050 758.400 ;
        RECT 562.800 757.950 564.900 758.400 ;
        RECT 566.100 759.600 568.200 760.050 ;
        RECT 584.400 759.600 585.600 761.400 ;
        RECT 595.950 760.950 598.050 761.400 ;
        RECT 601.950 761.100 607.050 763.050 ;
        RECT 603.000 760.950 607.050 761.100 ;
        RECT 673.950 760.950 676.050 764.400 ;
        RECT 688.950 764.400 715.050 765.600 ;
        RECT 688.950 763.950 691.050 764.400 ;
        RECT 712.950 763.950 715.050 764.400 ;
        RECT 730.950 765.600 733.050 766.050 ;
        RECT 748.950 765.600 751.050 766.050 ;
        RECT 730.950 764.400 751.050 765.600 ;
        RECT 730.950 763.950 733.050 764.400 ;
        RECT 748.950 763.950 751.050 764.400 ;
        RECT 682.950 762.600 685.050 763.050 ;
        RECT 778.950 762.600 781.050 763.200 ;
        RECT 796.950 762.600 799.050 763.050 ;
        RECT 682.950 762.000 696.600 762.600 ;
        RECT 682.950 761.400 697.050 762.000 ;
        RECT 682.950 760.950 685.050 761.400 ;
        RECT 566.100 758.400 585.600 759.600 ;
        RECT 586.950 759.600 589.050 760.050 ;
        RECT 601.950 759.600 604.050 759.900 ;
        RECT 586.950 758.400 604.050 759.600 ;
        RECT 566.100 757.950 568.200 758.400 ;
        RECT 586.950 757.950 589.050 758.400 ;
        RECT 601.950 757.800 604.050 758.400 ;
        RECT 694.950 757.950 697.050 761.400 ;
        RECT 734.400 761.400 799.050 762.600 ;
        RECT 727.950 759.600 730.050 760.050 ;
        RECT 734.400 759.600 735.600 761.400 ;
        RECT 778.950 761.100 781.050 761.400 ;
        RECT 796.950 760.950 799.050 761.400 ;
        RECT 805.950 762.600 808.050 763.050 ;
        RECT 814.950 762.600 817.050 763.050 ;
        RECT 805.950 761.400 817.050 762.600 ;
        RECT 805.950 760.950 808.050 761.400 ;
        RECT 814.950 760.950 817.050 761.400 ;
        RECT 793.950 759.600 796.050 760.050 ;
        RECT 727.950 758.400 735.600 759.600 ;
        RECT 779.400 759.000 796.050 759.600 ;
        RECT 778.950 758.400 796.050 759.000 ;
        RECT 727.950 757.950 730.050 758.400 ;
        RECT 31.950 756.600 34.050 757.050 ;
        RECT 46.950 756.600 49.050 757.050 ;
        RECT 16.950 756.000 49.050 756.600 ;
        RECT 17.400 755.400 49.050 756.000 ;
        RECT 31.950 754.950 34.050 755.400 ;
        RECT 46.950 754.950 49.050 755.400 ;
        RECT 58.950 756.600 64.050 757.050 ;
        RECT 79.950 756.600 82.050 757.050 ;
        RECT 58.950 755.400 82.050 756.600 ;
        RECT 58.950 754.950 64.050 755.400 ;
        RECT 79.950 754.950 82.050 755.400 ;
        RECT 100.950 756.600 103.050 756.900 ;
        RECT 127.950 756.600 130.050 757.050 ;
        RECT 100.950 755.400 130.050 756.600 ;
        RECT 100.950 754.800 103.050 755.400 ;
        RECT 127.950 754.950 130.050 755.400 ;
        RECT 181.950 756.600 184.050 757.050 ;
        RECT 190.950 756.600 193.050 757.050 ;
        RECT 181.950 755.400 193.050 756.600 ;
        RECT 181.950 754.950 184.050 755.400 ;
        RECT 190.950 754.950 193.050 755.400 ;
        RECT 268.800 756.000 270.900 757.050 ;
        RECT 268.800 754.950 271.050 756.000 ;
        RECT 272.100 754.950 277.050 757.050 ;
        RECT 418.950 756.600 421.050 757.050 ;
        RECT 529.950 756.600 532.050 757.050 ;
        RECT 418.950 755.400 483.600 756.600 ;
        RECT 512.400 756.000 532.050 756.600 ;
        RECT 418.950 754.950 421.050 755.400 ;
        RECT 103.950 753.600 106.050 754.050 ;
        RECT 112.950 753.600 115.050 754.050 ;
        RECT 268.950 753.600 271.050 754.950 ;
        RECT 343.950 753.600 346.050 754.050 ;
        RECT 103.950 752.400 115.050 753.600 ;
        RECT 103.950 751.950 106.050 752.400 ;
        RECT 112.950 751.950 115.050 752.400 ;
        RECT 194.400 752.400 346.050 753.600 ;
        RECT 67.950 750.600 70.050 751.050 ;
        RECT 106.950 750.600 109.050 751.050 ;
        RECT 67.950 749.400 109.050 750.600 ;
        RECT 67.950 748.950 70.050 749.400 ;
        RECT 106.950 748.950 109.050 749.400 ;
        RECT 187.950 750.600 190.050 751.050 ;
        RECT 194.400 750.600 195.600 752.400 ;
        RECT 343.950 751.950 346.050 752.400 ;
        RECT 349.950 753.600 352.050 754.050 ;
        RECT 370.950 753.600 373.050 753.900 ;
        RECT 349.950 752.400 373.050 753.600 ;
        RECT 349.950 751.950 352.050 752.400 ;
        RECT 370.950 751.800 373.050 752.400 ;
        RECT 388.950 753.600 391.050 754.050 ;
        RECT 421.950 753.600 424.050 754.050 ;
        RECT 433.800 753.600 435.900 754.050 ;
        RECT 388.950 752.400 435.900 753.600 ;
        RECT 388.950 751.950 391.050 752.400 ;
        RECT 421.950 751.950 424.050 752.400 ;
        RECT 433.800 751.950 435.900 752.400 ;
        RECT 437.100 753.600 439.200 754.050 ;
        RECT 451.950 753.600 454.050 754.050 ;
        RECT 437.100 752.400 454.050 753.600 ;
        RECT 437.100 751.950 439.200 752.400 ;
        RECT 451.950 751.950 454.050 752.400 ;
        RECT 457.950 753.600 460.050 754.050 ;
        RECT 475.950 753.600 478.050 754.050 ;
        RECT 457.950 752.400 478.050 753.600 ;
        RECT 482.400 753.600 483.600 755.400 ;
        RECT 511.950 755.400 532.050 756.000 ;
        RECT 493.950 753.600 496.050 754.050 ;
        RECT 482.400 752.400 496.050 753.600 ;
        RECT 457.950 751.950 460.050 752.400 ;
        RECT 475.950 751.950 478.050 752.400 ;
        RECT 493.950 751.950 496.050 752.400 ;
        RECT 511.950 751.950 514.050 755.400 ;
        RECT 529.950 754.950 532.050 755.400 ;
        RECT 673.950 756.600 676.050 757.050 ;
        RECT 700.950 756.600 703.050 757.050 ;
        RECT 706.950 756.600 709.050 757.050 ;
        RECT 673.950 755.400 709.050 756.600 ;
        RECT 673.950 754.950 676.050 755.400 ;
        RECT 700.950 754.950 703.050 755.400 ;
        RECT 706.950 754.950 709.050 755.400 ;
        RECT 739.950 756.600 742.050 757.050 ;
        RECT 748.950 756.600 751.050 757.050 ;
        RECT 739.950 755.400 751.050 756.600 ;
        RECT 739.950 754.950 742.050 755.400 ;
        RECT 748.950 754.950 751.050 755.400 ;
        RECT 778.950 754.950 781.050 758.400 ;
        RECT 793.950 757.950 796.050 758.400 ;
        RECT 544.950 753.600 547.050 754.050 ;
        RECT 568.950 753.600 571.050 754.050 ;
        RECT 544.950 752.400 571.050 753.600 ;
        RECT 544.950 751.950 547.050 752.400 ;
        RECT 568.950 751.950 571.050 752.400 ;
        RECT 691.950 753.600 694.050 754.050 ;
        RECT 703.950 753.600 706.050 754.050 ;
        RECT 691.950 752.400 706.050 753.600 ;
        RECT 691.950 751.950 694.050 752.400 ;
        RECT 703.950 751.950 706.050 752.400 ;
        RECT 187.950 749.400 195.600 750.600 ;
        RECT 253.950 750.600 256.050 751.200 ;
        RECT 280.950 750.600 283.050 751.050 ;
        RECT 292.950 750.600 295.050 751.050 ;
        RECT 253.950 749.400 295.050 750.600 ;
        RECT 187.950 748.950 190.050 749.400 ;
        RECT 253.950 749.100 256.050 749.400 ;
        RECT 280.950 748.950 283.050 749.400 ;
        RECT 292.950 748.950 295.050 749.400 ;
        RECT 556.950 750.600 559.050 751.050 ;
        RECT 577.950 750.600 580.050 751.050 ;
        RECT 556.950 749.400 580.050 750.600 ;
        RECT 556.950 748.950 559.050 749.400 ;
        RECT 577.950 748.950 580.050 749.400 ;
        RECT 601.950 750.600 604.050 751.050 ;
        RECT 634.950 750.600 637.050 751.050 ;
        RECT 658.950 750.600 661.050 751.050 ;
        RECT 601.950 749.400 661.050 750.600 ;
        RECT 601.950 748.950 604.050 749.400 ;
        RECT 634.950 748.950 637.050 749.400 ;
        RECT 658.950 748.950 661.050 749.400 ;
        RECT 775.950 750.600 778.050 751.050 ;
        RECT 826.950 750.600 829.050 751.050 ;
        RECT 775.950 749.400 829.050 750.600 ;
        RECT 775.950 748.950 778.050 749.400 ;
        RECT 826.950 748.950 829.050 749.400 ;
        RECT 139.950 747.600 142.050 748.050 ;
        RECT 151.950 747.600 154.050 748.050 ;
        RECT 139.950 746.400 154.050 747.600 ;
        RECT 139.950 745.950 142.050 746.400 ;
        RECT 151.950 745.950 154.050 746.400 ;
        RECT 157.950 747.600 160.050 748.050 ;
        RECT 178.950 747.600 181.050 748.050 ;
        RECT 157.950 746.400 181.050 747.600 ;
        RECT 157.950 745.950 160.050 746.400 ;
        RECT 178.950 745.950 181.050 746.400 ;
        RECT 244.950 747.600 247.050 748.050 ;
        RECT 253.950 747.600 256.050 747.900 ;
        RECT 244.950 746.400 256.050 747.600 ;
        RECT 244.950 745.950 247.050 746.400 ;
        RECT 253.950 745.800 256.050 746.400 ;
        RECT 340.950 747.600 343.050 748.050 ;
        RECT 364.950 747.600 367.050 748.050 ;
        RECT 403.950 747.600 406.050 748.050 ;
        RECT 340.950 746.400 406.050 747.600 ;
        RECT 340.950 745.950 343.050 746.400 ;
        RECT 364.950 745.950 367.050 746.400 ;
        RECT 403.950 745.950 406.050 746.400 ;
        RECT 712.950 747.600 715.050 748.050 ;
        RECT 712.950 746.400 774.600 747.600 ;
        RECT 712.950 745.950 715.050 746.400 ;
        RECT 220.950 744.600 223.050 745.050 ;
        RECT 238.950 744.600 241.050 745.050 ;
        RECT 337.950 744.600 340.050 745.050 ;
        RECT 220.950 743.400 340.050 744.600 ;
        RECT 220.950 742.950 223.050 743.400 ;
        RECT 238.950 742.950 241.050 743.400 ;
        RECT 337.950 742.950 340.050 743.400 ;
        RECT 475.950 744.600 478.050 745.050 ;
        RECT 559.950 744.600 562.050 745.050 ;
        RECT 475.950 743.400 562.050 744.600 ;
        RECT 475.950 742.950 478.050 743.400 ;
        RECT 559.950 742.950 562.050 743.400 ;
        RECT 577.950 744.600 580.050 745.050 ;
        RECT 589.950 744.600 592.050 745.050 ;
        RECT 577.950 743.400 592.050 744.600 ;
        RECT 577.950 742.950 580.050 743.400 ;
        RECT 589.950 742.950 592.050 743.400 ;
        RECT 595.950 744.600 598.050 745.050 ;
        RECT 628.950 744.600 631.050 745.050 ;
        RECT 643.950 744.600 646.050 745.050 ;
        RECT 595.950 743.400 646.050 744.600 ;
        RECT 773.400 744.600 774.600 746.400 ;
        RECT 814.950 744.600 817.050 745.050 ;
        RECT 773.400 743.400 817.050 744.600 ;
        RECT 595.950 742.950 598.050 743.400 ;
        RECT 628.950 742.950 631.050 743.400 ;
        RECT 643.950 742.950 646.050 743.400 ;
        RECT 814.950 742.950 817.050 743.400 ;
        RECT 115.950 741.600 118.050 742.050 ;
        RECT 193.950 741.600 196.050 742.050 ;
        RECT 226.950 741.600 229.050 742.050 ;
        RECT 244.950 741.600 247.050 742.050 ;
        RECT 115.950 740.400 247.050 741.600 ;
        RECT 115.950 739.950 118.050 740.400 ;
        RECT 193.950 739.950 196.050 740.400 ;
        RECT 226.950 739.950 229.050 740.400 ;
        RECT 244.950 739.950 247.050 740.400 ;
        RECT 298.950 741.600 301.050 742.050 ;
        RECT 304.950 741.600 307.050 742.050 ;
        RECT 298.950 740.400 307.050 741.600 ;
        RECT 298.950 739.950 301.050 740.400 ;
        RECT 304.950 739.950 307.050 740.400 ;
        RECT 415.950 741.600 418.050 742.050 ;
        RECT 436.950 741.600 439.050 742.050 ;
        RECT 415.950 740.400 439.050 741.600 ;
        RECT 415.950 739.950 418.050 740.400 ;
        RECT 436.950 739.950 439.050 740.400 ;
        RECT 457.950 741.600 460.050 742.050 ;
        RECT 466.950 741.600 469.050 742.050 ;
        RECT 457.950 740.400 469.050 741.600 ;
        RECT 457.950 739.950 460.050 740.400 ;
        RECT 466.950 739.950 469.050 740.400 ;
        RECT 523.950 741.600 526.050 742.050 ;
        RECT 550.950 741.600 553.050 742.050 ;
        RECT 583.950 741.600 586.050 742.050 ;
        RECT 523.950 740.400 586.050 741.600 ;
        RECT 523.950 739.950 526.050 740.400 ;
        RECT 550.950 739.950 553.050 740.400 ;
        RECT 583.950 739.950 586.050 740.400 ;
        RECT 733.950 741.600 736.050 742.050 ;
        RECT 745.950 741.600 748.050 742.050 ;
        RECT 733.950 740.400 748.050 741.600 ;
        RECT 733.950 739.950 736.050 740.400 ;
        RECT 745.950 739.950 748.050 740.400 ;
        RECT 49.950 738.600 52.050 739.050 ;
        RECT 76.950 738.600 79.050 739.050 ;
        RECT 49.950 737.400 79.050 738.600 ;
        RECT 49.950 736.950 52.050 737.400 ;
        RECT 76.950 736.950 79.050 737.400 ;
        RECT 121.950 738.600 124.050 739.050 ;
        RECT 136.950 738.600 139.050 739.050 ;
        RECT 121.950 737.400 139.050 738.600 ;
        RECT 121.950 736.950 124.050 737.400 ;
        RECT 136.950 736.950 139.050 737.400 ;
        RECT 166.950 738.600 169.050 739.050 ;
        RECT 451.950 738.600 454.050 739.050 ;
        RECT 166.950 737.400 454.050 738.600 ;
        RECT 166.950 736.950 169.050 737.400 ;
        RECT 451.950 736.950 454.050 737.400 ;
        RECT 526.950 738.600 529.050 739.050 ;
        RECT 547.950 738.600 550.050 739.200 ;
        RECT 526.950 737.400 550.050 738.600 ;
        RECT 526.950 736.950 529.050 737.400 ;
        RECT 547.950 737.100 550.050 737.400 ;
        RECT 634.950 738.600 637.050 739.050 ;
        RECT 676.950 738.600 679.050 739.050 ;
        RECT 685.950 738.600 688.050 739.050 ;
        RECT 634.950 737.400 688.050 738.600 ;
        RECT 634.950 736.950 637.050 737.400 ;
        RECT 676.950 736.950 679.050 737.400 ;
        RECT 685.950 736.950 688.050 737.400 ;
        RECT 184.950 735.600 187.050 736.050 ;
        RECT 196.950 735.600 199.050 736.050 ;
        RECT 184.950 734.400 199.050 735.600 ;
        RECT 184.950 733.950 187.050 734.400 ;
        RECT 196.950 733.950 199.050 734.400 ;
        RECT 205.950 735.600 208.050 736.200 ;
        RECT 217.950 735.600 220.050 736.050 ;
        RECT 205.950 734.400 220.050 735.600 ;
        RECT 205.950 734.100 208.050 734.400 ;
        RECT 217.950 733.950 220.050 734.400 ;
        RECT 223.950 735.600 226.050 736.050 ;
        RECT 235.950 735.600 238.050 736.050 ;
        RECT 241.950 735.600 244.050 736.050 ;
        RECT 223.950 734.400 244.050 735.600 ;
        RECT 223.950 733.950 226.050 734.400 ;
        RECT 235.950 733.950 238.050 734.400 ;
        RECT 241.950 733.950 244.050 734.400 ;
        RECT 295.950 735.600 298.050 736.050 ;
        RECT 307.950 735.600 310.050 736.050 ;
        RECT 325.950 735.600 328.050 736.050 ;
        RECT 295.950 734.400 328.050 735.600 ;
        RECT 295.950 733.950 298.050 734.400 ;
        RECT 307.950 733.950 310.050 734.400 ;
        RECT 325.950 733.950 328.050 734.400 ;
        RECT 367.950 735.600 370.050 736.050 ;
        RECT 385.950 735.600 388.050 736.050 ;
        RECT 367.950 734.400 388.050 735.600 ;
        RECT 367.950 733.950 370.050 734.400 ;
        RECT 385.950 733.950 388.050 734.400 ;
        RECT 466.950 735.600 469.050 736.050 ;
        RECT 472.950 735.600 475.050 736.050 ;
        RECT 466.950 734.400 475.050 735.600 ;
        RECT 466.950 733.950 469.050 734.400 ;
        RECT 472.950 733.950 475.050 734.400 ;
        RECT 547.950 735.600 550.050 735.900 ;
        RECT 553.950 735.600 556.050 736.050 ;
        RECT 547.950 734.400 556.050 735.600 ;
        RECT 547.950 733.800 550.050 734.400 ;
        RECT 553.950 733.950 556.050 734.400 ;
        RECT 691.950 735.600 694.050 736.050 ;
        RECT 799.950 735.600 802.050 736.050 ;
        RECT 823.950 735.600 826.050 736.050 ;
        RECT 691.950 734.400 826.050 735.600 ;
        RECT 691.950 733.950 694.050 734.400 ;
        RECT 799.950 733.950 802.050 734.400 ;
        RECT 823.950 733.950 826.050 734.400 ;
        RECT 133.950 732.600 136.050 733.050 ;
        RECT 151.950 732.600 154.050 733.050 ;
        RECT 160.950 732.600 163.050 733.050 ;
        RECT 133.950 731.400 163.050 732.600 ;
        RECT 133.950 730.950 136.050 731.400 ;
        RECT 151.950 730.950 154.050 731.400 ;
        RECT 160.950 730.950 163.050 731.400 ;
        RECT 469.950 732.600 474.000 733.050 ;
        RECT 469.950 730.950 474.600 732.600 ;
        RECT 16.950 730.050 19.050 730.200 ;
        RECT 13.950 729.600 16.050 730.050 ;
        RECT 16.950 729.600 21.000 730.050 ;
        RECT 28.950 729.600 31.050 730.050 ;
        RECT 34.950 729.600 37.050 730.050 ;
        RECT 13.950 728.400 21.600 729.600 ;
        RECT 28.950 728.400 37.050 729.600 ;
        RECT 13.950 727.950 16.050 728.400 ;
        RECT 16.950 728.100 21.000 728.400 ;
        RECT 18.000 727.950 21.000 728.100 ;
        RECT 28.950 727.950 31.050 728.400 ;
        RECT 34.950 727.950 37.050 728.400 ;
        RECT 199.950 729.600 202.050 730.050 ;
        RECT 208.950 729.600 211.050 730.050 ;
        RECT 199.950 728.400 211.050 729.600 ;
        RECT 199.950 727.950 202.050 728.400 ;
        RECT 208.950 727.950 211.050 728.400 ;
        RECT 217.950 729.600 220.050 730.050 ;
        RECT 238.950 729.600 241.050 730.050 ;
        RECT 217.950 728.400 241.050 729.600 ;
        RECT 217.950 727.950 220.050 728.400 ;
        RECT 238.950 727.950 241.050 728.400 ;
        RECT 292.950 729.600 295.050 730.050 ;
        RECT 304.950 729.600 307.050 730.050 ;
        RECT 358.950 729.600 361.050 730.050 ;
        RECT 292.950 728.400 361.050 729.600 ;
        RECT 292.950 727.950 295.050 728.400 ;
        RECT 304.950 727.950 307.050 728.400 ;
        RECT 358.950 727.950 361.050 728.400 ;
        RECT 391.950 729.600 394.050 730.050 ;
        RECT 427.950 729.600 430.050 730.050 ;
        RECT 433.950 729.600 436.050 730.050 ;
        RECT 391.950 729.000 408.600 729.600 ;
        RECT 391.950 728.400 409.050 729.000 ;
        RECT 391.950 727.950 394.050 728.400 ;
        RECT 16.950 726.600 19.050 726.900 ;
        RECT 25.950 726.600 28.050 727.050 ;
        RECT 16.950 725.400 28.050 726.600 ;
        RECT 16.950 724.800 19.050 725.400 ;
        RECT 25.950 724.950 28.050 725.400 ;
        RECT 43.950 726.600 46.050 727.050 ;
        RECT 52.950 726.600 55.050 727.050 ;
        RECT 43.950 725.400 55.050 726.600 ;
        RECT 43.950 724.950 46.050 725.400 ;
        RECT 52.950 724.950 55.050 725.400 ;
        RECT 88.950 726.600 91.050 727.050 ;
        RECT 97.950 726.600 100.050 727.050 ;
        RECT 124.950 726.600 127.050 727.050 ;
        RECT 88.950 725.400 127.050 726.600 ;
        RECT 88.950 724.950 91.050 725.400 ;
        RECT 97.950 724.950 100.050 725.400 ;
        RECT 124.950 724.950 127.050 725.400 ;
        RECT 139.950 726.600 142.050 727.050 ;
        RECT 145.950 726.600 148.050 727.200 ;
        RECT 139.950 725.400 148.050 726.600 ;
        RECT 139.950 724.950 142.050 725.400 ;
        RECT 145.950 725.100 148.050 725.400 ;
        RECT 181.950 726.600 184.050 727.050 ;
        RECT 190.950 726.600 193.050 727.050 ;
        RECT 181.950 725.400 193.050 726.600 ;
        RECT 181.950 724.950 184.050 725.400 ;
        RECT 190.950 724.950 193.050 725.400 ;
        RECT 265.950 726.600 268.050 727.050 ;
        RECT 271.950 726.600 274.050 727.050 ;
        RECT 349.950 726.600 352.050 727.050 ;
        RECT 265.950 725.400 274.050 726.600 ;
        RECT 335.400 726.000 352.050 726.600 ;
        RECT 265.950 724.950 268.050 725.400 ;
        RECT 271.950 724.950 274.050 725.400 ;
        RECT 334.950 725.400 352.050 726.000 ;
        RECT 61.950 723.600 64.050 724.050 ;
        RECT 67.950 723.600 70.050 724.050 ;
        RECT 61.950 722.400 70.050 723.600 ;
        RECT 61.950 721.950 64.050 722.400 ;
        RECT 67.950 721.950 70.050 722.400 ;
        RECT 109.950 723.600 112.050 724.050 ;
        RECT 121.950 723.600 124.050 724.050 ;
        RECT 109.950 722.400 124.050 723.600 ;
        RECT 109.950 721.950 112.050 722.400 ;
        RECT 121.950 721.950 124.050 722.400 ;
        RECT 175.950 723.600 178.050 724.050 ;
        RECT 184.950 723.600 187.050 724.050 ;
        RECT 175.950 722.400 187.050 723.600 ;
        RECT 175.950 721.950 178.050 722.400 ;
        RECT 184.950 721.950 187.050 722.400 ;
        RECT 196.950 723.600 199.050 724.050 ;
        RECT 208.950 723.600 211.050 723.900 ;
        RECT 196.950 722.400 211.050 723.600 ;
        RECT 196.950 721.950 199.050 722.400 ;
        RECT 208.950 721.800 211.050 722.400 ;
        RECT 214.950 723.600 217.050 724.050 ;
        RECT 223.950 723.600 226.050 724.050 ;
        RECT 214.950 722.400 226.050 723.600 ;
        RECT 214.950 721.950 217.050 722.400 ;
        RECT 223.950 721.950 226.050 722.400 ;
        RECT 250.950 723.600 253.050 724.050 ;
        RECT 259.950 723.600 262.050 724.050 ;
        RECT 250.950 722.400 262.050 723.600 ;
        RECT 250.950 721.950 253.050 722.400 ;
        RECT 259.950 721.950 262.050 722.400 ;
        RECT 277.950 723.600 280.050 724.050 ;
        RECT 283.950 723.600 286.050 724.050 ;
        RECT 277.950 722.400 286.050 723.600 ;
        RECT 277.950 721.950 280.050 722.400 ;
        RECT 283.950 721.950 286.050 722.400 ;
        RECT 334.950 721.950 337.050 725.400 ;
        RECT 349.950 724.950 352.050 725.400 ;
        RECT 370.950 723.600 373.050 727.050 ;
        RECT 406.950 724.950 409.050 728.400 ;
        RECT 427.950 728.400 436.050 729.600 ;
        RECT 473.400 729.600 474.600 730.950 ;
        RECT 490.950 729.600 493.050 730.050 ;
        RECT 523.950 729.600 526.050 730.050 ;
        RECT 473.400 728.400 526.050 729.600 ;
        RECT 427.950 727.950 430.050 728.400 ;
        RECT 433.950 727.950 436.050 728.400 ;
        RECT 490.950 727.950 493.050 728.400 ;
        RECT 523.950 727.950 526.050 728.400 ;
        RECT 574.950 729.600 577.050 730.050 ;
        RECT 583.950 729.600 586.050 730.050 ;
        RECT 607.950 729.600 610.050 733.050 ;
        RECT 703.950 732.600 706.050 733.050 ;
        RECT 718.950 732.600 721.050 733.050 ;
        RECT 703.950 731.400 721.050 732.600 ;
        RECT 703.950 730.950 706.050 731.400 ;
        RECT 718.950 730.950 721.050 731.400 ;
        RECT 574.950 729.000 610.050 729.600 ;
        RECT 658.950 729.600 661.050 730.050 ;
        RECT 682.950 729.600 685.050 730.050 ;
        RECT 688.950 729.600 691.050 730.050 ;
        RECT 574.950 728.400 609.600 729.000 ;
        RECT 658.950 728.400 691.050 729.600 ;
        RECT 574.950 727.950 577.050 728.400 ;
        RECT 583.950 727.950 586.050 728.400 ;
        RECT 658.950 727.950 661.050 728.400 ;
        RECT 682.950 727.950 685.050 728.400 ;
        RECT 688.950 727.950 691.050 728.400 ;
        RECT 745.950 729.600 748.050 730.050 ;
        RECT 775.950 729.600 778.050 730.050 ;
        RECT 745.950 728.400 778.050 729.600 ;
        RECT 745.950 727.950 748.050 728.400 ;
        RECT 775.950 727.950 778.050 728.400 ;
        RECT 460.950 726.600 463.050 727.200 ;
        RECT 481.950 726.600 484.050 727.050 ;
        RECT 519.000 726.600 523.050 727.050 ;
        RECT 541.950 726.600 544.050 727.050 ;
        RECT 559.950 726.600 562.050 727.050 ;
        RECT 460.950 725.400 484.050 726.600 ;
        RECT 518.400 725.400 562.050 726.600 ;
        RECT 460.950 725.100 463.050 725.400 ;
        RECT 481.950 724.950 484.050 725.400 ;
        RECT 519.000 724.950 523.050 725.400 ;
        RECT 541.950 724.950 544.050 725.400 ;
        RECT 559.950 724.950 562.050 725.400 ;
        RECT 595.950 726.600 598.050 727.050 ;
        RECT 634.950 726.600 637.050 726.900 ;
        RECT 595.950 725.400 637.050 726.600 ;
        RECT 595.950 724.950 598.050 725.400 ;
        RECT 634.950 724.800 637.050 725.400 ;
        RECT 667.950 726.600 670.050 727.050 ;
        RECT 685.950 726.600 688.050 727.050 ;
        RECT 667.950 725.400 688.050 726.600 ;
        RECT 667.950 724.950 670.050 725.400 ;
        RECT 685.950 724.950 688.050 725.400 ;
        RECT 787.950 724.950 793.050 727.050 ;
        RECT 820.950 726.600 823.050 727.200 ;
        RECT 826.950 726.600 829.050 727.050 ;
        RECT 820.950 725.400 829.050 726.600 ;
        RECT 820.950 725.100 823.050 725.400 ;
        RECT 826.950 724.950 829.050 725.400 ;
        RECT 382.950 723.600 385.050 724.050 ;
        RECT 388.950 723.600 391.050 723.900 ;
        RECT 409.950 723.600 412.050 724.050 ;
        RECT 370.950 723.000 412.050 723.600 ;
        RECT 371.400 722.400 412.050 723.000 ;
        RECT 382.950 721.950 385.050 722.400 ;
        RECT 388.950 721.800 391.050 722.400 ;
        RECT 409.950 721.950 412.050 722.400 ;
        RECT 430.950 723.600 433.050 724.050 ;
        RECT 439.950 723.600 442.050 724.050 ;
        RECT 430.950 722.400 442.050 723.600 ;
        RECT 430.950 721.950 433.050 722.400 ;
        RECT 439.950 721.950 442.050 722.400 ;
        RECT 451.950 723.600 454.050 724.050 ;
        RECT 460.950 723.600 463.050 723.900 ;
        RECT 451.950 722.400 463.050 723.600 ;
        RECT 451.950 721.950 454.050 722.400 ;
        RECT 460.950 721.800 463.050 722.400 ;
        RECT 502.950 723.600 505.050 724.050 ;
        RECT 535.950 723.600 538.050 724.050 ;
        RECT 502.950 722.400 538.050 723.600 ;
        RECT 502.950 721.950 505.050 722.400 ;
        RECT 535.950 721.950 538.050 722.400 ;
        RECT 640.950 723.600 643.050 724.050 ;
        RECT 646.950 723.600 649.050 724.050 ;
        RECT 658.950 723.600 661.050 724.050 ;
        RECT 640.950 722.400 661.050 723.600 ;
        RECT 640.950 721.950 643.050 722.400 ;
        RECT 646.950 721.950 649.050 722.400 ;
        RECT 658.950 721.950 661.050 722.400 ;
        RECT 331.950 720.600 334.050 721.050 ;
        RECT 340.950 720.600 343.050 721.050 ;
        RECT 331.950 719.400 343.050 720.600 ;
        RECT 331.950 718.950 334.050 719.400 ;
        RECT 340.950 718.950 343.050 719.400 ;
        RECT 424.950 720.600 427.050 721.050 ;
        RECT 448.950 720.600 451.050 721.050 ;
        RECT 424.950 719.400 451.050 720.600 ;
        RECT 424.950 718.950 427.050 719.400 ;
        RECT 448.950 718.950 451.050 719.400 ;
        RECT 469.950 720.600 472.050 721.050 ;
        RECT 487.950 720.600 490.050 721.050 ;
        RECT 469.950 719.400 490.050 720.600 ;
        RECT 469.950 718.950 472.050 719.400 ;
        RECT 487.950 718.950 490.050 719.400 ;
        RECT 505.950 720.600 508.050 721.050 ;
        RECT 523.950 720.600 526.050 721.050 ;
        RECT 544.950 720.600 547.050 721.050 ;
        RECT 505.950 719.400 547.050 720.600 ;
        RECT 505.950 718.950 508.050 719.400 ;
        RECT 523.950 718.950 526.050 719.400 ;
        RECT 544.950 718.950 547.050 719.400 ;
        RECT 550.950 720.600 553.050 721.050 ;
        RECT 568.950 720.600 571.050 721.050 ;
        RECT 550.950 719.400 571.050 720.600 ;
        RECT 550.950 718.950 553.050 719.400 ;
        RECT 568.950 718.950 571.050 719.400 ;
        RECT 583.950 720.600 586.050 721.050 ;
        RECT 625.950 720.600 628.050 721.050 ;
        RECT 583.950 719.400 628.050 720.600 ;
        RECT 583.950 718.950 586.050 719.400 ;
        RECT 625.950 718.950 628.050 719.400 ;
        RECT 643.950 720.600 646.050 721.050 ;
        RECT 664.950 720.600 667.050 724.050 ;
        RECT 739.950 723.600 742.050 724.050 ;
        RECT 757.950 723.600 760.050 724.050 ;
        RECT 778.950 723.600 781.050 724.050 ;
        RECT 739.950 722.400 781.050 723.600 ;
        RECT 739.950 721.950 742.050 722.400 ;
        RECT 757.950 721.950 760.050 722.400 ;
        RECT 778.950 721.950 781.050 722.400 ;
        RECT 643.950 720.000 667.050 720.600 ;
        RECT 643.950 719.400 666.600 720.000 ;
        RECT 643.950 718.950 646.050 719.400 ;
        RECT 22.950 717.600 25.050 718.050 ;
        RECT 112.950 717.600 115.050 718.050 ;
        RECT 22.950 716.400 115.050 717.600 ;
        RECT 22.950 715.950 25.050 716.400 ;
        RECT 112.950 715.950 115.050 716.400 ;
        RECT 133.950 717.600 136.050 718.050 ;
        RECT 169.950 717.600 172.050 718.050 ;
        RECT 199.950 717.600 202.050 718.050 ;
        RECT 133.950 716.400 202.050 717.600 ;
        RECT 133.950 715.950 136.050 716.400 ;
        RECT 169.950 715.950 172.050 716.400 ;
        RECT 199.950 715.950 202.050 716.400 ;
        RECT 286.950 717.600 289.050 718.050 ;
        RECT 298.950 717.600 301.050 718.050 ;
        RECT 286.950 716.400 301.050 717.600 ;
        RECT 286.950 715.950 289.050 716.400 ;
        RECT 298.950 715.950 301.050 716.400 ;
        RECT 334.950 717.600 337.050 718.050 ;
        RECT 370.950 717.600 373.050 718.050 ;
        RECT 334.950 716.400 373.050 717.600 ;
        RECT 334.950 715.950 337.050 716.400 ;
        RECT 370.950 715.950 373.050 716.400 ;
        RECT 535.950 717.600 538.050 718.050 ;
        RECT 577.950 717.600 580.050 718.050 ;
        RECT 535.950 716.400 580.050 717.600 ;
        RECT 535.950 715.950 538.050 716.400 ;
        RECT 577.950 715.950 580.050 716.400 ;
        RECT 721.950 717.600 724.050 718.050 ;
        RECT 760.950 717.600 763.050 718.050 ;
        RECT 721.950 716.400 763.050 717.600 ;
        RECT 721.950 715.950 724.050 716.400 ;
        RECT 760.950 715.950 763.050 716.400 ;
        RECT 805.950 717.600 808.050 718.050 ;
        RECT 814.950 717.600 817.050 718.050 ;
        RECT 820.950 717.600 823.050 718.050 ;
        RECT 805.950 716.400 823.050 717.600 ;
        RECT 805.950 715.950 808.050 716.400 ;
        RECT 814.950 715.950 817.050 716.400 ;
        RECT 820.950 715.950 823.050 716.400 ;
        RECT 115.950 714.600 118.050 715.050 ;
        RECT 127.950 714.600 130.050 715.050 ;
        RECT 115.950 713.400 130.050 714.600 ;
        RECT 115.950 712.950 118.050 713.400 ;
        RECT 127.950 712.950 130.050 713.400 ;
        RECT 208.950 714.600 211.050 715.050 ;
        RECT 271.950 714.600 274.050 715.050 ;
        RECT 208.950 713.400 274.050 714.600 ;
        RECT 208.950 712.950 211.050 713.400 ;
        RECT 271.950 712.950 274.050 713.400 ;
        RECT 322.950 714.600 325.050 715.050 ;
        RECT 335.400 714.600 336.600 715.950 ;
        RECT 322.950 713.400 336.600 714.600 ;
        RECT 496.950 714.600 499.050 715.050 ;
        RECT 505.950 714.600 508.050 715.050 ;
        RECT 496.950 713.400 508.050 714.600 ;
        RECT 322.950 712.950 325.050 713.400 ;
        RECT 496.950 712.950 499.050 713.400 ;
        RECT 505.950 712.950 508.050 713.400 ;
        RECT 580.950 714.600 583.050 715.050 ;
        RECT 604.950 714.600 607.050 715.050 ;
        RECT 580.950 713.400 607.050 714.600 ;
        RECT 580.950 712.950 583.050 713.400 ;
        RECT 604.950 712.950 607.050 713.400 ;
        RECT 634.950 714.600 637.050 715.050 ;
        RECT 703.950 714.600 706.050 715.050 ;
        RECT 634.950 713.400 706.050 714.600 ;
        RECT 634.950 712.950 637.050 713.400 ;
        RECT 703.950 712.950 706.050 713.400 ;
        RECT 46.950 711.600 49.050 712.050 ;
        RECT 133.950 711.600 136.050 712.050 ;
        RECT 46.950 710.400 136.050 711.600 ;
        RECT 46.950 709.950 49.050 710.400 ;
        RECT 133.950 709.950 136.050 710.400 ;
        RECT 400.950 711.600 403.050 712.050 ;
        RECT 652.950 711.600 655.050 712.050 ;
        RECT 673.950 711.600 676.050 712.050 ;
        RECT 697.950 711.600 700.050 712.050 ;
        RECT 400.950 710.400 420.600 711.600 ;
        RECT 400.950 709.950 403.050 710.400 ;
        RECT 61.950 708.600 64.050 709.050 ;
        RECT 136.950 708.600 139.050 709.050 ;
        RECT 61.950 707.400 139.050 708.600 ;
        RECT 61.950 706.950 64.050 707.400 ;
        RECT 136.950 706.950 139.050 707.400 ;
        RECT 163.950 708.600 166.050 709.050 ;
        RECT 223.950 708.600 226.050 709.050 ;
        RECT 163.950 707.400 226.050 708.600 ;
        RECT 163.950 706.950 166.050 707.400 ;
        RECT 223.950 706.950 226.050 707.400 ;
        RECT 253.950 708.600 256.050 709.050 ;
        RECT 352.950 708.600 355.050 709.050 ;
        RECT 253.950 707.400 355.050 708.600 ;
        RECT 253.950 706.950 256.050 707.400 ;
        RECT 352.950 706.950 355.050 707.400 ;
        RECT 358.950 708.600 361.050 709.050 ;
        RECT 385.950 708.600 388.050 709.050 ;
        RECT 415.950 708.600 418.050 709.050 ;
        RECT 358.950 707.400 418.050 708.600 ;
        RECT 419.400 708.600 420.600 710.400 ;
        RECT 652.950 710.400 700.050 711.600 ;
        RECT 652.950 709.950 655.050 710.400 ;
        RECT 673.950 709.950 676.050 710.400 ;
        RECT 697.950 709.950 700.050 710.400 ;
        RECT 502.950 708.600 505.050 709.050 ;
        RECT 419.400 707.400 505.050 708.600 ;
        RECT 358.950 706.950 361.050 707.400 ;
        RECT 385.950 706.950 388.050 707.400 ;
        RECT 415.950 706.950 418.050 707.400 ;
        RECT 502.950 706.950 505.050 707.400 ;
        RECT 550.950 708.600 553.050 709.050 ;
        RECT 721.950 708.600 724.050 709.050 ;
        RECT 550.950 707.400 724.050 708.600 ;
        RECT 550.950 706.950 553.050 707.400 ;
        RECT 721.950 706.950 724.050 707.400 ;
        RECT 178.950 705.600 181.050 706.050 ;
        RECT 271.950 705.600 274.050 706.050 ;
        RECT 178.950 704.400 201.600 705.600 ;
        RECT 178.950 703.950 181.050 704.400 ;
        RECT 25.950 702.600 28.050 703.050 ;
        RECT 118.950 702.600 121.050 703.050 ;
        RECT 25.950 701.400 121.050 702.600 ;
        RECT 25.950 700.950 28.050 701.400 ;
        RECT 118.950 700.950 121.050 701.400 ;
        RECT 139.950 702.600 142.050 703.050 ;
        RECT 175.950 702.600 178.050 703.050 ;
        RECT 139.950 701.400 178.050 702.600 ;
        RECT 200.400 702.600 201.600 704.400 ;
        RECT 257.400 704.400 274.050 705.600 ;
        RECT 257.400 702.600 258.600 704.400 ;
        RECT 271.950 703.950 274.050 704.400 ;
        RECT 463.950 705.600 466.050 706.050 ;
        RECT 484.950 705.600 487.050 706.050 ;
        RECT 511.950 705.600 514.050 706.050 ;
        RECT 463.950 704.400 514.050 705.600 ;
        RECT 463.950 703.950 466.050 704.400 ;
        RECT 484.950 703.950 487.050 704.400 ;
        RECT 511.950 703.950 514.050 704.400 ;
        RECT 535.950 705.600 538.050 706.050 ;
        RECT 589.950 705.600 592.050 706.050 ;
        RECT 619.950 705.600 622.050 706.050 ;
        RECT 535.950 704.400 622.050 705.600 ;
        RECT 535.950 703.950 538.050 704.400 ;
        RECT 589.950 703.950 592.050 704.400 ;
        RECT 619.950 703.950 622.050 704.400 ;
        RECT 694.950 705.600 697.050 706.050 ;
        RECT 733.950 705.600 736.050 706.050 ;
        RECT 694.950 704.400 736.050 705.600 ;
        RECT 694.950 703.950 697.050 704.400 ;
        RECT 733.950 703.950 736.050 704.400 ;
        RECT 200.400 701.400 258.600 702.600 ;
        RECT 493.950 702.600 496.050 703.050 ;
        RECT 550.950 702.600 553.050 703.050 ;
        RECT 493.950 701.400 553.050 702.600 ;
        RECT 139.950 700.950 142.050 701.400 ;
        RECT 175.950 700.950 178.050 701.400 ;
        RECT 493.950 700.950 496.050 701.400 ;
        RECT 550.950 700.950 553.050 701.400 ;
        RECT 634.950 702.600 637.050 703.050 ;
        RECT 715.950 702.600 718.050 703.050 ;
        RECT 634.950 701.400 718.050 702.600 ;
        RECT 634.950 700.950 637.050 701.400 ;
        RECT 715.950 700.950 718.050 701.400 ;
        RECT 76.950 699.600 79.050 700.050 ;
        RECT 160.950 699.600 163.050 700.050 ;
        RECT 76.950 698.400 163.050 699.600 ;
        RECT 76.950 697.950 79.050 698.400 ;
        RECT 160.950 697.950 163.050 698.400 ;
        RECT 274.950 699.600 277.050 700.050 ;
        RECT 313.950 699.600 316.050 700.050 ;
        RECT 346.950 699.600 349.050 700.050 ;
        RECT 274.950 698.400 349.050 699.600 ;
        RECT 274.950 697.950 277.050 698.400 ;
        RECT 313.950 697.950 316.050 698.400 ;
        RECT 346.950 697.950 349.050 698.400 ;
        RECT 418.950 699.600 421.050 700.050 ;
        RECT 487.950 699.600 490.050 700.050 ;
        RECT 418.950 698.400 490.050 699.600 ;
        RECT 418.950 697.950 421.050 698.400 ;
        RECT 487.950 697.950 490.050 698.400 ;
        RECT 511.950 699.600 514.050 700.050 ;
        RECT 553.950 699.600 556.050 700.050 ;
        RECT 559.950 699.600 562.050 700.050 ;
        RECT 511.950 698.400 562.050 699.600 ;
        RECT 511.950 697.950 514.050 698.400 ;
        RECT 553.950 697.950 556.050 698.400 ;
        RECT 559.950 697.950 562.050 698.400 ;
        RECT 574.950 699.600 577.050 700.050 ;
        RECT 622.950 699.600 625.050 700.050 ;
        RECT 574.950 698.400 625.050 699.600 ;
        RECT 716.400 699.600 717.600 700.950 ;
        RECT 736.950 699.600 739.050 700.050 ;
        RECT 748.950 699.600 751.050 700.050 ;
        RECT 716.400 698.400 751.050 699.600 ;
        RECT 574.950 697.950 577.050 698.400 ;
        RECT 622.950 697.950 625.050 698.400 ;
        RECT 736.950 697.950 739.050 698.400 ;
        RECT 748.950 697.950 751.050 698.400 ;
        RECT 103.950 696.600 106.050 697.050 ;
        RECT 142.950 696.600 145.050 697.050 ;
        RECT 103.950 695.400 145.050 696.600 ;
        RECT 103.950 694.950 106.050 695.400 ;
        RECT 142.950 694.950 145.050 695.400 ;
        RECT 184.950 696.600 187.050 697.050 ;
        RECT 211.950 696.600 214.050 697.050 ;
        RECT 232.950 696.600 235.050 697.050 ;
        RECT 184.950 695.400 198.600 696.600 ;
        RECT 184.950 694.950 187.050 695.400 ;
        RECT 197.400 694.050 198.600 695.400 ;
        RECT 211.950 695.400 235.050 696.600 ;
        RECT 211.950 694.950 214.050 695.400 ;
        RECT 232.950 694.950 235.050 695.400 ;
        RECT 271.950 696.600 274.050 697.050 ;
        RECT 304.950 696.600 307.050 697.050 ;
        RECT 379.950 696.600 382.050 697.050 ;
        RECT 271.950 695.400 382.050 696.600 ;
        RECT 271.950 694.950 274.050 695.400 ;
        RECT 304.950 694.950 307.050 695.400 ;
        RECT 379.950 694.950 382.050 695.400 ;
        RECT 451.950 696.600 454.050 697.050 ;
        RECT 472.950 696.600 475.050 697.050 ;
        RECT 451.950 695.400 475.050 696.600 ;
        RECT 451.950 694.950 454.050 695.400 ;
        RECT 472.950 694.950 475.050 695.400 ;
        RECT 820.950 696.600 823.050 697.050 ;
        RECT 826.950 696.600 829.050 697.050 ;
        RECT 820.950 695.400 829.050 696.600 ;
        RECT 820.950 694.950 823.050 695.400 ;
        RECT 826.950 694.950 829.050 695.400 ;
        RECT 31.950 693.600 34.050 694.050 ;
        RECT 70.950 693.600 73.050 694.050 ;
        RECT 31.950 692.400 73.050 693.600 ;
        RECT 31.950 691.950 34.050 692.400 ;
        RECT 70.950 691.950 73.050 692.400 ;
        RECT 196.950 693.600 199.050 694.050 ;
        RECT 256.950 693.600 259.050 694.050 ;
        RECT 196.950 692.400 259.050 693.600 ;
        RECT 196.950 691.950 199.050 692.400 ;
        RECT 256.950 691.950 259.050 692.400 ;
        RECT 295.950 693.600 298.050 694.050 ;
        RECT 301.950 693.600 304.050 694.050 ;
        RECT 295.950 692.400 304.050 693.600 ;
        RECT 295.950 691.950 298.050 692.400 ;
        RECT 301.950 691.950 304.050 692.400 ;
        RECT 388.950 693.600 391.050 694.050 ;
        RECT 403.950 693.600 406.050 694.050 ;
        RECT 388.950 692.400 406.050 693.600 ;
        RECT 388.950 691.950 391.050 692.400 ;
        RECT 403.950 691.950 406.050 692.400 ;
        RECT 415.950 693.600 418.050 694.050 ;
        RECT 436.950 693.600 439.050 694.050 ;
        RECT 415.950 692.400 439.050 693.600 ;
        RECT 415.950 691.950 418.050 692.400 ;
        RECT 436.950 691.950 439.050 692.400 ;
        RECT 706.950 693.600 709.050 694.050 ;
        RECT 829.950 693.600 832.050 694.050 ;
        RECT 706.950 692.400 832.050 693.600 ;
        RECT 706.950 691.950 709.050 692.400 ;
        RECT 829.950 691.950 832.050 692.400 ;
        RECT 88.950 690.600 91.050 691.050 ;
        RECT 106.950 690.600 109.050 691.050 ;
        RECT 88.950 689.400 109.050 690.600 ;
        RECT 88.950 688.950 91.050 689.400 ;
        RECT 106.950 688.950 109.050 689.400 ;
        RECT 22.950 687.600 25.050 688.050 ;
        RECT 37.950 687.600 40.050 688.050 ;
        RECT 52.950 687.600 55.050 688.050 ;
        RECT 22.950 686.400 55.050 687.600 ;
        RECT 22.950 685.950 25.050 686.400 ;
        RECT 37.950 685.950 40.050 686.400 ;
        RECT 52.950 685.950 55.050 686.400 ;
        RECT 28.950 684.600 31.050 685.200 ;
        RECT 34.950 684.600 37.050 685.050 ;
        RECT 28.950 683.400 37.050 684.600 ;
        RECT 28.950 683.100 31.050 683.400 ;
        RECT 34.950 682.950 37.050 683.400 ;
        RECT 97.950 682.950 103.050 685.050 ;
        RECT 121.950 684.600 124.050 688.050 ;
        RECT 127.950 687.600 130.050 688.050 ;
        RECT 139.950 687.600 142.050 691.050 ;
        RECT 178.950 690.600 181.050 691.050 ;
        RECT 190.950 690.600 193.050 691.050 ;
        RECT 202.950 690.600 205.050 691.050 ;
        RECT 178.950 689.400 205.050 690.600 ;
        RECT 178.950 688.950 181.050 689.400 ;
        RECT 190.950 688.950 193.050 689.400 ;
        RECT 202.950 688.950 205.050 689.400 ;
        RECT 220.950 690.600 223.050 691.050 ;
        RECT 229.950 690.600 232.050 691.200 ;
        RECT 238.950 690.600 241.050 691.050 ;
        RECT 265.950 690.600 268.050 691.050 ;
        RECT 220.950 689.400 268.050 690.600 ;
        RECT 220.950 688.950 223.050 689.400 ;
        RECT 229.950 689.100 232.050 689.400 ;
        RECT 238.950 688.950 241.050 689.400 ;
        RECT 265.950 688.950 268.050 689.400 ;
        RECT 277.950 690.600 280.050 691.050 ;
        RECT 343.950 690.600 346.050 691.050 ;
        RECT 277.950 689.400 346.050 690.600 ;
        RECT 277.950 688.950 280.050 689.400 ;
        RECT 343.950 688.950 346.050 689.400 ;
        RECT 364.950 690.600 367.050 691.050 ;
        RECT 409.950 690.600 412.050 691.050 ;
        RECT 364.950 689.400 412.050 690.600 ;
        RECT 364.950 688.950 367.050 689.400 ;
        RECT 409.950 688.950 412.050 689.400 ;
        RECT 541.950 690.600 544.050 691.050 ;
        RECT 565.950 690.600 568.050 691.050 ;
        RECT 541.950 689.400 568.050 690.600 ;
        RECT 541.950 688.950 544.050 689.400 ;
        RECT 565.950 688.950 568.050 689.400 ;
        RECT 586.950 690.600 589.050 691.050 ;
        RECT 598.950 690.600 601.050 691.050 ;
        RECT 586.950 689.400 601.050 690.600 ;
        RECT 586.950 688.950 589.050 689.400 ;
        RECT 598.950 688.950 601.050 689.400 ;
        RECT 127.950 687.000 142.050 687.600 ;
        RECT 241.950 687.600 244.050 688.050 ;
        RECT 247.950 687.600 250.050 688.050 ;
        RECT 127.950 686.400 141.600 687.000 ;
        RECT 241.950 686.400 250.050 687.600 ;
        RECT 127.950 685.950 130.050 686.400 ;
        RECT 241.950 685.950 244.050 686.400 ;
        RECT 247.950 685.950 250.050 686.400 ;
        RECT 421.950 687.600 424.050 688.050 ;
        RECT 430.950 687.600 433.050 688.050 ;
        RECT 421.950 686.400 433.050 687.600 ;
        RECT 421.950 685.950 424.050 686.400 ;
        RECT 430.950 685.950 433.050 686.400 ;
        RECT 445.950 687.600 448.050 688.050 ;
        RECT 481.950 687.600 484.050 688.050 ;
        RECT 445.950 686.400 484.050 687.600 ;
        RECT 445.950 685.950 448.050 686.400 ;
        RECT 481.950 685.950 484.050 686.400 ;
        RECT 517.950 687.600 520.050 688.050 ;
        RECT 517.950 686.400 543.600 687.600 ;
        RECT 517.950 685.950 520.050 686.400 ;
        RECT 133.950 684.600 138.000 685.050 ;
        RECT 214.950 684.600 217.050 685.050 ;
        RECT 242.400 684.600 243.600 685.950 ;
        RECT 385.950 685.050 388.050 685.200 ;
        RECT 274.950 684.600 277.050 685.050 ;
        RECT 121.950 684.000 138.600 684.600 ;
        RECT 122.400 683.400 138.600 684.000 ;
        RECT 133.950 682.950 138.600 683.400 ;
        RECT 214.950 683.400 243.600 684.600 ;
        RECT 257.400 683.400 277.050 684.600 ;
        RECT 214.950 682.950 217.050 683.400 ;
        RECT 10.950 681.600 13.050 682.050 ;
        RECT 25.950 681.600 28.050 682.050 ;
        RECT 10.950 680.400 28.050 681.600 ;
        RECT 137.400 681.600 138.600 682.950 ;
        RECT 160.950 681.600 163.050 681.900 ;
        RECT 169.950 681.600 172.050 682.050 ;
        RECT 137.400 680.400 156.600 681.600 ;
        RECT 10.950 679.950 13.050 680.400 ;
        RECT 25.950 679.950 28.050 680.400 ;
        RECT 49.950 678.600 52.050 679.050 ;
        RECT 64.950 678.600 67.050 679.050 ;
        RECT 49.950 677.400 67.050 678.600 ;
        RECT 49.950 676.950 52.050 677.400 ;
        RECT 64.950 676.950 67.050 677.400 ;
        RECT 94.950 678.600 97.050 679.050 ;
        RECT 100.950 678.600 103.050 679.050 ;
        RECT 94.950 677.400 103.050 678.600 ;
        RECT 155.400 678.600 156.600 680.400 ;
        RECT 160.950 680.400 172.050 681.600 ;
        RECT 160.950 679.800 163.050 680.400 ;
        RECT 169.950 679.950 172.050 680.400 ;
        RECT 181.950 681.600 184.050 682.050 ;
        RECT 193.950 681.600 196.050 682.050 ;
        RECT 181.950 680.400 196.050 681.600 ;
        RECT 181.950 679.950 184.050 680.400 ;
        RECT 193.950 679.950 196.050 680.400 ;
        RECT 223.950 681.600 226.050 682.050 ;
        RECT 232.950 681.600 235.050 682.050 ;
        RECT 223.950 680.400 235.050 681.600 ;
        RECT 223.950 679.950 226.050 680.400 ;
        RECT 232.950 679.950 235.050 680.400 ;
        RECT 257.400 679.050 258.600 683.400 ;
        RECT 274.950 682.950 277.050 683.400 ;
        RECT 280.950 682.950 286.050 685.050 ;
        RECT 322.950 684.600 325.050 685.050 ;
        RECT 331.950 684.600 334.050 685.050 ;
        RECT 322.950 683.400 334.050 684.600 ;
        RECT 322.950 682.950 325.050 683.400 ;
        RECT 331.950 682.950 334.050 683.400 ;
        RECT 346.950 684.600 349.050 685.050 ;
        RECT 355.950 684.600 358.050 685.050 ;
        RECT 346.950 683.400 358.050 684.600 ;
        RECT 346.950 682.950 349.050 683.400 ;
        RECT 355.950 682.950 358.050 683.400 ;
        RECT 370.950 684.600 373.050 685.050 ;
        RECT 385.950 684.600 391.050 685.050 ;
        RECT 370.950 683.400 391.050 684.600 ;
        RECT 370.950 682.950 373.050 683.400 ;
        RECT 385.950 683.100 391.050 683.400 ;
        RECT 387.000 682.950 391.050 683.100 ;
        RECT 394.950 684.600 397.050 685.050 ;
        RECT 415.950 684.600 418.050 685.050 ;
        RECT 394.950 683.400 418.050 684.600 ;
        RECT 394.950 682.950 397.050 683.400 ;
        RECT 415.950 682.950 418.050 683.400 ;
        RECT 487.950 684.600 490.050 685.050 ;
        RECT 514.950 684.600 517.050 685.050 ;
        RECT 487.950 683.400 517.050 684.600 ;
        RECT 487.950 682.950 490.050 683.400 ;
        RECT 514.950 682.950 517.050 683.400 ;
        RECT 364.950 681.600 367.050 682.050 ;
        RECT 382.950 681.600 385.050 681.900 ;
        RECT 364.950 680.400 385.050 681.600 ;
        RECT 364.950 679.950 367.050 680.400 ;
        RECT 382.950 679.800 385.050 680.400 ;
        RECT 424.950 681.600 427.050 682.050 ;
        RECT 445.950 681.600 448.050 681.900 ;
        RECT 454.950 681.600 457.050 682.050 ;
        RECT 424.950 680.400 457.050 681.600 ;
        RECT 424.950 679.950 427.050 680.400 ;
        RECT 445.950 679.800 448.050 680.400 ;
        RECT 454.950 679.950 457.050 680.400 ;
        RECT 520.950 681.600 523.050 682.050 ;
        RECT 535.950 681.600 538.050 682.050 ;
        RECT 542.400 681.900 543.600 686.400 ;
        RECT 583.950 685.950 586.050 688.050 ;
        RECT 700.950 687.600 703.050 688.200 ;
        RECT 709.950 687.600 712.050 688.050 ;
        RECT 700.950 686.400 712.050 687.600 ;
        RECT 700.950 686.100 703.050 686.400 ;
        RECT 709.950 685.950 712.050 686.400 ;
        RECT 739.950 687.600 742.050 688.050 ;
        RECT 751.950 687.600 754.050 688.050 ;
        RECT 739.950 686.400 754.050 687.600 ;
        RECT 739.950 685.950 742.050 686.400 ;
        RECT 751.950 685.950 754.050 686.400 ;
        RECT 787.800 687.000 789.900 688.050 ;
        RECT 791.100 687.600 793.200 688.050 ;
        RECT 799.950 687.600 802.050 688.050 ;
        RECT 787.800 685.950 790.050 687.000 ;
        RECT 791.100 686.400 802.050 687.600 ;
        RECT 791.100 685.950 793.200 686.400 ;
        RECT 799.950 685.950 802.050 686.400 ;
        RECT 584.400 682.050 585.600 685.950 ;
        RECT 652.950 684.600 655.050 685.050 ;
        RECT 661.950 684.600 664.050 685.050 ;
        RECT 652.950 683.400 664.050 684.600 ;
        RECT 652.950 682.950 655.050 683.400 ;
        RECT 661.950 682.950 664.050 683.400 ;
        RECT 682.950 684.600 685.050 685.200 ;
        RECT 700.950 684.600 703.050 684.900 ;
        RECT 682.950 683.400 703.050 684.600 ;
        RECT 682.950 683.100 685.050 683.400 ;
        RECT 700.950 682.800 703.050 683.400 ;
        RECT 772.950 684.600 775.050 685.050 ;
        RECT 787.950 684.600 790.050 685.950 ;
        RECT 808.950 684.600 811.050 685.050 ;
        RECT 772.950 683.400 783.600 684.600 ;
        RECT 787.950 684.000 811.050 684.600 ;
        RECT 788.250 683.400 811.050 684.000 ;
        RECT 772.950 682.950 775.050 683.400 ;
        RECT 782.400 682.050 783.600 683.400 ;
        RECT 808.950 682.950 811.050 683.400 ;
        RECT 520.950 680.400 538.050 681.600 ;
        RECT 520.950 679.950 523.050 680.400 ;
        RECT 535.950 679.950 538.050 680.400 ;
        RECT 541.950 679.800 544.050 681.900 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 631.950 681.600 634.050 681.900 ;
        RECT 670.950 681.600 673.050 682.050 ;
        RECT 682.950 681.600 685.050 681.900 ;
        RECT 703.950 681.600 706.050 681.900 ;
        RECT 631.950 681.000 648.600 681.600 ;
        RECT 631.950 680.400 649.050 681.000 ;
        RECT 631.950 679.800 634.050 680.400 ;
        RECT 241.950 678.600 244.050 679.050 ;
        RECT 155.400 677.400 244.050 678.600 ;
        RECT 94.950 676.950 97.050 677.400 ;
        RECT 100.950 676.950 103.050 677.400 ;
        RECT 241.950 676.950 244.050 677.400 ;
        RECT 256.950 676.950 259.050 679.050 ;
        RECT 277.950 678.600 280.050 679.050 ;
        RECT 295.950 678.600 298.050 679.050 ;
        RECT 277.950 677.400 298.050 678.600 ;
        RECT 277.950 676.950 280.050 677.400 ;
        RECT 295.950 676.950 298.050 677.400 ;
        RECT 334.950 678.600 337.050 678.900 ;
        RECT 349.950 678.600 352.050 679.050 ;
        RECT 334.950 677.400 352.050 678.600 ;
        RECT 334.950 676.800 337.050 677.400 ;
        RECT 349.950 676.950 352.050 677.400 ;
        RECT 391.950 678.600 394.050 679.050 ;
        RECT 412.950 678.600 415.050 679.050 ;
        RECT 391.950 677.400 415.050 678.600 ;
        RECT 391.950 676.950 394.050 677.400 ;
        RECT 412.950 676.950 415.050 677.400 ;
        RECT 571.950 678.600 574.050 679.050 ;
        RECT 586.950 678.600 589.050 679.050 ;
        RECT 571.950 677.400 589.050 678.600 ;
        RECT 571.950 676.950 574.050 677.400 ;
        RECT 586.950 676.950 589.050 677.400 ;
        RECT 592.950 678.600 595.050 679.050 ;
        RECT 613.950 678.600 616.050 679.050 ;
        RECT 625.950 678.600 628.050 679.200 ;
        RECT 592.950 677.400 628.050 678.600 ;
        RECT 592.950 676.950 595.050 677.400 ;
        RECT 613.950 676.950 616.050 677.400 ;
        RECT 625.950 677.100 628.050 677.400 ;
        RECT 646.950 678.600 649.050 680.400 ;
        RECT 670.950 680.400 706.050 681.600 ;
        RECT 670.950 679.950 673.050 680.400 ;
        RECT 682.950 679.800 685.050 680.400 ;
        RECT 703.950 679.800 706.050 680.400 ;
        RECT 781.950 681.600 784.050 682.050 ;
        RECT 823.950 681.600 826.050 682.050 ;
        RECT 781.950 680.400 826.050 681.600 ;
        RECT 781.950 679.950 784.050 680.400 ;
        RECT 823.950 679.950 826.050 680.400 ;
        RECT 658.950 678.600 661.050 679.050 ;
        RECT 646.950 677.400 661.050 678.600 ;
        RECT 646.950 676.950 649.050 677.400 ;
        RECT 658.950 676.950 661.050 677.400 ;
        RECT 712.950 678.600 715.050 679.050 ;
        RECT 736.950 678.600 739.050 679.050 ;
        RECT 747.000 678.600 751.050 679.050 ;
        RECT 760.950 678.600 763.050 679.050 ;
        RECT 712.950 677.400 739.050 678.600 ;
        RECT 746.400 677.400 763.050 678.600 ;
        RECT 712.950 676.950 715.050 677.400 ;
        RECT 736.950 676.950 739.050 677.400 ;
        RECT 747.000 676.950 751.050 677.400 ;
        RECT 760.950 676.950 763.050 677.400 ;
        RECT 766.950 678.600 769.050 679.050 ;
        RECT 775.950 678.600 778.050 679.050 ;
        RECT 766.950 677.400 778.050 678.600 ;
        RECT 766.950 676.950 769.050 677.400 ;
        RECT 775.950 676.950 778.050 677.400 ;
        RECT 28.950 675.600 31.050 676.050 ;
        RECT 46.950 675.600 49.050 676.050 ;
        RECT 28.950 674.400 49.050 675.600 ;
        RECT 28.950 673.950 31.050 674.400 ;
        RECT 46.950 673.950 49.050 674.400 ;
        RECT 151.950 675.600 154.050 676.050 ;
        RECT 259.950 675.600 262.050 676.050 ;
        RECT 151.950 674.400 262.050 675.600 ;
        RECT 151.950 673.950 154.050 674.400 ;
        RECT 259.950 673.950 262.050 674.400 ;
        RECT 268.950 675.600 271.050 676.050 ;
        RECT 292.950 675.600 295.050 676.050 ;
        RECT 367.950 675.600 370.050 676.050 ;
        RECT 268.950 674.400 295.050 675.600 ;
        RECT 268.950 673.950 271.050 674.400 ;
        RECT 292.950 673.950 295.050 674.400 ;
        RECT 353.400 674.400 370.050 675.600 ;
        RECT 106.950 672.600 109.050 673.050 ;
        RECT 136.950 672.600 139.050 673.050 ;
        RECT 106.950 671.400 139.050 672.600 ;
        RECT 106.950 670.950 109.050 671.400 ;
        RECT 136.950 670.950 139.050 671.400 ;
        RECT 343.950 672.600 346.050 673.050 ;
        RECT 353.400 672.600 354.600 674.400 ;
        RECT 367.950 673.950 370.050 674.400 ;
        RECT 541.950 675.600 544.050 676.050 ;
        RECT 565.950 675.600 568.050 676.200 ;
        RECT 541.950 674.400 568.050 675.600 ;
        RECT 541.950 673.950 544.050 674.400 ;
        RECT 565.950 674.100 568.050 674.400 ;
        RECT 625.950 675.600 628.050 675.900 ;
        RECT 676.950 675.600 679.050 676.050 ;
        RECT 625.950 674.400 679.050 675.600 ;
        RECT 625.950 673.800 628.050 674.400 ;
        RECT 676.950 673.950 679.050 674.400 ;
        RECT 343.950 671.400 354.600 672.600 ;
        RECT 424.950 672.600 427.050 673.050 ;
        RECT 436.950 672.600 439.050 673.050 ;
        RECT 424.950 671.400 439.050 672.600 ;
        RECT 343.950 670.950 346.050 671.400 ;
        RECT 424.950 670.950 427.050 671.400 ;
        RECT 436.950 670.950 439.050 671.400 ;
        RECT 517.950 672.600 520.050 673.050 ;
        RECT 538.950 672.600 541.050 673.050 ;
        RECT 544.950 672.600 547.050 673.050 ;
        RECT 517.950 671.400 547.050 672.600 ;
        RECT 517.950 670.950 520.050 671.400 ;
        RECT 538.950 670.950 541.050 671.400 ;
        RECT 544.950 670.950 547.050 671.400 ;
        RECT 568.950 672.600 571.050 672.900 ;
        RECT 607.800 672.600 609.900 673.050 ;
        RECT 568.950 671.400 609.900 672.600 ;
        RECT 568.950 670.800 571.050 671.400 ;
        RECT 607.800 670.950 609.900 671.400 ;
        RECT 611.100 672.600 613.200 673.050 ;
        RECT 640.950 672.600 643.050 673.050 ;
        RECT 611.100 671.400 643.050 672.600 ;
        RECT 677.400 672.600 678.600 673.950 ;
        RECT 718.950 672.600 721.050 673.050 ;
        RECT 677.400 671.400 721.050 672.600 ;
        RECT 611.100 670.950 613.200 671.400 ;
        RECT 640.950 670.950 643.050 671.400 ;
        RECT 718.950 670.950 721.050 671.400 ;
        RECT 229.950 669.600 232.050 670.050 ;
        RECT 262.950 669.600 265.050 670.050 ;
        RECT 229.950 668.400 265.050 669.600 ;
        RECT 229.950 667.950 232.050 668.400 ;
        RECT 262.950 667.950 265.050 668.400 ;
        RECT 553.950 669.600 556.050 670.050 ;
        RECT 598.950 669.600 601.050 670.050 ;
        RECT 553.950 668.400 601.050 669.600 ;
        RECT 553.950 667.950 556.050 668.400 ;
        RECT 598.950 667.950 601.050 668.400 ;
        RECT 163.950 666.600 166.050 667.050 ;
        RECT 230.400 666.600 231.600 667.950 ;
        RECT 163.950 665.400 231.600 666.600 ;
        RECT 370.950 666.600 373.050 667.050 ;
        RECT 490.950 666.600 493.050 667.050 ;
        RECT 370.950 665.400 493.050 666.600 ;
        RECT 163.950 664.950 166.050 665.400 ;
        RECT 370.950 664.950 373.050 665.400 ;
        RECT 490.950 664.950 493.050 665.400 ;
        RECT 532.950 666.600 535.050 667.050 ;
        RECT 538.950 666.600 541.050 667.050 ;
        RECT 532.950 665.400 541.050 666.600 ;
        RECT 532.950 664.950 535.050 665.400 ;
        RECT 538.950 664.950 541.050 665.400 ;
        RECT 547.950 666.600 550.050 667.050 ;
        RECT 580.950 666.600 583.050 667.050 ;
        RECT 547.950 665.400 583.050 666.600 ;
        RECT 547.950 664.950 550.050 665.400 ;
        RECT 580.950 664.950 583.050 665.400 ;
        RECT 607.950 666.600 610.050 667.050 ;
        RECT 634.950 666.600 637.050 667.050 ;
        RECT 607.950 665.400 637.050 666.600 ;
        RECT 607.950 664.950 610.050 665.400 ;
        RECT 634.950 664.950 637.050 665.400 ;
        RECT 103.950 663.600 106.050 664.050 ;
        RECT 130.950 663.600 133.050 664.050 ;
        RECT 103.950 662.400 133.050 663.600 ;
        RECT 103.950 661.950 106.050 662.400 ;
        RECT 130.950 661.950 133.050 662.400 ;
        RECT 148.950 663.600 151.050 664.050 ;
        RECT 169.950 663.600 172.050 664.050 ;
        RECT 148.950 662.400 172.050 663.600 ;
        RECT 148.950 661.950 151.050 662.400 ;
        RECT 169.950 661.950 172.050 662.400 ;
        RECT 217.950 663.600 220.050 664.050 ;
        RECT 280.950 663.600 283.050 664.050 ;
        RECT 217.950 662.400 283.050 663.600 ;
        RECT 217.950 661.950 220.050 662.400 ;
        RECT 280.950 661.950 283.050 662.400 ;
        RECT 307.950 663.600 310.050 664.050 ;
        RECT 319.950 663.600 322.050 664.050 ;
        RECT 328.950 663.600 331.050 664.050 ;
        RECT 307.950 662.400 331.050 663.600 ;
        RECT 307.950 661.950 310.050 662.400 ;
        RECT 319.950 661.950 322.050 662.400 ;
        RECT 328.950 661.950 331.050 662.400 ;
        RECT 364.950 663.600 367.050 664.050 ;
        RECT 391.950 663.600 394.050 664.050 ;
        RECT 364.950 662.400 394.050 663.600 ;
        RECT 364.950 661.950 367.050 662.400 ;
        RECT 391.950 661.950 394.050 662.400 ;
        RECT 667.950 663.600 670.050 664.050 ;
        RECT 697.950 663.600 700.050 664.050 ;
        RECT 667.950 662.400 700.050 663.600 ;
        RECT 667.950 661.950 670.050 662.400 ;
        RECT 697.950 661.950 700.050 662.400 ;
        RECT 151.950 660.600 154.050 661.050 ;
        RECT 163.950 660.600 166.050 661.050 ;
        RECT 151.950 659.400 166.050 660.600 ;
        RECT 151.950 658.950 154.050 659.400 ;
        RECT 163.950 658.950 166.050 659.400 ;
        RECT 175.950 660.600 178.050 661.050 ;
        RECT 256.950 660.600 259.050 661.050 ;
        RECT 175.950 659.400 259.050 660.600 ;
        RECT 175.950 658.950 178.050 659.400 ;
        RECT 256.950 658.950 259.050 659.400 ;
        RECT 460.950 660.600 463.050 661.050 ;
        RECT 499.950 660.600 502.050 661.050 ;
        RECT 460.950 659.400 502.050 660.600 ;
        RECT 460.950 658.950 463.050 659.400 ;
        RECT 499.950 658.950 502.050 659.400 ;
        RECT 511.950 660.600 514.050 661.050 ;
        RECT 529.950 660.600 532.050 661.050 ;
        RECT 553.950 660.600 556.050 661.050 ;
        RECT 511.950 659.400 556.050 660.600 ;
        RECT 511.950 658.950 514.050 659.400 ;
        RECT 529.950 658.950 532.050 659.400 ;
        RECT 553.950 658.950 556.050 659.400 ;
        RECT 571.950 660.600 574.050 661.050 ;
        RECT 625.800 660.600 627.900 661.050 ;
        RECT 571.950 659.400 627.900 660.600 ;
        RECT 571.950 658.950 574.050 659.400 ;
        RECT 625.800 658.950 627.900 659.400 ;
        RECT 629.100 660.600 631.200 661.050 ;
        RECT 634.950 660.600 637.050 661.050 ;
        RECT 629.100 659.400 637.050 660.600 ;
        RECT 629.100 658.950 631.200 659.400 ;
        RECT 634.950 658.950 637.050 659.400 ;
        RECT 643.950 660.600 646.050 661.050 ;
        RECT 721.950 660.600 724.050 661.050 ;
        RECT 730.950 660.600 733.050 661.050 ;
        RECT 805.950 660.600 808.050 661.050 ;
        RECT 643.950 659.400 808.050 660.600 ;
        RECT 643.950 658.950 646.050 659.400 ;
        RECT 721.950 658.950 724.050 659.400 ;
        RECT 730.950 658.950 733.050 659.400 ;
        RECT 805.950 658.950 808.050 659.400 ;
        RECT 46.950 657.600 49.050 658.050 ;
        RECT 55.950 657.600 58.050 658.050 ;
        RECT 46.950 656.400 58.050 657.600 ;
        RECT 46.950 655.950 49.050 656.400 ;
        RECT 55.950 655.950 58.050 656.400 ;
        RECT 64.950 657.600 67.050 658.050 ;
        RECT 70.950 657.600 73.050 658.200 ;
        RECT 64.950 656.400 73.050 657.600 ;
        RECT 64.950 655.950 67.050 656.400 ;
        RECT 70.950 656.100 73.050 656.400 ;
        RECT 145.950 657.600 148.050 658.050 ;
        RECT 172.950 657.600 175.050 658.050 ;
        RECT 145.950 656.400 175.050 657.600 ;
        RECT 145.950 655.950 148.050 656.400 ;
        RECT 172.950 655.950 175.050 656.400 ;
        RECT 211.950 657.600 214.050 658.200 ;
        RECT 229.950 657.600 232.050 658.050 ;
        RECT 211.950 656.400 232.050 657.600 ;
        RECT 211.950 656.100 214.050 656.400 ;
        RECT 229.950 655.950 232.050 656.400 ;
        RECT 295.950 657.600 298.050 658.050 ;
        RECT 316.950 657.600 319.050 658.050 ;
        RECT 295.950 656.400 319.050 657.600 ;
        RECT 295.950 655.950 298.050 656.400 ;
        RECT 316.950 655.950 319.050 656.400 ;
        RECT 367.950 657.600 370.050 658.050 ;
        RECT 421.950 657.600 424.050 658.050 ;
        RECT 451.950 657.600 454.050 658.050 ;
        RECT 367.950 656.400 454.050 657.600 ;
        RECT 367.950 655.950 370.050 656.400 ;
        RECT 421.950 655.950 424.050 656.400 ;
        RECT 451.950 655.950 454.050 656.400 ;
        RECT 502.950 657.600 505.050 658.050 ;
        RECT 568.950 657.600 571.050 658.050 ;
        RECT 502.950 656.400 571.050 657.600 ;
        RECT 502.950 655.950 505.050 656.400 ;
        RECT 568.950 655.950 571.050 656.400 ;
        RECT 574.950 657.600 577.050 658.050 ;
        RECT 586.950 657.600 589.050 658.050 ;
        RECT 574.950 656.400 589.050 657.600 ;
        RECT 574.950 655.950 577.050 656.400 ;
        RECT 586.950 655.950 589.050 656.400 ;
        RECT 604.950 657.600 607.050 658.050 ;
        RECT 616.950 657.600 619.050 658.050 ;
        RECT 604.950 656.400 619.050 657.600 ;
        RECT 604.950 655.950 607.050 656.400 ;
        RECT 616.950 655.950 619.050 656.400 ;
        RECT 673.950 657.600 676.050 658.050 ;
        RECT 682.950 657.600 685.050 658.050 ;
        RECT 673.950 656.400 685.050 657.600 ;
        RECT 673.950 655.950 676.050 656.400 ;
        RECT 682.950 655.950 685.050 656.400 ;
        RECT 13.950 654.600 16.050 655.050 ;
        RECT 52.950 654.600 55.050 655.050 ;
        RECT 70.950 654.600 73.050 654.900 ;
        RECT 13.950 653.400 73.050 654.600 ;
        RECT 13.950 652.950 16.050 653.400 ;
        RECT 52.950 652.950 55.050 653.400 ;
        RECT 70.950 652.800 73.050 653.400 ;
        RECT 127.950 651.600 130.050 655.200 ;
        RECT 202.950 654.600 205.050 655.200 ;
        RECT 211.950 654.600 214.050 654.900 ;
        RECT 202.950 653.400 214.050 654.600 ;
        RECT 202.950 653.100 205.050 653.400 ;
        RECT 211.950 652.800 214.050 653.400 ;
        RECT 289.950 654.600 292.050 655.050 ;
        RECT 301.950 654.600 304.050 655.050 ;
        RECT 289.950 653.400 304.050 654.600 ;
        RECT 289.950 652.950 292.050 653.400 ;
        RECT 301.950 652.950 304.050 653.400 ;
        RECT 472.950 654.600 475.050 655.050 ;
        RECT 499.950 654.600 502.050 655.050 ;
        RECT 472.950 653.400 502.050 654.600 ;
        RECT 472.950 652.950 475.050 653.400 ;
        RECT 499.950 652.950 502.050 653.400 ;
        RECT 739.950 654.600 742.050 655.050 ;
        RECT 784.950 654.600 787.050 655.050 ;
        RECT 739.950 653.400 787.050 654.600 ;
        RECT 739.950 652.950 742.050 653.400 ;
        RECT 784.950 652.950 787.050 653.400 ;
        RECT 133.950 651.600 136.050 652.050 ;
        RECT 127.950 651.000 136.050 651.600 ;
        RECT 128.400 650.400 136.050 651.000 ;
        RECT 133.950 649.950 136.050 650.400 ;
        RECT 343.950 651.600 346.050 652.200 ;
        RECT 352.950 651.600 355.050 652.050 ;
        RECT 343.950 650.400 355.050 651.600 ;
        RECT 343.950 650.100 346.050 650.400 ;
        RECT 352.950 649.950 355.050 650.400 ;
        RECT 388.950 651.600 391.050 652.050 ;
        RECT 394.950 651.600 397.050 652.050 ;
        RECT 388.950 650.400 397.050 651.600 ;
        RECT 388.950 649.950 391.050 650.400 ;
        RECT 394.950 649.950 397.050 650.400 ;
        RECT 451.950 651.600 454.050 652.050 ;
        RECT 463.950 651.600 466.050 652.200 ;
        RECT 451.950 650.400 466.050 651.600 ;
        RECT 500.400 651.600 501.600 652.950 ;
        RECT 514.950 651.600 517.050 652.050 ;
        RECT 550.950 651.600 553.050 652.050 ;
        RECT 568.950 651.600 571.050 652.050 ;
        RECT 622.950 651.600 625.050 652.050 ;
        RECT 500.400 650.400 517.050 651.600 ;
        RECT 451.950 649.950 454.050 650.400 ;
        RECT 463.950 650.100 466.050 650.400 ;
        RECT 514.950 649.950 517.050 650.400 ;
        RECT 524.400 650.400 571.050 651.600 ;
        RECT 614.400 651.000 625.050 651.600 ;
        RECT 145.950 649.050 148.050 649.200 ;
        RECT 19.950 648.600 22.050 649.050 ;
        RECT 19.950 648.000 33.600 648.600 ;
        RECT 19.950 647.400 34.050 648.000 ;
        RECT 19.950 646.950 22.050 647.400 ;
        RECT 31.950 643.950 34.050 647.400 ;
        RECT 142.950 647.100 148.050 649.050 ;
        RECT 313.950 648.600 316.050 649.050 ;
        RECT 340.800 648.600 342.900 648.900 ;
        RECT 313.950 647.400 342.900 648.600 ;
        RECT 142.950 646.950 147.000 647.100 ;
        RECT 313.950 646.950 316.050 647.400 ;
        RECT 340.800 646.800 342.900 647.400 ;
        RECT 344.100 648.600 346.200 648.900 ;
        RECT 382.950 648.600 385.050 649.050 ;
        RECT 344.100 647.400 385.050 648.600 ;
        RECT 344.100 646.800 346.200 647.400 ;
        RECT 382.950 646.950 385.050 647.400 ;
        RECT 403.950 648.600 406.050 649.050 ;
        RECT 436.950 648.600 439.050 649.050 ;
        RECT 403.950 647.400 439.050 648.600 ;
        RECT 403.950 646.950 406.050 647.400 ;
        RECT 436.950 646.950 439.050 647.400 ;
        RECT 463.950 648.600 466.050 648.900 ;
        RECT 478.950 648.600 481.050 649.200 ;
        RECT 524.400 648.600 525.600 650.400 ;
        RECT 550.950 649.950 553.050 650.400 ;
        RECT 568.950 649.950 571.050 650.400 ;
        RECT 613.950 650.400 625.050 651.000 ;
        RECT 463.950 647.400 481.050 648.600 ;
        RECT 463.950 646.800 466.050 647.400 ;
        RECT 478.950 647.100 481.050 647.400 ;
        RECT 521.400 647.400 525.600 648.600 ;
        RECT 580.950 648.600 583.050 649.050 ;
        RECT 601.950 648.600 604.050 649.050 ;
        RECT 580.950 647.400 604.050 648.600 ;
        RECT 52.950 645.600 55.050 645.900 ;
        RECT 64.800 645.600 66.900 646.050 ;
        RECT 52.950 644.400 66.900 645.600 ;
        RECT 52.950 643.800 55.050 644.400 ;
        RECT 64.800 643.950 66.900 644.400 ;
        RECT 68.100 645.600 70.200 646.050 ;
        RECT 82.950 645.600 85.050 646.050 ;
        RECT 68.100 644.400 85.050 645.600 ;
        RECT 68.100 643.950 70.200 644.400 ;
        RECT 82.950 643.950 85.050 644.400 ;
        RECT 106.950 645.600 109.050 646.050 ;
        RECT 127.950 645.600 130.050 646.050 ;
        RECT 151.800 645.600 153.900 646.200 ;
        RECT 277.950 646.050 280.050 646.200 ;
        RECT 106.950 644.400 153.900 645.600 ;
        RECT 106.950 643.950 109.050 644.400 ;
        RECT 127.950 643.950 130.050 644.400 ;
        RECT 112.950 642.600 115.050 643.050 ;
        RECT 118.950 642.600 121.050 643.050 ;
        RECT 112.950 641.400 121.050 642.600 ;
        RECT 112.950 640.950 115.050 641.400 ;
        RECT 118.950 640.950 121.050 641.400 ;
        RECT 145.950 640.800 148.050 644.400 ;
        RECT 151.800 644.100 153.900 644.400 ;
        RECT 163.950 645.600 166.050 646.050 ;
        RECT 190.950 645.600 193.050 646.050 ;
        RECT 163.950 644.400 193.050 645.600 ;
        RECT 163.950 643.950 166.050 644.400 ;
        RECT 190.950 643.950 193.050 644.400 ;
        RECT 253.950 645.600 256.050 646.050 ;
        RECT 277.950 645.600 283.050 646.050 ;
        RECT 253.950 644.400 283.050 645.600 ;
        RECT 253.950 643.950 256.050 644.400 ;
        RECT 277.950 644.100 283.050 644.400 ;
        RECT 279.000 643.950 283.050 644.100 ;
        RECT 319.950 645.600 322.050 645.900 ;
        RECT 328.950 645.600 331.050 646.050 ;
        RECT 319.950 644.400 331.050 645.600 ;
        RECT 319.950 643.800 322.050 644.400 ;
        RECT 328.950 643.950 331.050 644.400 ;
        RECT 400.950 645.600 403.050 646.050 ;
        RECT 430.950 645.600 433.050 646.050 ;
        RECT 451.950 645.600 454.050 646.050 ;
        RECT 400.950 645.000 411.600 645.600 ;
        RECT 400.950 644.400 412.050 645.000 ;
        RECT 400.950 643.950 403.050 644.400 ;
        RECT 181.950 642.600 184.050 643.050 ;
        RECT 226.950 642.600 229.050 643.050 ;
        RECT 181.950 641.400 229.050 642.600 ;
        RECT 181.950 640.950 184.050 641.400 ;
        RECT 226.950 640.950 229.050 641.400 ;
        RECT 310.950 642.600 313.050 643.050 ;
        RECT 325.950 642.600 328.050 643.050 ;
        RECT 310.950 641.400 328.050 642.600 ;
        RECT 310.950 640.950 313.050 641.400 ;
        RECT 325.950 640.950 328.050 641.400 ;
        RECT 409.950 640.950 412.050 644.400 ;
        RECT 430.950 644.400 454.050 645.600 ;
        RECT 430.950 643.950 433.050 644.400 ;
        RECT 451.950 643.950 454.050 644.400 ;
        RECT 508.950 645.600 511.050 646.050 ;
        RECT 521.400 645.600 522.600 647.400 ;
        RECT 580.950 646.950 583.050 647.400 ;
        RECT 601.950 646.950 604.050 647.400 ;
        RECT 613.950 646.950 616.050 650.400 ;
        RECT 622.950 649.950 625.050 650.400 ;
        RECT 658.950 651.600 661.050 652.050 ;
        RECT 670.950 651.600 673.050 652.050 ;
        RECT 688.950 651.600 691.050 652.050 ;
        RECT 658.950 650.400 691.050 651.600 ;
        RECT 658.950 649.950 661.050 650.400 ;
        RECT 670.950 649.950 673.050 650.400 ;
        RECT 688.950 649.950 691.050 650.400 ;
        RECT 712.950 648.600 715.050 649.050 ;
        RECT 724.950 648.600 727.050 649.200 ;
        RECT 733.950 648.600 736.050 652.050 ;
        RECT 742.950 651.600 745.050 652.050 ;
        RECT 775.950 651.600 778.050 652.050 ;
        RECT 742.950 650.400 778.050 651.600 ;
        RECT 742.950 649.950 745.050 650.400 ;
        RECT 775.950 649.950 778.050 650.400 ;
        RECT 712.950 648.000 736.050 648.600 ;
        RECT 712.950 647.400 735.600 648.000 ;
        RECT 712.950 646.950 715.050 647.400 ;
        RECT 724.950 647.100 727.050 647.400 ;
        RECT 778.950 646.950 784.050 649.050 ;
        RECT 787.950 648.600 790.050 649.050 ;
        RECT 796.950 648.600 799.050 649.050 ;
        RECT 787.950 647.400 799.050 648.600 ;
        RECT 787.950 646.950 790.050 647.400 ;
        RECT 796.950 646.950 799.050 647.400 ;
        RECT 823.950 646.950 829.050 649.050 ;
        RECT 508.950 644.400 522.600 645.600 ;
        RECT 526.950 645.600 529.050 646.050 ;
        RECT 532.950 645.600 535.050 646.050 ;
        RECT 526.950 644.400 535.050 645.600 ;
        RECT 508.950 643.950 511.050 644.400 ;
        RECT 526.950 643.950 529.050 644.400 ;
        RECT 532.950 643.950 535.050 644.400 ;
        RECT 544.950 645.600 547.050 646.050 ;
        RECT 589.950 645.600 592.050 646.050 ;
        RECT 544.950 644.400 592.050 645.600 ;
        RECT 544.950 643.950 547.050 644.400 ;
        RECT 589.950 643.950 592.050 644.400 ;
        RECT 598.950 645.600 601.050 646.050 ;
        RECT 607.950 645.600 610.050 646.050 ;
        RECT 598.950 644.400 610.050 645.600 ;
        RECT 598.950 643.950 601.050 644.400 ;
        RECT 607.950 643.950 610.050 644.400 ;
        RECT 757.950 645.600 760.050 646.050 ;
        RECT 769.950 645.600 772.050 646.050 ;
        RECT 757.950 644.400 772.050 645.600 ;
        RECT 757.950 643.950 760.050 644.400 ;
        RECT 769.950 643.950 772.050 644.400 ;
        RECT 523.950 642.600 526.050 643.050 ;
        RECT 541.950 642.600 544.050 643.050 ;
        RECT 523.950 641.400 544.050 642.600 ;
        RECT 523.950 640.950 526.050 641.400 ;
        RECT 541.950 640.950 544.050 641.400 ;
        RECT 550.950 642.600 553.050 643.050 ;
        RECT 574.950 642.600 577.050 643.050 ;
        RECT 550.950 641.400 577.050 642.600 ;
        RECT 550.950 640.950 553.050 641.400 ;
        RECT 574.950 640.950 577.050 641.400 ;
        RECT 628.950 642.600 631.050 643.050 ;
        RECT 637.950 642.600 640.050 643.050 ;
        RECT 628.950 641.400 640.050 642.600 ;
        RECT 628.950 640.950 631.050 641.400 ;
        RECT 637.950 640.950 640.050 641.400 ;
        RECT 670.950 642.600 673.050 643.050 ;
        RECT 676.950 642.600 679.050 643.050 ;
        RECT 694.950 642.600 697.050 643.050 ;
        RECT 670.950 641.400 697.050 642.600 ;
        RECT 670.950 640.950 673.050 641.400 ;
        RECT 676.950 640.950 679.050 641.400 ;
        RECT 694.950 640.950 697.050 641.400 ;
        RECT 760.950 642.600 763.050 643.050 ;
        RECT 766.950 642.600 769.050 643.050 ;
        RECT 772.950 642.600 775.050 643.050 ;
        RECT 760.950 641.400 775.050 642.600 ;
        RECT 760.950 640.950 763.050 641.400 ;
        RECT 766.950 640.950 769.050 641.400 ;
        RECT 772.950 640.950 775.050 641.400 ;
        RECT 799.950 642.600 802.050 643.050 ;
        RECT 817.950 642.600 820.050 643.050 ;
        RECT 799.950 641.400 820.050 642.600 ;
        RECT 799.950 640.950 802.050 641.400 ;
        RECT 817.950 640.950 820.050 641.400 ;
        RECT 94.950 639.600 97.050 640.050 ;
        RECT 205.950 639.600 208.050 640.050 ;
        RECT 94.950 638.400 208.050 639.600 ;
        RECT 94.950 637.950 97.050 638.400 ;
        RECT 205.950 637.950 208.050 638.400 ;
        RECT 286.950 639.600 289.050 640.050 ;
        RECT 433.950 639.600 436.050 640.050 ;
        RECT 445.800 639.600 447.900 640.050 ;
        RECT 286.950 639.000 315.600 639.600 ;
        RECT 286.950 638.400 316.050 639.000 ;
        RECT 286.950 637.950 289.050 638.400 ;
        RECT 292.950 636.600 295.050 637.050 ;
        RECT 301.950 636.600 304.050 637.050 ;
        RECT 292.950 635.400 304.050 636.600 ;
        RECT 292.950 634.950 295.050 635.400 ;
        RECT 301.950 634.950 304.050 635.400 ;
        RECT 313.950 634.950 316.050 638.400 ;
        RECT 433.950 638.400 447.900 639.600 ;
        RECT 433.950 637.950 436.050 638.400 ;
        RECT 445.800 637.950 447.900 638.400 ;
        RECT 449.100 639.600 451.200 640.050 ;
        RECT 526.950 639.600 529.050 640.050 ;
        RECT 449.100 638.400 529.050 639.600 ;
        RECT 449.100 637.950 451.200 638.400 ;
        RECT 526.950 637.950 529.050 638.400 ;
        RECT 553.950 639.600 556.050 640.050 ;
        RECT 559.950 639.600 562.050 640.050 ;
        RECT 553.950 638.400 562.050 639.600 ;
        RECT 553.950 637.950 556.050 638.400 ;
        RECT 559.950 637.950 562.050 638.400 ;
        RECT 586.950 639.600 589.050 640.050 ;
        RECT 610.950 639.600 613.050 640.050 ;
        RECT 586.950 638.400 613.050 639.600 ;
        RECT 586.950 637.950 589.050 638.400 ;
        RECT 610.950 637.950 613.050 638.400 ;
        RECT 805.950 639.600 808.050 640.050 ;
        RECT 811.950 639.600 814.050 640.050 ;
        RECT 805.950 638.400 814.050 639.600 ;
        RECT 805.950 637.950 808.050 638.400 ;
        RECT 811.950 637.950 814.050 638.400 ;
        RECT 319.950 636.600 322.050 637.050 ;
        RECT 346.950 636.600 349.050 637.050 ;
        RECT 319.950 635.400 349.050 636.600 ;
        RECT 319.950 634.950 322.050 635.400 ;
        RECT 346.950 634.950 349.050 635.400 ;
        RECT 517.950 636.600 520.050 637.050 ;
        RECT 532.950 636.600 535.050 637.050 ;
        RECT 517.950 635.400 535.050 636.600 ;
        RECT 517.950 634.950 520.050 635.400 ;
        RECT 532.950 634.950 535.050 635.400 ;
        RECT 541.950 636.600 544.050 637.050 ;
        RECT 574.950 636.600 577.050 637.050 ;
        RECT 541.950 635.400 577.050 636.600 ;
        RECT 541.950 634.950 544.050 635.400 ;
        RECT 574.950 634.950 577.050 635.400 ;
        RECT 745.950 636.600 748.050 637.050 ;
        RECT 799.950 636.600 802.050 637.050 ;
        RECT 745.950 635.400 802.050 636.600 ;
        RECT 745.950 634.950 748.050 635.400 ;
        RECT 799.950 634.950 802.050 635.400 ;
        RECT 91.950 633.600 94.050 634.050 ;
        RECT 103.950 633.600 106.050 634.050 ;
        RECT 91.950 632.400 106.050 633.600 ;
        RECT 91.950 631.950 94.050 632.400 ;
        RECT 103.950 631.950 106.050 632.400 ;
        RECT 232.950 633.600 235.050 634.050 ;
        RECT 355.950 633.600 358.050 634.050 ;
        RECT 370.950 633.600 373.050 634.050 ;
        RECT 544.950 633.600 547.050 634.050 ;
        RECT 232.950 632.400 373.050 633.600 ;
        RECT 232.950 631.950 235.050 632.400 ;
        RECT 355.950 631.950 358.050 632.400 ;
        RECT 370.950 631.950 373.050 632.400 ;
        RECT 500.400 632.400 547.050 633.600 ;
        RECT 500.400 631.050 501.600 632.400 ;
        RECT 544.950 631.950 547.050 632.400 ;
        RECT 268.950 630.600 271.050 631.050 ;
        RECT 319.800 630.600 321.900 631.050 ;
        RECT 268.950 629.400 321.900 630.600 ;
        RECT 268.950 628.950 271.050 629.400 ;
        RECT 319.800 628.950 321.900 629.400 ;
        RECT 323.100 630.600 325.200 631.050 ;
        RECT 343.950 630.600 346.050 631.050 ;
        RECT 323.100 629.400 346.050 630.600 ;
        RECT 323.100 628.950 325.200 629.400 ;
        RECT 343.950 628.950 346.050 629.400 ;
        RECT 415.950 630.600 418.050 631.050 ;
        RECT 454.950 630.600 457.050 631.050 ;
        RECT 463.950 630.600 466.050 631.050 ;
        RECT 499.800 630.600 501.900 631.050 ;
        RECT 415.950 629.400 501.900 630.600 ;
        RECT 415.950 628.950 418.050 629.400 ;
        RECT 454.950 628.950 457.050 629.400 ;
        RECT 463.950 628.950 466.050 629.400 ;
        RECT 499.800 628.950 501.900 629.400 ;
        RECT 640.950 630.600 643.050 631.050 ;
        RECT 664.950 630.600 667.050 631.050 ;
        RECT 670.950 630.600 673.050 631.050 ;
        RECT 640.950 629.400 673.050 630.600 ;
        RECT 640.950 628.950 643.050 629.400 ;
        RECT 664.950 628.950 667.050 629.400 ;
        RECT 670.950 628.950 673.050 629.400 ;
        RECT 70.950 627.600 73.050 628.050 ;
        RECT 106.950 627.600 109.050 628.050 ;
        RECT 70.950 626.400 109.050 627.600 ;
        RECT 70.950 625.950 73.050 626.400 ;
        RECT 106.950 625.950 109.050 626.400 ;
        RECT 154.950 627.600 157.050 628.050 ;
        RECT 175.950 627.600 178.050 628.050 ;
        RECT 154.950 626.400 178.050 627.600 ;
        RECT 154.950 625.950 157.050 626.400 ;
        RECT 175.950 625.950 178.050 626.400 ;
        RECT 202.950 627.600 205.050 628.050 ;
        RECT 232.950 627.600 235.050 628.050 ;
        RECT 202.950 626.400 235.050 627.600 ;
        RECT 202.950 625.950 205.050 626.400 ;
        RECT 232.950 625.950 235.050 626.400 ;
        RECT 238.950 627.600 241.050 628.050 ;
        RECT 364.950 627.600 367.050 628.050 ;
        RECT 373.950 627.600 376.050 628.050 ;
        RECT 580.950 627.600 583.050 628.050 ;
        RECT 238.950 626.400 583.050 627.600 ;
        RECT 238.950 625.950 241.050 626.400 ;
        RECT 364.950 625.950 367.050 626.400 ;
        RECT 373.950 625.950 376.050 626.400 ;
        RECT 580.950 625.950 583.050 626.400 ;
        RECT 703.950 627.600 706.050 628.050 ;
        RECT 796.950 627.600 799.050 628.050 ;
        RECT 703.950 626.400 799.050 627.600 ;
        RECT 703.950 625.950 706.050 626.400 ;
        RECT 796.950 625.950 799.050 626.400 ;
        RECT 133.950 624.600 136.050 625.050 ;
        RECT 253.950 624.600 256.050 625.050 ;
        RECT 133.950 623.400 256.050 624.600 ;
        RECT 133.950 622.950 136.050 623.400 ;
        RECT 253.950 622.950 256.050 623.400 ;
        RECT 340.950 624.600 343.050 625.050 ;
        RECT 415.950 624.600 418.050 625.050 ;
        RECT 340.950 623.400 418.050 624.600 ;
        RECT 340.950 622.950 343.050 623.400 ;
        RECT 415.950 622.950 418.050 623.400 ;
        RECT 535.950 624.600 538.050 625.050 ;
        RECT 622.950 624.600 625.050 625.050 ;
        RECT 535.950 623.400 625.050 624.600 ;
        RECT 535.950 622.950 538.050 623.400 ;
        RECT 622.950 622.950 625.050 623.400 ;
        RECT 679.950 624.600 682.050 625.050 ;
        RECT 754.950 624.600 757.050 625.050 ;
        RECT 679.950 623.400 757.050 624.600 ;
        RECT 679.950 622.950 682.050 623.400 ;
        RECT 754.950 622.950 757.050 623.400 ;
        RECT 787.950 624.600 790.050 625.050 ;
        RECT 811.950 624.600 814.050 625.050 ;
        RECT 787.950 623.400 814.050 624.600 ;
        RECT 787.950 622.950 790.050 623.400 ;
        RECT 811.950 622.950 814.050 623.400 ;
        RECT 160.950 621.600 163.050 622.050 ;
        RECT 178.950 621.600 181.050 622.050 ;
        RECT 202.950 621.600 205.050 622.050 ;
        RECT 418.950 621.600 421.050 622.050 ;
        RECT 160.950 620.400 192.600 621.600 ;
        RECT 160.950 619.950 163.050 620.400 ;
        RECT 178.950 619.950 181.050 620.400 ;
        RECT 64.950 618.600 67.050 619.050 ;
        RECT 112.950 618.600 115.050 619.050 ;
        RECT 64.950 617.400 115.050 618.600 ;
        RECT 191.400 618.600 192.600 620.400 ;
        RECT 202.950 620.400 421.050 621.600 ;
        RECT 202.950 619.950 205.050 620.400 ;
        RECT 418.950 619.950 421.050 620.400 ;
        RECT 490.950 621.600 493.050 622.050 ;
        RECT 523.950 621.600 526.050 622.050 ;
        RECT 490.950 620.400 526.050 621.600 ;
        RECT 490.950 619.950 493.050 620.400 ;
        RECT 523.950 619.950 526.050 620.400 ;
        RECT 532.950 621.600 535.050 622.050 ;
        RECT 556.950 621.600 559.050 622.050 ;
        RECT 532.950 620.400 559.050 621.600 ;
        RECT 532.950 619.950 535.050 620.400 ;
        RECT 556.950 619.950 559.050 620.400 ;
        RECT 577.950 621.600 580.050 622.050 ;
        RECT 601.950 621.600 604.050 622.050 ;
        RECT 577.950 620.400 604.050 621.600 ;
        RECT 577.950 619.950 580.050 620.400 ;
        RECT 601.950 619.950 604.050 620.400 ;
        RECT 751.950 621.600 754.050 622.050 ;
        RECT 760.950 621.600 763.050 622.050 ;
        RECT 751.950 620.400 763.050 621.600 ;
        RECT 751.950 619.950 754.050 620.400 ;
        RECT 760.950 619.950 763.050 620.400 ;
        RECT 199.950 618.600 202.050 619.050 ;
        RECT 277.950 618.600 280.050 619.050 ;
        RECT 283.950 618.600 286.050 619.050 ;
        RECT 191.400 617.400 286.050 618.600 ;
        RECT 64.950 616.950 67.050 617.400 ;
        RECT 112.950 616.950 115.050 617.400 ;
        RECT 199.950 616.950 202.050 617.400 ;
        RECT 277.950 616.950 280.050 617.400 ;
        RECT 283.950 616.950 286.050 617.400 ;
        RECT 706.950 618.600 709.050 619.050 ;
        RECT 766.950 618.600 769.050 619.050 ;
        RECT 790.950 618.600 793.050 619.050 ;
        RECT 706.950 617.400 793.050 618.600 ;
        RECT 706.950 616.950 709.050 617.400 ;
        RECT 766.950 616.950 769.050 617.400 ;
        RECT 790.950 616.950 793.050 617.400 ;
        RECT 79.950 615.600 82.050 616.050 ;
        RECT 109.950 615.600 112.050 616.050 ;
        RECT 79.950 614.400 112.050 615.600 ;
        RECT 79.950 613.950 82.050 614.400 ;
        RECT 109.950 613.950 112.050 614.400 ;
        RECT 157.950 615.600 160.050 616.050 ;
        RECT 187.950 615.600 190.050 616.050 ;
        RECT 157.950 614.400 190.050 615.600 ;
        RECT 157.950 613.950 160.050 614.400 ;
        RECT 187.950 613.950 190.050 614.400 ;
        RECT 211.950 615.600 214.050 616.050 ;
        RECT 217.950 615.600 220.050 616.200 ;
        RECT 211.950 614.400 220.050 615.600 ;
        RECT 211.950 613.950 214.050 614.400 ;
        RECT 217.950 614.100 220.050 614.400 ;
        RECT 223.950 615.600 226.050 616.050 ;
        RECT 244.950 615.600 247.050 616.050 ;
        RECT 223.950 614.400 247.050 615.600 ;
        RECT 223.950 613.950 226.050 614.400 ;
        RECT 244.950 613.950 247.050 614.400 ;
        RECT 325.950 615.600 328.050 616.050 ;
        RECT 340.950 615.600 343.050 616.050 ;
        RECT 325.950 614.400 343.050 615.600 ;
        RECT 325.950 613.950 328.050 614.400 ;
        RECT 340.950 613.950 343.050 614.400 ;
        RECT 517.950 615.600 520.050 616.050 ;
        RECT 529.950 615.600 532.050 616.050 ;
        RECT 517.950 614.400 532.050 615.600 ;
        RECT 517.950 613.950 520.050 614.400 ;
        RECT 529.950 613.950 532.050 614.400 ;
        RECT 550.950 615.600 553.050 616.050 ;
        RECT 562.950 615.600 565.050 616.050 ;
        RECT 550.950 614.400 565.050 615.600 ;
        RECT 550.950 613.950 553.050 614.400 ;
        RECT 562.950 613.950 565.050 614.400 ;
        RECT 607.950 615.600 610.050 616.050 ;
        RECT 667.950 615.600 670.050 616.050 ;
        RECT 688.950 615.600 691.050 616.050 ;
        RECT 607.950 614.400 691.050 615.600 ;
        RECT 607.950 613.950 610.050 614.400 ;
        RECT 667.950 613.950 670.050 614.400 ;
        RECT 688.950 613.950 691.050 614.400 ;
        RECT 28.950 612.600 31.050 613.050 ;
        RECT 40.950 612.600 43.050 613.050 ;
        RECT 20.400 611.400 43.050 612.600 ;
        RECT 20.400 610.050 21.600 611.400 ;
        RECT 28.950 610.950 31.050 611.400 ;
        RECT 40.950 610.950 43.050 611.400 ;
        RECT 46.950 612.600 49.050 613.050 ;
        RECT 76.950 612.600 79.050 613.050 ;
        RECT 46.950 611.400 79.050 612.600 ;
        RECT 46.950 610.950 49.050 611.400 ;
        RECT 76.950 610.950 79.050 611.400 ;
        RECT 82.950 612.600 85.050 613.050 ;
        RECT 100.950 612.600 103.050 613.050 ;
        RECT 82.950 611.400 103.050 612.600 ;
        RECT 82.950 610.950 85.050 611.400 ;
        RECT 100.950 610.950 103.050 611.400 ;
        RECT 16.950 608.400 21.600 610.050 ;
        RECT 34.950 609.600 37.050 610.050 ;
        RECT 47.400 609.600 48.600 610.950 ;
        RECT 34.950 608.400 48.600 609.600 ;
        RECT 115.950 609.600 118.050 610.050 ;
        RECT 127.950 609.600 130.050 613.050 ;
        RECT 193.950 612.600 196.050 613.050 ;
        RECT 202.950 612.600 205.050 613.050 ;
        RECT 193.950 611.400 205.050 612.600 ;
        RECT 193.950 610.950 196.050 611.400 ;
        RECT 202.950 610.950 205.050 611.400 ;
        RECT 217.950 612.600 220.050 612.900 ;
        RECT 226.950 612.600 229.050 613.050 ;
        RECT 217.950 611.400 229.050 612.600 ;
        RECT 217.950 610.800 220.050 611.400 ;
        RECT 226.950 610.950 229.050 611.400 ;
        RECT 310.950 612.600 313.050 613.200 ;
        RECT 478.950 612.600 481.050 613.050 ;
        RECT 553.950 612.600 556.050 613.050 ;
        RECT 310.950 611.400 327.600 612.600 ;
        RECT 310.950 611.100 313.050 611.400 ;
        RECT 115.950 609.000 130.050 609.600 ;
        RECT 115.950 608.400 129.600 609.000 ;
        RECT 16.950 607.950 21.000 608.400 ;
        RECT 34.950 607.950 37.050 608.400 ;
        RECT 115.950 607.950 118.050 608.400 ;
        RECT 25.950 606.600 28.050 607.050 ;
        RECT 58.950 606.600 61.050 607.050 ;
        RECT 25.950 605.400 61.050 606.600 ;
        RECT 25.950 604.950 28.050 605.400 ;
        RECT 58.950 604.950 61.050 605.400 ;
        RECT 70.950 606.600 73.050 607.050 ;
        RECT 97.950 606.600 103.050 607.050 ;
        RECT 70.950 605.400 103.050 606.600 ;
        RECT 70.950 604.950 73.050 605.400 ;
        RECT 97.950 604.950 103.050 605.400 ;
        RECT 166.950 606.600 172.050 607.050 ;
        RECT 181.950 606.600 184.050 610.050 ;
        RECT 238.950 609.600 241.050 610.050 ;
        RECT 259.950 609.600 262.050 610.050 ;
        RECT 238.950 608.400 262.050 609.600 ;
        RECT 238.950 607.950 241.050 608.400 ;
        RECT 259.950 607.950 262.050 608.400 ;
        RECT 289.950 609.600 292.050 610.200 ;
        RECT 295.950 609.600 298.050 610.050 ;
        RECT 289.950 608.400 298.050 609.600 ;
        RECT 289.950 608.100 292.050 608.400 ;
        RECT 295.950 607.950 298.050 608.400 ;
        RECT 310.950 609.600 313.050 609.900 ;
        RECT 322.950 609.600 325.050 610.050 ;
        RECT 310.950 608.400 325.050 609.600 ;
        RECT 326.400 609.600 327.600 611.400 ;
        RECT 478.950 611.400 556.050 612.600 ;
        RECT 478.950 610.950 481.050 611.400 ;
        RECT 553.950 610.950 556.050 611.400 ;
        RECT 418.950 609.600 421.050 610.050 ;
        RECT 451.950 609.600 454.050 610.050 ;
        RECT 326.400 608.400 333.600 609.600 ;
        RECT 310.950 607.800 313.050 608.400 ;
        RECT 322.950 607.950 325.050 608.400 ;
        RECT 166.950 606.000 184.050 606.600 ;
        RECT 220.950 606.600 223.050 607.200 ;
        RECT 332.400 607.050 333.600 608.400 ;
        RECT 418.950 608.400 454.050 609.600 ;
        RECT 418.950 607.950 421.050 608.400 ;
        RECT 451.950 607.950 454.050 608.400 ;
        RECT 457.950 609.600 460.050 610.050 ;
        RECT 466.950 609.600 469.050 610.050 ;
        RECT 457.950 608.400 469.050 609.600 ;
        RECT 601.950 609.600 604.050 613.050 ;
        RECT 742.950 612.600 745.050 613.050 ;
        RECT 757.950 612.600 760.050 613.050 ;
        RECT 742.950 611.400 760.050 612.600 ;
        RECT 742.950 610.950 745.050 611.400 ;
        RECT 757.950 610.950 760.050 611.400 ;
        RECT 625.950 609.600 628.050 610.050 ;
        RECT 601.950 609.000 628.050 609.600 ;
        RECT 602.400 608.400 628.050 609.000 ;
        RECT 457.950 607.950 460.050 608.400 ;
        RECT 466.950 607.950 469.050 608.400 ;
        RECT 625.950 607.950 628.050 608.400 ;
        RECT 631.950 609.600 634.050 610.050 ;
        RECT 652.950 609.600 655.050 610.050 ;
        RECT 631.950 608.400 655.050 609.600 ;
        RECT 631.950 607.950 634.050 608.400 ;
        RECT 652.950 607.950 655.050 608.400 ;
        RECT 232.950 606.600 235.050 607.050 ;
        RECT 166.950 605.400 183.600 606.000 ;
        RECT 220.950 605.400 235.050 606.600 ;
        RECT 166.950 604.950 172.050 605.400 ;
        RECT 220.950 605.100 223.050 605.400 ;
        RECT 232.950 604.950 235.050 605.400 ;
        RECT 268.950 606.600 271.050 606.900 ;
        RECT 292.950 606.600 295.050 607.050 ;
        RECT 268.950 605.400 295.050 606.600 ;
        RECT 332.400 605.400 337.050 607.050 ;
        RECT 268.950 604.800 271.050 605.400 ;
        RECT 292.950 604.950 295.050 605.400 ;
        RECT 333.000 604.950 337.050 605.400 ;
        RECT 376.950 606.600 379.050 607.050 ;
        RECT 388.950 606.600 391.050 607.050 ;
        RECT 415.950 606.600 418.050 607.050 ;
        RECT 376.950 605.400 418.050 606.600 ;
        RECT 376.950 604.950 379.050 605.400 ;
        RECT 388.950 604.950 391.050 605.400 ;
        RECT 415.950 604.950 418.050 605.400 ;
        RECT 427.950 606.600 430.050 607.200 ;
        RECT 514.950 606.600 517.050 607.200 ;
        RECT 520.950 606.600 523.050 607.050 ;
        RECT 427.950 605.400 441.600 606.600 ;
        RECT 427.950 605.100 430.050 605.400 ;
        RECT 109.950 601.950 115.050 604.050 ;
        RECT 136.950 603.600 139.050 604.200 ;
        RECT 116.400 602.400 139.050 603.600 ;
        RECT 7.950 600.600 10.050 601.050 ;
        RECT 19.950 600.600 22.050 601.050 ;
        RECT 7.950 599.400 22.050 600.600 ;
        RECT 7.950 598.950 10.050 599.400 ;
        RECT 19.950 598.950 22.050 599.400 ;
        RECT 88.950 600.600 91.050 601.050 ;
        RECT 116.400 600.600 117.600 602.400 ;
        RECT 136.950 602.100 139.050 602.400 ;
        RECT 175.950 603.600 178.050 604.050 ;
        RECT 184.950 603.600 187.050 604.200 ;
        RECT 175.950 602.400 187.050 603.600 ;
        RECT 175.950 601.950 178.050 602.400 ;
        RECT 184.950 602.100 187.050 602.400 ;
        RECT 190.950 603.600 193.050 604.050 ;
        RECT 205.950 603.600 208.050 604.050 ;
        RECT 190.950 602.400 208.050 603.600 ;
        RECT 190.950 601.950 193.050 602.400 ;
        RECT 205.950 601.950 208.050 602.400 ;
        RECT 256.950 603.600 259.050 604.050 ;
        RECT 277.950 603.600 280.050 604.050 ;
        RECT 256.950 602.400 280.050 603.600 ;
        RECT 256.950 601.950 259.050 602.400 ;
        RECT 277.950 601.950 280.050 602.400 ;
        RECT 289.950 603.600 292.050 604.050 ;
        RECT 304.950 603.600 307.050 604.050 ;
        RECT 289.950 602.400 307.050 603.600 ;
        RECT 289.950 601.950 292.050 602.400 ;
        RECT 304.950 601.950 307.050 602.400 ;
        RECT 328.950 603.600 331.050 604.050 ;
        RECT 343.950 603.600 346.050 604.050 ;
        RECT 328.950 602.400 346.050 603.600 ;
        RECT 328.950 601.950 331.050 602.400 ;
        RECT 343.950 601.950 346.050 602.400 ;
        RECT 367.950 603.600 370.050 604.050 ;
        RECT 373.950 603.600 376.050 604.050 ;
        RECT 367.950 602.400 376.050 603.600 ;
        RECT 367.950 601.950 370.050 602.400 ;
        RECT 373.950 601.950 376.050 602.400 ;
        RECT 385.950 603.600 388.050 604.050 ;
        RECT 391.950 603.600 394.050 604.050 ;
        RECT 385.950 602.400 394.050 603.600 ;
        RECT 385.950 601.950 388.050 602.400 ;
        RECT 391.950 601.950 394.050 602.400 ;
        RECT 421.950 603.600 424.050 604.200 ;
        RECT 440.400 604.050 441.600 605.400 ;
        RECT 514.950 605.400 523.050 606.600 ;
        RECT 514.950 605.100 517.050 605.400 ;
        RECT 520.950 604.950 523.050 605.400 ;
        RECT 529.950 606.600 532.050 607.050 ;
        RECT 538.950 606.600 541.050 607.200 ;
        RECT 529.950 605.400 541.050 606.600 ;
        RECT 529.950 604.950 532.050 605.400 ;
        RECT 538.950 605.100 541.050 605.400 ;
        RECT 544.950 606.600 547.050 607.050 ;
        RECT 556.950 606.600 559.050 607.050 ;
        RECT 544.950 605.400 559.050 606.600 ;
        RECT 544.950 604.950 547.050 605.400 ;
        RECT 556.950 604.950 559.050 605.400 ;
        RECT 634.950 606.600 637.050 607.050 ;
        RECT 643.950 606.600 646.050 607.050 ;
        RECT 634.950 605.400 646.050 606.600 ;
        RECT 634.950 604.950 637.050 605.400 ;
        RECT 643.950 604.950 646.050 605.400 ;
        RECT 670.950 606.600 673.050 607.050 ;
        RECT 688.950 606.600 691.050 607.200 ;
        RECT 670.950 605.400 691.050 606.600 ;
        RECT 670.950 604.950 673.050 605.400 ;
        RECT 688.950 605.100 691.050 605.400 ;
        RECT 724.950 606.600 727.050 607.050 ;
        RECT 733.950 606.600 736.050 607.050 ;
        RECT 724.950 605.400 736.050 606.600 ;
        RECT 724.950 604.950 727.050 605.400 ;
        RECT 733.950 604.950 736.050 605.400 ;
        RECT 742.950 606.600 745.050 607.050 ;
        RECT 748.950 606.600 751.050 607.050 ;
        RECT 742.950 605.400 751.050 606.600 ;
        RECT 742.950 604.950 745.050 605.400 ;
        RECT 748.950 604.950 751.050 605.400 ;
        RECT 796.950 606.600 799.050 607.050 ;
        RECT 814.950 606.600 817.050 610.050 ;
        RECT 796.950 606.000 817.050 606.600 ;
        RECT 796.950 605.400 816.600 606.000 ;
        RECT 796.950 604.950 799.050 605.400 ;
        RECT 427.950 603.600 430.050 603.900 ;
        RECT 421.950 602.400 430.050 603.600 ;
        RECT 421.950 602.100 424.050 602.400 ;
        RECT 427.950 601.800 430.050 602.400 ;
        RECT 439.950 603.600 442.050 604.050 ;
        RECT 460.950 603.600 463.050 604.050 ;
        RECT 439.950 602.400 463.050 603.600 ;
        RECT 439.950 601.950 442.050 602.400 ;
        RECT 460.950 601.950 463.050 602.400 ;
        RECT 688.950 603.600 691.050 603.900 ;
        RECT 715.950 603.600 718.050 604.050 ;
        RECT 754.950 603.600 757.050 604.050 ;
        RECT 772.950 603.600 775.050 604.050 ;
        RECT 688.950 602.400 775.050 603.600 ;
        RECT 688.950 601.800 691.050 602.400 ;
        RECT 715.950 601.950 718.050 602.400 ;
        RECT 754.950 601.950 757.050 602.400 ;
        RECT 772.950 601.950 775.050 602.400 ;
        RECT 784.950 603.600 787.050 604.050 ;
        RECT 790.950 603.600 793.050 603.900 ;
        RECT 784.950 602.400 793.050 603.600 ;
        RECT 784.950 601.950 787.050 602.400 ;
        RECT 790.950 601.800 793.050 602.400 ;
        RECT 88.950 599.400 117.600 600.600 ;
        RECT 259.950 600.600 262.050 601.050 ;
        RECT 271.950 600.600 274.050 601.050 ;
        RECT 259.950 599.400 274.050 600.600 ;
        RECT 88.950 598.950 91.050 599.400 ;
        RECT 259.950 598.950 262.050 599.400 ;
        RECT 271.950 598.950 274.050 599.400 ;
        RECT 349.950 600.600 352.050 601.050 ;
        RECT 379.950 600.600 384.000 601.050 ;
        RECT 442.950 600.600 445.050 601.050 ;
        RECT 481.950 600.600 484.050 601.050 ;
        RECT 499.950 600.600 502.050 601.050 ;
        RECT 349.950 599.400 384.600 600.600 ;
        RECT 442.950 600.000 456.600 600.600 ;
        RECT 442.950 599.400 457.050 600.000 ;
        RECT 349.950 598.950 352.050 599.400 ;
        RECT 379.950 598.950 384.000 599.400 ;
        RECT 442.950 598.950 445.050 599.400 ;
        RECT 22.950 597.600 25.050 598.050 ;
        RECT 31.950 597.600 34.050 598.050 ;
        RECT 22.950 596.400 34.050 597.600 ;
        RECT 22.950 595.950 25.050 596.400 ;
        RECT 31.950 595.950 34.050 596.400 ;
        RECT 136.950 597.600 139.050 598.050 ;
        RECT 160.950 597.600 163.050 598.050 ;
        RECT 136.950 596.400 163.050 597.600 ;
        RECT 136.950 595.950 139.050 596.400 ;
        RECT 160.950 595.950 163.050 596.400 ;
        RECT 205.950 597.600 208.050 598.050 ;
        RECT 220.950 597.600 223.050 598.050 ;
        RECT 205.950 596.400 223.050 597.600 ;
        RECT 205.950 595.950 208.050 596.400 ;
        RECT 220.950 595.950 223.050 596.400 ;
        RECT 298.950 597.600 301.050 598.050 ;
        RECT 313.950 597.600 316.050 598.050 ;
        RECT 298.950 596.400 316.050 597.600 ;
        RECT 298.950 595.950 301.050 596.400 ;
        RECT 313.950 595.950 316.050 596.400 ;
        RECT 394.950 597.600 397.050 598.050 ;
        RECT 409.950 597.600 412.050 598.050 ;
        RECT 394.950 596.400 412.050 597.600 ;
        RECT 394.950 595.950 397.050 596.400 ;
        RECT 409.950 595.950 412.050 596.400 ;
        RECT 454.950 595.950 457.050 599.400 ;
        RECT 481.950 599.400 502.050 600.600 ;
        RECT 481.950 598.950 484.050 599.400 ;
        RECT 499.950 598.950 502.050 599.400 ;
        RECT 505.950 600.600 508.050 601.050 ;
        RECT 583.950 600.600 586.050 601.050 ;
        RECT 505.950 599.400 586.050 600.600 ;
        RECT 505.950 598.950 508.050 599.400 ;
        RECT 583.950 598.950 586.050 599.400 ;
        RECT 628.950 600.600 631.050 601.050 ;
        RECT 646.950 600.600 649.050 601.050 ;
        RECT 628.950 599.400 649.050 600.600 ;
        RECT 628.950 598.950 631.050 599.400 ;
        RECT 646.950 598.950 649.050 599.400 ;
        RECT 460.950 597.600 463.050 597.900 ;
        RECT 478.950 597.600 481.050 598.050 ;
        RECT 460.950 596.400 481.050 597.600 ;
        RECT 460.950 595.800 463.050 596.400 ;
        RECT 478.950 595.950 481.050 596.400 ;
        RECT 502.950 597.600 505.050 598.050 ;
        RECT 514.950 597.600 517.050 598.050 ;
        RECT 502.950 596.400 517.050 597.600 ;
        RECT 502.950 595.950 505.050 596.400 ;
        RECT 514.950 595.950 517.050 596.400 ;
        RECT 532.950 597.600 535.050 598.050 ;
        RECT 586.950 597.600 589.050 598.050 ;
        RECT 532.950 596.400 589.050 597.600 ;
        RECT 532.950 595.950 535.050 596.400 ;
        RECT 586.950 595.950 589.050 596.400 ;
        RECT 610.950 597.600 613.050 598.050 ;
        RECT 625.950 597.600 628.050 598.050 ;
        RECT 610.950 596.400 628.050 597.600 ;
        RECT 610.950 595.950 613.050 596.400 ;
        RECT 625.950 595.950 628.050 596.400 ;
        RECT 664.950 597.600 667.050 598.050 ;
        RECT 733.950 597.600 736.050 598.050 ;
        RECT 787.950 597.600 790.050 598.050 ;
        RECT 664.950 596.400 790.050 597.600 ;
        RECT 664.950 595.950 667.050 596.400 ;
        RECT 733.950 595.950 736.050 596.400 ;
        RECT 787.950 595.950 790.050 596.400 ;
        RECT 169.950 594.600 172.050 595.050 ;
        RECT 184.950 594.600 187.050 595.050 ;
        RECT 169.950 593.400 187.050 594.600 ;
        RECT 169.950 592.950 172.050 593.400 ;
        RECT 184.950 592.950 187.050 593.400 ;
        RECT 196.950 594.600 199.050 595.050 ;
        RECT 217.950 594.600 220.050 595.050 ;
        RECT 196.950 593.400 220.050 594.600 ;
        RECT 196.950 592.950 199.050 593.400 ;
        RECT 217.950 592.950 220.050 593.400 ;
        RECT 241.950 594.600 244.050 595.050 ;
        RECT 358.950 594.600 361.050 595.050 ;
        RECT 241.950 593.400 361.050 594.600 ;
        RECT 241.950 592.950 244.050 593.400 ;
        RECT 358.950 592.950 361.050 593.400 ;
        RECT 370.950 594.600 373.050 595.050 ;
        RECT 415.950 594.600 418.050 595.050 ;
        RECT 448.950 594.600 451.050 595.050 ;
        RECT 370.950 593.400 451.050 594.600 ;
        RECT 370.950 592.950 373.050 593.400 ;
        RECT 415.950 592.950 418.050 593.400 ;
        RECT 448.950 592.950 451.050 593.400 ;
        RECT 466.950 594.600 469.050 595.050 ;
        RECT 487.950 594.600 490.050 595.050 ;
        RECT 466.950 593.400 490.050 594.600 ;
        RECT 466.950 592.950 469.050 593.400 ;
        RECT 487.950 592.950 490.050 593.400 ;
        RECT 706.950 594.600 709.050 595.050 ;
        RECT 718.950 594.600 721.050 595.050 ;
        RECT 817.950 594.600 820.050 595.050 ;
        RECT 706.950 593.400 721.050 594.600 ;
        RECT 706.950 592.950 709.050 593.400 ;
        RECT 718.950 592.950 721.050 593.400 ;
        RECT 797.400 593.400 820.050 594.600 ;
        RECT 91.950 591.600 94.050 592.050 ;
        RECT 136.950 591.600 139.050 592.050 ;
        RECT 91.950 590.400 139.050 591.600 ;
        RECT 91.950 589.950 94.050 590.400 ;
        RECT 136.950 589.950 139.050 590.400 ;
        RECT 166.950 591.600 169.050 592.050 ;
        RECT 187.950 591.600 190.050 592.050 ;
        RECT 166.950 590.400 190.050 591.600 ;
        RECT 166.950 589.950 169.050 590.400 ;
        RECT 187.950 589.950 190.050 590.400 ;
        RECT 220.950 591.600 223.050 592.050 ;
        RECT 271.950 591.600 274.050 592.050 ;
        RECT 220.950 590.400 274.050 591.600 ;
        RECT 220.950 589.950 223.050 590.400 ;
        RECT 271.950 589.950 274.050 590.400 ;
        RECT 331.950 591.600 334.050 592.050 ;
        RECT 385.950 591.600 388.050 592.050 ;
        RECT 397.800 591.600 399.900 592.050 ;
        RECT 331.950 590.400 388.050 591.600 ;
        RECT 331.950 589.950 334.050 590.400 ;
        RECT 385.950 589.950 388.050 590.400 ;
        RECT 389.400 590.400 399.900 591.600 ;
        RECT 277.950 588.600 280.050 589.050 ;
        RECT 295.950 588.600 298.050 589.050 ;
        RECT 337.950 588.600 340.050 589.050 ;
        RECT 389.400 588.600 390.600 590.400 ;
        RECT 397.800 589.950 399.900 590.400 ;
        RECT 401.100 591.600 403.200 592.050 ;
        RECT 421.950 591.600 424.050 592.050 ;
        RECT 401.100 590.400 424.050 591.600 ;
        RECT 401.100 589.950 403.200 590.400 ;
        RECT 421.950 589.950 424.050 590.400 ;
        RECT 472.950 591.600 475.050 592.050 ;
        RECT 490.950 591.600 493.050 592.050 ;
        RECT 748.950 591.600 751.050 592.050 ;
        RECT 787.950 591.600 790.050 592.050 ;
        RECT 797.400 591.600 798.600 593.400 ;
        RECT 817.950 592.950 820.050 593.400 ;
        RECT 472.950 590.400 493.050 591.600 ;
        RECT 472.950 589.950 475.050 590.400 ;
        RECT 490.950 589.950 493.050 590.400 ;
        RECT 593.400 590.400 609.600 591.600 ;
        RECT 430.950 588.600 433.050 589.050 ;
        RECT 277.950 587.400 390.600 588.600 ;
        RECT 398.400 587.400 433.050 588.600 ;
        RECT 277.950 586.950 280.050 587.400 ;
        RECT 295.950 586.950 298.050 587.400 ;
        RECT 337.950 586.950 340.050 587.400 ;
        RECT 178.950 585.600 181.050 586.050 ;
        RECT 193.950 585.600 196.050 586.050 ;
        RECT 178.950 584.400 196.050 585.600 ;
        RECT 178.950 583.950 181.050 584.400 ;
        RECT 193.950 583.950 196.050 584.400 ;
        RECT 286.950 585.600 289.050 586.050 ;
        RECT 298.950 585.600 301.050 586.050 ;
        RECT 310.950 585.600 313.050 586.050 ;
        RECT 286.950 584.400 313.050 585.600 ;
        RECT 286.950 583.950 289.050 584.400 ;
        RECT 298.950 583.950 301.050 584.400 ;
        RECT 310.950 583.950 313.050 584.400 ;
        RECT 382.950 585.600 385.050 586.050 ;
        RECT 398.400 585.600 399.600 587.400 ;
        RECT 430.950 586.950 433.050 587.400 ;
        RECT 445.950 588.600 448.050 589.050 ;
        RECT 457.950 588.600 460.050 589.050 ;
        RECT 517.950 588.600 520.050 589.050 ;
        RECT 593.400 588.600 594.600 590.400 ;
        RECT 445.950 587.400 520.050 588.600 ;
        RECT 445.950 586.950 448.050 587.400 ;
        RECT 457.950 586.950 460.050 587.400 ;
        RECT 517.950 586.950 520.050 587.400 ;
        RECT 554.400 587.400 594.600 588.600 ;
        RECT 608.400 588.600 609.600 590.400 ;
        RECT 748.950 590.400 798.600 591.600 ;
        RECT 748.950 589.950 751.050 590.400 ;
        RECT 787.950 589.950 790.050 590.400 ;
        RECT 634.950 588.600 637.050 589.050 ;
        RECT 608.400 587.400 637.050 588.600 ;
        RECT 382.950 584.400 399.600 585.600 ;
        RECT 400.950 585.600 403.050 586.050 ;
        RECT 412.950 585.600 415.050 586.050 ;
        RECT 400.950 584.400 415.050 585.600 ;
        RECT 382.950 583.950 385.050 584.400 ;
        RECT 400.950 583.950 403.050 584.400 ;
        RECT 412.950 583.950 415.050 584.400 ;
        RECT 475.950 585.600 478.050 586.050 ;
        RECT 502.950 585.600 505.050 586.050 ;
        RECT 475.950 584.400 505.050 585.600 ;
        RECT 475.950 583.950 478.050 584.400 ;
        RECT 502.950 583.950 505.050 584.400 ;
        RECT 508.950 585.600 511.050 586.050 ;
        RECT 538.950 585.600 541.050 586.050 ;
        RECT 508.950 584.400 541.050 585.600 ;
        RECT 508.950 583.950 511.050 584.400 ;
        RECT 538.950 583.950 541.050 584.400 ;
        RECT 544.950 585.600 547.050 586.050 ;
        RECT 554.400 585.600 555.600 587.400 ;
        RECT 634.950 586.950 637.050 587.400 ;
        RECT 649.950 588.600 652.050 589.050 ;
        RECT 676.950 588.600 679.050 589.050 ;
        RECT 694.950 588.600 697.050 589.050 ;
        RECT 649.950 587.400 697.050 588.600 ;
        RECT 649.950 586.950 652.050 587.400 ;
        RECT 676.950 586.950 679.050 587.400 ;
        RECT 694.950 586.950 697.050 587.400 ;
        RECT 799.950 588.600 802.050 589.050 ;
        RECT 823.950 588.600 826.050 589.050 ;
        RECT 799.950 587.400 826.050 588.600 ;
        RECT 799.950 586.950 802.050 587.400 ;
        RECT 823.950 586.950 826.050 587.400 ;
        RECT 544.950 584.400 555.600 585.600 ;
        RECT 544.950 583.950 547.050 584.400 ;
        RECT 88.950 582.600 91.050 583.050 ;
        RECT 103.950 582.600 106.050 583.050 ;
        RECT 142.950 582.600 145.050 583.050 ;
        RECT 88.950 581.400 145.050 582.600 ;
        RECT 88.950 580.950 91.050 581.400 ;
        RECT 103.950 580.950 106.050 581.400 ;
        RECT 142.950 580.950 145.050 581.400 ;
        RECT 184.950 582.600 187.050 583.050 ;
        RECT 199.950 582.600 202.050 583.050 ;
        RECT 184.950 581.400 202.050 582.600 ;
        RECT 184.950 580.950 187.050 581.400 ;
        RECT 199.950 580.950 202.050 581.400 ;
        RECT 208.950 582.600 211.050 583.050 ;
        RECT 277.950 582.600 280.050 583.050 ;
        RECT 208.950 581.400 280.050 582.600 ;
        RECT 208.950 580.950 211.050 581.400 ;
        RECT 277.950 580.950 280.050 581.400 ;
        RECT 289.950 582.600 292.050 583.050 ;
        RECT 301.950 582.600 304.050 583.050 ;
        RECT 334.950 582.600 337.050 583.050 ;
        RECT 370.950 582.600 373.050 583.050 ;
        RECT 289.950 581.400 373.050 582.600 ;
        RECT 289.950 580.950 292.050 581.400 ;
        RECT 301.950 580.950 304.050 581.400 ;
        RECT 334.950 580.950 337.050 581.400 ;
        RECT 370.950 580.950 373.050 581.400 ;
        RECT 442.950 582.600 445.050 583.050 ;
        RECT 472.950 582.600 475.050 583.050 ;
        RECT 442.950 581.400 475.050 582.600 ;
        RECT 442.950 580.950 445.050 581.400 ;
        RECT 472.950 580.950 475.050 581.400 ;
        RECT 481.950 582.600 484.050 583.050 ;
        RECT 532.950 582.600 535.050 583.050 ;
        RECT 481.950 581.400 535.050 582.600 ;
        RECT 481.950 580.950 484.050 581.400 ;
        RECT 532.950 580.950 535.050 581.400 ;
        RECT 559.950 582.600 562.050 583.050 ;
        RECT 595.950 582.600 598.050 583.050 ;
        RECT 619.950 582.600 622.050 583.050 ;
        RECT 559.950 581.400 622.050 582.600 ;
        RECT 559.950 580.950 562.050 581.400 ;
        RECT 595.950 580.950 598.050 581.400 ;
        RECT 619.950 580.950 622.050 581.400 ;
        RECT 739.950 582.600 742.050 583.050 ;
        RECT 751.950 582.600 754.050 583.050 ;
        RECT 739.950 581.400 754.050 582.600 ;
        RECT 739.950 580.950 742.050 581.400 ;
        RECT 751.950 580.950 754.050 581.400 ;
        RECT 49.950 579.600 52.050 580.050 ;
        RECT 61.950 579.600 64.050 580.050 ;
        RECT 49.950 578.400 64.050 579.600 ;
        RECT 49.950 577.950 52.050 578.400 ;
        RECT 61.950 577.950 64.050 578.400 ;
        RECT 271.950 579.600 274.050 580.050 ;
        RECT 295.950 579.600 298.050 580.050 ;
        RECT 271.950 578.400 298.050 579.600 ;
        RECT 271.950 577.950 274.050 578.400 ;
        RECT 295.950 577.950 298.050 578.400 ;
        RECT 565.950 579.600 568.050 580.050 ;
        RECT 574.950 579.600 577.050 580.050 ;
        RECT 565.950 578.400 577.050 579.600 ;
        RECT 565.950 577.950 568.050 578.400 ;
        RECT 574.950 577.950 577.050 578.400 ;
        RECT 712.950 579.600 715.050 580.050 ;
        RECT 775.950 579.600 778.050 580.050 ;
        RECT 808.950 579.600 811.050 580.050 ;
        RECT 712.950 578.400 811.050 579.600 ;
        RECT 712.950 577.950 715.050 578.400 ;
        RECT 775.950 577.950 778.050 578.400 ;
        RECT 808.950 577.950 811.050 578.400 ;
        RECT 10.950 576.600 13.050 577.050 ;
        RECT 34.950 576.600 37.050 577.050 ;
        RECT 10.950 575.400 37.050 576.600 ;
        RECT 10.950 574.950 13.050 575.400 ;
        RECT 34.950 574.950 37.050 575.400 ;
        RECT 79.950 576.600 82.050 577.200 ;
        RECT 85.950 576.600 88.050 577.050 ;
        RECT 79.950 575.400 88.050 576.600 ;
        RECT 79.950 575.100 82.050 575.400 ;
        RECT 85.950 574.950 88.050 575.400 ;
        RECT 127.950 576.600 130.050 577.050 ;
        RECT 142.950 576.600 145.050 577.050 ;
        RECT 166.950 576.600 169.050 577.050 ;
        RECT 127.950 575.400 169.050 576.600 ;
        RECT 127.950 574.950 130.050 575.400 ;
        RECT 142.950 574.950 145.050 575.400 ;
        RECT 166.950 574.950 169.050 575.400 ;
        RECT 262.950 576.600 265.050 577.050 ;
        RECT 292.950 576.600 295.050 577.050 ;
        RECT 262.950 575.400 295.050 576.600 ;
        RECT 262.950 574.950 265.050 575.400 ;
        RECT 292.950 574.950 295.050 575.400 ;
        RECT 361.950 574.950 364.050 577.050 ;
        RECT 367.950 574.950 370.050 577.050 ;
        RECT 436.950 576.600 439.050 577.050 ;
        RECT 562.950 576.600 565.050 577.050 ;
        RECT 580.950 576.600 583.050 577.200 ;
        RECT 436.950 575.400 456.600 576.600 ;
        RECT 436.950 574.950 439.050 575.400 ;
        RECT 16.950 573.600 19.050 574.050 ;
        RECT 25.950 573.600 28.050 574.050 ;
        RECT 16.950 572.400 28.050 573.600 ;
        RECT 16.950 571.950 19.050 572.400 ;
        RECT 25.950 571.950 28.050 572.400 ;
        RECT 298.950 573.600 301.050 574.050 ;
        RECT 304.950 573.600 307.050 574.050 ;
        RECT 298.950 572.400 307.050 573.600 ;
        RECT 298.950 571.950 301.050 572.400 ;
        RECT 304.950 571.950 307.050 572.400 ;
        RECT 34.950 570.600 37.050 570.900 ;
        RECT 49.950 570.600 52.050 571.050 ;
        RECT 34.950 569.400 52.050 570.600 ;
        RECT 34.950 568.800 37.050 569.400 ;
        RECT 49.950 568.950 52.050 569.400 ;
        RECT 175.950 570.600 178.050 571.200 ;
        RECT 362.400 571.050 363.600 574.950 ;
        RECT 368.400 571.050 369.600 574.950 ;
        RECT 181.950 570.600 184.050 571.050 ;
        RECT 175.950 569.400 184.050 570.600 ;
        RECT 175.950 569.100 178.050 569.400 ;
        RECT 181.950 568.950 184.050 569.400 ;
        RECT 211.950 570.600 214.050 571.050 ;
        RECT 220.950 570.600 223.050 571.050 ;
        RECT 211.950 569.400 223.050 570.600 ;
        RECT 211.950 568.950 214.050 569.400 ;
        RECT 220.950 568.950 223.050 569.400 ;
        RECT 316.950 570.600 319.050 571.050 ;
        RECT 346.950 570.600 349.050 571.050 ;
        RECT 316.950 569.400 349.050 570.600 ;
        RECT 316.950 568.950 319.050 569.400 ;
        RECT 346.950 568.950 349.050 569.400 ;
        RECT 358.950 569.400 363.600 571.050 ;
        RECT 358.950 568.950 363.000 569.400 ;
        RECT 367.950 568.950 370.050 571.050 ;
        RECT 397.950 570.600 400.050 571.200 ;
        RECT 406.950 570.600 409.050 571.050 ;
        RECT 397.950 569.400 409.050 570.600 ;
        RECT 424.950 570.600 427.050 574.050 ;
        RECT 455.400 573.600 456.600 575.400 ;
        RECT 562.950 575.400 583.050 576.600 ;
        RECT 562.950 574.950 565.050 575.400 ;
        RECT 580.950 575.100 583.050 575.400 ;
        RECT 475.950 573.600 478.050 574.050 ;
        RECT 455.400 572.400 478.050 573.600 ;
        RECT 475.950 571.950 478.050 572.400 ;
        RECT 484.950 573.600 487.050 574.050 ;
        RECT 514.950 573.600 517.050 573.900 ;
        RECT 523.950 573.600 526.050 574.050 ;
        RECT 484.950 572.400 526.050 573.600 ;
        RECT 484.950 571.950 487.050 572.400 ;
        RECT 514.950 571.800 517.050 572.400 ;
        RECT 523.950 571.950 526.050 572.400 ;
        RECT 568.950 573.600 571.050 574.050 ;
        RECT 574.950 573.600 577.050 574.050 ;
        RECT 568.950 572.400 577.050 573.600 ;
        RECT 568.950 571.950 571.050 572.400 ;
        RECT 574.950 571.950 577.050 572.400 ;
        RECT 586.950 573.600 589.050 574.050 ;
        RECT 652.950 573.600 655.050 574.050 ;
        RECT 586.950 572.400 655.050 573.600 ;
        RECT 586.950 571.950 589.050 572.400 ;
        RECT 652.950 571.950 655.050 572.400 ;
        RECT 709.950 573.600 712.050 574.050 ;
        RECT 718.950 573.600 721.050 574.050 ;
        RECT 709.950 572.400 721.050 573.600 ;
        RECT 709.950 571.950 712.050 572.400 ;
        RECT 718.950 571.950 721.050 572.400 ;
        RECT 436.950 570.600 439.050 571.050 ;
        RECT 424.950 570.000 439.050 570.600 ;
        RECT 425.400 569.400 439.050 570.000 ;
        RECT 397.950 569.100 400.050 569.400 ;
        RECT 406.950 568.950 409.050 569.400 ;
        RECT 436.950 568.950 439.050 569.400 ;
        RECT 19.950 565.950 25.050 568.050 ;
        RECT 97.950 567.600 100.050 568.200 ;
        RECT 109.950 567.600 112.050 568.050 ;
        RECT 97.950 566.400 112.050 567.600 ;
        RECT 97.950 566.100 100.050 566.400 ;
        RECT 109.950 565.950 112.050 566.400 ;
        RECT 124.950 567.600 127.050 568.050 ;
        RECT 145.950 567.600 148.050 568.050 ;
        RECT 124.950 566.400 148.050 567.600 ;
        RECT 124.950 565.950 127.050 566.400 ;
        RECT 31.950 564.600 34.050 565.050 ;
        RECT 52.950 564.600 55.050 565.050 ;
        RECT 70.950 564.600 73.050 565.050 ;
        RECT 31.950 563.400 73.050 564.600 ;
        RECT 31.950 562.950 34.050 563.400 ;
        RECT 52.950 562.950 55.050 563.400 ;
        RECT 70.950 562.950 73.050 563.400 ;
        RECT 137.400 562.050 138.600 566.400 ;
        RECT 145.950 565.950 148.050 566.400 ;
        RECT 217.950 567.600 220.050 568.050 ;
        RECT 223.950 567.600 226.050 568.050 ;
        RECT 217.950 566.400 226.050 567.600 ;
        RECT 217.950 565.950 220.050 566.400 ;
        RECT 223.950 565.950 226.050 566.400 ;
        RECT 235.950 567.600 238.050 568.050 ;
        RECT 277.950 567.600 280.050 568.050 ;
        RECT 352.950 567.600 355.050 568.200 ;
        RECT 235.950 567.000 264.600 567.600 ;
        RECT 235.950 566.400 265.050 567.000 ;
        RECT 235.950 565.950 238.050 566.400 ;
        RECT 262.950 562.800 265.050 566.400 ;
        RECT 277.950 566.400 355.050 567.600 ;
        RECT 277.950 565.950 280.050 566.400 ;
        RECT 352.950 566.100 355.050 566.400 ;
        RECT 382.950 567.600 385.050 568.050 ;
        RECT 397.950 567.600 400.050 567.900 ;
        RECT 382.950 566.400 400.050 567.600 ;
        RECT 407.400 567.600 408.600 568.950 ;
        RECT 442.950 567.600 445.050 571.050 ;
        RECT 571.950 570.600 574.050 571.050 ;
        RECT 615.000 570.600 619.050 571.050 ;
        RECT 628.950 570.600 631.050 571.050 ;
        RECT 643.950 570.600 646.050 571.050 ;
        RECT 571.950 569.400 591.600 570.600 ;
        RECT 614.400 569.400 646.050 570.600 ;
        RECT 781.950 570.600 784.050 574.050 ;
        RECT 796.950 573.600 799.050 574.050 ;
        RECT 802.950 573.600 805.050 574.050 ;
        RECT 796.950 572.400 805.050 573.600 ;
        RECT 796.950 571.950 799.050 572.400 ;
        RECT 802.950 571.950 805.050 572.400 ;
        RECT 823.950 573.600 826.050 574.050 ;
        RECT 829.950 573.600 832.050 574.050 ;
        RECT 823.950 572.400 832.050 573.600 ;
        RECT 823.950 571.950 826.050 572.400 ;
        RECT 829.950 571.950 832.050 572.400 ;
        RECT 790.950 570.600 793.050 571.200 ;
        RECT 781.950 570.000 793.050 570.600 ;
        RECT 782.400 569.400 793.050 570.000 ;
        RECT 571.950 568.950 574.050 569.400 ;
        RECT 407.400 567.000 445.050 567.600 ;
        RECT 499.950 567.600 502.050 568.050 ;
        RECT 526.950 567.600 529.050 568.050 ;
        RECT 538.950 567.600 541.050 568.200 ;
        RECT 590.400 568.050 591.600 569.400 ;
        RECT 615.000 568.950 619.050 569.400 ;
        RECT 628.950 568.950 631.050 569.400 ;
        RECT 643.950 568.950 646.050 569.400 ;
        RECT 790.950 569.100 793.050 569.400 ;
        RECT 407.400 566.400 444.600 567.000 ;
        RECT 499.950 566.400 516.600 567.600 ;
        RECT 382.950 565.950 385.050 566.400 ;
        RECT 397.950 565.800 400.050 566.400 ;
        RECT 499.950 565.950 502.050 566.400 ;
        RECT 343.950 564.600 346.050 565.050 ;
        RECT 361.950 564.600 364.050 565.050 ;
        RECT 343.950 563.400 364.050 564.600 ;
        RECT 343.950 562.950 346.050 563.400 ;
        RECT 361.950 562.950 364.050 563.400 ;
        RECT 415.950 564.600 418.050 565.050 ;
        RECT 508.950 564.600 511.050 565.050 ;
        RECT 415.950 563.400 511.050 564.600 ;
        RECT 515.400 564.600 516.600 566.400 ;
        RECT 526.950 566.400 541.050 567.600 ;
        RECT 526.950 565.950 529.050 566.400 ;
        RECT 538.950 566.100 541.050 566.400 ;
        RECT 589.950 567.600 592.050 568.050 ;
        RECT 598.950 567.600 601.050 568.050 ;
        RECT 589.950 566.400 601.050 567.600 ;
        RECT 589.950 565.950 592.050 566.400 ;
        RECT 598.950 565.950 601.050 566.400 ;
        RECT 625.950 567.600 628.050 568.050 ;
        RECT 706.950 567.600 709.050 568.050 ;
        RECT 712.950 567.600 715.050 568.050 ;
        RECT 625.950 567.000 666.600 567.600 ;
        RECT 625.950 566.400 667.050 567.000 ;
        RECT 625.950 565.950 628.050 566.400 ;
        RECT 529.950 564.600 532.050 565.050 ;
        RECT 538.950 564.600 541.050 564.900 ;
        RECT 515.400 563.400 541.050 564.600 ;
        RECT 415.950 562.950 418.050 563.400 ;
        RECT 508.950 562.950 511.050 563.400 ;
        RECT 529.950 562.950 532.050 563.400 ;
        RECT 538.950 562.800 541.050 563.400 ;
        RECT 592.950 564.600 595.050 565.050 ;
        RECT 622.950 564.600 625.050 565.050 ;
        RECT 592.950 563.400 625.050 564.600 ;
        RECT 592.950 562.950 595.050 563.400 ;
        RECT 622.950 562.950 625.050 563.400 ;
        RECT 664.950 562.950 667.050 566.400 ;
        RECT 706.950 566.400 715.050 567.600 ;
        RECT 706.950 565.950 709.050 566.400 ;
        RECT 712.950 565.950 715.050 566.400 ;
        RECT 718.950 567.600 721.050 568.050 ;
        RECT 727.950 567.600 730.050 568.050 ;
        RECT 718.950 566.400 730.050 567.600 ;
        RECT 718.950 565.950 721.050 566.400 ;
        RECT 727.950 565.950 730.050 566.400 ;
        RECT 736.950 567.600 739.050 568.050 ;
        RECT 793.950 567.600 796.050 567.900 ;
        RECT 814.950 567.600 817.050 568.050 ;
        RECT 736.950 566.400 817.050 567.600 ;
        RECT 736.950 565.950 739.050 566.400 ;
        RECT 793.950 565.800 796.050 566.400 ;
        RECT 814.950 565.950 817.050 566.400 ;
        RECT 82.950 561.600 85.050 562.050 ;
        RECT 100.950 561.600 103.050 562.050 ;
        RECT 106.950 561.600 109.050 562.050 ;
        RECT 82.950 560.400 109.050 561.600 ;
        RECT 82.950 559.950 85.050 560.400 ;
        RECT 100.950 559.950 103.050 560.400 ;
        RECT 106.950 559.950 109.050 560.400 ;
        RECT 136.950 559.950 139.050 562.050 ;
        RECT 169.950 561.600 172.050 562.050 ;
        RECT 184.950 561.600 187.050 562.050 ;
        RECT 169.950 560.400 187.050 561.600 ;
        RECT 169.950 559.950 172.050 560.400 ;
        RECT 184.950 559.950 187.050 560.400 ;
        RECT 199.950 561.600 202.050 562.050 ;
        RECT 226.950 561.600 229.050 562.050 ;
        RECT 199.950 560.400 229.050 561.600 ;
        RECT 199.950 559.950 202.050 560.400 ;
        RECT 226.950 559.950 229.050 560.400 ;
        RECT 235.950 561.600 238.050 562.050 ;
        RECT 298.950 561.600 301.050 562.050 ;
        RECT 235.950 560.400 301.050 561.600 ;
        RECT 235.950 559.950 238.050 560.400 ;
        RECT 298.950 559.950 301.050 560.400 ;
        RECT 352.950 561.600 355.050 562.050 ;
        RECT 370.950 561.600 373.050 562.050 ;
        RECT 352.950 560.400 373.050 561.600 ;
        RECT 352.950 559.950 355.050 560.400 ;
        RECT 370.950 559.950 373.050 560.400 ;
        RECT 424.950 561.600 427.050 562.050 ;
        RECT 478.950 561.600 481.050 562.050 ;
        RECT 424.950 560.400 481.050 561.600 ;
        RECT 424.950 559.950 427.050 560.400 ;
        RECT 478.950 559.950 481.050 560.400 ;
        RECT 568.950 561.600 571.050 562.050 ;
        RECT 574.950 561.600 577.050 562.050 ;
        RECT 568.950 560.400 577.050 561.600 ;
        RECT 568.950 559.950 571.050 560.400 ;
        RECT 574.950 559.950 577.050 560.400 ;
        RECT 580.950 561.600 583.050 562.050 ;
        RECT 634.950 561.600 637.050 562.050 ;
        RECT 580.950 560.400 637.050 561.600 ;
        RECT 580.950 559.950 583.050 560.400 ;
        RECT 634.950 559.950 637.050 560.400 ;
        RECT 28.950 558.600 31.050 559.050 ;
        RECT 46.950 558.600 49.050 559.050 ;
        RECT 28.950 557.400 49.050 558.600 ;
        RECT 28.950 556.950 31.050 557.400 ;
        RECT 46.950 556.950 49.050 557.400 ;
        RECT 190.950 558.600 193.050 559.050 ;
        RECT 247.950 558.600 250.050 559.050 ;
        RECT 190.950 557.400 250.050 558.600 ;
        RECT 190.950 556.950 193.050 557.400 ;
        RECT 247.950 556.950 250.050 557.400 ;
        RECT 350.100 558.600 352.200 559.050 ;
        RECT 367.950 558.600 370.050 559.050 ;
        RECT 350.100 557.400 370.050 558.600 ;
        RECT 350.100 556.950 352.200 557.400 ;
        RECT 367.950 556.950 370.050 557.400 ;
        RECT 508.950 558.600 511.050 559.050 ;
        RECT 553.950 558.600 556.050 559.050 ;
        RECT 559.950 558.600 562.050 559.050 ;
        RECT 508.950 557.400 562.050 558.600 ;
        RECT 508.950 556.950 511.050 557.400 ;
        RECT 553.950 556.950 556.050 557.400 ;
        RECT 559.950 556.950 562.050 557.400 ;
        RECT 565.950 558.600 568.050 559.050 ;
        RECT 628.950 558.600 631.050 559.050 ;
        RECT 565.950 557.400 631.050 558.600 ;
        RECT 565.950 556.950 568.050 557.400 ;
        RECT 628.950 556.950 631.050 557.400 ;
        RECT 664.950 558.600 667.050 559.050 ;
        RECT 691.800 558.600 693.900 559.050 ;
        RECT 664.950 557.400 693.900 558.600 ;
        RECT 664.950 556.950 667.050 557.400 ;
        RECT 691.800 556.950 693.900 557.400 ;
        RECT 695.100 558.600 697.200 559.050 ;
        RECT 784.950 558.600 787.050 559.050 ;
        RECT 695.100 557.400 787.050 558.600 ;
        RECT 695.100 556.950 697.200 557.400 ;
        RECT 784.950 556.950 787.050 557.400 ;
        RECT 64.950 555.600 67.050 556.050 ;
        RECT 184.950 555.600 187.050 556.050 ;
        RECT 64.950 554.400 187.050 555.600 ;
        RECT 64.950 553.950 67.050 554.400 ;
        RECT 184.950 553.950 187.050 554.400 ;
        RECT 196.950 555.600 199.050 556.050 ;
        RECT 235.950 555.600 238.050 556.050 ;
        RECT 388.950 555.600 391.050 556.050 ;
        RECT 196.950 554.400 238.050 555.600 ;
        RECT 196.950 553.950 199.050 554.400 ;
        RECT 235.950 553.950 238.050 554.400 ;
        RECT 305.400 554.400 391.050 555.600 ;
        RECT 67.950 552.600 70.050 553.050 ;
        RECT 197.400 552.600 198.600 553.950 ;
        RECT 67.950 551.400 198.600 552.600 ;
        RECT 253.950 552.600 256.050 553.050 ;
        RECT 265.950 552.600 268.050 553.050 ;
        RECT 305.400 552.600 306.600 554.400 ;
        RECT 388.950 553.950 391.050 554.400 ;
        RECT 253.950 551.400 306.600 552.600 ;
        RECT 478.950 552.600 481.050 553.050 ;
        RECT 556.950 552.600 559.050 553.050 ;
        RECT 610.950 552.600 613.050 553.050 ;
        RECT 478.950 551.400 613.050 552.600 ;
        RECT 67.950 550.950 70.050 551.400 ;
        RECT 253.950 550.950 256.050 551.400 ;
        RECT 265.950 550.950 268.050 551.400 ;
        RECT 478.950 550.950 481.050 551.400 ;
        RECT 556.950 550.950 559.050 551.400 ;
        RECT 610.950 550.950 613.050 551.400 ;
        RECT 640.950 552.600 643.050 553.050 ;
        RECT 679.950 552.600 682.050 553.050 ;
        RECT 640.950 551.400 682.050 552.600 ;
        RECT 640.950 550.950 643.050 551.400 ;
        RECT 679.950 550.950 682.050 551.400 ;
        RECT 745.950 552.600 748.050 553.050 ;
        RECT 766.950 552.600 769.050 553.050 ;
        RECT 745.950 551.400 769.050 552.600 ;
        RECT 745.950 550.950 748.050 551.400 ;
        RECT 766.950 550.950 769.050 551.400 ;
        RECT 10.950 549.600 13.050 550.050 ;
        RECT 70.950 549.600 73.050 550.050 ;
        RECT 10.950 548.400 73.050 549.600 ;
        RECT 10.950 547.950 13.050 548.400 ;
        RECT 70.950 547.950 73.050 548.400 ;
        RECT 194.100 549.600 196.200 550.050 ;
        RECT 205.950 549.600 208.050 550.050 ;
        RECT 313.950 549.600 316.050 550.200 ;
        RECT 376.950 549.600 379.050 550.050 ;
        RECT 194.100 548.400 379.050 549.600 ;
        RECT 194.100 547.950 196.200 548.400 ;
        RECT 205.950 547.950 208.050 548.400 ;
        RECT 313.950 548.100 316.050 548.400 ;
        RECT 376.950 547.950 379.050 548.400 ;
        RECT 433.950 549.600 436.050 550.050 ;
        RECT 523.950 549.600 526.050 550.050 ;
        RECT 574.950 549.600 577.050 550.050 ;
        RECT 433.950 548.400 577.050 549.600 ;
        RECT 433.950 547.950 436.050 548.400 ;
        RECT 523.950 547.950 526.050 548.400 ;
        RECT 574.950 547.950 577.050 548.400 ;
        RECT 604.950 549.600 607.050 550.050 ;
        RECT 724.950 549.600 727.050 550.050 ;
        RECT 604.950 548.400 727.050 549.600 ;
        RECT 604.950 547.950 607.050 548.400 ;
        RECT 724.950 547.950 727.050 548.400 ;
        RECT 55.950 546.600 58.050 547.050 ;
        RECT 67.950 546.600 70.050 547.050 ;
        RECT 55.950 545.400 70.050 546.600 ;
        RECT 55.950 544.950 58.050 545.400 ;
        RECT 67.950 544.950 70.050 545.400 ;
        RECT 109.950 546.600 112.050 547.050 ;
        RECT 139.950 546.600 142.050 547.050 ;
        RECT 166.950 546.600 169.050 547.050 ;
        RECT 109.950 545.400 169.050 546.600 ;
        RECT 109.950 544.950 112.050 545.400 ;
        RECT 139.950 544.950 142.050 545.400 ;
        RECT 166.950 544.950 169.050 545.400 ;
        RECT 196.950 546.600 199.050 547.050 ;
        RECT 265.950 546.600 268.050 547.050 ;
        RECT 196.950 545.400 268.050 546.600 ;
        RECT 196.950 544.950 199.050 545.400 ;
        RECT 265.950 544.950 268.050 545.400 ;
        RECT 292.950 546.600 295.050 547.050 ;
        RECT 313.950 546.600 316.050 546.900 ;
        RECT 292.950 545.400 316.050 546.600 ;
        RECT 292.950 544.950 295.050 545.400 ;
        RECT 313.950 544.800 316.050 545.400 ;
        RECT 589.950 546.600 592.050 547.050 ;
        RECT 670.950 546.600 673.050 547.050 ;
        RECT 589.950 545.400 673.050 546.600 ;
        RECT 589.950 544.950 592.050 545.400 ;
        RECT 670.950 544.950 673.050 545.400 ;
        RECT 736.950 546.600 739.050 547.050 ;
        RECT 748.950 546.600 751.050 547.050 ;
        RECT 736.950 545.400 751.050 546.600 ;
        RECT 736.950 544.950 739.050 545.400 ;
        RECT 748.950 544.950 751.050 545.400 ;
        RECT 583.950 543.600 586.050 544.050 ;
        RECT 658.950 543.600 661.050 544.050 ;
        RECT 583.950 542.400 661.050 543.600 ;
        RECT 583.950 541.950 586.050 542.400 ;
        RECT 658.950 541.950 661.050 542.400 ;
        RECT 751.950 543.600 754.050 544.050 ;
        RECT 763.950 543.600 766.050 544.050 ;
        RECT 751.950 542.400 766.050 543.600 ;
        RECT 751.950 541.950 754.050 542.400 ;
        RECT 763.950 541.950 766.050 542.400 ;
        RECT 46.950 540.600 49.050 541.050 ;
        RECT 55.950 540.600 58.050 541.050 ;
        RECT 46.950 539.400 58.050 540.600 ;
        RECT 46.950 538.950 49.050 539.400 ;
        RECT 55.950 538.950 58.050 539.400 ;
        RECT 166.950 540.600 169.050 541.050 ;
        RECT 178.950 540.600 181.050 541.050 ;
        RECT 187.950 540.600 190.050 541.050 ;
        RECT 166.950 539.400 177.600 540.600 ;
        RECT 166.950 538.950 169.050 539.400 ;
        RECT 133.950 537.600 136.050 538.050 ;
        RECT 169.950 537.600 172.050 538.050 ;
        RECT 133.950 536.400 172.050 537.600 ;
        RECT 176.400 537.600 177.600 539.400 ;
        RECT 178.950 539.400 190.050 540.600 ;
        RECT 178.950 538.950 181.050 539.400 ;
        RECT 187.950 538.950 190.050 539.400 ;
        RECT 259.950 540.600 262.050 541.050 ;
        RECT 298.950 540.600 301.050 541.050 ;
        RECT 259.950 539.400 301.050 540.600 ;
        RECT 259.950 538.950 262.050 539.400 ;
        RECT 298.950 538.950 301.050 539.400 ;
        RECT 307.950 540.600 310.050 541.050 ;
        RECT 319.950 540.600 322.050 541.050 ;
        RECT 340.950 540.600 343.050 541.050 ;
        RECT 307.950 539.400 343.050 540.600 ;
        RECT 307.950 538.950 310.050 539.400 ;
        RECT 319.950 538.950 322.050 539.400 ;
        RECT 340.950 538.950 343.050 539.400 ;
        RECT 499.950 540.600 502.050 541.050 ;
        RECT 586.950 540.600 589.050 541.050 ;
        RECT 625.950 540.600 628.050 541.050 ;
        RECT 499.950 539.400 510.600 540.600 ;
        RECT 499.950 538.950 502.050 539.400 ;
        RECT 196.950 537.600 199.050 538.200 ;
        RECT 176.400 536.400 199.050 537.600 ;
        RECT 133.950 535.950 136.050 536.400 ;
        RECT 169.950 535.950 172.050 536.400 ;
        RECT 196.950 536.100 199.050 536.400 ;
        RECT 220.950 537.600 223.050 538.050 ;
        RECT 235.950 537.600 238.050 538.050 ;
        RECT 220.950 536.400 238.050 537.600 ;
        RECT 220.950 535.950 223.050 536.400 ;
        RECT 235.950 535.950 238.050 536.400 ;
        RECT 301.950 537.600 304.050 538.200 ;
        RECT 352.950 537.600 355.050 538.050 ;
        RECT 301.950 536.400 355.050 537.600 ;
        RECT 509.400 537.600 510.600 539.400 ;
        RECT 586.950 539.400 628.050 540.600 ;
        RECT 586.950 538.950 589.050 539.400 ;
        RECT 625.950 538.950 628.050 539.400 ;
        RECT 724.950 540.600 727.050 541.050 ;
        RECT 742.950 540.600 745.050 541.050 ;
        RECT 724.950 539.400 745.050 540.600 ;
        RECT 724.950 538.950 727.050 539.400 ;
        RECT 742.950 538.950 745.050 539.400 ;
        RECT 547.950 537.600 550.050 538.050 ;
        RECT 509.400 536.400 550.050 537.600 ;
        RECT 301.950 536.100 304.050 536.400 ;
        RECT 352.950 535.950 355.050 536.400 ;
        RECT 547.950 535.950 550.050 536.400 ;
        RECT 565.950 537.600 568.050 538.200 ;
        RECT 571.950 537.600 574.050 538.050 ;
        RECT 565.950 536.400 574.050 537.600 ;
        RECT 565.950 536.100 568.050 536.400 ;
        RECT 571.950 535.950 574.050 536.400 ;
        RECT 637.950 537.600 640.050 538.050 ;
        RECT 670.950 537.600 673.050 538.050 ;
        RECT 682.950 537.600 685.050 538.050 ;
        RECT 637.950 536.400 685.050 537.600 ;
        RECT 637.950 535.950 640.050 536.400 ;
        RECT 670.950 535.950 673.050 536.400 ;
        RECT 682.950 535.950 685.050 536.400 ;
        RECT 751.950 537.600 754.050 538.050 ;
        RECT 757.950 537.600 760.050 538.050 ;
        RECT 751.950 536.400 760.050 537.600 ;
        RECT 751.950 535.950 754.050 536.400 ;
        RECT 757.950 535.950 760.050 536.400 ;
        RECT 13.950 534.600 16.050 535.050 ;
        RECT 31.950 534.600 34.050 535.200 ;
        RECT 46.950 534.600 49.050 535.050 ;
        RECT 13.950 533.400 49.050 534.600 ;
        RECT 13.950 532.950 16.050 533.400 ;
        RECT 31.950 533.100 34.050 533.400 ;
        RECT 46.950 532.950 49.050 533.400 ;
        RECT 31.950 531.600 34.050 531.900 ;
        RECT 88.950 531.600 91.050 532.050 ;
        RECT 17.250 530.400 91.050 531.600 ;
        RECT 17.250 526.050 18.450 530.400 ;
        RECT 31.950 529.800 34.050 530.400 ;
        RECT 61.950 528.600 64.050 529.050 ;
        RECT 50.400 528.000 64.050 528.600 ;
        RECT 88.950 528.600 91.050 530.400 ;
        RECT 115.950 531.600 118.050 532.200 ;
        RECT 142.950 531.600 145.050 535.050 ;
        RECT 181.950 534.600 184.050 535.050 ;
        RECT 196.950 534.600 199.050 534.900 ;
        RECT 181.950 533.400 199.050 534.600 ;
        RECT 181.950 532.950 184.050 533.400 ;
        RECT 196.950 532.800 199.050 533.400 ;
        RECT 268.950 534.600 271.050 535.050 ;
        RECT 295.950 534.600 298.050 535.050 ;
        RECT 301.950 534.600 304.050 534.900 ;
        RECT 268.950 533.400 304.050 534.600 ;
        RECT 268.950 532.950 271.050 533.400 ;
        RECT 295.950 532.950 298.050 533.400 ;
        RECT 301.950 532.800 304.050 533.400 ;
        RECT 316.950 534.600 319.050 535.050 ;
        RECT 322.950 534.600 325.050 535.050 ;
        RECT 316.950 533.400 325.050 534.600 ;
        RECT 316.950 532.950 319.050 533.400 ;
        RECT 322.950 532.950 325.050 533.400 ;
        RECT 409.950 534.600 412.050 535.050 ;
        RECT 481.950 534.600 484.050 535.050 ;
        RECT 502.950 534.600 505.050 535.050 ;
        RECT 409.950 533.400 505.050 534.600 ;
        RECT 409.950 532.950 412.050 533.400 ;
        RECT 481.950 532.950 484.050 533.400 ;
        RECT 502.950 532.950 505.050 533.400 ;
        RECT 565.950 534.600 568.050 534.900 ;
        RECT 589.950 534.600 592.050 535.050 ;
        RECT 565.950 533.400 592.050 534.600 ;
        RECT 565.950 532.800 568.050 533.400 ;
        RECT 589.950 532.950 592.050 533.400 ;
        RECT 739.950 534.600 742.050 535.050 ;
        RECT 748.950 534.600 751.050 535.050 ;
        RECT 739.950 533.400 751.050 534.600 ;
        RECT 739.950 532.950 742.050 533.400 ;
        RECT 748.950 532.950 751.050 533.400 ;
        RECT 775.950 534.600 778.050 535.050 ;
        RECT 802.950 534.600 805.050 535.050 ;
        RECT 775.950 533.400 805.050 534.600 ;
        RECT 775.950 532.950 778.050 533.400 ;
        RECT 802.950 532.950 805.050 533.400 ;
        RECT 823.950 534.600 826.050 535.050 ;
        RECT 829.950 534.600 832.050 535.050 ;
        RECT 823.950 533.400 832.050 534.600 ;
        RECT 823.950 532.950 826.050 533.400 ;
        RECT 829.950 532.950 832.050 533.400 ;
        RECT 115.950 530.400 177.600 531.600 ;
        RECT 115.950 530.100 118.050 530.400 ;
        RECT 176.400 529.050 177.600 530.400 ;
        RECT 97.950 528.600 100.050 529.050 ;
        RECT 151.950 528.600 154.050 529.050 ;
        RECT 88.950 528.000 100.050 528.600 ;
        RECT 122.400 528.000 154.050 528.600 ;
        RECT 49.950 527.400 64.050 528.000 ;
        RECT 89.400 527.400 100.050 528.000 ;
        RECT 49.950 526.050 52.050 527.400 ;
        RECT 61.950 526.950 64.050 527.400 ;
        RECT 97.950 526.950 100.050 527.400 ;
        RECT 121.950 527.400 154.050 528.000 ;
        RECT 176.400 527.400 181.050 529.050 ;
        RECT 16.800 523.950 18.900 526.050 ;
        RECT 20.100 525.600 22.200 526.050 ;
        RECT 31.950 525.600 34.050 525.900 ;
        RECT 20.100 524.400 34.050 525.600 ;
        RECT 20.100 523.950 22.200 524.400 ;
        RECT 31.950 523.800 34.050 524.400 ;
        RECT 49.800 525.000 52.050 526.050 ;
        RECT 53.100 525.600 55.200 526.050 ;
        RECT 64.950 525.600 67.050 526.200 ;
        RECT 79.950 525.600 82.050 525.900 ;
        RECT 49.800 523.950 51.900 525.000 ;
        RECT 53.100 524.400 82.050 525.600 ;
        RECT 53.100 523.950 55.200 524.400 ;
        RECT 64.950 524.100 67.050 524.400 ;
        RECT 79.950 523.800 82.050 524.400 ;
        RECT 106.950 525.600 109.050 526.050 ;
        RECT 121.950 525.600 124.050 527.400 ;
        RECT 151.950 526.950 154.050 527.400 ;
        RECT 177.000 526.950 181.050 527.400 ;
        RECT 229.950 526.950 235.050 529.050 ;
        RECT 238.950 528.600 241.050 529.050 ;
        RECT 259.950 528.600 262.050 532.050 ;
        RECT 327.000 531.600 331.050 532.050 ;
        RECT 326.400 529.950 331.050 531.600 ;
        RECT 364.950 531.600 367.050 532.050 ;
        RECT 373.950 531.600 376.050 532.050 ;
        RECT 364.950 530.400 376.050 531.600 ;
        RECT 364.950 529.950 367.050 530.400 ;
        RECT 373.950 529.950 376.050 530.400 ;
        RECT 238.950 528.000 262.050 528.600 ;
        RECT 295.950 528.600 298.050 528.900 ;
        RECT 326.400 528.600 327.600 529.950 ;
        RECT 238.950 527.400 261.600 528.000 ;
        RECT 295.950 527.400 327.600 528.600 ;
        RECT 370.950 528.600 373.050 528.900 ;
        RECT 382.950 528.600 385.050 529.050 ;
        RECT 370.950 527.400 385.050 528.600 ;
        RECT 238.950 526.950 241.050 527.400 ;
        RECT 295.950 526.800 298.050 527.400 ;
        RECT 370.950 526.800 373.050 527.400 ;
        RECT 382.950 526.950 385.050 527.400 ;
        RECT 439.950 528.600 442.050 529.050 ;
        RECT 454.950 528.600 457.050 529.200 ;
        RECT 439.950 527.400 457.050 528.600 ;
        RECT 439.950 526.950 442.050 527.400 ;
        RECT 454.950 527.100 457.050 527.400 ;
        RECT 106.950 524.400 124.050 525.600 ;
        RECT 106.950 523.950 109.050 524.400 ;
        RECT 121.950 523.950 124.050 524.400 ;
        RECT 454.950 525.600 457.050 525.900 ;
        RECT 475.950 525.600 478.050 529.050 ;
        RECT 532.950 528.600 535.050 529.050 ;
        RECT 565.950 528.600 568.050 529.050 ;
        RECT 532.950 527.400 568.050 528.600 ;
        RECT 532.950 526.950 535.050 527.400 ;
        RECT 565.950 526.950 568.050 527.400 ;
        RECT 574.950 528.600 577.050 529.050 ;
        RECT 592.950 528.600 595.050 529.050 ;
        RECT 574.950 527.400 595.050 528.600 ;
        RECT 574.950 526.950 577.050 527.400 ;
        RECT 592.950 526.950 595.050 527.400 ;
        RECT 619.950 528.600 622.050 529.050 ;
        RECT 634.950 528.600 637.050 532.050 ;
        RECT 658.950 531.600 661.050 532.050 ;
        RECT 673.950 531.600 676.050 532.050 ;
        RECT 658.950 530.400 676.050 531.600 ;
        RECT 658.950 529.950 661.050 530.400 ;
        RECT 673.950 529.950 676.050 530.400 ;
        RECT 784.950 531.600 787.050 532.050 ;
        RECT 799.950 531.600 802.050 532.050 ;
        RECT 784.950 530.400 802.050 531.600 ;
        RECT 784.950 529.950 787.050 530.400 ;
        RECT 799.950 529.950 802.050 530.400 ;
        RECT 619.950 528.000 637.050 528.600 ;
        RECT 619.950 527.400 636.600 528.000 ;
        RECT 619.950 526.950 622.050 527.400 ;
        RECT 454.950 525.000 478.050 525.600 ;
        RECT 454.950 524.400 477.600 525.000 ;
        RECT 454.950 523.800 457.050 524.400 ;
        RECT 43.950 522.600 46.050 523.050 ;
        RECT 82.950 522.600 85.050 523.050 ;
        RECT 43.950 521.400 85.050 522.600 ;
        RECT 43.950 520.950 46.050 521.400 ;
        RECT 82.950 520.950 85.050 521.400 ;
        RECT 340.950 522.600 343.050 523.050 ;
        RECT 403.950 522.600 406.050 523.050 ;
        RECT 340.950 521.400 406.050 522.600 ;
        RECT 340.950 520.950 343.050 521.400 ;
        RECT 403.950 520.950 406.050 521.400 ;
        RECT 466.950 522.600 469.050 523.050 ;
        RECT 493.950 522.600 496.050 526.050 ;
        RECT 502.950 525.600 505.050 526.050 ;
        RECT 514.950 525.600 517.050 526.050 ;
        RECT 502.950 524.400 517.050 525.600 ;
        RECT 502.950 523.950 505.050 524.400 ;
        RECT 514.950 523.950 517.050 524.400 ;
        RECT 499.950 522.600 502.050 523.050 ;
        RECT 466.950 521.400 502.050 522.600 ;
        RECT 466.950 520.950 469.050 521.400 ;
        RECT 499.950 520.950 502.050 521.400 ;
        RECT 520.950 522.600 523.050 523.050 ;
        RECT 529.950 522.600 532.050 526.050 ;
        RECT 586.950 525.600 589.050 526.050 ;
        RECT 581.400 525.000 589.050 525.600 ;
        RECT 580.950 524.400 589.050 525.000 ;
        RECT 556.950 522.600 559.050 522.900 ;
        RECT 520.950 521.400 559.050 522.600 ;
        RECT 520.950 520.950 523.050 521.400 ;
        RECT 556.950 520.800 559.050 521.400 ;
        RECT 580.950 520.950 583.050 524.400 ;
        RECT 586.950 523.950 589.050 524.400 ;
        RECT 637.950 525.600 640.050 526.050 ;
        RECT 652.950 525.600 655.050 526.050 ;
        RECT 637.950 524.400 655.050 525.600 ;
        RECT 637.950 523.950 640.050 524.400 ;
        RECT 652.950 523.950 655.050 524.400 ;
        RECT 658.950 525.600 661.050 526.050 ;
        RECT 676.950 525.600 679.050 526.050 ;
        RECT 685.950 525.600 688.050 526.050 ;
        RECT 658.950 524.400 688.050 525.600 ;
        RECT 658.950 523.950 661.050 524.400 ;
        RECT 676.950 523.950 679.050 524.400 ;
        RECT 685.950 523.950 688.050 524.400 ;
        RECT 715.950 525.600 718.050 525.900 ;
        RECT 757.950 525.600 760.050 526.050 ;
        RECT 715.950 524.400 760.050 525.600 ;
        RECT 715.950 523.800 718.050 524.400 ;
        RECT 757.950 523.950 760.050 524.400 ;
        RECT 769.950 525.600 772.050 526.050 ;
        RECT 778.950 525.600 781.050 526.050 ;
        RECT 769.950 524.400 781.050 525.600 ;
        RECT 769.950 523.950 772.050 524.400 ;
        RECT 778.950 523.950 781.050 524.400 ;
        RECT 796.950 525.600 799.050 526.050 ;
        RECT 817.950 525.600 820.050 526.050 ;
        RECT 796.950 524.400 820.050 525.600 ;
        RECT 796.950 523.950 799.050 524.400 ;
        RECT 817.950 523.950 820.050 524.400 ;
        RECT 703.950 522.600 706.050 523.050 ;
        RECT 727.800 522.600 729.900 523.050 ;
        RECT 703.950 521.400 729.900 522.600 ;
        RECT 703.950 520.950 706.050 521.400 ;
        RECT 727.800 520.950 729.900 521.400 ;
        RECT 731.100 522.600 733.200 523.050 ;
        RECT 739.950 522.600 742.050 523.050 ;
        RECT 754.950 522.600 757.050 523.050 ;
        RECT 731.100 521.400 757.050 522.600 ;
        RECT 731.100 520.950 733.200 521.400 ;
        RECT 739.950 520.950 742.050 521.400 ;
        RECT 754.950 520.950 757.050 521.400 ;
        RECT 55.950 519.600 58.050 520.050 ;
        RECT 70.950 519.600 73.050 520.050 ;
        RECT 55.950 518.400 73.050 519.600 ;
        RECT 55.950 517.950 58.050 518.400 ;
        RECT 70.950 517.950 73.050 518.400 ;
        RECT 163.950 519.600 166.050 520.050 ;
        RECT 202.950 519.600 205.050 520.050 ;
        RECT 163.950 518.400 205.050 519.600 ;
        RECT 163.950 517.950 166.050 518.400 ;
        RECT 202.950 517.950 205.050 518.400 ;
        RECT 259.950 519.600 262.050 520.050 ;
        RECT 586.950 519.600 589.050 520.050 ;
        RECT 598.950 519.600 601.050 520.050 ;
        RECT 604.950 519.600 607.050 520.050 ;
        RECT 259.950 518.400 342.600 519.600 ;
        RECT 259.950 517.950 262.050 518.400 ;
        RECT 76.950 516.600 79.050 517.050 ;
        RECT 106.950 516.600 109.050 517.050 ;
        RECT 76.950 515.400 109.050 516.600 ;
        RECT 76.950 514.950 79.050 515.400 ;
        RECT 106.950 514.950 109.050 515.400 ;
        RECT 232.950 516.600 235.050 517.050 ;
        RECT 256.950 516.600 259.050 517.050 ;
        RECT 232.950 515.400 259.050 516.600 ;
        RECT 341.400 516.600 342.600 518.400 ;
        RECT 586.950 518.400 607.050 519.600 ;
        RECT 586.950 517.950 589.050 518.400 ;
        RECT 598.950 517.950 601.050 518.400 ;
        RECT 604.950 517.950 607.050 518.400 ;
        RECT 709.950 519.600 712.050 520.050 ;
        RECT 742.950 519.600 745.050 520.050 ;
        RECT 709.950 518.400 745.050 519.600 ;
        RECT 709.950 517.950 712.050 518.400 ;
        RECT 742.950 517.950 745.050 518.400 ;
        RECT 757.950 519.600 760.050 520.050 ;
        RECT 769.950 519.600 772.050 520.050 ;
        RECT 757.950 518.400 772.050 519.600 ;
        RECT 757.950 517.950 760.050 518.400 ;
        RECT 769.950 517.950 772.050 518.400 ;
        RECT 358.950 516.600 361.050 517.050 ;
        RECT 341.400 515.400 361.050 516.600 ;
        RECT 232.950 514.950 235.050 515.400 ;
        RECT 256.950 514.950 259.050 515.400 ;
        RECT 358.950 514.950 361.050 515.400 ;
        RECT 376.950 516.600 379.050 517.050 ;
        RECT 385.950 516.600 388.050 517.050 ;
        RECT 376.950 515.400 388.050 516.600 ;
        RECT 376.950 514.950 379.050 515.400 ;
        RECT 385.950 514.950 388.050 515.400 ;
        RECT 463.950 516.600 466.050 517.050 ;
        RECT 517.950 516.600 520.050 517.050 ;
        RECT 463.950 515.400 520.050 516.600 ;
        RECT 463.950 514.950 466.050 515.400 ;
        RECT 517.950 514.950 520.050 515.400 ;
        RECT 556.950 516.600 559.050 517.050 ;
        RECT 607.950 516.600 610.050 517.050 ;
        RECT 556.950 515.400 610.050 516.600 ;
        RECT 556.950 514.950 559.050 515.400 ;
        RECT 607.950 514.950 610.050 515.400 ;
        RECT 760.950 516.600 763.050 517.050 ;
        RECT 790.950 516.600 793.050 517.050 ;
        RECT 760.950 515.400 793.050 516.600 ;
        RECT 760.950 514.950 763.050 515.400 ;
        RECT 790.950 514.950 793.050 515.400 ;
        RECT 271.950 513.600 274.050 514.050 ;
        RECT 322.950 513.600 325.050 514.050 ;
        RECT 271.950 512.400 325.050 513.600 ;
        RECT 271.950 511.950 274.050 512.400 ;
        RECT 322.950 511.950 325.050 512.400 ;
        RECT 460.950 513.600 463.050 514.050 ;
        RECT 499.950 513.600 502.050 514.050 ;
        RECT 460.950 512.400 502.050 513.600 ;
        RECT 460.950 511.950 463.050 512.400 ;
        RECT 499.950 511.950 502.050 512.400 ;
        RECT 547.950 513.600 550.050 514.050 ;
        RECT 601.950 513.600 604.050 514.050 ;
        RECT 547.950 512.400 604.050 513.600 ;
        RECT 547.950 511.950 550.050 512.400 ;
        RECT 601.950 511.950 604.050 512.400 ;
        RECT 679.950 513.600 682.050 514.050 ;
        RECT 697.950 513.600 700.050 514.050 ;
        RECT 679.950 512.400 700.050 513.600 ;
        RECT 679.950 511.950 682.050 512.400 ;
        RECT 697.950 511.950 700.050 512.400 ;
        RECT 718.950 513.600 721.050 514.050 ;
        RECT 757.950 513.600 760.050 514.050 ;
        RECT 718.950 512.400 760.050 513.600 ;
        RECT 718.950 511.950 721.050 512.400 ;
        RECT 757.950 511.950 760.050 512.400 ;
        RECT 769.950 513.600 772.050 514.050 ;
        RECT 805.950 513.600 808.050 514.050 ;
        RECT 769.950 512.400 808.050 513.600 ;
        RECT 769.950 511.950 772.050 512.400 ;
        RECT 805.950 511.950 808.050 512.400 ;
        RECT 112.950 510.600 115.050 511.050 ;
        RECT 130.950 510.600 133.050 511.050 ;
        RECT 199.950 510.600 202.050 511.050 ;
        RECT 208.950 510.600 211.050 511.050 ;
        RECT 112.950 509.400 147.600 510.600 ;
        RECT 112.950 508.950 115.050 509.400 ;
        RECT 130.950 508.950 133.050 509.400 ;
        RECT 146.400 508.050 147.600 509.400 ;
        RECT 199.950 509.400 211.050 510.600 ;
        RECT 199.950 508.950 202.050 509.400 ;
        RECT 208.950 508.950 211.050 509.400 ;
        RECT 352.950 510.600 355.050 511.050 ;
        RECT 421.950 510.600 424.050 511.050 ;
        RECT 352.950 509.400 424.050 510.600 ;
        RECT 352.950 508.950 355.050 509.400 ;
        RECT 421.950 508.950 424.050 509.400 ;
        RECT 472.950 510.600 475.050 511.050 ;
        RECT 500.400 510.600 501.600 511.950 ;
        RECT 625.950 510.600 628.050 511.050 ;
        RECT 472.950 509.400 483.600 510.600 ;
        RECT 500.400 509.400 628.050 510.600 ;
        RECT 472.950 508.950 475.050 509.400 ;
        RECT 145.950 507.600 148.050 508.050 ;
        RECT 163.950 507.600 166.050 508.050 ;
        RECT 145.950 506.400 166.050 507.600 ;
        RECT 145.950 505.950 148.050 506.400 ;
        RECT 163.950 505.950 166.050 506.400 ;
        RECT 235.950 507.600 238.050 508.050 ;
        RECT 265.950 507.600 268.050 508.050 ;
        RECT 286.950 507.600 289.050 508.050 ;
        RECT 235.950 506.400 289.050 507.600 ;
        RECT 235.950 505.950 238.050 506.400 ;
        RECT 265.950 505.950 268.050 506.400 ;
        RECT 286.950 505.950 289.050 506.400 ;
        RECT 328.950 507.600 331.050 508.050 ;
        RECT 361.950 507.600 364.050 508.050 ;
        RECT 328.950 506.400 364.050 507.600 ;
        RECT 482.400 507.600 483.600 509.400 ;
        RECT 625.950 508.950 628.050 509.400 ;
        RECT 712.950 510.600 715.050 511.050 ;
        RECT 763.950 510.600 766.050 511.050 ;
        RECT 712.950 509.400 766.050 510.600 ;
        RECT 712.950 508.950 715.050 509.400 ;
        RECT 763.950 508.950 766.050 509.400 ;
        RECT 511.950 507.600 514.050 508.050 ;
        RECT 482.400 506.400 514.050 507.600 ;
        RECT 328.950 505.950 331.050 506.400 ;
        RECT 361.950 505.950 364.050 506.400 ;
        RECT 511.950 505.950 514.050 506.400 ;
        RECT 694.950 507.600 697.050 508.050 ;
        RECT 709.950 507.600 712.050 508.050 ;
        RECT 694.950 506.400 712.050 507.600 ;
        RECT 694.950 505.950 697.050 506.400 ;
        RECT 709.950 505.950 712.050 506.400 ;
        RECT 787.950 507.600 790.050 508.050 ;
        RECT 823.950 507.600 826.050 508.050 ;
        RECT 787.950 506.400 826.050 507.600 ;
        RECT 787.950 505.950 790.050 506.400 ;
        RECT 823.950 505.950 826.050 506.400 ;
        RECT 148.950 504.600 151.050 505.050 ;
        RECT 199.950 504.600 202.050 505.050 ;
        RECT 148.950 503.400 202.050 504.600 ;
        RECT 148.950 502.950 151.050 503.400 ;
        RECT 199.950 502.950 202.050 503.400 ;
        RECT 232.950 504.600 235.050 505.050 ;
        RECT 268.950 504.600 271.050 505.050 ;
        RECT 232.950 503.400 271.050 504.600 ;
        RECT 232.950 502.950 235.050 503.400 ;
        RECT 268.950 502.950 271.050 503.400 ;
        RECT 313.950 504.600 316.050 505.050 ;
        RECT 358.950 504.600 361.050 505.050 ;
        RECT 391.950 504.600 394.050 505.050 ;
        RECT 454.950 504.600 457.050 505.050 ;
        RECT 313.950 503.400 457.050 504.600 ;
        RECT 313.950 502.950 316.050 503.400 ;
        RECT 358.950 502.950 361.050 503.400 ;
        RECT 391.950 502.950 394.050 503.400 ;
        RECT 454.950 502.950 457.050 503.400 ;
        RECT 514.950 504.600 517.050 505.050 ;
        RECT 532.950 504.600 535.050 505.050 ;
        RECT 514.950 503.400 535.050 504.600 ;
        RECT 514.950 502.950 517.050 503.400 ;
        RECT 532.950 502.950 535.050 503.400 ;
        RECT 538.950 504.600 541.050 505.050 ;
        RECT 580.950 504.600 583.050 505.050 ;
        RECT 538.950 503.400 583.050 504.600 ;
        RECT 538.950 502.950 541.050 503.400 ;
        RECT 580.950 502.950 583.050 503.400 ;
        RECT 625.950 504.600 628.050 505.050 ;
        RECT 646.950 504.600 649.050 505.050 ;
        RECT 625.950 503.400 649.050 504.600 ;
        RECT 625.950 502.950 628.050 503.400 ;
        RECT 646.950 502.950 649.050 503.400 ;
        RECT 43.950 501.600 46.050 502.050 ;
        RECT 64.950 501.600 67.050 502.050 ;
        RECT 43.950 500.400 67.050 501.600 ;
        RECT 43.950 499.950 46.050 500.400 ;
        RECT 64.950 499.950 67.050 500.400 ;
        RECT 97.950 501.600 100.050 502.050 ;
        RECT 103.950 501.600 106.050 502.050 ;
        RECT 127.950 501.600 130.050 502.050 ;
        RECT 142.950 501.600 145.050 502.050 ;
        RECT 97.950 500.400 145.050 501.600 ;
        RECT 97.950 499.950 100.050 500.400 ;
        RECT 103.950 499.950 106.050 500.400 ;
        RECT 127.950 499.950 130.050 500.400 ;
        RECT 142.950 499.950 145.050 500.400 ;
        RECT 184.950 501.600 187.050 502.050 ;
        RECT 223.950 501.600 226.050 502.050 ;
        RECT 184.950 500.400 226.050 501.600 ;
        RECT 184.950 499.950 187.050 500.400 ;
        RECT 223.950 499.950 226.050 500.400 ;
        RECT 283.950 501.600 286.050 502.050 ;
        RECT 388.950 501.600 391.050 502.050 ;
        RECT 283.950 500.400 391.050 501.600 ;
        RECT 283.950 499.950 286.050 500.400 ;
        RECT 388.950 499.950 391.050 500.400 ;
        RECT 478.950 501.600 481.050 502.050 ;
        RECT 526.950 501.600 529.050 502.050 ;
        RECT 478.950 500.400 529.050 501.600 ;
        RECT 478.950 499.950 481.050 500.400 ;
        RECT 526.950 499.950 529.050 500.400 ;
        RECT 691.950 501.600 694.050 502.050 ;
        RECT 703.950 501.600 706.050 502.050 ;
        RECT 691.950 500.400 706.050 501.600 ;
        RECT 691.950 499.950 694.050 500.400 ;
        RECT 703.950 499.950 706.050 500.400 ;
        RECT 754.950 501.600 757.050 502.050 ;
        RECT 766.950 501.600 769.050 502.050 ;
        RECT 754.950 500.400 769.050 501.600 ;
        RECT 754.950 499.950 757.050 500.400 ;
        RECT 766.950 499.950 769.050 500.400 ;
        RECT 205.950 498.600 208.050 499.050 ;
        RECT 229.950 498.600 232.050 499.050 ;
        RECT 205.950 497.400 232.050 498.600 ;
        RECT 205.950 496.950 208.050 497.400 ;
        RECT 229.950 496.950 232.050 497.400 ;
        RECT 82.950 495.600 85.050 496.050 ;
        RECT 109.950 495.600 112.050 496.050 ;
        RECT 118.950 495.600 121.050 496.050 ;
        RECT 82.950 494.400 121.050 495.600 ;
        RECT 82.950 493.950 85.050 494.400 ;
        RECT 109.950 493.950 112.050 494.400 ;
        RECT 118.950 493.950 121.050 494.400 ;
        RECT 196.950 495.600 199.050 496.050 ;
        RECT 238.950 495.600 241.050 496.050 ;
        RECT 259.950 495.600 262.050 496.050 ;
        RECT 196.950 494.400 241.050 495.600 ;
        RECT 254.400 495.000 262.050 495.600 ;
        RECT 196.950 493.950 199.050 494.400 ;
        RECT 238.950 493.950 241.050 494.400 ;
        RECT 253.950 494.400 262.050 495.000 ;
        RECT 130.950 492.600 133.050 493.200 ;
        RECT 139.950 492.600 142.050 493.200 ;
        RECT 130.950 491.400 142.050 492.600 ;
        RECT 130.950 491.100 133.050 491.400 ;
        RECT 139.950 491.100 142.050 491.400 ;
        RECT 154.950 492.600 157.050 493.050 ;
        RECT 160.950 492.600 163.050 493.050 ;
        RECT 154.950 491.400 163.050 492.600 ;
        RECT 154.950 490.950 157.050 491.400 ;
        RECT 160.950 490.950 163.050 491.400 ;
        RECT 169.950 492.600 172.050 493.050 ;
        RECT 175.950 492.600 178.050 493.050 ;
        RECT 169.950 491.400 178.050 492.600 ;
        RECT 169.950 490.950 172.050 491.400 ;
        RECT 175.950 490.950 178.050 491.400 ;
        RECT 199.950 492.600 202.050 493.050 ;
        RECT 232.950 492.600 235.050 493.050 ;
        RECT 199.950 491.400 235.050 492.600 ;
        RECT 199.950 490.950 202.050 491.400 ;
        RECT 232.950 490.950 235.050 491.400 ;
        RECT 253.950 490.950 256.050 494.400 ;
        RECT 259.950 493.950 262.050 494.400 ;
        RECT 268.950 495.600 271.050 496.050 ;
        RECT 298.950 495.600 301.050 496.050 ;
        RECT 310.950 495.600 313.050 496.050 ;
        RECT 268.950 494.400 313.050 495.600 ;
        RECT 346.950 495.600 349.050 499.050 ;
        RECT 604.950 498.600 607.050 499.050 ;
        RECT 655.950 498.600 658.050 499.050 ;
        RECT 604.950 497.400 658.050 498.600 ;
        RECT 604.950 496.950 607.050 497.400 ;
        RECT 655.950 496.950 658.050 497.400 ;
        RECT 733.950 498.600 736.050 499.050 ;
        RECT 748.950 498.600 751.050 499.050 ;
        RECT 733.950 497.400 751.050 498.600 ;
        RECT 733.950 496.950 736.050 497.400 ;
        RECT 748.950 496.950 751.050 497.400 ;
        RECT 784.950 498.600 787.050 499.050 ;
        RECT 814.950 498.600 817.050 499.050 ;
        RECT 784.950 497.400 817.050 498.600 ;
        RECT 784.950 496.950 787.050 497.400 ;
        RECT 814.950 496.950 817.050 497.400 ;
        RECT 358.950 495.600 361.050 496.200 ;
        RECT 346.950 495.000 361.050 495.600 ;
        RECT 347.400 494.400 361.050 495.000 ;
        RECT 268.950 493.950 271.050 494.400 ;
        RECT 298.950 493.950 301.050 494.400 ;
        RECT 310.950 493.950 313.050 494.400 ;
        RECT 358.950 494.100 361.050 494.400 ;
        RECT 502.950 495.600 505.050 496.050 ;
        RECT 508.950 495.600 511.050 496.050 ;
        RECT 502.950 494.400 511.050 495.600 ;
        RECT 502.950 493.950 505.050 494.400 ;
        RECT 508.950 493.950 511.050 494.400 ;
        RECT 607.950 495.600 610.050 496.050 ;
        RECT 625.950 495.600 628.050 496.050 ;
        RECT 607.950 494.400 628.050 495.600 ;
        RECT 607.950 493.950 610.050 494.400 ;
        RECT 625.950 493.950 628.050 494.400 ;
        RECT 697.950 495.600 700.050 496.050 ;
        RECT 706.950 495.600 709.050 496.050 ;
        RECT 697.950 494.400 709.050 495.600 ;
        RECT 697.950 493.950 700.050 494.400 ;
        RECT 706.950 493.950 709.050 494.400 ;
        RECT 727.950 495.600 730.050 496.050 ;
        RECT 736.950 495.600 739.050 496.050 ;
        RECT 727.950 494.400 739.050 495.600 ;
        RECT 727.950 493.950 730.050 494.400 ;
        RECT 736.950 493.950 739.050 494.400 ;
        RECT 751.950 495.600 754.050 496.050 ;
        RECT 769.950 495.600 775.050 496.050 ;
        RECT 751.950 494.400 775.050 495.600 ;
        RECT 751.950 493.950 754.050 494.400 ;
        RECT 769.950 493.950 775.050 494.400 ;
        RECT 796.950 495.600 799.050 496.050 ;
        RECT 817.950 495.600 820.050 496.050 ;
        RECT 796.950 494.400 820.050 495.600 ;
        RECT 796.950 493.950 799.050 494.400 ;
        RECT 817.950 493.950 820.050 494.400 ;
        RECT 364.950 492.600 367.050 493.050 ;
        RECT 391.950 492.600 394.050 493.050 ;
        RECT 364.950 491.400 394.050 492.600 ;
        RECT 364.950 490.950 367.050 491.400 ;
        RECT 391.950 490.950 394.050 491.400 ;
        RECT 433.950 492.600 436.050 493.050 ;
        RECT 490.950 492.600 493.050 493.050 ;
        RECT 433.950 491.400 493.050 492.600 ;
        RECT 433.950 490.950 436.050 491.400 ;
        RECT 490.950 490.950 493.050 491.400 ;
        RECT 535.950 492.600 538.050 493.050 ;
        RECT 568.950 492.600 574.050 493.050 ;
        RECT 535.950 491.400 574.050 492.600 ;
        RECT 535.950 490.950 538.050 491.400 ;
        RECT 568.950 490.950 574.050 491.400 ;
        RECT 619.950 492.600 622.050 493.050 ;
        RECT 649.950 492.600 652.050 493.050 ;
        RECT 664.950 492.600 667.050 493.050 ;
        RECT 679.950 492.600 682.050 493.050 ;
        RECT 619.950 491.400 645.600 492.600 ;
        RECT 619.950 490.950 622.050 491.400 ;
        RECT 10.950 489.600 13.050 490.200 ;
        RECT 19.950 489.600 22.050 490.050 ;
        RECT 10.950 488.400 22.050 489.600 ;
        RECT 10.950 488.100 13.050 488.400 ;
        RECT 19.950 487.950 22.050 488.400 ;
        RECT 184.950 489.600 187.050 490.050 ;
        RECT 196.950 489.600 199.050 490.050 ;
        RECT 184.950 488.400 199.050 489.600 ;
        RECT 184.950 487.950 187.050 488.400 ;
        RECT 196.950 487.950 199.050 488.400 ;
        RECT 304.950 489.600 307.050 490.050 ;
        RECT 319.950 489.600 322.050 490.050 ;
        RECT 304.950 488.400 322.050 489.600 ;
        RECT 304.950 487.950 307.050 488.400 ;
        RECT 319.950 487.950 322.050 488.400 ;
        RECT 397.950 487.950 403.050 490.050 ;
        RECT 448.950 489.600 451.050 490.050 ;
        RECT 466.950 489.600 469.050 490.050 ;
        RECT 448.950 488.400 469.050 489.600 ;
        RECT 448.950 487.950 451.050 488.400 ;
        RECT 466.950 487.950 469.050 488.400 ;
        RECT 514.950 489.600 517.050 490.050 ;
        RECT 526.950 489.600 529.050 490.050 ;
        RECT 514.950 488.400 529.050 489.600 ;
        RECT 514.950 487.950 517.050 488.400 ;
        RECT 526.950 487.950 529.050 488.400 ;
        RECT 628.950 489.600 631.050 490.050 ;
        RECT 637.950 489.600 640.050 490.050 ;
        RECT 628.950 488.400 640.050 489.600 ;
        RECT 644.400 489.600 645.600 491.400 ;
        RECT 649.950 491.400 667.050 492.600 ;
        RECT 649.950 490.950 652.050 491.400 ;
        RECT 664.950 490.950 667.050 491.400 ;
        RECT 674.400 491.400 682.050 492.600 ;
        RECT 655.950 489.600 658.050 490.050 ;
        RECT 670.950 489.600 673.050 490.200 ;
        RECT 644.400 488.400 673.050 489.600 ;
        RECT 628.950 487.950 631.050 488.400 ;
        RECT 637.950 487.950 640.050 488.400 ;
        RECT 655.950 487.950 658.050 488.400 ;
        RECT 670.950 488.100 673.050 488.400 ;
        RECT 674.400 487.050 675.600 491.400 ;
        RECT 679.950 490.950 682.050 491.400 ;
        RECT 739.950 492.600 742.050 493.050 ;
        RECT 748.950 492.600 751.050 493.050 ;
        RECT 739.950 491.400 751.050 492.600 ;
        RECT 739.950 490.950 742.050 491.400 ;
        RECT 748.950 490.950 751.050 491.400 ;
        RECT 724.950 487.950 730.050 490.050 ;
        RECT 754.950 489.600 757.050 490.050 ;
        RECT 766.950 489.600 769.050 490.050 ;
        RECT 754.950 488.400 769.050 489.600 ;
        RECT 754.950 487.950 757.050 488.400 ;
        RECT 766.950 487.950 769.050 488.400 ;
        RECT 7.950 486.600 10.050 486.900 ;
        RECT 13.950 486.600 16.050 487.050 ;
        RECT 7.950 485.400 16.050 486.600 ;
        RECT 7.950 484.800 10.050 485.400 ;
        RECT 13.950 484.950 16.050 485.400 ;
        RECT 82.950 486.600 85.050 487.050 ;
        RECT 103.950 486.600 106.050 487.050 ;
        RECT 118.950 486.600 121.050 487.050 ;
        RECT 139.950 486.600 142.050 487.050 ;
        RECT 253.950 486.600 256.050 487.050 ;
        RECT 82.950 485.400 142.050 486.600 ;
        RECT 218.400 486.000 256.050 486.600 ;
        RECT 82.950 484.950 85.050 485.400 ;
        RECT 103.950 484.950 106.050 485.400 ;
        RECT 118.950 484.950 121.050 485.400 ;
        RECT 139.950 484.950 142.050 485.400 ;
        RECT 217.950 485.400 256.050 486.000 ;
        RECT 100.950 483.600 103.050 484.050 ;
        RECT 109.950 483.600 112.050 484.050 ;
        RECT 130.950 483.600 133.050 484.050 ;
        RECT 100.950 482.400 133.050 483.600 ;
        RECT 100.950 481.950 103.050 482.400 ;
        RECT 109.950 481.950 112.050 482.400 ;
        RECT 130.950 481.950 133.050 482.400 ;
        RECT 217.950 482.100 220.050 485.400 ;
        RECT 253.950 484.950 256.050 485.400 ;
        RECT 274.950 486.600 277.050 487.050 ;
        RECT 283.950 486.600 286.050 487.050 ;
        RECT 274.950 485.400 286.050 486.600 ;
        RECT 274.950 484.950 277.050 485.400 ;
        RECT 283.950 484.950 286.050 485.400 ;
        RECT 340.950 486.600 343.050 487.050 ;
        RECT 475.950 486.600 478.050 487.050 ;
        RECT 340.950 485.400 478.050 486.600 ;
        RECT 340.950 484.950 343.050 485.400 ;
        RECT 475.950 484.950 478.050 485.400 ;
        RECT 538.950 486.600 541.050 487.050 ;
        RECT 592.950 486.600 595.050 487.050 ;
        RECT 616.950 486.600 619.050 487.050 ;
        RECT 622.950 486.600 625.050 487.050 ;
        RECT 672.000 486.900 675.600 487.050 ;
        RECT 538.950 485.400 625.050 486.600 ;
        RECT 538.950 484.950 541.050 485.400 ;
        RECT 592.950 484.950 595.050 485.400 ;
        RECT 616.950 484.950 619.050 485.400 ;
        RECT 622.950 484.950 625.050 485.400 ;
        RECT 670.950 485.400 675.600 486.900 ;
        RECT 682.950 486.600 685.050 487.050 ;
        RECT 700.950 486.600 703.050 486.900 ;
        RECT 682.950 485.400 703.050 486.600 ;
        RECT 670.950 484.950 675.000 485.400 ;
        RECT 682.950 484.950 685.050 485.400 ;
        RECT 670.950 484.800 673.050 484.950 ;
        RECT 700.950 484.800 703.050 485.400 ;
        RECT 706.950 486.600 709.050 487.050 ;
        RECT 718.950 486.600 721.050 487.050 ;
        RECT 706.950 485.400 721.050 486.600 ;
        RECT 706.950 484.950 709.050 485.400 ;
        RECT 718.950 484.950 721.050 485.400 ;
        RECT 781.950 486.600 784.050 487.200 ;
        RECT 787.950 486.600 790.050 490.050 ;
        RECT 781.950 486.000 790.050 486.600 ;
        RECT 781.950 485.400 789.600 486.000 ;
        RECT 781.950 485.100 784.050 485.400 ;
        RECT 412.950 483.600 415.050 484.050 ;
        RECT 427.950 483.600 430.050 484.050 ;
        RECT 436.950 483.600 439.050 483.900 ;
        RECT 412.950 482.400 439.050 483.600 ;
        RECT 412.950 481.950 415.050 482.400 ;
        RECT 427.950 481.950 430.050 482.400 ;
        RECT 436.950 481.800 439.050 482.400 ;
        RECT 553.950 483.600 556.050 484.050 ;
        RECT 715.950 483.600 718.050 484.050 ;
        RECT 553.950 482.400 718.050 483.600 ;
        RECT 553.950 481.950 556.050 482.400 ;
        RECT 715.950 481.950 718.050 482.400 ;
        RECT 775.950 483.600 778.050 484.050 ;
        RECT 808.950 483.600 811.050 484.050 ;
        RECT 775.950 482.400 811.050 483.600 ;
        RECT 775.950 481.950 778.050 482.400 ;
        RECT 808.950 481.950 811.050 482.400 ;
        RECT 46.950 480.600 49.050 481.050 ;
        RECT 58.950 480.600 61.050 481.050 ;
        RECT 46.950 479.400 61.050 480.600 ;
        RECT 46.950 478.950 49.050 479.400 ;
        RECT 58.950 478.950 61.050 479.400 ;
        RECT 133.950 480.600 136.050 481.050 ;
        RECT 178.950 480.600 181.050 481.050 ;
        RECT 133.950 479.400 181.050 480.600 ;
        RECT 133.950 478.950 136.050 479.400 ;
        RECT 178.950 478.950 181.050 479.400 ;
        RECT 217.950 480.600 220.050 480.900 ;
        RECT 226.950 480.600 229.050 481.050 ;
        RECT 217.950 479.400 229.050 480.600 ;
        RECT 217.950 478.800 220.050 479.400 ;
        RECT 226.950 478.950 229.050 479.400 ;
        RECT 244.950 480.600 247.050 481.050 ;
        RECT 256.950 480.600 259.050 481.050 ;
        RECT 244.950 479.400 259.050 480.600 ;
        RECT 244.950 478.950 247.050 479.400 ;
        RECT 256.950 478.950 259.050 479.400 ;
        RECT 298.950 480.600 301.050 481.050 ;
        RECT 313.950 480.600 316.050 481.050 ;
        RECT 382.950 480.600 385.050 481.050 ;
        RECT 298.950 479.400 385.050 480.600 ;
        RECT 437.400 480.600 438.600 481.800 ;
        RECT 460.950 480.600 463.050 481.050 ;
        RECT 493.950 480.600 496.050 481.050 ;
        RECT 437.400 479.400 496.050 480.600 ;
        RECT 298.950 478.950 301.050 479.400 ;
        RECT 313.950 478.950 316.050 479.400 ;
        RECT 382.950 478.950 385.050 479.400 ;
        RECT 460.950 478.950 463.050 479.400 ;
        RECT 493.950 478.950 496.050 479.400 ;
        RECT 502.950 480.600 505.050 481.050 ;
        RECT 544.950 480.600 547.050 481.050 ;
        RECT 502.950 479.400 547.050 480.600 ;
        RECT 502.950 478.950 505.050 479.400 ;
        RECT 544.950 478.950 547.050 479.400 ;
        RECT 691.950 480.600 694.050 481.050 ;
        RECT 745.950 480.600 748.050 481.050 ;
        RECT 691.950 479.400 748.050 480.600 ;
        RECT 691.950 478.950 694.050 479.400 ;
        RECT 745.950 478.950 748.050 479.400 ;
        RECT 187.950 477.600 190.050 478.050 ;
        RECT 205.800 477.600 207.900 478.050 ;
        RECT 187.950 476.400 207.900 477.600 ;
        RECT 187.950 475.950 190.050 476.400 ;
        RECT 205.800 475.950 207.900 476.400 ;
        RECT 209.100 477.600 211.200 478.050 ;
        RECT 229.950 477.600 232.050 478.050 ;
        RECT 271.950 477.600 274.050 478.050 ;
        RECT 209.100 476.400 274.050 477.600 ;
        RECT 209.100 475.950 211.200 476.400 ;
        RECT 229.950 475.950 232.050 476.400 ;
        RECT 271.950 475.950 274.050 476.400 ;
        RECT 280.950 477.600 283.050 478.050 ;
        RECT 403.950 477.600 406.050 478.050 ;
        RECT 280.950 476.400 406.050 477.600 ;
        RECT 494.400 477.600 495.600 478.950 ;
        RECT 508.950 477.600 511.050 478.050 ;
        RECT 494.400 476.400 511.050 477.600 ;
        RECT 280.950 475.950 283.050 476.400 ;
        RECT 403.950 475.950 406.050 476.400 ;
        RECT 508.950 475.950 511.050 476.400 ;
        RECT 808.950 477.600 811.050 478.050 ;
        RECT 826.950 477.600 829.050 478.050 ;
        RECT 808.950 476.400 829.050 477.600 ;
        RECT 808.950 475.950 811.050 476.400 ;
        RECT 826.950 475.950 829.050 476.400 ;
        RECT 451.950 474.600 454.050 475.050 ;
        RECT 475.950 474.600 478.050 475.050 ;
        RECT 784.950 474.600 787.050 475.050 ;
        RECT 451.950 473.400 478.050 474.600 ;
        RECT 451.950 472.950 454.050 473.400 ;
        RECT 475.950 472.950 478.050 473.400 ;
        RECT 518.400 473.400 787.050 474.600 ;
        RECT 55.950 471.600 58.050 472.050 ;
        RECT 64.950 471.600 67.050 472.050 ;
        RECT 73.950 471.600 76.050 472.050 ;
        RECT 217.950 471.600 220.050 472.050 ;
        RECT 55.950 470.400 220.050 471.600 ;
        RECT 55.950 469.950 58.050 470.400 ;
        RECT 64.950 469.950 67.050 470.400 ;
        RECT 73.950 469.950 76.050 470.400 ;
        RECT 217.950 469.950 220.050 470.400 ;
        RECT 352.950 471.600 355.050 472.050 ;
        RECT 358.950 471.600 361.050 472.050 ;
        RECT 352.950 470.400 361.050 471.600 ;
        RECT 352.950 469.950 355.050 470.400 ;
        RECT 358.950 469.950 361.050 470.400 ;
        RECT 496.950 471.600 499.050 472.050 ;
        RECT 518.400 471.600 519.600 473.400 ;
        RECT 784.950 472.950 787.050 473.400 ;
        RECT 496.950 470.400 519.600 471.600 ;
        RECT 685.950 471.600 688.050 472.050 ;
        RECT 694.950 471.600 697.050 472.050 ;
        RECT 685.950 470.400 697.050 471.600 ;
        RECT 496.950 469.950 499.050 470.400 ;
        RECT 685.950 469.950 688.050 470.400 ;
        RECT 694.950 469.950 697.050 470.400 ;
        RECT 1.950 468.600 4.050 469.050 ;
        RECT 22.950 468.600 25.050 469.050 ;
        RECT 1.950 467.400 25.050 468.600 ;
        RECT 1.950 466.950 4.050 467.400 ;
        RECT 22.950 466.950 25.050 467.400 ;
        RECT 328.950 468.600 331.050 469.050 ;
        RECT 712.950 468.600 715.050 469.050 ;
        RECT 748.950 468.600 751.050 469.050 ;
        RECT 328.950 467.400 751.050 468.600 ;
        RECT 328.950 466.950 331.050 467.400 ;
        RECT 712.950 466.950 715.050 467.400 ;
        RECT 748.950 466.950 751.050 467.400 ;
        RECT 766.950 468.600 769.050 469.050 ;
        RECT 778.950 468.600 781.050 469.050 ;
        RECT 766.950 467.400 781.050 468.600 ;
        RECT 766.950 466.950 769.050 467.400 ;
        RECT 778.950 466.950 781.050 467.400 ;
        RECT 40.950 465.600 43.050 466.050 ;
        RECT 64.800 465.600 66.900 466.050 ;
        RECT 40.950 464.400 66.900 465.600 ;
        RECT 40.950 463.950 43.050 464.400 ;
        RECT 64.800 463.950 66.900 464.400 ;
        RECT 68.100 465.600 70.200 466.050 ;
        RECT 82.950 465.600 85.050 466.050 ;
        RECT 68.100 464.400 85.050 465.600 ;
        RECT 68.100 463.950 70.200 464.400 ;
        RECT 82.950 463.950 85.050 464.400 ;
        RECT 100.950 465.600 103.050 466.050 ;
        RECT 160.950 465.600 163.050 466.050 ;
        RECT 190.950 465.600 193.050 466.050 ;
        RECT 100.950 464.400 193.050 465.600 ;
        RECT 100.950 463.950 103.050 464.400 ;
        RECT 160.950 463.950 163.050 464.400 ;
        RECT 190.950 463.950 193.050 464.400 ;
        RECT 202.950 465.600 205.050 466.050 ;
        RECT 217.950 465.600 220.050 466.050 ;
        RECT 202.950 464.400 220.050 465.600 ;
        RECT 202.950 463.950 205.050 464.400 ;
        RECT 217.950 463.950 220.050 464.400 ;
        RECT 355.950 465.600 358.050 466.050 ;
        RECT 370.950 465.600 373.050 466.050 ;
        RECT 355.950 464.400 373.050 465.600 ;
        RECT 355.950 463.950 358.050 464.400 ;
        RECT 370.950 463.950 373.050 464.400 ;
        RECT 403.950 465.600 406.050 466.050 ;
        RECT 499.950 465.600 502.050 466.050 ;
        RECT 403.950 464.400 502.050 465.600 ;
        RECT 403.950 463.950 406.050 464.400 ;
        RECT 499.950 463.950 502.050 464.400 ;
        RECT 505.950 465.600 508.050 466.050 ;
        RECT 523.950 465.600 526.050 466.050 ;
        RECT 559.950 465.600 562.050 466.050 ;
        RECT 505.950 464.400 562.050 465.600 ;
        RECT 505.950 463.950 508.050 464.400 ;
        RECT 523.950 463.950 526.050 464.400 ;
        RECT 559.950 463.950 562.050 464.400 ;
        RECT 580.950 465.600 583.050 466.050 ;
        RECT 688.950 465.600 691.050 466.050 ;
        RECT 580.950 464.400 691.050 465.600 ;
        RECT 580.950 463.950 583.050 464.400 ;
        RECT 688.950 463.950 691.050 464.400 ;
        RECT 10.950 462.600 13.050 463.050 ;
        RECT 22.950 462.600 25.050 463.050 ;
        RECT 91.950 462.600 94.050 463.050 ;
        RECT 121.950 462.600 124.050 463.050 ;
        RECT 10.950 461.400 124.050 462.600 ;
        RECT 10.950 460.950 13.050 461.400 ;
        RECT 22.950 460.950 25.050 461.400 ;
        RECT 91.950 460.950 94.050 461.400 ;
        RECT 121.950 460.950 124.050 461.400 ;
        RECT 151.950 462.600 154.050 463.050 ;
        RECT 166.950 462.600 169.050 463.050 ;
        RECT 220.950 462.600 223.050 463.050 ;
        RECT 151.950 461.400 223.050 462.600 ;
        RECT 151.950 460.950 154.050 461.400 ;
        RECT 166.950 460.950 169.050 461.400 ;
        RECT 220.950 460.950 223.050 461.400 ;
        RECT 232.950 462.600 235.050 463.050 ;
        RECT 238.950 462.600 241.050 463.050 ;
        RECT 232.950 461.400 241.050 462.600 ;
        RECT 232.950 460.950 235.050 461.400 ;
        RECT 238.950 460.950 241.050 461.400 ;
        RECT 325.950 462.600 328.050 463.050 ;
        RECT 502.950 462.600 505.050 463.050 ;
        RECT 325.950 461.400 505.050 462.600 ;
        RECT 325.950 460.950 328.050 461.400 ;
        RECT 502.950 460.950 505.050 461.400 ;
        RECT 718.950 462.600 721.050 463.050 ;
        RECT 778.950 462.600 781.050 463.050 ;
        RECT 718.950 461.400 781.050 462.600 ;
        RECT 718.950 460.950 721.050 461.400 ;
        RECT 778.950 460.950 781.050 461.400 ;
        RECT 811.950 462.600 814.050 463.050 ;
        RECT 829.950 462.600 832.050 463.050 ;
        RECT 811.950 461.400 832.050 462.600 ;
        RECT 811.950 460.950 814.050 461.400 ;
        RECT 829.950 460.950 832.050 461.400 ;
        RECT 193.950 459.600 196.050 460.050 ;
        RECT 214.950 459.600 217.050 460.050 ;
        RECT 193.950 458.400 217.050 459.600 ;
        RECT 193.950 457.950 196.050 458.400 ;
        RECT 214.950 457.950 217.050 458.400 ;
        RECT 301.950 459.600 304.050 460.050 ;
        RECT 307.950 459.600 310.050 460.050 ;
        RECT 301.950 458.400 310.050 459.600 ;
        RECT 301.950 457.950 304.050 458.400 ;
        RECT 307.950 457.950 310.050 458.400 ;
        RECT 424.950 459.600 427.050 460.050 ;
        RECT 442.950 459.600 445.050 460.050 ;
        RECT 424.950 458.400 445.050 459.600 ;
        RECT 424.950 457.950 427.050 458.400 ;
        RECT 442.950 457.950 445.050 458.400 ;
        RECT 484.950 459.600 487.050 460.050 ;
        RECT 511.950 459.600 514.050 460.050 ;
        RECT 484.950 458.400 514.050 459.600 ;
        RECT 484.950 457.950 487.050 458.400 ;
        RECT 511.950 457.950 514.050 458.400 ;
        RECT 667.950 459.600 670.050 460.050 ;
        RECT 679.950 459.600 682.050 460.050 ;
        RECT 715.950 459.600 718.050 460.050 ;
        RECT 667.950 458.400 682.050 459.600 ;
        RECT 667.950 457.950 670.050 458.400 ;
        RECT 679.950 457.950 682.050 458.400 ;
        RECT 686.400 458.400 718.050 459.600 ;
        RECT 686.400 457.050 687.600 458.400 ;
        RECT 715.950 457.950 718.050 458.400 ;
        RECT 37.950 456.600 40.050 457.050 ;
        RECT 52.950 456.600 55.050 457.050 ;
        RECT 37.950 455.400 55.050 456.600 ;
        RECT 37.950 454.950 40.050 455.400 ;
        RECT 52.950 454.950 55.050 455.400 ;
        RECT 217.950 456.600 220.050 457.050 ;
        RECT 238.950 456.600 241.050 457.050 ;
        RECT 217.950 455.400 241.050 456.600 ;
        RECT 217.950 454.950 220.050 455.400 ;
        RECT 238.950 454.950 241.050 455.400 ;
        RECT 499.950 456.600 502.050 457.050 ;
        RECT 541.950 456.600 544.050 457.050 ;
        RECT 499.950 455.400 544.050 456.600 ;
        RECT 499.950 454.950 502.050 455.400 ;
        RECT 541.950 454.950 544.050 455.400 ;
        RECT 640.950 456.600 643.050 457.050 ;
        RECT 685.950 456.600 688.050 457.050 ;
        RECT 640.950 455.400 688.050 456.600 ;
        RECT 640.950 454.950 643.050 455.400 ;
        RECT 685.950 454.950 688.050 455.400 ;
        RECT 694.950 456.600 697.050 457.050 ;
        RECT 730.950 456.600 733.050 457.050 ;
        RECT 694.950 455.400 733.050 456.600 ;
        RECT 694.950 454.950 697.050 455.400 ;
        RECT 730.950 454.950 733.050 455.400 ;
        RECT 1.950 454.050 4.050 454.200 ;
        RECT 0.000 453.600 4.050 454.050 ;
        RECT -0.600 452.100 4.050 453.600 ;
        RECT 13.950 453.600 16.050 454.050 ;
        RECT 94.950 453.600 97.050 454.050 ;
        RECT 13.950 452.400 97.050 453.600 ;
        RECT -0.600 451.950 3.000 452.100 ;
        RECT 13.950 451.950 16.050 452.400 ;
        RECT -0.600 447.600 0.600 451.950 ;
        RECT 1.950 450.600 4.050 450.900 ;
        RECT 7.950 450.600 10.050 451.200 ;
        RECT 1.950 449.400 10.050 450.600 ;
        RECT 1.950 448.800 4.050 449.400 ;
        RECT 7.950 449.100 10.050 449.400 ;
        RECT 26.400 448.050 27.600 452.400 ;
        RECT 94.950 451.950 97.050 452.400 ;
        RECT 112.950 453.600 115.050 454.050 ;
        RECT 127.950 453.600 130.050 454.050 ;
        RECT 157.950 453.600 160.050 454.050 ;
        RECT 112.950 452.400 160.050 453.600 ;
        RECT 112.950 451.950 115.050 452.400 ;
        RECT 127.950 451.950 130.050 452.400 ;
        RECT 157.950 451.950 160.050 452.400 ;
        RECT 169.950 453.600 172.050 454.050 ;
        RECT 181.950 453.600 184.050 454.050 ;
        RECT 169.950 452.400 184.050 453.600 ;
        RECT 169.950 451.950 172.050 452.400 ;
        RECT 181.950 451.950 184.050 452.400 ;
        RECT 265.950 453.600 268.050 454.200 ;
        RECT 289.950 453.600 292.050 454.050 ;
        RECT 265.950 452.400 292.050 453.600 ;
        RECT 265.950 452.100 268.050 452.400 ;
        RECT 289.950 451.950 292.050 452.400 ;
        RECT 295.950 453.600 298.050 454.050 ;
        RECT 325.950 453.600 328.050 454.200 ;
        RECT 331.950 453.600 334.050 454.050 ;
        RECT 295.950 452.400 321.600 453.600 ;
        RECT 295.950 451.950 298.050 452.400 ;
        RECT 320.400 451.050 321.600 452.400 ;
        RECT 325.950 452.400 334.050 453.600 ;
        RECT 325.950 452.100 328.050 452.400 ;
        RECT 331.950 451.950 334.050 452.400 ;
        RECT 322.950 451.050 325.050 451.200 ;
        RECT 73.950 450.600 76.050 451.050 ;
        RECT 79.950 450.600 82.050 451.050 ;
        RECT 73.950 449.400 82.050 450.600 ;
        RECT 73.950 448.950 76.050 449.400 ;
        RECT 79.950 448.950 82.050 449.400 ;
        RECT 88.950 450.600 91.050 451.050 ;
        RECT 106.950 450.600 109.050 451.050 ;
        RECT 88.950 449.400 109.050 450.600 ;
        RECT 88.950 448.950 91.050 449.400 ;
        RECT 106.950 448.950 109.050 449.400 ;
        RECT 187.950 450.600 190.050 451.050 ;
        RECT 232.950 450.600 235.050 451.050 ;
        RECT 187.950 449.400 235.050 450.600 ;
        RECT 187.950 448.950 190.050 449.400 ;
        RECT 232.950 448.950 235.050 449.400 ;
        RECT 265.950 450.600 268.050 450.900 ;
        RECT 271.950 450.600 274.050 451.050 ;
        RECT 292.950 450.600 295.050 451.050 ;
        RECT 265.950 449.400 295.050 450.600 ;
        RECT 265.950 448.800 268.050 449.400 ;
        RECT 271.950 448.950 274.050 449.400 ;
        RECT 292.950 448.950 295.050 449.400 ;
        RECT 319.950 449.100 325.050 451.050 ;
        RECT 379.950 450.600 382.050 451.050 ;
        RECT 400.950 450.600 403.050 454.050 ;
        RECT 637.950 453.600 640.050 454.050 ;
        RECT 667.950 453.600 670.050 454.050 ;
        RECT 637.950 452.400 670.050 453.600 ;
        RECT 637.950 451.950 640.050 452.400 ;
        RECT 667.950 451.950 670.050 452.400 ;
        RECT 709.950 453.600 712.050 454.050 ;
        RECT 718.950 453.600 721.050 454.050 ;
        RECT 709.950 452.400 721.050 453.600 ;
        RECT 709.950 451.950 712.050 452.400 ;
        RECT 718.950 451.950 721.050 452.400 ;
        RECT 379.950 450.000 403.050 450.600 ;
        RECT 439.950 450.600 442.050 451.050 ;
        RECT 505.950 450.600 508.050 451.050 ;
        RECT 379.950 449.400 402.600 450.000 ;
        RECT 439.950 449.400 508.050 450.600 ;
        RECT 319.950 448.950 324.000 449.100 ;
        RECT 379.950 448.950 382.050 449.400 ;
        RECT 439.950 448.950 442.050 449.400 ;
        RECT 505.950 448.950 508.050 449.400 ;
        RECT 574.950 450.600 577.050 451.050 ;
        RECT 628.950 450.600 631.050 451.050 ;
        RECT 574.950 449.400 631.050 450.600 ;
        RECT 574.950 448.950 577.050 449.400 ;
        RECT 628.950 448.950 631.050 449.400 ;
        RECT 661.950 449.100 664.050 451.200 ;
        RECT 670.950 450.600 673.050 451.050 ;
        RECT 691.950 450.600 694.050 451.050 ;
        RECT 670.950 449.400 694.050 450.600 ;
        RECT 7.950 447.600 10.050 447.900 ;
        RECT -0.600 446.400 10.050 447.600 ;
        RECT 7.950 445.800 10.050 446.400 ;
        RECT 25.950 445.950 28.050 448.050 ;
        RECT 34.950 447.600 37.050 448.050 ;
        RECT 52.950 447.600 55.050 448.050 ;
        RECT 34.950 446.400 55.050 447.600 ;
        RECT 34.950 445.950 37.050 446.400 ;
        RECT 52.950 445.950 55.050 446.400 ;
        RECT 64.950 447.600 67.050 448.050 ;
        RECT 133.950 447.600 136.050 448.050 ;
        RECT 157.950 447.600 160.050 448.050 ;
        RECT 64.950 446.400 160.050 447.600 ;
        RECT 64.950 445.950 67.050 446.400 ;
        RECT 133.950 445.950 136.050 446.400 ;
        RECT 157.950 445.950 160.050 446.400 ;
        RECT 220.950 447.600 223.050 448.050 ;
        RECT 235.950 447.600 238.050 448.050 ;
        RECT 220.950 446.400 238.050 447.600 ;
        RECT 220.950 445.950 223.050 446.400 ;
        RECT 235.950 445.950 238.050 446.400 ;
        RECT 301.950 447.600 304.050 448.050 ;
        RECT 322.950 447.600 325.050 447.900 ;
        RECT 301.950 446.400 325.050 447.600 ;
        RECT 301.950 445.950 304.050 446.400 ;
        RECT 322.950 445.800 325.050 446.400 ;
        RECT 493.950 447.600 496.050 448.050 ;
        RECT 502.950 447.600 505.050 448.050 ;
        RECT 493.950 446.400 505.050 447.600 ;
        RECT 493.950 445.950 496.050 446.400 ;
        RECT 502.950 445.950 505.050 446.400 ;
        RECT 67.950 444.600 70.050 445.050 ;
        RECT 73.950 444.600 76.050 445.050 ;
        RECT 67.950 443.400 76.050 444.600 ;
        RECT 67.950 442.950 70.050 443.400 ;
        RECT 73.950 442.950 76.050 443.400 ;
        RECT 115.950 444.600 118.050 445.050 ;
        RECT 121.950 444.600 124.050 445.050 ;
        RECT 115.950 443.400 124.050 444.600 ;
        RECT 115.950 442.950 118.050 443.400 ;
        RECT 121.950 442.950 124.050 443.400 ;
        RECT 178.950 444.600 181.050 445.200 ;
        RECT 211.950 444.600 214.050 445.050 ;
        RECT 178.950 443.400 214.050 444.600 ;
        RECT 178.950 443.100 181.050 443.400 ;
        RECT 211.950 442.950 214.050 443.400 ;
        RECT 259.950 444.600 262.050 445.050 ;
        RECT 355.950 444.600 358.050 445.050 ;
        RECT 259.950 443.400 358.050 444.600 ;
        RECT 259.950 442.950 262.050 443.400 ;
        RECT 355.950 442.950 358.050 443.400 ;
        RECT 373.950 444.600 376.050 445.050 ;
        RECT 406.950 444.600 409.050 445.050 ;
        RECT 460.950 444.600 463.050 445.050 ;
        RECT 373.950 443.400 463.050 444.600 ;
        RECT 373.950 442.950 376.050 443.400 ;
        RECT 406.950 442.950 409.050 443.400 ;
        RECT 460.950 442.950 463.050 443.400 ;
        RECT 475.950 444.600 478.050 445.050 ;
        RECT 520.950 444.600 523.050 445.050 ;
        RECT 475.950 443.400 523.050 444.600 ;
        RECT 475.950 442.950 478.050 443.400 ;
        RECT 520.950 442.950 523.050 443.400 ;
        RECT 562.950 444.600 565.050 445.050 ;
        RECT 586.950 444.600 589.050 445.050 ;
        RECT 562.950 443.400 589.050 444.600 ;
        RECT 562.950 442.950 565.050 443.400 ;
        RECT 586.950 442.950 589.050 443.400 ;
        RECT 643.950 444.600 646.050 445.050 ;
        RECT 662.400 444.600 663.600 449.100 ;
        RECT 670.950 448.950 673.050 449.400 ;
        RECT 691.950 448.950 694.050 449.400 ;
        RECT 724.950 447.600 727.050 448.050 ;
        RECT 736.950 447.600 739.050 451.050 ;
        RECT 748.950 450.600 751.050 451.050 ;
        RECT 757.950 450.600 760.050 451.050 ;
        RECT 748.950 449.400 760.050 450.600 ;
        RECT 748.950 448.950 751.050 449.400 ;
        RECT 757.950 448.950 760.050 449.400 ;
        RECT 781.950 450.600 784.050 451.050 ;
        RECT 796.950 450.600 799.050 451.050 ;
        RECT 781.950 449.400 799.050 450.600 ;
        RECT 781.950 448.950 784.050 449.400 ;
        RECT 796.950 448.950 799.050 449.400 ;
        RECT 724.950 447.000 739.050 447.600 ;
        RECT 724.950 446.400 738.600 447.000 ;
        RECT 724.950 445.950 727.050 446.400 ;
        RECT 688.950 444.600 691.050 445.050 ;
        RECT 694.950 444.600 697.050 445.050 ;
        RECT 643.950 443.400 697.050 444.600 ;
        RECT 643.950 442.950 646.050 443.400 ;
        RECT 688.950 442.950 691.050 443.400 ;
        RECT 694.950 442.950 697.050 443.400 ;
        RECT 766.950 444.600 769.050 445.050 ;
        RECT 772.950 444.600 775.050 445.050 ;
        RECT 766.950 443.400 775.050 444.600 ;
        RECT 766.950 442.950 769.050 443.400 ;
        RECT 772.950 442.950 775.050 443.400 ;
        RECT 16.950 441.600 19.050 442.050 ;
        RECT 31.950 441.600 34.050 442.050 ;
        RECT 64.950 441.600 67.050 442.050 ;
        RECT 16.950 440.400 67.050 441.600 ;
        RECT 16.950 439.950 19.050 440.400 ;
        RECT 31.950 439.950 34.050 440.400 ;
        RECT 64.950 439.950 67.050 440.400 ;
        RECT 70.950 441.600 73.050 442.050 ;
        RECT 82.950 441.600 85.050 442.050 ;
        RECT 70.950 440.400 85.050 441.600 ;
        RECT 70.950 439.950 73.050 440.400 ;
        RECT 82.950 439.950 85.050 440.400 ;
        RECT 148.950 441.600 151.050 442.050 ;
        RECT 169.950 441.600 172.050 442.050 ;
        RECT 190.950 441.600 193.050 442.050 ;
        RECT 148.950 440.400 193.050 441.600 ;
        RECT 148.950 439.950 151.050 440.400 ;
        RECT 169.950 439.950 172.050 440.400 ;
        RECT 190.950 439.950 193.050 440.400 ;
        RECT 256.950 441.600 259.050 442.050 ;
        RECT 286.950 441.600 289.050 442.050 ;
        RECT 307.950 441.600 310.050 442.050 ;
        RECT 256.950 440.400 310.050 441.600 ;
        RECT 256.950 439.950 259.050 440.400 ;
        RECT 286.950 439.950 289.050 440.400 ;
        RECT 307.950 439.950 310.050 440.400 ;
        RECT 316.950 441.600 319.050 442.050 ;
        RECT 340.950 441.600 343.050 442.050 ;
        RECT 316.950 440.400 343.050 441.600 ;
        RECT 316.950 439.950 319.050 440.400 ;
        RECT 340.950 439.950 343.050 440.400 ;
        RECT 376.950 441.600 379.050 442.050 ;
        RECT 427.950 441.600 430.050 442.050 ;
        RECT 376.950 440.400 430.050 441.600 ;
        RECT 376.950 439.950 379.050 440.400 ;
        RECT 427.950 439.950 430.050 440.400 ;
        RECT 655.950 441.600 658.050 442.050 ;
        RECT 661.950 441.600 664.050 442.050 ;
        RECT 655.950 440.400 664.050 441.600 ;
        RECT 655.950 439.950 658.050 440.400 ;
        RECT 661.950 439.950 664.050 440.400 ;
        RECT 67.950 438.600 70.050 439.050 ;
        RECT 205.950 438.600 208.050 439.050 ;
        RECT 67.950 437.400 208.050 438.600 ;
        RECT 67.950 436.950 70.050 437.400 ;
        RECT 205.950 436.950 208.050 437.400 ;
        RECT 541.950 438.600 544.050 439.050 ;
        RECT 577.950 438.600 580.050 439.050 ;
        RECT 541.950 437.400 580.050 438.600 ;
        RECT 541.950 436.950 544.050 437.400 ;
        RECT 577.950 436.950 580.050 437.400 ;
        RECT 1.950 435.600 4.050 436.050 ;
        RECT 19.950 435.600 22.050 436.050 ;
        RECT 1.950 434.400 22.050 435.600 ;
        RECT 1.950 433.950 4.050 434.400 ;
        RECT 19.950 433.950 22.050 434.400 ;
        RECT 73.950 435.600 76.050 436.050 ;
        RECT 130.950 435.600 133.050 436.050 ;
        RECT 73.950 434.400 133.050 435.600 ;
        RECT 73.950 433.950 76.050 434.400 ;
        RECT 130.950 433.950 133.050 434.400 ;
        RECT 166.950 435.600 169.050 436.050 ;
        RECT 175.950 435.600 178.050 436.050 ;
        RECT 199.950 435.600 202.050 436.050 ;
        RECT 166.950 434.400 202.050 435.600 ;
        RECT 166.950 433.950 169.050 434.400 ;
        RECT 175.950 433.950 178.050 434.400 ;
        RECT 199.950 433.950 202.050 434.400 ;
        RECT 211.950 435.600 214.050 436.050 ;
        RECT 241.950 435.600 244.050 436.050 ;
        RECT 211.950 434.400 244.050 435.600 ;
        RECT 211.950 433.950 214.050 434.400 ;
        RECT 241.950 433.950 244.050 434.400 ;
        RECT 262.950 435.600 265.050 436.050 ;
        RECT 310.950 435.600 313.050 436.050 ;
        RECT 262.950 434.400 313.050 435.600 ;
        RECT 262.950 433.950 265.050 434.400 ;
        RECT 310.950 433.950 313.050 434.400 ;
        RECT 382.950 435.600 385.050 436.050 ;
        RECT 487.950 435.600 490.050 436.050 ;
        RECT 817.950 435.600 820.050 436.050 ;
        RECT 382.950 434.400 490.050 435.600 ;
        RECT 382.950 433.950 385.050 434.400 ;
        RECT 487.950 433.950 490.050 434.400 ;
        RECT 581.400 434.400 820.050 435.600 ;
        RECT 508.950 432.600 511.050 433.050 ;
        RECT 581.400 432.600 582.600 434.400 ;
        RECT 817.950 433.950 820.050 434.400 ;
        RECT 508.950 431.400 582.600 432.600 ;
        RECT 508.950 430.950 511.050 431.400 ;
        RECT 28.950 429.600 31.050 430.050 ;
        RECT 43.950 429.600 46.050 430.050 ;
        RECT 94.950 429.600 97.050 430.050 ;
        RECT 28.950 428.400 97.050 429.600 ;
        RECT 28.950 427.950 31.050 428.400 ;
        RECT 43.950 427.950 46.050 428.400 ;
        RECT 94.950 427.950 97.050 428.400 ;
        RECT 217.950 429.600 220.050 430.050 ;
        RECT 256.950 429.600 259.050 430.200 ;
        RECT 217.950 428.400 259.050 429.600 ;
        RECT 217.950 427.950 220.050 428.400 ;
        RECT 256.950 428.100 259.050 428.400 ;
        RECT 724.950 429.600 727.050 430.050 ;
        RECT 769.950 429.600 772.050 430.050 ;
        RECT 724.950 428.400 772.050 429.600 ;
        RECT 724.950 427.950 727.050 428.400 ;
        RECT 769.950 427.950 772.050 428.400 ;
        RECT 256.950 426.600 259.050 426.900 ;
        RECT 265.950 426.600 268.050 427.050 ;
        RECT 256.950 425.400 268.050 426.600 ;
        RECT 256.950 424.800 259.050 425.400 ;
        RECT 265.950 424.950 268.050 425.400 ;
        RECT 646.950 426.600 649.050 427.050 ;
        RECT 658.950 426.600 661.050 427.050 ;
        RECT 646.950 425.400 661.050 426.600 ;
        RECT 646.950 424.950 649.050 425.400 ;
        RECT 658.950 424.950 661.050 425.400 ;
        RECT 733.950 426.600 736.050 427.050 ;
        RECT 748.950 426.600 751.050 427.050 ;
        RECT 733.950 425.400 751.050 426.600 ;
        RECT 733.950 424.950 736.050 425.400 ;
        RECT 748.950 424.950 751.050 425.400 ;
        RECT 118.950 423.600 121.050 424.050 ;
        RECT 154.950 423.600 157.050 424.050 ;
        RECT 178.950 423.600 181.050 424.050 ;
        RECT 118.950 422.400 181.050 423.600 ;
        RECT 118.950 421.950 121.050 422.400 ;
        RECT 154.950 421.950 157.050 422.400 ;
        RECT 178.950 421.950 181.050 422.400 ;
        RECT 223.950 423.600 226.050 424.050 ;
        RECT 232.950 423.600 235.050 424.050 ;
        RECT 268.950 423.600 271.050 424.050 ;
        RECT 223.950 422.400 271.050 423.600 ;
        RECT 223.950 421.950 226.050 422.400 ;
        RECT 232.950 421.950 235.050 422.400 ;
        RECT 268.950 421.950 271.050 422.400 ;
        RECT 286.950 423.600 289.050 424.050 ;
        RECT 298.950 423.600 301.050 424.050 ;
        RECT 286.950 422.400 301.050 423.600 ;
        RECT 286.950 421.950 289.050 422.400 ;
        RECT 298.950 421.950 301.050 422.400 ;
        RECT 460.950 423.600 463.050 424.050 ;
        RECT 511.950 423.600 514.050 424.050 ;
        RECT 460.950 422.400 514.050 423.600 ;
        RECT 460.950 421.950 463.050 422.400 ;
        RECT 511.950 421.950 514.050 422.400 ;
        RECT 613.950 423.600 616.050 424.050 ;
        RECT 679.950 423.600 682.050 424.050 ;
        RECT 613.950 422.400 682.050 423.600 ;
        RECT 613.950 421.950 616.050 422.400 ;
        RECT 679.950 421.950 682.050 422.400 ;
        RECT 796.950 423.600 799.050 424.050 ;
        RECT 823.950 423.600 826.050 424.050 ;
        RECT 796.950 422.400 826.050 423.600 ;
        RECT 796.950 421.950 799.050 422.400 ;
        RECT 823.950 421.950 826.050 422.400 ;
        RECT 61.950 420.600 64.050 421.200 ;
        RECT 76.950 420.600 79.050 421.050 ;
        RECT 61.950 419.400 79.050 420.600 ;
        RECT 61.950 419.100 64.050 419.400 ;
        RECT 76.950 418.950 79.050 419.400 ;
        RECT 121.950 420.600 124.050 421.050 ;
        RECT 139.950 420.600 142.050 421.200 ;
        RECT 121.950 419.400 142.050 420.600 ;
        RECT 121.950 418.950 124.050 419.400 ;
        RECT 139.950 419.100 142.050 419.400 ;
        RECT 4.950 417.600 7.050 418.050 ;
        RECT 10.950 417.600 13.050 418.050 ;
        RECT 46.950 417.600 49.050 418.050 ;
        RECT 4.950 416.400 49.050 417.600 ;
        RECT 4.950 415.950 7.050 416.400 ;
        RECT 10.950 415.950 13.050 416.400 ;
        RECT 46.950 415.950 49.050 416.400 ;
        RECT 106.950 417.600 109.050 418.050 ;
        RECT 122.400 417.600 123.600 418.950 ;
        RECT 106.950 416.400 123.600 417.600 ;
        RECT 151.950 417.600 154.050 418.050 ;
        RECT 157.950 417.600 160.050 421.050 ;
        RECT 208.950 420.600 211.050 421.050 ;
        RECT 244.950 420.600 247.050 421.200 ;
        RECT 259.950 420.600 262.050 421.050 ;
        RECT 208.950 419.400 262.050 420.600 ;
        RECT 208.950 418.950 211.050 419.400 ;
        RECT 244.950 419.100 247.050 419.400 ;
        RECT 259.950 418.950 262.050 419.400 ;
        RECT 274.950 420.600 277.050 421.050 ;
        RECT 283.950 420.600 286.050 421.050 ;
        RECT 274.950 419.400 286.050 420.600 ;
        RECT 274.950 418.950 277.050 419.400 ;
        RECT 283.950 418.950 286.050 419.400 ;
        RECT 355.950 420.600 358.050 421.050 ;
        RECT 382.950 420.600 385.050 421.050 ;
        RECT 355.950 419.400 385.050 420.600 ;
        RECT 355.950 418.950 358.050 419.400 ;
        RECT 151.950 417.000 160.050 417.600 ;
        RECT 247.950 418.050 250.050 418.200 ;
        RECT 151.950 416.400 159.600 417.000 ;
        RECT 106.950 415.950 109.050 416.400 ;
        RECT 151.950 415.950 154.050 416.400 ;
        RECT 247.950 416.100 253.050 418.050 ;
        RECT 249.000 415.950 253.050 416.100 ;
        RECT 265.950 417.600 268.050 418.050 ;
        RECT 292.950 417.600 295.050 418.050 ;
        RECT 265.950 416.400 295.050 417.600 ;
        RECT 265.950 415.950 268.050 416.400 ;
        RECT 292.950 415.950 295.050 416.400 ;
        RECT 319.950 417.600 322.050 418.050 ;
        RECT 346.950 417.600 349.050 418.050 ;
        RECT 319.950 416.400 349.050 417.600 ;
        RECT 319.950 415.950 322.050 416.400 ;
        RECT 346.950 415.950 349.050 416.400 ;
        RECT 364.950 415.950 367.050 419.400 ;
        RECT 382.950 418.950 385.050 419.400 ;
        RECT 430.950 420.600 433.050 421.050 ;
        RECT 454.950 420.600 457.050 421.200 ;
        RECT 430.950 419.400 457.050 420.600 ;
        RECT 512.400 420.600 513.600 421.950 ;
        RECT 547.950 420.600 550.050 421.050 ;
        RECT 512.400 419.400 550.050 420.600 ;
        RECT 430.950 418.950 433.050 419.400 ;
        RECT 454.950 419.100 457.050 419.400 ;
        RECT 547.950 418.950 550.050 419.400 ;
        RECT 637.950 420.600 640.050 421.050 ;
        RECT 649.950 420.600 652.050 421.050 ;
        RECT 637.950 419.400 652.050 420.600 ;
        RECT 637.950 418.950 640.050 419.400 ;
        RECT 649.950 418.950 652.050 419.400 ;
        RECT 661.950 418.050 664.050 421.050 ;
        RECT 577.950 417.600 580.050 418.050 ;
        RECT 586.950 417.600 589.050 418.050 ;
        RECT 577.950 416.400 589.050 417.600 ;
        RECT 661.950 417.000 667.050 418.050 ;
        RECT 662.400 416.400 667.050 417.000 ;
        RECT 577.950 415.950 580.050 416.400 ;
        RECT 586.950 415.950 589.050 416.400 ;
        RECT 663.000 415.950 667.050 416.400 ;
        RECT 709.950 417.600 712.050 418.050 ;
        RECT 745.950 417.600 748.050 421.050 ;
        RECT 709.950 417.000 748.050 417.600 ;
        RECT 790.950 417.600 793.050 421.050 ;
        RECT 802.950 417.600 805.050 418.050 ;
        RECT 790.950 417.000 805.050 417.600 ;
        RECT 709.950 416.400 747.600 417.000 ;
        RECT 791.400 416.400 805.050 417.000 ;
        RECT 709.950 415.950 712.050 416.400 ;
        RECT 802.950 415.950 805.050 416.400 ;
        RECT 31.950 414.600 34.050 415.050 ;
        RECT 37.950 414.600 40.050 415.050 ;
        RECT 31.950 413.400 40.050 414.600 ;
        RECT 31.950 412.950 34.050 413.400 ;
        RECT 37.950 412.950 40.050 413.400 ;
        RECT 19.950 409.950 25.050 412.050 ;
        RECT 124.950 411.600 127.050 415.050 ;
        RECT 139.950 414.600 142.050 415.050 ;
        RECT 148.950 414.600 151.050 415.050 ;
        RECT 139.950 413.400 151.050 414.600 ;
        RECT 139.950 412.950 142.050 413.400 ;
        RECT 148.950 412.950 151.050 413.400 ;
        RECT 172.950 414.600 175.050 415.050 ;
        RECT 181.950 414.600 184.050 415.050 ;
        RECT 172.950 413.400 184.050 414.600 ;
        RECT 172.950 412.950 175.050 413.400 ;
        RECT 181.950 412.950 184.050 413.400 ;
        RECT 205.950 414.600 208.050 415.200 ;
        RECT 217.800 414.600 219.900 415.050 ;
        RECT 205.950 413.400 219.900 414.600 ;
        RECT 221.100 414.000 223.200 415.050 ;
        RECT 205.950 413.100 208.050 413.400 ;
        RECT 217.800 412.950 219.900 413.400 ;
        RECT 220.950 412.950 223.200 414.000 ;
        RECT 130.950 411.600 133.050 412.050 ;
        RECT 124.950 411.000 133.050 411.600 ;
        RECT 125.400 410.400 133.050 411.000 ;
        RECT 130.950 409.950 133.050 410.400 ;
        RECT 211.950 411.600 214.050 412.050 ;
        RECT 220.950 411.600 223.050 412.950 ;
        RECT 211.950 411.000 223.050 411.600 ;
        RECT 241.950 411.600 244.050 412.050 ;
        RECT 247.950 411.600 250.050 414.900 ;
        RECT 484.950 414.600 487.050 415.050 ;
        RECT 523.950 414.600 526.050 415.050 ;
        RECT 541.950 414.600 544.050 415.050 ;
        RECT 484.950 414.000 507.600 414.600 ;
        RECT 484.950 413.400 508.050 414.000 ;
        RECT 484.950 412.950 487.050 413.400 ;
        RECT 241.950 411.000 250.050 411.600 ;
        RECT 307.950 411.600 310.050 412.050 ;
        RECT 316.950 411.600 319.050 412.050 ;
        RECT 211.950 410.400 222.600 411.000 ;
        RECT 241.950 410.400 249.600 411.000 ;
        RECT 307.950 410.400 319.050 411.600 ;
        RECT 211.950 409.950 214.050 410.400 ;
        RECT 241.950 409.950 244.050 410.400 ;
        RECT 307.950 409.950 310.050 410.400 ;
        RECT 316.950 409.950 319.050 410.400 ;
        RECT 352.950 411.600 355.050 412.050 ;
        RECT 373.950 411.600 376.050 412.050 ;
        RECT 352.950 410.400 376.050 411.600 ;
        RECT 352.950 409.950 355.050 410.400 ;
        RECT 373.950 409.950 376.050 410.400 ;
        RECT 457.950 411.600 460.050 412.050 ;
        RECT 478.950 411.600 481.050 412.050 ;
        RECT 457.950 410.400 481.050 411.600 ;
        RECT 457.950 409.950 460.050 410.400 ;
        RECT 478.950 409.950 481.050 410.400 ;
        RECT 505.950 409.950 508.050 413.400 ;
        RECT 523.950 413.400 544.050 414.600 ;
        RECT 523.950 412.950 526.050 413.400 ;
        RECT 541.950 411.600 544.050 413.400 ;
        RECT 556.950 414.600 559.050 415.050 ;
        RECT 571.950 414.600 574.050 415.050 ;
        RECT 556.950 413.400 574.050 414.600 ;
        RECT 556.950 412.950 559.050 413.400 ;
        RECT 571.950 412.950 574.050 413.400 ;
        RECT 622.950 414.600 625.050 415.050 ;
        RECT 634.950 414.600 637.050 414.900 ;
        RECT 622.950 413.400 637.050 414.600 ;
        RECT 622.950 412.950 625.050 413.400 ;
        RECT 634.950 412.800 637.050 413.400 ;
        RECT 751.950 414.600 754.050 415.050 ;
        RECT 772.950 414.600 775.050 415.050 ;
        RECT 751.950 413.400 775.050 414.600 ;
        RECT 751.950 412.950 754.050 413.400 ;
        RECT 772.950 412.950 775.050 413.400 ;
        RECT 580.950 411.600 583.050 412.050 ;
        RECT 541.950 411.000 583.050 411.600 ;
        RECT 542.400 410.400 583.050 411.000 ;
        RECT 580.950 409.950 583.050 410.400 ;
        RECT 640.950 411.600 643.050 412.050 ;
        RECT 682.950 411.600 685.050 412.050 ;
        RECT 640.950 410.400 685.050 411.600 ;
        RECT 640.950 409.950 643.050 410.400 ;
        RECT 682.950 409.950 685.050 410.400 ;
        RECT 718.950 409.950 724.050 412.050 ;
        RECT 730.950 411.600 733.050 412.050 ;
        RECT 745.950 411.600 748.050 412.050 ;
        RECT 730.950 410.400 748.050 411.600 ;
        RECT 730.950 409.950 733.050 410.400 ;
        RECT 745.950 409.950 748.050 410.400 ;
        RECT 31.950 405.600 34.050 406.050 ;
        RECT 46.950 405.600 49.050 406.050 ;
        RECT 31.950 404.400 49.050 405.600 ;
        RECT 31.950 403.950 34.050 404.400 ;
        RECT 46.950 403.950 49.050 404.400 ;
        RECT 70.950 405.600 73.050 406.050 ;
        RECT 85.950 405.600 88.050 406.050 ;
        RECT 70.950 404.400 88.050 405.600 ;
        RECT 106.950 405.600 109.050 409.050 ;
        RECT 259.950 408.600 262.050 409.050 ;
        RECT 298.950 408.600 301.050 409.050 ;
        RECT 259.950 407.400 301.050 408.600 ;
        RECT 259.950 406.950 262.050 407.400 ;
        RECT 298.950 406.950 301.050 407.400 ;
        RECT 487.950 408.600 490.050 409.050 ;
        RECT 538.950 408.600 541.050 409.050 ;
        RECT 544.950 408.600 547.050 409.050 ;
        RECT 487.950 407.400 547.050 408.600 ;
        RECT 487.950 406.950 490.050 407.400 ;
        RECT 538.950 406.950 541.050 407.400 ;
        RECT 544.950 406.950 547.050 407.400 ;
        RECT 706.950 408.600 709.050 409.050 ;
        RECT 754.950 408.600 757.050 409.050 ;
        RECT 706.950 407.400 757.050 408.600 ;
        RECT 706.950 406.950 709.050 407.400 ;
        RECT 754.950 406.950 757.050 407.400 ;
        RECT 124.950 405.600 127.050 406.050 ;
        RECT 106.950 405.000 127.050 405.600 ;
        RECT 107.400 404.400 127.050 405.000 ;
        RECT 70.950 403.950 73.050 404.400 ;
        RECT 85.950 403.950 88.050 404.400 ;
        RECT 124.950 403.950 127.050 404.400 ;
        RECT 292.950 405.600 295.050 406.050 ;
        RECT 301.950 405.600 304.050 406.050 ;
        RECT 322.950 405.600 325.050 406.050 ;
        RECT 292.950 404.400 325.050 405.600 ;
        RECT 292.950 403.950 295.050 404.400 ;
        RECT 301.950 403.950 304.050 404.400 ;
        RECT 322.950 403.950 325.050 404.400 ;
        RECT 760.950 405.600 763.050 406.050 ;
        RECT 781.950 405.600 784.050 406.050 ;
        RECT 802.950 405.600 805.050 406.050 ;
        RECT 760.950 404.400 805.050 405.600 ;
        RECT 760.950 403.950 763.050 404.400 ;
        RECT 781.950 403.950 784.050 404.400 ;
        RECT 802.950 403.950 805.050 404.400 ;
        RECT 814.950 405.600 817.050 406.050 ;
        RECT 823.950 405.600 826.050 406.050 ;
        RECT 814.950 404.400 826.050 405.600 ;
        RECT 814.950 403.950 817.050 404.400 ;
        RECT 823.950 403.950 826.050 404.400 ;
        RECT 406.950 402.600 409.050 403.050 ;
        RECT 412.950 402.600 415.050 403.050 ;
        RECT 424.950 402.600 427.050 403.050 ;
        RECT 433.950 402.600 436.050 403.050 ;
        RECT 406.950 401.400 436.050 402.600 ;
        RECT 406.950 400.950 409.050 401.400 ;
        RECT 412.950 400.950 415.050 401.400 ;
        RECT 424.950 400.950 427.050 401.400 ;
        RECT 433.950 400.950 436.050 401.400 ;
        RECT 451.950 399.600 454.050 400.050 ;
        RECT 490.950 399.600 493.050 400.050 ;
        RECT 511.950 399.600 514.050 400.050 ;
        RECT 574.950 399.600 577.050 400.050 ;
        RECT 451.950 398.400 577.050 399.600 ;
        RECT 451.950 397.950 454.050 398.400 ;
        RECT 490.950 397.950 493.050 398.400 ;
        RECT 511.950 397.950 514.050 398.400 ;
        RECT 574.950 397.950 577.050 398.400 ;
        RECT 643.950 399.600 646.050 400.050 ;
        RECT 682.950 399.600 685.050 400.050 ;
        RECT 709.950 399.600 712.050 400.050 ;
        RECT 793.950 399.600 796.050 400.050 ;
        RECT 805.950 399.600 808.050 400.050 ;
        RECT 817.950 399.600 820.050 400.050 ;
        RECT 643.950 398.400 820.050 399.600 ;
        RECT 643.950 397.950 646.050 398.400 ;
        RECT 682.950 397.950 685.050 398.400 ;
        RECT 709.950 397.950 712.050 398.400 ;
        RECT 793.950 397.950 796.050 398.400 ;
        RECT 805.950 397.950 808.050 398.400 ;
        RECT 817.950 397.950 820.050 398.400 ;
        RECT 367.950 396.600 370.050 397.050 ;
        RECT 469.950 396.600 472.050 397.050 ;
        RECT 367.950 395.400 472.050 396.600 ;
        RECT 367.950 394.950 370.050 395.400 ;
        RECT 469.950 394.950 472.050 395.400 ;
        RECT 607.950 396.600 610.050 397.050 ;
        RECT 622.950 396.600 625.050 397.050 ;
        RECT 607.950 395.400 625.050 396.600 ;
        RECT 607.950 394.950 610.050 395.400 ;
        RECT 622.950 394.950 625.050 395.400 ;
        RECT 73.950 393.600 76.050 394.050 ;
        RECT 82.950 393.600 85.050 394.050 ;
        RECT 73.950 392.400 85.050 393.600 ;
        RECT 73.950 391.950 76.050 392.400 ;
        RECT 82.950 391.950 85.050 392.400 ;
        RECT 139.950 393.600 142.050 394.050 ;
        RECT 190.950 393.600 193.050 394.050 ;
        RECT 139.950 392.400 193.050 393.600 ;
        RECT 139.950 391.950 142.050 392.400 ;
        RECT 190.950 391.950 193.050 392.400 ;
        RECT 199.950 393.600 202.050 394.050 ;
        RECT 241.950 393.600 244.050 394.050 ;
        RECT 199.950 392.400 244.050 393.600 ;
        RECT 199.950 391.950 202.050 392.400 ;
        RECT 241.950 391.950 244.050 392.400 ;
        RECT 691.950 393.600 694.050 394.050 ;
        RECT 742.950 393.600 745.050 394.050 ;
        RECT 691.950 392.400 745.050 393.600 ;
        RECT 691.950 391.950 694.050 392.400 ;
        RECT 742.950 391.950 745.050 392.400 ;
        RECT 808.950 393.600 811.050 394.050 ;
        RECT 826.950 393.600 829.050 394.050 ;
        RECT 808.950 392.400 829.050 393.600 ;
        RECT 808.950 391.950 811.050 392.400 ;
        RECT 826.950 391.950 829.050 392.400 ;
        RECT 64.950 390.600 67.050 391.050 ;
        RECT 79.950 390.600 82.050 391.050 ;
        RECT 64.950 389.400 82.050 390.600 ;
        RECT 64.950 388.950 67.050 389.400 ;
        RECT 79.950 388.950 82.050 389.400 ;
        RECT 121.950 390.600 124.050 391.050 ;
        RECT 202.950 390.600 205.050 391.050 ;
        RECT 121.950 389.400 205.050 390.600 ;
        RECT 121.950 388.950 124.050 389.400 ;
        RECT 202.950 388.950 205.050 389.400 ;
        RECT 658.950 390.600 661.050 391.050 ;
        RECT 730.950 390.600 733.050 391.050 ;
        RECT 658.950 389.400 733.050 390.600 ;
        RECT 658.950 388.950 661.050 389.400 ;
        RECT 730.950 388.950 733.050 389.400 ;
        RECT 784.950 390.600 787.050 391.050 ;
        RECT 802.950 390.600 805.050 391.050 ;
        RECT 784.950 389.400 805.050 390.600 ;
        RECT 784.950 388.950 787.050 389.400 ;
        RECT 802.950 388.950 805.050 389.400 ;
        RECT 88.950 387.600 91.050 388.050 ;
        RECT 103.950 387.600 106.050 388.050 ;
        RECT 145.950 387.600 148.050 388.050 ;
        RECT 88.950 386.400 148.050 387.600 ;
        RECT 88.950 385.950 91.050 386.400 ;
        RECT 103.950 385.950 106.050 386.400 ;
        RECT 145.950 385.950 148.050 386.400 ;
        RECT 688.950 387.600 691.050 388.050 ;
        RECT 700.950 387.600 703.050 388.050 ;
        RECT 688.950 386.400 703.050 387.600 ;
        RECT 688.950 385.950 691.050 386.400 ;
        RECT 700.950 385.950 703.050 386.400 ;
        RECT 727.950 387.600 730.050 388.050 ;
        RECT 739.950 387.600 742.050 388.050 ;
        RECT 727.950 386.400 742.050 387.600 ;
        RECT 727.950 385.950 730.050 386.400 ;
        RECT 739.950 385.950 742.050 386.400 ;
        RECT 772.950 387.600 775.050 388.050 ;
        RECT 811.950 387.600 814.050 388.050 ;
        RECT 772.950 386.400 814.050 387.600 ;
        RECT 772.950 385.950 775.050 386.400 ;
        RECT 811.950 385.950 814.050 386.400 ;
        RECT 202.950 384.600 205.050 385.050 ;
        RECT 244.950 384.600 247.050 385.050 ;
        RECT 202.950 383.400 247.050 384.600 ;
        RECT 202.950 382.950 205.050 383.400 ;
        RECT 244.950 382.950 247.050 383.400 ;
        RECT 469.950 384.600 472.050 385.050 ;
        RECT 646.950 384.600 649.050 385.050 ;
        RECT 469.950 383.400 649.050 384.600 ;
        RECT 469.950 382.950 472.050 383.400 ;
        RECT 646.950 382.950 649.050 383.400 ;
        RECT 34.950 381.600 37.050 382.050 ;
        RECT 40.950 381.600 43.050 382.200 ;
        RECT 34.950 380.400 43.050 381.600 ;
        RECT 34.950 379.950 37.050 380.400 ;
        RECT 40.950 380.100 43.050 380.400 ;
        RECT 82.950 381.600 85.050 382.050 ;
        RECT 109.950 381.600 112.050 382.050 ;
        RECT 82.950 380.400 112.050 381.600 ;
        RECT 82.950 379.950 85.050 380.400 ;
        RECT 109.950 379.950 112.050 380.400 ;
        RECT 160.950 381.600 163.050 382.050 ;
        RECT 292.950 381.600 295.050 382.050 ;
        RECT 160.950 380.400 295.050 381.600 ;
        RECT 160.950 379.950 163.050 380.400 ;
        RECT 292.950 379.950 295.050 380.400 ;
        RECT 790.950 381.600 793.050 382.050 ;
        RECT 802.950 381.600 805.050 382.050 ;
        RECT 811.950 381.600 814.050 382.050 ;
        RECT 790.950 380.400 814.050 381.600 ;
        RECT 790.950 379.950 793.050 380.400 ;
        RECT 802.950 379.950 805.050 380.400 ;
        RECT 811.950 379.950 814.050 380.400 ;
        RECT 70.950 378.600 73.050 379.050 ;
        RECT 97.950 378.600 100.050 379.050 ;
        RECT 70.950 377.400 100.050 378.600 ;
        RECT 70.950 376.950 73.050 377.400 ;
        RECT 97.950 376.950 100.050 377.400 ;
        RECT 112.950 378.600 115.050 379.200 ;
        RECT 118.950 378.600 121.050 379.050 ;
        RECT 169.950 378.600 172.050 379.050 ;
        RECT 112.950 377.400 172.050 378.600 ;
        RECT 112.950 377.100 115.050 377.400 ;
        RECT 118.950 376.950 121.050 377.400 ;
        RECT 169.950 376.950 172.050 377.400 ;
        RECT 493.950 378.600 496.050 379.050 ;
        RECT 529.950 378.600 532.050 379.050 ;
        RECT 568.950 378.600 571.050 379.050 ;
        RECT 592.950 378.600 595.050 379.050 ;
        RECT 610.950 378.600 613.050 379.050 ;
        RECT 493.950 377.400 613.050 378.600 ;
        RECT 493.950 376.950 496.050 377.400 ;
        RECT 529.950 376.950 532.050 377.400 ;
        RECT 568.950 376.950 571.050 377.400 ;
        RECT 592.950 376.950 595.050 377.400 ;
        RECT 610.950 376.950 613.050 377.400 ;
        RECT 664.950 378.600 667.050 379.050 ;
        RECT 670.950 378.600 673.050 379.050 ;
        RECT 754.950 378.600 757.050 379.050 ;
        RECT 778.950 378.600 781.050 379.050 ;
        RECT 664.950 377.400 673.050 378.600 ;
        RECT 664.950 376.950 667.050 377.400 ;
        RECT 670.950 376.950 673.050 377.400 ;
        RECT 695.400 377.400 781.050 378.600 ;
        RECT 13.950 375.600 16.050 376.050 ;
        RECT 40.950 375.600 43.050 376.050 ;
        RECT 13.950 374.400 43.050 375.600 ;
        RECT 13.950 373.950 16.050 374.400 ;
        RECT 40.950 373.950 43.050 374.400 ;
        RECT 22.950 372.600 25.050 373.050 ;
        RECT 37.950 372.600 40.050 373.050 ;
        RECT 22.950 371.400 40.050 372.600 ;
        RECT 22.950 370.950 25.050 371.400 ;
        RECT 37.950 370.950 40.050 371.400 ;
        RECT 94.950 372.600 97.050 373.050 ;
        RECT 106.950 372.600 109.050 376.050 ;
        RECT 112.950 375.600 115.050 375.900 ;
        RECT 133.950 375.600 136.050 376.050 ;
        RECT 112.950 374.400 136.050 375.600 ;
        RECT 112.950 373.800 115.050 374.400 ;
        RECT 133.950 373.950 136.050 374.400 ;
        RECT 178.950 375.600 181.050 376.050 ;
        RECT 214.950 375.600 217.050 376.050 ;
        RECT 178.950 374.400 217.050 375.600 ;
        RECT 178.950 373.950 181.050 374.400 ;
        RECT 214.950 373.950 217.050 374.400 ;
        RECT 235.950 375.600 238.050 376.050 ;
        RECT 265.950 375.600 268.050 376.050 ;
        RECT 235.950 374.400 268.050 375.600 ;
        RECT 235.950 373.950 238.050 374.400 ;
        RECT 265.950 373.950 268.050 374.400 ;
        RECT 310.950 375.600 313.050 376.050 ;
        RECT 379.950 375.600 382.050 376.050 ;
        RECT 310.950 374.400 382.050 375.600 ;
        RECT 310.950 373.950 313.050 374.400 ;
        RECT 379.950 373.950 382.050 374.400 ;
        RECT 424.950 375.600 427.050 376.050 ;
        RECT 430.950 375.600 433.050 376.050 ;
        RECT 424.950 374.400 433.050 375.600 ;
        RECT 424.950 373.950 427.050 374.400 ;
        RECT 430.950 373.950 433.050 374.400 ;
        RECT 625.950 375.600 628.050 376.050 ;
        RECT 637.950 375.600 640.050 376.050 ;
        RECT 625.950 374.400 640.050 375.600 ;
        RECT 625.950 373.950 628.050 374.400 ;
        RECT 637.950 373.950 640.050 374.400 ;
        RECT 679.950 375.600 682.050 376.200 ;
        RECT 695.400 376.050 696.600 377.400 ;
        RECT 754.950 376.950 757.050 377.400 ;
        RECT 778.950 376.950 781.050 377.400 ;
        RECT 799.950 376.050 802.050 376.200 ;
        RECT 694.950 375.600 697.050 376.050 ;
        RECT 679.950 374.400 697.050 375.600 ;
        RECT 679.950 374.100 682.050 374.400 ;
        RECT 694.950 373.950 697.050 374.400 ;
        RECT 712.950 375.600 715.050 376.050 ;
        RECT 721.950 375.600 724.050 376.050 ;
        RECT 798.000 375.600 802.050 376.050 ;
        RECT 712.950 374.400 724.050 375.600 ;
        RECT 797.400 375.000 802.050 375.600 ;
        RECT 712.950 373.950 715.050 374.400 ;
        RECT 721.950 373.950 724.050 374.400 ;
        RECT 796.950 374.100 802.050 375.000 ;
        RECT 814.950 375.600 817.050 376.050 ;
        RECT 820.950 375.600 823.050 376.050 ;
        RECT 814.950 374.400 823.050 375.600 ;
        RECT 796.950 373.950 801.000 374.100 ;
        RECT 814.950 373.950 817.050 374.400 ;
        RECT 820.950 373.950 823.050 374.400 ;
        RECT 94.950 372.000 109.050 372.600 ;
        RECT 205.950 372.600 208.050 373.050 ;
        RECT 211.950 372.600 214.050 373.050 ;
        RECT 94.950 371.400 108.600 372.000 ;
        RECT 205.950 371.400 214.050 372.600 ;
        RECT 94.950 370.950 97.050 371.400 ;
        RECT 205.950 370.950 208.050 371.400 ;
        RECT 211.950 370.950 214.050 371.400 ;
        RECT 292.950 372.600 295.050 373.050 ;
        RECT 352.950 372.600 355.050 373.050 ;
        RECT 292.950 371.400 355.050 372.600 ;
        RECT 292.950 370.950 295.050 371.400 ;
        RECT 352.950 370.950 355.050 371.400 ;
        RECT 415.950 372.600 418.050 373.050 ;
        RECT 442.950 372.600 445.050 373.050 ;
        RECT 415.950 371.400 445.050 372.600 ;
        RECT 415.950 370.950 418.050 371.400 ;
        RECT 442.950 370.950 445.050 371.400 ;
        RECT 472.950 372.600 475.050 373.050 ;
        RECT 490.950 372.600 493.050 373.050 ;
        RECT 472.950 371.400 493.050 372.600 ;
        RECT 472.950 370.950 475.050 371.400 ;
        RECT 490.950 370.950 493.050 371.400 ;
        RECT 640.950 370.950 646.050 373.050 ;
        RECT 673.950 372.600 676.050 373.050 ;
        RECT 679.950 372.600 682.050 372.900 ;
        RECT 673.950 371.400 682.050 372.600 ;
        RECT 673.950 370.950 676.050 371.400 ;
        RECT 679.950 370.800 682.050 371.400 ;
        RECT 796.950 370.950 799.050 373.950 ;
        RECT 40.950 369.600 43.050 370.050 ;
        RECT 52.950 369.600 55.050 370.050 ;
        RECT 61.950 369.600 64.050 370.050 ;
        RECT 40.950 368.400 64.050 369.600 ;
        RECT 40.950 367.950 43.050 368.400 ;
        RECT 52.950 367.950 55.050 368.400 ;
        RECT 61.950 367.950 64.050 368.400 ;
        RECT 19.950 366.600 22.050 367.050 ;
        RECT 34.950 366.600 37.050 367.050 ;
        RECT 19.950 365.400 37.050 366.600 ;
        RECT 19.950 364.950 22.050 365.400 ;
        RECT 34.950 364.950 37.050 365.400 ;
        RECT 55.950 366.600 58.050 367.050 ;
        RECT 76.950 366.600 79.050 370.050 ;
        RECT 127.950 369.600 130.050 370.050 ;
        RECT 133.950 369.600 136.050 370.050 ;
        RECT 127.950 368.400 136.050 369.600 ;
        RECT 127.950 367.950 130.050 368.400 ;
        RECT 133.950 367.950 136.050 368.400 ;
        RECT 142.950 369.600 145.050 370.050 ;
        RECT 175.950 369.600 178.050 370.050 ;
        RECT 193.950 369.600 196.050 370.050 ;
        RECT 223.950 369.600 226.050 370.050 ;
        RECT 241.950 369.600 244.050 370.050 ;
        RECT 268.950 369.600 271.050 370.050 ;
        RECT 142.950 368.400 271.050 369.600 ;
        RECT 142.950 367.950 145.050 368.400 ;
        RECT 175.950 367.950 178.050 368.400 ;
        RECT 193.950 367.950 196.050 368.400 ;
        RECT 223.950 367.950 226.050 368.400 ;
        RECT 241.950 367.950 244.050 368.400 ;
        RECT 268.950 367.950 271.050 368.400 ;
        RECT 379.950 369.600 382.050 370.050 ;
        RECT 400.950 369.600 403.050 370.050 ;
        RECT 379.950 368.400 403.050 369.600 ;
        RECT 379.950 367.950 382.050 368.400 ;
        RECT 400.950 367.950 403.050 368.400 ;
        RECT 433.950 369.600 436.050 370.050 ;
        RECT 454.950 369.600 457.050 370.050 ;
        RECT 463.950 369.600 466.050 370.050 ;
        RECT 433.950 368.400 466.050 369.600 ;
        RECT 433.950 367.950 436.050 368.400 ;
        RECT 454.950 367.950 457.050 368.400 ;
        RECT 463.950 367.950 466.050 368.400 ;
        RECT 55.950 366.000 79.050 366.600 ;
        RECT 88.950 366.600 91.050 367.050 ;
        RECT 94.950 366.600 97.050 367.050 ;
        RECT 55.950 365.400 78.600 366.000 ;
        RECT 88.950 365.400 97.050 366.600 ;
        RECT 55.950 364.950 58.050 365.400 ;
        RECT 88.950 364.950 91.050 365.400 ;
        RECT 94.950 364.950 97.050 365.400 ;
        RECT 208.950 364.950 214.050 367.050 ;
        RECT 292.950 366.600 295.050 367.050 ;
        RECT 343.950 366.600 346.050 367.050 ;
        RECT 292.950 365.400 346.050 366.600 ;
        RECT 292.950 364.950 295.050 365.400 ;
        RECT 343.950 364.950 346.050 365.400 ;
        RECT 385.950 366.600 388.050 367.050 ;
        RECT 436.950 366.600 439.050 367.050 ;
        RECT 385.950 365.400 439.050 366.600 ;
        RECT 385.950 364.950 388.050 365.400 ;
        RECT 436.950 364.950 439.050 365.400 ;
        RECT 496.950 366.600 499.050 367.050 ;
        RECT 496.950 366.000 507.600 366.600 ;
        RECT 496.950 365.400 508.050 366.000 ;
        RECT 496.950 364.950 499.050 365.400 ;
        RECT 196.950 363.600 199.050 364.050 ;
        RECT 205.950 363.600 208.050 364.050 ;
        RECT 196.950 362.400 208.050 363.600 ;
        RECT 196.950 361.950 199.050 362.400 ;
        RECT 205.950 361.950 208.050 362.400 ;
        RECT 316.950 363.600 319.050 364.050 ;
        RECT 331.950 363.600 334.050 364.050 ;
        RECT 316.950 362.400 334.050 363.600 ;
        RECT 316.950 361.950 319.050 362.400 ;
        RECT 331.950 361.950 334.050 362.400 ;
        RECT 346.950 363.600 349.050 364.050 ;
        RECT 460.950 363.600 463.050 364.050 ;
        RECT 346.950 362.400 463.050 363.600 ;
        RECT 346.950 361.950 349.050 362.400 ;
        RECT 460.950 361.950 463.050 362.400 ;
        RECT 505.950 361.950 508.050 365.400 ;
        RECT 544.950 364.950 550.050 367.050 ;
        RECT 556.950 366.600 559.050 367.050 ;
        RECT 576.000 366.600 580.050 367.050 ;
        RECT 556.950 365.400 580.050 366.600 ;
        RECT 634.950 366.600 637.050 370.050 ;
        RECT 664.950 366.600 667.050 367.050 ;
        RECT 634.950 366.000 667.050 366.600 ;
        RECT 635.400 365.400 667.050 366.000 ;
        RECT 556.950 364.950 559.050 365.400 ;
        RECT 574.950 364.950 580.050 365.400 ;
        RECT 664.950 364.950 667.050 365.400 ;
        RECT 712.950 366.600 715.050 367.200 ;
        RECT 724.950 366.600 727.050 370.050 ;
        RECT 730.950 366.600 733.050 367.050 ;
        RECT 712.950 365.400 733.050 366.600 ;
        RECT 712.950 365.100 715.050 365.400 ;
        RECT 730.950 364.950 733.050 365.400 ;
        RECT 748.950 366.600 751.050 367.050 ;
        RECT 814.950 366.600 817.050 370.050 ;
        RECT 748.950 366.000 817.050 366.600 ;
        RECT 748.950 365.400 816.600 366.000 ;
        RECT 748.950 364.950 751.050 365.400 ;
        RECT 574.950 361.950 577.050 364.950 ;
        RECT 589.950 363.600 592.050 364.050 ;
        RECT 610.950 363.600 613.050 364.050 ;
        RECT 589.950 362.400 613.050 363.600 ;
        RECT 589.950 361.950 592.050 362.400 ;
        RECT 610.950 361.950 613.050 362.400 ;
        RECT 706.950 363.600 709.050 364.050 ;
        RECT 712.950 363.600 715.050 363.900 ;
        RECT 706.950 362.400 715.050 363.600 ;
        RECT 706.950 361.950 709.050 362.400 ;
        RECT 712.950 361.800 715.050 362.400 ;
        RECT 73.950 360.600 76.050 361.050 ;
        RECT 82.950 360.600 85.050 361.050 ;
        RECT 73.950 359.400 85.050 360.600 ;
        RECT 73.950 358.950 76.050 359.400 ;
        RECT 82.950 358.950 85.050 359.400 ;
        RECT 286.950 360.600 289.050 361.050 ;
        RECT 295.950 360.600 298.050 361.050 ;
        RECT 286.950 359.400 298.050 360.600 ;
        RECT 286.950 358.950 289.050 359.400 ;
        RECT 295.950 358.950 298.050 359.400 ;
        RECT 397.950 360.600 400.050 361.050 ;
        RECT 421.800 360.600 423.900 361.050 ;
        RECT 397.950 359.400 423.900 360.600 ;
        RECT 397.950 358.950 400.050 359.400 ;
        RECT 421.800 358.950 423.900 359.400 ;
        RECT 425.100 360.600 427.200 361.050 ;
        RECT 442.950 360.600 445.050 361.050 ;
        RECT 425.100 359.400 445.050 360.600 ;
        RECT 425.100 358.950 427.200 359.400 ;
        RECT 442.950 358.950 445.050 359.400 ;
        RECT 769.950 360.600 772.050 361.050 ;
        RECT 802.950 360.600 805.050 361.050 ;
        RECT 769.950 359.400 805.050 360.600 ;
        RECT 769.950 358.950 772.050 359.400 ;
        RECT 802.950 358.950 805.050 359.400 ;
        RECT 37.950 357.600 40.050 358.050 ;
        RECT 187.950 357.600 190.050 358.050 ;
        RECT 37.950 356.400 190.050 357.600 ;
        RECT 37.950 355.950 40.050 356.400 ;
        RECT 187.950 355.950 190.050 356.400 ;
        RECT 598.950 357.600 601.050 358.050 ;
        RECT 685.950 357.600 688.050 358.050 ;
        RECT 598.950 356.400 688.050 357.600 ;
        RECT 598.950 355.950 601.050 356.400 ;
        RECT 685.950 355.950 688.050 356.400 ;
        RECT 49.950 354.600 52.050 355.050 ;
        RECT 58.950 354.600 61.050 355.050 ;
        RECT 49.950 353.400 61.050 354.600 ;
        RECT 49.950 352.950 52.050 353.400 ;
        RECT 58.950 352.950 61.050 353.400 ;
        RECT 97.950 354.600 100.050 355.050 ;
        RECT 286.950 354.600 289.050 355.050 ;
        RECT 97.950 353.400 289.050 354.600 ;
        RECT 97.950 352.950 100.050 353.400 ;
        RECT 286.950 352.950 289.050 353.400 ;
        RECT 460.950 354.600 463.050 355.050 ;
        RECT 484.950 354.600 487.050 355.050 ;
        RECT 460.950 353.400 487.050 354.600 ;
        RECT 460.950 352.950 463.050 353.400 ;
        RECT 484.950 352.950 487.050 353.400 ;
        RECT 709.950 354.600 712.050 355.050 ;
        RECT 772.950 354.600 775.050 355.050 ;
        RECT 709.950 353.400 775.050 354.600 ;
        RECT 709.950 352.950 712.050 353.400 ;
        RECT 772.950 352.950 775.050 353.400 ;
        RECT 100.950 351.600 103.050 352.050 ;
        RECT 151.950 351.600 154.050 352.050 ;
        RECT 214.950 351.600 217.050 352.050 ;
        RECT 232.950 351.600 235.050 352.050 ;
        RECT 100.950 350.400 183.600 351.600 ;
        RECT 100.950 349.950 103.050 350.400 ;
        RECT 151.950 349.950 154.050 350.400 ;
        RECT 182.400 348.600 183.600 350.400 ;
        RECT 214.950 350.400 235.050 351.600 ;
        RECT 214.950 349.950 217.050 350.400 ;
        RECT 232.950 349.950 235.050 350.400 ;
        RECT 298.950 351.600 301.050 352.050 ;
        RECT 310.950 351.600 313.050 352.050 ;
        RECT 298.950 350.400 313.050 351.600 ;
        RECT 298.950 349.950 301.050 350.400 ;
        RECT 310.950 349.950 313.050 350.400 ;
        RECT 325.950 351.600 328.050 352.050 ;
        RECT 361.950 351.600 364.050 352.050 ;
        RECT 325.950 350.400 364.050 351.600 ;
        RECT 325.950 349.950 328.050 350.400 ;
        RECT 361.950 349.950 364.050 350.400 ;
        RECT 382.950 351.600 385.050 352.050 ;
        RECT 388.950 351.600 391.050 352.050 ;
        RECT 382.950 350.400 391.050 351.600 ;
        RECT 382.950 349.950 385.050 350.400 ;
        RECT 388.950 349.950 391.050 350.400 ;
        RECT 466.950 351.600 469.050 352.050 ;
        RECT 478.950 351.600 481.050 352.050 ;
        RECT 679.950 351.600 682.050 352.050 ;
        RECT 466.950 350.400 481.050 351.600 ;
        RECT 466.950 349.950 469.050 350.400 ;
        RECT 478.950 349.950 481.050 350.400 ;
        RECT 599.400 350.400 682.050 351.600 ;
        RECT 599.400 349.050 600.600 350.400 ;
        RECT 679.950 349.950 682.050 350.400 ;
        RECT 703.950 351.600 706.050 352.050 ;
        RECT 730.950 351.600 733.050 352.050 ;
        RECT 703.950 350.400 733.050 351.600 ;
        RECT 703.950 349.950 706.050 350.400 ;
        RECT 730.950 349.950 733.050 350.400 ;
        RECT 754.950 351.600 757.050 352.050 ;
        RECT 766.950 351.600 769.050 352.050 ;
        RECT 754.950 350.400 769.050 351.600 ;
        RECT 754.950 349.950 757.050 350.400 ;
        RECT 766.950 349.950 769.050 350.400 ;
        RECT 349.950 348.600 352.050 349.050 ;
        RECT 182.400 347.400 352.050 348.600 ;
        RECT 349.950 346.950 352.050 347.400 ;
        RECT 571.950 348.600 574.050 349.050 ;
        RECT 598.950 348.600 601.050 349.050 ;
        RECT 571.950 347.400 601.050 348.600 ;
        RECT 571.950 346.950 574.050 347.400 ;
        RECT 598.950 346.950 601.050 347.400 ;
        RECT 784.950 348.600 787.050 349.050 ;
        RECT 799.950 348.600 802.050 349.050 ;
        RECT 784.950 347.400 802.050 348.600 ;
        RECT 784.950 346.950 787.050 347.400 ;
        RECT 799.950 346.950 802.050 347.400 ;
        RECT 178.950 345.600 181.050 346.050 ;
        RECT 355.950 345.600 358.050 346.050 ;
        RECT 367.950 345.600 370.050 346.050 ;
        RECT 178.950 344.400 370.050 345.600 ;
        RECT 178.950 343.950 181.050 344.400 ;
        RECT 355.950 343.950 358.050 344.400 ;
        RECT 367.950 343.950 370.050 344.400 ;
        RECT 454.950 345.600 457.050 346.050 ;
        RECT 466.950 345.600 469.050 346.050 ;
        RECT 454.950 344.400 469.050 345.600 ;
        RECT 454.950 343.950 457.050 344.400 ;
        RECT 466.950 343.950 469.050 344.400 ;
        RECT 496.950 345.600 499.050 346.050 ;
        RECT 631.950 345.600 634.050 346.050 ;
        RECT 496.950 344.400 634.050 345.600 ;
        RECT 496.950 343.950 499.050 344.400 ;
        RECT 631.950 343.950 634.050 344.400 ;
        RECT 652.950 345.600 655.050 346.050 ;
        RECT 736.950 345.600 739.050 346.050 ;
        RECT 652.950 344.400 739.050 345.600 ;
        RECT 652.950 343.950 655.050 344.400 ;
        RECT 736.950 343.950 739.050 344.400 ;
        RECT 796.950 345.600 799.050 346.050 ;
        RECT 811.950 345.600 814.050 346.050 ;
        RECT 796.950 344.400 814.050 345.600 ;
        RECT 796.950 343.950 799.050 344.400 ;
        RECT 811.950 343.950 814.050 344.400 ;
        RECT 7.950 342.600 10.050 343.050 ;
        RECT 46.950 342.600 49.050 343.050 ;
        RECT 58.950 342.600 61.050 343.050 ;
        RECT 7.950 341.400 61.050 342.600 ;
        RECT 7.950 340.950 10.050 341.400 ;
        RECT 46.950 340.950 49.050 341.400 ;
        RECT 58.950 340.950 61.050 341.400 ;
        RECT 103.950 342.600 106.050 343.050 ;
        RECT 112.950 342.600 115.050 343.050 ;
        RECT 103.950 341.400 115.050 342.600 ;
        RECT 103.950 340.950 106.050 341.400 ;
        RECT 112.950 340.950 115.050 341.400 ;
        RECT 421.950 342.600 424.050 343.050 ;
        RECT 445.950 342.600 448.050 343.050 ;
        RECT 421.950 341.400 448.050 342.600 ;
        RECT 421.950 340.950 424.050 341.400 ;
        RECT 445.950 340.950 448.050 341.400 ;
        RECT 523.950 342.600 526.050 343.050 ;
        RECT 529.950 342.600 532.050 343.050 ;
        RECT 523.950 341.400 532.050 342.600 ;
        RECT 523.950 340.950 526.050 341.400 ;
        RECT 529.950 340.950 532.050 341.400 ;
        RECT 562.950 342.600 565.050 343.050 ;
        RECT 592.950 342.600 595.050 343.050 ;
        RECT 562.950 341.400 595.050 342.600 ;
        RECT 562.950 340.950 565.050 341.400 ;
        RECT 592.950 340.950 595.050 341.400 ;
        RECT 43.950 339.600 46.050 340.050 ;
        RECT 61.950 339.600 64.050 340.050 ;
        RECT 43.950 338.400 64.050 339.600 ;
        RECT 43.950 337.950 46.050 338.400 ;
        RECT 61.950 337.950 64.050 338.400 ;
        RECT 130.950 339.600 133.050 340.050 ;
        RECT 145.950 339.600 148.050 340.050 ;
        RECT 130.950 338.400 148.050 339.600 ;
        RECT 130.950 337.950 133.050 338.400 ;
        RECT 145.950 337.950 148.050 338.400 ;
        RECT 157.950 339.600 160.050 340.050 ;
        RECT 163.950 339.600 166.050 340.050 ;
        RECT 157.950 338.400 166.050 339.600 ;
        RECT 157.950 337.950 160.050 338.400 ;
        RECT 163.950 337.950 166.050 338.400 ;
        RECT 235.950 339.600 238.050 340.050 ;
        RECT 241.950 339.600 244.050 340.050 ;
        RECT 235.950 338.400 244.050 339.600 ;
        RECT 235.950 337.950 238.050 338.400 ;
        RECT 241.950 337.950 244.050 338.400 ;
        RECT 280.950 337.950 286.050 340.050 ;
        RECT 304.950 339.600 307.050 340.050 ;
        RECT 328.950 339.600 331.050 340.050 ;
        RECT 304.950 338.400 331.050 339.600 ;
        RECT 304.950 337.950 307.050 338.400 ;
        RECT 328.950 337.950 331.050 338.400 ;
        RECT 340.950 337.950 346.050 340.050 ;
        RECT 349.950 339.600 352.050 340.050 ;
        RECT 430.950 339.600 433.050 340.050 ;
        RECT 349.950 338.400 433.050 339.600 ;
        RECT 349.950 337.950 352.050 338.400 ;
        RECT 430.950 337.950 433.050 338.400 ;
        RECT 511.950 339.600 514.050 340.050 ;
        RECT 532.950 339.600 535.050 340.050 ;
        RECT 511.950 338.400 535.050 339.600 ;
        RECT 511.950 337.950 514.050 338.400 ;
        RECT 532.950 337.950 535.050 338.400 ;
        RECT 661.950 339.600 664.050 340.050 ;
        RECT 670.950 339.600 673.050 340.050 ;
        RECT 715.950 339.600 718.050 340.050 ;
        RECT 661.950 338.400 673.050 339.600 ;
        RECT 707.400 339.000 718.050 339.600 ;
        RECT 661.950 337.950 664.050 338.400 ;
        RECT 670.950 337.950 673.050 338.400 ;
        RECT 706.950 338.400 718.050 339.000 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 85.950 336.600 88.050 337.050 ;
        RECT 91.950 336.600 94.050 337.050 ;
        RECT 85.950 335.400 94.050 336.600 ;
        RECT 85.950 334.950 88.050 335.400 ;
        RECT 91.950 334.950 94.050 335.400 ;
        RECT 112.950 334.950 118.050 337.050 ;
        RECT 151.950 336.600 154.050 337.050 ;
        RECT 172.950 336.600 175.050 337.050 ;
        RECT 151.950 335.400 175.050 336.600 ;
        RECT 151.950 334.950 154.050 335.400 ;
        RECT 172.950 334.950 175.050 335.400 ;
        RECT 244.950 336.600 247.050 337.050 ;
        RECT 256.950 336.600 259.050 337.050 ;
        RECT 244.950 335.400 259.050 336.600 ;
        RECT 244.950 334.950 247.050 335.400 ;
        RECT 256.950 334.950 259.050 335.400 ;
        RECT 7.950 330.600 10.050 334.050 ;
        RECT 41.400 331.050 42.600 334.950 ;
        RECT 64.950 333.600 67.050 334.050 ;
        RECT 79.950 333.600 82.050 334.050 ;
        RECT 136.950 333.600 139.050 334.050 ;
        RECT 166.950 333.600 169.050 334.050 ;
        RECT 64.950 332.400 139.050 333.600 ;
        RECT 158.400 333.000 169.050 333.600 ;
        RECT 64.950 331.950 67.050 332.400 ;
        RECT 79.950 331.950 82.050 332.400 ;
        RECT 136.950 331.950 139.050 332.400 ;
        RECT 157.950 332.400 169.050 333.000 ;
        RECT 25.950 330.600 28.050 331.050 ;
        RECT 7.950 330.000 28.050 330.600 ;
        RECT 8.400 329.400 28.050 330.000 ;
        RECT 25.950 328.950 28.050 329.400 ;
        RECT 40.950 328.950 43.050 331.050 ;
        RECT 145.950 330.600 148.050 331.050 ;
        RECT 151.950 330.600 154.050 331.050 ;
        RECT 145.950 329.400 154.050 330.600 ;
        RECT 145.950 328.950 148.050 329.400 ;
        RECT 151.950 328.950 154.050 329.400 ;
        RECT 157.950 328.950 160.050 332.400 ;
        RECT 166.950 331.950 169.050 332.400 ;
        RECT 271.950 333.600 277.050 334.050 ;
        RECT 334.950 333.600 337.050 337.050 ;
        RECT 367.950 336.600 370.050 337.050 ;
        RECT 376.950 336.600 379.050 337.050 ;
        RECT 367.950 335.400 379.050 336.600 ;
        RECT 367.950 334.950 370.050 335.400 ;
        RECT 376.950 334.950 379.050 335.400 ;
        RECT 457.950 336.600 460.050 337.050 ;
        RECT 463.950 336.600 466.050 337.050 ;
        RECT 478.950 336.600 481.050 337.050 ;
        RECT 490.950 336.600 493.050 337.050 ;
        RECT 457.950 335.400 493.050 336.600 ;
        RECT 457.950 334.950 460.050 335.400 ;
        RECT 463.950 334.950 466.050 335.400 ;
        RECT 478.950 334.950 481.050 335.400 ;
        RECT 490.950 334.950 493.050 335.400 ;
        RECT 580.950 336.600 583.050 337.050 ;
        RECT 613.950 336.600 616.050 337.050 ;
        RECT 580.950 335.400 616.050 336.600 ;
        RECT 580.950 334.950 583.050 335.400 ;
        RECT 613.950 334.950 616.050 335.400 ;
        RECT 667.950 336.600 670.050 337.050 ;
        RECT 667.950 336.000 690.600 336.600 ;
        RECT 667.950 335.400 691.050 336.000 ;
        RECT 667.950 334.950 670.050 335.400 ;
        RECT 271.950 333.000 337.050 333.600 ;
        RECT 271.950 332.400 336.600 333.000 ;
        RECT 271.950 331.950 277.050 332.400 ;
        RECT 520.950 331.950 526.050 334.050 ;
        RECT 619.950 333.600 622.050 333.900 ;
        RECT 628.950 333.600 631.050 334.050 ;
        RECT 619.950 332.400 631.050 333.600 ;
        RECT 619.950 331.800 622.050 332.400 ;
        RECT 628.950 331.950 631.050 332.400 ;
        RECT 640.950 333.600 643.050 334.050 ;
        RECT 661.950 333.600 664.050 334.050 ;
        RECT 640.950 332.400 664.050 333.600 ;
        RECT 640.950 331.950 643.050 332.400 ;
        RECT 661.950 331.950 664.050 332.400 ;
        RECT 688.950 331.950 691.050 335.400 ;
        RECT 706.950 334.950 709.050 338.400 ;
        RECT 715.950 337.950 718.050 338.400 ;
        RECT 739.950 336.600 742.050 337.050 ;
        RECT 760.950 336.600 763.050 337.050 ;
        RECT 739.950 335.400 763.050 336.600 ;
        RECT 739.950 334.950 742.050 335.400 ;
        RECT 760.950 334.950 763.050 335.400 ;
        RECT 769.950 336.600 772.050 337.050 ;
        RECT 778.950 336.600 781.050 337.050 ;
        RECT 769.950 335.400 781.050 336.600 ;
        RECT 769.950 334.950 772.050 335.400 ;
        RECT 778.950 334.950 781.050 335.400 ;
        RECT 787.950 336.600 790.050 337.050 ;
        RECT 805.950 336.600 808.050 337.050 ;
        RECT 787.950 335.400 808.050 336.600 ;
        RECT 787.950 334.950 790.050 335.400 ;
        RECT 805.950 334.950 808.050 335.400 ;
        RECT 730.950 331.950 736.050 334.050 ;
        RECT 808.950 333.600 811.050 334.050 ;
        RECT 820.950 333.600 823.050 334.050 ;
        RECT 808.950 332.400 823.050 333.600 ;
        RECT 808.950 331.950 811.050 332.400 ;
        RECT 820.950 331.950 823.050 332.400 ;
        RECT 196.950 330.600 199.050 331.050 ;
        RECT 304.950 330.600 307.050 331.050 ;
        RECT 343.950 330.600 346.050 331.050 ;
        RECT 358.950 330.600 361.050 331.050 ;
        RECT 196.950 329.400 361.050 330.600 ;
        RECT 196.950 328.950 199.050 329.400 ;
        RECT 304.950 328.950 307.050 329.400 ;
        RECT 343.950 328.950 346.050 329.400 ;
        RECT 358.950 328.950 361.050 329.400 ;
        RECT 388.950 330.600 391.050 331.050 ;
        RECT 427.950 330.600 430.050 331.050 ;
        RECT 388.950 329.400 430.050 330.600 ;
        RECT 388.950 328.950 391.050 329.400 ;
        RECT 427.950 328.950 430.050 329.400 ;
        RECT 442.950 330.600 445.050 331.050 ;
        RECT 469.950 330.600 472.050 331.050 ;
        RECT 505.950 330.600 508.050 331.050 ;
        RECT 442.950 329.400 508.050 330.600 ;
        RECT 442.950 328.950 445.050 329.400 ;
        RECT 469.950 328.950 472.050 329.400 ;
        RECT 505.950 328.950 508.050 329.400 ;
        RECT 532.950 330.600 535.050 331.050 ;
        RECT 544.950 330.600 547.050 331.050 ;
        RECT 586.950 330.600 589.050 331.050 ;
        RECT 532.950 329.400 589.050 330.600 ;
        RECT 620.400 330.600 621.600 331.800 ;
        RECT 634.950 330.600 637.050 331.050 ;
        RECT 620.400 329.400 637.050 330.600 ;
        RECT 532.950 328.950 535.050 329.400 ;
        RECT 544.950 328.950 547.050 329.400 ;
        RECT 586.950 328.950 589.050 329.400 ;
        RECT 634.950 328.950 637.050 329.400 ;
        RECT 49.950 327.600 52.050 328.050 ;
        RECT 58.950 327.600 61.050 328.050 ;
        RECT 73.950 327.600 76.050 328.050 ;
        RECT 49.950 326.400 76.050 327.600 ;
        RECT 49.950 325.950 52.050 326.400 ;
        RECT 58.950 325.950 61.050 326.400 ;
        RECT 73.950 325.950 76.050 326.400 ;
        RECT 133.950 327.600 136.050 328.050 ;
        RECT 190.950 327.600 193.050 328.050 ;
        RECT 133.950 326.400 193.050 327.600 ;
        RECT 133.950 325.950 136.050 326.400 ;
        RECT 190.950 325.950 193.050 326.400 ;
        RECT 220.950 327.600 223.050 328.050 ;
        RECT 250.950 327.600 253.050 328.050 ;
        RECT 220.950 326.400 253.050 327.600 ;
        RECT 220.950 325.950 223.050 326.400 ;
        RECT 250.950 325.950 253.050 326.400 ;
        RECT 547.950 327.600 550.050 328.050 ;
        RECT 646.950 327.600 649.050 328.050 ;
        RECT 547.950 326.400 649.050 327.600 ;
        RECT 547.950 325.950 550.050 326.400 ;
        RECT 646.950 325.950 649.050 326.400 ;
        RECT 712.950 327.600 715.050 328.050 ;
        RECT 742.950 327.600 745.050 328.050 ;
        RECT 712.950 326.400 745.050 327.600 ;
        RECT 712.950 325.950 715.050 326.400 ;
        RECT 742.950 325.950 745.050 326.400 ;
        RECT 13.950 324.600 16.050 325.050 ;
        RECT 37.950 324.600 40.050 325.050 ;
        RECT 13.950 323.400 40.050 324.600 ;
        RECT 13.950 322.950 16.050 323.400 ;
        RECT 37.950 322.950 40.050 323.400 ;
        RECT 373.950 324.600 376.050 325.050 ;
        RECT 448.950 324.600 451.050 325.050 ;
        RECT 373.950 323.400 451.050 324.600 ;
        RECT 373.950 322.950 376.050 323.400 ;
        RECT 448.950 322.950 451.050 323.400 ;
        RECT 583.950 324.600 586.050 325.050 ;
        RECT 613.950 324.600 616.050 325.050 ;
        RECT 583.950 323.400 616.050 324.600 ;
        RECT 583.950 322.950 586.050 323.400 ;
        RECT 613.950 322.950 616.050 323.400 ;
        RECT 88.950 321.600 91.050 322.050 ;
        RECT 160.950 321.600 163.050 322.050 ;
        RECT 88.950 320.400 163.050 321.600 ;
        RECT 88.950 319.950 91.050 320.400 ;
        RECT 160.950 319.950 163.050 320.400 ;
        RECT 202.950 321.600 205.050 322.050 ;
        RECT 253.950 321.600 256.050 322.050 ;
        RECT 202.950 320.400 256.050 321.600 ;
        RECT 202.950 319.950 205.050 320.400 ;
        RECT 253.950 319.950 256.050 320.400 ;
        RECT 457.950 321.600 460.050 322.050 ;
        RECT 484.950 321.600 487.050 322.050 ;
        RECT 697.950 321.600 700.050 322.050 ;
        RECT 457.950 320.400 700.050 321.600 ;
        RECT 457.950 319.950 460.050 320.400 ;
        RECT 484.950 319.950 487.050 320.400 ;
        RECT 697.950 319.950 700.050 320.400 ;
        RECT 394.950 318.600 397.050 319.050 ;
        RECT 403.950 318.600 406.050 319.050 ;
        RECT 394.950 317.400 406.050 318.600 ;
        RECT 394.950 316.950 397.050 317.400 ;
        RECT 403.950 316.950 406.050 317.400 ;
        RECT 430.950 318.600 433.050 319.050 ;
        RECT 436.950 318.600 439.050 319.050 ;
        RECT 430.950 317.400 439.050 318.600 ;
        RECT 430.950 316.950 433.050 317.400 ;
        RECT 436.950 316.950 439.050 317.400 ;
        RECT 715.950 318.600 718.050 319.050 ;
        RECT 757.950 318.600 760.050 319.050 ;
        RECT 715.950 317.400 760.050 318.600 ;
        RECT 715.950 316.950 718.050 317.400 ;
        RECT 757.950 316.950 760.050 317.400 ;
        RECT 193.950 315.600 196.050 316.050 ;
        RECT 220.950 315.600 223.050 316.050 ;
        RECT 229.950 315.600 232.050 316.050 ;
        RECT 193.950 314.400 232.050 315.600 ;
        RECT 193.950 313.950 196.050 314.400 ;
        RECT 220.950 313.950 223.050 314.400 ;
        RECT 229.950 313.950 232.050 314.400 ;
        RECT 427.950 315.600 430.050 316.050 ;
        RECT 472.950 315.600 475.050 316.050 ;
        RECT 427.950 314.400 475.050 315.600 ;
        RECT 427.950 313.950 430.050 314.400 ;
        RECT 472.950 313.950 475.050 314.400 ;
        RECT 352.950 312.600 355.050 313.050 ;
        RECT 388.950 312.600 391.050 313.050 ;
        RECT 352.950 311.400 391.050 312.600 ;
        RECT 352.950 310.950 355.050 311.400 ;
        RECT 388.950 310.950 391.050 311.400 ;
        RECT 439.950 312.600 442.050 313.050 ;
        RECT 460.950 312.600 463.050 313.050 ;
        RECT 541.950 312.600 544.050 313.050 ;
        RECT 439.950 311.400 544.050 312.600 ;
        RECT 439.950 310.950 442.050 311.400 ;
        RECT 460.950 310.950 463.050 311.400 ;
        RECT 541.950 310.950 544.050 311.400 ;
        RECT 670.950 312.600 673.050 313.050 ;
        RECT 706.950 312.600 709.050 313.050 ;
        RECT 718.950 312.600 721.050 313.050 ;
        RECT 670.950 311.400 721.050 312.600 ;
        RECT 670.950 310.950 673.050 311.400 ;
        RECT 706.950 310.950 709.050 311.400 ;
        RECT 718.950 310.950 721.050 311.400 ;
        RECT 796.950 312.600 799.050 313.050 ;
        RECT 802.950 312.600 805.050 313.050 ;
        RECT 796.950 311.400 805.050 312.600 ;
        RECT 796.950 310.950 799.050 311.400 ;
        RECT 802.950 310.950 805.050 311.400 ;
        RECT 4.950 309.600 7.050 310.050 ;
        RECT 13.950 309.600 16.050 310.050 ;
        RECT 4.950 308.400 16.050 309.600 ;
        RECT 4.950 307.950 7.050 308.400 ;
        RECT 13.950 307.950 16.050 308.400 ;
        RECT 34.950 309.600 37.050 310.050 ;
        RECT 100.950 309.600 103.050 310.050 ;
        RECT 34.950 308.400 103.050 309.600 ;
        RECT 34.950 307.950 37.050 308.400 ;
        RECT 100.950 307.950 103.050 308.400 ;
        RECT 217.950 309.600 220.050 310.050 ;
        RECT 226.950 309.600 229.050 310.050 ;
        RECT 217.950 308.400 229.050 309.600 ;
        RECT 217.950 307.950 220.050 308.400 ;
        RECT 226.950 307.950 229.050 308.400 ;
        RECT 241.950 309.600 244.050 310.050 ;
        RECT 283.950 309.600 286.050 310.050 ;
        RECT 241.950 308.400 286.050 309.600 ;
        RECT 241.950 307.950 244.050 308.400 ;
        RECT 283.950 307.950 286.050 308.400 ;
        RECT 367.950 309.600 370.050 310.050 ;
        RECT 397.950 309.600 400.050 310.050 ;
        RECT 367.950 308.400 400.050 309.600 ;
        RECT 367.950 307.950 370.050 308.400 ;
        RECT 397.950 307.950 400.050 308.400 ;
        RECT 550.950 309.600 553.050 310.050 ;
        RECT 598.950 309.600 601.050 310.050 ;
        RECT 550.950 308.400 601.050 309.600 ;
        RECT 550.950 307.950 553.050 308.400 ;
        RECT 598.950 307.950 601.050 308.400 ;
        RECT 46.950 306.600 49.050 307.050 ;
        RECT 97.950 306.600 100.050 307.050 ;
        RECT 46.950 305.400 100.050 306.600 ;
        RECT 46.950 304.950 49.050 305.400 ;
        RECT 97.950 304.950 100.050 305.400 ;
        RECT 655.950 306.600 658.050 307.050 ;
        RECT 715.950 306.600 718.050 307.050 ;
        RECT 655.950 305.400 718.050 306.600 ;
        RECT 655.950 304.950 658.050 305.400 ;
        RECT 715.950 304.950 718.050 305.400 ;
        RECT 376.950 303.600 379.050 304.050 ;
        RECT 424.950 303.600 427.050 304.050 ;
        RECT 376.950 302.400 427.050 303.600 ;
        RECT 376.950 301.950 379.050 302.400 ;
        RECT 424.950 301.950 427.050 302.400 ;
        RECT 451.950 303.600 454.050 304.050 ;
        RECT 469.950 303.600 472.050 304.050 ;
        RECT 451.950 302.400 472.050 303.600 ;
        RECT 451.950 301.950 454.050 302.400 ;
        RECT 469.950 301.950 472.050 302.400 ;
        RECT 592.950 303.600 595.050 304.050 ;
        RECT 622.950 303.600 625.050 304.050 ;
        RECT 592.950 302.400 625.050 303.600 ;
        RECT 592.950 301.950 595.050 302.400 ;
        RECT 622.950 301.950 625.050 302.400 ;
        RECT 637.950 303.600 640.050 304.050 ;
        RECT 745.950 303.600 748.050 304.050 ;
        RECT 637.950 302.400 748.050 303.600 ;
        RECT 637.950 301.950 640.050 302.400 ;
        RECT 745.950 301.950 748.050 302.400 ;
        RECT 763.950 303.600 766.050 304.050 ;
        RECT 799.950 303.600 802.050 304.050 ;
        RECT 763.950 302.400 802.050 303.600 ;
        RECT 763.950 301.950 766.050 302.400 ;
        RECT 799.950 301.950 802.050 302.400 ;
        RECT 4.950 300.600 7.050 301.050 ;
        RECT 13.950 300.600 16.050 301.050 ;
        RECT 4.950 299.400 16.050 300.600 ;
        RECT 4.950 298.950 7.050 299.400 ;
        RECT 13.950 298.950 16.050 299.400 ;
        RECT 40.950 300.600 43.050 301.200 ;
        RECT 52.950 300.600 55.050 301.050 ;
        RECT 40.950 299.400 55.050 300.600 ;
        RECT 40.950 299.100 43.050 299.400 ;
        RECT 52.950 298.950 55.050 299.400 ;
        RECT 280.950 300.600 283.050 301.050 ;
        RECT 289.950 300.600 292.050 301.050 ;
        RECT 280.950 299.400 292.050 300.600 ;
        RECT 280.950 298.950 283.050 299.400 ;
        RECT 289.950 298.950 292.050 299.400 ;
        RECT 223.950 296.100 226.050 298.200 ;
        RECT 298.950 297.600 301.050 298.050 ;
        RECT 340.950 297.600 343.050 298.050 ;
        RECT 298.950 296.400 343.050 297.600 ;
        RECT 136.950 295.050 139.050 295.200 ;
        RECT 43.950 294.600 46.050 295.050 ;
        RECT 52.950 294.600 55.050 295.050 ;
        RECT 43.950 293.400 55.050 294.600 ;
        RECT 43.950 292.950 46.050 293.400 ;
        RECT 52.950 292.950 55.050 293.400 ;
        RECT 73.950 291.600 76.050 295.050 ;
        RECT 94.950 294.600 97.050 295.050 ;
        RECT 121.950 294.600 124.050 295.050 ;
        RECT 94.950 293.400 124.050 294.600 ;
        RECT 94.950 292.950 97.050 293.400 ;
        RECT 121.950 292.950 124.050 293.400 ;
        RECT 136.950 293.100 142.050 295.050 ;
        RECT 138.000 292.950 142.050 293.100 ;
        RECT 100.950 291.600 103.050 292.050 ;
        RECT 73.950 291.000 103.050 291.600 ;
        RECT 74.400 290.400 103.050 291.000 ;
        RECT 100.950 289.950 103.050 290.400 ;
        RECT 49.950 286.950 55.050 289.050 ;
        RECT 136.950 288.600 139.050 291.900 ;
        RECT 142.950 288.600 145.050 292.050 ;
        RECT 151.950 291.600 154.050 292.050 ;
        RECT 193.950 291.600 196.050 292.050 ;
        RECT 224.400 291.900 225.600 296.100 ;
        RECT 298.950 295.950 301.050 296.400 ;
        RECT 340.950 295.950 343.050 296.400 ;
        RECT 415.950 297.600 418.050 298.050 ;
        RECT 427.950 297.600 430.050 301.050 ;
        RECT 553.950 300.600 556.050 301.050 ;
        RECT 649.950 300.600 652.050 301.050 ;
        RECT 553.950 299.400 652.050 300.600 ;
        RECT 553.950 298.950 556.050 299.400 ;
        RECT 649.950 298.950 652.050 299.400 ;
        RECT 676.950 300.600 679.050 301.050 ;
        RECT 688.950 300.600 691.050 301.050 ;
        RECT 676.950 299.400 691.050 300.600 ;
        RECT 676.950 298.950 679.050 299.400 ;
        RECT 688.950 298.950 691.050 299.400 ;
        RECT 727.950 300.600 730.050 301.050 ;
        RECT 739.950 300.600 742.050 301.050 ;
        RECT 727.950 299.400 742.050 300.600 ;
        RECT 727.950 298.950 730.050 299.400 ;
        RECT 739.950 298.950 742.050 299.400 ;
        RECT 805.950 300.600 808.050 301.050 ;
        RECT 817.950 300.600 820.050 301.050 ;
        RECT 805.950 299.400 820.050 300.600 ;
        RECT 805.950 298.950 808.050 299.400 ;
        RECT 817.950 298.950 820.050 299.400 ;
        RECT 415.950 297.000 430.050 297.600 ;
        RECT 505.950 297.600 508.050 298.050 ;
        RECT 523.950 297.600 526.050 298.050 ;
        RECT 415.950 296.400 429.600 297.000 ;
        RECT 505.950 296.400 526.050 297.600 ;
        RECT 415.950 295.950 418.050 296.400 ;
        RECT 505.950 295.950 508.050 296.400 ;
        RECT 523.950 295.950 526.050 296.400 ;
        RECT 571.950 297.600 574.050 298.050 ;
        RECT 586.950 297.600 589.050 298.050 ;
        RECT 571.950 296.400 589.050 297.600 ;
        RECT 571.950 295.950 574.050 296.400 ;
        RECT 586.950 295.950 589.050 296.400 ;
        RECT 604.950 297.600 607.050 298.050 ;
        RECT 637.950 297.600 640.050 298.050 ;
        RECT 604.950 296.400 640.050 297.600 ;
        RECT 604.950 295.950 607.050 296.400 ;
        RECT 637.950 295.950 640.050 296.400 ;
        RECT 646.950 297.600 649.050 298.050 ;
        RECT 652.950 297.600 655.050 298.050 ;
        RECT 646.950 296.400 655.050 297.600 ;
        RECT 646.950 295.950 649.050 296.400 ;
        RECT 652.950 295.950 655.050 296.400 ;
        RECT 712.950 297.600 715.050 298.050 ;
        RECT 724.950 297.600 727.050 298.050 ;
        RECT 748.950 297.600 751.050 298.050 ;
        RECT 775.950 297.600 778.050 298.050 ;
        RECT 712.950 296.400 778.050 297.600 ;
        RECT 712.950 295.950 715.050 296.400 ;
        RECT 724.950 295.950 727.050 296.400 ;
        RECT 748.950 295.950 751.050 296.400 ;
        RECT 775.950 295.950 778.050 296.400 ;
        RECT 799.950 297.600 802.050 298.050 ;
        RECT 808.950 297.600 811.050 298.050 ;
        RECT 799.950 296.400 811.050 297.600 ;
        RECT 799.950 295.950 802.050 296.400 ;
        RECT 808.950 295.950 811.050 296.400 ;
        RECT 256.950 292.950 262.050 295.050 ;
        RECT 274.950 294.600 277.050 295.050 ;
        RECT 316.950 294.600 319.050 295.050 ;
        RECT 367.950 294.600 370.050 295.050 ;
        RECT 274.950 293.400 370.050 294.600 ;
        RECT 274.950 292.950 277.050 293.400 ;
        RECT 316.950 292.950 319.050 293.400 ;
        RECT 367.950 292.950 370.050 293.400 ;
        RECT 400.950 294.600 403.050 295.050 ;
        RECT 409.950 294.600 412.050 295.050 ;
        RECT 400.950 293.400 412.050 294.600 ;
        RECT 400.950 292.950 403.050 293.400 ;
        RECT 409.950 292.950 412.050 293.400 ;
        RECT 418.950 294.600 421.050 295.050 ;
        RECT 442.950 294.600 445.050 295.050 ;
        RECT 537.000 294.600 541.050 295.050 ;
        RECT 418.950 293.400 445.050 294.600 ;
        RECT 418.950 292.950 421.050 293.400 ;
        RECT 442.950 292.950 445.050 293.400 ;
        RECT 536.400 292.950 541.050 294.600 ;
        RECT 610.950 294.600 616.050 295.050 ;
        RECT 619.950 294.600 622.050 295.050 ;
        RECT 610.950 293.400 622.050 294.600 ;
        RECT 610.950 292.950 616.050 293.400 ;
        RECT 619.950 292.950 622.050 293.400 ;
        RECT 796.950 294.600 799.050 295.050 ;
        RECT 811.950 294.600 814.050 295.050 ;
        RECT 796.950 293.400 814.050 294.600 ;
        RECT 796.950 292.950 799.050 293.400 ;
        RECT 811.950 292.950 814.050 293.400 ;
        RECT 151.950 290.400 196.050 291.600 ;
        RECT 151.950 289.950 154.050 290.400 ;
        RECT 193.950 289.950 196.050 290.400 ;
        RECT 223.950 289.800 226.050 291.900 ;
        RECT 451.950 291.600 454.050 291.900 ;
        RECT 478.950 291.600 481.050 292.050 ;
        RECT 451.950 290.400 481.050 291.600 ;
        RECT 451.950 289.800 454.050 290.400 ;
        RECT 478.950 289.950 481.050 290.400 ;
        RECT 526.950 291.600 529.050 292.050 ;
        RECT 536.400 291.600 537.600 292.950 ;
        RECT 526.950 290.400 537.600 291.600 ;
        RECT 541.950 291.600 544.050 292.050 ;
        RECT 574.950 291.600 577.050 292.050 ;
        RECT 541.950 290.400 577.050 291.600 ;
        RECT 526.950 289.950 529.050 290.400 ;
        RECT 541.950 289.950 544.050 290.400 ;
        RECT 574.950 289.950 577.050 290.400 ;
        RECT 652.950 291.600 655.050 292.050 ;
        RECT 679.950 291.600 682.050 292.050 ;
        RECT 691.950 291.600 694.050 292.050 ;
        RECT 652.950 290.400 694.050 291.600 ;
        RECT 652.950 289.950 655.050 290.400 ;
        RECT 679.950 289.950 682.050 290.400 ;
        RECT 691.950 289.950 694.050 290.400 ;
        RECT 751.950 291.600 754.050 292.050 ;
        RECT 772.950 291.900 777.000 292.050 ;
        RECT 772.950 291.600 778.050 291.900 ;
        RECT 751.950 290.400 778.050 291.600 ;
        RECT 751.950 289.950 754.050 290.400 ;
        RECT 772.950 289.950 778.050 290.400 ;
        RECT 775.950 289.800 778.050 289.950 ;
        RECT 136.950 288.000 145.050 288.600 ;
        RECT 253.950 288.600 256.050 289.050 ;
        RECT 295.950 288.600 298.050 289.050 ;
        RECT 137.400 287.400 144.600 288.000 ;
        RECT 253.950 287.400 298.050 288.600 ;
        RECT 253.950 286.950 256.050 287.400 ;
        RECT 295.950 286.950 298.050 287.400 ;
        RECT 313.950 288.600 316.050 289.050 ;
        RECT 319.950 288.600 322.050 289.050 ;
        RECT 325.950 288.600 328.050 289.050 ;
        RECT 313.950 287.400 328.050 288.600 ;
        RECT 313.950 286.950 316.050 287.400 ;
        RECT 319.950 286.950 322.050 287.400 ;
        RECT 325.950 286.950 328.050 287.400 ;
        RECT 346.950 288.600 349.050 289.050 ;
        RECT 376.950 288.600 379.050 289.050 ;
        RECT 346.950 287.400 379.050 288.600 ;
        RECT 346.950 286.950 349.050 287.400 ;
        RECT 376.950 286.950 379.050 287.400 ;
        RECT 424.950 288.600 427.050 289.050 ;
        RECT 430.950 288.600 433.050 289.050 ;
        RECT 424.950 287.400 433.050 288.600 ;
        RECT 424.950 286.950 427.050 287.400 ;
        RECT 430.950 286.950 433.050 287.400 ;
        RECT 517.950 288.600 520.050 289.050 ;
        RECT 529.950 288.600 532.050 289.050 ;
        RECT 517.950 287.400 532.050 288.600 ;
        RECT 517.950 286.950 520.050 287.400 ;
        RECT 529.950 286.950 532.050 287.400 ;
        RECT 613.950 288.600 616.050 289.050 ;
        RECT 631.950 288.600 634.050 289.050 ;
        RECT 613.950 287.400 634.050 288.600 ;
        RECT 613.950 286.950 616.050 287.400 ;
        RECT 631.950 286.950 634.050 287.400 ;
        RECT 661.950 288.600 664.050 289.050 ;
        RECT 673.950 288.600 676.050 289.050 ;
        RECT 661.950 287.400 676.050 288.600 ;
        RECT 661.950 286.950 664.050 287.400 ;
        RECT 673.950 286.950 676.050 287.400 ;
        RECT 715.950 288.600 718.050 289.200 ;
        RECT 784.950 288.600 787.050 289.050 ;
        RECT 807.000 288.900 811.050 289.050 ;
        RECT 715.950 287.400 787.050 288.600 ;
        RECT 715.950 287.100 718.050 287.400 ;
        RECT 784.950 286.950 787.050 287.400 ;
        RECT 805.950 286.950 811.050 288.900 ;
        RECT 805.950 286.800 808.050 286.950 ;
        RECT 4.950 285.600 7.050 286.050 ;
        RECT 13.950 285.600 16.050 286.050 ;
        RECT 4.950 284.400 16.050 285.600 ;
        RECT 4.950 283.950 7.050 284.400 ;
        RECT 13.950 283.950 16.050 284.400 ;
        RECT 433.950 285.600 436.050 286.050 ;
        RECT 451.950 285.600 454.050 285.900 ;
        RECT 460.950 285.600 463.050 286.050 ;
        RECT 433.950 284.400 463.050 285.600 ;
        RECT 433.950 283.950 436.050 284.400 ;
        RECT 451.950 283.800 454.050 284.400 ;
        RECT 460.950 283.950 463.050 284.400 ;
        RECT 565.950 285.600 568.050 286.050 ;
        RECT 580.950 285.600 583.050 286.050 ;
        RECT 565.950 284.400 583.050 285.600 ;
        RECT 565.950 283.950 568.050 284.400 ;
        RECT 580.950 283.950 583.050 284.400 ;
        RECT 664.950 285.600 667.050 286.050 ;
        RECT 685.950 285.600 688.050 286.050 ;
        RECT 664.950 284.400 688.050 285.600 ;
        RECT 664.950 283.950 667.050 284.400 ;
        RECT 685.950 283.950 688.050 284.400 ;
        RECT 742.950 285.600 745.050 286.050 ;
        RECT 751.950 285.600 754.050 286.050 ;
        RECT 742.950 284.400 754.050 285.600 ;
        RECT 742.950 283.950 745.050 284.400 ;
        RECT 751.950 283.950 754.050 284.400 ;
        RECT 19.950 282.600 22.050 283.050 ;
        RECT 67.950 282.600 70.050 283.050 ;
        RECT 19.950 281.400 70.050 282.600 ;
        RECT 19.950 280.950 22.050 281.400 ;
        RECT 67.950 280.950 70.050 281.400 ;
        RECT 208.950 282.600 211.050 283.050 ;
        RECT 250.950 282.600 253.050 283.050 ;
        RECT 208.950 281.400 253.050 282.600 ;
        RECT 208.950 280.950 211.050 281.400 ;
        RECT 250.950 280.950 253.050 281.400 ;
        RECT 418.950 282.600 421.050 283.050 ;
        RECT 424.950 282.600 427.050 283.050 ;
        RECT 418.950 281.400 427.050 282.600 ;
        RECT 418.950 280.950 421.050 281.400 ;
        RECT 424.950 280.950 427.050 281.400 ;
        RECT 478.950 282.600 481.050 283.050 ;
        RECT 490.950 282.600 493.050 283.050 ;
        RECT 517.950 282.600 520.050 283.050 ;
        RECT 478.950 281.400 520.050 282.600 ;
        RECT 478.950 280.950 481.050 281.400 ;
        RECT 490.950 280.950 493.050 281.400 ;
        RECT 517.950 280.950 520.050 281.400 ;
        RECT 697.950 282.600 700.050 283.050 ;
        RECT 805.950 282.600 808.050 283.050 ;
        RECT 697.950 281.400 808.050 282.600 ;
        RECT 697.950 280.950 700.050 281.400 ;
        RECT 805.950 280.950 808.050 281.400 ;
        RECT 457.950 279.600 460.050 280.050 ;
        RECT 469.800 279.600 471.900 280.050 ;
        RECT 457.950 278.400 471.900 279.600 ;
        RECT 457.950 277.950 460.050 278.400 ;
        RECT 469.800 277.950 471.900 278.400 ;
        RECT 473.100 279.600 475.200 280.050 ;
        RECT 532.950 279.600 535.050 280.050 ;
        RECT 473.100 278.400 535.050 279.600 ;
        RECT 473.100 277.950 475.200 278.400 ;
        RECT 532.950 277.950 535.050 278.400 ;
        RECT 634.950 279.600 637.050 280.050 ;
        RECT 667.950 279.600 670.050 280.050 ;
        RECT 634.950 278.400 670.050 279.600 ;
        RECT 634.950 277.950 637.050 278.400 ;
        RECT 667.950 277.950 670.050 278.400 ;
        RECT 700.950 279.600 703.050 280.050 ;
        RECT 760.950 279.600 763.050 280.050 ;
        RECT 700.950 278.400 763.050 279.600 ;
        RECT 700.950 277.950 703.050 278.400 ;
        RECT 760.950 277.950 763.050 278.400 ;
        RECT 82.950 276.600 85.050 277.050 ;
        RECT 94.950 276.600 97.050 277.050 ;
        RECT 82.950 275.400 97.050 276.600 ;
        RECT 82.950 274.950 85.050 275.400 ;
        RECT 94.950 274.950 97.050 275.400 ;
        RECT 265.950 276.600 268.050 277.050 ;
        RECT 298.950 276.600 301.050 277.050 ;
        RECT 328.950 276.600 331.050 277.050 ;
        RECT 265.950 275.400 331.050 276.600 ;
        RECT 265.950 274.950 268.050 275.400 ;
        RECT 298.950 274.950 301.050 275.400 ;
        RECT 328.950 274.950 331.050 275.400 ;
        RECT 355.950 276.600 358.050 277.050 ;
        RECT 370.950 276.600 373.050 277.050 ;
        RECT 415.950 276.600 418.050 277.050 ;
        RECT 496.950 276.600 499.050 277.050 ;
        RECT 355.950 275.400 499.050 276.600 ;
        RECT 355.950 274.950 358.050 275.400 ;
        RECT 370.950 274.950 373.050 275.400 ;
        RECT 415.950 274.950 418.050 275.400 ;
        RECT 496.950 274.950 499.050 275.400 ;
        RECT 802.950 276.600 805.050 277.050 ;
        RECT 811.950 276.600 814.050 277.050 ;
        RECT 802.950 275.400 814.050 276.600 ;
        RECT 802.950 274.950 805.050 275.400 ;
        RECT 811.950 274.950 814.050 275.400 ;
        RECT 13.950 273.600 16.050 274.050 ;
        RECT 8.400 272.400 16.050 273.600 ;
        RECT 8.400 270.600 9.600 272.400 ;
        RECT 13.950 271.950 16.050 272.400 ;
        RECT 22.950 273.600 25.050 274.050 ;
        RECT 37.950 273.600 40.050 274.050 ;
        RECT 55.950 273.600 58.050 274.050 ;
        RECT 97.950 273.600 100.050 274.050 ;
        RECT 22.950 272.400 100.050 273.600 ;
        RECT 22.950 271.950 25.050 272.400 ;
        RECT 37.950 271.950 40.050 272.400 ;
        RECT 55.950 271.950 58.050 272.400 ;
        RECT 97.950 271.950 100.050 272.400 ;
        RECT 5.400 269.400 9.600 270.600 ;
        RECT 100.950 270.600 103.050 271.050 ;
        RECT 106.950 270.600 109.050 271.050 ;
        RECT 100.950 269.400 109.050 270.600 ;
        RECT 5.400 265.050 6.600 269.400 ;
        RECT 100.950 268.950 103.050 269.400 ;
        RECT 106.950 268.950 109.050 269.400 ;
        RECT 229.950 270.600 232.050 271.050 ;
        RECT 256.950 270.600 259.050 271.050 ;
        RECT 229.950 269.400 259.050 270.600 ;
        RECT 229.950 268.950 232.050 269.400 ;
        RECT 256.950 268.950 259.050 269.400 ;
        RECT 367.950 270.600 370.050 271.050 ;
        RECT 385.950 270.600 388.050 274.050 ;
        RECT 595.950 273.600 598.050 274.050 ;
        RECT 676.950 273.600 679.050 274.050 ;
        RECT 700.950 273.600 703.050 274.050 ;
        RECT 798.000 273.600 802.050 274.050 ;
        RECT 595.950 272.400 669.600 273.600 ;
        RECT 595.950 271.950 598.050 272.400 ;
        RECT 367.950 270.000 388.050 270.600 ;
        RECT 427.950 270.600 430.050 271.050 ;
        RECT 454.950 270.600 457.050 271.050 ;
        RECT 367.950 269.400 387.600 270.000 ;
        RECT 427.950 269.400 457.050 270.600 ;
        RECT 367.950 268.950 370.050 269.400 ;
        RECT 427.950 268.950 430.050 269.400 ;
        RECT 454.950 268.950 457.050 269.400 ;
        RECT 574.950 270.600 577.050 271.050 ;
        RECT 640.950 270.600 643.050 271.050 ;
        RECT 574.950 269.400 643.050 270.600 ;
        RECT 668.400 270.600 669.600 272.400 ;
        RECT 676.950 272.400 703.050 273.600 ;
        RECT 676.950 271.950 679.050 272.400 ;
        RECT 700.950 271.950 703.050 272.400 ;
        RECT 797.400 271.950 802.050 273.600 ;
        RECT 724.950 270.600 727.050 271.050 ;
        RECT 668.400 269.400 727.050 270.600 ;
        RECT 574.950 268.950 577.050 269.400 ;
        RECT 640.950 268.950 643.050 269.400 ;
        RECT 724.950 268.950 727.050 269.400 ;
        RECT 781.950 270.600 784.050 271.050 ;
        RECT 790.950 270.600 793.050 271.050 ;
        RECT 781.950 269.400 793.050 270.600 ;
        RECT 781.950 268.950 784.050 269.400 ;
        RECT 790.950 268.950 793.050 269.400 ;
        RECT 13.950 267.600 16.050 268.050 ;
        RECT 46.950 267.600 49.050 268.050 ;
        RECT 13.950 266.400 49.050 267.600 ;
        RECT 13.950 265.950 16.050 266.400 ;
        RECT 46.950 265.950 49.050 266.400 ;
        RECT 121.950 267.600 124.050 268.050 ;
        RECT 178.950 267.600 181.050 268.050 ;
        RECT 121.950 266.400 181.050 267.600 ;
        RECT 121.950 265.950 124.050 266.400 ;
        RECT 178.950 265.950 181.050 266.400 ;
        RECT 232.950 267.600 235.050 268.050 ;
        RECT 280.950 267.600 283.050 268.050 ;
        RECT 232.950 266.400 283.050 267.600 ;
        RECT 232.950 265.950 235.050 266.400 ;
        RECT 280.950 265.950 283.050 266.400 ;
        RECT 499.950 267.600 502.050 268.050 ;
        RECT 553.950 267.600 556.050 268.050 ;
        RECT 499.950 266.400 556.050 267.600 ;
        RECT 499.950 265.950 502.050 266.400 ;
        RECT 553.950 265.950 556.050 266.400 ;
        RECT 577.950 267.600 580.050 268.050 ;
        RECT 601.950 267.600 604.050 268.050 ;
        RECT 622.950 267.600 625.050 268.050 ;
        RECT 577.950 266.400 625.050 267.600 ;
        RECT 577.950 265.950 580.050 266.400 ;
        RECT 601.950 265.950 604.050 266.400 ;
        RECT 622.950 265.950 625.050 266.400 ;
        RECT 757.950 267.600 760.050 268.050 ;
        RECT 763.950 267.600 766.050 268.050 ;
        RECT 757.950 266.400 766.050 267.600 ;
        RECT 757.950 265.950 760.050 266.400 ;
        RECT 763.950 265.950 766.050 266.400 ;
        RECT 797.400 265.050 798.600 271.950 ;
        RECT 4.950 262.950 7.050 265.050 ;
        RECT 67.950 264.600 70.050 265.050 ;
        RECT 109.950 264.600 112.050 265.050 ;
        RECT 67.950 263.400 112.050 264.600 ;
        RECT 67.950 262.950 70.050 263.400 ;
        RECT 109.950 262.950 112.050 263.400 ;
        RECT 34.950 261.600 37.050 262.050 ;
        RECT 40.950 261.600 43.050 262.050 ;
        RECT 61.950 261.600 64.050 262.050 ;
        RECT 34.950 260.400 64.050 261.600 ;
        RECT 118.950 261.600 121.050 265.050 ;
        RECT 151.950 264.600 154.050 265.050 ;
        RECT 184.950 264.600 187.050 265.050 ;
        RECT 151.950 263.400 187.050 264.600 ;
        RECT 151.950 262.950 154.050 263.400 ;
        RECT 184.950 262.950 187.050 263.400 ;
        RECT 235.950 264.600 238.050 265.050 ;
        RECT 268.950 264.600 271.050 265.050 ;
        RECT 235.950 263.400 271.050 264.600 ;
        RECT 235.950 262.950 238.050 263.400 ;
        RECT 268.950 262.950 271.050 263.400 ;
        RECT 127.950 261.600 130.050 262.050 ;
        RECT 118.950 261.000 130.050 261.600 ;
        RECT 119.400 260.400 130.050 261.000 ;
        RECT 34.950 259.950 37.050 260.400 ;
        RECT 40.950 259.950 43.050 260.400 ;
        RECT 61.950 259.950 64.050 260.400 ;
        RECT 127.950 259.950 130.050 260.400 ;
        RECT 292.950 261.600 295.050 262.050 ;
        RECT 310.950 261.600 313.050 265.050 ;
        RECT 340.950 264.600 343.050 265.050 ;
        RECT 370.950 264.600 373.050 265.050 ;
        RECT 340.950 263.400 373.050 264.600 ;
        RECT 340.950 262.950 343.050 263.400 ;
        RECT 370.950 262.950 373.050 263.400 ;
        RECT 406.950 264.600 409.050 265.050 ;
        RECT 436.950 264.600 439.050 265.050 ;
        RECT 442.950 264.600 445.050 265.050 ;
        RECT 469.950 264.600 472.050 265.050 ;
        RECT 406.950 263.400 472.050 264.600 ;
        RECT 406.950 262.950 409.050 263.400 ;
        RECT 436.950 262.950 439.050 263.400 ;
        RECT 442.950 262.950 445.050 263.400 ;
        RECT 469.950 262.950 472.050 263.400 ;
        RECT 292.950 261.000 313.050 261.600 ;
        RECT 505.950 261.600 508.050 262.050 ;
        RECT 520.950 261.600 523.050 265.050 ;
        RECT 565.950 264.600 568.050 265.050 ;
        RECT 574.950 264.600 577.050 265.050 ;
        RECT 565.950 263.400 577.050 264.600 ;
        RECT 565.950 262.950 568.050 263.400 ;
        RECT 574.950 262.950 577.050 263.400 ;
        RECT 715.950 264.600 718.050 265.050 ;
        RECT 739.950 264.600 742.050 265.050 ;
        RECT 754.950 264.600 757.050 265.050 ;
        RECT 715.950 263.400 738.600 264.600 ;
        RECT 715.950 262.950 718.050 263.400 ;
        RECT 505.950 261.000 523.050 261.600 ;
        RECT 589.950 261.600 592.050 262.050 ;
        RECT 607.950 261.600 610.050 262.050 ;
        RECT 292.950 260.400 312.600 261.000 ;
        RECT 505.950 260.400 522.600 261.000 ;
        RECT 589.950 260.400 610.050 261.600 ;
        RECT 292.950 259.950 295.050 260.400 ;
        RECT 505.950 259.950 508.050 260.400 ;
        RECT 589.950 259.950 592.050 260.400 ;
        RECT 607.950 259.950 610.050 260.400 ;
        RECT 637.950 261.600 640.050 262.050 ;
        RECT 658.950 261.600 661.050 262.050 ;
        RECT 637.950 260.400 661.050 261.600 ;
        RECT 737.400 261.600 738.600 263.400 ;
        RECT 739.950 263.400 757.050 264.600 ;
        RECT 739.950 262.950 742.050 263.400 ;
        RECT 754.950 262.950 757.050 263.400 ;
        RECT 796.950 262.950 799.050 265.050 ;
        RECT 763.950 261.600 766.050 262.050 ;
        RECT 737.400 260.400 766.050 261.600 ;
        RECT 637.950 259.950 640.050 260.400 ;
        RECT 658.950 259.950 661.050 260.400 ;
        RECT 763.950 259.950 766.050 260.400 ;
        RECT 109.950 258.600 112.050 259.050 ;
        RECT 154.950 258.600 157.050 259.050 ;
        RECT 109.950 257.400 157.050 258.600 ;
        RECT 109.950 256.950 112.050 257.400 ;
        RECT 154.950 256.950 157.050 257.400 ;
        RECT 169.950 258.600 172.050 259.050 ;
        RECT 205.950 258.600 208.050 259.050 ;
        RECT 169.950 257.400 208.050 258.600 ;
        RECT 169.950 256.950 172.050 257.400 ;
        RECT 205.950 256.950 208.050 257.400 ;
        RECT 223.950 256.950 229.050 259.050 ;
        RECT 244.950 258.600 247.050 259.050 ;
        RECT 250.950 258.600 253.050 259.050 ;
        RECT 244.950 257.400 253.050 258.600 ;
        RECT 244.950 256.950 247.050 257.400 ;
        RECT 250.950 256.950 253.050 257.400 ;
        RECT 271.950 258.600 274.050 259.050 ;
        RECT 280.950 258.600 283.050 259.050 ;
        RECT 271.950 257.400 283.050 258.600 ;
        RECT 271.950 256.950 274.050 257.400 ;
        RECT 280.950 256.950 283.050 257.400 ;
        RECT 322.950 258.600 325.050 259.200 ;
        RECT 328.950 258.600 331.050 258.900 ;
        RECT 322.950 257.400 331.050 258.600 ;
        RECT 322.950 257.100 325.050 257.400 ;
        RECT 328.950 256.800 331.050 257.400 ;
        RECT 376.950 258.600 379.050 259.050 ;
        RECT 415.950 258.600 418.050 259.050 ;
        RECT 376.950 257.400 418.050 258.600 ;
        RECT 376.950 256.950 379.050 257.400 ;
        RECT 415.950 256.950 418.050 257.400 ;
        RECT 463.950 258.600 466.050 259.200 ;
        RECT 469.950 258.600 472.050 259.050 ;
        RECT 463.950 257.400 472.050 258.600 ;
        RECT 463.950 257.100 466.050 257.400 ;
        RECT 469.950 256.950 472.050 257.400 ;
        RECT 499.950 258.600 502.050 258.900 ;
        RECT 514.950 258.600 517.050 259.050 ;
        RECT 499.950 257.400 517.050 258.600 ;
        RECT 499.950 256.800 502.050 257.400 ;
        RECT 514.950 256.950 517.050 257.400 ;
        RECT 37.950 255.600 40.050 256.200 ;
        RECT 43.950 255.600 46.050 256.050 ;
        RECT 37.950 254.400 46.050 255.600 ;
        RECT 37.950 254.100 40.050 254.400 ;
        RECT 43.950 253.950 46.050 254.400 ;
        RECT 55.950 255.600 58.050 256.050 ;
        RECT 67.950 255.600 70.050 256.050 ;
        RECT 55.950 254.400 70.050 255.600 ;
        RECT 55.950 253.950 58.050 254.400 ;
        RECT 67.950 253.950 70.050 254.400 ;
        RECT 124.950 255.600 127.050 256.050 ;
        RECT 130.950 255.600 133.050 256.050 ;
        RECT 124.950 254.400 133.050 255.600 ;
        RECT 124.950 253.950 127.050 254.400 ;
        RECT 130.950 253.950 133.050 254.400 ;
        RECT 184.950 255.600 187.050 256.050 ;
        RECT 202.950 255.600 205.050 256.050 ;
        RECT 324.000 255.900 328.050 256.050 ;
        RECT 184.950 254.400 205.050 255.600 ;
        RECT 184.950 253.950 187.050 254.400 ;
        RECT 202.950 253.950 205.050 254.400 ;
        RECT 322.950 253.950 328.050 255.900 ;
        RECT 322.950 253.800 325.050 253.950 ;
        RECT 208.950 252.600 211.050 253.050 ;
        RECT 241.950 252.600 244.050 253.050 ;
        RECT 208.950 251.400 244.050 252.600 ;
        RECT 208.950 250.950 211.050 251.400 ;
        RECT 241.950 250.950 244.050 251.400 ;
        RECT 250.950 252.600 253.050 253.050 ;
        RECT 304.950 252.600 307.050 253.050 ;
        RECT 340.950 252.600 343.050 253.050 ;
        RECT 250.950 251.400 343.050 252.600 ;
        RECT 358.950 252.600 361.050 256.050 ;
        RECT 394.950 255.600 397.050 256.050 ;
        RECT 406.950 255.600 409.050 256.050 ;
        RECT 394.950 254.400 409.050 255.600 ;
        RECT 394.950 253.950 397.050 254.400 ;
        RECT 406.950 253.950 409.050 254.400 ;
        RECT 427.950 255.600 430.050 256.200 ;
        RECT 439.950 255.600 442.050 256.050 ;
        RECT 427.950 254.400 442.050 255.600 ;
        RECT 427.950 254.100 430.050 254.400 ;
        RECT 439.950 253.950 442.050 254.400 ;
        RECT 460.950 255.600 463.050 256.050 ;
        RECT 475.950 255.600 478.050 256.050 ;
        RECT 460.950 254.400 478.050 255.600 ;
        RECT 460.950 253.950 463.050 254.400 ;
        RECT 475.950 253.950 478.050 254.400 ;
        RECT 517.950 255.600 520.050 256.050 ;
        RECT 553.950 255.600 556.050 256.050 ;
        RECT 577.950 255.600 580.050 256.050 ;
        RECT 517.950 254.400 556.050 255.600 ;
        RECT 517.950 253.950 520.050 254.400 ;
        RECT 553.950 253.950 556.050 254.400 ;
        RECT 563.400 254.400 580.050 255.600 ;
        RECT 563.400 253.050 564.600 254.400 ;
        RECT 577.950 253.950 580.050 254.400 ;
        RECT 604.950 253.950 610.050 256.050 ;
        RECT 652.950 255.600 655.050 259.050 ;
        RECT 682.950 258.600 685.050 259.050 ;
        RECT 706.800 258.600 708.900 259.050 ;
        RECT 682.950 257.400 708.900 258.600 ;
        RECT 682.950 256.950 685.050 257.400 ;
        RECT 706.800 256.950 708.900 257.400 ;
        RECT 710.100 258.600 712.200 259.200 ;
        RECT 715.950 258.600 718.050 259.050 ;
        RECT 710.100 257.400 718.050 258.600 ;
        RECT 710.100 257.100 712.200 257.400 ;
        RECT 715.950 256.950 718.050 257.400 ;
        RECT 772.950 258.600 775.050 259.050 ;
        RECT 784.950 258.600 787.050 259.200 ;
        RECT 772.950 257.400 787.050 258.600 ;
        RECT 772.950 256.950 775.050 257.400 ;
        RECT 784.950 257.100 787.050 257.400 ;
        RECT 644.400 255.000 655.050 255.600 ;
        RECT 679.950 255.600 682.050 256.050 ;
        RECT 688.950 255.600 691.050 256.050 ;
        RECT 727.950 255.600 730.050 256.050 ;
        RECT 742.950 255.600 745.050 256.050 ;
        RECT 643.950 254.400 654.600 255.000 ;
        RECT 679.950 254.400 691.050 255.600 ;
        RECT 370.950 252.600 373.050 253.050 ;
        RECT 391.950 252.600 394.050 253.050 ;
        RECT 358.950 252.000 394.050 252.600 ;
        RECT 359.400 251.400 394.050 252.000 ;
        RECT 250.950 250.950 253.050 251.400 ;
        RECT 304.950 250.950 307.050 251.400 ;
        RECT 340.950 250.950 343.050 251.400 ;
        RECT 370.950 250.950 373.050 251.400 ;
        RECT 391.950 250.950 394.050 251.400 ;
        RECT 403.950 252.600 406.050 253.050 ;
        RECT 418.950 252.600 421.050 253.050 ;
        RECT 403.950 251.400 421.050 252.600 ;
        RECT 403.950 250.950 406.050 251.400 ;
        RECT 418.950 250.950 421.050 251.400 ;
        RECT 427.950 252.600 430.050 252.900 ;
        RECT 469.950 252.600 472.050 253.050 ;
        RECT 427.950 251.400 472.050 252.600 ;
        RECT 427.950 250.800 430.050 251.400 ;
        RECT 469.950 250.950 472.050 251.400 ;
        RECT 481.950 252.600 484.050 253.050 ;
        RECT 562.950 252.600 565.050 253.050 ;
        RECT 481.950 251.400 565.050 252.600 ;
        RECT 481.950 250.950 484.050 251.400 ;
        RECT 562.950 250.950 565.050 251.400 ;
        RECT 571.950 252.600 574.050 253.050 ;
        RECT 619.950 252.600 622.050 253.050 ;
        RECT 571.950 251.400 622.050 252.600 ;
        RECT 571.950 250.950 574.050 251.400 ;
        RECT 619.950 250.950 622.050 251.400 ;
        RECT 643.950 250.950 646.050 254.400 ;
        RECT 679.950 253.950 682.050 254.400 ;
        RECT 688.950 253.950 691.050 254.400 ;
        RECT 713.400 254.400 745.050 255.600 ;
        RECT 713.400 253.050 714.600 254.400 ;
        RECT 727.950 253.950 730.050 254.400 ;
        RECT 742.950 253.950 745.050 254.400 ;
        RECT 664.950 252.600 667.050 253.050 ;
        RECT 694.950 252.600 697.050 253.050 ;
        RECT 664.950 251.400 697.050 252.600 ;
        RECT 664.950 250.950 667.050 251.400 ;
        RECT 694.950 250.950 697.050 251.400 ;
        RECT 709.950 251.400 714.600 253.050 ;
        RECT 709.950 250.950 714.000 251.400 ;
        RECT 4.950 249.600 7.050 250.050 ;
        RECT 13.950 249.600 16.050 250.050 ;
        RECT 4.950 248.400 16.050 249.600 ;
        RECT 4.950 247.950 7.050 248.400 ;
        RECT 13.950 247.950 16.050 248.400 ;
        RECT 34.950 249.600 37.050 250.050 ;
        RECT 49.950 249.600 52.050 250.050 ;
        RECT 79.950 249.600 82.050 250.050 ;
        RECT 34.950 248.400 82.050 249.600 ;
        RECT 34.950 247.950 37.050 248.400 ;
        RECT 49.950 247.950 52.050 248.400 ;
        RECT 79.950 247.950 82.050 248.400 ;
        RECT 127.950 249.600 130.050 250.050 ;
        RECT 133.950 249.600 136.050 250.050 ;
        RECT 127.950 248.400 136.050 249.600 ;
        RECT 127.950 247.950 130.050 248.400 ;
        RECT 133.950 247.950 136.050 248.400 ;
        RECT 448.950 249.600 451.050 250.050 ;
        RECT 472.950 249.600 475.050 250.050 ;
        RECT 448.950 248.400 475.050 249.600 ;
        RECT 448.950 247.950 451.050 248.400 ;
        RECT 472.950 247.950 475.050 248.400 ;
        RECT 700.950 249.600 703.050 250.050 ;
        RECT 712.950 249.600 715.050 250.050 ;
        RECT 700.950 248.400 715.050 249.600 ;
        RECT 700.950 247.950 703.050 248.400 ;
        RECT 712.950 247.950 715.050 248.400 ;
        RECT 187.950 246.600 190.050 247.050 ;
        RECT 337.950 246.600 340.050 247.050 ;
        RECT 187.950 245.400 340.050 246.600 ;
        RECT 187.950 244.950 190.050 245.400 ;
        RECT 337.950 244.950 340.050 245.400 ;
        RECT 430.950 246.600 433.050 247.050 ;
        RECT 535.950 246.600 538.050 247.050 ;
        RECT 430.950 245.400 538.050 246.600 ;
        RECT 430.950 244.950 433.050 245.400 ;
        RECT 535.950 244.950 538.050 245.400 ;
        RECT 556.950 246.600 559.050 247.050 ;
        RECT 634.950 246.600 637.050 247.050 ;
        RECT 556.950 245.400 637.050 246.600 ;
        RECT 556.950 244.950 559.050 245.400 ;
        RECT 634.950 244.950 637.050 245.400 ;
        RECT 694.950 246.600 697.050 247.050 ;
        RECT 748.950 246.600 751.050 247.050 ;
        RECT 694.950 245.400 751.050 246.600 ;
        RECT 694.950 244.950 697.050 245.400 ;
        RECT 748.950 244.950 751.050 245.400 ;
        RECT 283.950 243.600 286.050 244.050 ;
        RECT 289.950 243.600 292.050 244.050 ;
        RECT 313.950 243.600 316.050 244.050 ;
        RECT 283.950 242.400 316.050 243.600 ;
        RECT 283.950 241.950 286.050 242.400 ;
        RECT 289.950 241.950 292.050 242.400 ;
        RECT 313.950 241.950 316.050 242.400 ;
        RECT 571.950 243.600 574.050 244.050 ;
        RECT 631.950 243.600 634.050 244.050 ;
        RECT 571.950 242.400 634.050 243.600 ;
        RECT 571.950 241.950 574.050 242.400 ;
        RECT 631.950 241.950 634.050 242.400 ;
        RECT 139.950 240.600 142.050 241.050 ;
        RECT 145.950 240.600 148.050 241.050 ;
        RECT 139.950 239.400 148.050 240.600 ;
        RECT 139.950 238.950 142.050 239.400 ;
        RECT 145.950 238.950 148.050 239.400 ;
        RECT 421.950 240.600 424.050 241.050 ;
        RECT 433.950 240.600 436.050 241.050 ;
        RECT 421.950 239.400 436.050 240.600 ;
        RECT 421.950 238.950 424.050 239.400 ;
        RECT 433.950 238.950 436.050 239.400 ;
        RECT 649.950 240.600 652.050 241.050 ;
        RECT 661.950 240.600 664.050 241.050 ;
        RECT 649.950 239.400 664.050 240.600 ;
        RECT 649.950 238.950 652.050 239.400 ;
        RECT 661.950 238.950 664.050 239.400 ;
        RECT 676.950 240.600 679.050 241.050 ;
        RECT 703.950 240.600 706.050 241.050 ;
        RECT 676.950 239.400 706.050 240.600 ;
        RECT 676.950 238.950 679.050 239.400 ;
        RECT 703.950 238.950 706.050 239.400 ;
        RECT 730.950 240.600 733.050 241.050 ;
        RECT 751.950 240.600 754.050 241.050 ;
        RECT 730.950 239.400 754.050 240.600 ;
        RECT 730.950 238.950 733.050 239.400 ;
        RECT 751.950 238.950 754.050 239.400 ;
        RECT 241.950 237.600 244.050 238.050 ;
        RECT 286.950 237.600 289.050 238.050 ;
        RECT 367.950 237.600 370.050 238.050 ;
        RECT 241.950 236.400 289.050 237.600 ;
        RECT 241.950 235.950 244.050 236.400 ;
        RECT 286.950 235.950 289.050 236.400 ;
        RECT 320.400 236.400 370.050 237.600 ;
        RECT 115.950 234.600 118.050 235.050 ;
        RECT 320.400 234.600 321.600 236.400 ;
        RECT 367.950 235.950 370.050 236.400 ;
        RECT 409.950 237.600 412.050 238.050 ;
        RECT 427.800 237.600 429.900 238.050 ;
        RECT 409.950 236.400 429.900 237.600 ;
        RECT 409.950 235.950 412.050 236.400 ;
        RECT 427.800 235.950 429.900 236.400 ;
        RECT 431.100 237.600 433.200 238.050 ;
        RECT 445.950 237.600 448.050 238.050 ;
        RECT 431.100 236.400 448.050 237.600 ;
        RECT 431.100 235.950 433.200 236.400 ;
        RECT 445.950 235.950 448.050 236.400 ;
        RECT 550.950 237.600 553.050 238.050 ;
        RECT 601.950 237.600 604.050 238.050 ;
        RECT 550.950 236.400 604.050 237.600 ;
        RECT 550.950 235.950 553.050 236.400 ;
        RECT 601.950 235.950 604.050 236.400 ;
        RECT 607.950 237.600 610.050 238.050 ;
        RECT 646.950 237.600 649.050 238.050 ;
        RECT 607.950 236.400 649.050 237.600 ;
        RECT 607.950 235.950 610.050 236.400 ;
        RECT 646.950 235.950 649.050 236.400 ;
        RECT 115.950 233.400 321.600 234.600 ;
        RECT 406.950 234.600 409.050 235.050 ;
        RECT 460.950 234.600 463.050 235.050 ;
        RECT 406.950 233.400 463.050 234.600 ;
        RECT 115.950 232.950 118.050 233.400 ;
        RECT 406.950 232.950 409.050 233.400 ;
        RECT 460.950 232.950 463.050 233.400 ;
        RECT 490.950 234.600 493.050 235.050 ;
        RECT 551.400 234.600 552.600 235.950 ;
        RECT 490.950 233.400 552.600 234.600 ;
        RECT 604.950 234.600 607.050 235.050 ;
        RECT 643.950 234.600 646.050 235.050 ;
        RECT 604.950 233.400 646.050 234.600 ;
        RECT 490.950 232.950 493.050 233.400 ;
        RECT 604.950 232.950 607.050 233.400 ;
        RECT 643.950 232.950 646.050 233.400 ;
        RECT 130.950 228.600 133.050 229.050 ;
        RECT 172.950 228.600 175.050 229.050 ;
        RECT 130.950 227.400 175.050 228.600 ;
        RECT 130.950 226.950 133.050 227.400 ;
        RECT 172.950 226.950 175.050 227.400 ;
        RECT 283.950 228.600 286.050 229.050 ;
        RECT 328.950 228.600 331.050 229.050 ;
        RECT 283.950 227.400 331.050 228.600 ;
        RECT 283.950 226.950 286.050 227.400 ;
        RECT 328.950 226.950 331.050 227.400 ;
        RECT 358.950 228.600 361.050 229.050 ;
        RECT 370.950 228.600 373.050 229.050 ;
        RECT 358.950 227.400 373.050 228.600 ;
        RECT 358.950 226.950 361.050 227.400 ;
        RECT 370.950 226.950 373.050 227.400 ;
        RECT 535.950 228.600 538.050 229.050 ;
        RECT 598.950 228.600 601.050 229.050 ;
        RECT 535.950 227.400 601.050 228.600 ;
        RECT 535.950 226.950 538.050 227.400 ;
        RECT 598.950 226.950 601.050 227.400 ;
        RECT 631.950 228.600 634.050 229.050 ;
        RECT 676.950 228.600 679.050 229.050 ;
        RECT 631.950 227.400 679.050 228.600 ;
        RECT 631.950 226.950 634.050 227.400 ;
        RECT 676.950 226.950 679.050 227.400 ;
        RECT 688.950 228.600 691.050 229.050 ;
        RECT 697.950 228.600 700.050 229.050 ;
        RECT 688.950 227.400 700.050 228.600 ;
        RECT 688.950 226.950 691.050 227.400 ;
        RECT 697.950 226.950 700.050 227.400 ;
        RECT 448.950 225.600 451.050 226.050 ;
        RECT 493.950 225.600 496.050 226.050 ;
        RECT 448.950 224.400 496.050 225.600 ;
        RECT 448.950 223.950 451.050 224.400 ;
        RECT 493.950 223.950 496.050 224.400 ;
        RECT 610.950 225.600 613.050 226.050 ;
        RECT 616.950 225.600 619.050 226.050 ;
        RECT 700.950 225.600 703.050 226.050 ;
        RECT 610.950 224.400 703.050 225.600 ;
        RECT 610.950 223.950 613.050 224.400 ;
        RECT 616.950 223.950 619.050 224.400 ;
        RECT 700.950 223.950 703.050 224.400 ;
        RECT 67.950 222.600 70.050 223.050 ;
        RECT 73.950 222.600 76.050 223.050 ;
        RECT 67.950 221.400 76.050 222.600 ;
        RECT 67.950 220.950 70.050 221.400 ;
        RECT 73.950 220.950 76.050 221.400 ;
        RECT 88.950 222.600 91.050 223.050 ;
        RECT 109.950 222.600 112.050 223.050 ;
        RECT 88.950 221.400 112.050 222.600 ;
        RECT 88.950 220.950 91.050 221.400 ;
        RECT 109.950 220.950 112.050 221.400 ;
        RECT 127.950 222.600 130.050 223.050 ;
        RECT 157.950 222.600 160.050 223.050 ;
        RECT 175.950 222.600 178.050 223.050 ;
        RECT 127.950 221.400 178.050 222.600 ;
        RECT 127.950 220.950 130.050 221.400 ;
        RECT 157.950 220.950 160.050 221.400 ;
        RECT 175.950 220.950 178.050 221.400 ;
        RECT 211.950 222.600 214.050 223.050 ;
        RECT 229.950 222.600 232.050 223.050 ;
        RECT 286.950 222.600 289.050 223.050 ;
        RECT 211.950 221.400 289.050 222.600 ;
        RECT 211.950 220.950 214.050 221.400 ;
        RECT 229.950 220.950 232.050 221.400 ;
        RECT 286.950 220.950 289.050 221.400 ;
        RECT 355.950 222.600 358.050 223.200 ;
        RECT 361.950 222.600 364.050 223.050 ;
        RECT 355.950 221.400 364.050 222.600 ;
        RECT 355.950 221.100 358.050 221.400 ;
        RECT 361.950 220.950 364.050 221.400 ;
        RECT 370.950 222.600 373.050 223.050 ;
        RECT 424.950 222.600 427.050 223.050 ;
        RECT 370.950 221.400 427.050 222.600 ;
        RECT 370.950 220.950 373.050 221.400 ;
        RECT 424.950 220.950 427.050 221.400 ;
        RECT 622.950 222.600 625.050 223.050 ;
        RECT 637.950 222.600 640.050 223.050 ;
        RECT 622.950 221.400 640.050 222.600 ;
        RECT 622.950 220.950 625.050 221.400 ;
        RECT 637.950 220.950 640.050 221.400 ;
        RECT 691.950 222.600 694.050 223.050 ;
        RECT 730.950 222.600 733.050 223.050 ;
        RECT 691.950 221.400 733.050 222.600 ;
        RECT 691.950 220.950 694.050 221.400 ;
        RECT 730.950 220.950 733.050 221.400 ;
        RECT 37.950 219.600 40.050 220.050 ;
        RECT 49.950 219.600 52.050 220.050 ;
        RECT 37.950 218.400 52.050 219.600 ;
        RECT 37.950 217.950 40.050 218.400 ;
        RECT 49.950 217.950 52.050 218.400 ;
        RECT 262.950 219.600 265.050 220.200 ;
        RECT 268.950 219.600 271.050 220.050 ;
        RECT 262.950 218.400 271.050 219.600 ;
        RECT 262.950 218.100 265.050 218.400 ;
        RECT 268.950 217.950 271.050 218.400 ;
        RECT 466.950 219.600 469.050 220.050 ;
        RECT 484.950 219.600 487.050 220.050 ;
        RECT 499.950 219.600 502.050 220.050 ;
        RECT 466.950 218.400 502.050 219.600 ;
        RECT 466.950 217.950 469.050 218.400 ;
        RECT 484.950 217.950 487.050 218.400 ;
        RECT 499.950 217.950 502.050 218.400 ;
        RECT 574.950 219.600 577.050 220.050 ;
        RECT 682.950 219.600 685.050 220.050 ;
        RECT 574.950 218.400 685.050 219.600 ;
        RECT 574.950 217.950 577.050 218.400 ;
        RECT 682.950 217.950 685.050 218.400 ;
        RECT 739.950 219.600 742.050 220.050 ;
        RECT 754.800 219.600 756.900 220.050 ;
        RECT 739.950 218.400 756.900 219.600 ;
        RECT 739.950 217.950 742.050 218.400 ;
        RECT 754.800 217.950 756.900 218.400 ;
        RECT 758.100 219.600 760.200 220.050 ;
        RECT 781.950 219.600 784.050 220.050 ;
        RECT 758.100 218.400 784.050 219.600 ;
        RECT 758.100 217.950 760.200 218.400 ;
        RECT 781.950 217.950 784.050 218.400 ;
        RECT 790.950 219.600 793.050 220.200 ;
        RECT 796.950 219.600 799.050 220.050 ;
        RECT 790.950 218.400 799.050 219.600 ;
        RECT 790.950 218.100 793.050 218.400 ;
        RECT 796.950 217.950 799.050 218.400 ;
        RECT 1.950 216.600 4.050 217.050 ;
        RECT 10.950 216.600 13.050 217.050 ;
        RECT 1.950 215.400 13.050 216.600 ;
        RECT 1.950 214.950 4.050 215.400 ;
        RECT 10.950 214.950 13.050 215.400 ;
        RECT 67.950 216.600 70.050 217.050 ;
        RECT 82.950 216.600 85.050 217.200 ;
        RECT 67.950 215.400 85.050 216.600 ;
        RECT 67.950 214.950 70.050 215.400 ;
        RECT 82.950 215.100 85.050 215.400 ;
        RECT 172.950 216.600 175.050 217.050 ;
        RECT 181.950 216.600 184.050 217.050 ;
        RECT 172.950 215.400 184.050 216.600 ;
        RECT 172.950 214.950 175.050 215.400 ;
        RECT 181.950 214.950 184.050 215.400 ;
        RECT 193.950 214.950 199.050 217.050 ;
        RECT 202.950 216.600 205.050 217.050 ;
        RECT 220.950 216.600 223.050 217.050 ;
        RECT 202.950 215.400 223.050 216.600 ;
        RECT 202.950 214.950 205.050 215.400 ;
        RECT 220.950 214.950 223.050 215.400 ;
        RECT 232.950 216.600 235.050 217.050 ;
        RECT 262.950 216.600 265.050 216.900 ;
        RECT 273.000 216.600 277.050 217.050 ;
        RECT 232.950 215.400 265.050 216.600 ;
        RECT 232.950 214.950 235.050 215.400 ;
        RECT 262.950 214.800 265.050 215.400 ;
        RECT 272.400 214.950 277.050 216.600 ;
        RECT 292.950 216.600 295.050 217.050 ;
        RECT 298.950 216.600 301.050 217.050 ;
        RECT 292.950 215.400 301.050 216.600 ;
        RECT 292.950 214.950 295.050 215.400 ;
        RECT 298.950 214.950 301.050 215.400 ;
        RECT 325.950 216.600 328.050 217.050 ;
        RECT 373.950 216.600 376.050 217.050 ;
        RECT 325.950 215.400 376.050 216.600 ;
        RECT 325.950 214.950 328.050 215.400 ;
        RECT 373.950 214.950 376.050 215.400 ;
        RECT 418.950 216.600 421.050 217.050 ;
        RECT 433.950 216.600 436.050 217.050 ;
        RECT 418.950 215.400 436.050 216.600 ;
        RECT 418.950 214.950 421.050 215.400 ;
        RECT 433.950 214.950 436.050 215.400 ;
        RECT 508.950 216.600 511.050 217.200 ;
        RECT 520.950 216.600 523.050 217.050 ;
        RECT 508.950 215.400 523.050 216.600 ;
        RECT 508.950 215.100 511.050 215.400 ;
        RECT 520.950 214.950 523.050 215.400 ;
        RECT 655.950 216.600 658.050 217.050 ;
        RECT 670.950 216.600 673.050 217.050 ;
        RECT 655.950 215.400 673.050 216.600 ;
        RECT 655.950 214.950 658.050 215.400 ;
        RECT 670.950 214.950 673.050 215.400 ;
        RECT 697.950 216.600 700.050 217.050 ;
        RECT 706.950 216.600 709.050 217.050 ;
        RECT 697.950 215.400 709.050 216.600 ;
        RECT 697.950 214.950 700.050 215.400 ;
        RECT 706.950 214.950 709.050 215.400 ;
        RECT 733.950 216.600 736.050 217.050 ;
        RECT 778.950 216.600 781.050 217.200 ;
        RECT 733.950 215.400 781.050 216.600 ;
        RECT 733.950 214.950 736.050 215.400 ;
        RECT 778.950 215.100 781.050 215.400 ;
        RECT 94.950 213.600 97.050 214.050 ;
        RECT 103.950 213.600 106.050 214.200 ;
        RECT 94.950 212.400 106.050 213.600 ;
        RECT 94.950 211.950 97.050 212.400 ;
        RECT 103.950 212.100 106.050 212.400 ;
        RECT 223.950 213.600 226.050 214.050 ;
        RECT 272.400 213.600 273.600 214.950 ;
        RECT 223.950 212.400 273.600 213.600 ;
        RECT 283.950 213.600 286.050 213.900 ;
        RECT 289.950 213.600 292.050 214.200 ;
        RECT 283.950 212.400 292.050 213.600 ;
        RECT 223.950 211.950 226.050 212.400 ;
        RECT 283.950 211.800 286.050 212.400 ;
        RECT 289.950 212.100 292.050 212.400 ;
        RECT 496.950 213.600 499.050 214.050 ;
        RECT 508.950 213.600 511.050 213.900 ;
        RECT 496.950 212.400 511.050 213.600 ;
        RECT 496.950 211.950 499.050 212.400 ;
        RECT 508.950 211.800 511.050 212.400 ;
        RECT 565.950 213.600 568.050 214.050 ;
        RECT 571.950 213.600 574.050 214.050 ;
        RECT 565.950 212.400 574.050 213.600 ;
        RECT 565.950 211.950 568.050 212.400 ;
        RECT 571.950 211.950 574.050 212.400 ;
        RECT 613.950 213.600 616.050 214.050 ;
        RECT 751.950 213.600 754.050 214.050 ;
        RECT 613.950 212.400 754.050 213.600 ;
        RECT 613.950 211.950 616.050 212.400 ;
        RECT 751.950 211.950 754.050 212.400 ;
        RECT 760.950 213.600 763.050 214.050 ;
        RECT 781.950 213.600 784.050 214.050 ;
        RECT 760.950 212.400 784.050 213.600 ;
        RECT 760.950 211.950 763.050 212.400 ;
        RECT 781.950 211.950 784.050 212.400 ;
        RECT 1.950 210.600 4.050 211.050 ;
        RECT 13.950 210.600 16.050 211.050 ;
        RECT 1.950 209.400 16.050 210.600 ;
        RECT 1.950 208.950 4.050 209.400 ;
        RECT 13.950 208.950 16.050 209.400 ;
        RECT 25.950 210.600 28.050 211.050 ;
        RECT 46.950 210.600 49.050 211.050 ;
        RECT 25.950 209.400 49.050 210.600 ;
        RECT 25.950 208.950 28.050 209.400 ;
        RECT 46.950 208.950 49.050 209.400 ;
        RECT 103.950 210.600 106.050 210.900 ;
        RECT 115.950 210.600 118.050 211.050 ;
        RECT 103.950 209.400 118.050 210.600 ;
        RECT 103.950 208.800 106.050 209.400 ;
        RECT 115.950 208.950 118.050 209.400 ;
        RECT 136.950 210.600 139.050 211.050 ;
        RECT 148.950 210.600 151.050 211.050 ;
        RECT 136.950 209.400 151.050 210.600 ;
        RECT 136.950 208.950 139.050 209.400 ;
        RECT 148.950 208.950 151.050 209.400 ;
        RECT 163.950 210.600 166.050 211.050 ;
        RECT 205.950 210.600 208.050 211.050 ;
        RECT 214.950 210.600 217.050 211.050 ;
        RECT 163.950 209.400 217.050 210.600 ;
        RECT 163.950 208.950 166.050 209.400 ;
        RECT 205.950 208.950 208.050 209.400 ;
        RECT 214.950 208.950 217.050 209.400 ;
        RECT 256.950 210.600 259.050 211.050 ;
        RECT 277.950 210.600 280.050 211.050 ;
        RECT 256.950 209.400 280.050 210.600 ;
        RECT 256.950 208.950 259.050 209.400 ;
        RECT 277.950 208.950 280.050 209.400 ;
        RECT 397.950 210.600 400.050 211.050 ;
        RECT 406.950 210.600 412.050 211.050 ;
        RECT 397.950 209.400 412.050 210.600 ;
        RECT 397.950 208.950 400.050 209.400 ;
        RECT 406.950 208.950 412.050 209.400 ;
        RECT 484.950 208.950 490.050 211.050 ;
        RECT 550.950 210.600 553.050 211.050 ;
        RECT 556.950 210.600 559.050 211.050 ;
        RECT 550.950 209.400 559.050 210.600 ;
        RECT 550.950 208.950 553.050 209.400 ;
        RECT 556.950 208.950 559.050 209.400 ;
        RECT 631.950 210.600 634.050 211.050 ;
        RECT 667.950 210.600 670.050 211.050 ;
        RECT 718.950 210.600 721.050 211.050 ;
        RECT 631.950 209.400 670.050 210.600 ;
        RECT 713.400 210.000 721.050 210.600 ;
        RECT 631.950 208.950 634.050 209.400 ;
        RECT 667.950 208.950 670.050 209.400 ;
        RECT 712.950 209.400 721.050 210.000 ;
        RECT 154.950 207.600 157.050 208.050 ;
        RECT 172.950 207.600 175.050 208.050 ;
        RECT 154.950 206.400 175.050 207.600 ;
        RECT 154.950 205.950 157.050 206.400 ;
        RECT 172.950 205.950 175.050 206.400 ;
        RECT 340.950 207.600 343.050 208.050 ;
        RECT 349.950 207.600 352.050 208.050 ;
        RECT 385.950 207.600 388.050 208.050 ;
        RECT 340.950 206.400 388.050 207.600 ;
        RECT 340.950 205.950 343.050 206.400 ;
        RECT 349.950 205.950 352.050 206.400 ;
        RECT 385.950 205.950 388.050 206.400 ;
        RECT 616.950 207.600 619.050 208.050 ;
        RECT 622.950 207.600 625.050 208.050 ;
        RECT 616.950 206.400 625.050 207.600 ;
        RECT 616.950 205.950 619.050 206.400 ;
        RECT 622.950 205.950 625.050 206.400 ;
        RECT 703.950 207.600 706.050 208.050 ;
        RECT 712.950 207.600 715.050 209.400 ;
        RECT 718.950 208.950 721.050 209.400 ;
        RECT 736.950 210.600 739.050 211.050 ;
        RECT 787.950 210.600 790.050 211.050 ;
        RECT 811.950 210.600 814.050 211.200 ;
        RECT 736.950 210.000 744.600 210.600 ;
        RECT 736.950 209.400 745.050 210.000 ;
        RECT 736.950 208.950 739.050 209.400 ;
        RECT 703.950 206.400 715.050 207.600 ;
        RECT 703.950 205.950 706.050 206.400 ;
        RECT 712.950 205.950 715.050 206.400 ;
        RECT 742.950 205.950 745.050 209.400 ;
        RECT 787.950 209.400 814.050 210.600 ;
        RECT 787.950 208.950 790.050 209.400 ;
        RECT 811.950 209.100 814.050 209.400 ;
        RECT 220.950 204.600 223.050 205.050 ;
        RECT 232.950 204.600 235.050 205.050 ;
        RECT 220.950 203.400 235.050 204.600 ;
        RECT 220.950 202.950 223.050 203.400 ;
        RECT 232.950 202.950 235.050 203.400 ;
        RECT 304.950 204.600 307.050 205.050 ;
        RECT 325.950 204.600 328.050 205.050 ;
        RECT 304.950 203.400 328.050 204.600 ;
        RECT 304.950 202.950 307.050 203.400 ;
        RECT 325.950 202.950 328.050 203.400 ;
        RECT 451.950 204.600 454.050 205.050 ;
        RECT 493.950 204.600 496.050 205.050 ;
        RECT 451.950 203.400 496.050 204.600 ;
        RECT 451.950 202.950 454.050 203.400 ;
        RECT 493.950 202.950 496.050 203.400 ;
        RECT 226.950 201.600 229.050 202.050 ;
        RECT 253.950 201.600 256.050 202.050 ;
        RECT 289.950 201.600 292.050 202.050 ;
        RECT 226.950 200.400 292.050 201.600 ;
        RECT 226.950 199.950 229.050 200.400 ;
        RECT 253.950 199.950 256.050 200.400 ;
        RECT 289.950 199.950 292.050 200.400 ;
        RECT 601.950 201.600 604.050 202.050 ;
        RECT 634.950 201.600 637.050 202.050 ;
        RECT 601.950 200.400 637.050 201.600 ;
        RECT 601.950 199.950 604.050 200.400 ;
        RECT 634.950 199.950 637.050 200.400 ;
        RECT 703.950 201.600 706.050 202.050 ;
        RECT 772.950 201.600 775.050 202.050 ;
        RECT 703.950 200.400 775.050 201.600 ;
        RECT 703.950 199.950 706.050 200.400 ;
        RECT 772.950 199.950 775.050 200.400 ;
        RECT 166.950 198.600 169.050 199.050 ;
        RECT 181.950 198.600 184.050 199.050 ;
        RECT 217.950 198.600 220.050 199.050 ;
        RECT 166.950 197.400 220.050 198.600 ;
        RECT 166.950 196.950 169.050 197.400 ;
        RECT 181.950 196.950 184.050 197.400 ;
        RECT 217.950 196.950 220.050 197.400 ;
        RECT 307.950 198.600 310.050 199.050 ;
        RECT 529.950 198.600 532.050 199.050 ;
        RECT 574.950 198.600 577.050 199.050 ;
        RECT 307.950 197.400 577.050 198.600 ;
        RECT 307.950 196.950 310.050 197.400 ;
        RECT 529.950 196.950 532.050 197.400 ;
        RECT 574.950 196.950 577.050 197.400 ;
        RECT 595.950 198.600 598.050 199.050 ;
        RECT 763.950 198.600 766.050 199.050 ;
        RECT 793.950 198.600 796.050 199.050 ;
        RECT 595.950 197.400 796.050 198.600 ;
        RECT 595.950 196.950 598.050 197.400 ;
        RECT 763.950 196.950 766.050 197.400 ;
        RECT 793.950 196.950 796.050 197.400 ;
        RECT 67.950 195.600 70.050 196.050 ;
        RECT 88.950 195.600 91.050 196.050 ;
        RECT 67.950 194.400 91.050 195.600 ;
        RECT 67.950 193.950 70.050 194.400 ;
        RECT 88.950 193.950 91.050 194.400 ;
        RECT 100.950 195.600 103.050 196.050 ;
        RECT 130.950 195.600 133.050 196.050 ;
        RECT 100.950 194.400 133.050 195.600 ;
        RECT 100.950 193.950 103.050 194.400 ;
        RECT 130.950 193.950 133.050 194.400 ;
        RECT 271.950 195.600 274.050 196.050 ;
        RECT 295.950 195.600 298.050 196.050 ;
        RECT 271.950 194.400 298.050 195.600 ;
        RECT 271.950 193.950 274.050 194.400 ;
        RECT 295.950 193.950 298.050 194.400 ;
        RECT 589.950 195.600 592.050 196.050 ;
        RECT 622.950 195.600 625.050 196.050 ;
        RECT 589.950 194.400 625.050 195.600 ;
        RECT 589.950 193.950 592.050 194.400 ;
        RECT 622.950 193.950 625.050 194.400 ;
        RECT 34.950 192.600 37.050 193.050 ;
        RECT 61.950 192.600 64.050 193.050 ;
        RECT 34.950 191.400 64.050 192.600 ;
        RECT 34.950 190.950 37.050 191.400 ;
        RECT 61.950 190.950 64.050 191.400 ;
        RECT 193.950 192.600 196.050 193.050 ;
        RECT 220.950 192.600 223.050 193.050 ;
        RECT 193.950 191.400 223.050 192.600 ;
        RECT 193.950 190.950 196.050 191.400 ;
        RECT 220.950 190.950 223.050 191.400 ;
        RECT 388.950 192.600 391.050 193.050 ;
        RECT 421.950 192.600 424.050 193.050 ;
        RECT 388.950 191.400 424.050 192.600 ;
        RECT 388.950 190.950 391.050 191.400 ;
        RECT 421.950 190.950 424.050 191.400 ;
        RECT 529.950 192.600 532.050 193.050 ;
        RECT 553.950 192.600 556.050 193.050 ;
        RECT 529.950 191.400 556.050 192.600 ;
        RECT 529.950 190.950 532.050 191.400 ;
        RECT 553.950 190.950 556.050 191.400 ;
        RECT 631.950 192.600 634.050 193.050 ;
        RECT 736.950 192.600 739.050 193.050 ;
        RECT 631.950 191.400 739.050 192.600 ;
        RECT 631.950 190.950 634.050 191.400 ;
        RECT 736.950 190.950 739.050 191.400 ;
        RECT 70.950 189.600 73.050 190.050 ;
        RECT 100.950 189.600 103.050 190.050 ;
        RECT 70.950 188.400 103.050 189.600 ;
        RECT 70.950 187.950 73.050 188.400 ;
        RECT 100.950 187.950 103.050 188.400 ;
        RECT 142.950 189.600 145.050 190.050 ;
        RECT 169.950 189.600 172.050 190.050 ;
        RECT 142.950 188.400 172.050 189.600 ;
        RECT 142.950 187.950 145.050 188.400 ;
        RECT 169.950 187.950 172.050 188.400 ;
        RECT 214.950 189.600 219.000 190.050 ;
        RECT 367.950 189.600 370.050 190.050 ;
        RECT 451.950 189.600 454.050 190.050 ;
        RECT 214.950 187.950 219.600 189.600 ;
        RECT 367.950 188.400 454.050 189.600 ;
        RECT 367.950 187.950 370.050 188.400 ;
        RECT 451.950 187.950 454.050 188.400 ;
        RECT 523.950 189.600 526.050 190.050 ;
        RECT 556.950 189.600 559.050 190.050 ;
        RECT 523.950 188.400 559.050 189.600 ;
        RECT 523.950 187.950 526.050 188.400 ;
        RECT 556.950 187.950 559.050 188.400 ;
        RECT 604.950 189.600 607.050 190.050 ;
        RECT 643.950 189.600 646.050 190.050 ;
        RECT 604.950 188.400 646.050 189.600 ;
        RECT 604.950 187.950 607.050 188.400 ;
        RECT 643.950 187.950 646.050 188.400 ;
        RECT 751.950 189.600 754.050 190.050 ;
        RECT 769.950 189.600 772.050 190.050 ;
        RECT 775.950 189.600 778.050 190.050 ;
        RECT 751.950 188.400 778.050 189.600 ;
        RECT 751.950 187.950 754.050 188.400 ;
        RECT 769.950 187.950 772.050 188.400 ;
        RECT 775.950 187.950 778.050 188.400 ;
        RECT 43.950 183.600 46.050 184.050 ;
        RECT 55.950 183.600 58.050 187.050 ;
        RECT 82.950 186.600 85.050 187.050 ;
        RECT 112.950 186.600 115.050 187.050 ;
        RECT 82.950 185.400 115.050 186.600 ;
        RECT 82.950 184.950 85.050 185.400 ;
        RECT 112.950 184.950 115.050 185.400 ;
        RECT 151.950 186.600 154.050 187.050 ;
        RECT 211.950 186.600 214.050 187.050 ;
        RECT 151.950 185.400 214.050 186.600 ;
        RECT 218.400 186.600 219.600 187.950 ;
        RECT 295.950 186.600 298.050 187.050 ;
        RECT 218.400 185.400 298.050 186.600 ;
        RECT 151.950 184.950 154.050 185.400 ;
        RECT 211.950 184.950 214.050 185.400 ;
        RECT 295.950 184.950 298.050 185.400 ;
        RECT 526.950 186.600 529.050 187.050 ;
        RECT 532.950 186.600 535.050 187.050 ;
        RECT 526.950 185.400 535.050 186.600 ;
        RECT 526.950 184.950 529.050 185.400 ;
        RECT 532.950 184.950 535.050 185.400 ;
        RECT 568.950 186.600 571.050 187.050 ;
        RECT 595.950 186.600 598.050 187.050 ;
        RECT 568.950 185.400 598.050 186.600 ;
        RECT 568.950 184.950 571.050 185.400 ;
        RECT 595.950 184.950 598.050 185.400 ;
        RECT 43.950 183.000 58.050 183.600 ;
        RECT 73.950 183.600 76.050 184.200 ;
        RECT 91.950 183.600 94.050 184.050 ;
        RECT 43.950 182.400 57.600 183.000 ;
        RECT 73.950 182.400 94.050 183.600 ;
        RECT 43.950 181.950 46.050 182.400 ;
        RECT 73.950 182.100 76.050 182.400 ;
        RECT 91.950 181.950 94.050 182.400 ;
        RECT 169.950 181.950 175.050 184.050 ;
        RECT 301.950 183.600 304.050 184.050 ;
        RECT 307.950 183.600 310.050 184.050 ;
        RECT 301.950 182.400 310.050 183.600 ;
        RECT 301.950 181.950 304.050 182.400 ;
        RECT 307.950 181.950 310.050 182.400 ;
        RECT 340.950 183.600 343.050 184.200 ;
        RECT 355.950 183.600 358.050 184.050 ;
        RECT 340.950 182.400 358.050 183.600 ;
        RECT 340.950 182.100 343.050 182.400 ;
        RECT 355.950 181.950 358.050 182.400 ;
        RECT 376.950 183.600 379.050 184.050 ;
        RECT 403.950 183.600 408.000 184.050 ;
        RECT 424.950 183.600 427.050 184.050 ;
        RECT 430.950 183.600 433.050 184.200 ;
        RECT 376.950 182.400 408.600 183.600 ;
        RECT 424.950 182.400 433.050 183.600 ;
        RECT 376.950 181.950 379.050 182.400 ;
        RECT 403.950 181.950 408.000 182.400 ;
        RECT 424.950 181.950 427.050 182.400 ;
        RECT 430.950 182.100 433.050 182.400 ;
        RECT 514.950 183.600 517.050 184.050 ;
        RECT 535.950 183.600 538.050 184.050 ;
        RECT 514.950 182.400 538.050 183.600 ;
        RECT 514.950 181.950 517.050 182.400 ;
        RECT 535.950 181.950 538.050 182.400 ;
        RECT 604.950 183.600 607.050 184.050 ;
        RECT 616.950 183.600 619.050 184.050 ;
        RECT 604.950 182.400 619.050 183.600 ;
        RECT 664.950 183.600 667.050 187.050 ;
        RECT 679.950 186.600 682.050 187.050 ;
        RECT 688.950 186.600 691.050 187.050 ;
        RECT 679.950 185.400 691.050 186.600 ;
        RECT 679.950 184.950 682.050 185.400 ;
        RECT 688.950 184.950 691.050 185.400 ;
        RECT 772.950 186.600 775.050 187.050 ;
        RECT 790.950 186.600 793.050 187.050 ;
        RECT 772.950 185.400 793.050 186.600 ;
        RECT 772.950 184.950 775.050 185.400 ;
        RECT 790.950 184.950 793.050 185.400 ;
        RECT 703.950 183.600 706.050 184.050 ;
        RECT 664.950 183.000 706.050 183.600 ;
        RECT 665.400 182.400 706.050 183.000 ;
        RECT 604.950 181.950 607.050 182.400 ;
        RECT 616.950 181.950 619.050 182.400 ;
        RECT 703.950 181.950 706.050 182.400 ;
        RECT 754.950 183.600 757.050 184.050 ;
        RECT 808.950 183.600 811.050 184.050 ;
        RECT 754.950 182.400 811.050 183.600 ;
        RECT 754.950 181.950 757.050 182.400 ;
        RECT 808.950 181.950 811.050 182.400 ;
        RECT 7.950 177.600 10.050 178.050 ;
        RECT 43.950 177.600 46.050 178.050 ;
        RECT 7.950 176.400 46.050 177.600 ;
        RECT 58.950 177.600 61.050 181.050 ;
        RECT 79.950 180.600 82.050 181.050 ;
        RECT 85.950 180.600 88.050 181.050 ;
        RECT 79.950 179.400 88.050 180.600 ;
        RECT 79.950 178.950 82.050 179.400 ;
        RECT 85.950 178.950 88.050 179.400 ;
        RECT 127.950 180.600 130.050 181.050 ;
        RECT 190.950 180.600 193.050 181.050 ;
        RECT 226.950 180.600 229.050 181.050 ;
        RECT 127.950 179.400 229.050 180.600 ;
        RECT 127.950 178.950 130.050 179.400 ;
        RECT 190.950 178.950 193.050 179.400 ;
        RECT 226.950 178.950 229.050 179.400 ;
        RECT 232.950 180.600 235.050 181.050 ;
        RECT 271.950 180.600 274.050 181.050 ;
        RECT 232.950 179.400 274.050 180.600 ;
        RECT 232.950 178.950 235.050 179.400 ;
        RECT 271.950 178.950 274.050 179.400 ;
        RECT 286.950 180.600 289.050 181.200 ;
        RECT 313.950 180.600 316.050 181.050 ;
        RECT 286.950 179.400 316.050 180.600 ;
        RECT 286.950 179.100 289.050 179.400 ;
        RECT 313.950 178.950 316.050 179.400 ;
        RECT 328.950 180.600 331.050 181.200 ;
        RECT 373.950 180.600 376.050 181.050 ;
        RECT 412.950 180.600 415.050 181.050 ;
        RECT 433.950 180.600 436.050 181.200 ;
        RECT 328.950 179.400 436.050 180.600 ;
        RECT 328.950 179.100 331.050 179.400 ;
        RECT 373.950 178.950 376.050 179.400 ;
        RECT 412.950 178.950 415.050 179.400 ;
        RECT 433.950 179.100 436.050 179.400 ;
        RECT 685.950 180.600 688.050 181.050 ;
        RECT 697.950 180.600 700.050 181.200 ;
        RECT 685.950 179.400 700.050 180.600 ;
        RECT 685.950 178.950 688.050 179.400 ;
        RECT 697.950 179.100 700.050 179.400 ;
        RECT 715.950 180.600 718.050 181.050 ;
        RECT 733.950 180.600 736.050 181.050 ;
        RECT 715.950 179.400 736.050 180.600 ;
        RECT 76.950 177.600 79.050 178.050 ;
        RECT 58.950 177.000 79.050 177.600 ;
        RECT 59.400 176.400 79.050 177.000 ;
        RECT 7.950 175.950 10.050 176.400 ;
        RECT 43.950 175.950 46.050 176.400 ;
        RECT 76.950 175.950 79.050 176.400 ;
        RECT 88.950 177.600 91.050 178.050 ;
        RECT 94.950 177.600 97.050 178.050 ;
        RECT 88.950 176.400 97.050 177.600 ;
        RECT 88.950 175.950 91.050 176.400 ;
        RECT 94.950 175.950 97.050 176.400 ;
        RECT 280.950 175.950 286.050 178.050 ;
        RECT 304.950 175.950 310.050 178.050 ;
        RECT 316.950 177.600 319.050 178.050 ;
        RECT 325.950 177.600 328.050 177.900 ;
        RECT 316.950 176.400 328.050 177.600 ;
        RECT 316.950 175.950 319.050 176.400 ;
        RECT 325.950 175.800 328.050 176.400 ;
        RECT 337.950 175.950 342.900 178.050 ;
        RECT 344.100 177.600 346.200 178.050 ;
        RECT 358.950 177.600 361.050 178.050 ;
        RECT 391.950 177.600 394.050 178.050 ;
        RECT 344.100 176.400 394.050 177.600 ;
        RECT 344.100 175.950 346.200 176.400 ;
        RECT 358.950 175.950 361.050 176.400 ;
        RECT 391.950 175.950 394.050 176.400 ;
        RECT 400.950 177.600 403.050 178.050 ;
        RECT 406.950 177.600 409.050 178.050 ;
        RECT 424.950 177.600 427.050 178.050 ;
        RECT 433.950 177.600 436.050 177.900 ;
        RECT 400.950 176.400 436.050 177.600 ;
        RECT 400.950 175.950 403.050 176.400 ;
        RECT 406.950 175.950 409.050 176.400 ;
        RECT 424.950 175.950 427.050 176.400 ;
        RECT 433.950 175.800 436.050 176.400 ;
        RECT 517.950 175.950 523.050 178.050 ;
        RECT 589.950 177.600 592.050 178.050 ;
        RECT 601.950 177.600 604.050 178.050 ;
        RECT 589.950 176.400 604.050 177.600 ;
        RECT 589.950 175.950 592.050 176.400 ;
        RECT 601.950 175.950 604.050 176.400 ;
        RECT 610.950 177.600 613.050 178.050 ;
        RECT 616.950 177.600 619.050 178.050 ;
        RECT 610.950 176.400 619.050 177.600 ;
        RECT 610.950 175.950 613.050 176.400 ;
        RECT 616.950 175.950 619.050 176.400 ;
        RECT 628.950 177.600 631.050 178.050 ;
        RECT 640.950 177.600 643.050 178.050 ;
        RECT 628.950 176.400 643.050 177.600 ;
        RECT 628.950 175.950 631.050 176.400 ;
        RECT 640.950 175.950 643.050 176.400 ;
        RECT 667.950 177.600 670.050 178.050 ;
        RECT 676.950 177.600 679.050 178.050 ;
        RECT 667.950 176.400 679.050 177.600 ;
        RECT 667.950 175.950 670.050 176.400 ;
        RECT 676.950 175.950 679.050 176.400 ;
        RECT 709.950 177.600 712.050 178.050 ;
        RECT 715.950 177.600 718.050 179.400 ;
        RECT 733.950 178.950 736.050 179.400 ;
        RECT 778.950 180.600 781.050 181.050 ;
        RECT 802.950 180.600 805.050 181.050 ;
        RECT 778.950 179.400 805.050 180.600 ;
        RECT 778.950 178.950 781.050 179.400 ;
        RECT 802.950 178.950 805.050 179.400 ;
        RECT 811.950 180.600 814.050 181.050 ;
        RECT 820.950 180.600 823.050 181.050 ;
        RECT 811.950 179.400 823.050 180.600 ;
        RECT 811.950 178.950 814.050 179.400 ;
        RECT 820.950 178.950 823.050 179.400 ;
        RECT 709.950 177.000 718.050 177.600 ;
        RECT 709.950 176.400 717.600 177.000 ;
        RECT 709.950 175.950 712.050 176.400 ;
        RECT 52.950 174.600 55.050 175.050 ;
        RECT 64.950 174.600 67.050 175.050 ;
        RECT 52.950 173.400 67.050 174.600 ;
        RECT 52.950 172.950 55.050 173.400 ;
        RECT 64.950 172.950 67.050 173.400 ;
        RECT 691.950 174.600 694.050 175.050 ;
        RECT 697.950 174.600 700.050 174.900 ;
        RECT 691.950 173.400 700.050 174.600 ;
        RECT 691.950 172.950 694.050 173.400 ;
        RECT 697.950 172.800 700.050 173.400 ;
        RECT 763.950 174.600 766.050 175.050 ;
        RECT 778.950 174.600 781.050 175.050 ;
        RECT 763.950 173.400 781.050 174.600 ;
        RECT 763.950 172.950 766.050 173.400 ;
        RECT 778.950 172.950 781.050 173.400 ;
        RECT 76.950 171.600 79.050 172.050 ;
        RECT 151.950 171.600 154.050 172.050 ;
        RECT 184.950 171.600 187.050 172.050 ;
        RECT 76.950 170.400 187.050 171.600 ;
        RECT 76.950 169.950 79.050 170.400 ;
        RECT 151.950 169.950 154.050 170.400 ;
        RECT 184.950 169.950 187.050 170.400 ;
        RECT 262.950 171.600 265.050 172.050 ;
        RECT 337.950 171.600 340.050 172.050 ;
        RECT 262.950 170.400 340.050 171.600 ;
        RECT 262.950 169.950 265.050 170.400 ;
        RECT 337.950 169.950 340.050 170.400 ;
        RECT 409.950 171.600 412.050 172.050 ;
        RECT 418.950 171.600 421.050 172.050 ;
        RECT 409.950 170.400 421.050 171.600 ;
        RECT 409.950 169.950 412.050 170.400 ;
        RECT 418.950 169.950 421.050 170.400 ;
        RECT 220.950 168.600 223.050 169.050 ;
        RECT 352.950 168.600 355.050 169.050 ;
        RECT 220.950 167.400 355.050 168.600 ;
        RECT 220.950 166.950 223.050 167.400 ;
        RECT 352.950 166.950 355.050 167.400 ;
        RECT 580.950 168.600 583.050 169.050 ;
        RECT 598.950 168.600 601.050 169.050 ;
        RECT 580.950 167.400 601.050 168.600 ;
        RECT 580.950 166.950 583.050 167.400 ;
        RECT 598.950 166.950 601.050 167.400 ;
        RECT 736.950 168.600 739.050 169.050 ;
        RECT 805.950 168.600 808.050 169.050 ;
        RECT 736.950 167.400 808.050 168.600 ;
        RECT 736.950 166.950 739.050 167.400 ;
        RECT 805.950 166.950 808.050 167.400 ;
        RECT 472.950 165.600 475.050 166.050 ;
        RECT 526.950 165.600 529.050 166.050 ;
        RECT 472.950 164.400 529.050 165.600 ;
        RECT 472.950 163.950 475.050 164.400 ;
        RECT 526.950 163.950 529.050 164.400 ;
        RECT 673.950 165.600 676.050 166.050 ;
        RECT 715.950 165.600 718.050 166.050 ;
        RECT 673.950 164.400 718.050 165.600 ;
        RECT 673.950 163.950 676.050 164.400 ;
        RECT 715.950 163.950 718.050 164.400 ;
        RECT 241.950 162.600 244.050 163.050 ;
        RECT 343.950 162.600 346.050 163.050 ;
        RECT 241.950 161.400 346.050 162.600 ;
        RECT 241.950 160.950 244.050 161.400 ;
        RECT 343.950 160.950 346.050 161.400 ;
        RECT 562.950 162.600 565.050 163.050 ;
        RECT 577.950 162.600 580.050 163.050 ;
        RECT 562.950 161.400 580.050 162.600 ;
        RECT 562.950 160.950 565.050 161.400 ;
        RECT 577.950 160.950 580.050 161.400 ;
        RECT 685.950 162.600 688.050 163.050 ;
        RECT 736.950 162.600 739.050 163.050 ;
        RECT 775.950 162.600 778.050 163.050 ;
        RECT 685.950 161.400 778.050 162.600 ;
        RECT 685.950 160.950 688.050 161.400 ;
        RECT 736.950 160.950 739.050 161.400 ;
        RECT 775.950 160.950 778.050 161.400 ;
        RECT 103.950 159.600 106.050 160.050 ;
        RECT 121.950 159.600 124.050 160.050 ;
        RECT 103.950 158.400 124.050 159.600 ;
        RECT 103.950 157.950 106.050 158.400 ;
        RECT 121.950 157.950 124.050 158.400 ;
        RECT 301.950 159.600 304.050 160.050 ;
        RECT 331.950 159.600 334.050 160.050 ;
        RECT 301.950 158.400 334.050 159.600 ;
        RECT 301.950 157.950 304.050 158.400 ;
        RECT 331.950 157.950 334.050 158.400 ;
        RECT 430.950 159.600 433.050 160.050 ;
        RECT 448.950 159.600 451.050 160.050 ;
        RECT 430.950 158.400 451.050 159.600 ;
        RECT 430.950 157.950 433.050 158.400 ;
        RECT 448.950 157.950 451.050 158.400 ;
        RECT 496.950 159.600 499.050 160.050 ;
        RECT 631.950 159.600 634.050 160.050 ;
        RECT 496.950 158.400 634.050 159.600 ;
        RECT 496.950 157.950 499.050 158.400 ;
        RECT 631.950 157.950 634.050 158.400 ;
        RECT 19.950 156.600 22.050 157.050 ;
        RECT 28.950 156.600 31.050 157.050 ;
        RECT 19.950 155.400 31.050 156.600 ;
        RECT 19.950 154.950 22.050 155.400 ;
        RECT 28.950 154.950 31.050 155.400 ;
        RECT 451.950 156.600 454.050 157.050 ;
        RECT 694.950 156.600 697.050 157.050 ;
        RECT 757.950 156.600 760.050 157.050 ;
        RECT 451.950 155.400 760.050 156.600 ;
        RECT 451.950 154.950 454.050 155.400 ;
        RECT 694.950 154.950 697.050 155.400 ;
        RECT 757.950 154.950 760.050 155.400 ;
        RECT 7.950 153.600 10.050 154.050 ;
        RECT 37.950 153.600 40.050 154.050 ;
        RECT 7.950 152.400 40.050 153.600 ;
        RECT 7.950 151.950 10.050 152.400 ;
        RECT 37.950 151.950 40.050 152.400 ;
        RECT 280.950 153.600 283.050 154.050 ;
        RECT 301.950 153.600 304.050 154.050 ;
        RECT 280.950 152.400 304.050 153.600 ;
        RECT 280.950 151.950 283.050 152.400 ;
        RECT 301.950 151.950 304.050 152.400 ;
        RECT 472.950 153.600 475.050 154.050 ;
        RECT 505.950 153.600 508.050 154.050 ;
        RECT 544.950 153.600 547.050 154.050 ;
        RECT 472.950 152.400 547.050 153.600 ;
        RECT 472.950 151.950 475.050 152.400 ;
        RECT 505.950 151.950 508.050 152.400 ;
        RECT 544.950 151.950 547.050 152.400 ;
        RECT 550.950 153.600 553.050 154.050 ;
        RECT 556.950 153.600 559.050 154.050 ;
        RECT 637.950 153.600 640.050 154.050 ;
        RECT 550.950 152.400 640.050 153.600 ;
        RECT 550.950 151.950 553.050 152.400 ;
        RECT 556.950 151.950 559.050 152.400 ;
        RECT 637.950 151.950 640.050 152.400 ;
        RECT 787.950 153.600 790.050 154.050 ;
        RECT 811.950 153.600 814.050 154.050 ;
        RECT 820.950 153.600 823.050 154.050 ;
        RECT 787.950 152.400 823.050 153.600 ;
        RECT 787.950 151.950 790.050 152.400 ;
        RECT 811.950 151.950 814.050 152.400 ;
        RECT 820.950 151.950 823.050 152.400 ;
        RECT 49.950 150.600 52.050 151.050 ;
        RECT 97.950 150.600 100.050 151.050 ;
        RECT 109.950 150.600 112.050 151.050 ;
        RECT 49.950 149.400 112.050 150.600 ;
        RECT 49.950 148.950 52.050 149.400 ;
        RECT 97.950 148.950 100.050 149.400 ;
        RECT 109.950 148.950 112.050 149.400 ;
        RECT 289.950 150.600 292.050 151.050 ;
        RECT 295.950 150.600 298.050 151.050 ;
        RECT 289.950 149.400 298.050 150.600 ;
        RECT 289.950 148.950 292.050 149.400 ;
        RECT 295.950 148.950 298.050 149.400 ;
        RECT 394.950 150.600 397.050 151.050 ;
        RECT 430.950 150.600 433.050 151.050 ;
        RECT 394.950 149.400 433.050 150.600 ;
        RECT 394.950 148.950 397.050 149.400 ;
        RECT 430.950 148.950 433.050 149.400 ;
        RECT 766.950 150.600 769.050 151.050 ;
        RECT 784.950 150.600 787.050 151.050 ;
        RECT 766.950 149.400 787.050 150.600 ;
        RECT 766.950 148.950 769.050 149.400 ;
        RECT 784.950 148.950 787.050 149.400 ;
        RECT 64.950 147.600 67.050 148.050 ;
        RECT 76.950 147.600 79.050 148.050 ;
        RECT 64.950 146.400 79.050 147.600 ;
        RECT 64.950 145.950 67.050 146.400 ;
        RECT 76.950 145.950 79.050 146.400 ;
        RECT 142.950 147.600 145.050 148.050 ;
        RECT 157.950 147.600 160.050 148.050 ;
        RECT 142.950 146.400 160.050 147.600 ;
        RECT 142.950 145.950 145.050 146.400 ;
        RECT 157.950 145.950 160.050 146.400 ;
        RECT 388.950 147.600 391.050 148.050 ;
        RECT 445.950 147.600 448.050 148.050 ;
        RECT 451.950 147.600 454.050 148.050 ;
        RECT 388.950 146.400 399.600 147.600 ;
        RECT 388.950 145.950 391.050 146.400 ;
        RECT 88.950 144.600 91.050 145.050 ;
        RECT 127.950 144.600 130.050 145.050 ;
        RECT 88.950 143.400 130.050 144.600 ;
        RECT 88.950 142.950 91.050 143.400 ;
        RECT 127.950 142.950 130.050 143.400 ;
        RECT 244.950 144.600 247.050 145.050 ;
        RECT 256.950 144.600 259.050 145.050 ;
        RECT 295.950 144.600 298.050 145.050 ;
        RECT 244.950 143.400 298.050 144.600 ;
        RECT 244.950 142.950 247.050 143.400 ;
        RECT 256.950 142.950 259.050 143.400 ;
        RECT 295.950 142.950 298.050 143.400 ;
        RECT 70.950 141.600 73.050 142.200 ;
        RECT 398.400 142.050 399.600 146.400 ;
        RECT 445.950 146.400 454.050 147.600 ;
        RECT 445.950 145.950 448.050 146.400 ;
        RECT 451.950 145.950 454.050 146.400 ;
        RECT 610.950 147.600 613.050 148.050 ;
        RECT 643.950 147.600 646.050 148.050 ;
        RECT 610.950 146.400 646.050 147.600 ;
        RECT 610.950 145.950 613.050 146.400 ;
        RECT 643.950 145.950 646.050 146.400 ;
        RECT 790.950 147.600 793.050 148.050 ;
        RECT 796.950 147.600 799.050 148.050 ;
        RECT 790.950 146.400 799.050 147.600 ;
        RECT 790.950 145.950 793.050 146.400 ;
        RECT 796.950 145.950 799.050 146.400 ;
        RECT 526.950 144.600 529.050 145.050 ;
        RECT 619.950 144.600 622.050 145.050 ;
        RECT 526.950 143.400 622.050 144.600 ;
        RECT 526.950 142.950 529.050 143.400 ;
        RECT 619.950 142.950 622.050 143.400 ;
        RECT 703.950 144.600 706.050 145.050 ;
        RECT 712.950 144.600 715.050 145.050 ;
        RECT 703.950 143.400 715.050 144.600 ;
        RECT 703.950 142.950 706.050 143.400 ;
        RECT 712.950 142.950 715.050 143.400 ;
        RECT 718.950 144.600 721.050 145.050 ;
        RECT 727.950 144.600 730.050 145.050 ;
        RECT 718.950 143.400 730.050 144.600 ;
        RECT 718.950 142.950 721.050 143.400 ;
        RECT 727.950 142.950 730.050 143.400 ;
        RECT 742.950 144.600 745.050 145.050 ;
        RECT 784.950 144.600 787.050 145.050 ;
        RECT 742.950 143.400 787.050 144.600 ;
        RECT 742.950 142.950 745.050 143.400 ;
        RECT 784.950 142.950 787.050 143.400 ;
        RECT 85.950 141.600 88.050 142.050 ;
        RECT 70.950 140.400 88.050 141.600 ;
        RECT 70.950 140.100 73.050 140.400 ;
        RECT 85.950 139.950 88.050 140.400 ;
        RECT 151.950 141.600 154.050 142.050 ;
        RECT 160.950 141.600 163.050 142.050 ;
        RECT 175.950 141.600 178.050 142.050 ;
        RECT 190.950 141.600 193.050 142.050 ;
        RECT 151.950 140.400 193.050 141.600 ;
        RECT 151.950 139.950 154.050 140.400 ;
        RECT 160.950 139.950 163.050 140.400 ;
        RECT 175.950 139.950 178.050 140.400 ;
        RECT 190.950 139.950 193.050 140.400 ;
        RECT 211.950 141.600 214.050 142.050 ;
        RECT 247.950 141.600 250.050 142.050 ;
        RECT 298.950 141.600 301.050 142.050 ;
        RECT 211.950 140.400 301.050 141.600 ;
        RECT 211.950 139.950 214.050 140.400 ;
        RECT 247.950 139.950 250.050 140.400 ;
        RECT 298.950 139.950 301.050 140.400 ;
        RECT 397.950 139.950 400.050 142.050 ;
        RECT 52.950 138.600 58.050 139.050 ;
        RECT 67.950 138.600 70.050 138.900 ;
        RECT 52.950 137.400 70.050 138.600 ;
        RECT 52.950 136.950 58.050 137.400 ;
        RECT 67.950 136.800 70.050 137.400 ;
        RECT 220.950 138.600 223.050 139.050 ;
        RECT 232.950 138.600 235.050 139.050 ;
        RECT 220.950 137.400 235.050 138.600 ;
        RECT 220.950 136.950 223.050 137.400 ;
        RECT 232.950 136.950 235.050 137.400 ;
        RECT 262.950 138.600 265.050 139.050 ;
        RECT 286.950 138.600 289.050 139.050 ;
        RECT 361.950 138.600 364.050 139.050 ;
        RECT 367.950 138.600 370.050 139.200 ;
        RECT 262.950 138.000 294.600 138.600 ;
        RECT 262.950 137.400 295.050 138.000 ;
        RECT 262.950 136.950 265.050 137.400 ;
        RECT 286.950 136.950 289.050 137.400 ;
        RECT 16.950 135.600 19.050 136.050 ;
        RECT 196.950 135.600 199.050 136.050 ;
        RECT 238.950 135.600 241.050 136.050 ;
        RECT 16.950 134.400 51.600 135.600 ;
        RECT 16.950 133.950 19.050 134.400 ;
        RECT 50.400 132.600 51.600 134.400 ;
        RECT 196.950 134.400 241.050 135.600 ;
        RECT 196.950 133.950 199.050 134.400 ;
        RECT 238.950 133.950 241.050 134.400 ;
        RECT 292.950 133.950 295.050 137.400 ;
        RECT 361.950 137.400 370.050 138.600 ;
        RECT 361.950 136.950 364.050 137.400 ;
        RECT 367.950 137.100 370.050 137.400 ;
        RECT 379.950 136.950 385.050 139.050 ;
        RECT 442.950 138.600 445.050 142.050 ;
        RECT 490.950 141.600 493.050 142.050 ;
        RECT 490.950 141.000 498.600 141.600 ;
        RECT 490.950 140.400 499.050 141.000 ;
        RECT 490.950 139.950 493.050 140.400 ;
        RECT 454.950 138.600 457.050 139.050 ;
        RECT 442.950 138.000 457.050 138.600 ;
        RECT 443.400 137.400 457.050 138.000 ;
        RECT 454.950 136.950 457.050 137.400 ;
        RECT 496.950 136.950 499.050 140.400 ;
        RECT 511.950 138.600 514.050 142.050 ;
        RECT 544.950 141.600 547.050 142.050 ;
        RECT 577.950 141.600 580.050 142.050 ;
        RECT 589.950 141.600 592.050 142.050 ;
        RECT 544.950 140.400 592.050 141.600 ;
        RECT 544.950 139.950 547.050 140.400 ;
        RECT 577.950 139.950 580.050 140.400 ;
        RECT 589.950 139.950 592.050 140.400 ;
        RECT 634.950 139.950 640.050 142.050 ;
        RECT 649.950 139.950 655.050 142.050 ;
        RECT 526.950 138.600 529.050 139.050 ;
        RECT 511.950 138.000 529.050 138.600 ;
        RECT 512.400 137.400 529.050 138.000 ;
        RECT 526.950 136.950 529.050 137.400 ;
        RECT 595.950 138.600 598.050 139.050 ;
        RECT 613.950 138.600 616.050 139.050 ;
        RECT 595.950 137.400 616.050 138.600 ;
        RECT 673.950 138.600 676.050 142.050 ;
        RECT 772.950 141.600 775.050 142.050 ;
        RECT 790.950 141.600 793.050 142.050 ;
        RECT 772.950 140.400 793.050 141.600 ;
        RECT 772.950 139.950 775.050 140.400 ;
        RECT 790.950 139.950 793.050 140.400 ;
        RECT 799.950 141.600 802.050 142.050 ;
        RECT 811.950 141.600 814.050 142.050 ;
        RECT 799.950 140.400 814.050 141.600 ;
        RECT 799.950 139.950 802.050 140.400 ;
        RECT 811.950 139.950 814.050 140.400 ;
        RECT 691.950 138.600 694.050 139.050 ;
        RECT 673.950 138.000 694.050 138.600 ;
        RECT 674.400 137.400 694.050 138.000 ;
        RECT 595.950 136.950 598.050 137.400 ;
        RECT 613.950 136.950 616.050 137.400 ;
        RECT 691.950 136.950 694.050 137.400 ;
        RECT 706.950 136.950 712.050 139.050 ;
        RECT 724.950 138.600 727.050 139.050 ;
        RECT 745.950 138.600 748.050 139.050 ;
        RECT 724.950 137.400 748.050 138.600 ;
        RECT 724.950 136.950 727.050 137.400 ;
        RECT 745.950 136.950 748.050 137.400 ;
        RECT 322.950 135.600 325.050 136.050 ;
        RECT 331.950 135.600 334.050 136.050 ;
        RECT 322.950 134.400 334.050 135.600 ;
        RECT 322.950 133.950 325.050 134.400 ;
        RECT 331.950 133.950 334.050 134.400 ;
        RECT 367.950 135.600 370.050 135.900 ;
        RECT 388.950 135.600 391.050 136.050 ;
        RECT 367.950 134.400 391.050 135.600 ;
        RECT 367.950 133.800 370.050 134.400 ;
        RECT 388.950 133.950 391.050 134.400 ;
        RECT 409.950 135.600 412.050 135.900 ;
        RECT 451.950 135.600 454.050 136.050 ;
        RECT 409.950 134.400 454.050 135.600 ;
        RECT 409.950 133.800 412.050 134.400 ;
        RECT 451.950 133.950 454.050 134.400 ;
        RECT 493.950 135.600 496.050 136.050 ;
        RECT 505.950 135.600 508.050 136.050 ;
        RECT 556.950 135.600 559.050 136.050 ;
        RECT 493.950 134.400 559.050 135.600 ;
        RECT 493.950 133.950 496.050 134.400 ;
        RECT 505.950 133.950 508.050 134.400 ;
        RECT 556.950 133.950 559.050 134.400 ;
        RECT 766.950 135.600 769.050 136.200 ;
        RECT 778.950 135.600 781.050 136.050 ;
        RECT 766.950 134.400 781.050 135.600 ;
        RECT 766.950 134.100 769.050 134.400 ;
        RECT 778.950 133.950 781.050 134.400 ;
        RECT 433.950 133.050 436.050 133.200 ;
        RECT 91.950 132.600 94.050 133.050 ;
        RECT 103.950 132.600 106.050 133.050 ;
        RECT 50.400 131.400 66.600 132.600 ;
        RECT 65.400 129.600 66.600 131.400 ;
        RECT 91.950 131.400 106.050 132.600 ;
        RECT 91.950 130.950 94.050 131.400 ;
        RECT 103.950 130.950 106.050 131.400 ;
        RECT 115.950 132.600 118.050 133.050 ;
        RECT 157.950 132.600 160.050 133.050 ;
        RECT 115.950 131.400 160.050 132.600 ;
        RECT 115.950 130.950 118.050 131.400 ;
        RECT 157.950 130.950 160.050 131.400 ;
        RECT 433.950 131.100 439.050 133.050 ;
        RECT 447.000 132.600 451.050 133.050 ;
        RECT 481.950 132.600 484.050 133.050 ;
        RECT 446.400 131.400 484.050 132.600 ;
        RECT 435.000 130.950 439.050 131.100 ;
        RECT 447.000 130.950 451.050 131.400 ;
        RECT 481.950 130.950 484.050 131.400 ;
        RECT 595.950 132.600 598.050 133.050 ;
        RECT 610.950 132.600 613.050 133.050 ;
        RECT 595.950 131.400 613.050 132.600 ;
        RECT 595.950 130.950 598.050 131.400 ;
        RECT 610.950 130.950 613.050 131.400 ;
        RECT 652.950 132.600 655.050 133.050 ;
        RECT 688.950 132.600 691.050 133.050 ;
        RECT 652.950 131.400 691.050 132.600 ;
        RECT 652.950 130.950 655.050 131.400 ;
        RECT 688.950 130.950 691.050 131.400 ;
        RECT 724.950 132.600 727.050 133.050 ;
        RECT 733.950 132.600 736.050 133.050 ;
        RECT 724.950 131.400 736.050 132.600 ;
        RECT 724.950 130.950 727.050 131.400 ;
        RECT 733.950 130.950 736.050 131.400 ;
        RECT 748.950 132.600 751.050 133.050 ;
        RECT 790.950 132.600 793.050 133.050 ;
        RECT 748.950 131.400 793.050 132.600 ;
        RECT 748.950 130.950 751.050 131.400 ;
        RECT 790.950 130.950 793.050 131.400 ;
        RECT 796.950 132.600 799.050 133.050 ;
        RECT 817.950 132.600 820.050 133.050 ;
        RECT 796.950 131.400 820.050 132.600 ;
        RECT 796.950 130.950 799.050 131.400 ;
        RECT 817.950 130.950 820.050 131.400 ;
        RECT 73.950 129.600 76.050 130.050 ;
        RECT 65.400 128.400 76.050 129.600 ;
        RECT 73.950 127.950 76.050 128.400 ;
        RECT 385.950 129.600 388.050 130.050 ;
        RECT 412.950 129.600 415.050 130.050 ;
        RECT 385.950 128.400 415.050 129.600 ;
        RECT 385.950 127.950 388.050 128.400 ;
        RECT 412.950 127.950 415.050 128.400 ;
        RECT 493.950 129.600 496.050 130.050 ;
        RECT 529.950 129.600 532.050 130.050 ;
        RECT 493.950 128.400 532.050 129.600 ;
        RECT 493.950 127.950 496.050 128.400 ;
        RECT 529.950 127.950 532.050 128.400 ;
        RECT 691.950 129.600 694.050 130.050 ;
        RECT 706.950 129.600 709.050 130.050 ;
        RECT 691.950 128.400 709.050 129.600 ;
        RECT 691.950 127.950 694.050 128.400 ;
        RECT 706.950 127.950 709.050 128.400 ;
        RECT 751.950 129.600 754.050 130.050 ;
        RECT 787.950 129.600 790.050 130.050 ;
        RECT 751.950 128.400 790.050 129.600 ;
        RECT 751.950 127.950 754.050 128.400 ;
        RECT 787.950 127.950 790.050 128.400 ;
        RECT 538.950 126.600 541.050 127.050 ;
        RECT 652.950 126.600 655.050 127.050 ;
        RECT 538.950 125.400 655.050 126.600 ;
        RECT 538.950 124.950 541.050 125.400 ;
        RECT 652.950 124.950 655.050 125.400 ;
        RECT 16.950 123.600 19.050 124.050 ;
        RECT 34.950 123.600 37.050 124.050 ;
        RECT 55.950 123.600 58.050 124.050 ;
        RECT 16.950 122.400 58.050 123.600 ;
        RECT 16.950 121.950 19.050 122.400 ;
        RECT 34.950 121.950 37.050 122.400 ;
        RECT 55.950 121.950 58.050 122.400 ;
        RECT 151.950 123.600 154.050 124.050 ;
        RECT 325.950 123.600 328.050 124.050 ;
        RECT 337.950 123.600 340.050 124.050 ;
        RECT 151.950 122.400 340.050 123.600 ;
        RECT 151.950 121.950 154.050 122.400 ;
        RECT 325.950 121.950 328.050 122.400 ;
        RECT 337.950 121.950 340.050 122.400 ;
        RECT 391.950 123.600 394.050 124.050 ;
        RECT 415.950 123.600 418.050 124.050 ;
        RECT 391.950 122.400 418.050 123.600 ;
        RECT 391.950 121.950 394.050 122.400 ;
        RECT 415.950 121.950 418.050 122.400 ;
        RECT 664.950 123.600 667.050 124.050 ;
        RECT 700.950 123.600 703.050 124.050 ;
        RECT 664.950 122.400 703.050 123.600 ;
        RECT 664.950 121.950 667.050 122.400 ;
        RECT 700.950 121.950 703.050 122.400 ;
        RECT 424.950 120.600 427.050 121.050 ;
        RECT 454.950 120.600 457.050 121.050 ;
        RECT 424.950 119.400 457.050 120.600 ;
        RECT 424.950 118.950 427.050 119.400 ;
        RECT 454.950 118.950 457.050 119.400 ;
        RECT 460.950 120.600 463.050 121.050 ;
        RECT 508.950 120.600 511.050 121.050 ;
        RECT 529.950 120.600 532.050 121.050 ;
        RECT 460.950 119.400 532.050 120.600 ;
        RECT 460.950 118.950 463.050 119.400 ;
        RECT 508.950 118.950 511.050 119.400 ;
        RECT 529.950 118.950 532.050 119.400 ;
        RECT 544.950 120.600 547.050 121.050 ;
        RECT 550.950 120.600 553.050 121.050 ;
        RECT 544.950 119.400 553.050 120.600 ;
        RECT 544.950 118.950 547.050 119.400 ;
        RECT 550.950 118.950 553.050 119.400 ;
        RECT 580.950 120.600 583.050 121.050 ;
        RECT 595.950 120.600 598.050 121.050 ;
        RECT 580.950 119.400 598.050 120.600 ;
        RECT 580.950 118.950 583.050 119.400 ;
        RECT 595.950 118.950 598.050 119.400 ;
        RECT 619.950 120.600 622.050 121.050 ;
        RECT 739.950 120.600 742.050 121.050 ;
        RECT 619.950 119.400 742.050 120.600 ;
        RECT 619.950 118.950 622.050 119.400 ;
        RECT 739.950 118.950 742.050 119.400 ;
        RECT 775.950 120.600 778.050 121.050 ;
        RECT 808.950 120.600 811.050 121.050 ;
        RECT 775.950 119.400 811.050 120.600 ;
        RECT 775.950 118.950 778.050 119.400 ;
        RECT 808.950 118.950 811.050 119.400 ;
        RECT 46.950 117.600 49.050 118.050 ;
        RECT 35.400 116.400 49.050 117.600 ;
        RECT 13.950 114.600 16.050 115.050 ;
        RECT 35.400 114.600 36.600 116.400 ;
        RECT 46.950 115.950 49.050 116.400 ;
        RECT 397.950 117.600 400.050 118.050 ;
        RECT 406.950 117.600 409.050 118.050 ;
        RECT 397.950 116.400 409.050 117.600 ;
        RECT 397.950 115.950 400.050 116.400 ;
        RECT 406.950 115.950 409.050 116.400 ;
        RECT 667.950 117.600 670.050 118.050 ;
        RECT 679.950 117.600 682.050 118.050 ;
        RECT 667.950 116.400 682.050 117.600 ;
        RECT 667.950 115.950 670.050 116.400 ;
        RECT 679.950 115.950 682.050 116.400 ;
        RECT 724.950 117.600 727.050 118.050 ;
        RECT 766.950 117.600 769.050 118.050 ;
        RECT 724.950 116.400 769.050 117.600 ;
        RECT 724.950 115.950 727.050 116.400 ;
        RECT 766.950 115.950 769.050 116.400 ;
        RECT 13.950 113.400 36.600 114.600 ;
        RECT 286.950 114.600 289.050 115.050 ;
        RECT 322.950 114.600 325.050 115.050 ;
        RECT 286.950 113.400 325.050 114.600 ;
        RECT 13.950 112.950 16.050 113.400 ;
        RECT 286.950 112.950 289.050 113.400 ;
        RECT 322.950 112.950 325.050 113.400 ;
        RECT 31.950 111.600 34.050 112.050 ;
        RECT 37.950 111.600 40.050 112.200 ;
        RECT 31.950 110.400 40.050 111.600 ;
        RECT 31.950 109.950 34.050 110.400 ;
        RECT 37.950 110.100 40.050 110.400 ;
        RECT 172.950 111.600 175.050 112.050 ;
        RECT 337.950 111.600 340.050 112.050 ;
        RECT 172.950 110.400 340.050 111.600 ;
        RECT 172.950 109.950 175.050 110.400 ;
        RECT 337.950 109.950 340.050 110.400 ;
        RECT 418.950 111.600 421.050 112.050 ;
        RECT 472.950 111.600 475.050 112.050 ;
        RECT 418.950 110.400 475.050 111.600 ;
        RECT 418.950 109.950 421.050 110.400 ;
        RECT 472.950 109.950 475.050 110.400 ;
        RECT 490.950 111.600 493.050 112.050 ;
        RECT 514.950 111.600 517.050 112.050 ;
        RECT 490.950 110.400 517.050 111.600 ;
        RECT 490.950 109.950 493.050 110.400 ;
        RECT 514.950 109.950 517.050 110.400 ;
        RECT 556.950 111.600 559.050 112.050 ;
        RECT 583.950 111.600 586.050 112.050 ;
        RECT 556.950 110.400 586.050 111.600 ;
        RECT 556.950 109.950 559.050 110.400 ;
        RECT 583.950 109.950 586.050 110.400 ;
        RECT 607.950 111.600 610.050 112.050 ;
        RECT 664.950 111.600 667.050 112.050 ;
        RECT 607.950 110.400 667.050 111.600 ;
        RECT 607.950 109.950 610.050 110.400 ;
        RECT 664.950 109.950 667.050 110.400 ;
        RECT 715.950 111.600 718.050 112.050 ;
        RECT 745.950 111.600 748.050 112.050 ;
        RECT 715.950 110.400 748.050 111.600 ;
        RECT 715.950 109.950 718.050 110.400 ;
        RECT 745.950 109.950 748.050 110.400 ;
        RECT 214.950 108.600 217.050 109.050 ;
        RECT 232.950 108.600 235.050 109.050 ;
        RECT 214.950 107.400 235.050 108.600 ;
        RECT 214.950 106.950 217.050 107.400 ;
        RECT 232.950 106.950 235.050 107.400 ;
        RECT 370.950 108.600 373.050 109.050 ;
        RECT 412.950 108.600 415.050 109.050 ;
        RECT 370.950 107.400 415.050 108.600 ;
        RECT 370.950 106.950 373.050 107.400 ;
        RECT 412.950 106.950 415.050 107.400 ;
        RECT 511.950 108.600 514.050 109.050 ;
        RECT 559.950 108.600 562.050 109.050 ;
        RECT 511.950 107.400 562.050 108.600 ;
        RECT 511.950 106.950 514.050 107.400 ;
        RECT 559.950 106.950 562.050 107.400 ;
        RECT 37.950 105.600 40.050 106.050 ;
        RECT 46.950 105.600 49.050 106.050 ;
        RECT 61.950 105.600 64.050 106.050 ;
        RECT 79.950 105.600 82.050 106.050 ;
        RECT 37.950 104.400 82.050 105.600 ;
        RECT 37.950 103.950 40.050 104.400 ;
        RECT 46.950 103.950 49.050 104.400 ;
        RECT 61.950 103.950 64.050 104.400 ;
        RECT 79.950 103.950 82.050 104.400 ;
        RECT 130.950 105.600 133.050 106.050 ;
        RECT 241.950 105.600 244.050 106.050 ;
        RECT 262.950 105.600 265.050 106.050 ;
        RECT 130.950 105.000 144.600 105.600 ;
        RECT 130.950 104.400 145.050 105.000 ;
        RECT 130.950 103.950 133.050 104.400 ;
        RECT 106.950 102.600 109.050 103.050 ;
        RECT 136.950 102.600 139.050 103.050 ;
        RECT 106.950 101.400 139.050 102.600 ;
        RECT 106.950 100.950 109.050 101.400 ;
        RECT 136.950 100.950 139.050 101.400 ;
        RECT 142.950 100.950 145.050 104.400 ;
        RECT 241.950 104.400 265.050 105.600 ;
        RECT 241.950 103.950 244.050 104.400 ;
        RECT 262.950 103.950 265.050 104.400 ;
        RECT 157.950 102.600 160.050 103.050 ;
        RECT 166.950 102.600 169.050 103.050 ;
        RECT 157.950 101.400 169.050 102.600 ;
        RECT 295.950 102.600 298.050 106.050 ;
        RECT 313.950 103.950 319.050 106.050 ;
        RECT 340.950 105.600 343.050 106.050 ;
        RECT 355.950 105.600 358.050 106.050 ;
        RECT 367.950 105.600 370.050 106.050 ;
        RECT 340.950 104.400 370.050 105.600 ;
        RECT 340.950 103.950 343.050 104.400 ;
        RECT 355.950 103.950 358.050 104.400 ;
        RECT 367.950 103.950 370.050 104.400 ;
        RECT 307.950 102.600 310.050 103.050 ;
        RECT 295.950 102.000 310.050 102.600 ;
        RECT 296.400 101.400 310.050 102.000 ;
        RECT 157.950 100.950 160.050 101.400 ;
        RECT 166.950 100.950 169.050 101.400 ;
        RECT 307.950 100.950 310.050 101.400 ;
        RECT 31.950 99.600 34.050 100.050 ;
        RECT 43.950 99.600 46.050 100.050 ;
        RECT 31.950 98.400 46.050 99.600 ;
        RECT 31.950 97.950 34.050 98.400 ;
        RECT 43.950 97.950 46.050 98.400 ;
        RECT 55.950 99.600 58.050 100.050 ;
        RECT 64.950 99.600 67.050 100.050 ;
        RECT 85.950 99.600 88.050 100.050 ;
        RECT 55.950 98.400 88.050 99.600 ;
        RECT 55.950 97.950 58.050 98.400 ;
        RECT 64.950 97.950 67.050 98.400 ;
        RECT 85.950 97.950 88.050 98.400 ;
        RECT 115.950 99.600 118.050 100.050 ;
        RECT 121.950 99.600 124.050 100.050 ;
        RECT 115.950 98.400 124.050 99.600 ;
        RECT 115.950 97.950 118.050 98.400 ;
        RECT 121.950 97.950 124.050 98.400 ;
        RECT 106.950 96.600 109.050 97.050 ;
        RECT 142.950 96.600 145.050 97.050 ;
        RECT 106.950 95.400 145.050 96.600 ;
        RECT 106.950 94.950 109.050 95.400 ;
        RECT 142.950 94.950 145.050 95.400 ;
        RECT 160.950 96.600 163.050 97.050 ;
        RECT 172.950 96.600 175.050 99.900 ;
        RECT 226.950 99.600 229.050 100.050 ;
        RECT 232.950 99.600 235.050 100.050 ;
        RECT 226.950 98.400 235.050 99.600 ;
        RECT 226.950 97.950 229.050 98.400 ;
        RECT 232.950 97.950 235.050 98.400 ;
        RECT 244.950 97.950 250.050 100.050 ;
        RECT 298.950 99.600 301.050 100.050 ;
        RECT 328.950 99.600 331.050 103.050 ;
        RECT 298.950 99.000 331.050 99.600 ;
        RECT 337.950 99.600 340.050 100.050 ;
        RECT 358.950 99.600 361.050 100.050 ;
        RECT 298.950 98.400 330.600 99.000 ;
        RECT 337.950 98.400 361.050 99.600 ;
        RECT 298.950 97.950 301.050 98.400 ;
        RECT 337.950 97.950 340.050 98.400 ;
        RECT 358.950 97.950 361.050 98.400 ;
        RECT 364.950 99.600 367.050 100.050 ;
        RECT 385.950 99.600 388.050 103.050 ;
        RECT 442.950 102.600 445.050 106.050 ;
        RECT 526.950 105.600 529.050 106.050 ;
        RECT 518.400 104.400 529.050 105.600 ;
        RECT 565.950 105.600 568.050 109.050 ;
        RECT 586.950 108.600 589.050 109.050 ;
        RECT 601.950 108.600 604.050 109.050 ;
        RECT 586.950 107.400 604.050 108.600 ;
        RECT 586.950 106.950 589.050 107.400 ;
        RECT 601.950 106.950 604.050 107.400 ;
        RECT 736.950 108.600 739.050 109.050 ;
        RECT 748.950 108.600 751.050 109.050 ;
        RECT 736.950 107.400 751.050 108.600 ;
        RECT 736.950 106.950 739.050 107.400 ;
        RECT 748.950 106.950 751.050 107.400 ;
        RECT 781.950 108.600 784.050 109.050 ;
        RECT 808.950 108.600 811.050 109.050 ;
        RECT 781.950 107.400 811.050 108.600 ;
        RECT 781.950 106.950 784.050 107.400 ;
        RECT 808.950 106.950 811.050 107.400 ;
        RECT 583.950 105.600 586.050 106.050 ;
        RECT 667.950 105.600 670.050 106.050 ;
        RECT 565.950 105.000 586.050 105.600 ;
        RECT 635.400 105.000 670.050 105.600 ;
        RECT 566.400 104.400 586.050 105.000 ;
        RECT 518.400 103.050 519.600 104.400 ;
        RECT 526.950 103.950 529.050 104.400 ;
        RECT 583.950 103.950 586.050 104.400 ;
        RECT 634.950 104.400 670.050 105.000 ;
        RECT 460.950 102.600 463.050 103.050 ;
        RECT 517.950 102.600 520.050 103.050 ;
        RECT 442.950 102.000 463.050 102.600 ;
        RECT 443.400 101.400 463.050 102.000 ;
        RECT 460.950 100.950 463.050 101.400 ;
        RECT 506.400 101.400 520.050 102.600 ;
        RECT 506.400 100.050 507.600 101.400 ;
        RECT 517.950 100.950 520.050 101.400 ;
        RECT 559.950 102.600 562.050 103.050 ;
        RECT 598.950 102.600 601.050 103.050 ;
        RECT 559.950 101.400 601.050 102.600 ;
        RECT 559.950 100.950 562.050 101.400 ;
        RECT 598.950 100.950 601.050 101.400 ;
        RECT 634.950 100.800 637.050 104.400 ;
        RECT 667.950 103.950 670.050 104.400 ;
        RECT 679.950 105.600 682.050 106.050 ;
        RECT 775.950 105.600 778.050 106.050 ;
        RECT 679.950 104.400 778.050 105.600 ;
        RECT 679.950 103.950 682.050 104.400 ;
        RECT 775.950 103.950 778.050 104.400 ;
        RECT 685.950 102.600 688.050 103.050 ;
        RECT 709.950 102.600 712.050 103.050 ;
        RECT 685.950 101.400 712.050 102.600 ;
        RECT 685.950 100.950 688.050 101.400 ;
        RECT 709.950 100.950 712.050 101.400 ;
        RECT 715.950 102.600 718.050 103.200 ;
        RECT 751.950 102.600 756.000 103.050 ;
        RECT 793.950 102.600 796.050 103.050 ;
        RECT 805.950 102.600 808.050 103.200 ;
        RECT 715.950 101.400 756.600 102.600 ;
        RECT 793.950 101.400 808.050 102.600 ;
        RECT 715.950 101.100 718.050 101.400 ;
        RECT 751.950 100.950 756.000 101.400 ;
        RECT 793.950 100.950 796.050 101.400 ;
        RECT 805.950 101.100 808.050 101.400 ;
        RECT 610.950 100.050 613.050 100.200 ;
        RECT 364.950 99.000 388.050 99.600 ;
        RECT 403.950 99.600 406.050 100.050 ;
        RECT 412.950 99.600 415.050 99.900 ;
        RECT 424.950 99.600 427.050 100.050 ;
        RECT 364.950 98.400 387.600 99.000 ;
        RECT 403.950 98.400 427.050 99.600 ;
        RECT 364.950 97.950 367.050 98.400 ;
        RECT 403.950 97.950 406.050 98.400 ;
        RECT 412.950 97.800 415.050 98.400 ;
        RECT 424.950 97.950 427.050 98.400 ;
        RECT 478.950 99.600 481.050 100.050 ;
        RECT 496.950 99.600 499.050 100.050 ;
        RECT 478.950 98.400 499.050 99.600 ;
        RECT 478.950 97.950 481.050 98.400 ;
        RECT 496.950 97.950 499.050 98.400 ;
        RECT 502.950 98.400 507.600 100.050 ;
        RECT 502.950 97.950 507.000 98.400 ;
        RECT 607.950 98.100 613.050 100.050 ;
        RECT 715.950 99.600 718.050 99.900 ;
        RECT 721.950 99.600 724.050 100.050 ;
        RECT 715.950 98.400 724.050 99.600 ;
        RECT 607.950 97.950 612.000 98.100 ;
        RECT 715.950 97.800 718.050 98.400 ;
        RECT 721.950 97.950 724.050 98.400 ;
        RECT 160.950 96.000 175.050 96.600 ;
        RECT 289.950 96.600 292.050 97.050 ;
        RECT 301.950 96.600 304.050 97.050 ;
        RECT 160.950 95.400 174.600 96.000 ;
        RECT 289.950 95.400 304.050 96.600 ;
        RECT 160.950 94.950 163.050 95.400 ;
        RECT 289.950 94.950 292.050 95.400 ;
        RECT 301.950 94.950 304.050 95.400 ;
        RECT 481.950 96.600 484.050 97.050 ;
        RECT 493.950 96.600 496.050 97.050 ;
        RECT 481.950 95.400 496.050 96.600 ;
        RECT 481.950 94.950 484.050 95.400 ;
        RECT 493.950 94.950 496.050 95.400 ;
        RECT 565.950 96.600 568.050 97.050 ;
        RECT 577.950 96.600 580.050 97.050 ;
        RECT 565.950 95.400 580.050 96.600 ;
        RECT 565.950 94.950 568.050 95.400 ;
        RECT 577.950 94.950 580.050 95.400 ;
        RECT 598.950 96.600 601.050 97.050 ;
        RECT 619.950 96.600 622.050 97.050 ;
        RECT 598.950 95.400 622.050 96.600 ;
        RECT 598.950 94.950 601.050 95.400 ;
        RECT 619.950 94.950 622.050 95.400 ;
        RECT 706.950 96.600 709.050 97.050 ;
        RECT 733.950 96.600 736.050 97.050 ;
        RECT 706.950 95.400 736.050 96.600 ;
        RECT 706.950 94.950 709.050 95.400 ;
        RECT 733.950 94.950 736.050 95.400 ;
        RECT 76.950 93.600 79.050 94.050 ;
        RECT 100.950 93.600 103.050 94.050 ;
        RECT 76.950 92.400 103.050 93.600 ;
        RECT 76.950 91.950 79.050 92.400 ;
        RECT 100.950 91.950 103.050 92.400 ;
        RECT 130.950 93.600 133.050 94.050 ;
        RECT 136.950 93.600 139.050 94.050 ;
        RECT 130.950 92.400 139.050 93.600 ;
        RECT 130.950 91.950 133.050 92.400 ;
        RECT 136.950 91.950 139.050 92.400 ;
        RECT 556.950 93.600 559.050 94.050 ;
        RECT 583.950 93.600 586.050 94.050 ;
        RECT 556.950 92.400 586.050 93.600 ;
        RECT 556.950 91.950 559.050 92.400 ;
        RECT 583.950 91.950 586.050 92.400 ;
        RECT 241.950 90.600 244.050 91.050 ;
        RECT 319.950 90.600 322.050 91.050 ;
        RECT 241.950 89.400 322.050 90.600 ;
        RECT 241.950 88.950 244.050 89.400 ;
        RECT 319.950 88.950 322.050 89.400 ;
        RECT 484.950 90.600 487.050 91.050 ;
        RECT 499.950 90.600 502.050 91.050 ;
        RECT 505.800 90.600 507.900 91.050 ;
        RECT 484.950 89.400 507.900 90.600 ;
        RECT 484.950 88.950 487.050 89.400 ;
        RECT 499.950 88.950 502.050 89.400 ;
        RECT 505.800 88.950 507.900 89.400 ;
        RECT 509.100 90.600 511.200 91.050 ;
        RECT 550.950 90.600 553.050 91.050 ;
        RECT 509.100 89.400 553.050 90.600 ;
        RECT 509.100 88.950 511.200 89.400 ;
        RECT 550.950 88.950 553.050 89.400 ;
        RECT 349.950 87.600 352.050 88.050 ;
        RECT 463.950 87.600 466.050 88.050 ;
        RECT 652.950 87.600 655.050 88.050 ;
        RECT 349.950 86.400 655.050 87.600 ;
        RECT 349.950 85.950 352.050 86.400 ;
        RECT 463.950 85.950 466.050 86.400 ;
        RECT 652.950 85.950 655.050 86.400 ;
        RECT 67.950 84.600 70.050 85.050 ;
        RECT 79.950 84.600 82.050 85.050 ;
        RECT 67.950 83.400 82.050 84.600 ;
        RECT 67.950 82.950 70.050 83.400 ;
        RECT 79.950 82.950 82.050 83.400 ;
        RECT 205.950 84.600 208.050 85.050 ;
        RECT 268.950 84.600 271.050 85.050 ;
        RECT 205.950 83.400 271.050 84.600 ;
        RECT 205.950 82.950 208.050 83.400 ;
        RECT 268.950 82.950 271.050 83.400 ;
        RECT 274.950 84.600 277.050 85.050 ;
        RECT 350.400 84.600 351.600 85.950 ;
        RECT 274.950 83.400 351.600 84.600 ;
        RECT 478.950 84.600 481.050 85.050 ;
        RECT 640.950 84.600 643.050 85.050 ;
        RECT 478.950 83.400 643.050 84.600 ;
        RECT 274.950 82.950 277.050 83.400 ;
        RECT 478.950 82.950 481.050 83.400 ;
        RECT 640.950 82.950 643.050 83.400 ;
        RECT 739.950 84.600 742.050 85.050 ;
        RECT 808.950 84.600 811.050 85.050 ;
        RECT 739.950 83.400 811.050 84.600 ;
        RECT 739.950 82.950 742.050 83.400 ;
        RECT 808.950 82.950 811.050 83.400 ;
        RECT 124.950 81.600 127.050 82.050 ;
        RECT 154.950 81.600 157.050 82.050 ;
        RECT 124.950 80.400 157.050 81.600 ;
        RECT 124.950 79.950 127.050 80.400 ;
        RECT 154.950 79.950 157.050 80.400 ;
        RECT 577.950 81.600 580.050 82.050 ;
        RECT 595.950 81.600 598.050 82.050 ;
        RECT 577.950 80.400 598.050 81.600 ;
        RECT 577.950 79.950 580.050 80.400 ;
        RECT 595.950 79.950 598.050 80.400 ;
        RECT 79.950 78.600 82.050 79.050 ;
        RECT 166.950 78.600 169.050 79.050 ;
        RECT 79.950 77.400 169.050 78.600 ;
        RECT 79.950 76.950 82.050 77.400 ;
        RECT 166.950 76.950 169.050 77.400 ;
        RECT 268.950 78.600 271.050 79.050 ;
        RECT 412.950 78.600 415.050 79.050 ;
        RECT 535.950 78.600 538.050 79.050 ;
        RECT 631.950 78.600 634.050 79.050 ;
        RECT 268.950 77.400 415.050 78.600 ;
        RECT 268.950 76.950 271.050 77.400 ;
        RECT 412.950 76.950 415.050 77.400 ;
        RECT 524.400 77.400 634.050 78.600 ;
        RECT 524.400 76.050 525.600 77.400 ;
        RECT 535.950 76.950 538.050 77.400 ;
        RECT 631.950 76.950 634.050 77.400 ;
        RECT 724.950 78.600 727.050 79.050 ;
        RECT 745.950 78.600 748.050 79.050 ;
        RECT 817.950 78.600 820.050 79.050 ;
        RECT 724.950 77.400 748.050 78.600 ;
        RECT 724.950 76.950 727.050 77.400 ;
        RECT 745.950 76.950 748.050 77.400 ;
        RECT 803.400 77.400 820.050 78.600 ;
        RECT 40.950 75.600 43.050 76.050 ;
        RECT 76.950 75.600 79.050 76.050 ;
        RECT 40.950 74.400 79.050 75.600 ;
        RECT 40.950 73.950 43.050 74.400 ;
        RECT 76.950 73.950 79.050 74.400 ;
        RECT 184.950 75.600 187.050 76.050 ;
        RECT 190.950 75.600 193.050 76.050 ;
        RECT 184.950 74.400 193.050 75.600 ;
        RECT 184.950 73.950 187.050 74.400 ;
        RECT 190.950 73.950 193.050 74.400 ;
        RECT 232.950 75.600 235.050 76.050 ;
        RECT 262.950 75.600 265.050 76.050 ;
        RECT 232.950 74.400 265.050 75.600 ;
        RECT 232.950 73.950 235.050 74.400 ;
        RECT 262.950 73.950 265.050 74.400 ;
        RECT 379.950 75.600 382.050 76.050 ;
        RECT 391.950 75.600 394.050 76.050 ;
        RECT 397.950 75.600 400.050 76.050 ;
        RECT 379.950 74.400 400.050 75.600 ;
        RECT 379.950 73.950 382.050 74.400 ;
        RECT 391.950 73.950 394.050 74.400 ;
        RECT 397.950 73.950 400.050 74.400 ;
        RECT 457.950 75.600 460.050 76.050 ;
        RECT 523.950 75.600 526.050 76.050 ;
        RECT 457.950 74.400 526.050 75.600 ;
        RECT 457.950 73.950 460.050 74.400 ;
        RECT 523.950 73.950 526.050 74.400 ;
        RECT 529.950 75.600 532.050 76.050 ;
        RECT 544.950 75.600 547.050 76.050 ;
        RECT 529.950 74.400 547.050 75.600 ;
        RECT 529.950 73.950 532.050 74.400 ;
        RECT 544.950 73.950 547.050 74.400 ;
        RECT 796.950 75.600 799.050 76.050 ;
        RECT 803.400 75.600 804.600 77.400 ;
        RECT 817.950 76.950 820.050 77.400 ;
        RECT 796.950 74.400 804.600 75.600 ;
        RECT 796.950 73.950 799.050 74.400 ;
        RECT 286.950 72.600 289.050 73.050 ;
        RECT 301.950 72.600 304.050 73.050 ;
        RECT 340.950 72.600 343.050 73.050 ;
        RECT 286.950 71.400 343.050 72.600 ;
        RECT 286.950 70.950 289.050 71.400 ;
        RECT 301.950 70.950 304.050 71.400 ;
        RECT 340.950 70.950 343.050 71.400 ;
        RECT 610.950 72.600 613.050 73.050 ;
        RECT 682.950 72.600 685.050 73.050 ;
        RECT 610.950 71.400 685.050 72.600 ;
        RECT 610.950 70.950 613.050 71.400 ;
        RECT 682.950 70.950 685.050 71.400 ;
        RECT 724.950 72.600 727.050 73.050 ;
        RECT 748.950 72.600 751.050 73.050 ;
        RECT 805.950 72.600 808.050 73.050 ;
        RECT 724.950 71.400 808.050 72.600 ;
        RECT 724.950 70.950 727.050 71.400 ;
        RECT 748.950 70.950 751.050 71.400 ;
        RECT 805.950 70.950 808.050 71.400 ;
        RECT 112.950 69.600 115.050 70.050 ;
        RECT 184.950 69.600 187.050 70.050 ;
        RECT 112.950 68.400 187.050 69.600 ;
        RECT 112.950 67.950 115.050 68.400 ;
        RECT 184.950 67.950 187.050 68.400 ;
        RECT 199.950 69.600 202.050 70.050 ;
        RECT 214.950 69.600 217.050 70.050 ;
        RECT 256.950 69.600 259.050 70.050 ;
        RECT 199.950 68.400 259.050 69.600 ;
        RECT 199.950 67.950 202.050 68.400 ;
        RECT 214.950 67.950 217.050 68.400 ;
        RECT 256.950 67.950 259.050 68.400 ;
        RECT 406.950 69.600 409.050 70.050 ;
        RECT 433.950 69.600 436.050 70.050 ;
        RECT 406.950 68.400 436.050 69.600 ;
        RECT 406.950 67.950 409.050 68.400 ;
        RECT 433.950 67.950 436.050 68.400 ;
        RECT 460.950 69.600 463.050 70.050 ;
        RECT 499.950 69.600 502.050 70.050 ;
        RECT 460.950 68.400 502.050 69.600 ;
        RECT 460.950 67.950 463.050 68.400 ;
        RECT 499.950 67.950 502.050 68.400 ;
        RECT 673.950 69.600 676.050 70.050 ;
        RECT 679.950 69.600 682.050 70.050 ;
        RECT 673.950 68.400 682.050 69.600 ;
        RECT 673.950 67.950 676.050 68.400 ;
        RECT 679.950 67.950 682.050 68.400 ;
        RECT 730.950 69.600 733.050 70.050 ;
        RECT 742.950 69.600 745.050 70.050 ;
        RECT 730.950 68.400 745.050 69.600 ;
        RECT 730.950 67.950 733.050 68.400 ;
        RECT 742.950 67.950 745.050 68.400 ;
        RECT 4.950 66.600 7.050 67.050 ;
        RECT 13.950 66.600 16.050 67.050 ;
        RECT 4.950 65.400 16.050 66.600 ;
        RECT 4.950 64.950 7.050 65.400 ;
        RECT 13.950 64.950 16.050 65.400 ;
        RECT 277.950 66.600 280.050 67.050 ;
        RECT 283.950 66.600 286.050 67.050 ;
        RECT 277.950 65.400 286.050 66.600 ;
        RECT 277.950 64.950 280.050 65.400 ;
        RECT 283.950 64.950 286.050 65.400 ;
        RECT 130.950 63.600 133.050 64.050 ;
        RECT 253.950 63.600 256.050 64.050 ;
        RECT 286.950 63.600 289.050 64.050 ;
        RECT 130.950 62.400 256.050 63.600 ;
        RECT 266.400 63.000 289.050 63.600 ;
        RECT 130.950 61.950 133.050 62.400 ;
        RECT 253.950 61.950 256.050 62.400 ;
        RECT 265.950 62.400 289.050 63.000 ;
        RECT 1.950 60.600 4.050 61.050 ;
        RECT 16.950 60.600 19.050 61.050 ;
        RECT 1.950 59.400 19.050 60.600 ;
        RECT 1.950 58.950 4.050 59.400 ;
        RECT 16.950 58.950 19.050 59.400 ;
        RECT 163.950 60.600 166.050 61.200 ;
        RECT 202.950 60.600 205.050 61.050 ;
        RECT 163.950 59.400 205.050 60.600 ;
        RECT 163.950 59.100 166.050 59.400 ;
        RECT 202.950 58.950 205.050 59.400 ;
        RECT 241.950 60.600 244.050 61.050 ;
        RECT 250.950 60.600 253.050 61.050 ;
        RECT 241.950 59.400 253.050 60.600 ;
        RECT 241.950 58.950 244.050 59.400 ;
        RECT 250.950 58.950 253.050 59.400 ;
        RECT 265.950 58.950 268.050 62.400 ;
        RECT 286.950 61.950 289.050 62.400 ;
        RECT 274.950 60.600 277.050 61.050 ;
        RECT 292.950 60.600 295.050 61.050 ;
        RECT 274.950 59.400 295.050 60.600 ;
        RECT 274.950 58.950 277.050 59.400 ;
        RECT 292.950 58.950 295.050 59.400 ;
        RECT 328.950 60.600 331.050 61.050 ;
        RECT 343.950 60.600 346.050 64.050 ;
        RECT 328.950 60.000 346.050 60.600 ;
        RECT 355.950 60.600 358.050 61.050 ;
        RECT 373.950 60.600 376.050 64.050 ;
        RECT 394.950 63.600 397.050 64.050 ;
        RECT 406.950 63.600 409.050 64.050 ;
        RECT 394.950 62.400 409.050 63.600 ;
        RECT 394.950 61.950 397.050 62.400 ;
        RECT 406.950 61.950 409.050 62.400 ;
        RECT 496.950 63.600 499.050 64.050 ;
        RECT 520.950 63.600 523.050 64.050 ;
        RECT 496.950 62.400 523.050 63.600 ;
        RECT 496.950 61.950 499.050 62.400 ;
        RECT 520.950 61.950 523.050 62.400 ;
        RECT 538.950 63.600 541.050 64.050 ;
        RECT 568.950 63.600 571.050 64.050 ;
        RECT 538.950 62.400 571.050 63.600 ;
        RECT 538.950 61.950 541.050 62.400 ;
        RECT 568.950 61.950 571.050 62.400 ;
        RECT 589.950 63.600 592.050 64.050 ;
        RECT 616.950 63.600 619.050 64.050 ;
        RECT 589.950 62.400 619.050 63.600 ;
        RECT 589.950 61.950 592.050 62.400 ;
        RECT 616.950 61.950 619.050 62.400 ;
        RECT 628.950 63.600 631.050 64.200 ;
        RECT 649.950 63.600 652.050 64.050 ;
        RECT 688.950 63.600 691.050 67.050 ;
        RECT 727.950 66.600 730.050 67.050 ;
        RECT 781.950 66.600 784.050 67.050 ;
        RECT 799.950 66.600 802.050 67.050 ;
        RECT 814.950 66.600 817.050 67.050 ;
        RECT 716.400 65.400 817.050 66.600 ;
        RECT 716.400 64.050 717.600 65.400 ;
        RECT 727.950 64.950 730.050 65.400 ;
        RECT 781.950 64.950 784.050 65.400 ;
        RECT 799.950 64.950 802.050 65.400 ;
        RECT 814.950 64.950 817.050 65.400 ;
        RECT 715.950 63.600 718.050 64.050 ;
        RECT 628.950 62.400 718.050 63.600 ;
        RECT 628.950 62.100 631.050 62.400 ;
        RECT 649.950 61.950 652.050 62.400 ;
        RECT 715.950 61.950 718.050 62.400 ;
        RECT 721.950 63.600 724.050 64.050 ;
        RECT 751.950 63.600 754.050 64.050 ;
        RECT 757.950 63.600 760.050 64.050 ;
        RECT 721.950 62.400 760.050 63.600 ;
        RECT 721.950 61.950 724.050 62.400 ;
        RECT 751.950 61.950 754.050 62.400 ;
        RECT 757.950 61.950 760.050 62.400 ;
        RECT 355.950 60.000 376.050 60.600 ;
        RECT 424.950 60.600 427.050 61.050 ;
        RECT 487.950 60.600 490.050 61.050 ;
        RECT 328.950 59.400 345.600 60.000 ;
        RECT 355.950 59.400 375.600 60.000 ;
        RECT 424.950 59.400 490.050 60.600 ;
        RECT 328.950 58.950 331.050 59.400 ;
        RECT 355.950 58.950 358.050 59.400 ;
        RECT 424.950 58.950 427.050 59.400 ;
        RECT 487.950 58.950 490.050 59.400 ;
        RECT 643.950 60.600 646.050 61.050 ;
        RECT 652.950 60.600 655.050 61.050 ;
        RECT 661.950 60.600 664.050 61.050 ;
        RECT 643.950 59.400 664.050 60.600 ;
        RECT 643.950 58.950 646.050 59.400 ;
        RECT 652.950 58.950 655.050 59.400 ;
        RECT 661.950 58.950 664.050 59.400 ;
        RECT 766.950 60.600 769.050 61.050 ;
        RECT 775.950 60.600 778.050 61.050 ;
        RECT 787.950 60.600 790.050 61.050 ;
        RECT 766.950 59.400 790.050 60.600 ;
        RECT 766.950 58.950 769.050 59.400 ;
        RECT 775.950 58.950 778.050 59.400 ;
        RECT 787.950 58.950 790.050 59.400 ;
        RECT 49.950 57.600 52.050 58.050 ;
        RECT 112.950 57.600 115.050 58.050 ;
        RECT 20.400 57.000 115.050 57.600 ;
        RECT 19.950 56.400 115.050 57.000 ;
        RECT 4.950 54.600 7.050 55.050 ;
        RECT 13.950 54.600 16.050 55.050 ;
        RECT 4.950 53.400 16.050 54.600 ;
        RECT 4.950 52.950 7.050 53.400 ;
        RECT 13.950 52.950 16.050 53.400 ;
        RECT 19.950 52.950 22.050 56.400 ;
        RECT 49.950 55.950 52.050 56.400 ;
        RECT 112.950 55.950 115.050 56.400 ;
        RECT 163.950 57.600 166.050 57.900 ;
        RECT 178.950 57.600 181.050 58.050 ;
        RECT 163.950 56.400 181.050 57.600 ;
        RECT 163.950 55.800 166.050 56.400 ;
        RECT 178.950 55.950 181.050 56.400 ;
        RECT 127.950 52.950 133.050 55.050 ;
        RECT 196.950 54.600 199.050 58.050 ;
        RECT 253.950 57.600 256.050 58.050 ;
        RECT 313.950 57.600 316.050 58.050 ;
        RECT 253.950 56.400 316.050 57.600 ;
        RECT 253.950 55.950 256.050 56.400 ;
        RECT 313.950 55.950 316.050 56.400 ;
        RECT 322.950 57.600 325.050 58.050 ;
        RECT 403.950 57.600 406.050 58.050 ;
        RECT 409.950 57.600 412.050 58.200 ;
        RECT 322.950 56.400 412.050 57.600 ;
        RECT 322.950 55.950 325.050 56.400 ;
        RECT 403.950 55.950 406.050 56.400 ;
        RECT 409.950 56.100 412.050 56.400 ;
        RECT 205.950 54.600 208.050 55.050 ;
        RECT 196.950 54.000 208.050 54.600 ;
        RECT 197.400 53.400 208.050 54.000 ;
        RECT 205.950 52.950 208.050 53.400 ;
        RECT 337.950 54.600 340.050 55.050 ;
        RECT 355.800 54.600 357.900 55.050 ;
        RECT 394.950 54.600 397.050 55.050 ;
        RECT 337.950 53.400 357.900 54.600 ;
        RECT 359.400 54.000 397.050 54.600 ;
        RECT 337.950 52.950 340.050 53.400 ;
        RECT 355.800 52.950 357.900 53.400 ;
        RECT 358.950 53.400 397.050 54.000 ;
        RECT 16.950 51.600 19.050 52.050 ;
        RECT 31.950 51.600 34.050 52.050 ;
        RECT 16.950 50.400 34.050 51.600 ;
        RECT 16.950 49.950 19.050 50.400 ;
        RECT 31.950 49.950 34.050 50.400 ;
        RECT 58.950 51.600 61.050 52.050 ;
        RECT 85.950 51.600 88.050 52.050 ;
        RECT 58.950 50.400 88.050 51.600 ;
        RECT 58.950 49.950 61.050 50.400 ;
        RECT 85.950 49.950 88.050 50.400 ;
        RECT 142.950 51.600 145.050 52.050 ;
        RECT 151.950 51.600 154.050 52.050 ;
        RECT 199.950 51.600 202.050 52.050 ;
        RECT 142.950 50.400 202.050 51.600 ;
        RECT 142.950 49.950 145.050 50.400 ;
        RECT 151.950 49.950 154.050 50.400 ;
        RECT 199.950 49.950 202.050 50.400 ;
        RECT 232.950 51.600 235.050 52.050 ;
        RECT 238.950 51.600 241.050 52.050 ;
        RECT 343.950 51.600 346.050 52.050 ;
        RECT 232.950 50.400 346.050 51.600 ;
        RECT 232.950 49.950 235.050 50.400 ;
        RECT 238.950 49.950 241.050 50.400 ;
        RECT 343.950 49.950 346.050 50.400 ;
        RECT 358.950 49.950 361.050 53.400 ;
        RECT 394.950 52.950 397.050 53.400 ;
        RECT 418.950 54.600 424.050 55.050 ;
        RECT 448.950 54.600 451.050 55.200 ;
        RECT 418.950 53.400 451.050 54.600 ;
        RECT 418.950 52.950 424.050 53.400 ;
        RECT 448.950 53.100 451.050 53.400 ;
        RECT 466.950 54.600 469.050 55.050 ;
        RECT 472.950 54.600 475.050 55.050 ;
        RECT 466.950 53.400 475.050 54.600 ;
        RECT 508.950 54.600 511.050 58.050 ;
        RECT 544.950 57.600 547.050 58.050 ;
        RECT 592.950 57.600 595.050 58.050 ;
        RECT 544.950 56.400 595.050 57.600 ;
        RECT 544.950 55.950 547.050 56.400 ;
        RECT 592.950 55.950 595.050 56.400 ;
        RECT 628.950 57.600 631.050 58.050 ;
        RECT 727.950 57.600 732.000 58.050 ;
        RECT 736.950 57.600 739.050 58.050 ;
        RECT 754.950 57.600 757.050 58.050 ;
        RECT 628.950 56.400 732.600 57.600 ;
        RECT 736.950 56.400 757.050 57.600 ;
        RECT 628.950 55.950 631.050 56.400 ;
        RECT 727.950 55.950 732.000 56.400 ;
        RECT 736.950 55.950 739.050 56.400 ;
        RECT 754.950 55.950 757.050 56.400 ;
        RECT 520.950 54.600 523.050 55.050 ;
        RECT 565.950 54.600 568.050 55.050 ;
        RECT 508.950 54.000 523.050 54.600 ;
        RECT 557.400 54.000 568.050 54.600 ;
        RECT 509.400 53.400 523.050 54.000 ;
        RECT 466.950 52.950 469.050 53.400 ;
        RECT 472.950 52.950 475.050 53.400 ;
        RECT 520.950 52.950 523.050 53.400 ;
        RECT 556.950 53.400 568.050 54.000 ;
        RECT 448.950 51.600 451.050 51.900 ;
        RECT 460.950 51.600 463.050 52.050 ;
        RECT 448.950 50.400 463.050 51.600 ;
        RECT 448.950 49.800 451.050 50.400 ;
        RECT 460.950 49.950 463.050 50.400 ;
        RECT 493.950 51.600 496.050 52.050 ;
        RECT 508.950 51.600 511.050 51.900 ;
        RECT 493.950 50.400 511.050 51.600 ;
        RECT 493.950 49.950 496.050 50.400 ;
        RECT 508.950 49.800 511.050 50.400 ;
        RECT 556.950 49.950 559.050 53.400 ;
        RECT 565.950 52.950 568.050 53.400 ;
        RECT 760.950 54.600 763.050 55.050 ;
        RECT 802.950 54.600 805.050 55.050 ;
        RECT 760.950 53.400 805.050 54.600 ;
        RECT 760.950 52.950 763.050 53.400 ;
        RECT 802.950 52.950 805.050 53.400 ;
        RECT 631.950 51.600 634.050 52.050 ;
        RECT 649.950 51.600 652.050 52.050 ;
        RECT 667.950 51.600 670.050 52.050 ;
        RECT 706.950 51.600 709.050 52.050 ;
        RECT 631.950 50.400 709.050 51.600 ;
        RECT 631.950 49.950 634.050 50.400 ;
        RECT 649.950 49.950 652.050 50.400 ;
        RECT 667.950 49.950 670.050 50.400 ;
        RECT 706.950 49.950 709.050 50.400 ;
        RECT 769.950 51.600 772.050 52.050 ;
        RECT 775.950 51.600 778.050 52.050 ;
        RECT 769.950 50.400 778.050 51.600 ;
        RECT 769.950 49.950 772.050 50.400 ;
        RECT 775.950 49.950 778.050 50.400 ;
        RECT 409.950 48.600 412.050 49.050 ;
        RECT 418.950 48.600 421.050 49.050 ;
        RECT 409.950 47.400 421.050 48.600 ;
        RECT 409.950 46.950 412.050 47.400 ;
        RECT 418.950 46.950 421.050 47.400 ;
        RECT 13.950 45.600 16.050 46.050 ;
        RECT 19.950 45.600 22.050 46.050 ;
        RECT 13.950 44.400 22.050 45.600 ;
        RECT 13.950 43.950 16.050 44.400 ;
        RECT 19.950 43.950 22.050 44.400 ;
        RECT 127.950 45.600 130.050 46.050 ;
        RECT 145.950 45.600 148.050 46.050 ;
        RECT 127.950 44.400 148.050 45.600 ;
        RECT 127.950 43.950 130.050 44.400 ;
        RECT 145.950 43.950 148.050 44.400 ;
        RECT 208.950 45.600 211.050 46.050 ;
        RECT 259.950 45.600 262.050 46.050 ;
        RECT 208.950 44.400 262.050 45.600 ;
        RECT 208.950 43.950 211.050 44.400 ;
        RECT 259.950 43.950 262.050 44.400 ;
        RECT 292.950 45.600 295.050 46.050 ;
        RECT 322.950 45.600 325.050 46.050 ;
        RECT 292.950 44.400 325.050 45.600 ;
        RECT 292.950 43.950 295.050 44.400 ;
        RECT 322.950 43.950 325.050 44.400 ;
        RECT 421.950 45.600 424.050 46.050 ;
        RECT 439.950 45.600 442.050 46.050 ;
        RECT 421.950 44.400 442.050 45.600 ;
        RECT 421.950 43.950 424.050 44.400 ;
        RECT 439.950 43.950 442.050 44.400 ;
        RECT 685.950 45.600 688.050 46.050 ;
        RECT 772.950 45.600 775.050 46.050 ;
        RECT 685.950 44.400 775.050 45.600 ;
        RECT 685.950 43.950 688.050 44.400 ;
        RECT 772.950 43.950 775.050 44.400 ;
        RECT 37.950 42.600 40.050 43.050 ;
        RECT 43.950 42.600 46.050 43.050 ;
        RECT 37.950 41.400 46.050 42.600 ;
        RECT 37.950 40.950 40.050 41.400 ;
        RECT 43.950 40.950 46.050 41.400 ;
        RECT 61.950 42.600 64.050 43.050 ;
        RECT 82.950 42.600 85.050 43.050 ;
        RECT 61.950 41.400 85.050 42.600 ;
        RECT 61.950 40.950 64.050 41.400 ;
        RECT 82.950 40.950 85.050 41.400 ;
        RECT 373.950 42.600 376.050 43.050 ;
        RECT 529.950 42.600 532.050 43.050 ;
        RECT 577.950 42.600 580.050 43.050 ;
        RECT 373.950 41.400 580.050 42.600 ;
        RECT 373.950 40.950 376.050 41.400 ;
        RECT 529.950 40.950 532.050 41.400 ;
        RECT 577.950 40.950 580.050 41.400 ;
        RECT 745.950 42.600 748.050 42.900 ;
        RECT 787.950 42.600 790.050 43.050 ;
        RECT 745.950 41.400 790.050 42.600 ;
        RECT 745.950 40.800 748.050 41.400 ;
        RECT 787.950 40.950 790.050 41.400 ;
        RECT 88.950 39.600 91.050 40.050 ;
        RECT 187.950 39.600 190.050 40.050 ;
        RECT 88.950 38.400 190.050 39.600 ;
        RECT 88.950 37.950 91.050 38.400 ;
        RECT 187.950 37.950 190.050 38.400 ;
        RECT 247.950 39.600 250.050 40.050 ;
        RECT 256.950 39.600 259.050 40.050 ;
        RECT 247.950 38.400 259.050 39.600 ;
        RECT 247.950 37.950 250.050 38.400 ;
        RECT 256.950 37.950 259.050 38.400 ;
        RECT 481.950 39.600 484.050 40.050 ;
        RECT 493.950 39.600 496.050 40.050 ;
        RECT 481.950 38.400 496.050 39.600 ;
        RECT 481.950 37.950 484.050 38.400 ;
        RECT 493.950 37.950 496.050 38.400 ;
        RECT 262.950 36.600 265.050 37.050 ;
        RECT 268.950 36.600 271.050 37.050 ;
        RECT 262.950 35.400 271.050 36.600 ;
        RECT 262.950 34.950 265.050 35.400 ;
        RECT 268.950 34.950 271.050 35.400 ;
        RECT 316.950 36.600 319.050 37.050 ;
        RECT 367.950 36.600 370.050 37.050 ;
        RECT 316.950 35.400 370.050 36.600 ;
        RECT 316.950 34.950 319.050 35.400 ;
        RECT 367.950 34.950 370.050 35.400 ;
        RECT 607.950 36.600 610.050 37.050 ;
        RECT 619.950 36.600 622.050 37.050 ;
        RECT 607.950 35.400 622.050 36.600 ;
        RECT 607.950 34.950 610.050 35.400 ;
        RECT 619.950 34.950 622.050 35.400 ;
        RECT 742.950 36.600 745.050 37.050 ;
        RECT 781.950 36.600 784.050 37.050 ;
        RECT 742.950 35.400 784.050 36.600 ;
        RECT 742.950 34.950 745.050 35.400 ;
        RECT 781.950 34.950 784.050 35.400 ;
        RECT 787.950 36.600 790.050 37.050 ;
        RECT 808.950 36.600 811.050 37.050 ;
        RECT 787.950 35.400 811.050 36.600 ;
        RECT 787.950 34.950 790.050 35.400 ;
        RECT 808.950 34.950 811.050 35.400 ;
        RECT 304.950 33.600 307.050 34.050 ;
        RECT 310.950 33.600 313.050 34.050 ;
        RECT 322.950 33.600 325.050 34.050 ;
        RECT 379.950 33.600 382.050 34.050 ;
        RECT 304.950 32.400 382.050 33.600 ;
        RECT 304.950 31.950 307.050 32.400 ;
        RECT 310.950 31.950 313.050 32.400 ;
        RECT 322.950 31.950 325.050 32.400 ;
        RECT 379.950 31.950 382.050 32.400 ;
        RECT 487.950 33.600 490.050 34.050 ;
        RECT 538.950 33.600 541.050 34.050 ;
        RECT 487.950 32.400 541.050 33.600 ;
        RECT 487.950 31.950 490.050 32.400 ;
        RECT 538.950 31.950 541.050 32.400 ;
        RECT 559.950 33.600 562.050 34.050 ;
        RECT 574.950 33.600 577.050 34.050 ;
        RECT 559.950 32.400 577.050 33.600 ;
        RECT 559.950 31.950 562.050 32.400 ;
        RECT 574.950 31.950 577.050 32.400 ;
        RECT 19.950 30.600 22.050 31.050 ;
        RECT 49.950 30.600 52.050 31.050 ;
        RECT 19.950 29.400 52.050 30.600 ;
        RECT 19.950 28.950 22.050 29.400 ;
        RECT 49.950 28.950 52.050 29.400 ;
        RECT 76.950 30.600 79.050 31.050 ;
        RECT 118.950 30.600 121.050 31.050 ;
        RECT 133.950 30.600 136.050 31.050 ;
        RECT 76.950 29.400 136.050 30.600 ;
        RECT 76.950 28.950 79.050 29.400 ;
        RECT 118.950 28.950 121.050 29.400 ;
        RECT 133.950 28.950 136.050 29.400 ;
        RECT 391.950 30.600 394.050 31.050 ;
        RECT 415.950 30.600 418.050 31.050 ;
        RECT 391.950 29.400 418.050 30.600 ;
        RECT 391.950 28.950 394.050 29.400 ;
        RECT 415.950 28.950 418.050 29.400 ;
        RECT 13.950 25.950 19.050 28.050 ;
        RECT 37.950 27.600 40.050 28.050 ;
        RECT 64.950 27.600 67.050 28.050 ;
        RECT 106.950 27.600 109.050 28.050 ;
        RECT 112.950 27.600 115.050 28.050 ;
        RECT 37.950 26.400 115.050 27.600 ;
        RECT 37.950 25.950 40.050 26.400 ;
        RECT 64.950 25.950 67.050 26.400 ;
        RECT 106.950 25.950 109.050 26.400 ;
        RECT 112.950 25.950 115.050 26.400 ;
        RECT 283.950 27.600 286.050 28.050 ;
        RECT 289.950 27.600 292.050 28.050 ;
        RECT 283.950 26.400 292.050 27.600 ;
        RECT 283.950 25.950 286.050 26.400 ;
        RECT 289.950 25.950 292.050 26.400 ;
        RECT 316.950 27.600 319.050 28.050 ;
        RECT 325.950 27.600 328.050 28.050 ;
        RECT 421.950 27.600 424.050 28.050 ;
        RECT 316.950 26.400 328.050 27.600 ;
        RECT 410.400 27.000 424.050 27.600 ;
        RECT 316.950 25.950 319.050 26.400 ;
        RECT 325.950 25.950 328.050 26.400 ;
        RECT 409.950 26.400 424.050 27.000 ;
        RECT 70.950 24.600 73.050 25.050 ;
        RECT 88.950 24.600 91.050 25.050 ;
        RECT 70.950 23.400 91.050 24.600 ;
        RECT 70.950 22.950 73.050 23.400 ;
        RECT 88.950 22.950 91.050 23.400 ;
        RECT 142.950 24.600 145.050 25.050 ;
        RECT 154.950 24.600 157.050 25.050 ;
        RECT 142.950 23.400 157.050 24.600 ;
        RECT 142.950 22.950 145.050 23.400 ;
        RECT 154.950 22.950 157.050 23.400 ;
        RECT 184.950 24.600 187.050 25.050 ;
        RECT 202.950 24.600 205.050 25.050 ;
        RECT 184.950 23.400 205.050 24.600 ;
        RECT 184.950 22.950 187.050 23.400 ;
        RECT 202.950 22.950 205.050 23.400 ;
        RECT 211.950 24.600 214.050 25.050 ;
        RECT 226.950 24.600 229.050 25.050 ;
        RECT 211.950 23.400 229.050 24.600 ;
        RECT 211.950 22.950 214.050 23.400 ;
        RECT 226.950 22.950 229.050 23.400 ;
        RECT 232.950 24.600 235.050 25.050 ;
        RECT 271.950 24.600 274.050 25.050 ;
        RECT 232.950 23.400 274.050 24.600 ;
        RECT 232.950 22.950 235.050 23.400 ;
        RECT 271.950 22.950 274.050 23.400 ;
        RECT 343.950 24.600 346.050 25.050 ;
        RECT 397.950 24.600 400.050 25.050 ;
        RECT 343.950 23.400 400.050 24.600 ;
        RECT 343.950 22.950 346.050 23.400 ;
        RECT 397.950 22.950 400.050 23.400 ;
        RECT 409.950 22.950 412.050 26.400 ;
        RECT 421.950 25.950 424.050 26.400 ;
        RECT 436.950 27.600 439.050 28.050 ;
        RECT 442.950 27.600 445.050 28.050 ;
        RECT 436.950 26.400 445.050 27.600 ;
        RECT 451.950 27.600 454.050 31.050 ;
        RECT 709.950 30.600 712.050 31.050 ;
        RECT 715.950 30.600 718.050 31.050 ;
        RECT 709.950 29.400 718.050 30.600 ;
        RECT 709.950 28.950 712.050 29.400 ;
        RECT 715.950 28.950 718.050 29.400 ;
        RECT 778.950 30.600 781.050 31.050 ;
        RECT 802.950 30.600 805.050 31.050 ;
        RECT 778.950 29.400 805.050 30.600 ;
        RECT 778.950 28.950 781.050 29.400 ;
        RECT 802.950 28.950 805.050 29.400 ;
        RECT 466.950 27.600 469.050 28.050 ;
        RECT 451.950 27.000 469.050 27.600 ;
        RECT 452.400 26.400 469.050 27.000 ;
        RECT 436.950 25.950 439.050 26.400 ;
        RECT 442.950 25.950 445.050 26.400 ;
        RECT 466.950 25.950 469.050 26.400 ;
        RECT 472.950 27.600 475.050 28.050 ;
        RECT 478.950 27.600 481.050 28.050 ;
        RECT 565.950 27.600 568.050 28.050 ;
        RECT 472.950 26.400 481.050 27.600 ;
        RECT 472.950 25.950 475.050 26.400 ;
        RECT 478.950 25.950 481.050 26.400 ;
        RECT 539.400 26.400 568.050 27.600 ;
        RECT 539.400 25.050 540.600 26.400 ;
        RECT 565.950 25.950 568.050 26.400 ;
        RECT 571.950 27.600 574.050 28.050 ;
        RECT 601.950 27.600 604.050 28.050 ;
        RECT 673.950 27.600 676.050 28.050 ;
        RECT 763.950 27.600 766.050 28.050 ;
        RECT 571.950 26.400 582.600 27.600 ;
        RECT 571.950 25.950 574.050 26.400 ;
        RECT 526.950 24.600 529.050 25.050 ;
        RECT 538.950 24.600 541.050 25.050 ;
        RECT 526.950 23.400 541.050 24.600 ;
        RECT 526.950 22.950 529.050 23.400 ;
        RECT 538.950 22.950 541.050 23.400 ;
        RECT 547.950 24.600 550.050 25.050 ;
        RECT 577.950 24.600 580.050 25.050 ;
        RECT 547.950 23.400 580.050 24.600 ;
        RECT 547.950 22.950 550.050 23.400 ;
        RECT 577.950 22.950 580.050 23.400 ;
        RECT 10.950 21.600 13.050 22.050 ;
        RECT 19.950 21.600 22.050 22.050 ;
        RECT 10.950 20.400 22.050 21.600 ;
        RECT 10.950 19.950 13.050 20.400 ;
        RECT 19.950 19.950 22.050 20.400 ;
        RECT 34.950 21.600 37.050 22.050 ;
        RECT 43.950 21.600 46.050 22.050 ;
        RECT 34.950 20.400 46.050 21.600 ;
        RECT 34.950 19.950 37.050 20.400 ;
        RECT 43.950 19.950 46.050 20.400 ;
        RECT 166.950 21.600 169.050 22.200 ;
        RECT 581.400 22.050 582.600 26.400 ;
        RECT 601.950 26.400 766.050 27.600 ;
        RECT 601.950 25.950 604.050 26.400 ;
        RECT 673.950 25.950 676.050 26.400 ;
        RECT 763.950 25.950 766.050 26.400 ;
        RECT 589.950 24.600 592.050 25.050 ;
        RECT 625.950 24.600 628.050 25.050 ;
        RECT 589.950 23.400 628.050 24.600 ;
        RECT 589.950 22.950 592.050 23.400 ;
        RECT 625.950 22.950 628.050 23.400 ;
        RECT 655.950 24.600 658.050 25.050 ;
        RECT 661.950 24.600 664.050 25.050 ;
        RECT 655.950 23.400 664.050 24.600 ;
        RECT 655.950 22.950 658.050 23.400 ;
        RECT 661.950 22.950 664.050 23.400 ;
        RECT 181.950 21.600 184.050 22.050 ;
        RECT 166.950 20.400 184.050 21.600 ;
        RECT 166.950 20.100 169.050 20.400 ;
        RECT 181.950 19.950 184.050 20.400 ;
        RECT 289.950 19.950 295.050 22.050 ;
        RECT 313.950 21.600 316.050 22.050 ;
        RECT 337.950 21.600 340.050 22.050 ;
        RECT 361.950 21.600 364.050 22.050 ;
        RECT 313.950 20.400 340.050 21.600 ;
        RECT 347.400 21.000 364.050 21.600 ;
        RECT 313.950 19.950 316.050 20.400 ;
        RECT 337.950 19.950 340.050 20.400 ;
        RECT 346.950 20.400 364.050 21.000 ;
        RECT 40.950 18.600 43.050 19.050 ;
        RECT 61.950 18.600 64.050 19.050 ;
        RECT 40.950 17.400 64.050 18.600 ;
        RECT 40.950 16.950 43.050 17.400 ;
        RECT 61.950 16.950 64.050 17.400 ;
        RECT 100.950 18.600 103.050 19.050 ;
        RECT 124.950 18.600 127.050 19.050 ;
        RECT 148.950 18.600 151.050 19.050 ;
        RECT 100.950 17.400 151.050 18.600 ;
        RECT 100.950 16.950 103.050 17.400 ;
        RECT 124.950 16.950 127.050 17.400 ;
        RECT 148.950 16.950 151.050 17.400 ;
        RECT 163.950 18.900 168.000 19.050 ;
        RECT 163.950 16.950 169.050 18.900 ;
        RECT 247.950 18.600 250.050 19.050 ;
        RECT 301.950 18.600 304.050 19.050 ;
        RECT 247.950 17.400 304.050 18.600 ;
        RECT 247.950 16.950 250.050 17.400 ;
        RECT 301.950 16.950 304.050 17.400 ;
        RECT 346.950 16.950 349.050 20.400 ;
        RECT 361.950 19.950 364.050 20.400 ;
        RECT 379.950 21.600 382.050 22.050 ;
        RECT 391.950 21.600 394.050 22.050 ;
        RECT 379.950 20.400 394.050 21.600 ;
        RECT 379.950 19.950 382.050 20.400 ;
        RECT 391.950 19.950 394.050 20.400 ;
        RECT 580.950 19.950 583.050 22.050 ;
        RECT 586.950 21.600 589.050 22.050 ;
        RECT 656.400 21.600 657.600 22.950 ;
        RECT 586.950 20.400 657.600 21.600 ;
        RECT 679.950 21.600 682.050 25.050 ;
        RECT 724.950 24.600 727.050 25.050 ;
        RECT 739.950 24.600 742.050 25.050 ;
        RECT 724.950 23.400 742.050 24.600 ;
        RECT 724.950 22.950 727.050 23.400 ;
        RECT 739.950 22.950 742.050 23.400 ;
        RECT 745.950 24.600 748.050 25.050 ;
        RECT 751.950 24.600 754.050 25.050 ;
        RECT 745.950 23.400 754.050 24.600 ;
        RECT 745.950 22.950 748.050 23.400 ;
        RECT 751.950 22.950 754.050 23.400 ;
        RECT 793.950 24.600 796.050 25.050 ;
        RECT 811.950 24.600 814.050 25.050 ;
        RECT 793.950 23.400 814.050 24.600 ;
        RECT 793.950 22.950 796.050 23.400 ;
        RECT 811.950 22.950 814.050 23.400 ;
        RECT 694.950 21.600 697.050 22.050 ;
        RECT 679.950 21.000 697.050 21.600 ;
        RECT 680.400 20.400 697.050 21.000 ;
        RECT 586.950 19.950 589.050 20.400 ;
        RECT 694.950 19.950 697.050 20.400 ;
        RECT 448.950 18.600 451.050 19.050 ;
        RECT 550.950 18.600 553.050 19.050 ;
        RECT 448.950 17.400 553.050 18.600 ;
        RECT 448.950 16.950 451.050 17.400 ;
        RECT 550.950 16.950 553.050 17.400 ;
        RECT 568.950 16.950 574.050 19.050 ;
        RECT 631.950 18.600 634.050 19.050 ;
        RECT 649.950 18.600 652.050 19.050 ;
        RECT 631.950 17.400 652.050 18.600 ;
        RECT 631.950 16.950 634.050 17.400 ;
        RECT 649.950 16.950 652.050 17.400 ;
        RECT 796.950 18.600 799.050 19.050 ;
        RECT 802.950 18.600 805.050 19.050 ;
        RECT 796.950 17.400 805.050 18.600 ;
        RECT 796.950 16.950 799.050 17.400 ;
        RECT 802.950 16.950 805.050 17.400 ;
        RECT 166.950 16.800 169.050 16.950 ;
        RECT 112.950 15.600 115.050 16.050 ;
        RECT 142.950 15.600 145.050 16.050 ;
        RECT 112.950 14.400 145.050 15.600 ;
        RECT 112.950 13.950 115.050 14.400 ;
        RECT 142.950 13.950 145.050 14.400 ;
        RECT 187.950 15.600 190.050 16.050 ;
        RECT 316.950 15.600 319.050 16.050 ;
        RECT 187.950 14.400 319.050 15.600 ;
        RECT 187.950 13.950 190.050 14.400 ;
        RECT 316.950 13.950 319.050 14.400 ;
        RECT 364.950 15.600 367.050 16.050 ;
        RECT 442.950 15.600 445.050 16.050 ;
        RECT 364.950 14.400 445.050 15.600 ;
        RECT 364.950 13.950 367.050 14.400 ;
        RECT 442.950 13.950 445.050 14.400 ;
        RECT 565.950 15.600 568.050 16.050 ;
        RECT 625.950 15.600 628.050 16.050 ;
        RECT 565.950 14.400 628.050 15.600 ;
        RECT 565.950 13.950 568.050 14.400 ;
        RECT 625.950 13.950 628.050 14.400 ;
        RECT 730.950 15.600 733.050 16.050 ;
        RECT 742.950 15.600 745.050 16.050 ;
        RECT 778.950 15.600 781.050 16.050 ;
        RECT 730.950 14.400 781.050 15.600 ;
        RECT 730.950 13.950 733.050 14.400 ;
        RECT 742.950 13.950 745.050 14.400 ;
        RECT 778.950 13.950 781.050 14.400 ;
        RECT 58.950 12.600 61.050 13.050 ;
        RECT 70.950 12.600 73.050 13.050 ;
        RECT 58.950 11.400 73.050 12.600 ;
        RECT 58.950 10.950 61.050 11.400 ;
        RECT 70.950 10.950 73.050 11.400 ;
        RECT 82.950 12.600 85.050 13.050 ;
        RECT 175.950 12.600 178.050 13.050 ;
        RECT 82.950 11.400 178.050 12.600 ;
        RECT 82.950 10.950 85.050 11.400 ;
        RECT 175.950 10.950 178.050 11.400 ;
        RECT 337.950 12.600 340.050 13.050 ;
        RECT 370.950 12.600 373.050 13.050 ;
        RECT 337.950 11.400 373.050 12.600 ;
        RECT 337.950 10.950 340.050 11.400 ;
        RECT 370.950 10.950 373.050 11.400 ;
        RECT 646.950 12.600 649.050 13.050 ;
        RECT 700.950 12.600 703.050 13.050 ;
        RECT 646.950 11.400 703.050 12.600 ;
        RECT 646.950 10.950 649.050 11.400 ;
        RECT 700.950 10.950 703.050 11.400 ;
        RECT 736.950 12.600 739.050 13.050 ;
        RECT 781.950 12.600 784.050 13.050 ;
        RECT 736.950 11.400 784.050 12.600 ;
        RECT 736.950 10.950 739.050 11.400 ;
        RECT 781.950 10.950 784.050 11.400 ;
        RECT 298.950 9.600 301.050 10.050 ;
        RECT 364.950 9.600 367.050 10.050 ;
        RECT 298.950 8.400 367.050 9.600 ;
        RECT 298.950 7.950 301.050 8.400 ;
        RECT 364.950 7.950 367.050 8.400 ;
        RECT 367.950 6.600 370.050 7.050 ;
        RECT 478.950 6.600 481.050 7.050 ;
        RECT 367.950 5.400 481.050 6.600 ;
        RECT 367.950 4.950 370.050 5.400 ;
        RECT 478.950 4.950 481.050 5.400 ;
  END
END fir_pe
END LIBRARY

