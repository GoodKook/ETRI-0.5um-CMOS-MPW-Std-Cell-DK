magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect -34 78 124 159
<< nwell >>
rect -14 154 113 272
<< ntransistor >>
rect 22 14 26 34
rect 64 14 68 54
rect 74 14 78 54
<< ptransistor >>
rect 22 206 26 246
rect 64 166 68 246
rect 74 166 78 246
<< ndiffusion >>
rect 20 14 22 34
rect 26 14 28 34
rect 62 14 64 54
rect 68 14 74 54
rect 78 14 80 54
<< pdiffusion >>
rect 20 206 22 246
rect 26 206 28 246
rect 62 166 64 246
rect 68 166 74 246
rect 78 166 80 246
<< ndcontact >>
rect 8 14 20 34
rect 28 14 40 34
rect 50 14 62 54
rect 80 14 92 54
<< pdcontact >>
rect 8 206 20 246
rect 28 206 40 246
rect 50 166 62 246
rect 80 166 92 246
<< psubstratepcontact >>
rect -7 -6 107 6
<< nsubstratencontact >>
rect -7 254 107 266
<< polysilicon >>
rect 22 246 26 250
rect 64 246 68 250
rect 74 246 78 250
rect 22 128 26 206
rect 64 149 68 166
rect 46 145 68 149
rect 74 128 78 166
rect 20 116 26 128
rect 22 60 26 116
rect 22 56 68 60
rect 22 34 26 56
rect 64 54 68 56
rect 74 54 78 116
rect 22 10 26 14
rect 64 10 68 14
rect 74 10 78 14
<< polycontact >>
rect 34 145 46 157
rect 8 116 20 128
rect 72 116 84 128
<< metal1 >>
rect -7 266 107 268
rect -7 252 107 254
rect 8 246 20 252
rect 80 246 92 252
rect 34 157 40 206
rect 34 34 40 145
rect 53 117 60 166
rect 53 54 60 103
rect 8 8 20 14
rect 80 8 92 14
rect -7 6 107 8
rect -7 -8 107 -6
<< m2contact >>
rect 6 116 8 117
rect 8 116 20 117
rect 6 103 20 116
rect 46 103 60 117
rect 70 116 72 117
rect 72 116 84 117
rect 70 103 84 116
<< metal2 >>
rect 6 117 14 134
rect 46 117 54 134
rect 76 117 84 134
<< m1p >>
rect -7 252 107 268
rect -7 -8 107 8
<< m2p >>
rect 6 119 14 134
rect 46 119 54 134
rect 76 119 84 134
<< labels >>
rlabel metal2 80 131 80 131 7 A
port 1 n signal input
rlabel metal2 10 131 10 131 1 EN
port 2 n signal input
rlabel metal2 50 131 50 131 1 Y
port 3 n signal output
rlabel metal1 -7 252 107 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -7 -8 107 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
