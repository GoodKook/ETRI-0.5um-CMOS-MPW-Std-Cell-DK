magic
tech scmos
magscale 1 30
timestamp 1719895877
<< checkpaint >>
rect 47800 171700 61200 180850
rect 18300 145440 61200 171700
rect 18300 145200 44800 145440
rect 47800 145200 61200 145440
rect 61300 145200 74700 180850
rect 74800 145200 88200 180850
rect 88300 146970 101700 180850
rect 101900 146970 115100 180850
rect 88300 145200 115100 146970
rect 115300 145200 128700 180850
rect 128800 171700 142200 180850
rect 128800 145440 171700 171700
rect 128800 145200 142200 145440
rect 145200 145200 171700 145440
rect 18300 142200 44650 145200
rect 9150 128800 44800 142200
rect 101100 140200 103040 145200
rect 145440 142200 171700 145200
rect 145200 128800 180850 142200
rect 9150 115300 44800 128700
rect 145200 115300 180850 128700
rect 9150 101800 44800 115200
rect 145200 101800 180850 115200
rect 9150 88300 44800 101700
rect 145200 88300 180850 101700
rect 9150 74900 44800 88100
rect 45930 85530 47165 85855
rect 45055 77480 47165 85530
rect 145200 74800 180850 88200
rect 9150 61300 44800 74700
rect 145200 61300 180850 74700
rect 9150 47800 44800 61200
rect 145200 47800 180850 61200
rect 18300 44800 44560 47800
rect 97740 45875 100710 47165
rect 99000 45640 100610 45875
rect 145440 44800 171700 47800
rect 18300 44560 44800 44800
rect 47800 44560 61200 44800
rect 18300 18300 61200 44560
rect 47800 9150 61200 18300
rect 61300 9150 74700 44800
rect 74800 9150 88200 44800
rect 88300 9150 101700 44800
rect 101800 9150 115200 44800
rect 115300 9150 128700 44800
rect 128800 44560 142200 44800
rect 145200 44560 171700 44800
rect 128800 18300 171700 44560
rect 128800 9150 142200 18300
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI050
timestamp 1709081121
transform 0 -1 171100 -1 0 75646
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_1
timestamp 1709081121
transform 0 -1 171100 -1 0 62146
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_2
timestamp 1709081121
transform 0 -1 171100 -1 0 102646
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_3
timestamp 1709081121
transform 0 -1 171100 -1 0 89146
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_4
timestamp 1709081121
transform 0 -1 171100 -1 0 129646
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_5
timestamp 1709081121
transform 0 -1 171100 -1 0 116146
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_6
timestamp 1709081121
transform 1 0 73845 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_7
timestamp 1709081121
transform 1 0 60345 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_8
timestamp 1709081121
transform 1 0 100845 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_9
timestamp 1709081121
transform 1 0 87345 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_10
timestamp 1709081121
transform 1 0 127845 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_11
timestamp 1709081121
transform 1 0 114345 0 1 18900
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_12
timestamp 1709081121
transform 0 1 18900 -1 0 75655
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_13
timestamp 1709081121
transform 0 1 18900 -1 0 62155
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_14
timestamp 1709081121
transform 0 1 18900 -1 0 102655
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_15
timestamp 1709081121
transform 0 1 18900 -1 0 89155
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_16
timestamp 1709081121
transform 1 0 73845 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_17
timestamp 1709081121
transform 0 1 18900 -1 0 116155
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_18
timestamp 1709081121
transform 0 1 18900 -1 0 129655
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_19
timestamp 1709081121
transform 1 0 60345 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_20
timestamp 1709081121
transform 1 0 100845 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_21
timestamp 1709081121
transform 1 0 87345 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_22
timestamp 1709081121
transform 1 0 127845 0 -1 171099
box 0 0 1810 25060
use IOFILLER18  IOFILLER18_23
timestamp 1709081121
transform 1 0 114345 0 -1 171099
box 0 0 1810 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 43675 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1537935238
transform 1 0 141375 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1537935238
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1537935238
transform 1 0 43675 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1537935238
transform 0 1 18900 -1 0 48685
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1537935238
transform 0 1 18900 -1 0 146205
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1537935238
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1537935238
transform 0 -1 171100 -1 0 146325
box -35 0 5035 25060
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1537935238
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1537935238
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1537935238
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  CIN0_2 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN1_6
timestamp 1537935238
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN2_5
timestamp 1537935238
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN3_11
timestamp 1537935238
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use PIC  CIN4_15
timestamp 1537935238
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  CIN5_16
timestamp 1537935238
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC  CIN6_17
timestamp 1537935238
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC  CLK_4
timestamp 1537935238
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PIC  RDY_3
timestamp 1537935238
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  XIN0_12
timestamp 1537935238
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  XIN1_9
timestamp 1537935238
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN2_27
timestamp 1537935238
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  XIN3_13
timestamp 1537935238
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PIC  YIN0_1
timestamp 1537935238
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN1_0
timestamp 1537935238
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PIC  YIN2_7
timestamp 1537935238
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PIC  YIN3_8
timestamp 1537935238
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use POB8  VLD_14 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use POB8  XOUT0_24
timestamp 1537935238
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT1_23
timestamp 1537935238
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT2_21
timestamp 1537935238
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT3_20
timestamp 1537935238
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT0_19
timestamp 1537935238
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use POB8  YOUT1_18
timestamp 1537935238
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use POB8  YOUT2_25
timestamp 1537935238
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT3_26
timestamp 1537935238
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PVSS  PVSS_22 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 1 0 102500 0 -1 171100
box 0 -9150 12000 25300
use PVDD  PVDD_10 ~/ETRI050_DesignKit/devel/Ref_Design/FIR8/2_Splited_IO/MPW_Submit/2_Splited_IO/chiptop
timestamp 1537935238
transform 0 1 18900 -1 0 87500
box 0 -9150 12000 25300
<< end >>