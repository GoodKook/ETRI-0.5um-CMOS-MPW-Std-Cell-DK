magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -56 -56 164 164
<< diffusion >>
rect 5 5 103 103
<< metal1 >>
rect 4 4 104 104
<< end >>
