magic
tech scmos
magscale 1 2
timestamp 1702309798
<< nwell >>
rect -13 154 133 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 48 14 52 54
rect 68 14 72 54
rect 78 14 82 54
rect 98 14 102 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 48 166 52 246
rect 68 166 72 246
rect 78 166 82 246
rect 98 166 102 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 48 38 54
rect 22 14 24 48
rect 36 14 38 48
rect 42 14 48 54
rect 52 14 54 54
rect 66 14 68 54
rect 72 14 78 54
rect 82 48 98 54
rect 82 14 84 48
rect 96 14 98 48
rect 102 14 104 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 180 24 246
rect 36 180 38 246
rect 22 166 38 180
rect 42 166 48 246
rect 52 166 54 246
rect 66 166 68 246
rect 72 166 78 246
rect 82 180 84 246
rect 96 180 98 246
rect 82 166 98 180
rect 102 166 104 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 48
rect 54 14 66 54
rect 84 14 96 48
rect 104 14 116 54
<< pdcontact >>
rect 4 166 16 246
rect 24 180 36 246
rect 54 166 66 246
rect 84 180 96 246
rect 104 166 116 246
<< psubstratepcontact >>
rect -7 -6 127 6
<< nsubstratencontact >>
rect -7 254 127 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 48 246 52 250
rect 68 246 72 250
rect 78 246 82 250
rect 98 246 102 250
rect 18 54 22 166
rect 38 161 42 166
rect 27 157 42 161
rect 27 141 31 157
rect 48 153 52 166
rect 68 154 72 166
rect 78 164 82 166
rect 98 164 102 166
rect 78 159 102 164
rect 48 149 55 153
rect 68 150 85 154
rect 27 129 30 141
rect 27 63 31 129
rect 50 121 55 149
rect 53 115 55 121
rect 53 110 65 115
rect 81 111 85 150
rect 27 59 42 63
rect 38 54 42 59
rect 48 54 52 87
rect 61 62 65 110
rect 98 69 102 159
rect 78 64 102 69
rect 61 56 72 62
rect 68 54 72 56
rect 78 54 82 64
rect 98 54 102 64
rect 18 10 22 14
rect 38 10 42 14
rect 48 10 52 14
rect 68 10 72 14
rect 78 10 82 14
rect 98 10 102 14
<< polycontact >>
rect 6 105 18 117
rect 30 129 42 141
rect 41 109 53 121
rect 41 87 53 99
rect 73 99 85 111
rect 102 105 114 117
<< metal1 >>
rect -7 266 127 268
rect -7 252 127 254
rect 24 246 36 252
rect 84 246 96 252
rect 16 166 35 172
rect 59 156 66 166
rect 98 166 104 174
rect 59 149 74 156
rect 3 123 17 137
rect 63 137 74 149
rect 63 123 77 137
rect 103 123 117 137
rect 6 117 17 123
rect 18 109 41 117
rect 59 117 74 123
rect 103 117 114 123
rect 9 66 53 73
rect 9 54 16 66
rect 59 57 66 117
rect 59 54 77 57
rect 98 54 116 61
rect 66 43 77 54
rect 24 8 36 14
rect 84 8 96 14
rect -7 6 127 8
rect -7 -8 127 -6
<< m2contact >>
rect 21 152 35 166
rect 84 160 98 174
rect 42 129 56 143
rect 39 73 53 87
rect 72 85 86 99
rect 84 54 98 68
<< metal2 >>
rect 26 87 32 152
rect 50 118 56 129
rect 92 118 98 160
rect 50 112 98 118
rect 47 87 72 93
rect 26 80 39 87
rect 53 86 72 87
rect 92 68 98 112
<< m1p >>
rect -7 252 127 268
rect 3 123 17 137
rect 63 123 77 137
rect 103 123 117 137
rect 63 43 77 57
rect -7 -8 127 8
<< labels >>
rlabel nsubstratencontact 60 260 60 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 60 0 60 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 126 10 126 0 A
port 1 nsew signal input
rlabel metal1 70 130 70 130 0 Y
port 3 nsew signal output
rlabel metal1 110 130 110 130 0 B
port 2 nsew signal input
rlabel metal1 70 50 70 50 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
