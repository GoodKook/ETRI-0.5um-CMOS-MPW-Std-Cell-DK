magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect -17 39 57 79
rect 3 30 47 39
<< nwell >>
rect -6 77 47 136
<< ntransistor >>
rect 9 7 11 27
rect 14 7 16 27
rect 24 7 26 27
<< ptransistor >>
rect 9 103 11 123
rect 19 103 21 123
rect 29 83 31 123
<< ndiffusion >>
rect 8 7 9 27
rect 11 7 14 27
rect 16 7 17 27
rect 23 7 24 27
rect 26 7 27 27
<< pdiffusion >>
rect 8 103 9 123
rect 11 103 12 123
rect 18 103 19 123
rect 21 103 22 123
rect 28 85 29 123
rect 24 83 29 85
rect 31 83 32 123
<< ndcontact >>
rect 2 7 8 27
rect 17 7 23 27
rect 27 7 33 27
<< pdcontact >>
rect 2 103 8 123
rect 12 103 18 123
rect 22 85 28 123
rect 32 83 38 123
<< psubstratepcontact >>
rect -3 -3 43 3
<< nsubstratencontact >>
rect -3 127 43 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 9 102 11 103
rect 5 100 11 102
rect 5 51 7 100
rect 19 64 21 103
rect 5 31 7 45
rect 19 42 21 58
rect 14 40 21 42
rect 5 29 11 31
rect 9 27 11 29
rect 14 27 16 40
rect 29 36 31 83
rect 30 30 31 36
rect 24 27 26 30
rect 9 5 11 7
rect 14 5 16 7
rect 24 5 26 7
<< polycontact >>
rect 19 58 25 64
rect 2 45 8 51
rect 24 30 30 36
<< metal1 >>
rect -3 133 43 134
rect -3 126 43 127
rect 2 123 8 126
rect 22 123 28 126
rect 12 36 15 103
rect 33 58 36 83
rect 2 33 24 36
rect 2 27 8 33
rect 33 21 36 51
rect 17 4 23 7
rect -3 3 43 4
rect -3 -4 43 -3
<< m2contact >>
rect 2 51 9 58
rect 20 51 27 58
rect 31 51 38 58
<< metal2 >>
rect 3 58 7 67
rect 33 58 37 67
rect 23 43 27 51
<< m1p >>
rect -3 126 43 134
rect -3 -4 43 4
<< m2p >>
rect 3 59 7 67
rect 33 59 37 67
rect 23 43 27 50
<< labels >>
rlabel metal2 5 66 5 66 1 A
port 1 n signal input
rlabel metal2 25 44 25 44 1 B
port 2 n signal input
rlabel metal2 35 65 35 65 5 Y
port 3 n signal output
rlabel metal1 -3 126 43 134 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -3 -4 43 4 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 40 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
