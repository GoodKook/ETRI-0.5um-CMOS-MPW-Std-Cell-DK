magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -15 -15 505 505
<< nwell >>
rect 110 110 380 380
<< pdiffusion >>
rect 195 195 295 295
<< psubstratepdiff >>
rect 45 425 445 445
rect 45 65 65 425
rect 425 65 445 425
rect 45 45 445 65
<< nsubstratendiff >>
rect 130 340 360 360
rect 130 150 150 340
rect 340 150 360 340
rect 130 130 360 150
<< metal1 >>
rect 45 425 445 445
rect 45 65 65 425
rect 130 340 360 360
rect 130 150 150 340
rect 195 195 295 295
rect 340 150 360 340
rect 130 130 360 150
rect 425 65 445 425
rect 45 45 445 65
use ntap_CDNS_723012252911  ntap_CDNS_723012252911_0
timestamp 1723012252
transform 1 0 336 0 1 146
box 4 4 24 194
use ntap_CDNS_723012252911  ntap_CDNS_723012252911_1
timestamp 1723012252
transform 0 1 146 1 0 126
box 4 4 24 194
use ntap_CDNS_723012252911  ntap_CDNS_723012252911_2
timestamp 1723012252
transform 0 1 146 1 0 336
box 4 4 24 194
use ntap_CDNS_723012252911  ntap_CDNS_723012252911_3
timestamp 1723012252
transform 1 0 126 0 1 146
box 4 4 24 194
use ptap_CDNS_723012252912  ptap_CDNS_723012252912_0
timestamp 1723012252
transform 0 1 71 1 0 41
box 4 4 24 344
use ptap_CDNS_723012252912  ptap_CDNS_723012252912_1
timestamp 1723012252
transform 1 0 421 0 1 71
box 4 4 24 344
use ptap_CDNS_723012252912  ptap_CDNS_723012252912_2
timestamp 1723012252
transform 1 0 41 0 1 71
box 4 4 24 344
use ptap_CDNS_723012252912  ptap_CDNS_723012252912_3
timestamp 1723012252
transform 0 1 71 1 0 421
box 4 4 24 344
use ptap_CDNS_723012252913  ptap_CDNS_723012252913_0
timestamp 1723012252
transform 1 0 191 0 1 191
box 4 4 104 104
<< end >>
