magic
tech scmos
magscale 1 2
timestamp 1726836989
<< nwell >>
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 74
rect 30 14 34 74
rect 44 14 48 74
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 60 206 64 246
<< ndiffusion >>
rect 18 14 20 74
rect 24 14 30 74
rect 34 14 44 74
rect 48 72 62 74
rect 48 14 50 72
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 210 46 246
rect 58 210 60 246
rect 44 206 60 210
rect 64 206 66 246
<< ndcontact >>
rect 6 14 18 74
rect 50 14 62 72
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 46 210 58 246
rect 66 206 78 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 20 194 24 206
rect 40 194 44 206
rect 10 190 24 194
rect 30 190 44 194
rect 10 103 16 190
rect 30 129 34 190
rect 10 82 16 91
rect 10 78 24 82
rect 20 74 24 78
rect 30 74 34 117
rect 60 103 64 206
rect 56 91 64 103
rect 53 82 57 91
rect 44 78 57 82
rect 44 74 48 78
rect 20 10 24 14
rect 30 10 34 14
rect 44 10 48 14
<< polycontact >>
rect 24 117 36 129
rect 4 91 16 103
rect 44 91 56 103
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 6 246 18 252
rect 46 246 58 252
rect 28 204 38 206
rect 66 204 72 206
rect 28 198 72 204
rect 66 117 72 198
rect 66 78 72 103
rect 50 72 72 78
rect 62 70 72 72
rect 6 8 18 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
rect 43 103 57 117
rect 63 103 77 117
<< metal2 >>
rect 6 117 14 135
rect 46 117 54 135
rect 26 87 34 103
rect 66 87 74 103
<< m1p >>
rect -6 252 106 268
rect -6 -8 106 8
<< m2p >>
rect 6 119 14 135
rect 46 119 54 135
rect 26 87 34 101
rect 66 87 74 101
<< labels >>
rlabel metal1 -6 252 86 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal2 10 131 10 131 1 A
port 1 n signal input
rlabel metal2 30 91 30 91 5 B
port 2 n signal input
rlabel metal2 50 131 50 131 1 C
port 3 n signal input
rlabel metal2 70 89 70 89 5 Y
port 4 n signal output
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
