magic
tech scmos
magscale 1 2
timestamp 1702308645
<< nwell >>
rect -13 154 173 272
<< ntransistor >>
rect 38 14 42 34
rect 58 14 62 34
rect 78 14 82 34
<< ptransistor >>
rect 18 186 22 246
rect 38 186 42 246
rect 58 186 62 246
rect 78 186 82 246
rect 118 178 122 238
rect 138 178 142 238
<< ndiffusion >>
rect 36 14 38 34
rect 42 14 44 34
rect 56 14 58 34
rect 62 14 64 34
rect 76 14 78 34
rect 82 14 84 34
<< pdiffusion >>
rect 16 186 18 246
rect 22 186 24 246
rect 36 186 38 246
rect 42 186 44 246
rect 56 186 58 246
rect 62 234 78 246
rect 62 186 64 234
rect 76 186 78 234
rect 82 188 84 246
rect 82 186 88 188
rect 116 178 118 238
rect 122 234 138 238
rect 122 182 124 234
rect 136 182 138 234
rect 122 178 138 182
rect 142 178 144 238
<< ndcontact >>
rect 23 14 36 34
rect 44 14 56 34
rect 64 14 76 34
rect 84 14 96 34
<< pdcontact >>
rect 4 186 16 246
rect 24 186 36 246
rect 44 186 56 246
rect 64 186 76 234
rect 84 188 96 246
rect 104 178 116 238
rect 124 182 136 234
rect 144 178 156 238
<< psubstratepcontact >>
rect -7 -6 167 6
<< nsubstratencontact >>
rect -7 254 167 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 78 246 82 250
rect 118 238 122 242
rect 138 238 142 242
rect 18 184 22 186
rect 38 184 42 186
rect 18 180 42 184
rect 38 117 42 180
rect 37 105 42 117
rect 38 34 42 105
rect 58 184 62 186
rect 78 184 82 186
rect 58 180 82 184
rect 58 99 62 180
rect 118 176 122 178
rect 138 176 142 178
rect 118 172 142 176
rect 118 170 122 172
rect 58 34 62 87
rect 78 166 122 170
rect 78 105 83 166
rect 78 34 82 105
rect 38 10 42 14
rect 58 10 62 14
rect 78 10 82 14
<< polycontact >>
rect 25 105 37 117
rect 50 87 62 99
rect 83 105 95 117
<< metal1 >>
rect -7 266 167 268
rect -7 252 167 254
rect 24 246 36 252
rect 56 240 84 246
rect 4 180 16 186
rect 44 180 56 186
rect 4 174 56 180
rect 104 240 156 246
rect 104 238 116 240
rect 64 182 76 186
rect 64 178 104 182
rect 144 238 156 240
rect 64 176 116 178
rect 124 150 132 182
rect 106 143 132 150
rect 23 123 37 137
rect 25 117 37 123
rect 83 123 97 137
rect 83 117 95 123
rect 106 117 114 143
rect 43 103 57 117
rect 103 103 117 117
rect 46 99 57 103
rect 46 87 50 99
rect 106 47 114 103
rect 48 40 114 47
rect 48 34 54 40
rect 96 14 102 40
rect 23 8 36 14
rect 64 8 76 14
rect -7 6 167 8
rect -7 -8 167 -6
<< m1p >>
rect -7 252 167 268
rect 23 123 37 137
rect 83 123 97 137
rect 43 103 57 117
rect 103 103 117 117
rect -7 -8 167 8
<< labels >>
rlabel nsubstratencontact 80 260 80 260 0 vdd
port 5 nsew power bidirectional abutment
rlabel psubstratepcontact 80 0 80 0 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 30 127 30 127 0 A
port 1 nsew signal input
rlabel metal1 90 127 90 127 0 C
port 3 nsew signal input
rlabel metal1 50 107 50 107 0 B
port 2 nsew signal input
rlabel metal1 110 111 110 111 0 Y
port 4 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 160 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
