magic
tech scmos
magscale 1 2
timestamp 1726531033
<< nwell >>
rect -12 154 72 272
<< ntransistor >>
rect 20 14 24 34
<< ptransistor >>
rect 20 206 24 246
<< ndiffusion >>
rect 18 14 20 34
rect 24 14 26 34
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
<< ndcontact >>
rect 6 14 18 34
rect 26 14 38 34
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 20 246 24 250
rect 20 129 24 206
rect 16 117 24 129
rect 20 34 24 117
rect 20 10 24 14
<< polycontact >>
rect 4 117 16 129
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 6 246 18 252
rect 26 117 34 206
rect 26 34 34 103
rect 6 8 18 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
<< metal2 >>
rect 26 117 34 134
rect 6 86 14 103
<< m1p >>
rect -6 252 66 268
rect -6 -8 66 8
<< m2p >>
rect 26 119 34 134
rect 6 86 14 101
<< labels >>
rlabel metal1 -6 252 46 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 46 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal2 10 90 10 90 1 A
port 1 n signal input
rlabel metal2 28 128 28 128 1 Y
port 2 n signal output
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
