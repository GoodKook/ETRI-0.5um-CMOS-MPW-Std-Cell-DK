magic
tech scmos
magscale 1 30
timestamp 1569139307
<< checkpaint >>
rect -600 -600 12600 25900
<< metal1 >>
rect 5801 21703 6898 22103
rect 8011 21703 8531 22103
rect 500 20800 5610 21000
rect 1035 18300 2145 18500
rect 2295 18300 11700 18600
rect 600 7000 1420 7200
rect 1965 7000 11700 7300
<< metal2 >>
rect 11370 24010 11550 25300
rect 500 20800 930 21000
rect 1510 20800 2880 21000
rect 0 11300 400 19100
rect 60 7800 400 10800
rect 0 0 400 7800
rect 500 7200 600 20800
rect 1510 18300 1870 20800
rect 500 7000 975 7200
rect 1320 700 1860 18200
rect 2580 700 3120 18200
rect 3840 700 4380 18200
rect 5100 700 5640 18200
rect 6360 700 6900 22103
rect 7460 20600 7825 23855
rect 8010 23085 8610 23952
rect 8010 22860 9080 23085
rect 9620 22860 10490 23080
rect 8010 21703 8531 22860
rect 7460 19580 8710 20600
rect 7620 700 8160 18200
rect 8880 700 9420 18200
rect 10140 700 10680 18200
rect 11500 11300 12000 19100
rect 11500 8300 11940 11300
rect 1320 0 10680 700
rect 11500 0 12000 7800
use p2res_CDNS_704676826056  p2res_CDNS_704676826056_0
timestamp 1569139307
transform 1 0 5650 0 1 21625
box 80 80 2720 480
use VIA1  VIA1_0
timestamp 1569139307
transform 1 0 1770 0 1 18400
box -40 -40 40 40
use VIA1  VIA1_1
array 0 0 0 0 1 160
timestamp 1569139307
transform 1 0 8431 0 1 21818
box -40 -40 40 40
use VIA1  VIA1_2
timestamp 1569139307
transform 1 0 830 0 1 20900
box -40 -40 40 40
use VIA1  VIA1_3
timestamp 1569139307
transform 1 0 670 0 1 20900
box -40 -40 40 40
use VIA1  VIA1_4
array 0 1 160 0 1 160
timestamp 1569139307
transform 1 0 6536 0 1 21818
box -40 -40 40 40
use VIA1  VIA1_5
timestamp 1569139307
transform 1 0 1610 0 1 18400
box -40 -40 40 40
use VIA1  VIA1_6
array 0 1 160 0 0 0
timestamp 1569139307
transform 1 0 700 0 1 7100
box -40 -40 40 40
use VIA1  VIA1_7
array 0 1 180 0 4 180
timestamp 1569139307
transform 1 0 11625 0 1 8455
box -40 -40 40 40
use VIA1  VIA1_8
array 0 0 0 0 4 160
timestamp 1569139307
transform 1 0 225 0 1 9990
box -40 -40 40 40
use VIA1  VIA1_9
array 0 4 180 0 4 180
timestamp 1569139307
transform 1 0 7825 0 1 19735
box -40 -40 40 40
use VIA1  VIA1_10
array 0 0 0 0 1 160
timestamp 1569139307
transform 1 0 8111 0 1 21818
box -40 -40 40 40
use via1_array_CDNS_704676826051  via1_array_CDNS_704676826051_0
array 0 2 200 0 0 0
timestamp 1569139307
transform 1 0 8010 0 1 23752
box 0 0 200 200
use via1_CDNS_704676826054  via1_CDNS_704676826054_0
timestamp 1569139307
transform 1 0 5410 0 1 20800
box 0 0 200 200
use via1_CDNS_704676826054  via1_CDNS_704676826054_1
timestamp 1569139307
transform 1 0 5210 0 1 20800
box 0 0 200 200
use VIA2  VIA2_0
array 0 1 160 0 0 0
timestamp 1569139307
transform 1 0 7565 0 1 23735
box -40 -40 40 40
<< end >>
