** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-1_Inverter_XSchem/inverter_top.sch
**.subckt inverter_top A Y
*.ipin A
*.opin Y
X1 A Y VDD GND inverter
**.ends

* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-1_Inverter_XSchem/inverter.sym # of pins=4
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-1_Inverter_XSchem/inverter.sym
** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-1_Inverter_XSchem/inverter.sch
.subckt inverter A Y VP VN
*.ipin A
*.opin Y
*.iopin VP
*.iopin VN
M1 Y A VN VN nfet w=5u l=0.18u m=1
M2 Y A VP VP pfet w=5u l=0.18u m=1
.ends

.GLOBAL GND
.GLOBAL VDD
.end
