magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -140 -1950 2539 5180
<< metal2 >>
rect 433 5032 977 5060
rect 1076 5032 2020 5060
use DOUBLE_GUARD  DOUBLE_GUARD_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 0 0 1 1660
box -20 -20 2419 500
use METAL_RING  METAL_RING_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 0 0 1 0
box 0 0 2400 5012
use ndiode10_CDNS_7046768260510  ndiode10_CDNS_7046768260510_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
array 0 3 480 0 2 480
timestamp 1537935238
transform 1 0 230 0 1 51
box 20 20 480 480
use PAD_80  PAD_80_0
timestamp 1537935238
transform 1 0 1200 0 1 -980
box -850 -850 850 980
use PAD_METAL_ANA  PAD_METAL_ANA_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
timestamp 1537935238
transform 1 0 0 0 1 0
box 62 0 2337 5060
use pdiode10_CDNS_7046768260513  pdiode10_CDNS_7046768260513_0 ~/ETRI050_DesignKit/pads_ETRI050/GDS_Magic
array 0 3 480 0 2 480
timestamp 1537935238
transform 1 0 210 0 1 2314
box 0 0 540 540
<< labels >>
flabel space 1200 -980 1200 -980 0 FreeSans 1000 0 0 0 PAD
flabel m3p s 0 3061 0 3061 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 0 4358 0 4358 0 FreeSans 1000 0 0 0 VDD
flabel m3p s 1 4821 1 4821 0 FreeSans 1000 0 0 0 VSS
flabel m3p s 0 717 0 717 0 FreeSans 1000 0 0 0 VSS
flabel m2p s 744 5060 744 5060 0 FreeSans 400 0 0 0 PADR
flabel m2p s 1547 5060 1547 5060 0 FreeSans 400 0 0 0 PAD
<< end >>
