magic
tech scmos
magscale 1 2
timestamp 1727487319
<< nwell >>
rect -6 154 106 273
<< ntransistor >>
rect 20 14 24 54
rect 30 14 34 54
rect 50 14 54 54
<< ptransistor >>
rect 20 206 24 246
rect 40 206 44 246
rect 62 166 66 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 30 54
rect 34 14 36 54
rect 48 14 50 54
rect 54 14 56 54
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 40 246
rect 44 206 48 246
rect 60 166 62 246
rect 66 166 68 246
<< ndcontact >>
rect 6 14 18 54
rect 36 14 48 54
rect 56 14 68 54
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 48 166 60 246
rect 68 166 80 246
<< psubstratepcontact >>
rect 0 -6 100 6
<< nsubstratencontact >>
rect 0 254 100 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 62 246 66 250
rect 20 202 24 206
rect 40 202 44 206
rect 12 198 24 202
rect 30 198 44 202
rect 12 103 16 198
rect 12 72 16 91
rect 30 129 34 198
rect 62 161 66 166
rect 62 155 68 161
rect 30 117 44 129
rect 12 61 24 72
rect 20 54 24 61
rect 30 54 34 117
rect 64 72 68 155
rect 56 60 68 72
rect 50 54 54 60
rect 20 10 24 14
rect 30 10 34 14
rect 50 10 54 14
<< polycontact >>
rect 4 91 16 103
rect 44 117 56 129
rect 44 60 56 72
<< metal1 >>
rect 0 266 100 268
rect 0 252 100 254
rect 6 246 18 252
rect 48 246 60 252
rect 26 72 32 206
rect 68 117 74 166
rect 6 66 44 72
rect 6 54 18 66
rect 68 42 74 103
rect 36 8 48 14
rect 0 6 100 8
rect 0 -8 100 -6
<< m2contact >>
rect 3 103 17 117
rect 43 103 57 117
rect 63 103 77 117
<< metal2 >>
rect 3 117 17 137
rect 63 117 77 137
rect 43 83 57 103
<< m2p >>
rect 3 123 17 137
rect 63 123 77 137
rect 43 83 57 97
<< labels >>
rlabel metal2 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal2 43 83 57 97 0 B
port 1 nsew signal input
rlabel metal1 0 252 100 254 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 -8 100 -6 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal2 63 123 77 137 0 Y
port 2 nsew signal output
rlabel metal1 0 254 100 266 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 266 100 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 6 100 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -6 100 6 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
