magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -60 -60 78 152
<< polysilicon >>
rect 1 88 17 91
rect 1 4 3 88
rect 15 4 17 88
rect 1 1 17 4
<< polycontact >>
rect 3 4 15 88
<< metal1 >>
rect 0 88 18 92
rect 0 4 3 88
rect 15 4 18 88
rect 0 0 18 4
<< end >>
