magic
tech scmos
magscale 1 3
timestamp 1725342160
<< nwell >>
rect 110 110 300 300
<< diffusion >>
rect 76 346 334 364
rect 46 76 64 334
rect 151 261 259 279
rect 131 151 149 259
rect 196 196 214 214
rect 261 151 279 259
rect 151 131 259 149
rect 346 76 364 334
rect 76 46 334 64
<< pdiffusion >>
rect 195 214 215 215
rect 195 196 196 214
rect 214 196 215 214
rect 195 195 215 196
<< psubstratepdiff >>
rect 45 364 365 365
rect 45 346 76 364
rect 334 346 365 364
rect 45 345 365 346
rect 45 334 65 345
rect 45 76 46 334
rect 64 76 65 334
rect 345 334 365 345
rect 45 65 65 76
rect 345 76 346 334
rect 364 76 365 334
rect 345 65 365 76
rect 45 64 365 65
rect 45 46 76 64
rect 334 46 365 64
rect 45 45 365 46
<< nsubstratendiff >>
rect 130 279 280 280
rect 130 261 151 279
rect 259 261 280 279
rect 130 260 280 261
rect 130 259 150 260
rect 130 151 131 259
rect 149 151 150 259
rect 260 259 280 260
rect 130 150 150 151
rect 260 151 261 259
rect 279 151 280 259
rect 260 150 280 151
rect 130 149 280 150
rect 130 131 151 149
rect 259 131 280 149
rect 130 130 280 131
<< metal1 >>
rect 45 345 365 365
rect 45 65 65 345
rect 130 260 280 280
rect 130 150 150 260
rect 195 195 215 215
rect 260 150 280 260
rect 130 130 280 150
rect 345 65 365 345
rect 45 45 365 65
<< end >>
