* NGSPICE file created from fir_pe.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL vdd gnd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for XNOR2X1 abstract view
.subckt XNOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for XOR2X1 abstract view
.subckt XOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for INVX8 abstract view
.subckt INVX8 A Y vdd gnd
.ends

.subckt fir_pe gnd vdd Cin[5] Cin[4] Cin[3] Cin[2] Cin[1] Cin[0] Rdy Vld Xin[3] Xin[2]
+ Xin[1] Xin[0] Xout[3] Xout[2] Xout[1] Xout[0] Yin[3] Yin[2] Yin[1] Yin[0] Yout[3]
+ Yout[2] Yout[1] Yout[0] clk
XFILL_1__728_ vdd gnd FILL
XFILL86850x35250 vdd gnd FILL
XFILL_1__1104_ vdd gnd FILL
XFILL_2__992_ vdd gnd FILL
XFILL_1__1035_ vdd gnd FILL
XFILL_2__1213_ vdd gnd FILL
XFILL_0__815_ vdd gnd FILL
XFILL_2__1075_ vdd gnd FILL
XFILL_2__1144_ vdd gnd FILL
XFILL_0__746_ vdd gnd FILL
X_1270_ _1270_/A _1270_/B _1275_/C vdd gnd NAND2X1
XFILL_3__1253_ vdd gnd FILL
X_1468_ _804_/Y _1503_/CLK _802_/A vdd gnd DFFPOSX1
X_1399_ _738_/B _813_/A _1399_/C _1399_/D _1500_/D vdd gnd OAI22X1
XFILL_2__975_ vdd gnd FILL
XFILL_1__1018_ vdd gnd FILL
X_981_ _985_/A _985_/B _984_/A _982_/C vdd gnd OAI21X1
XFILL_3__742_ vdd gnd FILL
XFILL_0__1260_ vdd gnd FILL
XFILL_0__1191_ vdd gnd FILL
XFILL_2__1127_ vdd gnd FILL
XFILL_2__1058_ vdd gnd FILL
XFILL_0__729_ vdd gnd FILL
X_1253_ _1257_/B _1254_/A vdd gnd INVX1
X_1322_ _1322_/A _1329_/A _1324_/B vdd gnd XNOR2X1
XFILL_1__993_ vdd gnd FILL
X_1184_ _1370_/A _1184_/B _1184_/C _1481_/D vdd gnd OAI21X1
XFILL_0__1527_ vdd gnd FILL
XFILL_0__1389_ vdd gnd FILL
XFILL_2__760_ vdd gnd FILL
XFILL_2__958_ vdd gnd FILL
XFILL_2__889_ vdd gnd FILL
X_895_ _933_/D _895_/B _895_/C _904_/B vdd gnd OAI21X1
X_964_ _969_/D _969_/C _965_/A vdd gnd NAND2X1
XFILL_0__1243_ vdd gnd FILL
XFILL_0__1312_ vdd gnd FILL
XFILL_0__1174_ vdd gnd FILL
X_1236_ _1236_/A _1236_/B _1483_/D vdd gnd NAND2X1
X_1305_ _1307_/A _1306_/A _1309_/A vdd gnd NOR2X1
XFILL_1__976_ vdd gnd FILL
XFILL_1__1352_ vdd gnd FILL
XFILL_1__1421_ vdd gnd FILL
XBUFX2_insert0 _1526_/Q _786_/A vdd gnd BUFX2
XFILL_1__1283_ vdd gnd FILL
X_1098_ _1212_/B _1098_/B _1099_/B vdd gnd NAND2X1
X_1167_ _1202_/B _1173_/B _1174_/C _1192_/A vdd gnd NAND3X1
XFILL_2__743_ vdd gnd FILL
XFILL_2__812_ vdd gnd FILL
XFILL_2__1392_ vdd gnd FILL
XFILL_2__1530_ vdd gnd FILL
XFILL_0__994_ vdd gnd FILL
XFILL_1__761_ vdd gnd FILL
X_947_ _947_/A _947_/B _947_/C _952_/A vdd gnd AOI21X1
XFILL_1__830_ vdd gnd FILL
X_878_ _878_/A _915_/C vdd gnd INVX1
X_1021_ _974_/A _1089_/C _1036_/B _1025_/A vdd gnd NAND3X1
XFILL_0__1226_ vdd gnd FILL
XFILL_0__1157_ vdd gnd FILL
XFILL_0__1088_ vdd gnd FILL
XFILL_1__1404_ vdd gnd FILL
X_1219_ _1356_/B _812_/A _1219_/C _1482_/D vdd gnd OAI21X1
XFILL_1__959_ vdd gnd FILL
XFILL_1__1335_ vdd gnd FILL
XFILL_1__1266_ vdd gnd FILL
XFILL_2__726_ vdd gnd FILL
XFILL_1__1197_ vdd gnd FILL
X_732_ _732_/A _733_/B vdd gnd INVX1
X_801_ _807_/A _801_/B _801_/C _801_/Y vdd gnd OAI21X1
XFILL_2__1375_ vdd gnd FILL
XFILL_2__1444_ vdd gnd FILL
XFILL_0__1011_ vdd gnd FILL
XFILL_0__977_ vdd gnd FILL
XFILL_1__813_ vdd gnd FILL
XFILL_1__744_ vdd gnd FILL
XFILL87150x70350 vdd gnd FILL
XFILL87150x4050 vdd gnd FILL
X_1004_ _990_/A Cin[2] _998_/Y _999_/Y _1010_/B vdd gnd AOI22X1
XFILL_1__1120_ vdd gnd FILL
XFILL_0__1209_ vdd gnd FILL
XFILL_1__1051_ vdd gnd FILL
XFILL_2__1160_ vdd gnd FILL
XFILL_1__1249_ vdd gnd FILL
XFILL_0__762_ vdd gnd FILL
XFILL_1__1318_ vdd gnd FILL
XFILL_2__1091_ vdd gnd FILL
XFILL_0__900_ vdd gnd FILL
XFILL_0__831_ vdd gnd FILL
XFILL_2__1358_ vdd gnd FILL
XFILL_2__1289_ vdd gnd FILL
XFILL_2__1427_ vdd gnd FILL
X_1484_ _1484_/D _1503_/CLK _1484_/Q vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert25 vdd gnd FILL
XFILL_1__727_ vdd gnd FILL
XFILL_1__1034_ vdd gnd FILL
XFILL_1__1103_ vdd gnd FILL
XFILL_2__991_ vdd gnd FILL
XFILL_1_BUFX2_insert0 vdd gnd FILL
XFILL_2__1143_ vdd gnd FILL
XFILL_2__1212_ vdd gnd FILL
XFILL_0__745_ vdd gnd FILL
XFILL_0_CLKBUF1_insert7 vdd gnd FILL
XFILL_0__814_ vdd gnd FILL
XFILL_2__1074_ vdd gnd FILL
XFILL_3__1321_ vdd gnd FILL
X_1398_ _810_/B _1402_/B _813_/A _1399_/C vdd gnd OAI21X1
X_1467_ _801_/Y _1503_/CLK _799_/A vdd gnd DFFPOSX1
XFILL_1__1017_ vdd gnd FILL
XFILL_2__974_ vdd gnd FILL
XFILL_3__810_ vdd gnd FILL
XFILL85950x11850 vdd gnd FILL
X_980_ _980_/A Cin[4] _984_/A vdd gnd AND2X2
XFILL85650x46950 vdd gnd FILL
XFILL_0__1190_ vdd gnd FILL
XFILL_2__1126_ vdd gnd FILL
XFILL_0__728_ vdd gnd FILL
XFILL_2__1057_ vdd gnd FILL
X_1252_ _1252_/A _1252_/B _1252_/C _1254_/B vdd gnd AOI21X1
X_1321_ _1328_/B _1321_/B _1329_/A vdd gnd NOR2X1
XFILL_3__939_ vdd gnd FILL
XFILL_1__992_ vdd gnd FILL
X_1183_ _1481_/Q _1391_/B _1184_/C vdd gnd NAND2X1
XFILL_0__1388_ vdd gnd FILL
X_1519_ _1519_/D _1521_/CLK _977_/A vdd gnd DFFPOSX1
XFILL_2__957_ vdd gnd FILL
XFILL_2__888_ vdd gnd FILL
XFILL85950x23550 vdd gnd FILL
X_894_ _933_/C _894_/B _894_/C _904_/A vdd gnd NAND3X1
X_963_ _969_/A _969_/B _965_/B vdd gnd NAND2X1
XFILL_0__1311_ vdd gnd FILL
XFILL_0__1242_ vdd gnd FILL
XFILL_2__1109_ vdd gnd FILL
XFILL_0__1173_ vdd gnd FILL
XFILL_1__1420_ vdd gnd FILL
X_1304_ _1304_/A _1326_/C _1307_/A vdd gnd AND2X2
X_1235_ _807_/A _1235_/B _1235_/C _1236_/B vdd gnd NAND3X1
XBUFX2_insert1 _1526_/Q _807_/A vdd gnd BUFX2
XFILL_1__975_ vdd gnd FILL
X_1166_ _1193_/C _1169_/C _1169_/A _1202_/B vdd gnd NAND3X1
X_1097_ _1480_/Q _1391_/B _1147_/C vdd gnd NAND2X1
XFILL_2__811_ vdd gnd FILL
XFILL_1__1351_ vdd gnd FILL
XFILL_1__1282_ vdd gnd FILL
XFILL_2__742_ vdd gnd FILL
XFILL_2__1391_ vdd gnd FILL
XFILL_0__993_ vdd gnd FILL
XFILL_1__760_ vdd gnd FILL
X_877_ _877_/A _917_/A vdd gnd INVX1
X_1020_ _1020_/A _1020_/B _976_/Y _1036_/B vdd gnd OAI21X1
X_946_ _946_/A _989_/B _989_/A _952_/B vdd gnd AOI21X1
XFILL_3__1003_ vdd gnd FILL
XFILL_0__1225_ vdd gnd FILL
XFILL_0__1156_ vdd gnd FILL
XFILL_0__1087_ vdd gnd FILL
XFILL_1__1403_ vdd gnd FILL
X_1218_ _812_/A _1218_/B _1232_/C _1219_/C vdd gnd NAND3X1
X_1149_ _1191_/A _1214_/B _1149_/C _1182_/A vdd gnd AOI21X1
XFILL_1__958_ vdd gnd FILL
XFILL_1__889_ vdd gnd FILL
XFILL_1__1334_ vdd gnd FILL
XFILL_1__1265_ vdd gnd FILL
XFILL_1__1196_ vdd gnd FILL
XFILL_2__725_ vdd gnd FILL
X_731_ _743_/C _741_/A vdd gnd INVX1
X_800_ _812_/A _800_/B _801_/C vdd gnd NAND2X1
XFILL_2__1374_ vdd gnd FILL
XFILL_2__1443_ vdd gnd FILL
XFILL_0__976_ vdd gnd FILL
XFILL_0__1010_ vdd gnd FILL
XFILL_1__743_ vdd gnd FILL
XFILL_1__812_ vdd gnd FILL
X_1003_ _947_/C _1003_/B _946_/A _1078_/C vdd gnd OAI21X1
X_929_ _929_/A _929_/B _931_/C vdd gnd NAND2X1
XFILL_1__1050_ vdd gnd FILL
XFILL_0__1208_ vdd gnd FILL
XFILL_0__1139_ vdd gnd FILL
XFILL_1__1317_ vdd gnd FILL
XFILL_1__1248_ vdd gnd FILL
XFILL_0__761_ vdd gnd FILL
XFILL_1__1179_ vdd gnd FILL
XFILL_2__1090_ vdd gnd FILL
XFILL_0__830_ vdd gnd FILL
XFILL_2__1426_ vdd gnd FILL
XFILL_2__1288_ vdd gnd FILL
XFILL_2__1357_ vdd gnd FILL
XFILL_2_BUFX2_insert26 vdd gnd FILL
XFILL_0__959_ vdd gnd FILL
XFILL_2_BUFX2_insert15 vdd gnd FILL
X_1483_ _1483_/D _1503_/CLK _1483_/Q vdd gnd DFFPOSX1
XFILL_1__726_ vdd gnd FILL
XFILL_3__1397_ vdd gnd FILL
XFILL_2__990_ vdd gnd FILL
XFILL_1__1033_ vdd gnd FILL
XFILL_1__1102_ vdd gnd FILL
XFILL_1_BUFX2_insert1 vdd gnd FILL
XFILL_2__1211_ vdd gnd FILL
XFILL_2__1073_ vdd gnd FILL
XFILL_2__1142_ vdd gnd FILL
XFILL_0__813_ vdd gnd FILL
XFILL_0_CLKBUF1_insert8 vdd gnd FILL
XFILL_0__744_ vdd gnd FILL
XFILL_3__886_ vdd gnd FILL
XFILL_2__1409_ vdd gnd FILL
X_1535_ _745_/Y Yout[3] vdd gnd BUFX2
X_1397_ _808_/A _1401_/C _1399_/D vdd gnd NOR2X1
X_1466_ _798_/Y _1503_/CLK _796_/A vdd gnd DFFPOSX1
XFILL_2__973_ vdd gnd FILL
XFILL_1__1016_ vdd gnd FILL
XFILL_2__1056_ vdd gnd FILL
XFILL_2__1125_ vdd gnd FILL
XFILL_0__727_ vdd gnd FILL
X_1320_ _1328_/C _1321_/B vdd gnd INVX1
X_1251_ _1251_/A _1251_/B _1251_/C _1252_/C vdd gnd OAI21X1
X_1182_ _1182_/A _1214_/C _1184_/B vdd gnd XOR2X1
XFILL_1__991_ vdd gnd FILL
XFILL_0__1387_ vdd gnd FILL
X_1518_ _1518_/D _1523_/CLK _922_/A vdd gnd DFFPOSX1
X_1449_ _751_/A _979_/A _1449_/C _1520_/D vdd gnd OAI21X1
XFILL_2__887_ vdd gnd FILL
XFILL_2__956_ vdd gnd FILL
X_962_ _971_/A _971_/C _962_/C _969_/B vdd gnd NAND3X1
X_893_ _893_/A _893_/B _893_/C _904_/C vdd gnd AOI21X1
XFILL_0__1310_ vdd gnd FILL
XFILL_0__1241_ vdd gnd FILL
XFILL_2__1039_ vdd gnd FILL
XFILL_2__1108_ vdd gnd FILL
XFILL_0__1172_ vdd gnd FILL
X_1303_ _781_/A _966_/A _1326_/C vdd gnd NAND2X1
XFILL_1__974_ vdd gnd FILL
XFILL_1__1350_ vdd gnd FILL
X_1234_ _1241_/B _1234_/B _1235_/B vdd gnd NAND2X1
XBUFX2_insert2 _1526_/Q _815_/C vdd gnd BUFX2
X_1096_ _843_/B _1096_/B _1096_/C _1479_/D vdd gnd OAI21X1
X_1165_ _1165_/A _998_/B _1169_/C vdd gnd NOR2X1
XFILL_2__741_ vdd gnd FILL
XFILL_0__1439_ vdd gnd FILL
XFILL_2__810_ vdd gnd FILL
XFILL_1__1281_ vdd gnd FILL
XFILL_3__1079_ vdd gnd FILL
XFILL_2__1390_ vdd gnd FILL
XFILL_2__939_ vdd gnd FILL
XFILL_0__992_ vdd gnd FILL
X_945_ _951_/B _951_/C _952_/C _957_/B vdd gnd NAND3X1
X_876_ _876_/A _917_/B _876_/C _876_/D _876_/Y vdd gnd OAI22X1
XFILL_0__1224_ vdd gnd FILL
XFILL_0__1155_ vdd gnd FILL
XFILL_0__1086_ vdd gnd FILL
XFILL_1__957_ vdd gnd FILL
XFILL_1__1402_ vdd gnd FILL
X_1217_ _1217_/A _1252_/A _1217_/C _1232_/C vdd gnd OAI21X1
XFILL_1__1333_ vdd gnd FILL
X_1148_ _1214_/A _1149_/C vdd gnd INVX1
X_1079_ _987_/Y _1079_/B _1079_/C _1101_/C vdd gnd OAI21X1
XFILL_1__888_ vdd gnd FILL
XFILL_2__724_ vdd gnd FILL
XFILL_1__1264_ vdd gnd FILL
XFILL_1__1195_ vdd gnd FILL
X_730_ _730_/A _730_/B _730_/C _730_/Y vdd gnd OAI21X1
XFILL_2__1442_ vdd gnd FILL
XFILL_2__1373_ vdd gnd FILL
XFILL_0__975_ vdd gnd FILL
XFILL_1__811_ vdd gnd FILL
X_928_ _928_/A _931_/B vdd gnd INVX1
XFILL_1__742_ vdd gnd FILL
X_1002_ _990_/A _994_/B _994_/A _941_/B _1003_/B vdd gnd AOI22X1
X_859_ _859_/A _859_/B _859_/C _879_/C vdd gnd OAI21X1
XFILL_0__1207_ vdd gnd FILL
XFILL_0__1138_ vdd gnd FILL
XFILL_0__1069_ vdd gnd FILL
XFILL_1__1316_ vdd gnd FILL
XFILL_1__1247_ vdd gnd FILL
XFILL_0__760_ vdd gnd FILL
XFILL_1__1178_ vdd gnd FILL
XFILL_2__1356_ vdd gnd FILL
XFILL_2__1425_ vdd gnd FILL
XFILL_2__1287_ vdd gnd FILL
XFILL_0__958_ vdd gnd FILL
X_1482_ _1482_/D _1503_/CLK _1482_/Q vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert27 vdd gnd FILL
XFILL_0__889_ vdd gnd FILL
XFILL_2_BUFX2_insert16 vdd gnd FILL
XFILL_1__725_ vdd gnd FILL
XFILL_1__1101_ vdd gnd FILL
XFILL_1__1032_ vdd gnd FILL
XFILL_1_BUFX2_insert2 vdd gnd FILL
XFILL_2__1210_ vdd gnd FILL
XFILL_0__812_ vdd gnd FILL
XFILL_2__1141_ vdd gnd FILL
XFILL_2__1072_ vdd gnd FILL
XFILL_0_CLKBUF1_insert9 vdd gnd FILL
XFILL_0__743_ vdd gnd FILL
XFILL_3__954_ vdd gnd FILL
XFILL_2__1339_ vdd gnd FILL
XFILL_2__1408_ vdd gnd FILL
X_1534_ _741_/Y Yout[2] vdd gnd BUFX2
X_1465_ _795_/Y _1525_/CLK _793_/A vdd gnd DFFPOSX1
X_1396_ _1402_/B _1401_/C vdd gnd INVX1
XFILL_2__972_ vdd gnd FILL
XFILL_1__1015_ vdd gnd FILL
XFILL_2__1055_ vdd gnd FILL
XFILL_2__1124_ vdd gnd FILL
XFILL_0__726_ vdd gnd FILL
XFILL_1__990_ vdd gnd FILL
X_1250_ _1251_/B _1252_/B vdd gnd INVX1
X_1181_ _1189_/A _1188_/A _1214_/C vdd gnd AND2X2
XFILL_0__1386_ vdd gnd FILL
X_1517_ _1517_/D _1521_/CLK _776_/B vdd gnd DFFPOSX1
X_1448_ _757_/A Xin[2] _1449_/C vdd gnd NAND2X1
X_1379_ _1381_/A _1395_/A _1383_/A vdd gnd NOR2X1
XFILL86550x54750 vdd gnd FILL
XFILL_2__955_ vdd gnd FILL
XFILL_2__886_ vdd gnd FILL
X_961_ _961_/A _961_/B _961_/C _962_/C vdd gnd OAI21X1
X_892_ _905_/C _905_/B _905_/A _955_/B vdd gnd AOI21X1
XFILL_0__1240_ vdd gnd FILL
XFILL_2__1038_ vdd gnd FILL
XFILL_2__1107_ vdd gnd FILL
XFILL_0__1171_ vdd gnd FILL
X_1302_ _781_/A _966_/A _1304_/A vdd gnd OR2X2
X_1233_ _1233_/A _1242_/B _1241_/A _1234_/B vdd gnd OAI21X1
XFILL_1__973_ vdd gnd FILL
XBUFX2_insert3 _1526_/Q _817_/A vdd gnd BUFX2
XFILL_1__1280_ vdd gnd FILL
X_1095_ _1479_/Q _843_/B _1096_/C vdd gnd NAND2X1
X_1164_ _998_/B _1165_/A _1164_/C _1173_/B vdd gnd OAI21X1
XFILL_3__1147_ vdd gnd FILL
XFILL_0__1438_ vdd gnd FILL
XFILL_0__1369_ vdd gnd FILL
XFILL_2__740_ vdd gnd FILL
XFILL86550x66450 vdd gnd FILL
XFILL_0__991_ vdd gnd FILL
XFILL_2__938_ vdd gnd FILL
XFILL_2__869_ vdd gnd FILL
X_944_ _989_/A _989_/B _946_/A _951_/C vdd gnd NAND3X1
X_875_ _917_/B _878_/A _876_/D vdd gnd NAND2X1
XFILL_0__1223_ vdd gnd FILL
XFILL_0__1154_ vdd gnd FILL
XFILL_0__1085_ vdd gnd FILL
X_1216_ _1233_/A _1217_/C vdd gnd INVX1
XFILL_1__887_ vdd gnd FILL
XFILL_1__956_ vdd gnd FILL
X_1147_ _1404_/A _1147_/B _1147_/C _1480_/D vdd gnd OAI21X1
XFILL_1__1401_ vdd gnd FILL
XFILL_1__1263_ vdd gnd FILL
XFILL_1__1332_ vdd gnd FILL
X_1078_ _1078_/A _995_/Y _1078_/C _1079_/B vdd gnd AOI21X1
XFILL_2__723_ vdd gnd FILL
XFILL86850x43050 vdd gnd FILL
XFILL_1__1194_ vdd gnd FILL
XFILL86550x78150 vdd gnd FILL
XFILL_2__1372_ vdd gnd FILL
XFILL_2__1441_ vdd gnd FILL
XFILL_0__974_ vdd gnd FILL
XFILL_1__741_ vdd gnd FILL
XFILL_1__810_ vdd gnd FILL
X_927_ _928_/A _927_/B _927_/C _950_/A vdd gnd NAND3X1
X_858_ _879_/B _879_/A _871_/C _868_/B vdd gnd NAND3X1
XCLKBUF1_insert10 clk _1521_/CLK vdd gnd CLKBUF1
X_789_ _815_/C _789_/B _789_/C _789_/Y vdd gnd OAI21X1
X_1001_ _995_/Y _1078_/A _989_/Y _1016_/B vdd gnd NAND3X1
XFILL_0__1137_ vdd gnd FILL
XFILL_0__1206_ vdd gnd FILL
XFILL_0__1068_ vdd gnd FILL
XFILL_1__939_ vdd gnd FILL
XFILL_1__1246_ vdd gnd FILL
XFILL_1__1315_ vdd gnd FILL
XFILL_1__1177_ vdd gnd FILL
XFILL_2__1355_ vdd gnd FILL
XFILL_2__1424_ vdd gnd FILL
XFILL_2__1286_ vdd gnd FILL
XFILL_0__957_ vdd gnd FILL
X_1481_ _1481_/D _1526_/CLK _1481_/Q vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert28 vdd gnd FILL
XFILL_0__888_ vdd gnd FILL
XFILL_2_BUFX2_insert17 vdd gnd FILL
XFILL_1__724_ vdd gnd FILL
XFILL_1__1100_ vdd gnd FILL
XFILL_1__1031_ vdd gnd FILL
XFILL_1_BUFX2_insert3 vdd gnd FILL
XFILL_2__1140_ vdd gnd FILL
XFILL_0__811_ vdd gnd FILL
XFILL_0__742_ vdd gnd FILL
XFILL_1__1229_ vdd gnd FILL
XFILL_2__1071_ vdd gnd FILL
XFILL86550x7950 vdd gnd FILL
XFILL_2__1338_ vdd gnd FILL
XFILL_2__1269_ vdd gnd FILL
XFILL_2__1407_ vdd gnd FILL
X_1533_ _736_/Y Yout[1] vdd gnd BUFX2
X_1464_ _792_/Y _1515_/CLK _790_/A vdd gnd DFFPOSX1
X_1395_ _1395_/A _1395_/B _1395_/C _1402_/B vdd gnd AOI21X1
XFILL_2__971_ vdd gnd FILL
XFILL_1__1014_ vdd gnd FILL
XFILL_2__1123_ vdd gnd FILL
XFILL_0__725_ vdd gnd FILL
XFILL_2__1054_ vdd gnd FILL
X_1180_ _1192_/B _1180_/B _1180_/C _1188_/A vdd gnd NAND3X1
XFILL_0__1385_ vdd gnd FILL
XFILL_3__1094_ vdd gnd FILL
X_1516_ _1516_/D _1526_/CLK _773_/B vdd gnd DFFPOSX1
X_1378_ _1384_/C _1378_/B _1381_/A vdd gnd AND2X2
X_1447_ _751_/A _924_/A _1447_/C _1519_/D vdd gnd OAI21X1
XFILL_2__954_ vdd gnd FILL
XFILL_2__885_ vdd gnd FILL
X_960_ _970_/A _970_/B _970_/C _971_/C vdd gnd NAND3X1
X_891_ _933_/D _895_/B _933_/C _905_/C vdd gnd OAI21X1
XFILL_2__1106_ vdd gnd FILL
XFILL_0__1170_ vdd gnd FILL
XFILL_2__1037_ vdd gnd FILL
X_1232_ _1241_/A _1232_/B _1232_/C _1235_/C vdd gnd NAND3X1
X_1301_ _780_/B _917_/A _1301_/C _1306_/A vdd gnd OAI21X1
XFILL_1__972_ vdd gnd FILL
XFILL_0__1437_ vdd gnd FILL
XFILL_3__1215_ vdd gnd FILL
XBUFX2_insert4 _1526_/Q _917_/B vdd gnd BUFX2
X_1094_ _1094_/A _1100_/A _1096_/B vdd gnd XOR2X1
X_1163_ _1193_/C _1169_/A _1164_/C vdd gnd NAND2X1
XFILL_0__1299_ vdd gnd FILL
XFILL_0__1368_ vdd gnd FILL
XFILL_1_BUFX2_insert30 vdd gnd FILL
XFILL_0__990_ vdd gnd FILL
XFILL_2__937_ vdd gnd FILL
XFILL_2__799_ vdd gnd FILL
XFILL_2__868_ vdd gnd FILL
X_943_ _943_/A _999_/B _988_/A _989_/B vdd gnd OAI21X1
X_874_ _874_/A _874_/B _874_/C _878_/A vdd gnd NAND3X1
XFILL_0__1222_ vdd gnd FILL
XFILL_0__1153_ vdd gnd FILL
XFILL_0__1084_ vdd gnd FILL
XFILL_1__1400_ vdd gnd FILL
X_1146_ _1191_/A _1187_/B _1147_/B vdd gnd XOR2X1
X_1215_ _1215_/A _1215_/B _1215_/C _1252_/A vdd gnd AOI21X1
XFILL_1__955_ vdd gnd FILL
XFILL_1__886_ vdd gnd FILL
XFILL_1__1262_ vdd gnd FILL
XFILL_1__1331_ vdd gnd FILL
XFILL_1__1193_ vdd gnd FILL
X_1077_ _1101_/B _1101_/A _1085_/C _1091_/C vdd gnd NAND3X1
XFILL_2__1371_ vdd gnd FILL
XFILL_2__1440_ vdd gnd FILL
XFILL_1__1529_ vdd gnd FILL
XFILL_0__973_ vdd gnd FILL
XFILL_1__740_ vdd gnd FILL
X_788_ _815_/C _788_/B _789_/C vdd gnd NAND2X1
X_1000_ _999_/Y _996_/Y _998_/Y _1078_/A vdd gnd NAND3X1
X_857_ _893_/A _893_/B _881_/C _879_/B vdd gnd NAND3X1
X_926_ _979_/A _985_/B _929_/A _927_/C vdd gnd OAI21X1
XCLKBUF1_insert11 clk _1515_/CLK vdd gnd CLKBUF1
XFILL_0__1136_ vdd gnd FILL
XFILL_0__1205_ vdd gnd FILL
XFILL_0__1067_ vdd gnd FILL
X_1129_ _1129_/A _1129_/B _1129_/C _1130_/B vdd gnd AOI21X1
XFILL_1__938_ vdd gnd FILL
XFILL_1__869_ vdd gnd FILL
XFILL_1__1314_ vdd gnd FILL
XFILL_1__1245_ vdd gnd FILL
XFILL_1__1176_ vdd gnd FILL
XFILL_2__1423_ vdd gnd FILL
XFILL_2__1354_ vdd gnd FILL
XFILL_2__1285_ vdd gnd FILL
XFILL_0__887_ vdd gnd FILL
XFILL_0__956_ vdd gnd FILL
X_1480_ _1480_/D _1508_/CLK _1480_/Q vdd gnd DFFPOSX1
XFILL_3__1532_ vdd gnd FILL
XFILL_2_BUFX2_insert29 vdd gnd FILL
XFILL_2_BUFX2_insert18 vdd gnd FILL
XFILL_1__723_ vdd gnd FILL
X_909_ _909_/A _910_/C vdd gnd INVX1
XFILL_1__1030_ vdd gnd FILL
XFILL_0__1119_ vdd gnd FILL
XFILL_1_BUFX2_insert4 vdd gnd FILL
XFILL_0__741_ vdd gnd FILL
XFILL_0__810_ vdd gnd FILL
XFILL_1__1228_ vdd gnd FILL
XFILL_1__1159_ vdd gnd FILL
XFILL_2__1070_ vdd gnd FILL
XFILL85650x66450 vdd gnd FILL
XFILL_2__1406_ vdd gnd FILL
XFILL_2__1337_ vdd gnd FILL
XFILL_2__1268_ vdd gnd FILL
X_1532_ _730_/Y Yout[0] vdd gnd BUFX2
XFILL_2__1199_ vdd gnd FILL
XFILL_0__939_ vdd gnd FILL
X_1394_ _1394_/A _1394_/B _1395_/B vdd gnd NOR2X1
X_1463_ _789_/Y _1523_/CLK _787_/A vdd gnd DFFPOSX1
XFILL87150x7950 vdd gnd FILL
XFILL_2__970_ vdd gnd FILL
XFILL_1__1013_ vdd gnd FILL
XFILL_2__1053_ vdd gnd FILL
XFILL_2__1122_ vdd gnd FILL
XFILL_0__724_ vdd gnd FILL
XFILL_3__1162_ vdd gnd FILL
XFILL_0__1384_ vdd gnd FILL
X_1515_ _1515_/D _1515_/CLK _770_/B vdd gnd DFFPOSX1
X_1377_ _1392_/B _1384_/C vdd gnd INVX1
X_1446_ _751_/A Xin[1] _1447_/C vdd gnd NAND2X1
XFILL_2__953_ vdd gnd FILL
XFILL_2__884_ vdd gnd FILL
X_890_ _933_/A _988_/A _895_/B vdd gnd NOR2X1
XFILL_2__1105_ vdd gnd FILL
XFILL_2__1036_ vdd gnd FILL
X_1300_ _735_/D _967_/A _1309_/C vdd gnd NAND2X1
X_1231_ _1241_/B _1232_/B vdd gnd INVX1
XFILL_1__971_ vdd gnd FILL
X_1162_ _759_/A _1225_/B _1162_/C _1169_/A vdd gnd OAI21X1
XBUFX2_insert5 _1526_/Q _812_/A vdd gnd BUFX2
XFILL_0__1436_ vdd gnd FILL
X_1093_ _1212_/B _1212_/A _1100_/A vdd gnd NAND2X1
XFILL_0__1367_ vdd gnd FILL
XFILL_0__1298_ vdd gnd FILL
XFILL_1_BUFX2_insert20 vdd gnd FILL
X_1429_ _1437_/B _1435_/B _1429_/C _1510_/D vdd gnd OAI21X1
XFILL_1_BUFX2_insert31 vdd gnd FILL
XFILL_1_CLKBUF1_insert10 vdd gnd FILL
XFILL_2__936_ vdd gnd FILL
XFILL_2__798_ vdd gnd FILL
XFILL_2__867_ vdd gnd FILL
X_942_ _942_/A _998_/A _946_/A vdd gnd NAND2X1
X_873_ _874_/B _874_/C _874_/A _876_/C vdd gnd AOI21X1
XFILL_0__1221_ vdd gnd FILL
XFILL_0__1083_ vdd gnd FILL
XFILL_2__1019_ vdd gnd FILL
XFILL_0__1152_ vdd gnd FILL
XFILL_1__954_ vdd gnd FILL
XFILL_1__1330_ vdd gnd FILL
X_1145_ _1214_/A _1214_/B _1187_/B vdd gnd NAND2X1
X_1214_ _1214_/A _1214_/B _1214_/C _1215_/C vdd gnd NAND3X1
XFILL_1__885_ vdd gnd FILL
XFILL_0__1419_ vdd gnd FILL
XFILL_1__1192_ vdd gnd FILL
XFILL_1__1261_ vdd gnd FILL
X_1076_ _1130_/C _1106_/A _1106_/B _1101_/A vdd gnd NAND3X1
XFILL_2__1370_ vdd gnd FILL
XFILL_1__1528_ vdd gnd FILL
XFILL_0__972_ vdd gnd FILL
XFILL_2__919_ vdd gnd FILL
X_925_ Cin[3] _985_/B vdd gnd INVX2
X_787_ _787_/A _789_/B vdd gnd INVX1
X_856_ _881_/B _893_/B vdd gnd INVX1
XCLKBUF1_insert12 clk _1508_/CLK vdd gnd CLKBUF1
XFILL_0__1204_ vdd gnd FILL
XFILL_0__1135_ vdd gnd FILL
XFILL_0__1066_ vdd gnd FILL
XFILL_1__937_ vdd gnd FILL
XFILL_1__799_ vdd gnd FILL
XFILL_1__1313_ vdd gnd FILL
X_1128_ _1178_/A _1178_/B _1138_/C _1143_/A vdd gnd NAND3X1
X_1059_ _1120_/A _1113_/A vdd gnd INVX1
XFILL_1__868_ vdd gnd FILL
XFILL_1__1244_ vdd gnd FILL
XFILL_1__1175_ vdd gnd FILL
XFILL_2__1422_ vdd gnd FILL
XFILL_2__1353_ vdd gnd FILL
XFILL_2__1284_ vdd gnd FILL
XFILL_0__955_ vdd gnd FILL
XFILL_0__886_ vdd gnd FILL
XFILL_2_BUFX2_insert19 vdd gnd FILL
X_908_ _912_/A _908_/B _908_/C _969_/D vdd gnd NAND3X1
X_839_ _839_/A _874_/A vdd gnd INVX1
XFILL_0__1118_ vdd gnd FILL
XFILL_0__1049_ vdd gnd FILL
XFILL_1_BUFX2_insert5 vdd gnd FILL
XFILL_0__740_ vdd gnd FILL
XFILL_1__1227_ vdd gnd FILL
XFILL_1__1158_ vdd gnd FILL
XFILL_1__1089_ vdd gnd FILL
XFILL_2__1405_ vdd gnd FILL
XFILL_2__1336_ vdd gnd FILL
XFILL_2__1267_ vdd gnd FILL
XFILL_2__1198_ vdd gnd FILL
XFILL_0__938_ vdd gnd FILL
X_1462_ _786_/Y _1523_/CLK _784_/A vdd gnd DFFPOSX1
X_1531_ _757_/Y Xout[3] vdd gnd BUFX2
XFILL_0__869_ vdd gnd FILL
X_1393_ _1393_/A _1395_/C vdd gnd INVX1
XFILL_1__1012_ vdd gnd FILL
XFILL_2__1052_ vdd gnd FILL
XFILL_2__1121_ vdd gnd FILL
XFILL_0__723_ vdd gnd FILL
XFILL_0__1383_ vdd gnd FILL
XFILL_3__1230_ vdd gnd FILL
XFILL_2__1319_ vdd gnd FILL
X_1514_ _1514_/D _1526_/CLK _767_/A vdd gnd DFFPOSX1
X_1445_ _1523_/D _901_/A _1445_/C _1518_/D vdd gnd OAI21X1
X_1376_ _804_/B _1376_/B _1392_/B vdd gnd NOR2X1
XFILL_3__1359_ vdd gnd FILL
XFILL_2__952_ vdd gnd FILL
XFILL_2__883_ vdd gnd FILL
XFILL_2__1104_ vdd gnd FILL
XFILL_2__1035_ vdd gnd FILL
XFILL_1__970_ vdd gnd FILL
XBUFX2_insert6 _1526_/Q _813_/A vdd gnd BUFX2
X_1230_ _1239_/B _1239_/A _1241_/B vdd gnd XOR2X1
X_1161_ _1193_/A _1227_/B _1161_/C _1162_/C vdd gnd OAI21X1
X_1092_ _1092_/A _1092_/B _1092_/C _1212_/B vdd gnd NAND3X1
XFILL_3__848_ vdd gnd FILL
XFILL_0__1366_ vdd gnd FILL
XFILL_0__1435_ vdd gnd FILL
XFILL_0__1297_ vdd gnd FILL
XFILL_1_BUFX2_insert21 vdd gnd FILL
X_1428_ _728_/A _728_/B _779_/B _1429_/C vdd gnd OAI21X1
XFILL_1_BUFX2_insert32 vdd gnd FILL
XFILL_1_CLKBUF1_insert11 vdd gnd FILL
X_1359_ _1374_/B _1362_/A _1361_/B vdd gnd AND2X2
XFILL_2__935_ vdd gnd FILL
XFILL_2__866_ vdd gnd FILL
XFILL_2__797_ vdd gnd FILL
X_941_ _994_/A _941_/B _998_/A vdd gnd AND2X2
X_872_ _919_/B _909_/A _910_/B _874_/C vdd gnd NAND3X1
XFILL_0__1220_ vdd gnd FILL
XFILL_0__1082_ vdd gnd FILL
XFILL_2__1018_ vdd gnd FILL
XFILL_0__1151_ vdd gnd FILL
XFILL87150x150 vdd gnd FILL
X_1213_ _969_/Y _1213_/B _1213_/C _1215_/A vdd gnd NAND3X1
XFILL_1__953_ vdd gnd FILL
XFILL_1__1260_ vdd gnd FILL
X_1075_ _1075_/A _1133_/B _1075_/C _1106_/B vdd gnd OAI21X1
X_1144_ _1144_/A _1144_/B _1144_/C _1214_/B vdd gnd OAI21X1
XFILL_1__884_ vdd gnd FILL
XFILL_0__1349_ vdd gnd FILL
XFILL_0__1418_ vdd gnd FILL
XFILL_1__1191_ vdd gnd FILL
XFILL_1__1389_ vdd gnd FILL
XFILL_1__1527_ vdd gnd FILL
XFILL_0__971_ vdd gnd FILL
XFILL_2__849_ vdd gnd FILL
XFILL_2__918_ vdd gnd FILL
X_924_ _924_/A _979_/B _929_/B _927_/B vdd gnd OAI21X1
X_786_ _786_/A _786_/B _786_/C _786_/Y vdd gnd OAI21X1
X_855_ _865_/C _883_/A _881_/C vdd gnd NAND2X1
XCLKBUF1_insert13 clk _1526_/CLK vdd gnd CLKBUF1
XFILL_0__1203_ vdd gnd FILL
XFILL_0__1134_ vdd gnd FILL
XFILL_0__1065_ vdd gnd FILL
XFILL_1__936_ vdd gnd FILL
XFILL_1__867_ vdd gnd FILL
XFILL_1__798_ vdd gnd FILL
XFILL_1__1243_ vdd gnd FILL
XFILL_1__1312_ vdd gnd FILL
X_1127_ _1168_/B _1168_/A _1152_/C _1178_/B vdd gnd NAND3X1
X_1058_ _1120_/B _1133_/A _1120_/A _1129_/A vdd gnd OAI21X1
XFILL86550x50850 vdd gnd FILL
XFILL_1__1174_ vdd gnd FILL
XFILL_2__1352_ vdd gnd FILL
XFILL_2__1421_ vdd gnd FILL
XFILL_2__1283_ vdd gnd FILL
XFILL_0__954_ vdd gnd FILL
XFILL_0__885_ vdd gnd FILL
X_907_ _921_/B _955_/C _921_/A _912_/A vdd gnd NAND3X1
X_838_ _840_/C _840_/B _840_/A _839_/A vdd gnd NAND3X1
X_769_ _769_/A _771_/B vdd gnd INVX1
XFILL_0__1117_ vdd gnd FILL
XFILL_0__1048_ vdd gnd FILL
XFILL_1_BUFX2_insert6 vdd gnd FILL
XFILL_1__919_ vdd gnd FILL
XFILL_1__1226_ vdd gnd FILL
XFILL_1__1157_ vdd gnd FILL
XFILL_1__1088_ vdd gnd FILL
XFILL_2__1335_ vdd gnd FILL
XFILL_2__1404_ vdd gnd FILL
XFILL_2__1266_ vdd gnd FILL
XFILL_2__1197_ vdd gnd FILL
XFILL_0__937_ vdd gnd FILL
X_1392_ _1392_/A _1392_/B _1392_/C _1393_/A vdd gnd AOI21X1
XFILL_0__799_ vdd gnd FILL
X_1461_ _783_/Y _1525_/CLK _781_/A vdd gnd DFFPOSX1
X_1530_ _754_/Y Xout[2] vdd gnd BUFX2
XFILL_0__868_ vdd gnd FILL
XFILL_1__1011_ vdd gnd FILL
XFILL86550x74250 vdd gnd FILL
XFILL_1__1209_ vdd gnd FILL
XFILL_2__1120_ vdd gnd FILL
XFILL_2__1051_ vdd gnd FILL
XFILL_3__795_ vdd gnd FILL
XFILL_0__1382_ vdd gnd FILL
XFILL_2__1249_ vdd gnd FILL
XFILL_2__1318_ vdd gnd FILL
XFILL_0__1451_ vdd gnd FILL
X_1375_ _804_/B _1376_/B _1378_/B vdd gnd NAND2X1
X_1513_ _1513_/D _1521_/CLK _788_/B vdd gnd DFFPOSX1
X_1444_ _1523_/D Xin[0] _1445_/C vdd gnd NAND2X1
XFILL_3__1427_ vdd gnd FILL
XFILL_2__951_ vdd gnd FILL
XFILL_2__882_ vdd gnd FILL
XFILL_2__1103_ vdd gnd FILL
XFILL_2__1034_ vdd gnd FILL
XFILL_3__916_ vdd gnd FILL
X_1160_ _997_/A Cin[4] _1227_/B vdd gnd NAND2X1
X_1091_ _1102_/A _1091_/B _1091_/C _1092_/C vdd gnd NAND3X1
XFILL_0__1365_ vdd gnd FILL
XFILL_0__1296_ vdd gnd FILL
XFILL_0__1434_ vdd gnd FILL
X_1358_ _1373_/B _1362_/A vdd gnd INVX1
XFILL_1_BUFX2_insert22 vdd gnd FILL
X_1427_ _765_/B _1435_/B vdd gnd INVX1
XFILL_1_BUFX2_insert33 vdd gnd FILL
XFILL_1_CLKBUF1_insert12 vdd gnd FILL
X_1289_ _780_/B _917_/A _1291_/A vdd gnd NAND2X1
XFILL_2__796_ vdd gnd FILL
XFILL_2__934_ vdd gnd FILL
XFILL_2__865_ vdd gnd FILL
X_940_ _947_/C _989_/A vdd gnd INVX1
X_871_ _871_/A _871_/B _871_/C _910_/B vdd gnd OAI21X1
XFILL_0__1150_ vdd gnd FILL
XFILL_0__1081_ vdd gnd FILL
XFILL_2__1017_ vdd gnd FILL
X_1212_ _1212_/A _1212_/B _1213_/B vdd gnd AND2X2
XFILL_1__952_ vdd gnd FILL
XFILL_1__883_ vdd gnd FILL
XFILL_0__1417_ vdd gnd FILL
X_1143_ _1143_/A _1143_/B _1179_/A _1144_/B vdd gnd AOI21X1
X_1074_ _1129_/C _1129_/B _1129_/A _1130_/C vdd gnd NAND3X1
XFILL_0__1348_ vdd gnd FILL
XFILL_0__1279_ vdd gnd FILL
XFILL_1__1190_ vdd gnd FILL
XFILL_1__1388_ vdd gnd FILL
XFILL_0__970_ vdd gnd FILL
XFILL_2__917_ vdd gnd FILL
XFILL_2__779_ vdd gnd FILL
XFILL_2__848_ vdd gnd FILL
X_854_ _978_/A _884_/B _883_/A vdd gnd AND2X2
X_923_ _980_/A Cin[3] _929_/B vdd gnd AND2X2
X_785_ _815_/C _785_/B _786_/C vdd gnd NAND2X1
XCLKBUF1_insert14 clk _1523_/CLK vdd gnd CLKBUF1
XFILL_0__1202_ vdd gnd FILL
XFILL_0__1133_ vdd gnd FILL
XFILL_0__1064_ vdd gnd FILL
XFILL_1__797_ vdd gnd FILL
X_1126_ _1133_/C _1132_/B _1168_/B vdd gnd NAND2X1
XFILL_1__935_ vdd gnd FILL
XFILL_1__866_ vdd gnd FILL
XFILL_1__1311_ vdd gnd FILL
XFILL_1__1242_ vdd gnd FILL
X_1057_ _997_/A _997_/B _755_/A _993_/B _1120_/B vdd gnd AOI22X1
XFILL_3__1109_ vdd gnd FILL
XFILL_1__1173_ vdd gnd FILL
XFILL_2__1420_ vdd gnd FILL
XFILL_2__1351_ vdd gnd FILL
XFILL_2__1282_ vdd gnd FILL
XFILL_1_CLKBUF1_insert7 vdd gnd FILL
XFILL_0__953_ vdd gnd FILL
XFILL_0__884_ vdd gnd FILL
X_768_ _786_/A _768_/B _768_/C _768_/Y vdd gnd OAI21X1
X_906_ _955_/A _921_/B vdd gnd INVX1
X_837_ _847_/B _847_/A _859_/C _840_/B vdd gnd NAND3X1
XFILL_0__1116_ vdd gnd FILL
XFILL_0__1047_ vdd gnd FILL
XFILL86850x46950 vdd gnd FILL
XFILL_1__849_ vdd gnd FILL
X_1109_ _994_/A Cin[4] _1150_/B vdd gnd AND2X2
XFILL_1__918_ vdd gnd FILL
XFILL_1__1225_ vdd gnd FILL
XFILL_1__1156_ vdd gnd FILL
XFILL_1__1087_ vdd gnd FILL
XFILL_2__1334_ vdd gnd FILL
XFILL_2__1403_ vdd gnd FILL
XFILL_2__1265_ vdd gnd FILL
XFILL_2__1196_ vdd gnd FILL
XFILL_0__936_ vdd gnd FILL
XFILL_0__867_ vdd gnd FILL
X_1391_ _733_/B _1391_/B _1391_/C _1391_/D _1499_/D vdd gnd AOI22X1
XFILL_0__798_ vdd gnd FILL
X_1460_ _780_/Y _1522_/CLK _778_/A vdd gnd DFFPOSX1
XFILL_3__1374_ vdd gnd FILL
XFILL_1__1010_ vdd gnd FILL
XFILL86850x58650 vdd gnd FILL
XFILL_1__1208_ vdd gnd FILL
XFILL_1__1139_ vdd gnd FILL
XFILL_2__1050_ vdd gnd FILL
XFILL_3__863_ vdd gnd FILL
XFILL_0__1450_ vdd gnd FILL
XFILL_0__1381_ vdd gnd FILL
XFILL_2__1248_ vdd gnd FILL
XFILL_2__1317_ vdd gnd FILL
X_1512_ _1512_/D _1523_/CLK _785_/B vdd gnd DFFPOSX1
XFILL_2__1179_ vdd gnd FILL
XFILL_0__919_ vdd gnd FILL
X_1374_ _1374_/A _1374_/B _1374_/C _1395_/A vdd gnd OAI21X1
X_1443_ _728_/A _1443_/B _1443_/C _1517_/D vdd gnd AOI21X1
XFILL_2__950_ vdd gnd FILL
XFILL_2__881_ vdd gnd FILL
XFILL_2__1033_ vdd gnd FILL
XFILL_2__1102_ vdd gnd FILL
XFILL_0__1433_ vdd gnd FILL
X_1090_ _1090_/A _1102_/C _1090_/C _1092_/B vdd gnd NAND3X1
XFILL_0__1364_ vdd gnd FILL
XFILL_0__1295_ vdd gnd FILL
X_1288_ _729_/D _1350_/A _1299_/C vdd gnd NAND2X1
X_1357_ _1357_/A _1372_/B _1373_/B vdd gnd NOR2X1
XFILL_1_BUFX2_insert23 vdd gnd FILL
X_1426_ _1443_/B _1426_/B _1426_/C _1509_/D vdd gnd AOI21X1
XFILL_1_CLKBUF1_insert13 vdd gnd FILL
XFILL_2__933_ vdd gnd FILL
XFILL_2__795_ vdd gnd FILL
XFILL_2__864_ vdd gnd FILL
X_870_ _879_/C _879_/B _879_/A _909_/A vdd gnd NAND3X1
XFILL_0__1080_ vdd gnd FILL
XFILL_2__1016_ vdd gnd FILL
X_1211_ _1233_/A _1242_/B _1218_/B vdd gnd NAND2X1
XFILL_1__951_ vdd gnd FILL
X_1142_ _1142_/A _1179_/C _1142_/C _1144_/A vdd gnd AOI21X1
XFILL_1__882_ vdd gnd FILL
X_999_ _999_/A _999_/B _999_/C _999_/Y vdd gnd OAI21X1
XFILL_0__1416_ vdd gnd FILL
X_1073_ _1073_/A _1103_/B _1106_/A vdd gnd AND2X2
XFILL_0__1347_ vdd gnd FILL
XFILL_0__1278_ vdd gnd FILL
XFILL_3__1056_ vdd gnd FILL
X_1409_ Yin[1] _1439_/B vdd gnd INVX1
XFILL_1__1387_ vdd gnd FILL
XFILL_2__916_ vdd gnd FILL
XFILL_2__778_ vdd gnd FILL
XFILL_2__847_ vdd gnd FILL
X_784_ _784_/A _786_/B vdd gnd INVX1
X_853_ _881_/A _893_/A vdd gnd INVX1
X_922_ _922_/A Cin[5] _928_/A vdd gnd NAND2X1
XFILL_0__1201_ vdd gnd FILL
XFILL_0__1063_ vdd gnd FILL
XFILL_0__1132_ vdd gnd FILL
XFILL_1__934_ vdd gnd FILL
XFILL_1__796_ vdd gnd FILL
XFILL_1__1310_ vdd gnd FILL
X_1125_ _1133_/A _1133_/B _1132_/A _1152_/C vdd gnd OAI21X1
XFILL_1__865_ vdd gnd FILL
XFILL_1__1241_ vdd gnd FILL
X_1056_ _994_/C _1195_/A _1133_/A vdd gnd NOR2X1
XFILL_1__1172_ vdd gnd FILL
XFILL_2__1350_ vdd gnd FILL
XFILL_1__1439_ vdd gnd FILL
XFILL_2__1281_ vdd gnd FILL
XFILL_1_CLKBUF1_insert8 vdd gnd FILL
XFILL_0__952_ vdd gnd FILL
XFILL_0__883_ vdd gnd FILL
X_905_ _905_/A _905_/B _905_/C _955_/C vdd gnd NAND3X1
X_767_ _767_/A _815_/C _768_/C vdd gnd NAND2X1
X_836_ _924_/A _862_/B _836_/C _847_/B vdd gnd OAI21X1
XFILL_0__1046_ vdd gnd FILL
XFILL_0__1115_ vdd gnd FILL
XFILL_1__917_ vdd gnd FILL
XFILL_1__779_ vdd gnd FILL
X_1039_ _1079_/C _1040_/C vdd gnd INVX1
XFILL_1__848_ vdd gnd FILL
X_1108_ _985_/A _1225_/B _1150_/D vdd gnd NOR2X1
XFILL_1__1224_ vdd gnd FILL
XFILL_1__1155_ vdd gnd FILL
XFILL_1__1086_ vdd gnd FILL
XFILL_2__1402_ vdd gnd FILL
XFILL_2__1264_ vdd gnd FILL
XFILL_2__1333_ vdd gnd FILL
XFILL_2__1195_ vdd gnd FILL
XFILL_0__797_ vdd gnd FILL
XFILL_0__935_ vdd gnd FILL
XFILL_0__866_ vdd gnd FILL
X_1390_ _1390_/A _1394_/A _1391_/B _1391_/D vdd gnd AOI21X1
XFILL_3__1442_ vdd gnd FILL
X_819_ _977_/A _835_/B _826_/A vdd gnd NAND2X1
XFILL_0__1029_ vdd gnd FILL
XFILL_1__1138_ vdd gnd FILL
XFILL_1__1069_ vdd gnd FILL
XFILL_1__1207_ vdd gnd FILL
XFILL_3__931_ vdd gnd FILL
XFILL_0__1380_ vdd gnd FILL
XFILL_2__1316_ vdd gnd FILL
XFILL_2__1247_ vdd gnd FILL
XFILL_2__1178_ vdd gnd FILL
X_1511_ _1511_/D _1523_/CLK _782_/B vdd gnd DFFPOSX1
X_1442_ _728_/A _776_/B _1443_/C vdd gnd NOR2X1
XFILL_0__849_ vdd gnd FILL
XFILL_0__918_ vdd gnd FILL
X_1373_ _1373_/A _1373_/B _1374_/A vdd gnd NAND2X1
XFILL_2__880_ vdd gnd FILL
XFILL_2__1032_ vdd gnd FILL
XFILL_2__1101_ vdd gnd FILL
XFILL_0__1363_ vdd gnd FILL
XFILL_0__1432_ vdd gnd FILL
XFILL_0__1294_ vdd gnd FILL
X_1425_ _800_/B _1426_/B _1426_/C vdd gnd NOR2X1
XFILL_1_BUFX2_insert24 vdd gnd FILL
X_1356_ _798_/B _1356_/B _1372_/B vdd gnd NOR2X1
X_1287_ _843_/B _1287_/B _1287_/C _1489_/D vdd gnd OAI21X1
XFILL_1_CLKBUF1_insert14 vdd gnd FILL
XFILL_2__932_ vdd gnd FILL
XFILL_2__863_ vdd gnd FILL
XFILL_2__794_ vdd gnd FILL
XFILL85950x46950 vdd gnd FILL
XFILL_2__1015_ vdd gnd FILL
XFILL_1__950_ vdd gnd FILL
X_1210_ _1241_/A _1241_/C _1233_/A vdd gnd NAND2X1
X_1141_ _1141_/A _1144_/C vdd gnd INVX1
X_1072_ _1130_/A _1081_/B _1081_/A _1101_/B vdd gnd NAND3X1
X_998_ _998_/A _998_/B _998_/Y vdd gnd NAND2X1
XFILL_1__881_ vdd gnd FILL
XFILL_0__1415_ vdd gnd FILL
XFILL_0__1346_ vdd gnd FILL
XFILL_3__1124_ vdd gnd FILL
XFILL_0__1277_ vdd gnd FILL
X_1408_ _1437_/B _1417_/B _1408_/C _1502_/D vdd gnd OAI21X1
X_1339_ _1339_/A _1352_/B vdd gnd INVX1
XFILL_1__1386_ vdd gnd FILL
XFILL_2__915_ vdd gnd FILL
XFILL_2__846_ vdd gnd FILL
XFILL_2__777_ vdd gnd FILL
X_921_ _921_/A _921_/B _921_/C _961_/C vdd gnd AOI21X1
X_783_ _817_/A _783_/B _783_/C _783_/Y vdd gnd OAI21X1
X_852_ _881_/B _893_/C _881_/A _879_/A vdd gnd OAI21X1
XFILL_0__1200_ vdd gnd FILL
XFILL_0__1131_ vdd gnd FILL
XFILL_0__1062_ vdd gnd FILL
XFILL_1__933_ vdd gnd FILL
XFILL_1__795_ vdd gnd FILL
XFILL_1__864_ vdd gnd FILL
X_1055_ _755_/A _997_/B _1195_/A vdd gnd NAND2X1
X_1124_ _1150_/C _1150_/D _1168_/A vdd gnd XOR2X1
XFILL_0__1329_ vdd gnd FILL
XFILL_1__1240_ vdd gnd FILL
XFILL_1__1171_ vdd gnd FILL
XFILL_1__1438_ vdd gnd FILL
XFILL_1__1369_ vdd gnd FILL
XFILL_2__1280_ vdd gnd FILL
XFILL_0__951_ vdd gnd FILL
XFILL_1_CLKBUF1_insert9 vdd gnd FILL
XFILL_0__882_ vdd gnd FILL
XFILL_2__829_ vdd gnd FILL
X_904_ _904_/A _904_/B _904_/C _921_/A vdd gnd NAND3X1
X_766_ _766_/A _768_/B vdd gnd INVX1
X_835_ _980_/A _835_/B _836_/C vdd gnd NAND2X1
XFILL_0__1114_ vdd gnd FILL
XFILL_0__1045_ vdd gnd FILL
XFILL_1__847_ vdd gnd FILL
XFILL_1__916_ vdd gnd FILL
XFILL_1__778_ vdd gnd FILL
XFILL_1__1223_ vdd gnd FILL
X_1038_ _1090_/A _1102_/A vdd gnd INVX1
X_1107_ Cin[5] _1225_/B vdd gnd INVX2
XFILL_1__1085_ vdd gnd FILL
XFILL_1__1154_ vdd gnd FILL
XFILL_2__1401_ vdd gnd FILL
XFILL_2__1332_ vdd gnd FILL
XFILL_2__1263_ vdd gnd FILL
XFILL_2__1194_ vdd gnd FILL
XFILL_0__934_ vdd gnd FILL
XFILL_0__796_ vdd gnd FILL
XFILL_0__865_ vdd gnd FILL
X_818_ _922_/A _834_/A _823_/A vdd gnd NAND2X1
X_749_ _994_/A _943_/A vdd gnd INVX1
XFILL_0__1028_ vdd gnd FILL
XFILL_1__1206_ vdd gnd FILL
XFILL_1__1137_ vdd gnd FILL
XFILL_1__1068_ vdd gnd FILL
XFILL_2__1315_ vdd gnd FILL
XFILL_2__1246_ vdd gnd FILL
XFILL_2__1177_ vdd gnd FILL
XFILL_0__917_ vdd gnd FILL
X_1441_ _728_/A _1441_/B _1441_/C _1516_/D vdd gnd AOI21X1
X_1510_ _1510_/D _1526_/CLK _779_/B vdd gnd DFFPOSX1
XFILL_0__779_ vdd gnd FILL
XFILL_0__848_ vdd gnd FILL
XFILL87150x19650 vdd gnd FILL
X_1372_ _1373_/A _1372_/B _1372_/C _1374_/C vdd gnd AOI21X1
XFILL_2__1031_ vdd gnd FILL
XFILL_2__1100_ vdd gnd FILL
XFILL_0__1362_ vdd gnd FILL
XFILL_0__1431_ vdd gnd FILL
XFILL_0__1293_ vdd gnd FILL
XFILL_2__1229_ vdd gnd FILL
XFILL_3__1140_ vdd gnd FILL
XFILL_3__1071_ vdd gnd FILL
X_1355_ _796_/A _1482_/Q _1357_/A vdd gnd NOR2X1
X_1424_ _1441_/B _1426_/B _1424_/C _1508_/D vdd gnd AOI21X1
XFILL_1_BUFX2_insert25 vdd gnd FILL
X_1286_ _744_/B _843_/B _1287_/C vdd gnd NAND2X1
XFILL_2__793_ vdd gnd FILL
XFILL_2__862_ vdd gnd FILL
XFILL_2__931_ vdd gnd FILL
XFILL_2__1014_ vdd gnd FILL
XFILL_1__880_ vdd gnd FILL
X_997_ _997_/A _997_/B _998_/B vdd gnd AND2X2
X_1140_ _1141_/A _1177_/B _1140_/C _1214_/A vdd gnd NAND3X1
X_1071_ _1075_/A _1133_/B _1129_/C _1081_/A vdd gnd OAI21X1
XFILL_0__1345_ vdd gnd FILL
XFILL_0__1414_ vdd gnd FILL
XFILL_0__1276_ vdd gnd FILL
X_1338_ _1354_/A _1342_/B vdd gnd INVX1
X_1407_ _803_/B _1417_/B _1408_/C vdd gnd NAND2X1
XFILL_1__1385_ vdd gnd FILL
X_1269_ _1271_/B _1271_/A _1270_/B vdd gnd NOR2X1
XFILL_2__776_ vdd gnd FILL
XFILL_2__845_ vdd gnd FILL
XFILL_2__914_ vdd gnd FILL
X_920_ _971_/A _959_/A vdd gnd INVX1
X_851_ _980_/A _938_/B _978_/A _884_/B _881_/B vdd gnd AOI22X1
X_782_ _815_/C _782_/B _783_/C vdd gnd NAND2X1
XFILL_0__1130_ vdd gnd FILL
XFILL_0__1061_ vdd gnd FILL
XFILL_1__932_ vdd gnd FILL
XFILL_1__863_ vdd gnd FILL
XFILL_1__794_ vdd gnd FILL
X_1054_ _994_/A Cin[2] _1120_/A vdd gnd NAND2X1
X_1123_ _1152_/A _1168_/C _1152_/B _1178_/A vdd gnd OAI21X1
XFILL_0__1259_ vdd gnd FILL
XFILL_0__1328_ vdd gnd FILL
XFILL_1__1170_ vdd gnd FILL
XFILL_1__1368_ vdd gnd FILL
XFILL_1__1437_ vdd gnd FILL
XFILL_0__950_ vdd gnd FILL
XFILL_1__1299_ vdd gnd FILL
XFILL_2__759_ vdd gnd FILL
XFILL_0__881_ vdd gnd FILL
XFILL_2__828_ vdd gnd FILL
X_903_ _955_/B _921_/C _955_/A _908_/C vdd gnd OAI21X1
X_834_ _834_/A _862_/B vdd gnd INVX1
X_765_ _765_/A _765_/B _765_/C _765_/Y vdd gnd OAI21X1
XFILL_0__1113_ vdd gnd FILL
XFILL_0__1044_ vdd gnd FILL
XFILL_1__777_ vdd gnd FILL
X_1106_ _1106_/A _1106_/B _1106_/C _1138_/C vdd gnd AOI21X1
XFILL_1__915_ vdd gnd FILL
XFILL_1__846_ vdd gnd FILL
XFILL_1__1222_ vdd gnd FILL
XFILL_1__1153_ vdd gnd FILL
X_1037_ _986_/C _987_/A _1090_/A vdd gnd NAND2X1
XFILL_1__1084_ vdd gnd FILL
XFILL_2__1400_ vdd gnd FILL
XFILL_2__1262_ vdd gnd FILL
XFILL_2__1331_ vdd gnd FILL
XFILL_2__1193_ vdd gnd FILL
XFILL_0__933_ vdd gnd FILL
XFILL_0__864_ vdd gnd FILL
XFILL_0__795_ vdd gnd FILL
X_817_ _817_/A _817_/Y vdd gnd INVX8
XFILL_2__1529_ vdd gnd FILL
X_748_ _751_/A _759_/A _748_/C _748_/Y vdd gnd OAI21X1
XFILL_0__1027_ vdd gnd FILL
XFILL_1__829_ vdd gnd FILL
XFILL_1__1136_ vdd gnd FILL
XFILL_1__1205_ vdd gnd FILL
XFILL_1__1067_ vdd gnd FILL
XFILL_2__1314_ vdd gnd FILL
XFILL_2__1245_ vdd gnd FILL
XFILL_2__1176_ vdd gnd FILL
XFILL_0__847_ vdd gnd FILL
XFILL_0__916_ vdd gnd FILL
X_1371_ _723_/B _1404_/A _1383_/C vdd gnd NAND2X1
X_1440_ _728_/A _773_/B _1441_/C vdd gnd NOR2X1
XFILL_0__778_ vdd gnd FILL
XFILL_2__1030_ vdd gnd FILL
XFILL_1__1119_ vdd gnd FILL
XFILL_0__1430_ vdd gnd FILL
XFILL_0__1361_ vdd gnd FILL
XFILL_0__1292_ vdd gnd FILL
XFILL_2__1228_ vdd gnd FILL
XFILL_2__1159_ vdd gnd FILL
X_1423_ _797_/B _1426_/B _1424_/C vdd gnd NOR2X1
X_1354_ _1354_/A _1354_/B _1354_/C _1374_/B vdd gnd AOI21X1
X_1285_ _1294_/B _1285_/B _1287_/B vdd gnd XOR2X1
XFILL_1_BUFX2_insert26 vdd gnd FILL
XFILL_1_BUFX2_insert15 vdd gnd FILL
XFILL_2__930_ vdd gnd FILL
XFILL_2__792_ vdd gnd FILL
XFILL_3__1268_ vdd gnd FILL
XFILL_2__861_ vdd gnd FILL
XFILL_2__1013_ vdd gnd FILL
X_996_ _996_/A _996_/Y vdd gnd INVX1
XFILL_0__1413_ vdd gnd FILL
X_1070_ _1070_/A _1070_/B _1120_/A _1133_/B vdd gnd AOI21X1
XFILL_3__757_ vdd gnd FILL
XFILL_0__1275_ vdd gnd FILL
XFILL_0__1344_ vdd gnd FILL
X_1337_ _1339_/A _1354_/A _1341_/A vdd gnd NOR2X1
X_1268_ _769_/A _821_/A _1271_/B vdd gnd NOR2X1
X_1406_ _1526_/D _743_/A _743_/C _1417_/B vdd gnd NAND3X1
XFILL_1__1384_ vdd gnd FILL
XFILL86850x54750 vdd gnd FILL
X_1199_ _1223_/A _1224_/C _1199_/C _1223_/D vdd gnd OAI21X1
XFILL_2__913_ vdd gnd FILL
XFILL_2__775_ vdd gnd FILL
XFILL_2__844_ vdd gnd FILL
X_781_ _781_/A _783_/B vdd gnd INVX1
X_850_ _850_/A _933_/A _893_/C vdd gnd NOR2X1
XFILL_0__1060_ vdd gnd FILL
XFILL_1__793_ vdd gnd FILL
X_1122_ _1122_/A _1132_/A _1152_/A vdd gnd NOR2X1
XFILL_1__862_ vdd gnd FILL
XFILL_1__931_ vdd gnd FILL
X_979_ _979_/A _979_/B _984_/B _982_/B vdd gnd OAI21X1
X_1053_ _998_/A _998_/B _999_/Y _996_/Y _1075_/C vdd gnd AOI22X1
XFILL_0__1258_ vdd gnd FILL
XFILL_0__1189_ vdd gnd FILL
XFILL_0__1327_ vdd gnd FILL
XFILL86850x66450 vdd gnd FILL
XFILL_1__1367_ vdd gnd FILL
XFILL_1__1298_ vdd gnd FILL
XFILL_1__1436_ vdd gnd FILL
XFILL_0__880_ vdd gnd FILL
XFILL_2__758_ vdd gnd FILL
XFILL_2__827_ vdd gnd FILL
X_764_ Xin[3] _765_/B _765_/C vdd gnd NAND2X1
X_902_ _902_/A _930_/C _902_/C _955_/A vdd gnd OAI21X1
X_833_ _977_/A _924_/A vdd gnd INVX1
XFILL_0__1112_ vdd gnd FILL
XFILL_0__1043_ vdd gnd FILL
XFILL_1__914_ vdd gnd FILL
XFILL_1__776_ vdd gnd FILL
XFILL_1__845_ vdd gnd FILL
X_1105_ _1130_/C _1106_/C vdd gnd INVX1
XFILL_1__1221_ vdd gnd FILL
X_1036_ _974_/A _1036_/B _1036_/C _1087_/C vdd gnd AOI21X1
XFILL_1__1152_ vdd gnd FILL
XFILL_1__1083_ vdd gnd FILL
XFILL86850x78150 vdd gnd FILL
XFILL_1__1419_ vdd gnd FILL
XFILL_2__1261_ vdd gnd FILL
XFILL_2__1330_ vdd gnd FILL
XFILL_2__1192_ vdd gnd FILL
XFILL_0__932_ vdd gnd FILL
XFILL_0__863_ vdd gnd FILL
XFILL_0__794_ vdd gnd FILL
X_816_ _816_/A _917_/B _816_/C _816_/Y vdd gnd OAI21X1
XFILL_2__1528_ vdd gnd FILL
X_747_ _751_/A _922_/A _748_/C vdd gnd NAND2X1
XFILL_0__1026_ vdd gnd FILL
XFILL_1__759_ vdd gnd FILL
X_1019_ _1088_/B _1088_/C _1088_/A _1089_/C vdd gnd NAND3X1
XFILL_1__828_ vdd gnd FILL
XFILL_1__1204_ vdd gnd FILL
XFILL_1__1135_ vdd gnd FILL
XFILL_1__1066_ vdd gnd FILL
XFILL_2__1313_ vdd gnd FILL
XFILL_2__1244_ vdd gnd FILL
XFILL_2__1175_ vdd gnd FILL
XFILL_0__777_ vdd gnd FILL
XFILL_0__915_ vdd gnd FILL
XFILL_0__846_ vdd gnd FILL
X_1370_ _1370_/A _1370_/B _1370_/C _1497_/D vdd gnd OAI21X1
XFILL_0__1009_ vdd gnd FILL
X_1499_ _1499_/D _1508_/CLK _732_/A vdd gnd DFFPOSX1
XFILL_1__1118_ vdd gnd FILL
XFILL_1__1049_ vdd gnd FILL
XFILL_0__1360_ vdd gnd FILL
XFILL_0__1291_ vdd gnd FILL
XFILL_2__1227_ vdd gnd FILL
XFILL_2__1158_ vdd gnd FILL
X_1422_ _1439_/B _1426_/B _1422_/C _1507_/D vdd gnd AOI21X1
XFILL_2__1089_ vdd gnd FILL
XFILL_0__829_ vdd gnd FILL
X_1353_ _1353_/A _1353_/B _1353_/C _1354_/C vdd gnd OAI21X1
X_1284_ _1294_/A _1293_/A _1285_/B vdd gnd NOR2X1
XFILL_1_BUFX2_insert27 vdd gnd FILL
XFILL_1_BUFX2_insert16 vdd gnd FILL
XFILL_3__1336_ vdd gnd FILL
XFILL_2__860_ vdd gnd FILL
XFILL_2__791_ vdd gnd FILL
XFILL_2__1012_ vdd gnd FILL
XFILL_2__989_ vdd gnd FILL
XBUFX2_insert30 Cin[1] _834_/A vdd gnd BUFX2
X_995_ _996_/A _995_/B _995_/C _995_/Y vdd gnd NAND3X1
XFILL_3__825_ vdd gnd FILL
XFILL_0__1412_ vdd gnd FILL
XFILL_0__1343_ vdd gnd FILL
XFILL_0__1274_ vdd gnd FILL
X_1405_ Yin[0] _1437_/B vdd gnd INVX1
X_1336_ _1336_/A _1353_/A _1339_/A vdd gnd AND2X2
X_1267_ _771_/B _1275_/B _1271_/A vdd gnd NOR2X1
X_1198_ _755_/A Cin[4] _1224_/C vdd gnd NAND2X1
XFILL_1__1383_ vdd gnd FILL
XFILL_2__843_ vdd gnd FILL
XFILL_2__912_ vdd gnd FILL
XFILL_2__774_ vdd gnd FILL
X_780_ _786_/A _780_/B _780_/C _780_/Y vdd gnd OAI21X1
XFILL_1__930_ vdd gnd FILL
XFILL_1__792_ vdd gnd FILL
X_1052_ _1103_/B _1073_/A _1130_/A vdd gnd NAND2X1
X_1121_ _1195_/A _1195_/B _1132_/A vdd gnd XOR2X1
XFILL_1__861_ vdd gnd FILL
X_978_ _978_/A Cin[3] _984_/B vdd gnd AND2X2
XFILL_0__1326_ vdd gnd FILL
XFILL_0__1257_ vdd gnd FILL
XFILL_0__1188_ vdd gnd FILL
XFILL_1__1435_ vdd gnd FILL
X_1319_ _787_/A _1479_/Q _1328_/C vdd gnd NAND2X1
XFILL_1__1366_ vdd gnd FILL
XFILL_1__1297_ vdd gnd FILL
XFILL_2__826_ vdd gnd FILL
X_901_ _901_/A _979_/B _973_/A _902_/C vdd gnd OAI21X1
XFILL_2__757_ vdd gnd FILL
X_763_ _999_/A _765_/B _763_/C _763_/Y vdd gnd OAI21X1
X_832_ _832_/A _865_/C _859_/C vdd gnd NAND2X1
XFILL_0__1111_ vdd gnd FILL
XFILL_0__1042_ vdd gnd FILL
XFILL_1__913_ vdd gnd FILL
XFILL_1__775_ vdd gnd FILL
XFILL_1__844_ vdd gnd FILL
X_1104_ _1142_/C _1179_/A vdd gnd INVX1
X_1035_ _1089_/C _1036_/C vdd gnd INVX1
XFILL_1__1220_ vdd gnd FILL
XFILL_0__1309_ vdd gnd FILL
XFILL_1__1082_ vdd gnd FILL
XFILL_3__1018_ vdd gnd FILL
XFILL_1__1151_ vdd gnd FILL
XFILL_1__1349_ vdd gnd FILL
XFILL_1__1418_ vdd gnd FILL
XFILL_2__1260_ vdd gnd FILL
XFILL_2__1191_ vdd gnd FILL
XFILL_0__931_ vdd gnd FILL
XFILL_2__809_ vdd gnd FILL
XFILL_0__793_ vdd gnd FILL
XFILL_0__862_ vdd gnd FILL
XFILL_2__1527_ vdd gnd FILL
X_815_ _922_/A _835_/B _815_/C _816_/C vdd gnd NAND3X1
X_746_ _990_/A _759_/A vdd gnd INVX2
XFILL_2__1389_ vdd gnd FILL
XFILL_0__1025_ vdd gnd FILL
XFILL_1__827_ vdd gnd FILL
XFILL_1__1203_ vdd gnd FILL
XFILL_1__758_ vdd gnd FILL
X_1018_ _974_/Y _1029_/B _1029_/A _1025_/B vdd gnd NAND3X1
XFILL_1__1134_ vdd gnd FILL
XFILL_1__1065_ vdd gnd FILL
XFILL_2__1312_ vdd gnd FILL
XFILL_2__1243_ vdd gnd FILL
XFILL_0__914_ vdd gnd FILL
XFILL_2__1174_ vdd gnd FILL
XFILL_0__776_ vdd gnd FILL
XFILL_0__845_ vdd gnd FILL
X_729_ _744_/A _729_/B _765_/B _729_/D _730_/C vdd gnd AOI22X1
XFILL_3__1352_ vdd gnd FILL
XFILL_3__1283_ vdd gnd FILL
XFILL_0__1008_ vdd gnd FILL
X_1498_ _1498_/D _1503_/CLK _723_/B vdd gnd DFFPOSX1
XFILL_3_BUFX2_insert3 vdd gnd FILL
XFILL_1__1117_ vdd gnd FILL
XFILL_1__1048_ vdd gnd FILL
XFILL_3__772_ vdd gnd FILL
XFILL_3__841_ vdd gnd FILL
XFILL85950x66450 vdd gnd FILL
XFILL_0__1290_ vdd gnd FILL
XFILL_2__1226_ vdd gnd FILL
XFILL_2__1157_ vdd gnd FILL
XFILL_2__1088_ vdd gnd FILL
X_1421_ _794_/B _1426_/B _1422_/C vdd gnd NOR2X1
XFILL_0__759_ vdd gnd FILL
XFILL_0__828_ vdd gnd FILL
X_1352_ _1352_/A _1352_/B _1354_/B vdd gnd NOR2X1
XFILL_3__1404_ vdd gnd FILL
X_1283_ _777_/B _876_/A _1293_/A vdd gnd NOR2X1
XFILL_1_BUFX2_insert28 vdd gnd FILL
XFILL_1_BUFX2_insert17 vdd gnd FILL
XFILL_2__790_ vdd gnd FILL
XBUFX2_insert20 _817_/Y _967_/A vdd gnd BUFX2
XFILL_2__1011_ vdd gnd FILL
XFILL_2__988_ vdd gnd FILL
XBUFX2_insert31 Cin[1] _997_/B vdd gnd BUFX2
XFILL85950x78150 vdd gnd FILL
X_994_ _994_/A _994_/B _994_/C _995_/C vdd gnd NAND3X1
XFILL_0__1273_ vdd gnd FILL
XFILL_0__1342_ vdd gnd FILL
XFILL_0__1411_ vdd gnd FILL
XFILL_2__1209_ vdd gnd FILL
X_1335_ _790_/A _1480_/Q _1353_/A vdd gnd NAND2X1
X_1404_ _1404_/A _1404_/B _1404_/C _1501_/D vdd gnd OAI21X1
XFILL_1__1382_ vdd gnd FILL
X_1266_ _821_/A _1275_/B vdd gnd INVX1
X_1197_ _765_/A _985_/B _1227_/B _1199_/C vdd gnd OAI21X1
XFILL_1__1451_ vdd gnd FILL
XFILL_2__773_ vdd gnd FILL
XFILL_2__842_ vdd gnd FILL
XFILL_2__911_ vdd gnd FILL
XFILL_1__860_ vdd gnd FILL
X_977_ _977_/A Cin[5] _983_/A vdd gnd NAND2X1
XFILL_1__791_ vdd gnd FILL
X_1120_ _1120_/A _1120_/B _1120_/C _1122_/A vdd gnd OAI21X1
XFILL87150x15750 vdd gnd FILL
X_1051_ _1051_/A _1051_/B _1103_/A _1103_/B vdd gnd NAND3X1
XFILL_0__1325_ vdd gnd FILL
XFILL_0__1256_ vdd gnd FILL
XFILL_3__1034_ vdd gnd FILL
XFILL_0__1187_ vdd gnd FILL
X_1318_ _787_/A _1479_/Q _1328_/B vdd gnd NOR2X1
XFILL_1__989_ vdd gnd FILL
XFILL_1__1365_ vdd gnd FILL
X_1249_ _1257_/B _1257_/A _1255_/C vdd gnd NOR2X1
XFILL_1__1434_ vdd gnd FILL
XFILL_1__1296_ vdd gnd FILL
XFILL_2__825_ vdd gnd FILL
XFILL_2__756_ vdd gnd FILL
X_900_ _977_/A Cin[3] _973_/A vdd gnd NAND2X1
X_831_ _980_/A _834_/A _865_/C vdd gnd AND2X2
X_762_ Xin[2] _765_/B _763_/C vdd gnd NAND2X1
XFILL_0__1110_ vdd gnd FILL
XFILL_0__1041_ vdd gnd FILL
XFILL_1__843_ vdd gnd FILL
XFILL_1__912_ vdd gnd FILL
XFILL87150x27450 vdd gnd FILL
XFILL_1__774_ vdd gnd FILL
X_1034_ _1034_/A _1034_/B _1100_/B _1094_/A vdd gnd OAI21X1
X_1103_ _1103_/A _1103_/B _1142_/C vdd gnd NAND2X1
XFILL_0__1308_ vdd gnd FILL
XFILL_0__1239_ vdd gnd FILL
XFILL_1__1081_ vdd gnd FILL
XFILL_1__1150_ vdd gnd FILL
XFILL_0_BUFX2_insert30 vdd gnd FILL
XFILL_1__1348_ vdd gnd FILL
XFILL_1__1417_ vdd gnd FILL
XFILL_2__1190_ vdd gnd FILL
XFILL_0__930_ vdd gnd FILL
XFILL_0__792_ vdd gnd FILL
XFILL_2__808_ vdd gnd FILL
XFILL_2__739_ vdd gnd FILL
XFILL_1__1279_ vdd gnd FILL
XFILL_0__861_ vdd gnd FILL
X_814_ _814_/A _816_/A vdd gnd INVX1
X_745_ _745_/A _745_/B _745_/C _745_/Y vdd gnd OAI21X1
XFILL_2__1388_ vdd gnd FILL
XFILL87150x39150 vdd gnd FILL
XFILL_0__1024_ vdd gnd FILL
XFILL_1__826_ vdd gnd FILL
XFILL_1__1202_ vdd gnd FILL
X_1017_ _1020_/A _1020_/B _1088_/C _1029_/B vdd gnd OAI21X1
XFILL_1__757_ vdd gnd FILL
XFILL_1__1064_ vdd gnd FILL
XFILL_1__1133_ vdd gnd FILL
XFILL_2__1311_ vdd gnd FILL
XFILL_2__1242_ vdd gnd FILL
XFILL_0__844_ vdd gnd FILL
XFILL_0__913_ vdd gnd FILL
XFILL_2__1173_ vdd gnd FILL
XFILL_0__775_ vdd gnd FILL
XFILL_3__1420_ vdd gnd FILL
X_728_ _728_/A _728_/B _765_/B vdd gnd NOR2X1
XFILL_0_BUFX2_insert0 vdd gnd FILL
XFILL_0__1007_ vdd gnd FILL
X_1497_ _1497_/D _1526_/CLK _743_/B vdd gnd DFFPOSX1
XFILL_1__809_ vdd gnd FILL
XFILL_1__1116_ vdd gnd FILL
XFILL_1__1047_ vdd gnd FILL
XFILL_2__1225_ vdd gnd FILL
XFILL_2__1156_ vdd gnd FILL
XFILL_2__1087_ vdd gnd FILL
XFILL_0__827_ vdd gnd FILL
X_1420_ _1437_/B _1426_/B _1420_/C _1506_/D vdd gnd AOI21X1
X_1351_ _739_/B _1404_/A _1361_/C vdd gnd NAND2X1
XFILL_1_BUFX2_insert29 vdd gnd FILL
XFILL_0__758_ vdd gnd FILL
XFILL_1_BUFX2_insert18 vdd gnd FILL
X_1282_ _775_/A _845_/A _1294_/A vdd gnd NOR2X1
XFILL_3__969_ vdd gnd FILL
XBUFX2_insert21 _817_/Y _1370_/A vdd gnd BUFX2
XFILL_2__1010_ vdd gnd FILL
XBUFX2_insert32 Cin[1] _994_/B vdd gnd BUFX2
XFILL_2__987_ vdd gnd FILL
X_993_ _997_/A _993_/B _994_/C vdd gnd NAND2X1
XFILL_0__1410_ vdd gnd FILL
XFILL_0__1341_ vdd gnd FILL
XFILL_0__1272_ vdd gnd FILL
XFILL_2__1208_ vdd gnd FILL
XFILL_2__1139_ vdd gnd FILL
X_1334_ _790_/A _1480_/Q _1336_/A vdd gnd OR2X2
X_1403_ _1403_/A _1403_/B _1404_/B vdd gnd NAND2X1
X_1265_ _967_/A _1265_/B _1265_/C _1486_/D vdd gnd OAI21X1
XFILL_1__1381_ vdd gnd FILL
X_1196_ _943_/A _1225_/B _1222_/A vdd gnd NOR2X1
XFILL_1__1450_ vdd gnd FILL
XFILL_2__910_ vdd gnd FILL
XFILL_2__772_ vdd gnd FILL
XFILL_2__841_ vdd gnd FILL
XFILL_2_CLKBUF1_insert7 vdd gnd FILL
XFILL_1__790_ vdd gnd FILL
X_976_ _976_/A _976_/B _976_/C _976_/Y vdd gnd AOI21X1
XFILL_3__1102_ vdd gnd FILL
X_1050_ _985_/A _979_/B _1050_/C _1051_/A vdd gnd OAI21X1
XFILL_0__1255_ vdd gnd FILL
XFILL_0__1324_ vdd gnd FILL
XFILL_0__1186_ vdd gnd FILL
X_1248_ _1258_/A _1248_/B _1257_/B vdd gnd AND2X2
X_1317_ _786_/B _968_/Y _1317_/C _1322_/A vdd gnd OAI21X1
XFILL_1__988_ vdd gnd FILL
XFILL_1__1364_ vdd gnd FILL
XFILL_1__1295_ vdd gnd FILL
XFILL_1__1433_ vdd gnd FILL
X_1179_ _1179_/A _1179_/B _1179_/C _1180_/C vdd gnd OAI21X1
XFILL_2__755_ vdd gnd FILL
XFILL_2__824_ vdd gnd FILL
X_761_ _943_/A _765_/B _761_/C _761_/Y vdd gnd OAI21X1
X_830_ _977_/A _884_/B _832_/A vdd gnd AND2X2
XFILL_0__1040_ vdd gnd FILL
XFILL_1__773_ vdd gnd FILL
XFILL_1__842_ vdd gnd FILL
X_1102_ _1102_/A _1102_/B _1102_/C _1141_/A vdd gnd OAI21X1
X_959_ _959_/A _959_/B _959_/C _969_/A vdd gnd NAND3X1
XFILL_1__911_ vdd gnd FILL
X_1033_ _968_/Y _917_/B _1033_/C _1033_/D _1478_/D vdd gnd OAI22X1
XFILL_0__1307_ vdd gnd FILL
XFILL_0__1238_ vdd gnd FILL
XFILL_1__1080_ vdd gnd FILL
XFILL_0__1169_ vdd gnd FILL
XFILL_0_BUFX2_insert20 vdd gnd FILL
XFILL_0_BUFX2_insert31 vdd gnd FILL
XFILL_1__1347_ vdd gnd FILL
XFILL_1__1278_ vdd gnd FILL
XFILL_1__1416_ vdd gnd FILL
XFILL_0__860_ vdd gnd FILL
XFILL_0__791_ vdd gnd FILL
XFILL_2__807_ vdd gnd FILL
XFILL_2__738_ vdd gnd FILL
X_813_ _813_/A _813_/B _813_/C _813_/Y vdd gnd OAI21X1
X_744_ _744_/A _744_/B _765_/B _744_/D _745_/C vdd gnd AOI22X1
XFILL_2__1387_ vdd gnd FILL
XFILL_0__1023_ vdd gnd FILL
XFILL_0__989_ vdd gnd FILL
XFILL_1__825_ vdd gnd FILL
XFILL_1__756_ vdd gnd FILL
XFILL_1__1201_ vdd gnd FILL
X_1016_ _1016_/A _1016_/B _987_/Y _1020_/B vdd gnd AOI21X1
XFILL_1__1132_ vdd gnd FILL
XFILL86850x50850 vdd gnd FILL
XFILL_1__1063_ vdd gnd FILL
XFILL_2__1310_ vdd gnd FILL
XFILL_2__1241_ vdd gnd FILL
XFILL_0__843_ vdd gnd FILL
XFILL_0__912_ vdd gnd FILL
XFILL_2__1172_ vdd gnd FILL
XFILL_0__774_ vdd gnd FILL
X_727_ _727_/A _728_/B vdd gnd INVX2
XFILL_2__1439_ vdd gnd FILL
XFILL_0_BUFX2_insert1 vdd gnd FILL
XFILL_0__1006_ vdd gnd FILL
X_1496_ _1496_/D _1515_/CLK _739_/B vdd gnd DFFPOSX1
XFILL_1__808_ vdd gnd FILL
XFILL_1__739_ vdd gnd FILL
XFILL_1__1046_ vdd gnd FILL
XFILL_1__1115_ vdd gnd FILL
XFILL_2__1224_ vdd gnd FILL
XFILL_2__1155_ vdd gnd FILL
XFILL_2__1086_ vdd gnd FILL
XFILL_0__826_ vdd gnd FILL
XFILL_0__757_ vdd gnd FILL
X_1350_ _1350_/A _1350_/B _1350_/C _1495_/D vdd gnd OAI21X1
XFILL_1_BUFX2_insert19 vdd gnd FILL
X_1281_ _1281_/A _1281_/B _1281_/C _1294_/B vdd gnd AOI21X1
X_1479_ _1479_/D _1523_/CLK _1479_/Q vdd gnd DFFPOSX1
XFILL86250x27450 vdd gnd FILL
XFILL86850x74250 vdd gnd FILL
XBUFX2_insert22 _817_/Y _1350_/A vdd gnd BUFX2
XFILL_1__1029_ vdd gnd FILL
XBUFX2_insert33 Cin[1] _938_/B vdd gnd BUFX2
XFILL_2__986_ vdd gnd FILL
X_992_ _997_/A _993_/B _999_/C _995_/B vdd gnd NAND3X1
XFILL_0__1340_ vdd gnd FILL
XFILL_0__1271_ vdd gnd FILL
XFILL_2__1138_ vdd gnd FILL
XFILL_2__1207_ vdd gnd FILL
X_1402_ _810_/B _1402_/B _813_/B _1403_/A vdd gnd OAI21X1
XFILL_0__809_ vdd gnd FILL
XFILL_2__1069_ vdd gnd FILL
X_1264_ _729_/B _967_/A _1265_/C vdd gnd NAND2X1
X_1333_ _1333_/A _1333_/B _1354_/A vdd gnd NAND2X1
XFILL_1__1380_ vdd gnd FILL
X_1195_ _1195_/A _1195_/B _1202_/A vdd gnd OR2X2
XFILL_2__771_ vdd gnd FILL
XFILL_2__840_ vdd gnd FILL
XFILL_2_CLKBUF1_insert8 vdd gnd FILL
XFILL_2__969_ vdd gnd FILL
XCLKBUF1_insert7 clk _1522_/CLK vdd gnd CLKBUF1
X_975_ _975_/A _976_/C vdd gnd INVX1
XFILL_0__1323_ vdd gnd FILL
XFILL_0__1185_ vdd gnd FILL
XFILL_0__1254_ vdd gnd FILL
X_1316_ _1316_/A _1316_/B _1316_/C _1492_/D vdd gnd OAI21X1
X_1247_ _1247_/A _1257_/C _1247_/C _1248_/B vdd gnd OAI21X1
XFILL_1__1432_ vdd gnd FILL
X_1178_ _1178_/A _1178_/B _1178_/C _1179_/B vdd gnd AOI21X1
XFILL_1__987_ vdd gnd FILL
XFILL_1__1363_ vdd gnd FILL
XFILL_1__1294_ vdd gnd FILL
XFILL_2__823_ vdd gnd FILL
XFILL_2__754_ vdd gnd FILL
X_760_ Xin[1] _765_/B _761_/C vdd gnd NAND2X1
XFILL_1__910_ vdd gnd FILL
XFILL_1__772_ vdd gnd FILL
X_1032_ _917_/B _1100_/B _1033_/C vdd gnd NAND2X1
X_1101_ _1101_/A _1101_/B _1101_/C _1102_/B vdd gnd AOI21X1
X_958_ _961_/A _961_/B _970_/C _959_/C vdd gnd OAI21X1
X_889_ _990_/A _994_/B _988_/A vdd gnd NAND2X1
XFILL_1__841_ vdd gnd FILL
XFILL_0__1306_ vdd gnd FILL
XFILL_0__1237_ vdd gnd FILL
XFILL_0__1099_ vdd gnd FILL
XFILL_0__1168_ vdd gnd FILL
XFILL_1__1415_ vdd gnd FILL
XFILL_0_BUFX2_insert21 vdd gnd FILL
XFILL_0_BUFX2_insert32 vdd gnd FILL
XFILL_0__790_ vdd gnd FILL
XFILL_2__806_ vdd gnd FILL
XFILL_1__1346_ vdd gnd FILL
XFILL_1__1277_ vdd gnd FILL
XFILL_2__737_ vdd gnd FILL
X_743_ _743_/A _743_/B _743_/C _745_/B vdd gnd OAI21X1
X_812_ _812_/A _812_/B _813_/C vdd gnd NAND2X1
XFILL_2__1386_ vdd gnd FILL
XFILL_0__1022_ vdd gnd FILL
XFILL_0__988_ vdd gnd FILL
X_1015_ _1040_/B _1079_/C _1040_/A _1020_/A vdd gnd AOI21X1
XFILL_1__755_ vdd gnd FILL
XFILL_1__824_ vdd gnd FILL
XFILL_1__1200_ vdd gnd FILL
XFILL_1__1131_ vdd gnd FILL
XFILL_1__1062_ vdd gnd FILL
XFILL_2__1240_ vdd gnd FILL
XFILL_2__1171_ vdd gnd FILL
XFILL_0__773_ vdd gnd FILL
XFILL_1__1329_ vdd gnd FILL
XFILL_0__842_ vdd gnd FILL
XFILL_0__911_ vdd gnd FILL
XFILL_3__984_ vdd gnd FILL
X_726_ _743_/A _726_/B _743_/C _730_/B vdd gnd OAI21X1
XFILL_2__1438_ vdd gnd FILL
XFILL_0_BUFX2_insert2 vdd gnd FILL
XFILL_2__1369_ vdd gnd FILL
XFILL_0__1005_ vdd gnd FILL
X_1495_ _1495_/D _1508_/CLK _734_/B vdd gnd DFFPOSX1
XFILL_1__807_ vdd gnd FILL
XFILL_1__738_ vdd gnd FILL
XFILL_1__1114_ vdd gnd FILL
XFILL_1__1045_ vdd gnd FILL
XFILL_2__1223_ vdd gnd FILL
XFILL_2__1154_ vdd gnd FILL
XFILL_2__1085_ vdd gnd FILL
XFILL_0__825_ vdd gnd FILL
XFILL_0__756_ vdd gnd FILL
X_1280_ _774_/B _843_/A _1281_/C vdd gnd NOR2X1
X_1478_ _1478_/D _1522_/CLK _968_/A vdd gnd DFFPOSX1
XFILL_2__985_ vdd gnd FILL
XBUFX2_insert23 _817_/Y _1404_/A vdd gnd BUFX2
XFILL_1__1028_ vdd gnd FILL
X_991_ _994_/A _994_/B _999_/C vdd gnd NAND2X1
XFILL_0__1270_ vdd gnd FILL
XFILL_2__1137_ vdd gnd FILL
XFILL_2__1068_ vdd gnd FILL
XFILL_2__1206_ vdd gnd FILL
XFILL_0__808_ vdd gnd FILL
X_1401_ _808_/A _811_/A _1401_/C _1403_/B vdd gnd NAND3X1
XFILL_0__739_ vdd gnd FILL
X_1263_ _1263_/A _1271_/C _1265_/B vdd gnd NAND2X1
X_1332_ _1332_/A _1332_/B _1332_/C _1333_/B vdd gnd NAND3X1
X_1194_ _1221_/A _1204_/C vdd gnd INVX1
XFILL_3__1246_ vdd gnd FILL
XFILL_3__1177_ vdd gnd FILL
XFILL_2__770_ vdd gnd FILL
XFILL_0__1399_ vdd gnd FILL
XFILL_2_CLKBUF1_insert9 vdd gnd FILL
XFILL_2__968_ vdd gnd FILL
XCLKBUF1_insert8 clk _1525_/CLK vdd gnd CLKBUF1
XFILL_2__899_ vdd gnd FILL
XFILL_3__735_ vdd gnd FILL
X_974_ _974_/A _974_/Y vdd gnd INVX1
XFILL_0__1322_ vdd gnd FILL
XFILL_0__1184_ vdd gnd FILL
XFILL_0__1253_ vdd gnd FILL
X_1315_ _786_/A _1317_/C _1316_/B vdd gnd NAND2X1
XFILL_1__986_ vdd gnd FILL
XFILL_1__1362_ vdd gnd FILL
XFILL_1__1431_ vdd gnd FILL
X_1246_ _1246_/A _1257_/C vdd gnd INVX1
X_1177_ _1179_/C _1177_/B _1177_/C _1189_/A vdd gnd NAND3X1
XFILL_2__822_ vdd gnd FILL
XFILL_1__1293_ vdd gnd FILL
XFILL_2__753_ vdd gnd FILL
X_957_ _957_/A _957_/B _957_/C _961_/B vdd gnd AOI21X1
XFILL_1__840_ vdd gnd FILL
XFILL_1__771_ vdd gnd FILL
X_1031_ _1098_/B _969_/Y _1031_/C _1100_/B vdd gnd NAND3X1
X_888_ _895_/C _894_/B _894_/C _905_/B vdd gnd NAND3X1
X_1100_ _1100_/A _1100_/B _1215_/B _1191_/A vdd gnd OAI21X1
XFILL_0__1236_ vdd gnd FILL
XFILL_0__1305_ vdd gnd FILL
XFILL_0__1098_ vdd gnd FILL
XFILL_0__1167_ vdd gnd FILL
XFILL_0_BUFX2_insert22 vdd gnd FILL
XFILL_1__969_ vdd gnd FILL
XFILL_0_BUFX2_insert33 vdd gnd FILL
XFILL_1__1345_ vdd gnd FILL
XFILL_1__1414_ vdd gnd FILL
X_1229_ _1243_/B _1243_/A _1239_/B vdd gnd XNOR2X1
XFILL_2__736_ vdd gnd FILL
XFILL_2__805_ vdd gnd FILL
XFILL_1__1276_ vdd gnd FILL
X_811_ _811_/A _813_/B vdd gnd INVX1
X_742_ _742_/A _742_/B _745_/A vdd gnd NOR2X1
XFILL_2__1385_ vdd gnd FILL
XFILL_0__1021_ vdd gnd FILL
XFILL_0__987_ vdd gnd FILL
XFILL_1__823_ vdd gnd FILL
XFILL_1__754_ vdd gnd FILL
X_1014_ _957_/C _1014_/B _975_/A _1088_/C vdd gnd OAI21X1
XFILL_0__1219_ vdd gnd FILL
XFILL_1__1130_ vdd gnd FILL
XFILL_1__1061_ vdd gnd FILL
XFILL_1__1328_ vdd gnd FILL
XFILL_0__910_ vdd gnd FILL
XFILL_2__1170_ vdd gnd FILL
XFILL_1__1259_ vdd gnd FILL
XFILL_0__772_ vdd gnd FILL
XFILL_0__841_ vdd gnd FILL
X_725_ _727_/A _744_/A _743_/C vdd gnd NOR2X1
XFILL_0_BUFX2_insert3 vdd gnd FILL
XFILL_2__1437_ vdd gnd FILL
XFILL_2__1299_ vdd gnd FILL
XFILL_2__1368_ vdd gnd FILL
XFILL87150x11850 vdd gnd FILL
X_1494_ _1494_/D _1515_/CLK _726_/B vdd gnd DFFPOSX1
XFILL_0__1004_ vdd gnd FILL
XFILL_1__806_ vdd gnd FILL
XFILL_1__737_ vdd gnd FILL
XFILL_1__1113_ vdd gnd FILL
XFILL_1__1044_ vdd gnd FILL
XFILL_2__1222_ vdd gnd FILL
XFILL_2__1153_ vdd gnd FILL
XFILL_2__1084_ vdd gnd FILL
XFILL_0__824_ vdd gnd FILL
XFILL_0__755_ vdd gnd FILL
XFILL_3__1193_ vdd gnd FILL
XFILL87150x23550 vdd gnd FILL
X_1477_ _967_/Y _1525_/CLK _966_/A vdd gnd DFFPOSX1
XBUFX2_insert24 _817_/Y _1391_/B vdd gnd BUFX2
XFILL_2__984_ vdd gnd FILL
XFILL_1__1027_ vdd gnd FILL
X_990_ _990_/A Cin[2] _996_/A vdd gnd NAND2X1
XFILL_2__1205_ vdd gnd FILL
XFILL_0__807_ vdd gnd FILL
XFILL_2__1136_ vdd gnd FILL
XFILL_2__1067_ vdd gnd FILL
XFILL_0__738_ vdd gnd FILL
X_1400_ _742_/B _1404_/A _1404_/C vdd gnd NAND2X1
X_1331_ _1331_/A _1331_/B _1332_/A vdd gnd NOR2X1
X_1262_ _768_/B _816_/A _1263_/A vdd gnd NAND2X1
XFILL_3__1314_ vdd gnd FILL
XFILL87150x35250 vdd gnd FILL
X_1193_ _1193_/A _1227_/B _1193_/C _1221_/A vdd gnd OAI21X1
XFILL_0__1398_ vdd gnd FILL
X_1529_ _751_/Y Xout[1] vdd gnd BUFX2
XFILL_2__967_ vdd gnd FILL
XFILL_2__898_ vdd gnd FILL
XCLKBUF1_insert9 clk _1503_/CLK vdd gnd CLKBUF1
X_973_ _973_/A _985_/C _973_/C _974_/A vdd gnd OAI21X1
XFILL_3__803_ vdd gnd FILL
XFILL_0__1252_ vdd gnd FILL
XFILL_0__1321_ vdd gnd FILL
XFILL_0__1183_ vdd gnd FILL
XFILL_2__1119_ vdd gnd FILL
X_1314_ _1329_/B _1314_/B _1317_/C vdd gnd NAND2X1
XFILL_1__985_ vdd gnd FILL
XFILL_1__1361_ vdd gnd FILL
XFILL_1__1430_ vdd gnd FILL
X_1245_ _1247_/C _1245_/B _1258_/A vdd gnd OR2X2
X_1176_ _1192_/B _1180_/B _1177_/C vdd gnd NAND2X1
XFILL_2__821_ vdd gnd FILL
XFILL_1__1292_ vdd gnd FILL
XFILL_2__752_ vdd gnd FILL
XFILL_1__770_ vdd gnd FILL
X_956_ _976_/B _975_/A _976_/A _961_/A vdd gnd AOI21X1
X_887_ _933_/C _895_/C vdd gnd INVX1
X_1030_ _1030_/A _1030_/B _1034_/A _1031_/C vdd gnd OAI21X1
XFILL_0__1304_ vdd gnd FILL
XFILL_0__1235_ vdd gnd FILL
XFILL_0__1166_ vdd gnd FILL
XFILL_0__1097_ vdd gnd FILL
XFILL_0_BUFX2_insert23 vdd gnd FILL
X_1228_ _1246_/A _1228_/B _1243_/B vdd gnd AND2X2
XFILL_1__899_ vdd gnd FILL
XFILL_1__968_ vdd gnd FILL
XFILL_1__1275_ vdd gnd FILL
XFILL_1__1344_ vdd gnd FILL
XFILL_1__1413_ vdd gnd FILL
X_1159_ _994_/A Cin[3] _1193_/A vdd gnd NAND2X1
XFILL_2__804_ vdd gnd FILL
XFILL_2__735_ vdd gnd FILL
X_810_ _813_/A _810_/B _810_/C _810_/Y vdd gnd OAI21X1
XFILL_2__1384_ vdd gnd FILL
X_741_ _741_/A _741_/B _741_/C _741_/Y vdd gnd OAI21X1
XFILL_0__1020_ vdd gnd FILL
XFILL_0__986_ vdd gnd FILL
XFILL_1__822_ vdd gnd FILL
XFILL_1__753_ vdd gnd FILL
X_939_ _947_/C _947_/A _947_/B _951_/B vdd gnd NAND3X1
X_1013_ _951_/C _951_/B _951_/A _1014_/B vdd gnd AOI21X1
XFILL_0__1218_ vdd gnd FILL
XFILL_0__1149_ vdd gnd FILL
XFILL_1__1060_ vdd gnd FILL
XFILL_1__1258_ vdd gnd FILL
XFILL_1__1327_ vdd gnd FILL
XFILL_0__840_ vdd gnd FILL
XFILL_0__771_ vdd gnd FILL
XFILL_1__1189_ vdd gnd FILL
X_724_ _742_/A _743_/A vdd gnd INVX2
XFILL_2__1367_ vdd gnd FILL
XFILL_2__1436_ vdd gnd FILL
XFILL_0_BUFX2_insert4 vdd gnd FILL
XFILL_2__1298_ vdd gnd FILL
XFILL_0__1003_ vdd gnd FILL
XFILL_0__969_ vdd gnd FILL
X_1493_ _1493_/D _1525_/CLK _744_/D vdd gnd DFFPOSX1
XFILL_1__736_ vdd gnd FILL
XFILL_1__805_ vdd gnd FILL
XFILL_1__1112_ vdd gnd FILL
XFILL_1__1043_ vdd gnd FILL
XFILL_2__1221_ vdd gnd FILL
XFILL_2__1083_ vdd gnd FILL
XFILL_2__1152_ vdd gnd FILL
XFILL_0__823_ vdd gnd FILL
XFILL_0__754_ vdd gnd FILL
XFILL_2__1419_ vdd gnd FILL
XFILL_3__1261_ vdd gnd FILL
X_1476_ _917_/Y _1522_/CLK _877_/A vdd gnd DFFPOSX1
XBUFX2_insert25 _1522_/Q _757_/A vdd gnd BUFX2
XFILL_2__983_ vdd gnd FILL
XFILL_1__1026_ vdd gnd FILL
XFILL_3__750_ vdd gnd FILL
XFILL_2__1204_ vdd gnd FILL
XFILL_2__1135_ vdd gnd FILL
XFILL_0__737_ vdd gnd FILL
XFILL_0__806_ vdd gnd FILL
XFILL_2__1066_ vdd gnd FILL
X_1261_ _1270_/A _1271_/C vdd gnd INVX1
X_1330_ _1330_/A _1332_/B _1330_/C _1333_/A vdd gnd AOI21X1
XFILL_0__1535_ vdd gnd FILL
X_1192_ _1192_/A _1192_/B _1209_/B vdd gnd NAND2X1
XFILL_0__1397_ vdd gnd FILL
X_1459_ _777_/Y _1522_/CLK _775_/A vdd gnd DFFPOSX1
X_1528_ _748_/Y Xout[0] vdd gnd BUFX2
XFILL_2__966_ vdd gnd FILL
XFILL_1__1009_ vdd gnd FILL
XFILL_2__897_ vdd gnd FILL
X_972_ _980_/A Cin[4] _985_/C vdd gnd NAND2X1
XFILL_0__1251_ vdd gnd FILL
XFILL_0__1182_ vdd gnd FILL
XFILL_0__1320_ vdd gnd FILL
XFILL_2__1118_ vdd gnd FILL
XFILL_2__1049_ vdd gnd FILL
X_1313_ _1329_/B _1314_/B _1316_/A vdd gnd NOR2X1
X_1244_ _999_/A _979_/B _1244_/C _1245_/B vdd gnd OAI21X1
XFILL_1__984_ vdd gnd FILL
XFILL_1__1360_ vdd gnd FILL
XFILL_1__1291_ vdd gnd FILL
X_1175_ _1175_/A _1175_/B _1175_/C _1180_/B vdd gnd NAND3X1
XFILL_2__820_ vdd gnd FILL
XFILL86250x11850 vdd gnd FILL
XFILL_2__751_ vdd gnd FILL
XFILL_0__1449_ vdd gnd FILL
XFILL86850x4050 vdd gnd FILL
XFILL_2__949_ vdd gnd FILL
X_955_ _955_/A _955_/B _955_/C _970_/C vdd gnd OAI21X1
X_886_ _980_/A Cin[2] _933_/C vdd gnd NAND2X1
XFILL_0__1303_ vdd gnd FILL
XFILL_0__1234_ vdd gnd FILL
XFILL_0__1165_ vdd gnd FILL
XFILL_0__1096_ vdd gnd FILL
XFILL_1__1412_ vdd gnd FILL
XFILL_0_BUFX2_insert24 vdd gnd FILL
XFILL_1__967_ vdd gnd FILL
X_1227_ _1247_/A _1227_/B _1246_/A vdd gnd OR2X2
XFILL_1__898_ vdd gnd FILL
X_1158_ _1158_/A _1161_/C _1158_/C _1193_/C vdd gnd NAND3X1
XFILL_1__1274_ vdd gnd FILL
XFILL_1__1343_ vdd gnd FILL
XFILL_2__803_ vdd gnd FILL
X_1089_ _974_/Y _1089_/B _1089_/C _1092_/A vdd gnd OAI21X1
XFILL86250x23550 vdd gnd FILL
XFILL_2__734_ vdd gnd FILL
X_740_ _744_/A _740_/B _765_/B _740_/D _741_/C vdd gnd AOI22X1
XFILL_2__1383_ vdd gnd FILL
XFILL_0__985_ vdd gnd FILL
XFILL_1__821_ vdd gnd FILL
XFILL_1__752_ vdd gnd FILL
X_1012_ _1088_/B _1088_/A _976_/Y _1029_/A vdd gnd NAND3X1
X_938_ _990_/A _938_/B _988_/B _947_/B vdd gnd NAND3X1
X_869_ _902_/A _919_/B vdd gnd INVX1
XFILL_0__1217_ vdd gnd FILL
XFILL_0__1148_ vdd gnd FILL
XFILL_0__1079_ vdd gnd FILL
XFILL_0__770_ vdd gnd FILL
XFILL_1__1257_ vdd gnd FILL
XFILL_1__1326_ vdd gnd FILL
XFILL_1__1188_ vdd gnd FILL
X_723_ _742_/A _723_/B _730_/A vdd gnd NOR2X1
XFILL_2__1366_ vdd gnd FILL
XFILL_2__1297_ vdd gnd FILL
XFILL_0_BUFX2_insert5 vdd gnd FILL
XFILL_2__1435_ vdd gnd FILL
XFILL_0__899_ vdd gnd FILL
XFILL_0__968_ vdd gnd FILL
XFILL_0__1002_ vdd gnd FILL
X_1492_ _1492_/D _1522_/CLK _740_/D vdd gnd DFFPOSX1
XFILL_1__804_ vdd gnd FILL
XFILL_1__735_ vdd gnd FILL
XFILL_1__1111_ vdd gnd FILL
XFILL_1__1042_ vdd gnd FILL
XFILL_2__1220_ vdd gnd FILL
XFILL_2__1151_ vdd gnd FILL
XFILL_0__822_ vdd gnd FILL
XFILL_1__1309_ vdd gnd FILL
XFILL_0__753_ vdd gnd FILL
XFILL_2__1082_ vdd gnd FILL
XFILL_2__1418_ vdd gnd FILL
XFILL_2__1349_ vdd gnd FILL
X_1475_ _876_/Y _1522_/CLK _845_/A vdd gnd DFFPOSX1
XFILL_3__1389_ vdd gnd FILL
XFILL_2__982_ vdd gnd FILL
XBUFX2_insert26 _1522_/Q _728_/A vdd gnd BUFX2
XFILL_1__1025_ vdd gnd FILL
XBUFX2_insert15 Cin[0] _993_/B vdd gnd BUFX2
XFILL_2__1203_ vdd gnd FILL
XFILL_2__1134_ vdd gnd FILL
XFILL_0__736_ vdd gnd FILL
XFILL_0__805_ vdd gnd FILL
XFILL_2__1065_ vdd gnd FILL
X_1260_ _768_/B _816_/A _1270_/A vdd gnd NOR2X1
X_1191_ _1191_/A _1191_/B _1217_/A _1242_/B vdd gnd AOI21X1
XFILL_3__947_ vdd gnd FILL
XFILL_3__878_ vdd gnd FILL
XFILL_0__1534_ vdd gnd FILL
XFILL_0__1396_ vdd gnd FILL
X_1527_ _786_/A Vld vdd gnd BUFX2
X_1389_ _1390_/A _1394_/A _1391_/C vdd gnd OR2X2
X_1458_ _774_/Y _1523_/CLK _772_/A vdd gnd DFFPOSX1
XFILL_2__965_ vdd gnd FILL
XFILL_2__896_ vdd gnd FILL
XFILL_1__1008_ vdd gnd FILL
X_971_ _971_/A _971_/B _971_/C _971_/Y vdd gnd OAI21X1
XFILL_0__1250_ vdd gnd FILL
XFILL_0__1181_ vdd gnd FILL
XFILL_2__1117_ vdd gnd FILL
XFILL_2__1048_ vdd gnd FILL
X_1243_ _1243_/A _1243_/B _1247_/C vdd gnd NAND2X1
X_1312_ _784_/A _968_/A _1329_/B vdd gnd XOR2X1
XFILL_1__983_ vdd gnd FILL
X_1174_ _1174_/A _1174_/B _1174_/C _1175_/C vdd gnd OAI21X1
XFILL_1__1290_ vdd gnd FILL
XFILL_0__1448_ vdd gnd FILL
XFILL_0__1379_ vdd gnd FILL
XFILL_2__750_ vdd gnd FILL
XFILL_2__948_ vdd gnd FILL
XFILL_2__879_ vdd gnd FILL
X_954_ _970_/A _970_/B _961_/C _959_/B vdd gnd NAND3X1
X_885_ _933_/D _894_/B vdd gnd INVX1
XFILL_0__1302_ vdd gnd FILL
XFILL_3__1011_ vdd gnd FILL
XFILL_0__1233_ vdd gnd FILL
XFILL_2_CLKBUF1_insert10 vdd gnd FILL
XFILL_0__1095_ vdd gnd FILL
XFILL_0__1164_ vdd gnd FILL
XFILL_1__966_ vdd gnd FILL
XFILL_1__1342_ vdd gnd FILL
XFILL_1__1411_ vdd gnd FILL
X_1226_ _1244_/C _1247_/A vdd gnd INVX1
XFILL_0_BUFX2_insert25 vdd gnd FILL
X_1157_ _999_/A _985_/B _1157_/C _1161_/C vdd gnd OAI21X1
XFILL_1__897_ vdd gnd FILL
XFILL_1__1273_ vdd gnd FILL
XFILL_2__802_ vdd gnd FILL
X_1088_ _1088_/A _1088_/B _1088_/C _1089_/B vdd gnd AOI21X1
XFILL_2__733_ vdd gnd FILL
XFILL_2__1451_ vdd gnd FILL
XFILL_2__1382_ vdd gnd FILL
XFILL_0__984_ vdd gnd FILL
XFILL_1__820_ vdd gnd FILL
X_799_ _799_/A _801_/B vdd gnd INVX1
X_1011_ _1079_/C _1040_/B _1040_/A _1088_/A vdd gnd NAND3X1
X_937_ _994_/A _941_/B _988_/B vdd gnd NAND2X1
X_868_ _902_/A _868_/B _868_/C _874_/B vdd gnd NAND3X1
XFILL_1__751_ vdd gnd FILL
XFILL_0__1216_ vdd gnd FILL
XFILL_0__1147_ vdd gnd FILL
XFILL_0__1078_ vdd gnd FILL
XFILL_1__949_ vdd gnd FILL
XFILL_1__1325_ vdd gnd FILL
X_1209_ _1209_/A _1209_/B _1241_/C vdd gnd OR2X2
XFILL_1__1256_ vdd gnd FILL
XFILL_1__1187_ vdd gnd FILL
XFILL_2__1434_ vdd gnd FILL
XFILL_2__1365_ vdd gnd FILL
XFILL_2__1296_ vdd gnd FILL
XFILL_0_BUFX2_insert6 vdd gnd FILL
XFILL_0__967_ vdd gnd FILL
XFILL_0__898_ vdd gnd FILL
XFILL_0__1001_ vdd gnd FILL
X_1491_ _1491_/D _1525_/CLK _735_/D vdd gnd DFFPOSX1
XFILL_1__803_ vdd gnd FILL
XFILL_1__734_ vdd gnd FILL
XFILL_1__1110_ vdd gnd FILL
XFILL_1__1041_ vdd gnd FILL
XFILL_1__1308_ vdd gnd FILL
XFILL_2__1081_ vdd gnd FILL
XFILL_2__1150_ vdd gnd FILL
XFILL_0__821_ vdd gnd FILL
XFILL_1__1239_ vdd gnd FILL
XFILL_0__752_ vdd gnd FILL
XFILL_3__894_ vdd gnd FILL
XFILL_2__1417_ vdd gnd FILL
XFILL_2__1348_ vdd gnd FILL
XFILL_2__1279_ vdd gnd FILL
X_1474_ _844_/Y _1523_/CLK _842_/A vdd gnd DFFPOSX1
XFILL_2__981_ vdd gnd FILL
XBUFX2_insert27 _1522_/Q _1523_/D vdd gnd BUFX2
XFILL_1__1024_ vdd gnd FILL
XBUFX2_insert16 Cin[0] _884_/B vdd gnd BUFX2
XFILL_0__804_ vdd gnd FILL
XFILL_2__1202_ vdd gnd FILL
XFILL_2__1064_ vdd gnd FILL
XFILL_2__1133_ vdd gnd FILL
XFILL_0__735_ vdd gnd FILL
X_1190_ _1251_/A _1217_/A vdd gnd INVX1
XFILL_0__1533_ vdd gnd FILL
XFILL_0__1395_ vdd gnd FILL
X_1457_ _771_/Y _1515_/CLK _769_/A vdd gnd DFFPOSX1
X_1526_ _1526_/D _1526_/CLK _1526_/Q vdd gnd DFFPOSX1
X_1388_ _1392_/A _1394_/A vdd gnd INVX1
XFILL_2__895_ vdd gnd FILL
XFILL_2__964_ vdd gnd FILL
X_970_ _970_/A _970_/B _970_/C _971_/B vdd gnd AOI21X1
XFILL_1__1007_ vdd gnd FILL
XFILL_2__1116_ vdd gnd FILL
XFILL_2__1047_ vdd gnd FILL
XFILL_0__1180_ vdd gnd FILL
X_1311_ _1331_/A _1311_/B _1326_/C _1314_/B vdd gnd OAI21X1
XFILL_1__982_ vdd gnd FILL
X_1242_ _1251_/B _1242_/B _1251_/C _1257_/A vdd gnd OAI21X1
X_1173_ _1202_/B _1173_/B _1173_/C _1175_/B vdd gnd NAND3X1
XFILL_0__1378_ vdd gnd FILL
XFILL_3__1087_ vdd gnd FILL
XFILL_0__1447_ vdd gnd FILL
X_1509_ _1509_/D _1526_/CLK _800_/B vdd gnd DFFPOSX1
XFILL_2__947_ vdd gnd FILL
XFILL_2__878_ vdd gnd FILL
X_953_ _975_/A _976_/A _976_/B _970_/B vdd gnd NAND3X1
X_884_ _990_/A _884_/B _978_/A _938_/B _933_/D vdd gnd AOI22X1
XFILL_0__1232_ vdd gnd FILL
XFILL_0__1301_ vdd gnd FILL
XFILL_2_CLKBUF1_insert11 vdd gnd FILL
XFILL_0__1094_ vdd gnd FILL
XFILL_0__1163_ vdd gnd FILL
XFILL_0_BUFX2_insert15 vdd gnd FILL
XFILL_1__965_ vdd gnd FILL
XFILL_1__1341_ vdd gnd FILL
XFILL_1__1410_ vdd gnd FILL
XFILL_0_BUFX2_insert26 vdd gnd FILL
X_1225_ _765_/A _1225_/B _1244_/C vdd gnd NOR2X1
X_1156_ _1157_/C _1223_/A _1158_/C vdd gnd OR2X2
XFILL_1__896_ vdd gnd FILL
X_1087_ _1087_/A _1087_/B _1087_/C _1212_/A vdd gnd OAI21X1
XFILL_2__732_ vdd gnd FILL
XFILL_1__1272_ vdd gnd FILL
XFILL_2__801_ vdd gnd FILL
XFILL_3__1208_ vdd gnd FILL
XFILL_2__1450_ vdd gnd FILL
XFILL_2__1381_ vdd gnd FILL
XFILL_0__983_ vdd gnd FILL
X_936_ _994_/A _941_/B _988_/A _947_/A vdd gnd NAND3X1
X_798_ _812_/A _798_/B _798_/C _798_/Y vdd gnd OAI21X1
X_1010_ _1010_/A _1010_/B _989_/Y _1040_/B vdd gnd OAI21X1
X_867_ _871_/A _871_/B _879_/C _868_/C vdd gnd OAI21X1
XFILL_1__750_ vdd gnd FILL
XFILL_0__1215_ vdd gnd FILL
XFILL87150x31350 vdd gnd FILL
XFILL_0__1146_ vdd gnd FILL
XFILL_0__1077_ vdd gnd FILL
X_1208_ _1209_/B _1209_/A _1241_/A vdd gnd NAND2X1
XFILL_1__948_ vdd gnd FILL
XFILL_1__879_ vdd gnd FILL
XFILL_1__1255_ vdd gnd FILL
XFILL_1__1324_ vdd gnd FILL
X_1139_ _1142_/C _1179_/C _1142_/A _1177_/B vdd gnd NAND3X1
XFILL_1__1186_ vdd gnd FILL
XFILL_2__1364_ vdd gnd FILL
XFILL_2__1433_ vdd gnd FILL
XFILL_2__1295_ vdd gnd FILL
XFILL_0__966_ vdd gnd FILL
XFILL_0__1000_ vdd gnd FILL
X_1490_ _1490_/D _1515_/CLK _729_/D vdd gnd DFFPOSX1
XFILL_0__897_ vdd gnd FILL
XFILL_1__733_ vdd gnd FILL
XFILL_1__802_ vdd gnd FILL
X_919_ _929_/A _919_/B _971_/A vdd gnd NAND2X1
XFILL87150x43050 vdd gnd FILL
XFILL_1__1040_ vdd gnd FILL
XFILL_0__1129_ vdd gnd FILL
XFILL_1__1307_ vdd gnd FILL
XFILL_1__1238_ vdd gnd FILL
XFILL_0__820_ vdd gnd FILL
XFILL_2__1080_ vdd gnd FILL
XFILL_0__751_ vdd gnd FILL
XFILL_1__1169_ vdd gnd FILL
XFILL_3__962_ vdd gnd FILL
XFILL_2__1347_ vdd gnd FILL
XFILL_2__1416_ vdd gnd FILL
XFILL_2__1278_ vdd gnd FILL
XFILL_0__949_ vdd gnd FILL
X_1473_ _822_/Y _1525_/CLK _821_/A vdd gnd DFFPOSX1
XFILL_2__980_ vdd gnd FILL
XBUFX2_insert28 _1522_/Q _751_/A vdd gnd BUFX2
XFILL_1__1023_ vdd gnd FILL
XBUFX2_insert17 Cin[0] _941_/B vdd gnd BUFX2
XFILL_2__1201_ vdd gnd FILL
XFILL_0__803_ vdd gnd FILL
XFILL_2__1063_ vdd gnd FILL
XFILL_2__1132_ vdd gnd FILL
XFILL_0__734_ vdd gnd FILL
XFILL_0__1532_ vdd gnd FILL
XFILL_0__1394_ vdd gnd FILL
X_1387_ _1387_/A _1392_/C _1392_/A vdd gnd NOR2X1
X_1525_ _742_/A _1525_/CLK _1526_/D vdd gnd DFFPOSX1
X_1456_ _768_/Y _1522_/CLK _766_/A vdd gnd DFFPOSX1
XFILL_2__894_ vdd gnd FILL
XFILL_2__963_ vdd gnd FILL
XFILL_1__1006_ vdd gnd FILL
XFILL_2__1115_ vdd gnd FILL
XFILL_2__1046_ vdd gnd FILL
X_1310_ _740_/D _843_/B _1316_/C vdd gnd NAND2X1
X_1241_ _1241_/A _1241_/B _1241_/C _1251_/B vdd gnd NAND3X1
XFILL_1__981_ vdd gnd FILL
X_1172_ _1172_/A _1192_/A _1172_/C _1192_/B vdd gnd NAND3X1
XFILL_0__1377_ vdd gnd FILL
XFILL_3__1155_ vdd gnd FILL
XFILL_0__1446_ vdd gnd FILL
X_1439_ _744_/A _1439_/B _1439_/C _1515_/D vdd gnd AOI21X1
X_1508_ _1508_/D _1508_/CLK _797_/B vdd gnd DFFPOSX1
XFILL_2__877_ vdd gnd FILL
XFILL_2__946_ vdd gnd FILL
X_952_ _952_/A _952_/B _952_/C _976_/B vdd gnd OAI21X1
X_883_ _883_/A _942_/A _894_/C vdd gnd NAND2X1
XFILL_0__1300_ vdd gnd FILL
XFILL_0__1231_ vdd gnd FILL
XFILL_0__1162_ vdd gnd FILL
XFILL_2_CLKBUF1_insert12 vdd gnd FILL
XFILL_0__1093_ vdd gnd FILL
XFILL_2__1029_ vdd gnd FILL
X_1224_ _999_/A _1225_/B _1224_/C _1228_/B vdd gnd OAI21X1
XFILL_0_BUFX2_insert27 vdd gnd FILL
XFILL_1__895_ vdd gnd FILL
XFILL_1__964_ vdd gnd FILL
XFILL_0_BUFX2_insert16 vdd gnd FILL
XFILL_1__1340_ vdd gnd FILL
XFILL_1__1271_ vdd gnd FILL
X_1155_ _997_/A Cin[3] _1223_/A vdd gnd NAND2X1
X_1086_ _1090_/C _1102_/C _1090_/A _1087_/A vdd gnd AOI21X1
XFILL_2__731_ vdd gnd FILL
XFILL_2__800_ vdd gnd FILL
XFILL_0__1429_ vdd gnd FILL
XFILL_2__1380_ vdd gnd FILL
XFILL_0__982_ vdd gnd FILL
XFILL_2__929_ vdd gnd FILL
X_935_ _978_/A Cin[2] _947_/C vdd gnd NAND2X1
X_866_ _866_/A _866_/B _881_/A _871_/B vdd gnd AOI21X1
X_797_ _812_/A _797_/B _798_/C vdd gnd NAND2X1
XFILL_0__1145_ vdd gnd FILL
XFILL_0__1214_ vdd gnd FILL
XFILL_0__1076_ vdd gnd FILL
XFILL_1__947_ vdd gnd FILL
XFILL_1__878_ vdd gnd FILL
X_1207_ _1207_/A _1207_/B _1209_/A vdd gnd AND2X2
XFILL_1__1323_ vdd gnd FILL
XFILL_1__1254_ vdd gnd FILL
X_1138_ _1138_/A _1138_/B _1138_/C _1142_/A vdd gnd OAI21X1
X_1069_ _765_/A _999_/B _998_/B _1070_/B vdd gnd OAI21X1
XFILL_1__1185_ vdd gnd FILL
XFILL_2__1363_ vdd gnd FILL
XFILL_2__1294_ vdd gnd FILL
XFILL_2__1432_ vdd gnd FILL
XFILL_0__896_ vdd gnd FILL
XFILL_0__965_ vdd gnd FILL
XFILL_1__732_ vdd gnd FILL
XFILL_1__801_ vdd gnd FILL
X_849_ _978_/A _884_/B _933_/A vdd gnd NAND2X1
X_918_ _977_/A Cin[4] _929_/A vdd gnd AND2X2
XFILL_0__1128_ vdd gnd FILL
XFILL_0__1059_ vdd gnd FILL
XFILL_1__1237_ vdd gnd FILL
XFILL_1__1306_ vdd gnd FILL
XFILL_1__1168_ vdd gnd FILL
XFILL_0__750_ vdd gnd FILL
XFILL_1__1099_ vdd gnd FILL
XFILL_2__1415_ vdd gnd FILL
XFILL_2__1346_ vdd gnd FILL
XFILL_2__1277_ vdd gnd FILL
XFILL_0__948_ vdd gnd FILL
XFILL_0__879_ vdd gnd FILL
X_1472_ _816_/Y _1522_/CLK _814_/A vdd gnd DFFPOSX1
XBUFX2_insert29 _1522_/Q _744_/A vdd gnd BUFX2
XFILL_1__1022_ vdd gnd FILL
XBUFX2_insert18 Cin[0] _835_/B vdd gnd BUFX2
XFILL_2__1200_ vdd gnd FILL
XFILL_2__1131_ vdd gnd FILL
XFILL_0__733_ vdd gnd FILL
XFILL_0__802_ vdd gnd FILL
XFILL_2__1062_ vdd gnd FILL
XFILL_0__1531_ vdd gnd FILL
XFILL_0__1393_ vdd gnd FILL
XFILL_2__1329_ vdd gnd FILL
X_1524_ _727_/A _1525_/CLK _742_/A vdd gnd DFFPOSX1
X_1386_ _807_/B _1386_/B _1392_/C vdd gnd NOR2X1
X_1455_ _765_/Y _1521_/CLK _755_/A vdd gnd DFFPOSX1
XFILL_2__962_ vdd gnd FILL
XFILL_1__1005_ vdd gnd FILL
XFILL_2__893_ vdd gnd FILL
XFILL_2__1114_ vdd gnd FILL
XFILL_2__1045_ vdd gnd FILL
X_1240_ _1240_/A _1240_/B _1251_/C vdd gnd NOR2X1
XFILL_1__980_ vdd gnd FILL
X_1171_ _1174_/A _1174_/B _1173_/C _1172_/C vdd gnd OAI21X1
XFILL_3__1223_ vdd gnd FILL
XFILL_0__1445_ vdd gnd FILL
XFILL_0__1376_ vdd gnd FILL
X_1507_ _1507_/D _1525_/CLK _794_/B vdd gnd DFFPOSX1
X_1438_ _744_/A _770_/B _1439_/C vdd gnd NOR2X1
X_1369_ _743_/B _1370_/A _1370_/C vdd gnd NAND2X1
XFILL_2__945_ vdd gnd FILL
XFILL_2__876_ vdd gnd FILL
X_951_ _951_/A _951_/B _951_/C _975_/A vdd gnd NAND3X1
X_882_ _990_/A _938_/B _942_/A vdd gnd AND2X2
XFILL_0__1230_ vdd gnd FILL
XFILL_0__1161_ vdd gnd FILL
XFILL_0__1092_ vdd gnd FILL
XFILL_2__1028_ vdd gnd FILL
XFILL_2_CLKBUF1_insert13 vdd gnd FILL
XFILL_0_BUFX2_insert28 vdd gnd FILL
X_1223_ _1223_/A _1224_/C _1223_/C _1223_/D _1243_/A vdd gnd OAI22X1
XFILL_1__894_ vdd gnd FILL
XFILL_0_BUFX2_insert17 vdd gnd FILL
XFILL_1__963_ vdd gnd FILL
X_1154_ _994_/A Cin[4] _1157_/C vdd gnd NAND2X1
XFILL_1__1270_ vdd gnd FILL
XFILL_0__1428_ vdd gnd FILL
X_1085_ _1085_/A _1085_/B _1085_/C _1090_/C vdd gnd OAI21X1
XFILL_2__730_ vdd gnd FILL
XFILL_0__1359_ vdd gnd FILL
XFILL_1__1399_ vdd gnd FILL
XFILL_2__928_ vdd gnd FILL
XFILL_0__981_ vdd gnd FILL
XFILL_2__859_ vdd gnd FILL
X_796_ _796_/A _798_/B vdd gnd INVX1
X_934_ _951_/A _952_/C vdd gnd INVX1
X_865_ _985_/A _999_/B _865_/C _866_/B vdd gnd OAI21X1
XFILL_0__1213_ vdd gnd FILL
XFILL_0__1075_ vdd gnd FILL
XFILL_0__1144_ vdd gnd FILL
XFILL_1__877_ vdd gnd FILL
XFILL_1__946_ vdd gnd FILL
X_1137_ _1178_/B _1178_/A _1178_/C _1179_/C vdd gnd NAND3X1
X_1206_ _1221_/A _1221_/B _1206_/C _1207_/B vdd gnd NAND3X1
XFILL_1__1184_ vdd gnd FILL
XFILL_1__1253_ vdd gnd FILL
XFILL_1__1322_ vdd gnd FILL
X_1068_ _999_/A _862_/B _1068_/C _1070_/A vdd gnd OAI21X1
XFILL_2__1431_ vdd gnd FILL
XFILL_2__1362_ vdd gnd FILL
XFILL_2__1293_ vdd gnd FILL
XFILL86850x7950 vdd gnd FILL
XFILL_0__895_ vdd gnd FILL
XFILL_0__964_ vdd gnd FILL
XFILL_1__800_ vdd gnd FILL
XFILL_1__731_ vdd gnd FILL
X_779_ _786_/A _779_/B _780_/C vdd gnd NAND2X1
X_848_ _977_/A Cin[2] _881_/A vdd gnd NAND2X1
X_917_ _917_/A _917_/B _917_/C _917_/D _917_/Y vdd gnd OAI22X1
XFILL_0__1127_ vdd gnd FILL
XFILL_0__1058_ vdd gnd FILL
XFILL_1__929_ vdd gnd FILL
XFILL_1__1305_ vdd gnd FILL
XFILL_1__1236_ vdd gnd FILL
XFILL_1__1098_ vdd gnd FILL
XFILL_1__1167_ vdd gnd FILL
XFILL_2__1414_ vdd gnd FILL
XFILL_2__1345_ vdd gnd FILL
XFILL_2__1276_ vdd gnd FILL
XFILL_0__947_ vdd gnd FILL
XFILL_0__878_ vdd gnd FILL
X_1471_ _813_/Y _1508_/CLK _811_/A vdd gnd DFFPOSX1
XBUFX2_insert19 _817_/Y _843_/B vdd gnd BUFX2
XFILL_1__1021_ vdd gnd FILL
XFILL_2__1130_ vdd gnd FILL
XFILL_2__1061_ vdd gnd FILL
XFILL_0__732_ vdd gnd FILL
XFILL_0__801_ vdd gnd FILL
XFILL_1__1219_ vdd gnd FILL
XFILL_0__1530_ vdd gnd FILL
XFILL_3__1170_ vdd gnd FILL
XFILL_0__1392_ vdd gnd FILL
XFILL_2__1259_ vdd gnd FILL
XFILL_2__1328_ vdd gnd FILL
X_1523_ _1523_/D _1523_/CLK _727_/A vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert0 vdd gnd FILL
X_1454_ _763_/Y _1521_/CLK _997_/A vdd gnd DFFPOSX1
X_1385_ _805_/A _1485_/Q _1387_/A vdd gnd NOR2X1
XFILL_3__1299_ vdd gnd FILL
XFILL_2__961_ vdd gnd FILL
XFILL_2__892_ vdd gnd FILL
XFILL_1__1004_ vdd gnd FILL
XFILL_2__1113_ vdd gnd FILL
XFILL_2__1044_ vdd gnd FILL
XFILL_3__788_ vdd gnd FILL
X_1170_ _1202_/B _1174_/B vdd gnd INVX1
XFILL_0__1375_ vdd gnd FILL
XFILL_0__1444_ vdd gnd FILL
X_1506_ _1506_/D _1515_/CLK _791_/B vdd gnd DFFPOSX1
X_1437_ _728_/A _1437_/B _1437_/C _1514_/D vdd gnd AOI21X1
X_1299_ _1350_/A _1299_/B _1299_/C _1490_/D vdd gnd OAI21X1
X_1368_ _1368_/A _1373_/A _1370_/B vdd gnd XOR2X1
XFILL86550x27450 vdd gnd FILL
XFILL_2__944_ vdd gnd FILL
XFILL_2__875_ vdd gnd FILL
X_950_ _950_/A _973_/C _976_/A vdd gnd AND2X2
X_881_ _881_/A _881_/B _881_/C _905_/A vdd gnd OAI21X1
XFILL_2_CLKBUF1_insert14 vdd gnd FILL
XFILL_0__1160_ vdd gnd FILL
XFILL_0__1091_ vdd gnd FILL
XFILL_2__1027_ vdd gnd FILL
XFILL_1__962_ vdd gnd FILL
XFILL_0_BUFX2_insert29 vdd gnd FILL
X_1222_ _1222_/A _1223_/C vdd gnd INVX1
X_1153_ _759_/A _1225_/B _1158_/A vdd gnd NOR2X1
X_1084_ _1101_/C _1101_/B _1101_/A _1102_/C vdd gnd NAND3X1
XFILL_1__893_ vdd gnd FILL
XFILL_3__909_ vdd gnd FILL
XFILL_0_BUFX2_insert18 vdd gnd FILL
XFILL_0__1358_ vdd gnd FILL
XFILL_0__1427_ vdd gnd FILL
XFILL_0__1289_ vdd gnd FILL
XFILL86550x39150 vdd gnd FILL
XFILL_1__1398_ vdd gnd FILL
XFILL_0__980_ vdd gnd FILL
XFILL_2__927_ vdd gnd FILL
XFILL_2__858_ vdd gnd FILL
XFILL_2__789_ vdd gnd FILL
X_933_ _933_/A _988_/A _933_/C _933_/D _951_/A vdd gnd OAI22X1
X_795_ _813_/A _795_/B _795_/C _795_/Y vdd gnd OAI21X1
X_864_ _941_/B _999_/B vdd gnd INVX1
XFILL_0__1212_ vdd gnd FILL
XFILL_0__1143_ vdd gnd FILL
XFILL_0__1074_ vdd gnd FILL
XFILL_1__945_ vdd gnd FILL
XFILL_1__1321_ vdd gnd FILL
X_1136_ _1179_/A _1143_/B _1143_/A _1140_/C vdd gnd NAND3X1
X_1205_ _1221_/C _1206_/C vdd gnd INVX1
X_1067_ _1120_/C _1113_/B _1113_/A _1075_/A vdd gnd AOI21X1
XFILL_1__876_ vdd gnd FILL
XFILL_1__1183_ vdd gnd FILL
XFILL_1__1252_ vdd gnd FILL
XFILL_2__1430_ vdd gnd FILL
XFILL_2__1361_ vdd gnd FILL
XFILL_2__1292_ vdd gnd FILL
XFILL_0__894_ vdd gnd FILL
XFILL_0__963_ vdd gnd FILL
X_916_ _917_/B _969_/C _917_/D vdd gnd NAND2X1
XFILL_1__730_ vdd gnd FILL
X_778_ _778_/A _780_/B vdd gnd INVX1
X_847_ _847_/A _847_/B _847_/C _871_/C vdd gnd AOI21X1
XFILL_0__1126_ vdd gnd FILL
XFILL_3_BUFX2_insert33 vdd gnd FILL
XFILL_0__1057_ vdd gnd FILL
XFILL_1__859_ vdd gnd FILL
XFILL_1__928_ vdd gnd FILL
XFILL_1__1304_ vdd gnd FILL
XFILL_1__1235_ vdd gnd FILL
X_1119_ _1133_/C _1132_/B _1168_/C vdd gnd NOR2X1
XFILL_1__1097_ vdd gnd FILL
XFILL_1__1166_ vdd gnd FILL
XFILL_2__1344_ vdd gnd FILL
XFILL_2__1413_ vdd gnd FILL
XFILL_2__1275_ vdd gnd FILL
XFILL_0__946_ vdd gnd FILL
X_1470_ _810_/Y _1508_/CLK _808_/A vdd gnd DFFPOSX1
XFILL_0__877_ vdd gnd FILL
XFILL_1__1020_ vdd gnd FILL
XFILL_0__1109_ vdd gnd FILL
XFILL_0__800_ vdd gnd FILL
XFILL_1__1218_ vdd gnd FILL
XFILL_2__1060_ vdd gnd FILL
XFILL_0__731_ vdd gnd FILL
XFILL_1__1149_ vdd gnd FILL
XFILL_0__1391_ vdd gnd FILL
XFILL_2__1327_ vdd gnd FILL
XFILL_2__1258_ vdd gnd FILL
XFILL_2__1189_ vdd gnd FILL
XFILL_0__929_ vdd gnd FILL
XFILL_2_BUFX2_insert1 vdd gnd FILL
X_1522_ Rdy _1522_/CLK _1522_/Q vdd gnd DFFPOSX1
X_1453_ _761_/Y _1521_/CLK _994_/A vdd gnd DFFPOSX1
X_1384_ _1394_/B _1384_/B _1384_/C _1390_/A vdd gnd OAI21X1
XFILL_3__1367_ vdd gnd FILL
XFILL_2__960_ vdd gnd FILL
XFILL_2__891_ vdd gnd FILL
XFILL_1__1003_ vdd gnd FILL
XFILL_2__1112_ vdd gnd FILL
XFILL_2__1043_ vdd gnd FILL
XFILL_3__856_ vdd gnd FILL
XFILL_0__1374_ vdd gnd FILL
XFILL_0__1443_ vdd gnd FILL
X_1367_ _1367_/A _1372_/C _1373_/A vdd gnd NOR2X1
X_1505_ _1505_/D _1526_/CLK _812_/B vdd gnd DFFPOSX1
X_1436_ _1523_/D _767_/A _1437_/C vdd gnd NOR2X1
X_1298_ _1301_/C _1298_/B _1299_/B vdd gnd NAND2X1
XFILL_2__943_ vdd gnd FILL
XFILL_2__874_ vdd gnd FILL
X_880_ _902_/A _880_/B _909_/A _908_/B vdd gnd OAI21X1
XFILL_0__1090_ vdd gnd FILL
XFILL_2__1026_ vdd gnd FILL
X_1221_ _1221_/A _1221_/B _1221_/C _1239_/A vdd gnd AOI21X1
XFILL_1__961_ vdd gnd FILL
XFILL_1__892_ vdd gnd FILL
XFILL_0_BUFX2_insert19 vdd gnd FILL
X_1083_ _1091_/C _1091_/B _1102_/A _1087_/B vdd gnd AOI21X1
X_1152_ _1152_/A _1152_/B _1152_/C _1174_/C vdd gnd OAI21X1
XFILL_0__1288_ vdd gnd FILL
XFILL_0__1357_ vdd gnd FILL
XFILL_0__1426_ vdd gnd FILL
X_1419_ _791_/B _1426_/B _1420_/C vdd gnd NOR2X1
XFILL_1__1535_ vdd gnd FILL
XFILL_1__1397_ vdd gnd FILL
XFILL_2__788_ vdd gnd FILL
XFILL_2__857_ vdd gnd FILL
XFILL_2__926_ vdd gnd FILL
X_932_ _973_/C _950_/A _957_/C vdd gnd NAND2X1
X_863_ _978_/A _985_/A vdd gnd INVX2
X_794_ _813_/A _794_/B _795_/C vdd gnd NAND2X1
XFILL_0__1211_ vdd gnd FILL
XFILL_0__1142_ vdd gnd FILL
XFILL_0__1073_ vdd gnd FILL
XFILL_2__1009_ vdd gnd FILL
X_1204_ _1221_/C _1204_/B _1204_/C _1207_/A vdd gnd OAI21X1
XFILL_1__944_ vdd gnd FILL
XFILL_1__875_ vdd gnd FILL
XFILL_1__1251_ vdd gnd FILL
XFILL_1__1320_ vdd gnd FILL
X_1135_ _1138_/A _1138_/B _1178_/C _1143_/B vdd gnd OAI21X1
X_1066_ _996_/A _1066_/B _998_/Y _1129_/C vdd gnd OAI21X1
XFILL_0__1409_ vdd gnd FILL
XFILL_1__1182_ vdd gnd FILL
XFILL_3__1049_ vdd gnd FILL
XFILL_2__1360_ vdd gnd FILL
XFILL_2__1291_ vdd gnd FILL
XFILL_0__962_ vdd gnd FILL
XFILL_1__1449_ vdd gnd FILL
XFILL_0__893_ vdd gnd FILL
XFILL_2__909_ vdd gnd FILL
X_915_ _969_/D _915_/B _915_/C _969_/C vdd gnd NAND3X1
X_846_ _922_/A Cin[3] _902_/A vdd gnd NAND2X1
X_777_ _786_/A _777_/B _777_/C _777_/Y vdd gnd OAI21X1
XFILL_0__1125_ vdd gnd FILL
XFILL_0__1056_ vdd gnd FILL
XFILL_1__927_ vdd gnd FILL
XFILL_1__858_ vdd gnd FILL
XFILL_1__1303_ vdd gnd FILL
XFILL_1__1234_ vdd gnd FILL
XFILL_1__789_ vdd gnd FILL
X_1118_ _1118_/A _1165_/A _1118_/C _1133_/C vdd gnd OAI21X1
X_1049_ _990_/A Cin[3] _1050_/C vdd gnd NAND2X1
XFILL_1__1096_ vdd gnd FILL
XFILL_1__1165_ vdd gnd FILL
XFILL_2__1412_ vdd gnd FILL
XFILL_2__1274_ vdd gnd FILL
XFILL_2__1343_ vdd gnd FILL
XFILL85650x27450 vdd gnd FILL
XFILL_0__945_ vdd gnd FILL
XFILL_0__876_ vdd gnd FILL
X_829_ _859_/A _847_/A vdd gnd INVX1
XFILL_0__1039_ vdd gnd FILL
XFILL_0__1108_ vdd gnd FILL
XFILL_0__730_ vdd gnd FILL
XFILL_1__1217_ vdd gnd FILL
XFILL_1__1148_ vdd gnd FILL
XFILL_1__1079_ vdd gnd FILL
XFILL_0__1390_ vdd gnd FILL
XFILL_2__1257_ vdd gnd FILL
XFILL_2__1326_ vdd gnd FILL
XFILL_2__1188_ vdd gnd FILL
XFILL_0__859_ vdd gnd FILL
XFILL_0__928_ vdd gnd FILL
X_1383_ _1383_/A _1383_/B _1383_/C _1498_/D vdd gnd OAI21X1
XFILL_2_BUFX2_insert2 vdd gnd FILL
XFILL87150x46950 vdd gnd FILL
X_1452_ _759_/Y _1521_/CLK _990_/A vdd gnd DFFPOSX1
X_1521_ _1521_/D _1521_/CLK _978_/A vdd gnd DFFPOSX1
XFILL_3__1435_ vdd gnd FILL
XFILL_2__890_ vdd gnd FILL
XFILL_1__1002_ vdd gnd FILL
XFILL_2__1111_ vdd gnd FILL
XFILL_2__1042_ vdd gnd FILL
XFILL_3__924_ vdd gnd FILL
XFILL_0__1373_ vdd gnd FILL
XFILL_2__1309_ vdd gnd FILL
XFILL_0__1442_ vdd gnd FILL
X_1504_ _1504_/D _1508_/CLK _809_/B vdd gnd DFFPOSX1
XFILL87150x58650 vdd gnd FILL
X_1366_ _1366_/A _1372_/C vdd gnd INVX1
X_1435_ _1443_/B _1435_/B _1435_/C _1513_/D vdd gnd OAI21X1
X_1297_ _1297_/A _1332_/C _1301_/C vdd gnd NAND2X1
XFILL_2__942_ vdd gnd FILL
XFILL_2__873_ vdd gnd FILL
XFILL_2__1025_ vdd gnd FILL
X_1220_ _1483_/Q _1391_/B _1236_/A vdd gnd NAND2X1
XFILL_1__960_ vdd gnd FILL
XFILL_1__891_ vdd gnd FILL
X_1151_ _1175_/A _1172_/A vdd gnd INVX1
XFILL_0__1425_ vdd gnd FILL
X_1082_ _1085_/A _1085_/B _1101_/C _1091_/B vdd gnd OAI21X1
XFILL_0__1356_ vdd gnd FILL
XFILL_0__1287_ vdd gnd FILL
XFILL_1__1534_ vdd gnd FILL
X_1349_ _734_/B _1404_/A _1350_/C vdd gnd NAND2X1
X_1418_ _743_/A _741_/A _1426_/B vdd gnd NOR2X1
XFILL_1__1396_ vdd gnd FILL
XFILL_2__925_ vdd gnd FILL
XFILL_2__787_ vdd gnd FILL
XFILL_2__856_ vdd gnd FILL
X_862_ _979_/A _862_/B _883_/A _866_/A vdd gnd OAI21X1
X_931_ _931_/A _931_/B _931_/C _973_/C vdd gnd NAND3X1
X_793_ _793_/A _795_/B vdd gnd INVX1
XFILL_0__1210_ vdd gnd FILL
XFILL_0__1141_ vdd gnd FILL
XFILL_0__1072_ vdd gnd FILL
XFILL_2__1008_ vdd gnd FILL
X_1203_ _1221_/B _1204_/B vdd gnd INVX1
XFILL_1__943_ vdd gnd FILL
X_1134_ _1134_/A _1134_/B _1152_/B _1138_/B vdd gnd AOI21X1
XFILL_1__874_ vdd gnd FILL
XFILL_0__1408_ vdd gnd FILL
XFILL_1__1250_ vdd gnd FILL
XFILL_1__1181_ vdd gnd FILL
X_1065_ _994_/A _997_/B _997_/A _993_/B _1066_/B vdd gnd AOI22X1
XFILL_3__1117_ vdd gnd FILL
XFILL_0__1339_ vdd gnd FILL
XFILL_2__1290_ vdd gnd FILL
XFILL_1__1379_ vdd gnd FILL
XFILL_0__961_ vdd gnd FILL
XFILL_0__892_ vdd gnd FILL
XFILL_2__908_ vdd gnd FILL
XFILL_1__1448_ vdd gnd FILL
XFILL_2__839_ vdd gnd FILL
X_776_ _815_/C _776_/B _777_/C vdd gnd NAND2X1
X_845_ _845_/A _876_/A vdd gnd INVX1
X_914_ _969_/D _915_/B _915_/C _917_/C vdd gnd AOI21X1
XFILL_0__1055_ vdd gnd FILL
XFILL_0__1124_ vdd gnd FILL
XFILL_1__788_ vdd gnd FILL
XFILL_1__857_ vdd gnd FILL
X_1117_ _765_/A _862_/B _1195_/B _1118_/C vdd gnd OAI21X1
XFILL_1__926_ vdd gnd FILL
XFILL_1__1302_ vdd gnd FILL
XFILL_1__1233_ vdd gnd FILL
XFILL_1__1164_ vdd gnd FILL
X_1048_ _1048_/A _1150_/A _1103_/A vdd gnd NAND2X1
XFILL_1__1095_ vdd gnd FILL
XFILL_2__1411_ vdd gnd FILL
XFILL_2__1273_ vdd gnd FILL
XFILL_2__1342_ vdd gnd FILL
XFILL_0__944_ vdd gnd FILL
XFILL_0__875_ vdd gnd FILL
XFILL_3__1382_ vdd gnd FILL
X_759_ _759_/A _765_/B _759_/C _759_/Y vdd gnd OAI21X1
X_828_ _859_/B _847_/C _859_/A _840_/A vdd gnd OAI21X1
XFILL_0__1038_ vdd gnd FILL
XFILL_0__1107_ vdd gnd FILL
XFILL_1__909_ vdd gnd FILL
XFILL_1__1147_ vdd gnd FILL
XFILL_1__1216_ vdd gnd FILL
XFILL_1__1078_ vdd gnd FILL
XFILL_3__871_ vdd gnd FILL
XFILL_2__1325_ vdd gnd FILL
XFILL_2__1256_ vdd gnd FILL
XFILL_2__1187_ vdd gnd FILL
XFILL_0__789_ vdd gnd FILL
XFILL_0__927_ vdd gnd FILL
XFILL_0__858_ vdd gnd FILL
X_1520_ _1520_/D _1521_/CLK _980_/A vdd gnd DFFPOSX1
X_1382_ _1394_/B _1384_/B _807_/A _1383_/B vdd gnd OAI21X1
XFILL_2_BUFX2_insert3 vdd gnd FILL
X_1451_ _757_/A _985_/A _1451_/C _1521_/D vdd gnd OAI21X1
XFILL_1__1001_ vdd gnd FILL
XFILL_2__1110_ vdd gnd FILL
XFILL_2__1041_ vdd gnd FILL
XFILL_0__1441_ vdd gnd FILL
XFILL_0__1372_ vdd gnd FILL
XFILL_2__1308_ vdd gnd FILL
XFILL_2__1239_ vdd gnd FILL
X_1503_ _1503_/D _1503_/CLK _806_/B vdd gnd DFFPOSX1
X_1365_ _799_/A _1483_/Q _1366_/A vdd gnd NAND2X1
X_1296_ _1331_/B _1296_/B _1298_/B vdd gnd NAND2X1
X_1434_ _1523_/D _728_/B _788_/B _1435_/C vdd gnd OAI21X1
XFILL_2__941_ vdd gnd FILL
XFILL_2__872_ vdd gnd FILL
XFILL_2__1024_ vdd gnd FILL
XFILL_0_CLKBUF1_insert10 vdd gnd FILL
XFILL_1__890_ vdd gnd FILL
X_1150_ _1150_/A _1150_/B _1150_/C _1150_/D _1175_/A vdd gnd AOI22X1
XFILL_0__1355_ vdd gnd FILL
XFILL_0__1424_ vdd gnd FILL
X_1081_ _1081_/A _1081_/B _1130_/A _1085_/B vdd gnd AOI21X1
XFILL_0__1286_ vdd gnd FILL
XFILL_3__1064_ vdd gnd FILL
X_1417_ _1443_/B _1417_/B _1417_/C _1505_/D vdd gnd OAI21X1
XFILL_1__1533_ vdd gnd FILL
X_1348_ _1348_/A _1352_/A _1350_/B vdd gnd XOR2X1
X_1279_ _843_/B _1279_/B _1279_/C _1488_/D vdd gnd OAI21X1
XFILL_1__1395_ vdd gnd FILL
XFILL_2__855_ vdd gnd FILL
XFILL_2__924_ vdd gnd FILL
XFILL_2__786_ vdd gnd FILL
X_930_ _979_/A _985_/B _930_/C _931_/A vdd gnd OAI21X1
X_792_ _817_/A _792_/B _792_/C _792_/Y vdd gnd OAI21X1
X_861_ _980_/A _979_/A vdd gnd INVX2
XFILL_0__1140_ vdd gnd FILL
XFILL_2__1007_ vdd gnd FILL
XFILL_0__1071_ vdd gnd FILL
XFILL_1__942_ vdd gnd FILL
X_1202_ _1202_/A _1202_/B _1202_/C _1221_/B vdd gnd NAND3X1
XFILL86850x150 vdd gnd FILL
X_1064_ _1129_/B _1075_/C _1129_/A _1081_/B vdd gnd NAND3X1
X_1133_ _1133_/A _1133_/B _1133_/C _1134_/A vdd gnd OAI21X1
XFILL_1__873_ vdd gnd FILL
XFILL_0__1338_ vdd gnd FILL
XFILL_0__1407_ vdd gnd FILL
XFILL_1__1180_ vdd gnd FILL
XFILL_0__1269_ vdd gnd FILL
XFILL86550x11850 vdd gnd FILL
XFILL86250x46950 vdd gnd FILL
XFILL_1__1447_ vdd gnd FILL
XFILL_1__1378_ vdd gnd FILL
XFILL_0__960_ vdd gnd FILL
XFILL_2__907_ vdd gnd FILL
XFILL_0__891_ vdd gnd FILL
XFILL_2__838_ vdd gnd FILL
XFILL_2__769_ vdd gnd FILL
X_913_ _913_/A _913_/B _913_/C _915_/B vdd gnd OAI21X1
X_775_ _775_/A _777_/B vdd gnd INVX1
X_844_ _844_/A _844_/B _844_/Y vdd gnd AND2X2
XFILL_0__1054_ vdd gnd FILL
XFILL_0__1123_ vdd gnd FILL
XFILL_1__925_ vdd gnd FILL
XFILL_1__1301_ vdd gnd FILL
XFILL_1__787_ vdd gnd FILL
XFILL_1__856_ vdd gnd FILL
X_1116_ _997_/A Cin[2] _1195_/B vdd gnd NAND2X1
X_1047_ _1047_/A _1051_/B vdd gnd INVX1
XFILL_1__1232_ vdd gnd FILL
XFILL_1__1094_ vdd gnd FILL
XFILL86550x23550 vdd gnd FILL
XFILL_1__1163_ vdd gnd FILL
XFILL_2__1410_ vdd gnd FILL
XFILL_2__1341_ vdd gnd FILL
XFILL_2__1272_ vdd gnd FILL
XFILL_0__943_ vdd gnd FILL
XFILL_0__874_ vdd gnd FILL
XFILL_3__1450_ vdd gnd FILL
X_758_ Xin[0] _765_/B _759_/C vdd gnd NAND2X1
X_827_ _977_/A _834_/A _980_/A _835_/B _859_/B vdd gnd AOI22X1
XFILL_0__1106_ vdd gnd FILL
XFILL_0__1037_ vdd gnd FILL
XFILL_1__908_ vdd gnd FILL
XFILL_1__1215_ vdd gnd FILL
XFILL86550x35250 vdd gnd FILL
XFILL_1__839_ vdd gnd FILL
XFILL_1__1146_ vdd gnd FILL
XFILL_1__1077_ vdd gnd FILL
XFILL_2__1324_ vdd gnd FILL
XFILL_2__1255_ vdd gnd FILL
XFILL_2__1186_ vdd gnd FILL
XFILL_0__926_ vdd gnd FILL
XFILL_0__788_ vdd gnd FILL
XFILL_2_BUFX2_insert4 vdd gnd FILL
X_1450_ _757_/A Xin[3] _1451_/C vdd gnd NAND2X1
XFILL_0__857_ vdd gnd FILL
X_1381_ _1381_/A _1394_/B vdd gnd INVX1
XFILL_3__999_ vdd gnd FILL
XFILL_1__1000_ vdd gnd FILL
XFILL_2__1040_ vdd gnd FILL
XFILL_1__1129_ vdd gnd FILL
XFILL_0__1371_ vdd gnd FILL
XFILL_2__1307_ vdd gnd FILL
XFILL_0__1440_ vdd gnd FILL
XFILL_2__1238_ vdd gnd FILL
XFILL_0__909_ vdd gnd FILL
XFILL_2__1169_ vdd gnd FILL
X_1502_ _1502_/D _1526_/CLK _803_/B vdd gnd DFFPOSX1
X_1433_ _1441_/B _1435_/B _1433_/C _1512_/D vdd gnd OAI21X1
X_1364_ _799_/A _1483_/Q _1367_/A vdd gnd NOR2X1
X_1295_ _1332_/C _1296_/B vdd gnd INVX1
XFILL_2__940_ vdd gnd FILL
XFILL_2__871_ vdd gnd FILL
XFILL_2__1023_ vdd gnd FILL
XFILL_0_CLKBUF1_insert11 vdd gnd FILL
X_1080_ _1106_/B _1130_/C _1106_/A _1085_/A vdd gnd AOI21X1
XFILL_0__1423_ vdd gnd FILL
XFILL_0__1354_ vdd gnd FILL
XFILL_3__1132_ vdd gnd FILL
XFILL_0__1285_ vdd gnd FILL
X_1347_ _1347_/A _1352_/A vdd gnd INVX1
X_1416_ _812_/B _1417_/B _1417_/C vdd gnd NAND2X1
XFILL_1__1532_ vdd gnd FILL
XFILL_1__1394_ vdd gnd FILL
X_1278_ _740_/B _1370_/A _1279_/C vdd gnd NAND2X1
XFILL_2__854_ vdd gnd FILL
XFILL_2__923_ vdd gnd FILL
XFILL_2__785_ vdd gnd FILL
X_791_ _817_/A _791_/B _792_/C vdd gnd NAND2X1
X_860_ _881_/C _893_/B _893_/A _871_/A vdd gnd AOI21X1
XFILL_2__1006_ vdd gnd FILL
XFILL_0__1070_ vdd gnd FILL
X_1201_ _1202_/A _1202_/B _1202_/C _1221_/C vdd gnd AOI21X1
XFILL_1__941_ vdd gnd FILL
XFILL_1__872_ vdd gnd FILL
X_989_ _989_/A _989_/B _989_/C _989_/Y vdd gnd AOI21X1
X_1063_ _1113_/A _1113_/B _1120_/C _1129_/B vdd gnd NAND3X1
X_1132_ _1132_/A _1132_/B _1134_/B vdd gnd NAND2X1
XFILL_0__1337_ vdd gnd FILL
XFILL_0__1268_ vdd gnd FILL
XFILL_0__1406_ vdd gnd FILL
XFILL_0__1199_ vdd gnd FILL
XFILL_1__1377_ vdd gnd FILL
XFILL_1__1446_ vdd gnd FILL
XFILL_2__768_ vdd gnd FILL
XFILL_0__890_ vdd gnd FILL
XFILL_2__906_ vdd gnd FILL
XFILL_2__837_ vdd gnd FILL
X_843_ _843_/A _843_/B _844_/B vdd gnd NAND2X1
X_912_ _912_/A _913_/B vdd gnd INVX1
X_774_ _786_/A _774_/B _774_/C _774_/Y vdd gnd OAI21X1
XFILL_0__1122_ vdd gnd FILL
XFILL_3_BUFX2_insert26 vdd gnd FILL
XFILL_0__1053_ vdd gnd FILL
XFILL_1__855_ vdd gnd FILL
XFILL_1__924_ vdd gnd FILL
XFILL_1__1300_ vdd gnd FILL
XFILL_1__1231_ vdd gnd FILL
XFILL_1__786_ vdd gnd FILL
X_1046_ _1047_/A _1046_/B _1046_/C _1073_/A vdd gnd NAND3X1
X_1115_ _755_/A Cin[2] _1165_/A vdd gnd NAND2X1
XFILL_1__1093_ vdd gnd FILL
XFILL_1__1162_ vdd gnd FILL
XFILL_2__1340_ vdd gnd FILL
XFILL_2__1271_ vdd gnd FILL
XFILL_1__1429_ vdd gnd FILL
XFILL_0__942_ vdd gnd FILL
XFILL_0__873_ vdd gnd FILL
X_826_ _826_/A _850_/A _847_/C vdd gnd NOR2X1
X_757_ _757_/A _765_/A _757_/C _757_/Y vdd gnd OAI21X1
XFILL_0__1105_ vdd gnd FILL
XFILL_0__1036_ vdd gnd FILL
XFILL_1__907_ vdd gnd FILL
XFILL_1__838_ vdd gnd FILL
XFILL_1__769_ vdd gnd FILL
XFILL_1__1214_ vdd gnd FILL
X_1029_ _1029_/A _1029_/B _974_/Y _1030_/B vdd gnd AOI21X1
XFILL_1__1145_ vdd gnd FILL
XFILL_1__1076_ vdd gnd FILL
XFILL_2__1323_ vdd gnd FILL
XFILL_2__1185_ vdd gnd FILL
XFILL_2__1254_ vdd gnd FILL
XFILL_0__925_ vdd gnd FILL
X_1380_ _1395_/A _1384_/B vdd gnd INVX1
XFILL_2_BUFX2_insert5 vdd gnd FILL
XFILL_0__787_ vdd gnd FILL
XFILL_0__856_ vdd gnd FILL
X_809_ _813_/A _809_/B _810_/C vdd gnd NAND2X1
XFILL_0__1019_ vdd gnd FILL
XFILL_1__1128_ vdd gnd FILL
XFILL_1__1059_ vdd gnd FILL
XFILL_2__1237_ vdd gnd FILL
XFILL_0__1370_ vdd gnd FILL
XFILL_2__1306_ vdd gnd FILL
XFILL_2__1099_ vdd gnd FILL
XFILL_2__1168_ vdd gnd FILL
XFILL_0__908_ vdd gnd FILL
XFILL_0__839_ vdd gnd FILL
X_1363_ _1372_/B _1363_/B _1368_/A vdd gnd NOR2X1
X_1501_ _1501_/D _1508_/CLK _742_/B vdd gnd DFFPOSX1
X_1432_ _1523_/D _728_/B _785_/B _1433_/C vdd gnd OAI21X1
X_1294_ _1294_/A _1294_/B _1294_/C _1332_/C vdd gnd OAI21X1
XFILL_2__870_ vdd gnd FILL
XFILL_2__1022_ vdd gnd FILL
XFILL_2__999_ vdd gnd FILL
XFILL85650x23550 vdd gnd FILL
XFILL_0_CLKBUF1_insert12 vdd gnd FILL
XFILL_3__1200_ vdd gnd FILL
XFILL_0__1353_ vdd gnd FILL
XFILL_0__1422_ vdd gnd FILL
XFILL_0__1284_ vdd gnd FILL
X_1415_ Yin[3] _1443_/B vdd gnd INVX1
X_1346_ _1353_/B _1346_/B _1347_/A vdd gnd NOR2X1
XFILL_1__1531_ vdd gnd FILL
XFILL_1__1393_ vdd gnd FILL
X_1277_ _1281_/A _1281_/B _1279_/B vdd gnd XNOR2X1
XFILL_3__1329_ vdd gnd FILL
XFILL_2__922_ vdd gnd FILL
XFILL_2__784_ vdd gnd FILL
XFILL_2__853_ vdd gnd FILL
X_790_ _790_/A _792_/B vdd gnd INVX1
XFILL_2__1005_ vdd gnd FILL
X_1200_ _1223_/D _1222_/A _1202_/C vdd gnd XOR2X1
XFILL_1__940_ vdd gnd FILL
X_988_ _988_/A _988_/B _989_/C vdd gnd NOR2X1
XFILL_1__871_ vdd gnd FILL
XFILL_3__818_ vdd gnd FILL
XFILL_0__1405_ vdd gnd FILL
X_1131_ _1152_/C _1168_/B _1168_/A _1138_/A vdd gnd AOI21X1
X_1062_ _1120_/B _1113_/B vdd gnd INVX1
XFILL_0__1336_ vdd gnd FILL
XFILL_0__1267_ vdd gnd FILL
XFILL_0__1198_ vdd gnd FILL
X_1329_ _1329_/A _1329_/B _1332_/B vdd gnd AND2X2
XFILL_1__1376_ vdd gnd FILL
XFILL_1__1445_ vdd gnd FILL
XFILL_2__905_ vdd gnd FILL
XFILL_2__767_ vdd gnd FILL
XFILL_2__836_ vdd gnd FILL
X_842_ _842_/A _843_/A vdd gnd INVX1
X_911_ _921_/A _955_/C _921_/B _913_/A vdd gnd AOI21X1
X_773_ _815_/C _773_/B _774_/C vdd gnd NAND2X1
XFILL_0__1052_ vdd gnd FILL
XFILL_0__1121_ vdd gnd FILL
XFILL87150x54750 vdd gnd FILL
XFILL_1__785_ vdd gnd FILL
XFILL_1__854_ vdd gnd FILL
X_1114_ _997_/A _997_/B _1118_/A vdd gnd NAND2X1
XFILL_1__923_ vdd gnd FILL
XFILL_1__1230_ vdd gnd FILL
XFILL_1__1161_ vdd gnd FILL
X_1045_ _759_/A _985_/B _1048_/A _1046_/C vdd gnd OAI21X1
XFILL_0__1319_ vdd gnd FILL
XFILL_1__1092_ vdd gnd FILL
XFILL_2__1270_ vdd gnd FILL
XFILL_1__1359_ vdd gnd FILL
XFILL_1__1428_ vdd gnd FILL
XFILL_0__941_ vdd gnd FILL
XFILL_0__872_ vdd gnd FILL
XFILL_2__819_ vdd gnd FILL
X_825_ _980_/A _834_/A _850_/A vdd gnd NAND2X1
X_756_ _757_/A _978_/A _757_/C vdd gnd NAND2X1
XFILL_2__1399_ vdd gnd FILL
XFILL_0__1104_ vdd gnd FILL
XFILL_0__1035_ vdd gnd FILL
XFILL87150x66450 vdd gnd FILL
XFILL_1__768_ vdd gnd FILL
XFILL_1__906_ vdd gnd FILL
XFILL_1__837_ vdd gnd FILL
XFILL_1__1213_ vdd gnd FILL
X_1028_ _1036_/B _1089_/C _974_/A _1030_/A vdd gnd AOI21X1
XFILL_1__1144_ vdd gnd FILL
XFILL_1__1075_ vdd gnd FILL
XFILL_2__1253_ vdd gnd FILL
XFILL_2__1322_ vdd gnd FILL
XFILL_2__1184_ vdd gnd FILL
XFILL_0__855_ vdd gnd FILL
XFILL_0__924_ vdd gnd FILL
XFILL_2_BUFX2_insert6 vdd gnd FILL
XFILL_0__786_ vdd gnd FILL
X_808_ _808_/A _810_/B vdd gnd INVX1
X_739_ _743_/A _739_/B _739_/C _741_/B vdd gnd OAI21X1
XFILL87150x78150 vdd gnd FILL
XFILL_0__1018_ vdd gnd FILL
XFILL_1__1127_ vdd gnd FILL
XFILL_1__1058_ vdd gnd FILL
XFILL_2__1236_ vdd gnd FILL
XFILL_2__1305_ vdd gnd FILL
XFILL_2__1167_ vdd gnd FILL
XFILL_0__769_ vdd gnd FILL
X_1500_ _1500_/D _1508_/CLK _737_/A vdd gnd DFFPOSX1
XFILL_2__1098_ vdd gnd FILL
XFILL_0__907_ vdd gnd FILL
XFILL_0__838_ vdd gnd FILL
X_1362_ _1362_/A _1374_/B _1363_/B vdd gnd NOR2X1
X_1431_ _1439_/B _1435_/B _1431_/C _1511_/D vdd gnd OAI21X1
X_1293_ _1293_/A _1294_/C vdd gnd INVX1
XFILL_3__1276_ vdd gnd FILL
XFILL_2__1021_ vdd gnd FILL
XFILL_2__998_ vdd gnd FILL
XFILL_0_CLKBUF1_insert13 vdd gnd FILL
XFILL_0__1421_ vdd gnd FILL
XFILL_3__765_ vdd gnd FILL
XFILL_0__1352_ vdd gnd FILL
XFILL_2__1219_ vdd gnd FILL
XFILL_0__1283_ vdd gnd FILL
X_1345_ _1353_/C _1346_/B vdd gnd INVX1
X_1414_ _1441_/B _1417_/B _1414_/C _1504_/D vdd gnd OAI21X1
X_1276_ _772_/A _842_/A _1281_/B vdd gnd XOR2X1
XFILL_1__1530_ vdd gnd FILL
XFILL_1__1392_ vdd gnd FILL
XFILL_2__921_ vdd gnd FILL
XFILL_2__783_ vdd gnd FILL
XFILL_2__852_ vdd gnd FILL
XFILL_2__1004_ vdd gnd FILL
X_1130_ _1130_/A _1130_/B _1130_/C _1178_/C vdd gnd OAI21X1
X_987_ _987_/A _987_/B _987_/Y vdd gnd NAND2X1
XFILL_1__870_ vdd gnd FILL
XFILL_0__1335_ vdd gnd FILL
XFILL_0__1404_ vdd gnd FILL
X_1061_ _998_/B _1068_/C _1120_/C vdd gnd NAND2X1
XFILL_0__1266_ vdd gnd FILL
XFILL_0__1197_ vdd gnd FILL
X_1259_ _1386_/B _1391_/B _1259_/C _1259_/D _1485_/D vdd gnd AOI22X1
X_1328_ _1328_/A _1328_/B _1328_/C _1330_/C vdd gnd OAI21X1
XFILL_1__1444_ vdd gnd FILL
XFILL_1__999_ vdd gnd FILL
XFILL_1__1375_ vdd gnd FILL
XFILL_2__904_ vdd gnd FILL
XFILL_2__835_ vdd gnd FILL
XFILL_2__766_ vdd gnd FILL
X_772_ _772_/A _774_/B vdd gnd INVX1
X_910_ _919_/B _910_/B _910_/C _913_/C vdd gnd AOI21X1
X_841_ _841_/A _874_/A _917_/B _844_/A vdd gnd OAI21X1
XFILL_0__1120_ vdd gnd FILL
XFILL_0__1051_ vdd gnd FILL
XFILL_1__922_ vdd gnd FILL
XFILL_1__784_ vdd gnd FILL
X_1113_ _1113_/A _1113_/B _1133_/A _1132_/B vdd gnd AOI21X1
XFILL_1__853_ vdd gnd FILL
X_1044_ _978_/A Cin[4] _1048_/A vdd gnd AND2X2
XFILL_1__1160_ vdd gnd FILL
XFILL_0__1318_ vdd gnd FILL
XFILL_1__1091_ vdd gnd FILL
XFILL_0__1249_ vdd gnd FILL
XFILL_1__1427_ vdd gnd FILL
XFILL_1__1358_ vdd gnd FILL
XFILL_1__1289_ vdd gnd FILL
XFILL_0__940_ vdd gnd FILL
XFILL_0__871_ vdd gnd FILL
XFILL_2__818_ vdd gnd FILL
XFILL_2__749_ vdd gnd FILL
X_755_ _755_/A _765_/A vdd gnd INVX2
X_824_ _922_/A Cin[2] _859_/A vdd gnd NAND2X1
XFILL_2__1398_ vdd gnd FILL
XFILL_0__1034_ vdd gnd FILL
XFILL_0__1103_ vdd gnd FILL
XFILL_1__905_ vdd gnd FILL
XFILL_1__767_ vdd gnd FILL
X_1027_ _959_/A _962_/C _1027_/C _1034_/A vdd gnd AOI21X1
XFILL_1__836_ vdd gnd FILL
XFILL_1__1143_ vdd gnd FILL
XFILL_1__1212_ vdd gnd FILL
XFILL_1__1074_ vdd gnd FILL
XFILL_2__1183_ vdd gnd FILL
XFILL_2__1252_ vdd gnd FILL
XFILL_2__1321_ vdd gnd FILL
XFILL_0__785_ vdd gnd FILL
XFILL_0__854_ vdd gnd FILL
XFILL_0__923_ vdd gnd FILL
X_807_ _807_/A _807_/B _807_/C _807_/Y vdd gnd OAI21X1
X_738_ _743_/A _738_/B _739_/C vdd gnd NAND2X1
XFILL_0__1017_ vdd gnd FILL
XFILL_1__819_ vdd gnd FILL
XFILL_1__1126_ vdd gnd FILL
XFILL_1__1057_ vdd gnd FILL
XFILL_2__1304_ vdd gnd FILL
XFILL_2__1235_ vdd gnd FILL
XFILL_0__906_ vdd gnd FILL
XFILL_2__1166_ vdd gnd FILL
XFILL_2__1097_ vdd gnd FILL
XFILL_0__768_ vdd gnd FILL
X_1430_ _1523_/D _728_/B _782_/B _1431_/C vdd gnd OAI21X1
XFILL_0__837_ vdd gnd FILL
X_1361_ _1361_/A _1361_/B _1361_/C _1496_/D vdd gnd OAI21X1
X_1292_ _1297_/A _1331_/B vdd gnd INVX1
XFILL_3__1344_ vdd gnd FILL
XFILL_2_BUFX2_insert30 vdd gnd FILL
XFILL_2__1020_ vdd gnd FILL
XFILL_2__997_ vdd gnd FILL
XFILL_1__1109_ vdd gnd FILL
XFILL_0_CLKBUF1_insert14 vdd gnd FILL
XFILL_3__833_ vdd gnd FILL
XFILL_0__1420_ vdd gnd FILL
XFILL_0__1351_ vdd gnd FILL
XFILL_2__1218_ vdd gnd FILL
XFILL_2__1149_ vdd gnd FILL
XFILL_0__1282_ vdd gnd FILL
X_1413_ _809_/B _1417_/B _1414_/C vdd gnd NAND2X1
X_1275_ _771_/B _1275_/B _1275_/C _1281_/A vdd gnd OAI21X1
X_1344_ _793_/A _1481_/Q _1353_/C vdd gnd NAND2X1
XFILL_1__1391_ vdd gnd FILL
XFILL_2__920_ vdd gnd FILL
XFILL_2__851_ vdd gnd FILL
XFILL_2__782_ vdd gnd FILL
XFILL86250x66450 vdd gnd FILL
XFILL_2__1003_ vdd gnd FILL
X_1060_ _755_/A _993_/B _1068_/C vdd gnd AND2X2
X_986_ _986_/A _986_/B _986_/C _987_/A vdd gnd NAND3X1
XFILL_0__1334_ vdd gnd FILL
XFILL_0__1403_ vdd gnd FILL
XFILL_0__1265_ vdd gnd FILL
XFILL_0__1196_ vdd gnd FILL
X_1258_ _1258_/A _812_/A _1259_/D vdd gnd AND2X2
X_1189_ _1189_/A _1189_/B _1251_/A vdd gnd NAND2X1
XFILL_1__1443_ vdd gnd FILL
X_1327_ _784_/A _968_/A _1328_/A vdd gnd NAND2X1
XFILL_1__998_ vdd gnd FILL
XFILL_1__1374_ vdd gnd FILL
XFILL_2__903_ vdd gnd FILL
XFILL_2__834_ vdd gnd FILL
XFILL86250x78150 vdd gnd FILL
XFILL_2__765_ vdd gnd FILL
X_771_ _817_/A _771_/B _771_/C _771_/Y vdd gnd OAI21X1
X_840_ _840_/A _840_/B _840_/C _841_/A vdd gnd AOI21X1
XFILL_0__1050_ vdd gnd FILL
XFILL_3_BUFX2_insert18 vdd gnd FILL
XFILL_1__921_ vdd gnd FILL
XFILL_1__852_ vdd gnd FILL
XFILL_1__783_ vdd gnd FILL
X_969_ _969_/A _969_/B _969_/C _969_/D _969_/Y vdd gnd AOI22X1
X_1112_ _1150_/C _1150_/D _1152_/B vdd gnd XNOR2X1
X_1043_ _985_/A _979_/B _1150_/A _1046_/B vdd gnd OAI21X1
XFILL_0__1248_ vdd gnd FILL
XFILL_0__1317_ vdd gnd FILL
XFILL_1__1090_ vdd gnd FILL
XFILL_3__1026_ vdd gnd FILL
XFILL_0__1179_ vdd gnd FILL
XFILL_1__1357_ vdd gnd FILL
XFILL_1__1426_ vdd gnd FILL
XFILL_1__1288_ vdd gnd FILL
XFILL_2__817_ vdd gnd FILL
XFILL_0__870_ vdd gnd FILL
XFILL_2__748_ vdd gnd FILL
X_823_ _823_/A _826_/A _840_/C vdd gnd NOR2X1
XFILL_2__1535_ vdd gnd FILL
X_754_ _757_/A _999_/A _754_/C _754_/Y vdd gnd OAI21X1
XFILL_2__1397_ vdd gnd FILL
XFILL_0__1102_ vdd gnd FILL
XFILL_0__1033_ vdd gnd FILL
XFILL_0__999_ vdd gnd FILL
XFILL_1__904_ vdd gnd FILL
XFILL_1__835_ vdd gnd FILL
XFILL_1__1211_ vdd gnd FILL
XFILL_1__766_ vdd gnd FILL
X_1026_ _971_/C _1027_/C vdd gnd INVX1
XFILL_1__1073_ vdd gnd FILL
XFILL_1__1142_ vdd gnd FILL
XFILL_2__1320_ vdd gnd FILL
XFILL_1__1409_ vdd gnd FILL
XFILL_2__1251_ vdd gnd FILL
XFILL_2__1182_ vdd gnd FILL
XFILL_0__922_ vdd gnd FILL
XFILL_0__784_ vdd gnd FILL
XFILL_0__853_ vdd gnd FILL
X_806_ _807_/A _806_/B _807_/C vdd gnd NAND2X1
X_737_ _737_/A _738_/B vdd gnd INVX1
XFILL_3__1291_ vdd gnd FILL
XFILL_2__1449_ vdd gnd FILL
XFILL_0__1016_ vdd gnd FILL
XFILL_1__818_ vdd gnd FILL
X_1009_ _995_/Y _1078_/C _1078_/A _1079_/C vdd gnd NAND3X1
XFILL_1__749_ vdd gnd FILL
XFILL_1__1056_ vdd gnd FILL
XFILL_1__1125_ vdd gnd FILL
XFILL_3__780_ vdd gnd FILL
XFILL_2__1303_ vdd gnd FILL
XFILL_2__1234_ vdd gnd FILL
XFILL_2__1096_ vdd gnd FILL
XFILL_0__905_ vdd gnd FILL
XFILL_2__1165_ vdd gnd FILL
X_1360_ _1362_/A _1374_/B _813_/A _1361_/A vdd gnd OAI21X1
XFILL_0__767_ vdd gnd FILL
XFILL_0__836_ vdd gnd FILL
XFILL_3__1412_ vdd gnd FILL
X_1291_ _1291_/A _1326_/A _1297_/A vdd gnd AND2X2
XFILL_2_BUFX2_insert20 vdd gnd FILL
X_1489_ _1489_/D _1522_/CLK _744_/B vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert31 vdd gnd FILL
XFILL_2__996_ vdd gnd FILL
XFILL_1__1108_ vdd gnd FILL
XFILL_1__1039_ vdd gnd FILL
XFILL_3__901_ vdd gnd FILL
XFILL_0__1350_ vdd gnd FILL
XFILL_2__1217_ vdd gnd FILL
XFILL_0__1281_ vdd gnd FILL
XFILL_2__1148_ vdd gnd FILL
XFILL_2__1079_ vdd gnd FILL
XFILL_0__819_ vdd gnd FILL
X_1412_ Yin[2] _1441_/B vdd gnd INVX1
X_1343_ _793_/A _1481_/Q _1353_/B vdd gnd NOR2X1
XFILL_1__1390_ vdd gnd FILL
X_1274_ _1350_/A _1274_/B _1274_/C _1487_/D vdd gnd OAI21X1
XFILL_2__781_ vdd gnd FILL
XFILL_2__850_ vdd gnd FILL
XFILL_2__1002_ vdd gnd FILL
XFILL_2__979_ vdd gnd FILL
X_985_ _985_/A _985_/B _985_/C _986_/A vdd gnd OAI21X1
XFILL_0__1402_ vdd gnd FILL
XFILL_0__1264_ vdd gnd FILL
XFILL_0__1333_ vdd gnd FILL
XFILL_0__1195_ vdd gnd FILL
X_1326_ _1326_/A _1331_/A _1326_/C _1330_/A vdd gnd OAI21X1
XFILL_1__997_ vdd gnd FILL
XFILL_1__1373_ vdd gnd FILL
X_1257_ _1257_/A _1257_/B _1257_/C _1259_/C vdd gnd AOI21X1
X_1188_ _1188_/A _1214_/A _1189_/B vdd gnd NAND2X1
XFILL_1__1442_ vdd gnd FILL
XFILL86850x27450 vdd gnd FILL
XFILL_2__764_ vdd gnd FILL
XFILL_2__902_ vdd gnd FILL
XFILL_2__833_ vdd gnd FILL
X_770_ _817_/A _770_/B _771_/C vdd gnd NAND2X1
X_968_ _968_/A _968_/Y vdd gnd INVX1
XFILL_1__920_ vdd gnd FILL
XFILL_1__851_ vdd gnd FILL
XFILL_1__782_ vdd gnd FILL
X_899_ Cin[4] _979_/B vdd gnd INVX2
X_1111_ _1150_/A _1150_/B _1111_/C _1150_/C vdd gnd AOI21X1
X_1042_ _990_/A Cin[3] _1150_/A vdd gnd AND2X2
XFILL_0__1316_ vdd gnd FILL
XFILL_0__1247_ vdd gnd FILL
XFILL_0__1178_ vdd gnd FILL
X_1309_ _1309_/A _1309_/B _1309_/C _1491_/D vdd gnd OAI21X1
XFILL86850x39150 vdd gnd FILL
XFILL_1__1356_ vdd gnd FILL
XFILL_1__1425_ vdd gnd FILL
XFILL_1__1287_ vdd gnd FILL
XFILL_2__816_ vdd gnd FILL
XFILL_2__747_ vdd gnd FILL
X_822_ _967_/A _822_/B _822_/C _822_/Y vdd gnd OAI21X1
XFILL_2__1534_ vdd gnd FILL
XFILL_2__1396_ vdd gnd FILL
X_753_ _757_/A _980_/A _754_/C vdd gnd NAND2X1
XFILL_0__1032_ vdd gnd FILL
XFILL_0__1101_ vdd gnd FILL
XFILL_0__998_ vdd gnd FILL
XFILL_1__765_ vdd gnd FILL
XFILL_1__903_ vdd gnd FILL
XFILL_1__834_ vdd gnd FILL
XFILL_1__1210_ vdd gnd FILL
XFILL_1__1141_ vdd gnd FILL
X_1025_ _1025_/A _1025_/B _971_/Y _1098_/B vdd gnd NAND3X1
XFILL_1__1072_ vdd gnd FILL
XFILL_2__1250_ vdd gnd FILL
XFILL_1__1339_ vdd gnd FILL
XFILL_1__1408_ vdd gnd FILL
XFILL_2__1181_ vdd gnd FILL
XFILL_0__921_ vdd gnd FILL
XFILL_0__852_ vdd gnd FILL
XFILL_0__783_ vdd gnd FILL
X_736_ _741_/A _736_/B _736_/C _736_/Y vdd gnd OAI21X1
X_805_ _805_/A _807_/B vdd gnd INVX1
XFILL_2__1379_ vdd gnd FILL
XFILL_2__1448_ vdd gnd FILL
XFILL_0__1015_ vdd gnd FILL
XFILL_1__817_ vdd gnd FILL
XFILL_1__748_ vdd gnd FILL
X_1008_ _987_/B _987_/A _1040_/A vdd gnd AND2X2
XFILL_1__1124_ vdd gnd FILL
XFILL_1__1055_ vdd gnd FILL
XFILL_2__1302_ vdd gnd FILL
XFILL_2__1233_ vdd gnd FILL
XFILL_2__1095_ vdd gnd FILL
XFILL_0__904_ vdd gnd FILL
XFILL_2__1164_ vdd gnd FILL
XFILL_0__835_ vdd gnd FILL
XFILL_0__766_ vdd gnd FILL
XFILL_3__977_ vdd gnd FILL
X_1290_ _778_/A _877_/A _1326_/A vdd gnd NAND2X1
XFILL87150x50850 vdd gnd FILL
X_1488_ _1488_/D _1525_/CLK _740_/B vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert21 vdd gnd FILL
XFILL_2_BUFX2_insert32 vdd gnd FILL
XFILL_2__995_ vdd gnd FILL
XFILL_1__1107_ vdd gnd FILL
XFILL_1__1038_ vdd gnd FILL
XFILL_2__1216_ vdd gnd FILL
XFILL_0__1280_ vdd gnd FILL
XFILL_2__1147_ vdd gnd FILL
XFILL_2__1078_ vdd gnd FILL
XFILL_0__818_ vdd gnd FILL
X_1273_ _735_/B _1350_/A _1274_/C vdd gnd NAND2X1
X_1342_ _1352_/B _1342_/B _1353_/A _1348_/A vdd gnd OAI21X1
X_1411_ _1439_/B _1417_/B _1411_/C _1503_/D vdd gnd OAI21X1
XFILL_0__749_ vdd gnd FILL
XFILL_2__780_ vdd gnd FILL
XFILL_2__1001_ vdd gnd FILL
XFILL_2__978_ vdd gnd FILL
X_984_ _984_/A _984_/B _986_/C vdd gnd NAND2X1
XFILL_0__1401_ vdd gnd FILL
XFILL_0__1263_ vdd gnd FILL
XFILL_0__1332_ vdd gnd FILL
XFILL_0__1194_ vdd gnd FILL
XFILL_3__1041_ vdd gnd FILL
XFILL87150x74250 vdd gnd FILL
X_1325_ _726_/B _1350_/A _1341_/C vdd gnd NAND2X1
X_1256_ _1485_/Q _1386_/B vdd gnd INVX1
XFILL_1__996_ vdd gnd FILL
XFILL_1__1372_ vdd gnd FILL
XFILL_1__1441_ vdd gnd FILL
X_1187_ _1187_/A _1187_/B _1191_/B vdd gnd NOR2X1
XFILL_2__901_ vdd gnd FILL
XFILL_2__763_ vdd gnd FILL
XFILL_2__832_ vdd gnd FILL
XFILL_1__781_ vdd gnd FILL
X_967_ _967_/A _967_/B _967_/C _967_/Y vdd gnd OAI21X1
X_898_ _922_/A _901_/A vdd gnd INVX1
XFILL_1__850_ vdd gnd FILL
X_1110_ _990_/A Cin[4] _994_/A Cin[3] _1111_/C vdd gnd AOI22X1
X_1041_ _980_/A Cin[5] _1047_/A vdd gnd NAND2X1
XFILL_0__1246_ vdd gnd FILL
XFILL_0__1315_ vdd gnd FILL
XFILL_0__1177_ vdd gnd FILL
XFILL_1__1424_ vdd gnd FILL
X_1308_ _1331_/A _1311_/B _817_/A _1309_/B vdd gnd OAI21X1
X_1239_ _1239_/A _1239_/B _1241_/A _1240_/B vdd gnd AOI21X1
XFILL_1__979_ vdd gnd FILL
XFILL_1__1355_ vdd gnd FILL
XFILL_1__1286_ vdd gnd FILL
XFILL_2__815_ vdd gnd FILL
XFILL_2__746_ vdd gnd FILL
XFILL_2__1533_ vdd gnd FILL
X_821_ _821_/A _967_/A _822_/C vdd gnd NAND2X1
X_752_ _997_/A _999_/A vdd gnd INVX2
XFILL_2__1395_ vdd gnd FILL
XFILL_0__1031_ vdd gnd FILL
XFILL_0__997_ vdd gnd FILL
XFILL_0__1100_ vdd gnd FILL
XFILL_1__902_ vdd gnd FILL
XFILL_1__764_ vdd gnd FILL
X_1024_ _969_/Y _1213_/C _1033_/D vdd gnd NOR2X1
XFILL_1__833_ vdd gnd FILL
XFILL_1__1140_ vdd gnd FILL
XFILL_0__1229_ vdd gnd FILL
XFILL_1__1071_ vdd gnd FILL
XFILL_1__1407_ vdd gnd FILL
XFILL_2__1180_ vdd gnd FILL
XFILL_1__1338_ vdd gnd FILL
XFILL_1__1269_ vdd gnd FILL
XFILL_0__782_ vdd gnd FILL
XFILL_0__920_ vdd gnd FILL
XFILL_0__851_ vdd gnd FILL
XFILL_2__729_ vdd gnd FILL
X_804_ _807_/A _804_/B _804_/C _804_/Y vdd gnd OAI21X1
X_735_ _744_/A _735_/B _765_/B _735_/D _736_/C vdd gnd AOI22X1
XFILL_2__1378_ vdd gnd FILL
XFILL_2__1447_ vdd gnd FILL
XFILL_0__1014_ vdd gnd FILL
XFILL_1__816_ vdd gnd FILL
X_1007_ _987_/Y _1016_/B _1016_/A _1088_/B vdd gnd NAND3X1
XFILL_1__747_ vdd gnd FILL
XFILL_1__1054_ vdd gnd FILL
XFILL_1__1123_ vdd gnd FILL
XFILL_2__1232_ vdd gnd FILL
XFILL_2__1301_ vdd gnd FILL
XFILL_2__1163_ vdd gnd FILL
XFILL85950x27450 vdd gnd FILL
XFILL_0__765_ vdd gnd FILL
XFILL_0__903_ vdd gnd FILL
XFILL_2__1094_ vdd gnd FILL
XFILL_0__834_ vdd gnd FILL
XFILL_2_BUFX2_insert22 vdd gnd FILL
XFILL_2_BUFX2_insert33 vdd gnd FILL
X_1487_ _1487_/D _1515_/CLK _735_/B vdd gnd DFFPOSX1
XFILL_2__994_ vdd gnd FILL
XFILL_1__1106_ vdd gnd FILL
XFILL_1__1037_ vdd gnd FILL
XFILL_2__1146_ vdd gnd FILL
XFILL_2__1215_ vdd gnd FILL
X_1410_ _806_/B _1417_/B _1411_/C vdd gnd NAND2X1
XFILL_0__817_ vdd gnd FILL
XFILL_2__1077_ vdd gnd FILL
XFILL_0__748_ vdd gnd FILL
X_1341_ _1341_/A _1341_/B _1341_/C _1494_/D vdd gnd OAI21X1
X_1272_ _1272_/A _1275_/C _1274_/B vdd gnd NAND2X1
XFILL_2__1000_ vdd gnd FILL
XFILL_2__977_ vdd gnd FILL
X_983_ _983_/A _986_/B vdd gnd INVX1
XFILL_0__1400_ vdd gnd FILL
XFILL_0__1331_ vdd gnd FILL
XFILL_0__1262_ vdd gnd FILL
XFILL_0__1193_ vdd gnd FILL
XFILL_2__1129_ vdd gnd FILL
X_1255_ _1376_/B _807_/A _1255_/C _1255_/D _1484_/D vdd gnd OAI22X1
X_1324_ _1370_/A _1324_/B _1324_/C _1493_/D vdd gnd OAI21X1
XFILL_1__1440_ vdd gnd FILL
X_1186_ _1188_/A _1189_/A _1187_/A vdd gnd NAND2X1
XFILL_1__995_ vdd gnd FILL
XFILL_1__1371_ vdd gnd FILL
XFILL_3__1238_ vdd gnd FILL
XFILL_0__1529_ vdd gnd FILL
XFILL_2__900_ vdd gnd FILL
XFILL_2__831_ vdd gnd FILL
XFILL_2__762_ vdd gnd FILL
X_966_ _966_/A _967_/A _967_/C vdd gnd NAND2X1
XFILL_3__727_ vdd gnd FILL
XFILL_1__780_ vdd gnd FILL
X_1040_ _1040_/A _1040_/B _1040_/C _1085_/C vdd gnd AOI21X1
X_897_ _977_/A Cin[4] _930_/C vdd gnd NAND2X1
XFILL_0__1314_ vdd gnd FILL
XFILL_0__1245_ vdd gnd FILL
XFILL_0__1176_ vdd gnd FILL
XFILL_1__1423_ vdd gnd FILL
X_1307_ _1307_/A _1331_/A vdd gnd INVX1
X_1238_ _1239_/A _1239_/B _1240_/A vdd gnd NOR2X1
XFILL_1__978_ vdd gnd FILL
X_1169_ _1169_/A _1193_/C _1169_/C _1174_/A vdd gnd AOI21X1
XFILL_1__1354_ vdd gnd FILL
XFILL_1__1285_ vdd gnd FILL
XFILL_2__814_ vdd gnd FILL
XFILL_2__745_ vdd gnd FILL
XFILL_2__1532_ vdd gnd FILL
X_820_ _823_/A _826_/A _822_/B vdd gnd XNOR2X1
X_751_ _751_/A _943_/A _751_/C _751_/Y vdd gnd OAI21X1
XFILL_2__1394_ vdd gnd FILL
XFILL_0__1030_ vdd gnd FILL
XFILL_0__996_ vdd gnd FILL
XFILL_1__832_ vdd gnd FILL
XFILL_1__901_ vdd gnd FILL
XFILL_1__763_ vdd gnd FILL
X_949_ _957_/C _957_/B _957_/A _970_/A vdd gnd NAND3X1
X_1023_ _1034_/B _971_/Y _1213_/C vdd gnd XNOR2X1
XFILL_0__1228_ vdd gnd FILL
XFILL_1__1070_ vdd gnd FILL
XFILL_0__1159_ vdd gnd FILL
XFILL_1__1337_ vdd gnd FILL
XFILL_1__1406_ vdd gnd FILL
XFILL_1__1268_ vdd gnd FILL
XFILL_0__781_ vdd gnd FILL
XFILL_2__728_ vdd gnd FILL
XFILL_1__1199_ vdd gnd FILL
XFILL_0__850_ vdd gnd FILL
XFILL_3__992_ vdd gnd FILL
X_734_ _743_/A _734_/B _734_/C _736_/B vdd gnd OAI21X1
X_803_ _807_/A _803_/B _804_/C vdd gnd NAND2X1
XFILL_2__1446_ vdd gnd FILL
XFILL_2__1377_ vdd gnd FILL
XFILL_0__1013_ vdd gnd FILL
XFILL_0__979_ vdd gnd FILL
XFILL_1__815_ vdd gnd FILL
X_1006_ _1010_/A _1010_/B _1078_/C _1016_/A vdd gnd OAI21X1
XFILL_1__746_ vdd gnd FILL
XFILL_1__1053_ vdd gnd FILL
XFILL_1__1122_ vdd gnd FILL
XFILL86250x74250 vdd gnd FILL
XFILL_2__1300_ vdd gnd FILL
XFILL_2__1231_ vdd gnd FILL
XFILL_2__1093_ vdd gnd FILL
XFILL_0__902_ vdd gnd FILL
XFILL_2__1162_ vdd gnd FILL
XFILL_0__764_ vdd gnd FILL
XFILL_0__833_ vdd gnd FILL
XFILL_2__1429_ vdd gnd FILL
XFILL_2_BUFX2_insert23 vdd gnd FILL
X_1486_ _1486_/D _1515_/CLK _729_/B vdd gnd DFFPOSX1
XFILL_1__729_ vdd gnd FILL
XFILL_2__993_ vdd gnd FILL
XFILL_1__1105_ vdd gnd FILL
XFILL_1__1036_ vdd gnd FILL
XFILL_2__1145_ vdd gnd FILL
XFILL_2__1214_ vdd gnd FILL
XFILL_2__1076_ vdd gnd FILL
X_1340_ _1352_/B _1342_/B _817_/A _1341_/B vdd gnd OAI21X1
XFILL_0__816_ vdd gnd FILL
XFILL_0__747_ vdd gnd FILL
X_1271_ _1271_/A _1271_/B _1271_/C _1272_/A vdd gnd OAI21X1
XFILL_3__1185_ vdd gnd FILL
X_1469_ _807_/Y _1503_/CLK _805_/A vdd gnd DFFPOSX1
XFILL_2__976_ vdd gnd FILL
XFILL_1__1019_ vdd gnd FILL
X_982_ _983_/A _982_/B _982_/C _987_/B vdd gnd NAND3X1
XFILL_0__1261_ vdd gnd FILL
XFILL_0__1330_ vdd gnd FILL
XFILL_0__1192_ vdd gnd FILL
XFILL_2__1128_ vdd gnd FILL
XFILL_2__1059_ vdd gnd FILL
X_1323_ _744_/D _1370_/A _1324_/C vdd gnd NAND2X1
XFILL_1__994_ vdd gnd FILL
X_1185_ _1482_/Q _1356_/B vdd gnd INVX1
XFILL_1__1370_ vdd gnd FILL
XFILL_3__1306_ vdd gnd FILL
X_1254_ _1254_/A _1254_/B _812_/A _1255_/D vdd gnd OAI21X1
XFILL_2__761_ vdd gnd FILL
XFILL_0__1528_ vdd gnd FILL
XFILL_2__830_ vdd gnd FILL
XFILL_2__959_ vdd gnd FILL
X_965_ _965_/A _965_/B _967_/B vdd gnd XNOR2X1
X_896_ _904_/B _904_/A _904_/C _921_/C vdd gnd AOI21X1
XFILL_0__1313_ vdd gnd FILL
XFILL_0__1244_ vdd gnd FILL
XFILL_0__1175_ vdd gnd FILL
X_1306_ _1306_/A _1311_/B vdd gnd INVX1
XFILL_1__977_ vdd gnd FILL
X_1237_ _1484_/Q _1376_/B vdd gnd INVX1
XFILL_1__1353_ vdd gnd FILL
XFILL_1__1422_ vdd gnd FILL
X_1099_ _1212_/A _1099_/B _1215_/B vdd gnd NAND2X1
X_1168_ _1168_/A _1168_/B _1168_/C _1173_/C vdd gnd AOI21X1
XFILL_2__813_ vdd gnd FILL
XFILL_2__744_ vdd gnd FILL
XFILL_1__1284_ vdd gnd FILL
XFILL_3_CLKBUF1_insert11 vdd gnd FILL
XFILL_2__1531_ vdd gnd FILL
X_750_ _751_/A _977_/A _751_/C vdd gnd NAND2X1
XFILL_2__1393_ vdd gnd FILL
XFILL_0__995_ vdd gnd FILL
X_948_ _952_/A _952_/B _951_/A _957_/A vdd gnd OAI21X1
XFILL_1__900_ vdd gnd FILL
XFILL_1__831_ vdd gnd FILL
XFILL_1__762_ vdd gnd FILL
X_1022_ _1025_/A _1025_/B _1034_/B vdd gnd NAND2X1
X_879_ _879_/A _879_/B _879_/C _880_/B vdd gnd AOI21X1
XFILL_0__1227_ vdd gnd FILL
XFILL_0__1158_ vdd gnd FILL
XFILL_0__1089_ vdd gnd FILL
XFILL86850x11850 vdd gnd FILL
XFILL86550x46950 vdd gnd FILL
XFILL_1__1405_ vdd gnd FILL
XFILL_1__1336_ vdd gnd FILL
XFILL_1__1267_ vdd gnd FILL
XFILL_2__727_ vdd gnd FILL
XFILL_0__780_ vdd gnd FILL
XFILL_1__1198_ vdd gnd FILL
X_802_ _802_/A _804_/B vdd gnd INVX1
XFILL_2__1376_ vdd gnd FILL
X_733_ _743_/A _733_/B _734_/C vdd gnd NAND2X1
XFILL_2__1445_ vdd gnd FILL
XFILL_0__978_ vdd gnd FILL
XFILL_0__1012_ vdd gnd FILL
XFILL_1__745_ vdd gnd FILL
XFILL_1__814_ vdd gnd FILL
X_1005_ _995_/B _995_/C _996_/A _1010_/A vdd gnd AOI21X1
XFILL_1__1121_ vdd gnd FILL
XFILL_1__1052_ vdd gnd FILL
XFILL86850x23550 vdd gnd FILL
XFILL_2__1230_ vdd gnd FILL
XFILL_1__1319_ vdd gnd FILL
XFILL_2__1161_ vdd gnd FILL
XFILL_2__1092_ vdd gnd FILL
XFILL_0__832_ vdd gnd FILL
XFILL_0__901_ vdd gnd FILL
XFILL_0__763_ vdd gnd FILL
XFILL_2__1359_ vdd gnd FILL
XFILL_2__1428_ vdd gnd FILL
X_1485_ _1485_/D _1503_/CLK _1485_/Q vdd gnd DFFPOSX1
XFILL_2_BUFX2_insert24 vdd gnd FILL
.ends

