magic
tech scmos
magscale 1 30
timestamp 1719958228
<< checkpaint >>
rect 41700 43460 146540 146600
<< metal1 >>
rect 106100 145925 113245 146000
rect 106100 145835 106207 145925
rect 106297 145835 106387 145925
rect 106477 145835 106567 145925
rect 106657 145835 106747 145925
rect 106837 145835 106927 145925
rect 107017 145835 107107 145925
rect 107197 145835 107287 145925
rect 107377 145835 107467 145925
rect 107557 145835 107647 145925
rect 107737 145835 107827 145925
rect 107917 145835 108007 145925
rect 108097 145835 108187 145925
rect 108277 145835 108367 145925
rect 108457 145835 108547 145925
rect 108637 145835 108727 145925
rect 108817 145835 108907 145925
rect 108997 145835 109087 145925
rect 109177 145835 109267 145925
rect 109357 145835 109447 145925
rect 109537 145835 109627 145925
rect 109717 145835 109807 145925
rect 109897 145835 109987 145925
rect 110077 145835 110167 145925
rect 110257 145835 110347 145925
rect 110437 145835 110527 145925
rect 110617 145835 110707 145925
rect 110797 145835 110887 145925
rect 110977 145835 111067 145925
rect 111157 145835 111247 145925
rect 111337 145835 111427 145925
rect 111517 145835 111607 145925
rect 111697 145835 111787 145925
rect 111877 145835 111967 145925
rect 112057 145835 112147 145925
rect 112237 145835 112327 145925
rect 112417 145835 112507 145925
rect 112597 145835 112687 145925
rect 112777 145835 112867 145925
rect 112957 145835 113047 145925
rect 113137 145835 113245 145925
rect 106100 145745 113245 145835
rect 106100 145655 106207 145745
rect 106297 145655 106387 145745
rect 106477 145655 106567 145745
rect 106657 145655 106747 145745
rect 106837 145655 106927 145745
rect 107017 145655 107107 145745
rect 107197 145655 107287 145745
rect 107377 145655 107467 145745
rect 107557 145655 107647 145745
rect 107737 145655 107827 145745
rect 107917 145655 108007 145745
rect 108097 145655 108187 145745
rect 108277 145655 108367 145745
rect 108457 145655 108547 145745
rect 108637 145655 108727 145745
rect 108817 145655 108907 145745
rect 108997 145655 109087 145745
rect 109177 145655 109267 145745
rect 109357 145655 109447 145745
rect 109537 145655 109627 145745
rect 109717 145655 109807 145745
rect 109897 145655 109987 145745
rect 110077 145655 110167 145745
rect 110257 145655 110347 145745
rect 110437 145655 110527 145745
rect 110617 145655 110707 145745
rect 110797 145655 110887 145745
rect 110977 145655 111067 145745
rect 111157 145655 111247 145745
rect 111337 145655 111427 145745
rect 111517 145655 111607 145745
rect 111697 145655 111787 145745
rect 111877 145655 111967 145745
rect 112057 145655 112147 145745
rect 112237 145655 112327 145745
rect 112417 145655 112507 145745
rect 112597 145655 112687 145745
rect 112777 145655 112867 145745
rect 112957 145655 113047 145745
rect 113137 145655 113245 145745
rect 106100 145565 113245 145655
rect 106100 145475 106207 145565
rect 106297 145475 106387 145565
rect 106477 145475 106567 145565
rect 106657 145475 106747 145565
rect 106837 145475 106927 145565
rect 107017 145475 107107 145565
rect 107197 145475 107287 145565
rect 107377 145475 107467 145565
rect 107557 145475 107647 145565
rect 107737 145475 107827 145565
rect 107917 145475 108007 145565
rect 108097 145475 108187 145565
rect 108277 145475 108367 145565
rect 108457 145475 108547 145565
rect 108637 145475 108727 145565
rect 108817 145475 108907 145565
rect 108997 145475 109087 145565
rect 109177 145475 109267 145565
rect 109357 145475 109447 145565
rect 109537 145475 109627 145565
rect 109717 145475 109807 145565
rect 109897 145475 109987 145565
rect 110077 145475 110167 145565
rect 110257 145475 110347 145565
rect 110437 145475 110527 145565
rect 110617 145475 110707 145565
rect 110797 145475 110887 145565
rect 110977 145475 111067 145565
rect 111157 145475 111247 145565
rect 111337 145475 111427 145565
rect 111517 145475 111607 145565
rect 111697 145475 111787 145565
rect 111877 145475 111967 145565
rect 112057 145475 112147 145565
rect 112237 145475 112327 145565
rect 112417 145475 112507 145565
rect 112597 145475 112687 145565
rect 112777 145475 112867 145565
rect 112957 145475 113047 145565
rect 113137 145475 113245 145565
rect 106100 145385 113245 145475
rect 106100 145295 106207 145385
rect 106297 145295 106387 145385
rect 106477 145295 106567 145385
rect 106657 145295 106747 145385
rect 106837 145295 106927 145385
rect 107017 145295 107107 145385
rect 107197 145295 107287 145385
rect 107377 145295 107467 145385
rect 107557 145295 107647 145385
rect 107737 145295 107827 145385
rect 107917 145295 108007 145385
rect 108097 145295 108187 145385
rect 108277 145295 108367 145385
rect 108457 145295 108547 145385
rect 108637 145295 108727 145385
rect 108817 145295 108907 145385
rect 108997 145295 109087 145385
rect 109177 145295 109267 145385
rect 109357 145295 109447 145385
rect 109537 145295 109627 145385
rect 109717 145295 109807 145385
rect 109897 145295 109987 145385
rect 110077 145295 110167 145385
rect 110257 145295 110347 145385
rect 110437 145295 110527 145385
rect 110617 145295 110707 145385
rect 110797 145295 110887 145385
rect 110977 145295 111067 145385
rect 111157 145295 111247 145385
rect 111337 145295 111427 145385
rect 111517 145295 111607 145385
rect 111697 145295 111787 145385
rect 111877 145295 111967 145385
rect 112057 145295 112147 145385
rect 112237 145295 112327 145385
rect 112417 145295 112507 145385
rect 112597 145295 112687 145385
rect 112777 145295 112867 145385
rect 112957 145295 113047 145385
rect 113137 145295 113245 145385
rect 106100 145205 113245 145295
rect 106100 145115 106207 145205
rect 106297 145115 106387 145205
rect 106477 145115 106567 145205
rect 106657 145115 106747 145205
rect 106837 145115 106927 145205
rect 107017 145115 107107 145205
rect 107197 145115 107287 145205
rect 107377 145115 107467 145205
rect 107557 145115 107647 145205
rect 107737 145115 107827 145205
rect 107917 145115 108007 145205
rect 108097 145115 108187 145205
rect 108277 145115 108367 145205
rect 108457 145115 108547 145205
rect 108637 145115 108727 145205
rect 108817 145115 108907 145205
rect 108997 145115 109087 145205
rect 109177 145115 109267 145205
rect 109357 145115 109447 145205
rect 109537 145115 109627 145205
rect 109717 145115 109807 145205
rect 109897 145115 109987 145205
rect 110077 145115 110167 145205
rect 110257 145115 110347 145205
rect 110437 145115 110527 145205
rect 110617 145115 110707 145205
rect 110797 145115 110887 145205
rect 110977 145115 111067 145205
rect 111157 145115 111247 145205
rect 111337 145115 111427 145205
rect 111517 145115 111607 145205
rect 111697 145115 111787 145205
rect 111877 145115 111967 145205
rect 112057 145115 112147 145205
rect 112237 145115 112327 145205
rect 112417 145115 112507 145205
rect 112597 145115 112687 145205
rect 112777 145115 112867 145205
rect 112957 145115 113047 145205
rect 113137 145115 113245 145205
rect 106100 145025 113245 145115
rect 106100 144935 106207 145025
rect 106297 144935 106387 145025
rect 106477 144935 106567 145025
rect 106657 144935 106747 145025
rect 106837 144935 106927 145025
rect 107017 144935 107107 145025
rect 107197 144935 107287 145025
rect 107377 144935 107467 145025
rect 107557 144935 107647 145025
rect 107737 144935 107827 145025
rect 107917 144935 108007 145025
rect 108097 144935 108187 145025
rect 108277 144935 108367 145025
rect 108457 144935 108547 145025
rect 108637 144935 108727 145025
rect 108817 144935 108907 145025
rect 108997 144935 109087 145025
rect 109177 144935 109267 145025
rect 109357 144935 109447 145025
rect 109537 144935 109627 145025
rect 109717 144935 109807 145025
rect 109897 144935 109987 145025
rect 110077 144935 110167 145025
rect 110257 144935 110347 145025
rect 110437 144935 110527 145025
rect 110617 144935 110707 145025
rect 110797 144935 110887 145025
rect 110977 144935 111067 145025
rect 111157 144935 111247 145025
rect 111337 144935 111427 145025
rect 111517 144935 111607 145025
rect 111697 144935 111787 145025
rect 111877 144935 111967 145025
rect 112057 144935 112147 145025
rect 112237 144935 112327 145025
rect 112417 144935 112507 145025
rect 112597 144935 112687 145025
rect 112777 144935 112867 145025
rect 112957 144935 113047 145025
rect 113137 144935 113245 145025
rect 106100 144845 113245 144935
rect 106100 144755 106207 144845
rect 106297 144755 106387 144845
rect 106477 144755 106567 144845
rect 106657 144755 106747 144845
rect 106837 144755 106927 144845
rect 107017 144755 107107 144845
rect 107197 144755 107287 144845
rect 107377 144755 107467 144845
rect 107557 144755 107647 144845
rect 107737 144755 107827 144845
rect 107917 144755 108007 144845
rect 108097 144755 108187 144845
rect 108277 144755 108367 144845
rect 108457 144755 108547 144845
rect 108637 144755 108727 144845
rect 108817 144755 108907 144845
rect 108997 144755 109087 144845
rect 109177 144755 109267 144845
rect 109357 144755 109447 144845
rect 109537 144755 109627 144845
rect 109717 144755 109807 144845
rect 109897 144755 109987 144845
rect 110077 144755 110167 144845
rect 110257 144755 110347 144845
rect 110437 144755 110527 144845
rect 110617 144755 110707 144845
rect 110797 144755 110887 144845
rect 110977 144755 111067 144845
rect 111157 144755 111247 144845
rect 111337 144755 111427 144845
rect 111517 144755 111607 144845
rect 111697 144755 111787 144845
rect 111877 144755 111967 144845
rect 112057 144755 112147 144845
rect 112237 144755 112327 144845
rect 112417 144755 112507 144845
rect 112597 144755 112687 144845
rect 112777 144755 112867 144845
rect 112957 144755 113047 144845
rect 113137 144755 113245 144845
rect 106100 144665 113245 144755
rect 106100 144575 106207 144665
rect 106297 144575 106387 144665
rect 106477 144575 106567 144665
rect 106657 144575 106747 144665
rect 106837 144575 106927 144665
rect 107017 144575 107107 144665
rect 107197 144575 107287 144665
rect 107377 144575 107467 144665
rect 107557 144575 107647 144665
rect 107737 144575 107827 144665
rect 107917 144575 108007 144665
rect 108097 144575 108187 144665
rect 108277 144575 108367 144665
rect 108457 144575 108547 144665
rect 108637 144575 108727 144665
rect 108817 144575 108907 144665
rect 108997 144575 109087 144665
rect 109177 144575 109267 144665
rect 109357 144575 109447 144665
rect 109537 144575 109627 144665
rect 109717 144575 109807 144665
rect 109897 144575 109987 144665
rect 110077 144575 110167 144665
rect 110257 144575 110347 144665
rect 110437 144575 110527 144665
rect 110617 144575 110707 144665
rect 110797 144575 110887 144665
rect 110977 144575 111067 144665
rect 111157 144575 111247 144665
rect 111337 144575 111427 144665
rect 111517 144575 111607 144665
rect 111697 144575 111787 144665
rect 111877 144575 111967 144665
rect 112057 144575 112147 144665
rect 112237 144575 112327 144665
rect 112417 144575 112507 144665
rect 112597 144575 112687 144665
rect 112777 144575 112867 144665
rect 112957 144575 113047 144665
rect 113137 144575 113245 144665
rect 106100 144500 113245 144575
rect 103800 143060 104500 144200
rect 106100 143700 144145 144500
rect 143245 140000 144145 143700
rect 143440 116155 143860 116260
rect 143440 116065 143515 116155
rect 143605 116065 143695 116155
rect 143785 116065 143860 116155
rect 143440 115960 143860 116065
rect 143650 114035 143860 114460
rect 143650 113320 144075 113530
rect 145400 103205 145940 103320
rect 145400 103115 145535 103205
rect 145625 103115 145715 103205
rect 145805 103115 145940 103205
rect 145400 103000 145940 103115
rect 145400 87120 145650 103000
rect 145395 86800 145910 87120
rect 45655 84790 46530 84930
rect 45655 84700 45777 84790
rect 45867 84700 45957 84790
rect 46047 84700 46137 84790
rect 46227 84700 46317 84790
rect 46407 84700 46530 84790
rect 45655 84610 46530 84700
rect 45655 84520 45777 84610
rect 45867 84520 45957 84610
rect 46047 84520 46137 84610
rect 46227 84520 46317 84610
rect 46407 84520 46530 84610
rect 45655 84430 46530 84520
rect 45655 84340 45777 84430
rect 45867 84340 45957 84430
rect 46047 84340 46137 84430
rect 46227 84340 46317 84430
rect 46407 84340 46530 84430
rect 45655 84250 46530 84340
rect 45655 84160 45777 84250
rect 45867 84160 45957 84250
rect 46047 84160 46137 84250
rect 46227 84160 46317 84250
rect 46407 84160 46530 84250
rect 45655 84070 46530 84160
rect 45655 83980 45777 84070
rect 45867 83980 45957 84070
rect 46047 83980 46137 84070
rect 46227 83980 46317 84070
rect 46407 83980 46530 84070
rect 45655 83890 46530 83980
rect 45655 83800 45777 83890
rect 45867 83800 45957 83890
rect 46047 83800 46137 83890
rect 46227 83800 46317 83890
rect 46407 83800 46530 83890
rect 45655 83710 46530 83800
rect 45655 83620 45777 83710
rect 45867 83620 45957 83710
rect 46047 83620 46137 83710
rect 46227 83620 46317 83710
rect 46407 83620 46530 83710
rect 45655 83530 46530 83620
rect 45655 83440 45777 83530
rect 45867 83440 45957 83530
rect 46047 83440 46137 83530
rect 46227 83440 46317 83530
rect 46407 83440 46530 83530
rect 45655 83350 46530 83440
rect 45655 83260 45777 83350
rect 45867 83260 45957 83350
rect 46047 83260 46137 83350
rect 46227 83260 46317 83350
rect 46407 83260 46530 83350
rect 45655 83170 46530 83260
rect 45655 83080 45777 83170
rect 45867 83080 45957 83170
rect 46047 83080 46137 83170
rect 46227 83080 46317 83170
rect 46407 83080 46530 83170
rect 45655 82990 46530 83080
rect 45655 82900 45777 82990
rect 45867 82900 45957 82990
rect 46047 82900 46137 82990
rect 46227 82900 46317 82990
rect 46407 82900 46530 82990
rect 45655 82810 46530 82900
rect 45655 82720 45777 82810
rect 45867 82720 45957 82810
rect 46047 82720 46137 82810
rect 46227 82720 46317 82810
rect 46407 82720 46530 82810
rect 45655 82630 46530 82720
rect 45655 82540 45777 82630
rect 45867 82540 45957 82630
rect 46047 82540 46137 82630
rect 46227 82540 46317 82630
rect 46407 82540 46530 82630
rect 45655 82450 46530 82540
rect 45655 82360 45777 82450
rect 45867 82360 45957 82450
rect 46047 82360 46137 82450
rect 46227 82360 46317 82450
rect 46407 82360 46530 82450
rect 45655 82270 46530 82360
rect 45655 82180 45777 82270
rect 45867 82180 45957 82270
rect 46047 82180 46137 82270
rect 46227 82180 46317 82270
rect 46407 82180 46530 82270
rect 45655 82090 46530 82180
rect 45655 82000 45777 82090
rect 45867 82000 45957 82090
rect 46047 82000 46137 82090
rect 46227 82000 46317 82090
rect 46407 82000 46530 82090
rect 45655 81910 46530 82000
rect 45655 81820 45777 81910
rect 45867 81820 45957 81910
rect 46047 81820 46137 81910
rect 46227 81820 46317 81910
rect 46407 81820 46530 81910
rect 45655 81730 46530 81820
rect 45655 81640 45777 81730
rect 45867 81640 45957 81730
rect 46047 81640 46137 81730
rect 46227 81640 46317 81730
rect 46407 81640 46530 81730
rect 45655 81550 46530 81640
rect 45655 81460 45777 81550
rect 45867 81460 45957 81550
rect 46047 81460 46137 81550
rect 46227 81460 46317 81550
rect 46407 81460 46530 81550
rect 45655 81370 46530 81460
rect 45655 81280 45777 81370
rect 45867 81280 45957 81370
rect 46047 81280 46137 81370
rect 46227 81280 46317 81370
rect 46407 81280 46530 81370
rect 45655 81190 46530 81280
rect 45655 81100 45777 81190
rect 45867 81100 45957 81190
rect 46047 81100 46137 81190
rect 46227 81100 46317 81190
rect 46407 81100 46530 81190
rect 45655 81010 46530 81100
rect 45655 80920 45777 81010
rect 45867 80920 45957 81010
rect 46047 80920 46137 81010
rect 46227 80920 46317 81010
rect 46407 80920 46530 81010
rect 45655 80830 46530 80920
rect 45655 80740 45777 80830
rect 45867 80740 45957 80830
rect 46047 80740 46137 80830
rect 46227 80740 46317 80830
rect 46407 80740 46530 80830
rect 45655 80650 46530 80740
rect 45655 80560 45777 80650
rect 45867 80560 45957 80650
rect 46047 80560 46137 80650
rect 46227 80560 46317 80650
rect 46407 80560 46530 80650
rect 45655 80470 46530 80560
rect 45655 80380 45777 80470
rect 45867 80380 45957 80470
rect 46047 80380 46137 80470
rect 46227 80380 46317 80470
rect 46407 80380 46530 80470
rect 45655 80290 46530 80380
rect 45655 80200 45777 80290
rect 45867 80200 45957 80290
rect 46047 80200 46137 80290
rect 46227 80200 46317 80290
rect 46407 80200 46530 80290
rect 45655 80110 46530 80200
rect 45655 80020 45777 80110
rect 45867 80020 45957 80110
rect 46047 80020 46137 80110
rect 46227 80020 46317 80110
rect 46407 80020 46530 80110
rect 45655 79930 46530 80020
rect 45655 79840 45777 79930
rect 45867 79840 45957 79930
rect 46047 79840 46137 79930
rect 46227 79840 46317 79930
rect 46407 79840 46530 79930
rect 45655 79750 46530 79840
rect 45655 79660 45777 79750
rect 45867 79660 45957 79750
rect 46047 79660 46137 79750
rect 46227 79660 46317 79750
rect 46407 79660 46530 79750
rect 45655 79570 46530 79660
rect 45655 79480 45777 79570
rect 45867 79480 45957 79570
rect 46047 79480 46137 79570
rect 46227 79480 46317 79570
rect 46407 79480 46530 79570
rect 45655 79390 46530 79480
rect 45655 79300 45777 79390
rect 45867 79300 45957 79390
rect 46047 79300 46137 79390
rect 46227 79300 46317 79390
rect 46407 79300 46530 79390
rect 45655 79210 46530 79300
rect 45655 79120 45777 79210
rect 45867 79120 45957 79210
rect 46047 79120 46137 79210
rect 46227 79120 46317 79210
rect 46407 79120 46530 79210
rect 45655 79030 46530 79120
rect 45655 78940 45777 79030
rect 45867 78940 45957 79030
rect 46047 78940 46137 79030
rect 46227 78940 46317 79030
rect 46407 78940 46530 79030
rect 45655 78850 46530 78940
rect 45655 78760 45777 78850
rect 45867 78760 45957 78850
rect 46047 78760 46137 78850
rect 46227 78760 46317 78850
rect 46407 78760 46530 78850
rect 45655 78670 46530 78760
rect 45655 78580 45777 78670
rect 45867 78580 45957 78670
rect 46047 78580 46137 78670
rect 46227 78580 46317 78670
rect 46407 78580 46530 78670
rect 45655 78490 46530 78580
rect 45655 78400 45777 78490
rect 45867 78400 45957 78490
rect 46047 78400 46137 78490
rect 46227 78400 46317 78490
rect 46407 78400 46530 78490
rect 45655 78310 46530 78400
rect 45655 78220 45777 78310
rect 45867 78220 45957 78310
rect 46047 78220 46137 78310
rect 46227 78220 46317 78310
rect 46407 78220 46530 78310
rect 45655 78080 46530 78220
rect 45955 75940 46235 76360
rect 143690 59375 143900 59815
rect 143740 57040 144260 57255
rect 145400 56675 145650 86800
rect 143740 56440 144260 56655
rect 145400 56585 145480 56675
rect 145570 56585 145650 56675
rect 145400 56440 145650 56585
rect 98400 46402 100050 46475
rect 98400 46312 99690 46402
rect 99780 46312 99870 46402
rect 99960 46312 100050 46402
rect 98400 46240 100050 46312
rect 98400 45900 98700 46240
rect 59800 45807 98700 45900
rect 59800 45717 59915 45807
rect 60005 45717 98700 45807
rect 59800 45627 98700 45717
rect 59800 45537 59915 45627
rect 60005 45600 98700 45627
rect 99000 45795 106945 45900
rect 99000 45705 106615 45795
rect 106705 45705 106795 45795
rect 106885 45705 106945 45795
rect 99000 45600 106945 45705
rect 60005 45537 60120 45600
rect 59800 45445 60120 45537
rect 99000 45300 99300 45600
rect 73300 45195 99300 45300
rect 73300 45105 73415 45195
rect 73505 45105 99300 45195
rect 73300 45000 99300 45105
rect 73300 44135 73620 45000
<< m2contact >>
rect 106207 145835 106297 145925
rect 106387 145835 106477 145925
rect 106567 145835 106657 145925
rect 106747 145835 106837 145925
rect 106927 145835 107017 145925
rect 107107 145835 107197 145925
rect 107287 145835 107377 145925
rect 107467 145835 107557 145925
rect 107647 145835 107737 145925
rect 107827 145835 107917 145925
rect 108007 145835 108097 145925
rect 108187 145835 108277 145925
rect 108367 145835 108457 145925
rect 108547 145835 108637 145925
rect 108727 145835 108817 145925
rect 108907 145835 108997 145925
rect 109087 145835 109177 145925
rect 109267 145835 109357 145925
rect 109447 145835 109537 145925
rect 109627 145835 109717 145925
rect 109807 145835 109897 145925
rect 109987 145835 110077 145925
rect 110167 145835 110257 145925
rect 110347 145835 110437 145925
rect 110527 145835 110617 145925
rect 110707 145835 110797 145925
rect 110887 145835 110977 145925
rect 111067 145835 111157 145925
rect 111247 145835 111337 145925
rect 111427 145835 111517 145925
rect 111607 145835 111697 145925
rect 111787 145835 111877 145925
rect 111967 145835 112057 145925
rect 112147 145835 112237 145925
rect 112327 145835 112417 145925
rect 112507 145835 112597 145925
rect 112687 145835 112777 145925
rect 112867 145835 112957 145925
rect 113047 145835 113137 145925
rect 106207 145655 106297 145745
rect 106387 145655 106477 145745
rect 106567 145655 106657 145745
rect 106747 145655 106837 145745
rect 106927 145655 107017 145745
rect 107107 145655 107197 145745
rect 107287 145655 107377 145745
rect 107467 145655 107557 145745
rect 107647 145655 107737 145745
rect 107827 145655 107917 145745
rect 108007 145655 108097 145745
rect 108187 145655 108277 145745
rect 108367 145655 108457 145745
rect 108547 145655 108637 145745
rect 108727 145655 108817 145745
rect 108907 145655 108997 145745
rect 109087 145655 109177 145745
rect 109267 145655 109357 145745
rect 109447 145655 109537 145745
rect 109627 145655 109717 145745
rect 109807 145655 109897 145745
rect 109987 145655 110077 145745
rect 110167 145655 110257 145745
rect 110347 145655 110437 145745
rect 110527 145655 110617 145745
rect 110707 145655 110797 145745
rect 110887 145655 110977 145745
rect 111067 145655 111157 145745
rect 111247 145655 111337 145745
rect 111427 145655 111517 145745
rect 111607 145655 111697 145745
rect 111787 145655 111877 145745
rect 111967 145655 112057 145745
rect 112147 145655 112237 145745
rect 112327 145655 112417 145745
rect 112507 145655 112597 145745
rect 112687 145655 112777 145745
rect 112867 145655 112957 145745
rect 113047 145655 113137 145745
rect 106207 145475 106297 145565
rect 106387 145475 106477 145565
rect 106567 145475 106657 145565
rect 106747 145475 106837 145565
rect 106927 145475 107017 145565
rect 107107 145475 107197 145565
rect 107287 145475 107377 145565
rect 107467 145475 107557 145565
rect 107647 145475 107737 145565
rect 107827 145475 107917 145565
rect 108007 145475 108097 145565
rect 108187 145475 108277 145565
rect 108367 145475 108457 145565
rect 108547 145475 108637 145565
rect 108727 145475 108817 145565
rect 108907 145475 108997 145565
rect 109087 145475 109177 145565
rect 109267 145475 109357 145565
rect 109447 145475 109537 145565
rect 109627 145475 109717 145565
rect 109807 145475 109897 145565
rect 109987 145475 110077 145565
rect 110167 145475 110257 145565
rect 110347 145475 110437 145565
rect 110527 145475 110617 145565
rect 110707 145475 110797 145565
rect 110887 145475 110977 145565
rect 111067 145475 111157 145565
rect 111247 145475 111337 145565
rect 111427 145475 111517 145565
rect 111607 145475 111697 145565
rect 111787 145475 111877 145565
rect 111967 145475 112057 145565
rect 112147 145475 112237 145565
rect 112327 145475 112417 145565
rect 112507 145475 112597 145565
rect 112687 145475 112777 145565
rect 112867 145475 112957 145565
rect 113047 145475 113137 145565
rect 106207 145295 106297 145385
rect 106387 145295 106477 145385
rect 106567 145295 106657 145385
rect 106747 145295 106837 145385
rect 106927 145295 107017 145385
rect 107107 145295 107197 145385
rect 107287 145295 107377 145385
rect 107467 145295 107557 145385
rect 107647 145295 107737 145385
rect 107827 145295 107917 145385
rect 108007 145295 108097 145385
rect 108187 145295 108277 145385
rect 108367 145295 108457 145385
rect 108547 145295 108637 145385
rect 108727 145295 108817 145385
rect 108907 145295 108997 145385
rect 109087 145295 109177 145385
rect 109267 145295 109357 145385
rect 109447 145295 109537 145385
rect 109627 145295 109717 145385
rect 109807 145295 109897 145385
rect 109987 145295 110077 145385
rect 110167 145295 110257 145385
rect 110347 145295 110437 145385
rect 110527 145295 110617 145385
rect 110707 145295 110797 145385
rect 110887 145295 110977 145385
rect 111067 145295 111157 145385
rect 111247 145295 111337 145385
rect 111427 145295 111517 145385
rect 111607 145295 111697 145385
rect 111787 145295 111877 145385
rect 111967 145295 112057 145385
rect 112147 145295 112237 145385
rect 112327 145295 112417 145385
rect 112507 145295 112597 145385
rect 112687 145295 112777 145385
rect 112867 145295 112957 145385
rect 113047 145295 113137 145385
rect 106207 145115 106297 145205
rect 106387 145115 106477 145205
rect 106567 145115 106657 145205
rect 106747 145115 106837 145205
rect 106927 145115 107017 145205
rect 107107 145115 107197 145205
rect 107287 145115 107377 145205
rect 107467 145115 107557 145205
rect 107647 145115 107737 145205
rect 107827 145115 107917 145205
rect 108007 145115 108097 145205
rect 108187 145115 108277 145205
rect 108367 145115 108457 145205
rect 108547 145115 108637 145205
rect 108727 145115 108817 145205
rect 108907 145115 108997 145205
rect 109087 145115 109177 145205
rect 109267 145115 109357 145205
rect 109447 145115 109537 145205
rect 109627 145115 109717 145205
rect 109807 145115 109897 145205
rect 109987 145115 110077 145205
rect 110167 145115 110257 145205
rect 110347 145115 110437 145205
rect 110527 145115 110617 145205
rect 110707 145115 110797 145205
rect 110887 145115 110977 145205
rect 111067 145115 111157 145205
rect 111247 145115 111337 145205
rect 111427 145115 111517 145205
rect 111607 145115 111697 145205
rect 111787 145115 111877 145205
rect 111967 145115 112057 145205
rect 112147 145115 112237 145205
rect 112327 145115 112417 145205
rect 112507 145115 112597 145205
rect 112687 145115 112777 145205
rect 112867 145115 112957 145205
rect 113047 145115 113137 145205
rect 106207 144935 106297 145025
rect 106387 144935 106477 145025
rect 106567 144935 106657 145025
rect 106747 144935 106837 145025
rect 106927 144935 107017 145025
rect 107107 144935 107197 145025
rect 107287 144935 107377 145025
rect 107467 144935 107557 145025
rect 107647 144935 107737 145025
rect 107827 144935 107917 145025
rect 108007 144935 108097 145025
rect 108187 144935 108277 145025
rect 108367 144935 108457 145025
rect 108547 144935 108637 145025
rect 108727 144935 108817 145025
rect 108907 144935 108997 145025
rect 109087 144935 109177 145025
rect 109267 144935 109357 145025
rect 109447 144935 109537 145025
rect 109627 144935 109717 145025
rect 109807 144935 109897 145025
rect 109987 144935 110077 145025
rect 110167 144935 110257 145025
rect 110347 144935 110437 145025
rect 110527 144935 110617 145025
rect 110707 144935 110797 145025
rect 110887 144935 110977 145025
rect 111067 144935 111157 145025
rect 111247 144935 111337 145025
rect 111427 144935 111517 145025
rect 111607 144935 111697 145025
rect 111787 144935 111877 145025
rect 111967 144935 112057 145025
rect 112147 144935 112237 145025
rect 112327 144935 112417 145025
rect 112507 144935 112597 145025
rect 112687 144935 112777 145025
rect 112867 144935 112957 145025
rect 113047 144935 113137 145025
rect 106207 144755 106297 144845
rect 106387 144755 106477 144845
rect 106567 144755 106657 144845
rect 106747 144755 106837 144845
rect 106927 144755 107017 144845
rect 107107 144755 107197 144845
rect 107287 144755 107377 144845
rect 107467 144755 107557 144845
rect 107647 144755 107737 144845
rect 107827 144755 107917 144845
rect 108007 144755 108097 144845
rect 108187 144755 108277 144845
rect 108367 144755 108457 144845
rect 108547 144755 108637 144845
rect 108727 144755 108817 144845
rect 108907 144755 108997 144845
rect 109087 144755 109177 144845
rect 109267 144755 109357 144845
rect 109447 144755 109537 144845
rect 109627 144755 109717 144845
rect 109807 144755 109897 144845
rect 109987 144755 110077 144845
rect 110167 144755 110257 144845
rect 110347 144755 110437 144845
rect 110527 144755 110617 144845
rect 110707 144755 110797 144845
rect 110887 144755 110977 144845
rect 111067 144755 111157 144845
rect 111247 144755 111337 144845
rect 111427 144755 111517 144845
rect 111607 144755 111697 144845
rect 111787 144755 111877 144845
rect 111967 144755 112057 144845
rect 112147 144755 112237 144845
rect 112327 144755 112417 144845
rect 112507 144755 112597 144845
rect 112687 144755 112777 144845
rect 112867 144755 112957 144845
rect 113047 144755 113137 144845
rect 106207 144575 106297 144665
rect 106387 144575 106477 144665
rect 106567 144575 106657 144665
rect 106747 144575 106837 144665
rect 106927 144575 107017 144665
rect 107107 144575 107197 144665
rect 107287 144575 107377 144665
rect 107467 144575 107557 144665
rect 107647 144575 107737 144665
rect 107827 144575 107917 144665
rect 108007 144575 108097 144665
rect 108187 144575 108277 144665
rect 108367 144575 108457 144665
rect 108547 144575 108637 144665
rect 108727 144575 108817 144665
rect 108907 144575 108997 144665
rect 109087 144575 109177 144665
rect 109267 144575 109357 144665
rect 109447 144575 109537 144665
rect 109627 144575 109717 144665
rect 109807 144575 109897 144665
rect 109987 144575 110077 144665
rect 110167 144575 110257 144665
rect 110347 144575 110437 144665
rect 110527 144575 110617 144665
rect 110707 144575 110797 144665
rect 110887 144575 110977 144665
rect 111067 144575 111157 144665
rect 111247 144575 111337 144665
rect 111427 144575 111517 144665
rect 111607 144575 111697 144665
rect 111787 144575 111877 144665
rect 111967 144575 112057 144665
rect 112147 144575 112237 144665
rect 112327 144575 112417 144665
rect 112507 144575 112597 144665
rect 112687 144575 112777 144665
rect 112867 144575 112957 144665
rect 113047 144575 113137 144665
rect 143515 116065 143605 116155
rect 143695 116065 143785 116155
rect 145535 103115 145625 103205
rect 145715 103115 145805 103205
rect 45777 84700 45867 84790
rect 45957 84700 46047 84790
rect 46137 84700 46227 84790
rect 46317 84700 46407 84790
rect 45777 84520 45867 84610
rect 45957 84520 46047 84610
rect 46137 84520 46227 84610
rect 46317 84520 46407 84610
rect 45777 84340 45867 84430
rect 45957 84340 46047 84430
rect 46137 84340 46227 84430
rect 46317 84340 46407 84430
rect 45777 84160 45867 84250
rect 45957 84160 46047 84250
rect 46137 84160 46227 84250
rect 46317 84160 46407 84250
rect 45777 83980 45867 84070
rect 45957 83980 46047 84070
rect 46137 83980 46227 84070
rect 46317 83980 46407 84070
rect 45777 83800 45867 83890
rect 45957 83800 46047 83890
rect 46137 83800 46227 83890
rect 46317 83800 46407 83890
rect 45777 83620 45867 83710
rect 45957 83620 46047 83710
rect 46137 83620 46227 83710
rect 46317 83620 46407 83710
rect 45777 83440 45867 83530
rect 45957 83440 46047 83530
rect 46137 83440 46227 83530
rect 46317 83440 46407 83530
rect 45777 83260 45867 83350
rect 45957 83260 46047 83350
rect 46137 83260 46227 83350
rect 46317 83260 46407 83350
rect 45777 83080 45867 83170
rect 45957 83080 46047 83170
rect 46137 83080 46227 83170
rect 46317 83080 46407 83170
rect 45777 82900 45867 82990
rect 45957 82900 46047 82990
rect 46137 82900 46227 82990
rect 46317 82900 46407 82990
rect 45777 82720 45867 82810
rect 45957 82720 46047 82810
rect 46137 82720 46227 82810
rect 46317 82720 46407 82810
rect 45777 82540 45867 82630
rect 45957 82540 46047 82630
rect 46137 82540 46227 82630
rect 46317 82540 46407 82630
rect 45777 82360 45867 82450
rect 45957 82360 46047 82450
rect 46137 82360 46227 82450
rect 46317 82360 46407 82450
rect 45777 82180 45867 82270
rect 45957 82180 46047 82270
rect 46137 82180 46227 82270
rect 46317 82180 46407 82270
rect 45777 82000 45867 82090
rect 45957 82000 46047 82090
rect 46137 82000 46227 82090
rect 46317 82000 46407 82090
rect 45777 81820 45867 81910
rect 45957 81820 46047 81910
rect 46137 81820 46227 81910
rect 46317 81820 46407 81910
rect 45777 81640 45867 81730
rect 45957 81640 46047 81730
rect 46137 81640 46227 81730
rect 46317 81640 46407 81730
rect 45777 81460 45867 81550
rect 45957 81460 46047 81550
rect 46137 81460 46227 81550
rect 46317 81460 46407 81550
rect 45777 81280 45867 81370
rect 45957 81280 46047 81370
rect 46137 81280 46227 81370
rect 46317 81280 46407 81370
rect 45777 81100 45867 81190
rect 45957 81100 46047 81190
rect 46137 81100 46227 81190
rect 46317 81100 46407 81190
rect 45777 80920 45867 81010
rect 45957 80920 46047 81010
rect 46137 80920 46227 81010
rect 46317 80920 46407 81010
rect 45777 80740 45867 80830
rect 45957 80740 46047 80830
rect 46137 80740 46227 80830
rect 46317 80740 46407 80830
rect 45777 80560 45867 80650
rect 45957 80560 46047 80650
rect 46137 80560 46227 80650
rect 46317 80560 46407 80650
rect 45777 80380 45867 80470
rect 45957 80380 46047 80470
rect 46137 80380 46227 80470
rect 46317 80380 46407 80470
rect 45777 80200 45867 80290
rect 45957 80200 46047 80290
rect 46137 80200 46227 80290
rect 46317 80200 46407 80290
rect 45777 80020 45867 80110
rect 45957 80020 46047 80110
rect 46137 80020 46227 80110
rect 46317 80020 46407 80110
rect 45777 79840 45867 79930
rect 45957 79840 46047 79930
rect 46137 79840 46227 79930
rect 46317 79840 46407 79930
rect 45777 79660 45867 79750
rect 45957 79660 46047 79750
rect 46137 79660 46227 79750
rect 46317 79660 46407 79750
rect 45777 79480 45867 79570
rect 45957 79480 46047 79570
rect 46137 79480 46227 79570
rect 46317 79480 46407 79570
rect 45777 79300 45867 79390
rect 45957 79300 46047 79390
rect 46137 79300 46227 79390
rect 46317 79300 46407 79390
rect 45777 79120 45867 79210
rect 45957 79120 46047 79210
rect 46137 79120 46227 79210
rect 46317 79120 46407 79210
rect 45777 78940 45867 79030
rect 45957 78940 46047 79030
rect 46137 78940 46227 79030
rect 46317 78940 46407 79030
rect 45777 78760 45867 78850
rect 45957 78760 46047 78850
rect 46137 78760 46227 78850
rect 46317 78760 46407 78850
rect 45777 78580 45867 78670
rect 45957 78580 46047 78670
rect 46137 78580 46227 78670
rect 46317 78580 46407 78670
rect 45777 78400 45867 78490
rect 45957 78400 46047 78490
rect 46137 78400 46227 78490
rect 46317 78400 46407 78490
rect 45777 78220 45867 78310
rect 45957 78220 46047 78310
rect 46137 78220 46227 78310
rect 46317 78220 46407 78310
rect 145480 56585 145570 56675
rect 99690 46312 99780 46402
rect 99870 46312 99960 46402
rect 59915 45717 60005 45807
rect 59915 45537 60005 45627
rect 106615 45705 106705 45795
rect 106795 45705 106885 45795
rect 73415 45105 73505 45195
<< metal2 >>
rect 49000 145510 49320 145940
rect 49000 145420 50845 145510
rect 49000 145330 49067 145420
rect 49157 145330 49247 145420
rect 49337 145330 49427 145420
rect 49517 145330 49607 145420
rect 49697 145330 49787 145420
rect 49877 145330 49967 145420
rect 50057 145330 50147 145420
rect 50237 145330 50327 145420
rect 50417 145330 50507 145420
rect 50597 145330 50687 145420
rect 50777 145330 50845 145420
rect 49000 145240 50845 145330
rect 49000 145150 49067 145240
rect 49157 145150 49247 145240
rect 49337 145150 49427 145240
rect 49517 145150 49607 145240
rect 49697 145150 49787 145240
rect 49877 145150 49967 145240
rect 50057 145150 50147 145240
rect 50237 145150 50327 145240
rect 50417 145150 50507 145240
rect 50597 145150 50687 145240
rect 50777 145150 50845 145240
rect 49000 145060 50845 145150
rect 49000 144970 49067 145060
rect 49157 144970 49247 145060
rect 49337 144970 49427 145060
rect 49517 144970 49607 145060
rect 49697 144970 49787 145060
rect 49877 144970 49967 145060
rect 50057 144970 50147 145060
rect 50237 144970 50327 145060
rect 50417 144970 50507 145060
rect 50597 144970 50687 145060
rect 50777 144970 50845 145060
rect 49000 144880 50845 144970
rect 49000 144790 49067 144880
rect 49157 144790 49247 144880
rect 49337 144790 49427 144880
rect 49517 144790 49607 144880
rect 49697 144790 49787 144880
rect 49877 144790 49967 144880
rect 50057 144790 50147 144880
rect 50237 144790 50327 144880
rect 50417 144790 50507 144880
rect 50597 144790 50687 144880
rect 50777 144790 50845 144880
rect 49000 144700 50845 144790
rect 62500 144205 62820 145940
rect 62500 144117 64455 144205
rect 62500 144027 62622 144117
rect 62712 144027 62802 144117
rect 62892 144027 62982 144117
rect 63072 144027 63162 144117
rect 63252 144027 63342 144117
rect 63432 144027 63522 144117
rect 63612 144027 63702 144117
rect 63792 144027 63882 144117
rect 63972 144027 64062 144117
rect 64152 144027 64242 144117
rect 64332 144027 64455 144117
rect 62500 143937 64455 144027
rect 62500 143847 62622 143937
rect 62712 143847 62802 143937
rect 62892 143847 62982 143937
rect 63072 143847 63162 143937
rect 63252 143847 63342 143937
rect 63432 143847 63522 143937
rect 63612 143847 63702 143937
rect 63792 143847 63882 143937
rect 63972 143847 64062 143937
rect 64152 143847 64242 143937
rect 64332 143847 64455 143937
rect 62500 143757 64455 143847
rect 62500 143667 62622 143757
rect 62712 143667 62802 143757
rect 62892 143667 62982 143757
rect 63072 143667 63162 143757
rect 63252 143667 63342 143757
rect 63432 143667 63522 143757
rect 63612 143667 63702 143757
rect 63792 143667 63882 143757
rect 63972 143667 64062 143757
rect 64152 143667 64242 143757
rect 64332 143667 64455 143757
rect 62500 143577 64455 143667
rect 62500 143487 62622 143577
rect 62712 143487 62802 143577
rect 62892 143487 62982 143577
rect 63072 143487 63162 143577
rect 63252 143487 63342 143577
rect 63432 143487 63522 143577
rect 63612 143487 63702 143577
rect 63792 143487 63882 143577
rect 63972 143487 64062 143577
rect 64152 143487 64242 143577
rect 64332 143487 64455 143577
rect 62500 143400 64455 143487
rect 76000 142900 76320 145940
rect 76000 142100 79780 142900
rect 77850 141260 78750 141350
rect 77850 141170 77985 141260
rect 78075 141170 78165 141260
rect 78255 141170 78345 141260
rect 78435 141170 78525 141260
rect 78615 141170 78750 141260
rect 77850 141080 78750 141170
rect 77850 140990 77985 141080
rect 78075 140990 78165 141080
rect 78255 140990 78345 141080
rect 78435 140990 78525 141080
rect 78615 140990 78750 141080
rect 77850 140900 78750 140990
rect 79235 140900 79780 142100
rect 89500 141350 89820 145940
rect 106100 145925 113245 146000
rect 106100 145835 106207 145925
rect 106297 145835 106387 145925
rect 106477 145835 106567 145925
rect 106657 145835 106747 145925
rect 106837 145835 106927 145925
rect 107017 145835 107107 145925
rect 107197 145835 107287 145925
rect 107377 145835 107467 145925
rect 107557 145835 107647 145925
rect 107737 145835 107827 145925
rect 107917 145835 108007 145925
rect 108097 145835 108187 145925
rect 108277 145835 108367 145925
rect 108457 145835 108547 145925
rect 108637 145835 108727 145925
rect 108817 145835 108907 145925
rect 108997 145835 109087 145925
rect 109177 145835 109267 145925
rect 109357 145835 109447 145925
rect 109537 145835 109627 145925
rect 109717 145835 109807 145925
rect 109897 145835 109987 145925
rect 110077 145835 110167 145925
rect 110257 145835 110347 145925
rect 110437 145835 110527 145925
rect 110617 145835 110707 145925
rect 110797 145835 110887 145925
rect 110977 145835 111067 145925
rect 111157 145835 111247 145925
rect 111337 145835 111427 145925
rect 111517 145835 111607 145925
rect 111697 145835 111787 145925
rect 111877 145835 111967 145925
rect 112057 145835 112147 145925
rect 112237 145835 112327 145925
rect 112417 145835 112507 145925
rect 112597 145835 112687 145925
rect 112777 145835 112867 145925
rect 112957 145835 113047 145925
rect 113137 145835 113245 145925
rect 106100 145745 113245 145835
rect 106100 145655 106207 145745
rect 106297 145655 106387 145745
rect 106477 145655 106567 145745
rect 106657 145655 106747 145745
rect 106837 145655 106927 145745
rect 107017 145655 107107 145745
rect 107197 145655 107287 145745
rect 107377 145655 107467 145745
rect 107557 145655 107647 145745
rect 107737 145655 107827 145745
rect 107917 145655 108007 145745
rect 108097 145655 108187 145745
rect 108277 145655 108367 145745
rect 108457 145655 108547 145745
rect 108637 145655 108727 145745
rect 108817 145655 108907 145745
rect 108997 145655 109087 145745
rect 109177 145655 109267 145745
rect 109357 145655 109447 145745
rect 109537 145655 109627 145745
rect 109717 145655 109807 145745
rect 109897 145655 109987 145745
rect 110077 145655 110167 145745
rect 110257 145655 110347 145745
rect 110437 145655 110527 145745
rect 110617 145655 110707 145745
rect 110797 145655 110887 145745
rect 110977 145655 111067 145745
rect 111157 145655 111247 145745
rect 111337 145655 111427 145745
rect 111517 145655 111607 145745
rect 111697 145655 111787 145745
rect 111877 145655 111967 145745
rect 112057 145655 112147 145745
rect 112237 145655 112327 145745
rect 112417 145655 112507 145745
rect 112597 145655 112687 145745
rect 112777 145655 112867 145745
rect 112957 145655 113047 145745
rect 113137 145655 113245 145745
rect 106100 145565 113245 145655
rect 106100 145475 106207 145565
rect 106297 145475 106387 145565
rect 106477 145475 106567 145565
rect 106657 145475 106747 145565
rect 106837 145475 106927 145565
rect 107017 145475 107107 145565
rect 107197 145475 107287 145565
rect 107377 145475 107467 145565
rect 107557 145475 107647 145565
rect 107737 145475 107827 145565
rect 107917 145475 108007 145565
rect 108097 145475 108187 145565
rect 108277 145475 108367 145565
rect 108457 145475 108547 145565
rect 108637 145475 108727 145565
rect 108817 145475 108907 145565
rect 108997 145475 109087 145565
rect 109177 145475 109267 145565
rect 109357 145475 109447 145565
rect 109537 145475 109627 145565
rect 109717 145475 109807 145565
rect 109897 145475 109987 145565
rect 110077 145475 110167 145565
rect 110257 145475 110347 145565
rect 110437 145475 110527 145565
rect 110617 145475 110707 145565
rect 110797 145475 110887 145565
rect 110977 145475 111067 145565
rect 111157 145475 111247 145565
rect 111337 145475 111427 145565
rect 111517 145475 111607 145565
rect 111697 145475 111787 145565
rect 111877 145475 111967 145565
rect 112057 145475 112147 145565
rect 112237 145475 112327 145565
rect 112417 145475 112507 145565
rect 112597 145475 112687 145565
rect 112777 145475 112867 145565
rect 112957 145475 113047 145565
rect 113137 145475 113245 145565
rect 106100 145385 113245 145475
rect 106100 145295 106207 145385
rect 106297 145295 106387 145385
rect 106477 145295 106567 145385
rect 106657 145295 106747 145385
rect 106837 145295 106927 145385
rect 107017 145295 107107 145385
rect 107197 145295 107287 145385
rect 107377 145295 107467 145385
rect 107557 145295 107647 145385
rect 107737 145295 107827 145385
rect 107917 145295 108007 145385
rect 108097 145295 108187 145385
rect 108277 145295 108367 145385
rect 108457 145295 108547 145385
rect 108637 145295 108727 145385
rect 108817 145295 108907 145385
rect 108997 145295 109087 145385
rect 109177 145295 109267 145385
rect 109357 145295 109447 145385
rect 109537 145295 109627 145385
rect 109717 145295 109807 145385
rect 109897 145295 109987 145385
rect 110077 145295 110167 145385
rect 110257 145295 110347 145385
rect 110437 145295 110527 145385
rect 110617 145295 110707 145385
rect 110797 145295 110887 145385
rect 110977 145295 111067 145385
rect 111157 145295 111247 145385
rect 111337 145295 111427 145385
rect 111517 145295 111607 145385
rect 111697 145295 111787 145385
rect 111877 145295 111967 145385
rect 112057 145295 112147 145385
rect 112237 145295 112327 145385
rect 112417 145295 112507 145385
rect 112597 145295 112687 145385
rect 112777 145295 112867 145385
rect 112957 145295 113047 145385
rect 113137 145295 113245 145385
rect 106100 145205 113245 145295
rect 106100 145115 106207 145205
rect 106297 145115 106387 145205
rect 106477 145115 106567 145205
rect 106657 145115 106747 145205
rect 106837 145115 106927 145205
rect 107017 145115 107107 145205
rect 107197 145115 107287 145205
rect 107377 145115 107467 145205
rect 107557 145115 107647 145205
rect 107737 145115 107827 145205
rect 107917 145115 108007 145205
rect 108097 145115 108187 145205
rect 108277 145115 108367 145205
rect 108457 145115 108547 145205
rect 108637 145115 108727 145205
rect 108817 145115 108907 145205
rect 108997 145115 109087 145205
rect 109177 145115 109267 145205
rect 109357 145115 109447 145205
rect 109537 145115 109627 145205
rect 109717 145115 109807 145205
rect 109897 145115 109987 145205
rect 110077 145115 110167 145205
rect 110257 145115 110347 145205
rect 110437 145115 110527 145205
rect 110617 145115 110707 145205
rect 110797 145115 110887 145205
rect 110977 145115 111067 145205
rect 111157 145115 111247 145205
rect 111337 145115 111427 145205
rect 111517 145115 111607 145205
rect 111697 145115 111787 145205
rect 111877 145115 111967 145205
rect 112057 145115 112147 145205
rect 112237 145115 112327 145205
rect 112417 145115 112507 145205
rect 112597 145115 112687 145205
rect 112777 145115 112867 145205
rect 112957 145115 113047 145205
rect 113137 145115 113245 145205
rect 106100 145025 113245 145115
rect 106100 144935 106207 145025
rect 106297 144935 106387 145025
rect 106477 144935 106567 145025
rect 106657 144935 106747 145025
rect 106837 144935 106927 145025
rect 107017 144935 107107 145025
rect 107197 144935 107287 145025
rect 107377 144935 107467 145025
rect 107557 144935 107647 145025
rect 107737 144935 107827 145025
rect 107917 144935 108007 145025
rect 108097 144935 108187 145025
rect 108277 144935 108367 145025
rect 108457 144935 108547 145025
rect 108637 144935 108727 145025
rect 108817 144935 108907 145025
rect 108997 144935 109087 145025
rect 109177 144935 109267 145025
rect 109357 144935 109447 145025
rect 109537 144935 109627 145025
rect 109717 144935 109807 145025
rect 109897 144935 109987 145025
rect 110077 144935 110167 145025
rect 110257 144935 110347 145025
rect 110437 144935 110527 145025
rect 110617 144935 110707 145025
rect 110797 144935 110887 145025
rect 110977 144935 111067 145025
rect 111157 144935 111247 145025
rect 111337 144935 111427 145025
rect 111517 144935 111607 145025
rect 111697 144935 111787 145025
rect 111877 144935 111967 145025
rect 112057 144935 112147 145025
rect 112237 144935 112327 145025
rect 112417 144935 112507 145025
rect 112597 144935 112687 145025
rect 112777 144935 112867 145025
rect 112957 144935 113047 145025
rect 113137 144935 113245 145025
rect 106100 144845 113245 144935
rect 106100 144755 106207 144845
rect 106297 144755 106387 144845
rect 106477 144755 106567 144845
rect 106657 144755 106747 144845
rect 106837 144755 106927 144845
rect 107017 144755 107107 144845
rect 107197 144755 107287 144845
rect 107377 144755 107467 144845
rect 107557 144755 107647 144845
rect 107737 144755 107827 144845
rect 107917 144755 108007 144845
rect 108097 144755 108187 144845
rect 108277 144755 108367 144845
rect 108457 144755 108547 144845
rect 108637 144755 108727 144845
rect 108817 144755 108907 144845
rect 108997 144755 109087 144845
rect 109177 144755 109267 144845
rect 109357 144755 109447 144845
rect 109537 144755 109627 144845
rect 109717 144755 109807 144845
rect 109897 144755 109987 144845
rect 110077 144755 110167 144845
rect 110257 144755 110347 144845
rect 110437 144755 110527 144845
rect 110617 144755 110707 144845
rect 110797 144755 110887 144845
rect 110977 144755 111067 144845
rect 111157 144755 111247 144845
rect 111337 144755 111427 144845
rect 111517 144755 111607 144845
rect 111697 144755 111787 144845
rect 111877 144755 111967 144845
rect 112057 144755 112147 144845
rect 112237 144755 112327 144845
rect 112417 144755 112507 144845
rect 112597 144755 112687 144845
rect 112777 144755 112867 144845
rect 112957 144755 113047 144845
rect 113137 144755 113245 144845
rect 106100 144665 113245 144755
rect 106100 144575 106207 144665
rect 106297 144575 106387 144665
rect 106477 144575 106567 144665
rect 106657 144575 106747 144665
rect 106837 144575 106927 144665
rect 107017 144575 107107 144665
rect 107197 144575 107287 144665
rect 107377 144575 107467 144665
rect 107557 144575 107647 144665
rect 107737 144575 107827 144665
rect 107917 144575 108007 144665
rect 108097 144575 108187 144665
rect 108277 144575 108367 144665
rect 108457 144575 108547 144665
rect 108637 144575 108727 144665
rect 108817 144575 108907 144665
rect 108997 144575 109087 144665
rect 109177 144575 109267 144665
rect 109357 144575 109447 144665
rect 109537 144575 109627 144665
rect 109717 144575 109807 144665
rect 109897 144575 109987 144665
rect 110077 144575 110167 144665
rect 110257 144575 110347 144665
rect 110437 144575 110527 144665
rect 110617 144575 110707 144665
rect 110797 144575 110887 144665
rect 110977 144575 111067 144665
rect 111157 144575 111247 144665
rect 111337 144575 111427 144665
rect 111517 144575 111607 144665
rect 111697 144575 111787 144665
rect 111877 144575 111967 144665
rect 112057 144575 112147 144665
rect 112237 144575 112327 144665
rect 112417 144575 112507 144665
rect 112597 144575 112687 144665
rect 112777 144575 112867 144665
rect 112957 144575 113047 144665
rect 113137 144575 113245 144665
rect 106100 144500 113245 144575
rect 88400 141260 89820 141350
rect 88400 141170 88525 141260
rect 88615 141170 88705 141260
rect 88795 141170 88885 141260
rect 88975 141170 89065 141260
rect 89155 141170 89245 141260
rect 89335 141170 89425 141260
rect 89515 141170 89605 141260
rect 89695 141170 89820 141260
rect 88400 141080 89820 141170
rect 88400 140990 88525 141080
rect 88615 140990 88705 141080
rect 88795 140990 88885 141080
rect 88975 140990 89065 141080
rect 89155 140990 89245 141080
rect 89335 140990 89425 141080
rect 89515 140990 89605 141080
rect 89695 140990 89820 141080
rect 88400 140900 89820 140990
rect 101700 144080 102440 144200
rect 101700 143990 101845 144080
rect 101935 143990 102025 144080
rect 102115 143990 102205 144080
rect 102295 143990 102440 144080
rect 101700 143900 102440 143990
rect 101700 143810 101845 143900
rect 101935 143810 102025 143900
rect 102115 143810 102205 143900
rect 102295 143810 102440 143900
rect 101700 143720 102440 143810
rect 101700 143630 101845 143720
rect 101935 143630 102025 143720
rect 102115 143630 102205 143720
rect 102295 143630 102440 143720
rect 101700 143540 102440 143630
rect 101700 143450 101845 143540
rect 101935 143450 102025 143540
rect 102115 143450 102205 143540
rect 102295 143450 102440 143540
rect 101700 143360 102440 143450
rect 101700 143270 101845 143360
rect 101935 143270 102025 143360
rect 102115 143270 102205 143360
rect 102295 143270 102440 143360
rect 101700 143180 102440 143270
rect 101700 143090 101845 143180
rect 101935 143090 102025 143180
rect 102115 143090 102205 143180
rect 102295 143090 102440 143180
rect 101700 140800 102440 143090
rect 103800 144125 104500 144200
rect 103800 144035 103925 144125
rect 104015 144035 104105 144125
rect 104195 144035 104285 144125
rect 104375 144035 104500 144125
rect 103800 143945 104500 144035
rect 103800 143855 103925 143945
rect 104015 143855 104105 143945
rect 104195 143855 104285 143945
rect 104375 143855 104500 143945
rect 103800 143765 104500 143855
rect 103800 143675 103925 143765
rect 104015 143675 104105 143765
rect 104195 143675 104285 143765
rect 104375 143675 104500 143765
rect 103800 143585 104500 143675
rect 103800 143495 103925 143585
rect 104015 143495 104105 143585
rect 104195 143495 104285 143585
rect 104375 143495 104500 143585
rect 103800 143405 104500 143495
rect 103800 143315 103925 143405
rect 104015 143315 104105 143405
rect 104195 143315 104285 143405
rect 104375 143315 104500 143405
rect 103800 143225 104500 143315
rect 103800 143135 103925 143225
rect 104015 143135 104105 143225
rect 104195 143135 104285 143225
rect 104375 143135 104500 143225
rect 103800 140800 104500 143135
rect 116500 141800 116820 145940
rect 130000 143100 130320 145940
rect 130000 142400 135745 143100
rect 116500 141100 133045 141800
rect 135300 141000 135745 142400
rect 44060 129880 45500 130200
rect 44060 116380 44900 116700
rect 44500 105272 44900 116380
rect 45100 105872 45500 129880
rect 144900 130000 145940 130320
rect 144400 116725 144650 116820
rect 144400 116635 144480 116725
rect 144570 116635 144650 116725
rect 144400 116545 144650 116635
rect 144400 116455 144480 116545
rect 144570 116455 144650 116545
rect 143440 116155 143860 116260
rect 143440 116065 143515 116155
rect 143605 116065 143695 116155
rect 143785 116065 143860 116155
rect 143440 115885 143860 116065
rect 143440 115795 143515 115885
rect 143605 115795 143695 115885
rect 143785 115795 143860 115885
rect 143440 115705 143860 115795
rect 143440 115615 143515 115705
rect 143605 115615 143695 115705
rect 143785 115615 143860 115705
rect 143440 115540 143860 115615
rect 143650 114382 143860 114460
rect 143650 114292 143710 114382
rect 143800 114292 143860 114382
rect 143650 114202 143860 114292
rect 143650 114112 143710 114202
rect 143800 114112 143860 114202
rect 143650 113530 143860 114112
rect 143650 113470 144075 113530
rect 143650 113380 143727 113470
rect 143817 113380 143907 113470
rect 143997 113380 144075 113470
rect 143650 113320 144075 113380
rect 45100 105782 45165 105872
rect 45255 105782 45345 105872
rect 45435 105782 45500 105872
rect 45100 105640 45500 105782
rect 44500 105182 44565 105272
rect 44655 105182 44745 105272
rect 44835 105182 44900 105272
rect 44500 105160 44900 105182
rect 44500 105040 45720 105160
rect 44500 104417 44900 104560
rect 44500 104327 44565 104417
rect 44655 104327 44745 104417
rect 44835 104327 44900 104417
rect 44500 103200 44900 104327
rect 44060 102880 44900 103200
rect 45100 103840 45996 103960
rect 45100 103817 45500 103840
rect 45100 103727 45165 103817
rect 45255 103727 45345 103817
rect 45435 103727 45500 103817
rect 45100 102500 45500 103727
rect 44500 102100 45500 102500
rect 44500 89699 44900 102100
rect 44060 89379 44900 89699
rect 42300 84790 46530 84930
rect 42300 84700 45777 84790
rect 45867 84700 45957 84790
rect 46047 84700 46137 84790
rect 46227 84700 46317 84790
rect 46407 84700 46530 84790
rect 42300 84610 46530 84700
rect 42300 84520 45777 84610
rect 45867 84520 45957 84610
rect 46047 84520 46137 84610
rect 46227 84520 46317 84610
rect 46407 84520 46530 84610
rect 42300 84430 46530 84520
rect 42300 84340 45777 84430
rect 45867 84340 45957 84430
rect 46047 84340 46137 84430
rect 46227 84340 46317 84430
rect 46407 84340 46530 84430
rect 42300 84250 46530 84340
rect 42300 84160 45777 84250
rect 45867 84160 45957 84250
rect 46047 84160 46137 84250
rect 46227 84160 46317 84250
rect 46407 84160 46530 84250
rect 42300 84070 46530 84160
rect 42300 83980 45777 84070
rect 45867 83980 45957 84070
rect 46047 83980 46137 84070
rect 46227 83980 46317 84070
rect 46407 83980 46530 84070
rect 42300 83890 46530 83980
rect 42300 83800 45777 83890
rect 45867 83800 45957 83890
rect 46047 83800 46137 83890
rect 46227 83800 46317 83890
rect 46407 83800 46530 83890
rect 42300 83710 46530 83800
rect 42300 83620 45777 83710
rect 45867 83620 45957 83710
rect 46047 83620 46137 83710
rect 46227 83620 46317 83710
rect 46407 83620 46530 83710
rect 42300 83530 46530 83620
rect 42300 83440 45777 83530
rect 45867 83440 45957 83530
rect 46047 83440 46137 83530
rect 46227 83440 46317 83530
rect 46407 83440 46530 83530
rect 42300 83350 46530 83440
rect 42300 83260 45777 83350
rect 45867 83260 45957 83350
rect 46047 83260 46137 83350
rect 46227 83260 46317 83350
rect 46407 83260 46530 83350
rect 42300 83170 46530 83260
rect 42300 83080 45777 83170
rect 45867 83080 45957 83170
rect 46047 83080 46137 83170
rect 46227 83080 46317 83170
rect 46407 83080 46530 83170
rect 42300 82990 46530 83080
rect 42300 82900 45777 82990
rect 45867 82900 45957 82990
rect 46047 82900 46137 82990
rect 46227 82900 46317 82990
rect 46407 82900 46530 82990
rect 42300 82810 46530 82900
rect 42300 82720 45777 82810
rect 45867 82720 45957 82810
rect 46047 82720 46137 82810
rect 46227 82720 46317 82810
rect 46407 82720 46530 82810
rect 42300 82630 46530 82720
rect 42300 82540 45777 82630
rect 45867 82540 45957 82630
rect 46047 82540 46137 82630
rect 46227 82540 46317 82630
rect 46407 82540 46530 82630
rect 42300 82450 46530 82540
rect 42300 82360 45777 82450
rect 45867 82360 45957 82450
rect 46047 82360 46137 82450
rect 46227 82360 46317 82450
rect 46407 82360 46530 82450
rect 42300 82270 46530 82360
rect 42300 82180 45777 82270
rect 45867 82180 45957 82270
rect 46047 82180 46137 82270
rect 46227 82180 46317 82270
rect 46407 82180 46530 82270
rect 42300 82090 46530 82180
rect 42300 82000 45777 82090
rect 45867 82000 45957 82090
rect 46047 82000 46137 82090
rect 46227 82000 46317 82090
rect 46407 82000 46530 82090
rect 42300 81910 46530 82000
rect 42300 81820 45777 81910
rect 45867 81820 45957 81910
rect 46047 81820 46137 81910
rect 46227 81820 46317 81910
rect 46407 81820 46530 81910
rect 42300 81730 46530 81820
rect 42300 81640 45777 81730
rect 45867 81640 45957 81730
rect 46047 81640 46137 81730
rect 46227 81640 46317 81730
rect 46407 81640 46530 81730
rect 42300 81550 46530 81640
rect 42300 81460 45777 81550
rect 45867 81460 45957 81550
rect 46047 81460 46137 81550
rect 46227 81460 46317 81550
rect 46407 81460 46530 81550
rect 42300 81370 46530 81460
rect 42300 81280 45777 81370
rect 45867 81280 45957 81370
rect 46047 81280 46137 81370
rect 46227 81280 46317 81370
rect 46407 81280 46530 81370
rect 42300 81190 46530 81280
rect 42300 81100 45777 81190
rect 45867 81100 45957 81190
rect 46047 81100 46137 81190
rect 46227 81100 46317 81190
rect 46407 81100 46530 81190
rect 42300 81010 46530 81100
rect 42300 80920 45777 81010
rect 45867 80920 45957 81010
rect 46047 80920 46137 81010
rect 46227 80920 46317 81010
rect 46407 80920 46530 81010
rect 42300 80830 46530 80920
rect 42300 80740 45777 80830
rect 45867 80740 45957 80830
rect 46047 80740 46137 80830
rect 46227 80740 46317 80830
rect 46407 80740 46530 80830
rect 42300 80650 46530 80740
rect 42300 80560 45777 80650
rect 45867 80560 45957 80650
rect 46047 80560 46137 80650
rect 46227 80560 46317 80650
rect 46407 80560 46530 80650
rect 42300 80470 46530 80560
rect 42300 80380 45777 80470
rect 45867 80380 45957 80470
rect 46047 80380 46137 80470
rect 46227 80380 46317 80470
rect 46407 80380 46530 80470
rect 42300 80290 46530 80380
rect 42300 80200 45777 80290
rect 45867 80200 45957 80290
rect 46047 80200 46137 80290
rect 46227 80200 46317 80290
rect 46407 80200 46530 80290
rect 42300 80110 46530 80200
rect 42300 80020 45777 80110
rect 45867 80020 45957 80110
rect 46047 80020 46137 80110
rect 46227 80020 46317 80110
rect 46407 80020 46530 80110
rect 42300 79930 46530 80020
rect 42300 79840 45777 79930
rect 45867 79840 45957 79930
rect 46047 79840 46137 79930
rect 46227 79840 46317 79930
rect 46407 79840 46530 79930
rect 42300 79750 46530 79840
rect 42300 79660 45777 79750
rect 45867 79660 45957 79750
rect 46047 79660 46137 79750
rect 46227 79660 46317 79750
rect 46407 79660 46530 79750
rect 42300 79570 46530 79660
rect 42300 79480 45777 79570
rect 45867 79480 45957 79570
rect 46047 79480 46137 79570
rect 46227 79480 46317 79570
rect 46407 79480 46530 79570
rect 42300 79390 46530 79480
rect 42300 79300 45777 79390
rect 45867 79300 45957 79390
rect 46047 79300 46137 79390
rect 46227 79300 46317 79390
rect 46407 79300 46530 79390
rect 42300 79210 46530 79300
rect 42300 79120 45777 79210
rect 45867 79120 45957 79210
rect 46047 79120 46137 79210
rect 46227 79120 46317 79210
rect 46407 79120 46530 79210
rect 42300 79030 46530 79120
rect 42300 78940 45777 79030
rect 45867 78940 45957 79030
rect 46047 78940 46137 79030
rect 46227 78940 46317 79030
rect 46407 78940 46530 79030
rect 42300 78850 46530 78940
rect 42300 78760 45777 78850
rect 45867 78760 45957 78850
rect 46047 78760 46137 78850
rect 46227 78760 46317 78850
rect 46407 78760 46530 78850
rect 42300 78670 46530 78760
rect 42300 78580 45777 78670
rect 45867 78580 45957 78670
rect 46047 78580 46137 78670
rect 46227 78580 46317 78670
rect 46407 78580 46530 78670
rect 42300 78490 46530 78580
rect 42300 78400 45777 78490
rect 45867 78400 45957 78490
rect 46047 78400 46137 78490
rect 46227 78400 46317 78490
rect 46407 78400 46530 78490
rect 42300 78310 46530 78400
rect 42300 78220 45777 78310
rect 45867 78220 45957 78310
rect 46047 78220 46137 78310
rect 46227 78220 46317 78310
rect 46407 78220 46530 78310
rect 42300 78080 46530 78220
rect 44500 76285 46360 76360
rect 44500 76195 46022 76285
rect 46112 76195 46202 76285
rect 46292 76195 46360 76285
rect 44500 76105 46360 76195
rect 44500 76015 46022 76105
rect 46112 76015 46202 76105
rect 46292 76015 46360 76105
rect 44500 75940 46360 76015
rect 44500 62700 44900 75940
rect 44060 62380 44900 62700
rect 143690 59730 143900 59815
rect 143690 59640 143750 59730
rect 143840 59640 143900 59730
rect 143690 59585 143900 59640
rect 144400 59585 144650 116455
rect 143690 59550 144650 59585
rect 143690 59460 143750 59550
rect 143840 59460 144650 59550
rect 143690 59375 144650 59460
rect 144900 57255 145150 130000
rect 145440 116705 145940 116820
rect 145440 116615 145555 116705
rect 145645 116615 145735 116705
rect 145825 116615 145940 116705
rect 145440 116500 145940 116615
rect 145400 103205 145940 103320
rect 145400 103115 145535 103205
rect 145625 103115 145715 103205
rect 145805 103115 145940 103205
rect 145400 103000 145940 103115
rect 145650 100827 145940 100905
rect 145650 100737 145750 100827
rect 145840 100737 145940 100827
rect 145650 100647 145940 100737
rect 145650 100557 145750 100647
rect 145840 100557 145940 100647
rect 145650 100467 145940 100557
rect 145650 100377 145750 100467
rect 145840 100377 145940 100467
rect 145650 100300 145940 100377
rect 145395 87005 145940 87120
rect 145395 86915 145532 87005
rect 145622 86915 145712 87005
rect 145802 86915 145940 87005
rect 145395 86800 145940 86915
rect 145360 73505 145940 73620
rect 145360 73415 145425 73505
rect 145515 73415 145605 73505
rect 145695 73415 145785 73505
rect 145875 73415 145940 73505
rect 145360 73300 145940 73415
rect 145545 60005 145940 60120
rect 145545 59915 145607 60005
rect 145697 59915 145787 60005
rect 145877 59915 145940 60005
rect 145545 59800 145940 59915
rect 143740 57192 145150 57255
rect 143740 57102 143865 57192
rect 143955 57102 144045 57192
rect 144135 57102 145150 57192
rect 143740 57040 145150 57102
rect 145400 56675 145650 56820
rect 145400 56655 145480 56675
rect 143740 56592 145480 56655
rect 143740 56502 143865 56592
rect 143955 56502 144045 56592
rect 144135 56585 145480 56592
rect 145570 56585 145650 56675
rect 144135 56502 145650 56585
rect 143740 56440 145650 56502
rect 45100 49282 45500 49415
rect 45100 49200 45165 49282
rect 44060 49192 45165 49200
rect 45255 49192 45345 49282
rect 45435 49192 45500 49282
rect 44060 49102 45500 49192
rect 44060 49012 45165 49102
rect 45255 49012 45345 49102
rect 45435 49012 45500 49102
rect 44060 48880 45500 49012
rect 99600 46402 100050 46475
rect 59800 45807 60120 45900
rect 59800 45717 59915 45807
rect 60005 45717 60120 45807
rect 59800 45627 60120 45717
rect 59800 45537 59915 45627
rect 60005 45537 60120 45627
rect 59800 44060 60120 45537
rect 67540 45000 67645 46265
rect 94240 45600 94505 46345
rect 94840 46200 94945 46365
rect 99600 46312 99690 46402
rect 99780 46312 99870 46402
rect 99960 46312 100050 46402
rect 99600 46240 100050 46312
rect 94840 46095 95325 46200
rect 94840 46005 94947 46095
rect 95037 46005 95127 46095
rect 95217 46005 95325 46095
rect 94840 45900 95325 46005
rect 106840 45900 106945 46350
rect 106555 45795 106945 45900
rect 106555 45705 106615 45795
rect 106705 45705 106795 45795
rect 106885 45705 106945 45795
rect 106555 45600 106945 45705
rect 94240 45495 94725 45600
rect 94240 45405 94347 45495
rect 94437 45405 94527 45495
rect 94617 45405 94725 45495
rect 94240 45300 94725 45405
rect 107440 45300 107545 46285
rect 73300 45195 73620 45300
rect 73300 45105 73415 45195
rect 73505 45105 73620 45195
rect 67540 44895 68070 45000
rect 67540 44805 67670 44895
rect 67760 44805 67850 44895
rect 67940 44805 68070 44895
rect 67540 44700 68070 44805
rect 73300 44135 73620 45105
rect 99600 45000 107545 45300
rect 99600 44400 99900 45000
rect 108640 44400 108745 46465
rect 140800 46122 141120 46200
rect 140800 46032 140915 46122
rect 141005 46032 141120 46122
rect 140800 45942 141120 46032
rect 140800 45852 140915 45942
rect 141005 45852 141120 45942
rect 127300 45535 127620 45600
rect 127300 45445 127415 45535
rect 127505 45445 127620 45535
rect 127300 45355 127620 45445
rect 127300 45265 127415 45355
rect 127505 45265 127620 45355
rect 86800 44100 99900 44400
rect 100300 44100 108745 44400
rect 113800 44902 114120 45000
rect 113800 44812 113915 44902
rect 114005 44812 114120 44902
rect 113800 44722 114120 44812
rect 113800 44632 113915 44722
rect 114005 44632 114120 44722
rect 113800 44060 114120 44632
rect 127300 44060 127620 45265
rect 140800 44060 141120 45852
<< m3contact >>
rect 49067 145330 49157 145420
rect 49247 145330 49337 145420
rect 49427 145330 49517 145420
rect 49607 145330 49697 145420
rect 49787 145330 49877 145420
rect 49967 145330 50057 145420
rect 50147 145330 50237 145420
rect 50327 145330 50417 145420
rect 50507 145330 50597 145420
rect 50687 145330 50777 145420
rect 49067 145150 49157 145240
rect 49247 145150 49337 145240
rect 49427 145150 49517 145240
rect 49607 145150 49697 145240
rect 49787 145150 49877 145240
rect 49967 145150 50057 145240
rect 50147 145150 50237 145240
rect 50327 145150 50417 145240
rect 50507 145150 50597 145240
rect 50687 145150 50777 145240
rect 49067 144970 49157 145060
rect 49247 144970 49337 145060
rect 49427 144970 49517 145060
rect 49607 144970 49697 145060
rect 49787 144970 49877 145060
rect 49967 144970 50057 145060
rect 50147 144970 50237 145060
rect 50327 144970 50417 145060
rect 50507 144970 50597 145060
rect 50687 144970 50777 145060
rect 49067 144790 49157 144880
rect 49247 144790 49337 144880
rect 49427 144790 49517 144880
rect 49607 144790 49697 144880
rect 49787 144790 49877 144880
rect 49967 144790 50057 144880
rect 50147 144790 50237 144880
rect 50327 144790 50417 144880
rect 50507 144790 50597 144880
rect 50687 144790 50777 144880
rect 62622 144027 62712 144117
rect 62802 144027 62892 144117
rect 62982 144027 63072 144117
rect 63162 144027 63252 144117
rect 63342 144027 63432 144117
rect 63522 144027 63612 144117
rect 63702 144027 63792 144117
rect 63882 144027 63972 144117
rect 64062 144027 64152 144117
rect 64242 144027 64332 144117
rect 62622 143847 62712 143937
rect 62802 143847 62892 143937
rect 62982 143847 63072 143937
rect 63162 143847 63252 143937
rect 63342 143847 63432 143937
rect 63522 143847 63612 143937
rect 63702 143847 63792 143937
rect 63882 143847 63972 143937
rect 64062 143847 64152 143937
rect 64242 143847 64332 143937
rect 62622 143667 62712 143757
rect 62802 143667 62892 143757
rect 62982 143667 63072 143757
rect 63162 143667 63252 143757
rect 63342 143667 63432 143757
rect 63522 143667 63612 143757
rect 63702 143667 63792 143757
rect 63882 143667 63972 143757
rect 64062 143667 64152 143757
rect 64242 143667 64332 143757
rect 62622 143487 62712 143577
rect 62802 143487 62892 143577
rect 62982 143487 63072 143577
rect 63162 143487 63252 143577
rect 63342 143487 63432 143577
rect 63522 143487 63612 143577
rect 63702 143487 63792 143577
rect 63882 143487 63972 143577
rect 64062 143487 64152 143577
rect 64242 143487 64332 143577
rect 77985 141170 78075 141260
rect 78165 141170 78255 141260
rect 78345 141170 78435 141260
rect 78525 141170 78615 141260
rect 77985 140990 78075 141080
rect 78165 140990 78255 141080
rect 78345 140990 78435 141080
rect 78525 140990 78615 141080
rect 88525 141170 88615 141260
rect 88705 141170 88795 141260
rect 88885 141170 88975 141260
rect 89065 141170 89155 141260
rect 89245 141170 89335 141260
rect 89425 141170 89515 141260
rect 89605 141170 89695 141260
rect 88525 140990 88615 141080
rect 88705 140990 88795 141080
rect 88885 140990 88975 141080
rect 89065 140990 89155 141080
rect 89245 140990 89335 141080
rect 89425 140990 89515 141080
rect 89605 140990 89695 141080
rect 101845 143990 101935 144080
rect 102025 143990 102115 144080
rect 102205 143990 102295 144080
rect 101845 143810 101935 143900
rect 102025 143810 102115 143900
rect 102205 143810 102295 143900
rect 101845 143630 101935 143720
rect 102025 143630 102115 143720
rect 102205 143630 102295 143720
rect 101845 143450 101935 143540
rect 102025 143450 102115 143540
rect 102205 143450 102295 143540
rect 101845 143270 101935 143360
rect 102025 143270 102115 143360
rect 102205 143270 102295 143360
rect 101845 143090 101935 143180
rect 102025 143090 102115 143180
rect 102205 143090 102295 143180
rect 103925 144035 104015 144125
rect 104105 144035 104195 144125
rect 104285 144035 104375 144125
rect 103925 143855 104015 143945
rect 104105 143855 104195 143945
rect 104285 143855 104375 143945
rect 103925 143675 104015 143765
rect 104105 143675 104195 143765
rect 104285 143675 104375 143765
rect 103925 143495 104015 143585
rect 104105 143495 104195 143585
rect 104285 143495 104375 143585
rect 103925 143315 104015 143405
rect 104105 143315 104195 143405
rect 104285 143315 104375 143405
rect 103925 143135 104015 143225
rect 104105 143135 104195 143225
rect 104285 143135 104375 143225
rect 144480 116635 144570 116725
rect 144480 116455 144570 116545
rect 143515 115795 143605 115885
rect 143695 115795 143785 115885
rect 143515 115615 143605 115705
rect 143695 115615 143785 115705
rect 143710 114292 143800 114382
rect 143710 114112 143800 114202
rect 143727 113380 143817 113470
rect 143907 113380 143997 113470
rect 45165 105782 45255 105872
rect 45345 105782 45435 105872
rect 44565 105182 44655 105272
rect 44745 105182 44835 105272
rect 44565 104327 44655 104417
rect 44745 104327 44835 104417
rect 45165 103727 45255 103817
rect 45345 103727 45435 103817
rect 46022 76195 46112 76285
rect 46202 76195 46292 76285
rect 46022 76015 46112 76105
rect 46202 76015 46292 76105
rect 143750 59640 143840 59730
rect 143750 59460 143840 59550
rect 145555 116615 145645 116705
rect 145735 116615 145825 116705
rect 145750 100737 145840 100827
rect 145750 100557 145840 100647
rect 145750 100377 145840 100467
rect 145532 86915 145622 87005
rect 145712 86915 145802 87005
rect 145425 73415 145515 73505
rect 145605 73415 145695 73505
rect 145785 73415 145875 73505
rect 145607 59915 145697 60005
rect 145787 59915 145877 60005
rect 143865 57102 143955 57192
rect 144045 57102 144135 57192
rect 143865 56502 143955 56592
rect 144045 56502 144135 56592
rect 45165 49192 45255 49282
rect 45345 49192 45435 49282
rect 45165 49012 45255 49102
rect 45345 49012 45435 49102
rect 94947 46005 95037 46095
rect 95127 46005 95217 46095
rect 94347 45405 94437 45495
rect 94527 45405 94617 45495
rect 67670 44805 67760 44895
rect 67850 44805 67940 44895
rect 140915 46032 141005 46122
rect 140915 45852 141005 45942
rect 127415 45445 127505 45535
rect 127415 45265 127505 45355
rect 113915 44812 114005 44902
rect 113915 44632 114005 44722
<< metal3 >>
rect 49000 145500 50845 145510
rect 49000 145420 104500 145500
rect 49000 145330 49067 145420
rect 49157 145330 49247 145420
rect 49337 145330 49427 145420
rect 49517 145330 49607 145420
rect 49697 145330 49787 145420
rect 49877 145330 49967 145420
rect 50057 145330 50147 145420
rect 50237 145330 50327 145420
rect 50417 145330 50507 145420
rect 50597 145330 50687 145420
rect 50777 145330 104500 145420
rect 49000 145240 104500 145330
rect 49000 145150 49067 145240
rect 49157 145150 49247 145240
rect 49337 145150 49427 145240
rect 49517 145150 49607 145240
rect 49697 145150 49787 145240
rect 49877 145150 49967 145240
rect 50057 145150 50147 145240
rect 50237 145150 50327 145240
rect 50417 145150 50507 145240
rect 50597 145150 50687 145240
rect 50777 145150 104500 145240
rect 49000 145060 104500 145150
rect 49000 144970 49067 145060
rect 49157 144970 49247 145060
rect 49337 144970 49427 145060
rect 49517 144970 49607 145060
rect 49697 144970 49787 145060
rect 49877 144970 49967 145060
rect 50057 144970 50147 145060
rect 50237 144970 50327 145060
rect 50417 144970 50507 145060
rect 50597 144970 50687 145060
rect 50777 144970 104500 145060
rect 49000 144880 104500 144970
rect 49000 144790 49067 144880
rect 49157 144790 49247 144880
rect 49337 144790 49427 144880
rect 49517 144790 49607 144880
rect 49697 144790 49787 144880
rect 49877 144790 49967 144880
rect 50057 144790 50147 144880
rect 50237 144790 50327 144880
rect 50417 144790 50507 144880
rect 50597 144790 50687 144880
rect 50777 144790 104500 144880
rect 49000 144700 104500 144790
rect 62500 144200 64455 144205
rect 62500 144117 102440 144200
rect 62500 144027 62622 144117
rect 62712 144027 62802 144117
rect 62892 144027 62982 144117
rect 63072 144027 63162 144117
rect 63252 144027 63342 144117
rect 63432 144027 63522 144117
rect 63612 144027 63702 144117
rect 63792 144027 63882 144117
rect 63972 144027 64062 144117
rect 64152 144027 64242 144117
rect 64332 144080 102440 144117
rect 64332 144027 101845 144080
rect 62500 143990 101845 144027
rect 101935 143990 102025 144080
rect 102115 143990 102205 144080
rect 102295 143990 102440 144080
rect 62500 143937 102440 143990
rect 62500 143847 62622 143937
rect 62712 143847 62802 143937
rect 62892 143847 62982 143937
rect 63072 143847 63162 143937
rect 63252 143847 63342 143937
rect 63432 143847 63522 143937
rect 63612 143847 63702 143937
rect 63792 143847 63882 143937
rect 63972 143847 64062 143937
rect 64152 143847 64242 143937
rect 64332 143900 102440 143937
rect 64332 143847 101845 143900
rect 62500 143810 101845 143847
rect 101935 143810 102025 143900
rect 102115 143810 102205 143900
rect 102295 143810 102440 143900
rect 62500 143757 102440 143810
rect 62500 143667 62622 143757
rect 62712 143667 62802 143757
rect 62892 143667 62982 143757
rect 63072 143667 63162 143757
rect 63252 143667 63342 143757
rect 63432 143667 63522 143757
rect 63612 143667 63702 143757
rect 63792 143667 63882 143757
rect 63972 143667 64062 143757
rect 64152 143667 64242 143757
rect 64332 143720 102440 143757
rect 64332 143667 101845 143720
rect 62500 143630 101845 143667
rect 101935 143630 102025 143720
rect 102115 143630 102205 143720
rect 102295 143630 102440 143720
rect 62500 143577 102440 143630
rect 62500 143487 62622 143577
rect 62712 143487 62802 143577
rect 62892 143487 62982 143577
rect 63072 143487 63162 143577
rect 63252 143487 63342 143577
rect 63432 143487 63522 143577
rect 63612 143487 63702 143577
rect 63792 143487 63882 143577
rect 63972 143487 64062 143577
rect 64152 143487 64242 143577
rect 64332 143540 102440 143577
rect 64332 143487 101845 143540
rect 62500 143450 101845 143487
rect 101935 143450 102025 143540
rect 102115 143450 102205 143540
rect 102295 143450 102440 143540
rect 62500 143400 102440 143450
rect 101700 143360 102440 143400
rect 101700 143270 101845 143360
rect 101935 143270 102025 143360
rect 102115 143270 102205 143360
rect 102295 143270 102440 143360
rect 101700 143180 102440 143270
rect 101700 143090 101845 143180
rect 101935 143090 102025 143180
rect 102115 143090 102205 143180
rect 102295 143090 102440 143180
rect 101700 142970 102440 143090
rect 103800 144125 104500 144700
rect 103800 144035 103925 144125
rect 104015 144035 104105 144125
rect 104195 144035 104285 144125
rect 104375 144035 104500 144125
rect 103800 143945 104500 144035
rect 103800 143855 103925 143945
rect 104015 143855 104105 143945
rect 104195 143855 104285 143945
rect 104375 143855 104500 143945
rect 103800 143765 104500 143855
rect 103800 143675 103925 143765
rect 104015 143675 104105 143765
rect 104195 143675 104285 143765
rect 104375 143675 104500 143765
rect 103800 143585 104500 143675
rect 103800 143495 103925 143585
rect 104015 143495 104105 143585
rect 104195 143495 104285 143585
rect 104375 143495 104500 143585
rect 103800 143405 104500 143495
rect 103800 143315 103925 143405
rect 104015 143315 104105 143405
rect 104195 143315 104285 143405
rect 104375 143315 104500 143405
rect 103800 143225 104500 143315
rect 103800 143135 103925 143225
rect 104015 143135 104105 143225
rect 104195 143135 104285 143225
rect 104375 143135 104500 143225
rect 103800 143060 104500 143135
rect 77850 141260 89820 141350
rect 77850 141170 77985 141260
rect 78075 141170 78165 141260
rect 78255 141170 78345 141260
rect 78435 141170 78525 141260
rect 78615 141170 88525 141260
rect 88615 141170 88705 141260
rect 88795 141170 88885 141260
rect 88975 141170 89065 141260
rect 89155 141170 89245 141260
rect 89335 141170 89425 141260
rect 89515 141170 89605 141260
rect 89695 141170 89820 141260
rect 77850 141080 89820 141170
rect 77850 140990 77985 141080
rect 78075 140990 78165 141080
rect 78255 140990 78345 141080
rect 78435 140990 78525 141080
rect 78615 140990 88525 141080
rect 88615 140990 88705 141080
rect 88795 140990 88885 141080
rect 88975 140990 89065 141080
rect 89155 140990 89245 141080
rect 89335 140990 89425 141080
rect 89515 140990 89605 141080
rect 89695 140990 89820 141080
rect 77850 140900 89820 140990
rect 144400 116725 145940 116820
rect 144400 116635 144480 116725
rect 144570 116705 145940 116725
rect 144570 116635 145555 116705
rect 144400 116615 145555 116635
rect 145645 116615 145735 116705
rect 145825 116615 145940 116705
rect 144400 116545 145940 116615
rect 144400 116455 144480 116545
rect 144570 116500 145940 116545
rect 144570 116455 144650 116500
rect 144400 116360 144650 116455
rect 143440 115885 143860 115960
rect 143440 115795 143515 115885
rect 143605 115795 143695 115885
rect 143785 115795 143860 115885
rect 143440 115705 143860 115795
rect 143440 115615 143515 115705
rect 143605 115615 143695 115705
rect 143785 115615 143860 115705
rect 143440 115540 143860 115615
rect 143650 114382 143860 114460
rect 143650 114292 143710 114382
rect 143800 114292 143860 114382
rect 143650 114202 143860 114292
rect 143650 114112 143710 114202
rect 143800 114112 143860 114202
rect 143650 114035 143860 114112
rect 144105 113740 145900 113950
rect 143650 113470 145400 113530
rect 143650 113380 143727 113470
rect 143817 113380 143907 113470
rect 143997 113380 145400 113470
rect 143650 113320 145400 113380
rect 143695 112240 144900 112360
rect 143840 111640 144400 111760
rect 45100 105872 45500 106015
rect 45100 105782 45165 105872
rect 45255 105782 45345 105872
rect 45435 105782 45500 105872
rect 45100 105760 45500 105782
rect 45100 105640 46315 105760
rect 44500 105272 44900 105415
rect 44500 105182 44565 105272
rect 44655 105182 44745 105272
rect 44835 105182 44900 105272
rect 44500 105160 44900 105182
rect 44500 105040 46590 105160
rect 44500 104440 46785 104560
rect 44500 104417 44900 104440
rect 44500 104327 44565 104417
rect 44655 104327 44745 104417
rect 44835 104327 44900 104417
rect 44500 104185 44900 104327
rect 45100 103840 46530 103960
rect 45100 103817 45500 103840
rect 45100 103727 45165 103817
rect 45255 103727 45345 103817
rect 45435 103727 45500 103817
rect 45100 103585 45500 103727
rect 45100 101440 47970 101561
rect 45100 49282 45500 101440
rect 45955 76285 46360 76360
rect 45955 76195 46022 76285
rect 46112 76195 46202 76285
rect 46292 76195 46360 76285
rect 45955 76105 46360 76195
rect 45955 76015 46022 76105
rect 46112 76015 46202 76105
rect 46292 76015 46360 76105
rect 45955 75940 46360 76015
rect 143690 59730 143900 60460
rect 144150 60120 144400 111640
rect 144650 73620 144900 112240
rect 145150 87120 145400 113320
rect 145650 100905 145900 113740
rect 145650 100827 145940 100905
rect 145650 100737 145750 100827
rect 145840 100737 145940 100827
rect 145650 100647 145940 100737
rect 145650 100557 145750 100647
rect 145840 100557 145940 100647
rect 145650 100467 145940 100557
rect 145650 100377 145750 100467
rect 145840 100377 145940 100467
rect 145650 100300 145940 100377
rect 145150 87005 145940 87120
rect 145150 86915 145532 87005
rect 145622 86915 145712 87005
rect 145802 86915 145940 87005
rect 145150 86800 145940 86915
rect 144650 73505 145940 73620
rect 144650 73415 145425 73505
rect 145515 73415 145605 73505
rect 145695 73415 145785 73505
rect 145875 73415 145940 73505
rect 144650 73300 145940 73415
rect 144150 60005 145940 60120
rect 144150 59915 145607 60005
rect 145697 59915 145787 60005
rect 145877 59915 145940 60005
rect 144150 59800 145940 59915
rect 143690 59640 143750 59730
rect 143840 59640 143900 59730
rect 143690 59550 143900 59640
rect 143690 59460 143750 59550
rect 143840 59460 143900 59550
rect 143690 59375 143900 59460
rect 143740 57192 144260 57255
rect 143740 57102 143865 57192
rect 143955 57102 144045 57192
rect 144135 57102 144260 57192
rect 143740 57040 144260 57102
rect 143740 56592 144260 56655
rect 143740 56502 143865 56592
rect 143955 56502 144045 56592
rect 144135 56502 144260 56592
rect 143740 56440 144260 56502
rect 45100 49192 45165 49282
rect 45255 49192 45345 49282
rect 45435 49192 45500 49282
rect 45100 49102 45500 49192
rect 45100 49012 45165 49102
rect 45255 49012 45345 49102
rect 45435 49012 45500 49102
rect 45100 48880 45500 49012
rect 94840 46122 141120 46200
rect 94840 46095 140915 46122
rect 94840 46005 94947 46095
rect 95037 46005 95127 46095
rect 95217 46032 140915 46095
rect 141005 46032 141120 46122
rect 95217 46005 141120 46032
rect 94840 45942 141120 46005
rect 94840 45900 140915 45942
rect 140800 45852 140915 45900
rect 141005 45852 141120 45942
rect 140800 45775 141120 45852
rect 94240 45535 127620 45600
rect 94240 45495 127415 45535
rect 94240 45405 94347 45495
rect 94437 45405 94527 45495
rect 94617 45445 127415 45495
rect 127505 45445 127620 45535
rect 94617 45405 127620 45445
rect 94240 45355 127620 45405
rect 94240 45300 127415 45355
rect 127300 45265 127415 45300
rect 127505 45265 127620 45355
rect 127300 45200 127620 45265
rect 67540 44902 114120 45000
rect 67540 44895 113915 44902
rect 67540 44805 67670 44895
rect 67760 44805 67850 44895
rect 67940 44812 113915 44895
rect 114005 44812 114120 44902
rect 67940 44805 114120 44812
rect 67540 44722 114120 44805
rect 67540 44700 113915 44722
rect 113800 44632 113915 44700
rect 114005 44632 114120 44722
rect 113800 44535 114120 44632
<< end >>
