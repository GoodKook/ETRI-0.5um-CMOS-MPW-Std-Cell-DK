magic
tech scmos
magscale 1 2
timestamp 1727424219
<< nwell >>
rect 87 272 112 273
rect -12 154 112 272
<< ntransistor >>
rect 20 14 24 54
rect 30 14 34 54
rect 50 14 54 54
<< ptransistor >>
rect 20 206 24 246
rect 42 206 46 246
rect 64 166 68 246
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 30 54
rect 34 14 36 54
rect 48 14 50 54
rect 54 14 56 54
<< pdiffusion >>
rect 18 206 20 246
rect 24 206 26 246
rect 38 206 42 246
rect 46 206 50 246
rect 62 166 64 246
rect 68 166 70 246
<< ndcontact >>
rect 6 14 18 54
rect 36 14 48 54
rect 56 14 68 54
<< pdcontact >>
rect 6 206 18 246
rect 26 206 38 246
rect 50 166 62 246
rect 70 166 82 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 20 246 24 250
rect 42 246 46 250
rect 64 246 68 250
rect 20 129 24 206
rect 16 117 24 129
rect 42 123 46 206
rect 20 54 24 117
rect 30 111 44 123
rect 30 54 34 111
rect 64 72 68 166
rect 56 60 68 72
rect 50 54 54 60
rect 20 10 24 14
rect 30 10 34 14
rect 50 10 54 14
<< polycontact >>
rect 4 117 16 129
rect 44 111 56 123
rect 44 60 56 72
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 6 246 18 252
rect 50 246 62 252
rect 3 103 17 117
rect 26 72 33 206
rect 43 123 57 137
rect 70 97 77 166
rect 63 83 77 97
rect 6 66 44 72
rect 6 54 18 66
rect 63 54 69 83
rect 68 42 69 54
rect 36 8 48 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect 43 123 57 137
rect 3 103 17 117
rect 63 83 77 97
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 63 83 77 97 0 Y
port 2 nsew signal output
rlabel metal1 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal1 43 123 57 137 0 B
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
