magic
tech scmos
magscale 1 2
timestamp 1702307383
<< nwell >>
rect -14 154 114 272
<< ntransistor >>
rect 22 14 26 54
rect 32 14 36 54
rect 52 14 56 54
rect 62 14 66 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 58 166 62 246
rect 78 166 82 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 32 54
rect 36 14 38 54
rect 50 14 52 54
rect 56 14 62 54
rect 66 14 68 54
<< pdiffusion >>
rect 16 169 18 246
rect 4 166 18 169
rect 22 181 24 246
rect 36 181 38 246
rect 22 166 38 181
rect 42 169 44 246
rect 56 169 58 246
rect 42 166 58 169
rect 62 234 78 246
rect 62 166 64 234
rect 76 166 78 234
rect 82 166 84 246
<< ndcontact >>
rect 8 14 20 54
rect 38 14 50 54
rect 68 14 80 54
<< pdcontact >>
rect 4 169 16 246
rect 24 181 36 246
rect 44 169 56 246
rect 64 166 76 234
rect 84 166 96 246
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 254 106 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 78 246 82 250
rect 18 144 22 166
rect 13 138 22 144
rect 13 117 18 138
rect 17 105 18 117
rect 13 63 18 105
rect 38 85 42 166
rect 58 94 62 166
rect 78 114 82 166
rect 78 102 83 114
rect 13 58 26 63
rect 22 54 26 58
rect 32 54 36 85
rect 52 82 58 94
rect 52 54 56 82
rect 78 63 82 102
rect 62 59 82 63
rect 62 54 66 59
rect 22 10 26 14
rect 32 10 36 14
rect 52 10 56 14
rect 62 10 66 14
<< polycontact >>
rect 5 105 17 117
rect 26 85 38 97
rect 83 102 95 114
rect 58 82 70 94
<< metal1 >>
rect -6 266 106 268
rect -6 252 106 254
rect 24 246 36 252
rect 16 169 44 175
rect 56 240 84 246
rect 64 161 76 166
rect 46 155 76 161
rect 46 137 54 155
rect 3 123 17 137
rect 43 123 57 137
rect 83 123 97 137
rect 5 117 17 123
rect 23 103 37 117
rect 26 97 37 103
rect 44 54 50 123
rect 63 103 77 117
rect 83 114 95 123
rect 63 94 74 103
rect 70 82 74 94
rect 8 8 20 14
rect 68 8 80 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m1p >>
rect -6 252 106 268
rect 3 123 17 137
rect 43 123 57 137
rect 83 123 97 137
rect 23 103 37 117
rect 63 103 77 117
rect -6 -8 106 8
<< labels >>
rlabel nsubstratencontact 51 260 51 260 0 vdd
port 6 nsew power bidirectional abutment
rlabel psubstratepcontact 51 0 51 0 0 gnd
port 7 nsew ground bidirectional abutment
rlabel metal1 10 128 10 128 0 A
port 1 nsew signal input
rlabel metal1 50 131 50 131 0 Y
port 5 nsew signal output
rlabel metal1 90 131 90 131 0 C
port 3 nsew signal input
rlabel metal1 30 110 30 110 0 B
port 2 nsew signal input
rlabel metal1 70 110 70 110 0 D
port 4 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 100 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
