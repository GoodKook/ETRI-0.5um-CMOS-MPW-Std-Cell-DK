magic
tech scmos
magscale 1 2
timestamp 0
<< metal1 >>
<< metal1 >>
rect 55 12 56 13
rect 54 12 55 13
rect 53 12 54 13
rect 52 12 53 13
rect 51 12 52 13
rect 50 12 51 13
rect 49 12 50 13
rect 48 12 49 13
rect 47 12 48 13
rect 46 12 47 13
rect 45 12 46 13
rect 44 12 45 13
rect 43 12 44 13
rect 42 12 43 13
rect 59 13 60 14
rect 58 13 59 14
rect 57 13 58 14
rect 56 13 57 14
rect 55 13 56 14
rect 54 13 55 14
rect 53 13 54 14
rect 52 13 53 14
rect 51 13 52 14
rect 50 13 51 14
rect 49 13 50 14
rect 48 13 49 14
rect 47 13 48 14
rect 46 13 47 14
rect 45 13 46 14
rect 44 13 45 14
rect 43 13 44 14
rect 42 13 43 14
rect 41 13 42 14
rect 40 13 41 14
rect 39 13 40 14
rect 38 13 39 14
rect 37 13 38 14
rect 62 14 63 15
rect 61 14 62 15
rect 60 14 61 15
rect 59 14 60 15
rect 58 14 59 15
rect 57 14 58 15
rect 56 14 57 15
rect 55 14 56 15
rect 54 14 55 15
rect 53 14 54 15
rect 52 14 53 15
rect 51 14 52 15
rect 50 14 51 15
rect 49 14 50 15
rect 48 14 49 15
rect 47 14 48 15
rect 46 14 47 15
rect 45 14 46 15
rect 44 14 45 15
rect 43 14 44 15
rect 42 14 43 15
rect 41 14 42 15
rect 40 14 41 15
rect 39 14 40 15
rect 38 14 39 15
rect 37 14 38 15
rect 36 14 37 15
rect 35 14 36 15
rect 34 14 35 15
rect 64 15 65 16
rect 63 15 64 16
rect 62 15 63 16
rect 61 15 62 16
rect 60 15 61 16
rect 59 15 60 16
rect 58 15 59 16
rect 57 15 58 16
rect 56 15 57 16
rect 55 15 56 16
rect 54 15 55 16
rect 53 15 54 16
rect 52 15 53 16
rect 51 15 52 16
rect 50 15 51 16
rect 49 15 50 16
rect 48 15 49 16
rect 47 15 48 16
rect 46 15 47 16
rect 45 15 46 16
rect 44 15 45 16
rect 43 15 44 16
rect 42 15 43 16
rect 41 15 42 16
rect 40 15 41 16
rect 39 15 40 16
rect 38 15 39 16
rect 37 15 38 16
rect 36 15 37 16
rect 35 15 36 16
rect 34 15 35 16
rect 33 15 34 16
rect 32 15 33 16
rect 66 16 67 17
rect 65 16 66 17
rect 64 16 65 17
rect 63 16 64 17
rect 62 16 63 17
rect 61 16 62 17
rect 60 16 61 17
rect 59 16 60 17
rect 58 16 59 17
rect 57 16 58 17
rect 56 16 57 17
rect 55 16 56 17
rect 54 16 55 17
rect 53 16 54 17
rect 52 16 53 17
rect 51 16 52 17
rect 50 16 51 17
rect 49 16 50 17
rect 48 16 49 17
rect 47 16 48 17
rect 46 16 47 17
rect 45 16 46 17
rect 44 16 45 17
rect 43 16 44 17
rect 42 16 43 17
rect 41 16 42 17
rect 40 16 41 17
rect 39 16 40 17
rect 38 16 39 17
rect 37 16 38 17
rect 36 16 37 17
rect 35 16 36 17
rect 34 16 35 17
rect 33 16 34 17
rect 32 16 33 17
rect 31 16 32 17
rect 30 16 31 17
rect 68 17 69 18
rect 67 17 68 18
rect 66 17 67 18
rect 65 17 66 18
rect 64 17 65 18
rect 63 17 64 18
rect 62 17 63 18
rect 61 17 62 18
rect 60 17 61 18
rect 59 17 60 18
rect 58 17 59 18
rect 57 17 58 18
rect 56 17 57 18
rect 55 17 56 18
rect 54 17 55 18
rect 53 17 54 18
rect 52 17 53 18
rect 51 17 52 18
rect 50 17 51 18
rect 49 17 50 18
rect 48 17 49 18
rect 47 17 48 18
rect 46 17 47 18
rect 45 17 46 18
rect 44 17 45 18
rect 43 17 44 18
rect 42 17 43 18
rect 41 17 42 18
rect 40 17 41 18
rect 39 17 40 18
rect 38 17 39 18
rect 37 17 38 18
rect 36 17 37 18
rect 35 17 36 18
rect 34 17 35 18
rect 33 17 34 18
rect 32 17 33 18
rect 31 17 32 18
rect 30 17 31 18
rect 29 17 30 18
rect 69 18 70 19
rect 68 18 69 19
rect 67 18 68 19
rect 66 18 67 19
rect 65 18 66 19
rect 64 18 65 19
rect 63 18 64 19
rect 62 18 63 19
rect 61 18 62 19
rect 60 18 61 19
rect 59 18 60 19
rect 58 18 59 19
rect 57 18 58 19
rect 56 18 57 19
rect 55 18 56 19
rect 54 18 55 19
rect 53 18 54 19
rect 52 18 53 19
rect 51 18 52 19
rect 50 18 51 19
rect 49 18 50 19
rect 48 18 49 19
rect 47 18 48 19
rect 46 18 47 19
rect 45 18 46 19
rect 44 18 45 19
rect 43 18 44 19
rect 42 18 43 19
rect 41 18 42 19
rect 40 18 41 19
rect 39 18 40 19
rect 38 18 39 19
rect 37 18 38 19
rect 36 18 37 19
rect 35 18 36 19
rect 34 18 35 19
rect 33 18 34 19
rect 32 18 33 19
rect 31 18 32 19
rect 30 18 31 19
rect 29 18 30 19
rect 28 18 29 19
rect 27 18 28 19
rect 70 19 71 20
rect 69 19 70 20
rect 68 19 69 20
rect 67 19 68 20
rect 66 19 67 20
rect 65 19 66 20
rect 64 19 65 20
rect 63 19 64 20
rect 62 19 63 20
rect 61 19 62 20
rect 60 19 61 20
rect 59 19 60 20
rect 58 19 59 20
rect 57 19 58 20
rect 56 19 57 20
rect 55 19 56 20
rect 54 19 55 20
rect 53 19 54 20
rect 52 19 53 20
rect 51 19 52 20
rect 50 19 51 20
rect 49 19 50 20
rect 48 19 49 20
rect 47 19 48 20
rect 46 19 47 20
rect 45 19 46 20
rect 44 19 45 20
rect 43 19 44 20
rect 42 19 43 20
rect 41 19 42 20
rect 40 19 41 20
rect 39 19 40 20
rect 38 19 39 20
rect 37 19 38 20
rect 36 19 37 20
rect 35 19 36 20
rect 34 19 35 20
rect 33 19 34 20
rect 32 19 33 20
rect 31 19 32 20
rect 30 19 31 20
rect 29 19 30 20
rect 28 19 29 20
rect 27 19 28 20
rect 26 19 27 20
rect 71 20 72 21
rect 70 20 71 21
rect 69 20 70 21
rect 68 20 69 21
rect 67 20 68 21
rect 66 20 67 21
rect 65 20 66 21
rect 64 20 65 21
rect 63 20 64 21
rect 62 20 63 21
rect 61 20 62 21
rect 60 20 61 21
rect 59 20 60 21
rect 58 20 59 21
rect 57 20 58 21
rect 56 20 57 21
rect 55 20 56 21
rect 54 20 55 21
rect 53 20 54 21
rect 52 20 53 21
rect 51 20 52 21
rect 50 20 51 21
rect 49 20 50 21
rect 48 20 49 21
rect 47 20 48 21
rect 46 20 47 21
rect 45 20 46 21
rect 44 20 45 21
rect 43 20 44 21
rect 42 20 43 21
rect 41 20 42 21
rect 40 20 41 21
rect 39 20 40 21
rect 38 20 39 21
rect 37 20 38 21
rect 36 20 37 21
rect 35 20 36 21
rect 34 20 35 21
rect 33 20 34 21
rect 32 20 33 21
rect 31 20 32 21
rect 30 20 31 21
rect 29 20 30 21
rect 28 20 29 21
rect 27 20 28 21
rect 26 20 27 21
rect 25 20 26 21
rect 72 21 73 22
rect 71 21 72 22
rect 70 21 71 22
rect 69 21 70 22
rect 68 21 69 22
rect 67 21 68 22
rect 66 21 67 22
rect 65 21 66 22
rect 64 21 65 22
rect 63 21 64 22
rect 62 21 63 22
rect 61 21 62 22
rect 60 21 61 22
rect 59 21 60 22
rect 58 21 59 22
rect 57 21 58 22
rect 56 21 57 22
rect 55 21 56 22
rect 54 21 55 22
rect 53 21 54 22
rect 52 21 53 22
rect 51 21 52 22
rect 50 21 51 22
rect 49 21 50 22
rect 48 21 49 22
rect 47 21 48 22
rect 46 21 47 22
rect 45 21 46 22
rect 44 21 45 22
rect 43 21 44 22
rect 42 21 43 22
rect 41 21 42 22
rect 40 21 41 22
rect 39 21 40 22
rect 38 21 39 22
rect 37 21 38 22
rect 36 21 37 22
rect 35 21 36 22
rect 34 21 35 22
rect 33 21 34 22
rect 32 21 33 22
rect 31 21 32 22
rect 30 21 31 22
rect 29 21 30 22
rect 28 21 29 22
rect 27 21 28 22
rect 26 21 27 22
rect 25 21 26 22
rect 24 21 25 22
rect 23 21 24 22
rect 73 22 74 23
rect 72 22 73 23
rect 71 22 72 23
rect 70 22 71 23
rect 69 22 70 23
rect 68 22 69 23
rect 67 22 68 23
rect 66 22 67 23
rect 65 22 66 23
rect 64 22 65 23
rect 63 22 64 23
rect 62 22 63 23
rect 61 22 62 23
rect 60 22 61 23
rect 59 22 60 23
rect 58 22 59 23
rect 57 22 58 23
rect 56 22 57 23
rect 55 22 56 23
rect 54 22 55 23
rect 53 22 54 23
rect 52 22 53 23
rect 51 22 52 23
rect 50 22 51 23
rect 49 22 50 23
rect 48 22 49 23
rect 47 22 48 23
rect 46 22 47 23
rect 45 22 46 23
rect 44 22 45 23
rect 43 22 44 23
rect 42 22 43 23
rect 41 22 42 23
rect 40 22 41 23
rect 39 22 40 23
rect 38 22 39 23
rect 37 22 38 23
rect 36 22 37 23
rect 35 22 36 23
rect 34 22 35 23
rect 33 22 34 23
rect 32 22 33 23
rect 31 22 32 23
rect 30 22 31 23
rect 29 22 30 23
rect 28 22 29 23
rect 27 22 28 23
rect 26 22 27 23
rect 25 22 26 23
rect 24 22 25 23
rect 23 22 24 23
rect 22 22 23 23
rect 74 23 75 24
rect 73 23 74 24
rect 72 23 73 24
rect 71 23 72 24
rect 70 23 71 24
rect 69 23 70 24
rect 68 23 69 24
rect 67 23 68 24
rect 66 23 67 24
rect 65 23 66 24
rect 64 23 65 24
rect 63 23 64 24
rect 62 23 63 24
rect 61 23 62 24
rect 60 23 61 24
rect 59 23 60 24
rect 58 23 59 24
rect 57 23 58 24
rect 56 23 57 24
rect 55 23 56 24
rect 54 23 55 24
rect 53 23 54 24
rect 52 23 53 24
rect 51 23 52 24
rect 50 23 51 24
rect 49 23 50 24
rect 48 23 49 24
rect 47 23 48 24
rect 46 23 47 24
rect 45 23 46 24
rect 44 23 45 24
rect 43 23 44 24
rect 42 23 43 24
rect 41 23 42 24
rect 40 23 41 24
rect 39 23 40 24
rect 38 23 39 24
rect 37 23 38 24
rect 36 23 37 24
rect 35 23 36 24
rect 34 23 35 24
rect 33 23 34 24
rect 32 23 33 24
rect 31 23 32 24
rect 30 23 31 24
rect 29 23 30 24
rect 28 23 29 24
rect 27 23 28 24
rect 26 23 27 24
rect 25 23 26 24
rect 24 23 25 24
rect 23 23 24 24
rect 22 23 23 24
rect 75 24 76 25
rect 74 24 75 25
rect 73 24 74 25
rect 72 24 73 25
rect 71 24 72 25
rect 70 24 71 25
rect 69 24 70 25
rect 68 24 69 25
rect 67 24 68 25
rect 66 24 67 25
rect 65 24 66 25
rect 64 24 65 25
rect 63 24 64 25
rect 62 24 63 25
rect 61 24 62 25
rect 60 24 61 25
rect 59 24 60 25
rect 58 24 59 25
rect 57 24 58 25
rect 56 24 57 25
rect 55 24 56 25
rect 54 24 55 25
rect 53 24 54 25
rect 52 24 53 25
rect 51 24 52 25
rect 50 24 51 25
rect 49 24 50 25
rect 48 24 49 25
rect 47 24 48 25
rect 46 24 47 25
rect 45 24 46 25
rect 44 24 45 25
rect 43 24 44 25
rect 42 24 43 25
rect 41 24 42 25
rect 40 24 41 25
rect 39 24 40 25
rect 38 24 39 25
rect 37 24 38 25
rect 36 24 37 25
rect 35 24 36 25
rect 34 24 35 25
rect 33 24 34 25
rect 32 24 33 25
rect 31 24 32 25
rect 30 24 31 25
rect 29 24 30 25
rect 28 24 29 25
rect 27 24 28 25
rect 26 24 27 25
rect 25 24 26 25
rect 24 24 25 25
rect 23 24 24 25
rect 22 24 23 25
rect 21 24 22 25
rect 76 25 77 26
rect 75 25 76 26
rect 74 25 75 26
rect 73 25 74 26
rect 72 25 73 26
rect 71 25 72 26
rect 70 25 71 26
rect 69 25 70 26
rect 68 25 69 26
rect 67 25 68 26
rect 66 25 67 26
rect 65 25 66 26
rect 64 25 65 26
rect 63 25 64 26
rect 62 25 63 26
rect 61 25 62 26
rect 60 25 61 26
rect 59 25 60 26
rect 58 25 59 26
rect 57 25 58 26
rect 56 25 57 26
rect 55 25 56 26
rect 54 25 55 26
rect 53 25 54 26
rect 52 25 53 26
rect 51 25 52 26
rect 50 25 51 26
rect 49 25 50 26
rect 48 25 49 26
rect 47 25 48 26
rect 46 25 47 26
rect 45 25 46 26
rect 44 25 45 26
rect 43 25 44 26
rect 42 25 43 26
rect 41 25 42 26
rect 40 25 41 26
rect 39 25 40 26
rect 38 25 39 26
rect 37 25 38 26
rect 36 25 37 26
rect 35 25 36 26
rect 34 25 35 26
rect 33 25 34 26
rect 32 25 33 26
rect 31 25 32 26
rect 30 25 31 26
rect 29 25 30 26
rect 28 25 29 26
rect 27 25 28 26
rect 26 25 27 26
rect 25 25 26 26
rect 24 25 25 26
rect 23 25 24 26
rect 22 25 23 26
rect 21 25 22 26
rect 20 25 21 26
rect 76 26 77 27
rect 75 26 76 27
rect 74 26 75 27
rect 73 26 74 27
rect 72 26 73 27
rect 71 26 72 27
rect 70 26 71 27
rect 69 26 70 27
rect 68 26 69 27
rect 67 26 68 27
rect 66 26 67 27
rect 65 26 66 27
rect 64 26 65 27
rect 63 26 64 27
rect 62 26 63 27
rect 61 26 62 27
rect 60 26 61 27
rect 59 26 60 27
rect 58 26 59 27
rect 57 26 58 27
rect 56 26 57 27
rect 55 26 56 27
rect 54 26 55 27
rect 53 26 54 27
rect 52 26 53 27
rect 51 26 52 27
rect 50 26 51 27
rect 49 26 50 27
rect 48 26 49 27
rect 47 26 48 27
rect 46 26 47 27
rect 45 26 46 27
rect 44 26 45 27
rect 43 26 44 27
rect 42 26 43 27
rect 41 26 42 27
rect 40 26 41 27
rect 39 26 40 27
rect 38 26 39 27
rect 37 26 38 27
rect 36 26 37 27
rect 35 26 36 27
rect 34 26 35 27
rect 33 26 34 27
rect 32 26 33 27
rect 31 26 32 27
rect 30 26 31 27
rect 29 26 30 27
rect 28 26 29 27
rect 27 26 28 27
rect 26 26 27 27
rect 25 26 26 27
rect 24 26 25 27
rect 23 26 24 27
rect 22 26 23 27
rect 21 26 22 27
rect 20 26 21 27
rect 19 26 20 27
rect 77 27 78 28
rect 76 27 77 28
rect 75 27 76 28
rect 74 27 75 28
rect 73 27 74 28
rect 72 27 73 28
rect 71 27 72 28
rect 70 27 71 28
rect 69 27 70 28
rect 68 27 69 28
rect 67 27 68 28
rect 66 27 67 28
rect 65 27 66 28
rect 64 27 65 28
rect 63 27 64 28
rect 62 27 63 28
rect 61 27 62 28
rect 60 27 61 28
rect 59 27 60 28
rect 58 27 59 28
rect 57 27 58 28
rect 56 27 57 28
rect 55 27 56 28
rect 54 27 55 28
rect 53 27 54 28
rect 52 27 53 28
rect 51 27 52 28
rect 50 27 51 28
rect 49 27 50 28
rect 48 27 49 28
rect 47 27 48 28
rect 46 27 47 28
rect 45 27 46 28
rect 44 27 45 28
rect 43 27 44 28
rect 42 27 43 28
rect 41 27 42 28
rect 40 27 41 28
rect 39 27 40 28
rect 38 27 39 28
rect 37 27 38 28
rect 36 27 37 28
rect 35 27 36 28
rect 34 27 35 28
rect 33 27 34 28
rect 32 27 33 28
rect 31 27 32 28
rect 30 27 31 28
rect 29 27 30 28
rect 28 27 29 28
rect 27 27 28 28
rect 26 27 27 28
rect 25 27 26 28
rect 24 27 25 28
rect 23 27 24 28
rect 22 27 23 28
rect 21 27 22 28
rect 20 27 21 28
rect 19 27 20 28
rect 77 28 78 29
rect 76 28 77 29
rect 75 28 76 29
rect 74 28 75 29
rect 73 28 74 29
rect 72 28 73 29
rect 71 28 72 29
rect 70 28 71 29
rect 69 28 70 29
rect 68 28 69 29
rect 67 28 68 29
rect 66 28 67 29
rect 65 28 66 29
rect 64 28 65 29
rect 63 28 64 29
rect 62 28 63 29
rect 61 28 62 29
rect 60 28 61 29
rect 59 28 60 29
rect 58 28 59 29
rect 57 28 58 29
rect 56 28 57 29
rect 55 28 56 29
rect 54 28 55 29
rect 53 28 54 29
rect 52 28 53 29
rect 51 28 52 29
rect 50 28 51 29
rect 49 28 50 29
rect 48 28 49 29
rect 47 28 48 29
rect 46 28 47 29
rect 45 28 46 29
rect 44 28 45 29
rect 43 28 44 29
rect 42 28 43 29
rect 41 28 42 29
rect 40 28 41 29
rect 39 28 40 29
rect 38 28 39 29
rect 37 28 38 29
rect 36 28 37 29
rect 35 28 36 29
rect 34 28 35 29
rect 33 28 34 29
rect 32 28 33 29
rect 31 28 32 29
rect 30 28 31 29
rect 29 28 30 29
rect 28 28 29 29
rect 27 28 28 29
rect 26 28 27 29
rect 25 28 26 29
rect 24 28 25 29
rect 23 28 24 29
rect 22 28 23 29
rect 21 28 22 29
rect 20 28 21 29
rect 19 28 20 29
rect 18 28 19 29
rect 78 29 79 30
rect 77 29 78 30
rect 76 29 77 30
rect 75 29 76 30
rect 74 29 75 30
rect 73 29 74 30
rect 72 29 73 30
rect 71 29 72 30
rect 70 29 71 30
rect 69 29 70 30
rect 68 29 69 30
rect 67 29 68 30
rect 66 29 67 30
rect 65 29 66 30
rect 64 29 65 30
rect 63 29 64 30
rect 62 29 63 30
rect 61 29 62 30
rect 60 29 61 30
rect 59 29 60 30
rect 58 29 59 30
rect 57 29 58 30
rect 56 29 57 30
rect 55 29 56 30
rect 54 29 55 30
rect 53 29 54 30
rect 52 29 53 30
rect 51 29 52 30
rect 50 29 51 30
rect 49 29 50 30
rect 48 29 49 30
rect 47 29 48 30
rect 46 29 47 30
rect 45 29 46 30
rect 44 29 45 30
rect 43 29 44 30
rect 42 29 43 30
rect 41 29 42 30
rect 40 29 41 30
rect 39 29 40 30
rect 38 29 39 30
rect 37 29 38 30
rect 36 29 37 30
rect 35 29 36 30
rect 34 29 35 30
rect 33 29 34 30
rect 32 29 33 30
rect 31 29 32 30
rect 30 29 31 30
rect 29 29 30 30
rect 28 29 29 30
rect 27 29 28 30
rect 26 29 27 30
rect 25 29 26 30
rect 24 29 25 30
rect 23 29 24 30
rect 22 29 23 30
rect 21 29 22 30
rect 20 29 21 30
rect 19 29 20 30
rect 18 29 19 30
rect 78 30 79 31
rect 77 30 78 31
rect 76 30 77 31
rect 75 30 76 31
rect 74 30 75 31
rect 73 30 74 31
rect 72 30 73 31
rect 71 30 72 31
rect 70 30 71 31
rect 69 30 70 31
rect 68 30 69 31
rect 67 30 68 31
rect 66 30 67 31
rect 65 30 66 31
rect 64 30 65 31
rect 63 30 64 31
rect 62 30 63 31
rect 61 30 62 31
rect 60 30 61 31
rect 59 30 60 31
rect 58 30 59 31
rect 57 30 58 31
rect 56 30 57 31
rect 55 30 56 31
rect 54 30 55 31
rect 53 30 54 31
rect 52 30 53 31
rect 51 30 52 31
rect 50 30 51 31
rect 49 30 50 31
rect 48 30 49 31
rect 47 30 48 31
rect 46 30 47 31
rect 45 30 46 31
rect 44 30 45 31
rect 43 30 44 31
rect 42 30 43 31
rect 41 30 42 31
rect 40 30 41 31
rect 39 30 40 31
rect 38 30 39 31
rect 37 30 38 31
rect 36 30 37 31
rect 35 30 36 31
rect 34 30 35 31
rect 33 30 34 31
rect 32 30 33 31
rect 31 30 32 31
rect 30 30 31 31
rect 29 30 30 31
rect 28 30 29 31
rect 27 30 28 31
rect 26 30 27 31
rect 25 30 26 31
rect 24 30 25 31
rect 23 30 24 31
rect 22 30 23 31
rect 21 30 22 31
rect 20 30 21 31
rect 19 30 20 31
rect 18 30 19 31
rect 17 30 18 31
rect 142 31 143 32
rect 141 31 142 32
rect 140 31 141 32
rect 139 31 140 32
rect 138 31 139 32
rect 137 31 138 32
rect 79 31 80 32
rect 78 31 79 32
rect 77 31 78 32
rect 76 31 77 32
rect 75 31 76 32
rect 74 31 75 32
rect 73 31 74 32
rect 72 31 73 32
rect 71 31 72 32
rect 70 31 71 32
rect 69 31 70 32
rect 68 31 69 32
rect 67 31 68 32
rect 66 31 67 32
rect 65 31 66 32
rect 64 31 65 32
rect 63 31 64 32
rect 62 31 63 32
rect 61 31 62 32
rect 60 31 61 32
rect 59 31 60 32
rect 58 31 59 32
rect 57 31 58 32
rect 56 31 57 32
rect 55 31 56 32
rect 54 31 55 32
rect 53 31 54 32
rect 52 31 53 32
rect 51 31 52 32
rect 50 31 51 32
rect 49 31 50 32
rect 48 31 49 32
rect 47 31 48 32
rect 46 31 47 32
rect 45 31 46 32
rect 44 31 45 32
rect 43 31 44 32
rect 42 31 43 32
rect 41 31 42 32
rect 40 31 41 32
rect 39 31 40 32
rect 38 31 39 32
rect 37 31 38 32
rect 36 31 37 32
rect 35 31 36 32
rect 34 31 35 32
rect 33 31 34 32
rect 32 31 33 32
rect 31 31 32 32
rect 30 31 31 32
rect 29 31 30 32
rect 28 31 29 32
rect 27 31 28 32
rect 26 31 27 32
rect 25 31 26 32
rect 24 31 25 32
rect 23 31 24 32
rect 22 31 23 32
rect 21 31 22 32
rect 20 31 21 32
rect 19 31 20 32
rect 18 31 19 32
rect 17 31 18 32
rect 142 32 143 33
rect 141 32 142 33
rect 140 32 141 33
rect 139 32 140 33
rect 138 32 139 33
rect 137 32 138 33
rect 136 32 137 33
rect 135 32 136 33
rect 122 32 123 33
rect 121 32 122 33
rect 120 32 121 33
rect 119 32 120 33
rect 79 32 80 33
rect 78 32 79 33
rect 77 32 78 33
rect 76 32 77 33
rect 75 32 76 33
rect 74 32 75 33
rect 73 32 74 33
rect 72 32 73 33
rect 71 32 72 33
rect 70 32 71 33
rect 69 32 70 33
rect 68 32 69 33
rect 67 32 68 33
rect 66 32 67 33
rect 65 32 66 33
rect 64 32 65 33
rect 63 32 64 33
rect 62 32 63 33
rect 61 32 62 33
rect 60 32 61 33
rect 59 32 60 33
rect 58 32 59 33
rect 57 32 58 33
rect 56 32 57 33
rect 55 32 56 33
rect 54 32 55 33
rect 53 32 54 33
rect 52 32 53 33
rect 51 32 52 33
rect 50 32 51 33
rect 49 32 50 33
rect 48 32 49 33
rect 47 32 48 33
rect 46 32 47 33
rect 45 32 46 33
rect 44 32 45 33
rect 43 32 44 33
rect 42 32 43 33
rect 41 32 42 33
rect 40 32 41 33
rect 39 32 40 33
rect 38 32 39 33
rect 37 32 38 33
rect 36 32 37 33
rect 35 32 36 33
rect 34 32 35 33
rect 33 32 34 33
rect 32 32 33 33
rect 31 32 32 33
rect 30 32 31 33
rect 29 32 30 33
rect 28 32 29 33
rect 27 32 28 33
rect 26 32 27 33
rect 25 32 26 33
rect 24 32 25 33
rect 23 32 24 33
rect 22 32 23 33
rect 21 32 22 33
rect 20 32 21 33
rect 19 32 20 33
rect 18 32 19 33
rect 17 32 18 33
rect 16 32 17 33
rect 142 33 143 34
rect 141 33 142 34
rect 140 33 141 34
rect 139 33 140 34
rect 138 33 139 34
rect 137 33 138 34
rect 136 33 137 34
rect 135 33 136 34
rect 134 33 135 34
rect 122 33 123 34
rect 121 33 122 34
rect 120 33 121 34
rect 119 33 120 34
rect 118 33 119 34
rect 79 33 80 34
rect 78 33 79 34
rect 77 33 78 34
rect 76 33 77 34
rect 75 33 76 34
rect 74 33 75 34
rect 73 33 74 34
rect 72 33 73 34
rect 71 33 72 34
rect 70 33 71 34
rect 69 33 70 34
rect 68 33 69 34
rect 67 33 68 34
rect 66 33 67 34
rect 65 33 66 34
rect 64 33 65 34
rect 63 33 64 34
rect 62 33 63 34
rect 61 33 62 34
rect 60 33 61 34
rect 59 33 60 34
rect 58 33 59 34
rect 57 33 58 34
rect 56 33 57 34
rect 55 33 56 34
rect 54 33 55 34
rect 53 33 54 34
rect 52 33 53 34
rect 51 33 52 34
rect 43 33 44 34
rect 42 33 43 34
rect 41 33 42 34
rect 40 33 41 34
rect 39 33 40 34
rect 38 33 39 34
rect 37 33 38 34
rect 36 33 37 34
rect 35 33 36 34
rect 34 33 35 34
rect 33 33 34 34
rect 32 33 33 34
rect 31 33 32 34
rect 30 33 31 34
rect 29 33 30 34
rect 28 33 29 34
rect 27 33 28 34
rect 26 33 27 34
rect 25 33 26 34
rect 24 33 25 34
rect 23 33 24 34
rect 22 33 23 34
rect 21 33 22 34
rect 20 33 21 34
rect 19 33 20 34
rect 18 33 19 34
rect 17 33 18 34
rect 16 33 17 34
rect 142 34 143 35
rect 141 34 142 35
rect 140 34 141 35
rect 139 34 140 35
rect 138 34 139 35
rect 137 34 138 35
rect 136 34 137 35
rect 135 34 136 35
rect 134 34 135 35
rect 133 34 134 35
rect 121 34 122 35
rect 120 34 121 35
rect 119 34 120 35
rect 118 34 119 35
rect 79 34 80 35
rect 78 34 79 35
rect 77 34 78 35
rect 76 34 77 35
rect 75 34 76 35
rect 74 34 75 35
rect 73 34 74 35
rect 72 34 73 35
rect 71 34 72 35
rect 70 34 71 35
rect 69 34 70 35
rect 68 34 69 35
rect 67 34 68 35
rect 66 34 67 35
rect 65 34 66 35
rect 64 34 65 35
rect 63 34 64 35
rect 62 34 63 35
rect 61 34 62 35
rect 60 34 61 35
rect 59 34 60 35
rect 58 34 59 35
rect 57 34 58 35
rect 56 34 57 35
rect 55 34 56 35
rect 39 34 40 35
rect 38 34 39 35
rect 37 34 38 35
rect 36 34 37 35
rect 35 34 36 35
rect 34 34 35 35
rect 33 34 34 35
rect 32 34 33 35
rect 31 34 32 35
rect 30 34 31 35
rect 29 34 30 35
rect 28 34 29 35
rect 27 34 28 35
rect 26 34 27 35
rect 25 34 26 35
rect 24 34 25 35
rect 23 34 24 35
rect 22 34 23 35
rect 21 34 22 35
rect 20 34 21 35
rect 19 34 20 35
rect 18 34 19 35
rect 17 34 18 35
rect 16 34 17 35
rect 15 34 16 35
rect 142 35 143 36
rect 141 35 142 36
rect 140 35 141 36
rect 139 35 140 36
rect 138 35 139 36
rect 137 35 138 36
rect 136 35 137 36
rect 135 35 136 36
rect 134 35 135 36
rect 133 35 134 36
rect 132 35 133 36
rect 121 35 122 36
rect 120 35 121 36
rect 119 35 120 36
rect 118 35 119 36
rect 80 35 81 36
rect 79 35 80 36
rect 78 35 79 36
rect 77 35 78 36
rect 76 35 77 36
rect 75 35 76 36
rect 74 35 75 36
rect 73 35 74 36
rect 72 35 73 36
rect 71 35 72 36
rect 70 35 71 36
rect 69 35 70 36
rect 68 35 69 36
rect 67 35 68 36
rect 66 35 67 36
rect 65 35 66 36
rect 64 35 65 36
rect 63 35 64 36
rect 62 35 63 36
rect 61 35 62 36
rect 60 35 61 36
rect 59 35 60 36
rect 58 35 59 36
rect 57 35 58 36
rect 37 35 38 36
rect 36 35 37 36
rect 35 35 36 36
rect 34 35 35 36
rect 33 35 34 36
rect 32 35 33 36
rect 31 35 32 36
rect 30 35 31 36
rect 29 35 30 36
rect 28 35 29 36
rect 27 35 28 36
rect 26 35 27 36
rect 25 35 26 36
rect 24 35 25 36
rect 23 35 24 36
rect 22 35 23 36
rect 21 35 22 36
rect 20 35 21 36
rect 19 35 20 36
rect 18 35 19 36
rect 17 35 18 36
rect 16 35 17 36
rect 15 35 16 36
rect 142 36 143 37
rect 141 36 142 37
rect 140 36 141 37
rect 139 36 140 37
rect 138 36 139 37
rect 137 36 138 37
rect 136 36 137 37
rect 135 36 136 37
rect 134 36 135 37
rect 133 36 134 37
rect 132 36 133 37
rect 121 36 122 37
rect 120 36 121 37
rect 119 36 120 37
rect 118 36 119 37
rect 117 36 118 37
rect 80 36 81 37
rect 79 36 80 37
rect 78 36 79 37
rect 77 36 78 37
rect 76 36 77 37
rect 75 36 76 37
rect 74 36 75 37
rect 73 36 74 37
rect 72 36 73 37
rect 71 36 72 37
rect 70 36 71 37
rect 69 36 70 37
rect 68 36 69 37
rect 67 36 68 37
rect 66 36 67 37
rect 65 36 66 37
rect 64 36 65 37
rect 63 36 64 37
rect 62 36 63 37
rect 61 36 62 37
rect 60 36 61 37
rect 59 36 60 37
rect 58 36 59 37
rect 36 36 37 37
rect 35 36 36 37
rect 34 36 35 37
rect 33 36 34 37
rect 32 36 33 37
rect 31 36 32 37
rect 30 36 31 37
rect 29 36 30 37
rect 28 36 29 37
rect 27 36 28 37
rect 26 36 27 37
rect 25 36 26 37
rect 24 36 25 37
rect 23 36 24 37
rect 22 36 23 37
rect 21 36 22 37
rect 20 36 21 37
rect 19 36 20 37
rect 18 36 19 37
rect 17 36 18 37
rect 16 36 17 37
rect 15 36 16 37
rect 142 37 143 38
rect 141 37 142 38
rect 140 37 141 38
rect 139 37 140 38
rect 138 37 139 38
rect 136 37 137 38
rect 135 37 136 38
rect 134 37 135 38
rect 133 37 134 38
rect 132 37 133 38
rect 131 37 132 38
rect 120 37 121 38
rect 119 37 120 38
rect 118 37 119 38
rect 117 37 118 38
rect 80 37 81 38
rect 79 37 80 38
rect 78 37 79 38
rect 77 37 78 38
rect 76 37 77 38
rect 75 37 76 38
rect 74 37 75 38
rect 73 37 74 38
rect 72 37 73 38
rect 71 37 72 38
rect 70 37 71 38
rect 69 37 70 38
rect 68 37 69 38
rect 67 37 68 38
rect 66 37 67 38
rect 65 37 66 38
rect 64 37 65 38
rect 63 37 64 38
rect 62 37 63 38
rect 61 37 62 38
rect 60 37 61 38
rect 34 37 35 38
rect 33 37 34 38
rect 32 37 33 38
rect 31 37 32 38
rect 30 37 31 38
rect 29 37 30 38
rect 28 37 29 38
rect 27 37 28 38
rect 26 37 27 38
rect 25 37 26 38
rect 24 37 25 38
rect 23 37 24 38
rect 22 37 23 38
rect 21 37 22 38
rect 20 37 21 38
rect 19 37 20 38
rect 18 37 19 38
rect 17 37 18 38
rect 16 37 17 38
rect 15 37 16 38
rect 14 37 15 38
rect 142 38 143 39
rect 141 38 142 39
rect 140 38 141 39
rect 139 38 140 39
rect 138 38 139 39
rect 135 38 136 39
rect 134 38 135 39
rect 133 38 134 39
rect 132 38 133 39
rect 131 38 132 39
rect 130 38 131 39
rect 120 38 121 39
rect 119 38 120 39
rect 118 38 119 39
rect 117 38 118 39
rect 80 38 81 39
rect 79 38 80 39
rect 78 38 79 39
rect 77 38 78 39
rect 76 38 77 39
rect 75 38 76 39
rect 74 38 75 39
rect 73 38 74 39
rect 72 38 73 39
rect 71 38 72 39
rect 70 38 71 39
rect 69 38 70 39
rect 68 38 69 39
rect 67 38 68 39
rect 66 38 67 39
rect 65 38 66 39
rect 64 38 65 39
rect 63 38 64 39
rect 62 38 63 39
rect 61 38 62 39
rect 33 38 34 39
rect 32 38 33 39
rect 31 38 32 39
rect 30 38 31 39
rect 29 38 30 39
rect 28 38 29 39
rect 27 38 28 39
rect 26 38 27 39
rect 25 38 26 39
rect 24 38 25 39
rect 23 38 24 39
rect 22 38 23 39
rect 21 38 22 39
rect 20 38 21 39
rect 19 38 20 39
rect 18 38 19 39
rect 17 38 18 39
rect 16 38 17 39
rect 15 38 16 39
rect 14 38 15 39
rect 142 39 143 40
rect 141 39 142 40
rect 140 39 141 40
rect 139 39 140 40
rect 138 39 139 40
rect 134 39 135 40
rect 133 39 134 40
rect 132 39 133 40
rect 131 39 132 40
rect 130 39 131 40
rect 129 39 130 40
rect 121 39 122 40
rect 120 39 121 40
rect 119 39 120 40
rect 118 39 119 40
rect 117 39 118 40
rect 80 39 81 40
rect 79 39 80 40
rect 78 39 79 40
rect 77 39 78 40
rect 76 39 77 40
rect 75 39 76 40
rect 74 39 75 40
rect 73 39 74 40
rect 72 39 73 40
rect 71 39 72 40
rect 70 39 71 40
rect 69 39 70 40
rect 68 39 69 40
rect 67 39 68 40
rect 66 39 67 40
rect 65 39 66 40
rect 64 39 65 40
rect 63 39 64 40
rect 62 39 63 40
rect 32 39 33 40
rect 31 39 32 40
rect 30 39 31 40
rect 29 39 30 40
rect 28 39 29 40
rect 27 39 28 40
rect 26 39 27 40
rect 25 39 26 40
rect 24 39 25 40
rect 23 39 24 40
rect 22 39 23 40
rect 21 39 22 40
rect 20 39 21 40
rect 19 39 20 40
rect 18 39 19 40
rect 17 39 18 40
rect 16 39 17 40
rect 15 39 16 40
rect 14 39 15 40
rect 142 40 143 41
rect 141 40 142 41
rect 140 40 141 41
rect 139 40 140 41
rect 138 40 139 41
rect 133 40 134 41
rect 132 40 133 41
rect 131 40 132 41
rect 130 40 131 41
rect 129 40 130 41
rect 128 40 129 41
rect 121 40 122 41
rect 120 40 121 41
rect 119 40 120 41
rect 118 40 119 41
rect 117 40 118 41
rect 81 40 82 41
rect 80 40 81 41
rect 79 40 80 41
rect 78 40 79 41
rect 77 40 78 41
rect 76 40 77 41
rect 75 40 76 41
rect 74 40 75 41
rect 73 40 74 41
rect 72 40 73 41
rect 71 40 72 41
rect 70 40 71 41
rect 69 40 70 41
rect 68 40 69 41
rect 67 40 68 41
rect 66 40 67 41
rect 65 40 66 41
rect 64 40 65 41
rect 63 40 64 41
rect 62 40 63 41
rect 32 40 33 41
rect 31 40 32 41
rect 30 40 31 41
rect 29 40 30 41
rect 28 40 29 41
rect 27 40 28 41
rect 26 40 27 41
rect 25 40 26 41
rect 24 40 25 41
rect 23 40 24 41
rect 22 40 23 41
rect 21 40 22 41
rect 20 40 21 41
rect 19 40 20 41
rect 18 40 19 41
rect 17 40 18 41
rect 16 40 17 41
rect 15 40 16 41
rect 14 40 15 41
rect 142 41 143 42
rect 141 41 142 42
rect 140 41 141 42
rect 139 41 140 42
rect 138 41 139 42
rect 133 41 134 42
rect 132 41 133 42
rect 131 41 132 42
rect 130 41 131 42
rect 129 41 130 42
rect 128 41 129 42
rect 127 41 128 42
rect 122 41 123 42
rect 121 41 122 42
rect 120 41 121 42
rect 119 41 120 42
rect 118 41 119 42
rect 117 41 118 42
rect 81 41 82 42
rect 80 41 81 42
rect 79 41 80 42
rect 78 41 79 42
rect 77 41 78 42
rect 76 41 77 42
rect 75 41 76 42
rect 74 41 75 42
rect 73 41 74 42
rect 72 41 73 42
rect 71 41 72 42
rect 70 41 71 42
rect 69 41 70 42
rect 68 41 69 42
rect 67 41 68 42
rect 66 41 67 42
rect 65 41 66 42
rect 64 41 65 42
rect 63 41 64 42
rect 31 41 32 42
rect 30 41 31 42
rect 29 41 30 42
rect 28 41 29 42
rect 27 41 28 42
rect 26 41 27 42
rect 25 41 26 42
rect 24 41 25 42
rect 23 41 24 42
rect 22 41 23 42
rect 21 41 22 42
rect 20 41 21 42
rect 19 41 20 42
rect 18 41 19 42
rect 17 41 18 42
rect 16 41 17 42
rect 15 41 16 42
rect 14 41 15 42
rect 142 42 143 43
rect 141 42 142 43
rect 140 42 141 43
rect 139 42 140 43
rect 138 42 139 43
rect 132 42 133 43
rect 131 42 132 43
rect 130 42 131 43
rect 129 42 130 43
rect 128 42 129 43
rect 127 42 128 43
rect 126 42 127 43
rect 125 42 126 43
rect 124 42 125 43
rect 123 42 124 43
rect 122 42 123 43
rect 121 42 122 43
rect 120 42 121 43
rect 119 42 120 43
rect 118 42 119 43
rect 117 42 118 43
rect 81 42 82 43
rect 80 42 81 43
rect 79 42 80 43
rect 78 42 79 43
rect 77 42 78 43
rect 76 42 77 43
rect 75 42 76 43
rect 74 42 75 43
rect 73 42 74 43
rect 72 42 73 43
rect 71 42 72 43
rect 70 42 71 43
rect 69 42 70 43
rect 68 42 69 43
rect 67 42 68 43
rect 66 42 67 43
rect 65 42 66 43
rect 64 42 65 43
rect 63 42 64 43
rect 31 42 32 43
rect 30 42 31 43
rect 29 42 30 43
rect 28 42 29 43
rect 27 42 28 43
rect 26 42 27 43
rect 25 42 26 43
rect 24 42 25 43
rect 23 42 24 43
rect 22 42 23 43
rect 21 42 22 43
rect 20 42 21 43
rect 19 42 20 43
rect 18 42 19 43
rect 17 42 18 43
rect 16 42 17 43
rect 15 42 16 43
rect 14 42 15 43
rect 13 42 14 43
rect 142 43 143 44
rect 141 43 142 44
rect 140 43 141 44
rect 139 43 140 44
rect 138 43 139 44
rect 131 43 132 44
rect 130 43 131 44
rect 129 43 130 44
rect 128 43 129 44
rect 127 43 128 44
rect 126 43 127 44
rect 125 43 126 44
rect 124 43 125 44
rect 123 43 124 44
rect 122 43 123 44
rect 121 43 122 44
rect 120 43 121 44
rect 119 43 120 44
rect 118 43 119 44
rect 81 43 82 44
rect 80 43 81 44
rect 79 43 80 44
rect 78 43 79 44
rect 77 43 78 44
rect 76 43 77 44
rect 75 43 76 44
rect 74 43 75 44
rect 73 43 74 44
rect 72 43 73 44
rect 71 43 72 44
rect 70 43 71 44
rect 69 43 70 44
rect 68 43 69 44
rect 67 43 68 44
rect 66 43 67 44
rect 65 43 66 44
rect 64 43 65 44
rect 30 43 31 44
rect 29 43 30 44
rect 28 43 29 44
rect 27 43 28 44
rect 26 43 27 44
rect 25 43 26 44
rect 24 43 25 44
rect 23 43 24 44
rect 22 43 23 44
rect 21 43 22 44
rect 20 43 21 44
rect 19 43 20 44
rect 18 43 19 44
rect 17 43 18 44
rect 16 43 17 44
rect 15 43 16 44
rect 14 43 15 44
rect 13 43 14 44
rect 142 44 143 45
rect 141 44 142 45
rect 140 44 141 45
rect 139 44 140 45
rect 138 44 139 45
rect 130 44 131 45
rect 129 44 130 45
rect 128 44 129 45
rect 127 44 128 45
rect 126 44 127 45
rect 125 44 126 45
rect 124 44 125 45
rect 123 44 124 45
rect 122 44 123 45
rect 121 44 122 45
rect 120 44 121 45
rect 119 44 120 45
rect 118 44 119 45
rect 81 44 82 45
rect 80 44 81 45
rect 79 44 80 45
rect 78 44 79 45
rect 77 44 78 45
rect 76 44 77 45
rect 75 44 76 45
rect 74 44 75 45
rect 73 44 74 45
rect 72 44 73 45
rect 71 44 72 45
rect 70 44 71 45
rect 69 44 70 45
rect 68 44 69 45
rect 67 44 68 45
rect 66 44 67 45
rect 65 44 66 45
rect 64 44 65 45
rect 30 44 31 45
rect 29 44 30 45
rect 28 44 29 45
rect 27 44 28 45
rect 26 44 27 45
rect 25 44 26 45
rect 24 44 25 45
rect 23 44 24 45
rect 22 44 23 45
rect 21 44 22 45
rect 20 44 21 45
rect 19 44 20 45
rect 18 44 19 45
rect 17 44 18 45
rect 16 44 17 45
rect 15 44 16 45
rect 14 44 15 45
rect 13 44 14 45
rect 142 45 143 46
rect 141 45 142 46
rect 140 45 141 46
rect 139 45 140 46
rect 138 45 139 46
rect 129 45 130 46
rect 128 45 129 46
rect 127 45 128 46
rect 126 45 127 46
rect 125 45 126 46
rect 124 45 125 46
rect 123 45 124 46
rect 122 45 123 46
rect 121 45 122 46
rect 120 45 121 46
rect 119 45 120 46
rect 81 45 82 46
rect 80 45 81 46
rect 79 45 80 46
rect 78 45 79 46
rect 77 45 78 46
rect 76 45 77 46
rect 75 45 76 46
rect 74 45 75 46
rect 73 45 74 46
rect 72 45 73 46
rect 71 45 72 46
rect 70 45 71 46
rect 69 45 70 46
rect 68 45 69 46
rect 67 45 68 46
rect 66 45 67 46
rect 65 45 66 46
rect 64 45 65 46
rect 30 45 31 46
rect 29 45 30 46
rect 28 45 29 46
rect 27 45 28 46
rect 26 45 27 46
rect 25 45 26 46
rect 24 45 25 46
rect 23 45 24 46
rect 22 45 23 46
rect 21 45 22 46
rect 20 45 21 46
rect 19 45 20 46
rect 18 45 19 46
rect 17 45 18 46
rect 16 45 17 46
rect 15 45 16 46
rect 14 45 15 46
rect 13 45 14 46
rect 142 46 143 47
rect 141 46 142 47
rect 140 46 141 47
rect 139 46 140 47
rect 138 46 139 47
rect 128 46 129 47
rect 127 46 128 47
rect 126 46 127 47
rect 125 46 126 47
rect 124 46 125 47
rect 123 46 124 47
rect 122 46 123 47
rect 121 46 122 47
rect 120 46 121 47
rect 81 46 82 47
rect 80 46 81 47
rect 79 46 80 47
rect 78 46 79 47
rect 77 46 78 47
rect 76 46 77 47
rect 75 46 76 47
rect 74 46 75 47
rect 73 46 74 47
rect 72 46 73 47
rect 71 46 72 47
rect 70 46 71 47
rect 69 46 70 47
rect 68 46 69 47
rect 67 46 68 47
rect 66 46 67 47
rect 65 46 66 47
rect 29 46 30 47
rect 28 46 29 47
rect 27 46 28 47
rect 26 46 27 47
rect 25 46 26 47
rect 24 46 25 47
rect 23 46 24 47
rect 22 46 23 47
rect 21 46 22 47
rect 20 46 21 47
rect 19 46 20 47
rect 18 46 19 47
rect 17 46 18 47
rect 16 46 17 47
rect 15 46 16 47
rect 14 46 15 47
rect 13 46 14 47
rect 142 47 143 48
rect 141 47 142 48
rect 140 47 141 48
rect 139 47 140 48
rect 138 47 139 48
rect 125 47 126 48
rect 124 47 125 48
rect 123 47 124 48
rect 81 47 82 48
rect 80 47 81 48
rect 79 47 80 48
rect 78 47 79 48
rect 77 47 78 48
rect 76 47 77 48
rect 75 47 76 48
rect 74 47 75 48
rect 73 47 74 48
rect 72 47 73 48
rect 71 47 72 48
rect 70 47 71 48
rect 69 47 70 48
rect 68 47 69 48
rect 67 47 68 48
rect 66 47 67 48
rect 65 47 66 48
rect 29 47 30 48
rect 28 47 29 48
rect 27 47 28 48
rect 26 47 27 48
rect 25 47 26 48
rect 24 47 25 48
rect 23 47 24 48
rect 22 47 23 48
rect 21 47 22 48
rect 20 47 21 48
rect 19 47 20 48
rect 18 47 19 48
rect 17 47 18 48
rect 16 47 17 48
rect 15 47 16 48
rect 14 47 15 48
rect 13 47 14 48
rect 81 48 82 49
rect 80 48 81 49
rect 79 48 80 49
rect 78 48 79 49
rect 77 48 78 49
rect 76 48 77 49
rect 75 48 76 49
rect 74 48 75 49
rect 73 48 74 49
rect 72 48 73 49
rect 71 48 72 49
rect 70 48 71 49
rect 69 48 70 49
rect 68 48 69 49
rect 67 48 68 49
rect 66 48 67 49
rect 65 48 66 49
rect 29 48 30 49
rect 28 48 29 49
rect 27 48 28 49
rect 26 48 27 49
rect 25 48 26 49
rect 24 48 25 49
rect 23 48 24 49
rect 22 48 23 49
rect 21 48 22 49
rect 20 48 21 49
rect 19 48 20 49
rect 18 48 19 49
rect 17 48 18 49
rect 16 48 17 49
rect 15 48 16 49
rect 14 48 15 49
rect 13 48 14 49
rect 81 49 82 50
rect 80 49 81 50
rect 79 49 80 50
rect 78 49 79 50
rect 77 49 78 50
rect 76 49 77 50
rect 75 49 76 50
rect 74 49 75 50
rect 73 49 74 50
rect 72 49 73 50
rect 71 49 72 50
rect 70 49 71 50
rect 69 49 70 50
rect 68 49 69 50
rect 67 49 68 50
rect 66 49 67 50
rect 65 49 66 50
rect 29 49 30 50
rect 28 49 29 50
rect 27 49 28 50
rect 26 49 27 50
rect 25 49 26 50
rect 24 49 25 50
rect 23 49 24 50
rect 22 49 23 50
rect 21 49 22 50
rect 20 49 21 50
rect 19 49 20 50
rect 18 49 19 50
rect 17 49 18 50
rect 16 49 17 50
rect 15 49 16 50
rect 14 49 15 50
rect 13 49 14 50
rect 81 50 82 51
rect 80 50 81 51
rect 79 50 80 51
rect 78 50 79 51
rect 77 50 78 51
rect 76 50 77 51
rect 75 50 76 51
rect 74 50 75 51
rect 73 50 74 51
rect 72 50 73 51
rect 71 50 72 51
rect 70 50 71 51
rect 69 50 70 51
rect 68 50 69 51
rect 67 50 68 51
rect 66 50 67 51
rect 65 50 66 51
rect 29 50 30 51
rect 28 50 29 51
rect 27 50 28 51
rect 26 50 27 51
rect 25 50 26 51
rect 24 50 25 51
rect 23 50 24 51
rect 22 50 23 51
rect 21 50 22 51
rect 20 50 21 51
rect 19 50 20 51
rect 18 50 19 51
rect 17 50 18 51
rect 16 50 17 51
rect 15 50 16 51
rect 14 50 15 51
rect 13 50 14 51
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 78 51 79 52
rect 77 51 78 52
rect 76 51 77 52
rect 75 51 76 52
rect 74 51 75 52
rect 73 51 74 52
rect 72 51 73 52
rect 71 51 72 52
rect 70 51 71 52
rect 69 51 70 52
rect 68 51 69 52
rect 67 51 68 52
rect 66 51 67 52
rect 65 51 66 52
rect 29 51 30 52
rect 28 51 29 52
rect 27 51 28 52
rect 26 51 27 52
rect 25 51 26 52
rect 24 51 25 52
rect 23 51 24 52
rect 22 51 23 52
rect 21 51 22 52
rect 20 51 21 52
rect 19 51 20 52
rect 18 51 19 52
rect 17 51 18 52
rect 16 51 17 52
rect 15 51 16 52
rect 14 51 15 52
rect 13 51 14 52
rect 135 52 136 53
rect 134 52 135 53
rect 133 52 134 53
rect 132 52 133 53
rect 131 52 132 53
rect 130 52 131 53
rect 129 52 130 53
rect 128 52 129 53
rect 127 52 128 53
rect 126 52 127 53
rect 125 52 126 53
rect 124 52 125 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 77 52 78 53
rect 76 52 77 53
rect 75 52 76 53
rect 74 52 75 53
rect 73 52 74 53
rect 72 52 73 53
rect 71 52 72 53
rect 70 52 71 53
rect 69 52 70 53
rect 68 52 69 53
rect 67 52 68 53
rect 66 52 67 53
rect 65 52 66 53
rect 29 52 30 53
rect 28 52 29 53
rect 27 52 28 53
rect 26 52 27 53
rect 25 52 26 53
rect 24 52 25 53
rect 23 52 24 53
rect 22 52 23 53
rect 21 52 22 53
rect 20 52 21 53
rect 19 52 20 53
rect 18 52 19 53
rect 17 52 18 53
rect 16 52 17 53
rect 15 52 16 53
rect 14 52 15 53
rect 13 52 14 53
rect 138 53 139 54
rect 137 53 138 54
rect 136 53 137 54
rect 135 53 136 54
rect 134 53 135 54
rect 133 53 134 54
rect 132 53 133 54
rect 131 53 132 54
rect 130 53 131 54
rect 129 53 130 54
rect 128 53 129 54
rect 127 53 128 54
rect 126 53 127 54
rect 125 53 126 54
rect 124 53 125 54
rect 123 53 124 54
rect 122 53 123 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 76 53 77 54
rect 75 53 76 54
rect 74 53 75 54
rect 73 53 74 54
rect 72 53 73 54
rect 71 53 72 54
rect 70 53 71 54
rect 69 53 70 54
rect 68 53 69 54
rect 67 53 68 54
rect 66 53 67 54
rect 65 53 66 54
rect 29 53 30 54
rect 28 53 29 54
rect 27 53 28 54
rect 26 53 27 54
rect 25 53 26 54
rect 24 53 25 54
rect 23 53 24 54
rect 22 53 23 54
rect 21 53 22 54
rect 20 53 21 54
rect 19 53 20 54
rect 18 53 19 54
rect 17 53 18 54
rect 16 53 17 54
rect 15 53 16 54
rect 14 53 15 54
rect 13 53 14 54
rect 139 54 140 55
rect 138 54 139 55
rect 137 54 138 55
rect 136 54 137 55
rect 135 54 136 55
rect 134 54 135 55
rect 133 54 134 55
rect 132 54 133 55
rect 131 54 132 55
rect 130 54 131 55
rect 129 54 130 55
rect 128 54 129 55
rect 127 54 128 55
rect 126 54 127 55
rect 125 54 126 55
rect 124 54 125 55
rect 123 54 124 55
rect 122 54 123 55
rect 121 54 122 55
rect 120 54 121 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 75 54 76 55
rect 74 54 75 55
rect 73 54 74 55
rect 72 54 73 55
rect 71 54 72 55
rect 70 54 71 55
rect 69 54 70 55
rect 68 54 69 55
rect 67 54 68 55
rect 66 54 67 55
rect 65 54 66 55
rect 29 54 30 55
rect 28 54 29 55
rect 27 54 28 55
rect 26 54 27 55
rect 25 54 26 55
rect 24 54 25 55
rect 23 54 24 55
rect 22 54 23 55
rect 21 54 22 55
rect 20 54 21 55
rect 19 54 20 55
rect 18 54 19 55
rect 17 54 18 55
rect 16 54 17 55
rect 15 54 16 55
rect 14 54 15 55
rect 13 54 14 55
rect 140 55 141 56
rect 139 55 140 56
rect 138 55 139 56
rect 137 55 138 56
rect 136 55 137 56
rect 135 55 136 56
rect 134 55 135 56
rect 133 55 134 56
rect 132 55 133 56
rect 131 55 132 56
rect 130 55 131 56
rect 129 55 130 56
rect 128 55 129 56
rect 127 55 128 56
rect 126 55 127 56
rect 125 55 126 56
rect 124 55 125 56
rect 123 55 124 56
rect 122 55 123 56
rect 121 55 122 56
rect 120 55 121 56
rect 119 55 120 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 75 55 76 56
rect 74 55 75 56
rect 73 55 74 56
rect 72 55 73 56
rect 71 55 72 56
rect 70 55 71 56
rect 69 55 70 56
rect 68 55 69 56
rect 67 55 68 56
rect 66 55 67 56
rect 65 55 66 56
rect 29 55 30 56
rect 28 55 29 56
rect 27 55 28 56
rect 26 55 27 56
rect 25 55 26 56
rect 24 55 25 56
rect 23 55 24 56
rect 22 55 23 56
rect 21 55 22 56
rect 20 55 21 56
rect 19 55 20 56
rect 18 55 19 56
rect 17 55 18 56
rect 16 55 17 56
rect 15 55 16 56
rect 14 55 15 56
rect 13 55 14 56
rect 141 56 142 57
rect 140 56 141 57
rect 139 56 140 57
rect 138 56 139 57
rect 137 56 138 57
rect 136 56 137 57
rect 135 56 136 57
rect 134 56 135 57
rect 133 56 134 57
rect 132 56 133 57
rect 131 56 132 57
rect 130 56 131 57
rect 129 56 130 57
rect 128 56 129 57
rect 127 56 128 57
rect 126 56 127 57
rect 125 56 126 57
rect 124 56 125 57
rect 123 56 124 57
rect 122 56 123 57
rect 121 56 122 57
rect 120 56 121 57
rect 119 56 120 57
rect 118 56 119 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 74 56 75 57
rect 73 56 74 57
rect 72 56 73 57
rect 71 56 72 57
rect 70 56 71 57
rect 69 56 70 57
rect 68 56 69 57
rect 67 56 68 57
rect 66 56 67 57
rect 65 56 66 57
rect 64 56 65 57
rect 29 56 30 57
rect 28 56 29 57
rect 27 56 28 57
rect 26 56 27 57
rect 25 56 26 57
rect 24 56 25 57
rect 23 56 24 57
rect 22 56 23 57
rect 21 56 22 57
rect 20 56 21 57
rect 19 56 20 57
rect 18 56 19 57
rect 17 56 18 57
rect 16 56 17 57
rect 15 56 16 57
rect 14 56 15 57
rect 141 57 142 58
rect 140 57 141 58
rect 139 57 140 58
rect 138 57 139 58
rect 137 57 138 58
rect 136 57 137 58
rect 135 57 136 58
rect 134 57 135 58
rect 133 57 134 58
rect 126 57 127 58
rect 125 57 126 58
rect 124 57 125 58
rect 123 57 124 58
rect 122 57 123 58
rect 121 57 122 58
rect 120 57 121 58
rect 119 57 120 58
rect 118 57 119 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 73 57 74 58
rect 72 57 73 58
rect 71 57 72 58
rect 70 57 71 58
rect 69 57 70 58
rect 68 57 69 58
rect 67 57 68 58
rect 66 57 67 58
rect 65 57 66 58
rect 64 57 65 58
rect 30 57 31 58
rect 29 57 30 58
rect 28 57 29 58
rect 27 57 28 58
rect 26 57 27 58
rect 25 57 26 58
rect 24 57 25 58
rect 23 57 24 58
rect 22 57 23 58
rect 21 57 22 58
rect 20 57 21 58
rect 19 57 20 58
rect 18 57 19 58
rect 17 57 18 58
rect 16 57 17 58
rect 15 57 16 58
rect 14 57 15 58
rect 142 58 143 59
rect 141 58 142 59
rect 140 58 141 59
rect 139 58 140 59
rect 138 58 139 59
rect 137 58 138 59
rect 122 58 123 59
rect 121 58 122 59
rect 120 58 121 59
rect 119 58 120 59
rect 118 58 119 59
rect 117 58 118 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 73 58 74 59
rect 72 58 73 59
rect 71 58 72 59
rect 70 58 71 59
rect 69 58 70 59
rect 68 58 69 59
rect 67 58 68 59
rect 66 58 67 59
rect 65 58 66 59
rect 64 58 65 59
rect 30 58 31 59
rect 29 58 30 59
rect 28 58 29 59
rect 27 58 28 59
rect 26 58 27 59
rect 25 58 26 59
rect 24 58 25 59
rect 23 58 24 59
rect 22 58 23 59
rect 21 58 22 59
rect 20 58 21 59
rect 19 58 20 59
rect 18 58 19 59
rect 17 58 18 59
rect 16 58 17 59
rect 15 58 16 59
rect 14 58 15 59
rect 142 59 143 60
rect 141 59 142 60
rect 140 59 141 60
rect 139 59 140 60
rect 138 59 139 60
rect 121 59 122 60
rect 120 59 121 60
rect 119 59 120 60
rect 118 59 119 60
rect 117 59 118 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 72 59 73 60
rect 71 59 72 60
rect 70 59 71 60
rect 69 59 70 60
rect 68 59 69 60
rect 67 59 68 60
rect 66 59 67 60
rect 65 59 66 60
rect 64 59 65 60
rect 30 59 31 60
rect 29 59 30 60
rect 28 59 29 60
rect 27 59 28 60
rect 26 59 27 60
rect 25 59 26 60
rect 24 59 25 60
rect 23 59 24 60
rect 22 59 23 60
rect 21 59 22 60
rect 20 59 21 60
rect 19 59 20 60
rect 18 59 19 60
rect 17 59 18 60
rect 16 59 17 60
rect 15 59 16 60
rect 14 59 15 60
rect 142 60 143 61
rect 141 60 142 61
rect 140 60 141 61
rect 139 60 140 61
rect 120 60 121 61
rect 119 60 120 61
rect 118 60 119 61
rect 117 60 118 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 72 60 73 61
rect 71 60 72 61
rect 70 60 71 61
rect 69 60 70 61
rect 68 60 69 61
rect 67 60 68 61
rect 66 60 67 61
rect 65 60 66 61
rect 64 60 65 61
rect 63 60 64 61
rect 31 60 32 61
rect 30 60 31 61
rect 29 60 30 61
rect 28 60 29 61
rect 27 60 28 61
rect 26 60 27 61
rect 25 60 26 61
rect 24 60 25 61
rect 23 60 24 61
rect 22 60 23 61
rect 21 60 22 61
rect 20 60 21 61
rect 19 60 20 61
rect 18 60 19 61
rect 17 60 18 61
rect 16 60 17 61
rect 15 60 16 61
rect 14 60 15 61
rect 142 61 143 62
rect 141 61 142 62
rect 140 61 141 62
rect 139 61 140 62
rect 120 61 121 62
rect 119 61 120 62
rect 118 61 119 62
rect 117 61 118 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 71 61 72 62
rect 70 61 71 62
rect 69 61 70 62
rect 68 61 69 62
rect 67 61 68 62
rect 66 61 67 62
rect 65 61 66 62
rect 64 61 65 62
rect 63 61 64 62
rect 31 61 32 62
rect 30 61 31 62
rect 29 61 30 62
rect 28 61 29 62
rect 27 61 28 62
rect 26 61 27 62
rect 25 61 26 62
rect 24 61 25 62
rect 23 61 24 62
rect 22 61 23 62
rect 21 61 22 62
rect 20 61 21 62
rect 19 61 20 62
rect 18 61 19 62
rect 17 61 18 62
rect 16 61 17 62
rect 15 61 16 62
rect 14 61 15 62
rect 142 62 143 63
rect 141 62 142 63
rect 140 62 141 63
rect 139 62 140 63
rect 138 62 139 63
rect 121 62 122 63
rect 120 62 121 63
rect 119 62 120 63
rect 118 62 119 63
rect 117 62 118 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 71 62 72 63
rect 70 62 71 63
rect 69 62 70 63
rect 68 62 69 63
rect 67 62 68 63
rect 66 62 67 63
rect 65 62 66 63
rect 64 62 65 63
rect 63 62 64 63
rect 31 62 32 63
rect 30 62 31 63
rect 29 62 30 63
rect 28 62 29 63
rect 27 62 28 63
rect 26 62 27 63
rect 25 62 26 63
rect 24 62 25 63
rect 23 62 24 63
rect 22 62 23 63
rect 21 62 22 63
rect 20 62 21 63
rect 19 62 20 63
rect 18 62 19 63
rect 17 62 18 63
rect 16 62 17 63
rect 15 62 16 63
rect 14 62 15 63
rect 142 63 143 64
rect 141 63 142 64
rect 140 63 141 64
rect 139 63 140 64
rect 138 63 139 64
rect 137 63 138 64
rect 122 63 123 64
rect 121 63 122 64
rect 120 63 121 64
rect 119 63 120 64
rect 118 63 119 64
rect 117 63 118 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 70 63 71 64
rect 69 63 70 64
rect 68 63 69 64
rect 67 63 68 64
rect 66 63 67 64
rect 65 63 66 64
rect 64 63 65 64
rect 63 63 64 64
rect 62 63 63 64
rect 32 63 33 64
rect 31 63 32 64
rect 30 63 31 64
rect 29 63 30 64
rect 28 63 29 64
rect 27 63 28 64
rect 26 63 27 64
rect 25 63 26 64
rect 24 63 25 64
rect 23 63 24 64
rect 22 63 23 64
rect 21 63 22 64
rect 20 63 21 64
rect 19 63 20 64
rect 18 63 19 64
rect 17 63 18 64
rect 16 63 17 64
rect 15 63 16 64
rect 141 64 142 65
rect 140 64 141 65
rect 139 64 140 65
rect 138 64 139 65
rect 137 64 138 65
rect 136 64 137 65
rect 135 64 136 65
rect 134 64 135 65
rect 125 64 126 65
rect 124 64 125 65
rect 123 64 124 65
rect 122 64 123 65
rect 121 64 122 65
rect 120 64 121 65
rect 119 64 120 65
rect 118 64 119 65
rect 117 64 118 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 70 64 71 65
rect 69 64 70 65
rect 68 64 69 65
rect 67 64 68 65
rect 66 64 67 65
rect 65 64 66 65
rect 64 64 65 65
rect 63 64 64 65
rect 62 64 63 65
rect 32 64 33 65
rect 31 64 32 65
rect 30 64 31 65
rect 29 64 30 65
rect 28 64 29 65
rect 27 64 28 65
rect 26 64 27 65
rect 25 64 26 65
rect 24 64 25 65
rect 23 64 24 65
rect 22 64 23 65
rect 21 64 22 65
rect 20 64 21 65
rect 19 64 20 65
rect 18 64 19 65
rect 17 64 18 65
rect 16 64 17 65
rect 15 64 16 65
rect 141 65 142 66
rect 140 65 141 66
rect 139 65 140 66
rect 138 65 139 66
rect 137 65 138 66
rect 136 65 137 66
rect 135 65 136 66
rect 134 65 135 66
rect 133 65 134 66
rect 132 65 133 66
rect 131 65 132 66
rect 130 65 131 66
rect 129 65 130 66
rect 128 65 129 66
rect 127 65 128 66
rect 126 65 127 66
rect 125 65 126 66
rect 124 65 125 66
rect 123 65 124 66
rect 122 65 123 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 118 65 119 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 69 65 70 66
rect 68 65 69 66
rect 67 65 68 66
rect 66 65 67 66
rect 65 65 66 66
rect 64 65 65 66
rect 63 65 64 66
rect 62 65 63 66
rect 61 65 62 66
rect 33 65 34 66
rect 32 65 33 66
rect 31 65 32 66
rect 30 65 31 66
rect 29 65 30 66
rect 28 65 29 66
rect 27 65 28 66
rect 26 65 27 66
rect 25 65 26 66
rect 24 65 25 66
rect 23 65 24 66
rect 22 65 23 66
rect 21 65 22 66
rect 20 65 21 66
rect 19 65 20 66
rect 18 65 19 66
rect 17 65 18 66
rect 16 65 17 66
rect 15 65 16 66
rect 140 66 141 67
rect 139 66 140 67
rect 138 66 139 67
rect 137 66 138 67
rect 136 66 137 67
rect 135 66 136 67
rect 134 66 135 67
rect 133 66 134 67
rect 132 66 133 67
rect 131 66 132 67
rect 130 66 131 67
rect 129 66 130 67
rect 128 66 129 67
rect 127 66 128 67
rect 126 66 127 67
rect 125 66 126 67
rect 124 66 125 67
rect 123 66 124 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 118 66 119 67
rect 139 67 140 68
rect 138 67 139 68
rect 137 67 138 68
rect 136 67 137 68
rect 135 67 136 68
rect 134 67 135 68
rect 133 67 134 68
rect 132 67 133 68
rect 131 67 132 68
rect 130 67 131 68
rect 129 67 130 68
rect 128 67 129 68
rect 127 67 128 68
rect 126 67 127 68
rect 125 67 126 68
rect 124 67 125 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 119 67 120 68
rect 138 68 139 69
rect 137 68 138 69
rect 136 68 137 69
rect 135 68 136 69
rect 134 68 135 69
rect 133 68 134 69
rect 132 68 133 69
rect 131 68 132 69
rect 130 68 131 69
rect 129 68 130 69
rect 128 68 129 69
rect 127 68 128 69
rect 126 68 127 69
rect 125 68 126 69
rect 124 68 125 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 136 69 137 70
rect 135 69 136 70
rect 134 69 135 70
rect 133 69 134 70
rect 132 69 133 70
rect 131 69 132 70
rect 130 69 131 70
rect 129 69 130 70
rect 128 69 129 70
rect 127 69 128 70
rect 126 69 127 70
rect 125 69 126 70
rect 124 69 125 70
rect 123 69 124 70
rect 142 74 143 75
rect 141 74 142 75
rect 140 74 141 75
rect 139 74 140 75
rect 138 74 139 75
rect 137 74 138 75
rect 142 75 143 76
rect 141 75 142 76
rect 140 75 141 76
rect 139 75 140 76
rect 138 75 139 76
rect 137 75 138 76
rect 136 75 137 76
rect 135 75 136 76
rect 122 75 123 76
rect 121 75 122 76
rect 120 75 121 76
rect 119 75 120 76
rect 142 76 143 77
rect 141 76 142 77
rect 140 76 141 77
rect 139 76 140 77
rect 138 76 139 77
rect 137 76 138 77
rect 136 76 137 77
rect 135 76 136 77
rect 134 76 135 77
rect 122 76 123 77
rect 121 76 122 77
rect 120 76 121 77
rect 119 76 120 77
rect 118 76 119 77
rect 80 76 81 77
rect 79 76 80 77
rect 78 76 79 77
rect 77 76 78 77
rect 76 76 77 77
rect 75 76 76 77
rect 74 76 75 77
rect 73 76 74 77
rect 72 76 73 77
rect 71 76 72 77
rect 70 76 71 77
rect 69 76 70 77
rect 68 76 69 77
rect 67 76 68 77
rect 66 76 67 77
rect 65 76 66 77
rect 64 76 65 77
rect 63 76 64 77
rect 62 76 63 77
rect 61 76 62 77
rect 60 76 61 77
rect 59 76 60 77
rect 58 76 59 77
rect 57 76 58 77
rect 56 76 57 77
rect 55 76 56 77
rect 54 76 55 77
rect 53 76 54 77
rect 52 76 53 77
rect 51 76 52 77
rect 50 76 51 77
rect 49 76 50 77
rect 48 76 49 77
rect 47 76 48 77
rect 46 76 47 77
rect 45 76 46 77
rect 44 76 45 77
rect 43 76 44 77
rect 42 76 43 77
rect 41 76 42 77
rect 40 76 41 77
rect 39 76 40 77
rect 38 76 39 77
rect 37 76 38 77
rect 36 76 37 77
rect 35 76 36 77
rect 34 76 35 77
rect 33 76 34 77
rect 32 76 33 77
rect 31 76 32 77
rect 30 76 31 77
rect 29 76 30 77
rect 28 76 29 77
rect 27 76 28 77
rect 26 76 27 77
rect 25 76 26 77
rect 24 76 25 77
rect 23 76 24 77
rect 22 76 23 77
rect 21 76 22 77
rect 20 76 21 77
rect 19 76 20 77
rect 18 76 19 77
rect 17 76 18 77
rect 16 76 17 77
rect 15 76 16 77
rect 14 76 15 77
rect 142 77 143 78
rect 141 77 142 78
rect 140 77 141 78
rect 139 77 140 78
rect 138 77 139 78
rect 137 77 138 78
rect 136 77 137 78
rect 135 77 136 78
rect 134 77 135 78
rect 133 77 134 78
rect 121 77 122 78
rect 120 77 121 78
rect 119 77 120 78
rect 118 77 119 78
rect 80 77 81 78
rect 79 77 80 78
rect 78 77 79 78
rect 77 77 78 78
rect 76 77 77 78
rect 75 77 76 78
rect 74 77 75 78
rect 73 77 74 78
rect 72 77 73 78
rect 71 77 72 78
rect 70 77 71 78
rect 69 77 70 78
rect 68 77 69 78
rect 67 77 68 78
rect 66 77 67 78
rect 65 77 66 78
rect 64 77 65 78
rect 63 77 64 78
rect 62 77 63 78
rect 61 77 62 78
rect 60 77 61 78
rect 59 77 60 78
rect 58 77 59 78
rect 57 77 58 78
rect 56 77 57 78
rect 55 77 56 78
rect 54 77 55 78
rect 53 77 54 78
rect 52 77 53 78
rect 51 77 52 78
rect 50 77 51 78
rect 49 77 50 78
rect 48 77 49 78
rect 47 77 48 78
rect 46 77 47 78
rect 45 77 46 78
rect 44 77 45 78
rect 43 77 44 78
rect 42 77 43 78
rect 41 77 42 78
rect 40 77 41 78
rect 39 77 40 78
rect 38 77 39 78
rect 37 77 38 78
rect 36 77 37 78
rect 35 77 36 78
rect 34 77 35 78
rect 33 77 34 78
rect 32 77 33 78
rect 31 77 32 78
rect 30 77 31 78
rect 29 77 30 78
rect 28 77 29 78
rect 27 77 28 78
rect 26 77 27 78
rect 25 77 26 78
rect 24 77 25 78
rect 23 77 24 78
rect 22 77 23 78
rect 21 77 22 78
rect 20 77 21 78
rect 19 77 20 78
rect 18 77 19 78
rect 17 77 18 78
rect 16 77 17 78
rect 15 77 16 78
rect 14 77 15 78
rect 142 78 143 79
rect 141 78 142 79
rect 140 78 141 79
rect 139 78 140 79
rect 138 78 139 79
rect 137 78 138 79
rect 136 78 137 79
rect 135 78 136 79
rect 134 78 135 79
rect 133 78 134 79
rect 132 78 133 79
rect 121 78 122 79
rect 120 78 121 79
rect 119 78 120 79
rect 118 78 119 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 66 78 67 79
rect 65 78 66 79
rect 64 78 65 79
rect 63 78 64 79
rect 62 78 63 79
rect 61 78 62 79
rect 60 78 61 79
rect 59 78 60 79
rect 58 78 59 79
rect 57 78 58 79
rect 56 78 57 79
rect 55 78 56 79
rect 54 78 55 79
rect 53 78 54 79
rect 52 78 53 79
rect 51 78 52 79
rect 50 78 51 79
rect 49 78 50 79
rect 48 78 49 79
rect 47 78 48 79
rect 46 78 47 79
rect 45 78 46 79
rect 44 78 45 79
rect 43 78 44 79
rect 42 78 43 79
rect 41 78 42 79
rect 40 78 41 79
rect 39 78 40 79
rect 38 78 39 79
rect 37 78 38 79
rect 36 78 37 79
rect 35 78 36 79
rect 34 78 35 79
rect 33 78 34 79
rect 32 78 33 79
rect 31 78 32 79
rect 30 78 31 79
rect 29 78 30 79
rect 28 78 29 79
rect 27 78 28 79
rect 26 78 27 79
rect 25 78 26 79
rect 24 78 25 79
rect 23 78 24 79
rect 22 78 23 79
rect 21 78 22 79
rect 20 78 21 79
rect 19 78 20 79
rect 18 78 19 79
rect 17 78 18 79
rect 16 78 17 79
rect 15 78 16 79
rect 14 78 15 79
rect 142 79 143 80
rect 141 79 142 80
rect 140 79 141 80
rect 139 79 140 80
rect 138 79 139 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 134 79 135 80
rect 133 79 134 80
rect 132 79 133 80
rect 121 79 122 80
rect 120 79 121 80
rect 119 79 120 80
rect 118 79 119 80
rect 117 79 118 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 65 79 66 80
rect 64 79 65 80
rect 63 79 64 80
rect 62 79 63 80
rect 61 79 62 80
rect 60 79 61 80
rect 59 79 60 80
rect 58 79 59 80
rect 57 79 58 80
rect 56 79 57 80
rect 55 79 56 80
rect 54 79 55 80
rect 53 79 54 80
rect 52 79 53 80
rect 51 79 52 80
rect 50 79 51 80
rect 49 79 50 80
rect 48 79 49 80
rect 47 79 48 80
rect 46 79 47 80
rect 45 79 46 80
rect 44 79 45 80
rect 43 79 44 80
rect 42 79 43 80
rect 41 79 42 80
rect 40 79 41 80
rect 39 79 40 80
rect 38 79 39 80
rect 37 79 38 80
rect 36 79 37 80
rect 35 79 36 80
rect 34 79 35 80
rect 33 79 34 80
rect 32 79 33 80
rect 31 79 32 80
rect 30 79 31 80
rect 29 79 30 80
rect 28 79 29 80
rect 27 79 28 80
rect 26 79 27 80
rect 25 79 26 80
rect 24 79 25 80
rect 23 79 24 80
rect 22 79 23 80
rect 21 79 22 80
rect 20 79 21 80
rect 19 79 20 80
rect 18 79 19 80
rect 17 79 18 80
rect 16 79 17 80
rect 15 79 16 80
rect 14 79 15 80
rect 142 80 143 81
rect 141 80 142 81
rect 140 80 141 81
rect 139 80 140 81
rect 138 80 139 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 133 80 134 81
rect 132 80 133 81
rect 131 80 132 81
rect 120 80 121 81
rect 119 80 120 81
rect 118 80 119 81
rect 117 80 118 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 61 80 62 81
rect 60 80 61 81
rect 59 80 60 81
rect 58 80 59 81
rect 57 80 58 81
rect 56 80 57 81
rect 55 80 56 81
rect 54 80 55 81
rect 53 80 54 81
rect 52 80 53 81
rect 51 80 52 81
rect 50 80 51 81
rect 49 80 50 81
rect 48 80 49 81
rect 47 80 48 81
rect 46 80 47 81
rect 45 80 46 81
rect 44 80 45 81
rect 43 80 44 81
rect 42 80 43 81
rect 41 80 42 81
rect 40 80 41 81
rect 39 80 40 81
rect 38 80 39 81
rect 37 80 38 81
rect 36 80 37 81
rect 35 80 36 81
rect 34 80 35 81
rect 33 80 34 81
rect 32 80 33 81
rect 31 80 32 81
rect 30 80 31 81
rect 29 80 30 81
rect 28 80 29 81
rect 27 80 28 81
rect 26 80 27 81
rect 25 80 26 81
rect 24 80 25 81
rect 23 80 24 81
rect 22 80 23 81
rect 21 80 22 81
rect 20 80 21 81
rect 19 80 20 81
rect 18 80 19 81
rect 17 80 18 81
rect 16 80 17 81
rect 15 80 16 81
rect 14 80 15 81
rect 142 81 143 82
rect 141 81 142 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 135 81 136 82
rect 134 81 135 82
rect 133 81 134 82
rect 132 81 133 82
rect 131 81 132 82
rect 130 81 131 82
rect 120 81 121 82
rect 119 81 120 82
rect 118 81 119 82
rect 117 81 118 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 61 81 62 82
rect 60 81 61 82
rect 59 81 60 82
rect 58 81 59 82
rect 57 81 58 82
rect 56 81 57 82
rect 55 81 56 82
rect 54 81 55 82
rect 53 81 54 82
rect 52 81 53 82
rect 51 81 52 82
rect 50 81 51 82
rect 49 81 50 82
rect 48 81 49 82
rect 47 81 48 82
rect 46 81 47 82
rect 45 81 46 82
rect 44 81 45 82
rect 43 81 44 82
rect 42 81 43 82
rect 41 81 42 82
rect 40 81 41 82
rect 39 81 40 82
rect 38 81 39 82
rect 37 81 38 82
rect 36 81 37 82
rect 35 81 36 82
rect 34 81 35 82
rect 33 81 34 82
rect 32 81 33 82
rect 31 81 32 82
rect 30 81 31 82
rect 29 81 30 82
rect 28 81 29 82
rect 27 81 28 82
rect 26 81 27 82
rect 25 81 26 82
rect 24 81 25 82
rect 23 81 24 82
rect 22 81 23 82
rect 21 81 22 82
rect 20 81 21 82
rect 19 81 20 82
rect 18 81 19 82
rect 17 81 18 82
rect 16 81 17 82
rect 15 81 16 82
rect 14 81 15 82
rect 142 82 143 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 134 82 135 83
rect 133 82 134 83
rect 132 82 133 83
rect 131 82 132 83
rect 130 82 131 83
rect 129 82 130 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 118 82 119 83
rect 117 82 118 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 60 82 61 83
rect 59 82 60 83
rect 58 82 59 83
rect 57 82 58 83
rect 56 82 57 83
rect 55 82 56 83
rect 54 82 55 83
rect 53 82 54 83
rect 52 82 53 83
rect 51 82 52 83
rect 50 82 51 83
rect 49 82 50 83
rect 48 82 49 83
rect 47 82 48 83
rect 46 82 47 83
rect 45 82 46 83
rect 44 82 45 83
rect 43 82 44 83
rect 42 82 43 83
rect 41 82 42 83
rect 40 82 41 83
rect 39 82 40 83
rect 38 82 39 83
rect 37 82 38 83
rect 36 82 37 83
rect 35 82 36 83
rect 34 82 35 83
rect 33 82 34 83
rect 32 82 33 83
rect 31 82 32 83
rect 30 82 31 83
rect 29 82 30 83
rect 28 82 29 83
rect 27 82 28 83
rect 26 82 27 83
rect 25 82 26 83
rect 24 82 25 83
rect 23 82 24 83
rect 22 82 23 83
rect 21 82 22 83
rect 20 82 21 83
rect 19 82 20 83
rect 18 82 19 83
rect 17 82 18 83
rect 16 82 17 83
rect 15 82 16 83
rect 14 82 15 83
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 133 83 134 84
rect 132 83 133 84
rect 131 83 132 84
rect 130 83 131 84
rect 129 83 130 84
rect 128 83 129 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 118 83 119 84
rect 117 83 118 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 59 83 60 84
rect 58 83 59 84
rect 57 83 58 84
rect 56 83 57 84
rect 55 83 56 84
rect 54 83 55 84
rect 53 83 54 84
rect 52 83 53 84
rect 51 83 52 84
rect 50 83 51 84
rect 49 83 50 84
rect 48 83 49 84
rect 47 83 48 84
rect 46 83 47 84
rect 45 83 46 84
rect 44 83 45 84
rect 43 83 44 84
rect 42 83 43 84
rect 41 83 42 84
rect 40 83 41 84
rect 39 83 40 84
rect 38 83 39 84
rect 37 83 38 84
rect 36 83 37 84
rect 35 83 36 84
rect 34 83 35 84
rect 33 83 34 84
rect 32 83 33 84
rect 31 83 32 84
rect 30 83 31 84
rect 29 83 30 84
rect 28 83 29 84
rect 27 83 28 84
rect 26 83 27 84
rect 25 83 26 84
rect 24 83 25 84
rect 23 83 24 84
rect 22 83 23 84
rect 21 83 22 84
rect 20 83 21 84
rect 19 83 20 84
rect 18 83 19 84
rect 17 83 18 84
rect 16 83 17 84
rect 15 83 16 84
rect 14 83 15 84
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 130 84 131 85
rect 129 84 130 85
rect 128 84 129 85
rect 127 84 128 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 118 84 119 85
rect 117 84 118 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 59 84 60 85
rect 58 84 59 85
rect 57 84 58 85
rect 56 84 57 85
rect 55 84 56 85
rect 54 84 55 85
rect 53 84 54 85
rect 52 84 53 85
rect 51 84 52 85
rect 50 84 51 85
rect 49 84 50 85
rect 48 84 49 85
rect 47 84 48 85
rect 46 84 47 85
rect 45 84 46 85
rect 44 84 45 85
rect 43 84 44 85
rect 42 84 43 85
rect 41 84 42 85
rect 40 84 41 85
rect 39 84 40 85
rect 38 84 39 85
rect 37 84 38 85
rect 36 84 37 85
rect 35 84 36 85
rect 34 84 35 85
rect 33 84 34 85
rect 32 84 33 85
rect 31 84 32 85
rect 30 84 31 85
rect 29 84 30 85
rect 28 84 29 85
rect 27 84 28 85
rect 26 84 27 85
rect 25 84 26 85
rect 24 84 25 85
rect 23 84 24 85
rect 22 84 23 85
rect 21 84 22 85
rect 20 84 21 85
rect 19 84 20 85
rect 18 84 19 85
rect 17 84 18 85
rect 16 84 17 85
rect 15 84 16 85
rect 14 84 15 85
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 139 85 140 86
rect 138 85 139 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 129 85 130 86
rect 128 85 129 86
rect 127 85 128 86
rect 126 85 127 86
rect 125 85 126 86
rect 124 85 125 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 118 85 119 86
rect 117 85 118 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 58 85 59 86
rect 57 85 58 86
rect 56 85 57 86
rect 55 85 56 86
rect 54 85 55 86
rect 53 85 54 86
rect 52 85 53 86
rect 51 85 52 86
rect 50 85 51 86
rect 49 85 50 86
rect 48 85 49 86
rect 47 85 48 86
rect 46 85 47 86
rect 45 85 46 86
rect 44 85 45 86
rect 43 85 44 86
rect 42 85 43 86
rect 41 85 42 86
rect 40 85 41 86
rect 39 85 40 86
rect 38 85 39 86
rect 37 85 38 86
rect 36 85 37 86
rect 35 85 36 86
rect 34 85 35 86
rect 33 85 34 86
rect 32 85 33 86
rect 31 85 32 86
rect 30 85 31 86
rect 29 85 30 86
rect 28 85 29 86
rect 27 85 28 86
rect 26 85 27 86
rect 25 85 26 86
rect 24 85 25 86
rect 23 85 24 86
rect 22 85 23 86
rect 21 85 22 86
rect 20 85 21 86
rect 19 85 20 86
rect 18 85 19 86
rect 17 85 18 86
rect 16 85 17 86
rect 15 85 16 86
rect 14 85 15 86
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 139 86 140 87
rect 138 86 139 87
rect 131 86 132 87
rect 130 86 131 87
rect 129 86 130 87
rect 128 86 129 87
rect 127 86 128 87
rect 126 86 127 87
rect 125 86 126 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 118 86 119 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 57 86 58 87
rect 56 86 57 87
rect 55 86 56 87
rect 54 86 55 87
rect 53 86 54 87
rect 52 86 53 87
rect 51 86 52 87
rect 50 86 51 87
rect 49 86 50 87
rect 48 86 49 87
rect 47 86 48 87
rect 46 86 47 87
rect 45 86 46 87
rect 44 86 45 87
rect 43 86 44 87
rect 42 86 43 87
rect 41 86 42 87
rect 40 86 41 87
rect 39 86 40 87
rect 38 86 39 87
rect 37 86 38 87
rect 36 86 37 87
rect 35 86 36 87
rect 34 86 35 87
rect 33 86 34 87
rect 32 86 33 87
rect 31 86 32 87
rect 30 86 31 87
rect 29 86 30 87
rect 28 86 29 87
rect 27 86 28 87
rect 26 86 27 87
rect 25 86 26 87
rect 24 86 25 87
rect 23 86 24 87
rect 22 86 23 87
rect 21 86 22 87
rect 20 86 21 87
rect 19 86 20 87
rect 18 86 19 87
rect 17 86 18 87
rect 16 86 17 87
rect 15 86 16 87
rect 14 86 15 87
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 139 87 140 88
rect 138 87 139 88
rect 130 87 131 88
rect 129 87 130 88
rect 128 87 129 88
rect 127 87 128 88
rect 126 87 127 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 118 87 119 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 57 87 58 88
rect 56 87 57 88
rect 55 87 56 88
rect 54 87 55 88
rect 53 87 54 88
rect 52 87 53 88
rect 51 87 52 88
rect 50 87 51 88
rect 49 87 50 88
rect 48 87 49 88
rect 47 87 48 88
rect 46 87 47 88
rect 45 87 46 88
rect 44 87 45 88
rect 43 87 44 88
rect 42 87 43 88
rect 41 87 42 88
rect 40 87 41 88
rect 39 87 40 88
rect 38 87 39 88
rect 37 87 38 88
rect 36 87 37 88
rect 35 87 36 88
rect 34 87 35 88
rect 33 87 34 88
rect 32 87 33 88
rect 31 87 32 88
rect 30 87 31 88
rect 29 87 30 88
rect 28 87 29 88
rect 27 87 28 88
rect 26 87 27 88
rect 25 87 26 88
rect 24 87 25 88
rect 23 87 24 88
rect 22 87 23 88
rect 21 87 22 88
rect 20 87 21 88
rect 19 87 20 88
rect 18 87 19 88
rect 17 87 18 88
rect 16 87 17 88
rect 15 87 16 88
rect 14 87 15 88
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 139 88 140 89
rect 138 88 139 89
rect 129 88 130 89
rect 128 88 129 89
rect 127 88 128 89
rect 126 88 127 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 119 88 120 89
rect 80 88 81 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 56 88 57 89
rect 55 88 56 89
rect 54 88 55 89
rect 53 88 54 89
rect 52 88 53 89
rect 51 88 52 89
rect 50 88 51 89
rect 49 88 50 89
rect 48 88 49 89
rect 47 88 48 89
rect 46 88 47 89
rect 45 88 46 89
rect 44 88 45 89
rect 43 88 44 89
rect 42 88 43 89
rect 41 88 42 89
rect 40 88 41 89
rect 39 88 40 89
rect 38 88 39 89
rect 37 88 38 89
rect 36 88 37 89
rect 35 88 36 89
rect 34 88 35 89
rect 33 88 34 89
rect 32 88 33 89
rect 31 88 32 89
rect 30 88 31 89
rect 29 88 30 89
rect 28 88 29 89
rect 27 88 28 89
rect 26 88 27 89
rect 25 88 26 89
rect 24 88 25 89
rect 23 88 24 89
rect 22 88 23 89
rect 21 88 22 89
rect 20 88 21 89
rect 19 88 20 89
rect 18 88 19 89
rect 17 88 18 89
rect 16 88 17 89
rect 15 88 16 89
rect 14 88 15 89
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 139 89 140 90
rect 138 89 139 90
rect 128 89 129 90
rect 127 89 128 90
rect 126 89 127 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 80 89 81 90
rect 79 89 80 90
rect 78 89 79 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 55 89 56 90
rect 54 89 55 90
rect 53 89 54 90
rect 52 89 53 90
rect 51 89 52 90
rect 50 89 51 90
rect 49 89 50 90
rect 48 89 49 90
rect 47 89 48 90
rect 46 89 47 90
rect 45 89 46 90
rect 44 89 45 90
rect 43 89 44 90
rect 42 89 43 90
rect 41 89 42 90
rect 40 89 41 90
rect 39 89 40 90
rect 38 89 39 90
rect 37 89 38 90
rect 36 89 37 90
rect 35 89 36 90
rect 34 89 35 90
rect 33 89 34 90
rect 32 89 33 90
rect 31 89 32 90
rect 30 89 31 90
rect 29 89 30 90
rect 28 89 29 90
rect 27 89 28 90
rect 26 89 27 90
rect 25 89 26 90
rect 24 89 25 90
rect 23 89 24 90
rect 22 89 23 90
rect 21 89 22 90
rect 20 89 21 90
rect 19 89 20 90
rect 18 89 19 90
rect 17 89 18 90
rect 16 89 17 90
rect 15 89 16 90
rect 14 89 15 90
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 139 90 140 91
rect 138 90 139 91
rect 125 90 126 91
rect 124 90 125 91
rect 123 90 124 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 77 90 78 91
rect 76 90 77 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 55 90 56 91
rect 54 90 55 91
rect 53 90 54 91
rect 52 90 53 91
rect 51 90 52 91
rect 50 90 51 91
rect 49 90 50 91
rect 48 90 49 91
rect 47 90 48 91
rect 46 90 47 91
rect 45 90 46 91
rect 44 90 45 91
rect 43 90 44 91
rect 42 90 43 91
rect 41 90 42 91
rect 40 90 41 91
rect 39 90 40 91
rect 38 90 39 91
rect 37 90 38 91
rect 36 90 37 91
rect 35 90 36 91
rect 34 90 35 91
rect 33 90 34 91
rect 32 90 33 91
rect 31 90 32 91
rect 30 90 31 91
rect 29 90 30 91
rect 28 90 29 91
rect 27 90 28 91
rect 26 90 27 91
rect 25 90 26 91
rect 24 90 25 91
rect 23 90 24 91
rect 22 90 23 91
rect 21 90 22 91
rect 20 90 21 91
rect 19 90 20 91
rect 18 90 19 91
rect 17 90 18 91
rect 16 90 17 91
rect 15 90 16 91
rect 14 90 15 91
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 74 91 75 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 54 91 55 92
rect 53 91 54 92
rect 52 91 53 92
rect 51 91 52 92
rect 50 91 51 92
rect 49 91 50 92
rect 48 91 49 92
rect 47 91 48 92
rect 46 91 47 92
rect 45 91 46 92
rect 44 91 45 92
rect 43 91 44 92
rect 42 91 43 92
rect 41 91 42 92
rect 40 91 41 92
rect 39 91 40 92
rect 38 91 39 92
rect 37 91 38 92
rect 36 91 37 92
rect 35 91 36 92
rect 34 91 35 92
rect 33 91 34 92
rect 32 91 33 92
rect 31 91 32 92
rect 30 91 31 92
rect 29 91 30 92
rect 28 91 29 92
rect 27 91 28 92
rect 26 91 27 92
rect 25 91 26 92
rect 24 91 25 92
rect 23 91 24 92
rect 22 91 23 92
rect 21 91 22 92
rect 20 91 21 92
rect 19 91 20 92
rect 18 91 19 92
rect 17 91 18 92
rect 16 91 17 92
rect 15 91 16 92
rect 14 91 15 92
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 72 92 73 93
rect 71 92 72 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 53 92 54 93
rect 52 92 53 93
rect 51 92 52 93
rect 50 92 51 93
rect 49 92 50 93
rect 48 92 49 93
rect 47 92 48 93
rect 46 92 47 93
rect 45 92 46 93
rect 44 92 45 93
rect 43 92 44 93
rect 42 92 43 93
rect 41 92 42 93
rect 40 92 41 93
rect 39 92 40 93
rect 38 92 39 93
rect 37 92 38 93
rect 36 92 37 93
rect 35 92 36 93
rect 34 92 35 93
rect 33 92 34 93
rect 32 92 33 93
rect 31 92 32 93
rect 30 92 31 93
rect 29 92 30 93
rect 28 92 29 93
rect 27 92 28 93
rect 26 92 27 93
rect 25 92 26 93
rect 24 92 25 93
rect 23 92 24 93
rect 22 92 23 93
rect 21 92 22 93
rect 20 92 21 93
rect 19 92 20 93
rect 18 92 19 93
rect 17 92 18 93
rect 16 92 17 93
rect 15 92 16 93
rect 14 92 15 93
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 70 93 71 94
rect 69 93 70 94
rect 68 93 69 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 52 93 53 94
rect 51 93 52 94
rect 50 93 51 94
rect 49 93 50 94
rect 48 93 49 94
rect 47 93 48 94
rect 46 93 47 94
rect 45 93 46 94
rect 44 93 45 94
rect 43 93 44 94
rect 42 93 43 94
rect 41 93 42 94
rect 40 93 41 94
rect 39 93 40 94
rect 38 93 39 94
rect 37 93 38 94
rect 36 93 37 94
rect 35 93 36 94
rect 34 93 35 94
rect 33 93 34 94
rect 32 93 33 94
rect 31 93 32 94
rect 30 93 31 94
rect 29 93 30 94
rect 28 93 29 94
rect 27 93 28 94
rect 26 93 27 94
rect 25 93 26 94
rect 24 93 25 94
rect 23 93 24 94
rect 22 93 23 94
rect 21 93 22 94
rect 20 93 21 94
rect 19 93 20 94
rect 18 93 19 94
rect 17 93 18 94
rect 16 93 17 94
rect 15 93 16 94
rect 14 93 15 94
rect 137 94 138 95
rect 136 94 137 95
rect 135 94 136 95
rect 134 94 135 95
rect 133 94 134 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 68 94 69 95
rect 67 94 68 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 51 94 52 95
rect 50 94 51 95
rect 49 94 50 95
rect 48 94 49 95
rect 47 94 48 95
rect 46 94 47 95
rect 45 94 46 95
rect 44 94 45 95
rect 43 94 44 95
rect 42 94 43 95
rect 41 94 42 95
rect 40 94 41 95
rect 39 94 40 95
rect 38 94 39 95
rect 37 94 38 95
rect 36 94 37 95
rect 35 94 36 95
rect 34 94 35 95
rect 33 94 34 95
rect 32 94 33 95
rect 31 94 32 95
rect 30 94 31 95
rect 29 94 30 95
rect 28 94 29 95
rect 27 94 28 95
rect 26 94 27 95
rect 25 94 26 95
rect 24 94 25 95
rect 23 94 24 95
rect 22 94 23 95
rect 21 94 22 95
rect 20 94 21 95
rect 19 94 20 95
rect 18 94 19 95
rect 17 94 18 95
rect 16 94 17 95
rect 15 94 16 95
rect 14 94 15 95
rect 137 95 138 96
rect 136 95 137 96
rect 135 95 136 96
rect 134 95 135 96
rect 133 95 134 96
rect 132 95 133 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 72 95 73 96
rect 71 95 72 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 67 95 68 96
rect 66 95 67 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 50 95 51 96
rect 49 95 50 96
rect 48 95 49 96
rect 47 95 48 96
rect 46 95 47 96
rect 45 95 46 96
rect 44 95 45 96
rect 43 95 44 96
rect 42 95 43 96
rect 41 95 42 96
rect 40 95 41 96
rect 39 95 40 96
rect 38 95 39 96
rect 37 95 38 96
rect 36 95 37 96
rect 35 95 36 96
rect 34 95 35 96
rect 33 95 34 96
rect 32 95 33 96
rect 31 95 32 96
rect 30 95 31 96
rect 29 95 30 96
rect 28 95 29 96
rect 27 95 28 96
rect 26 95 27 96
rect 25 95 26 96
rect 24 95 25 96
rect 23 95 24 96
rect 22 95 23 96
rect 21 95 22 96
rect 20 95 21 96
rect 19 95 20 96
rect 18 95 19 96
rect 17 95 18 96
rect 16 95 17 96
rect 15 95 16 96
rect 14 95 15 96
rect 137 96 138 97
rect 136 96 137 97
rect 135 96 136 97
rect 134 96 135 97
rect 133 96 134 97
rect 132 96 133 97
rect 131 96 132 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 49 96 50 97
rect 48 96 49 97
rect 47 96 48 97
rect 46 96 47 97
rect 45 96 46 97
rect 27 96 28 97
rect 26 96 27 97
rect 25 96 26 97
rect 24 96 25 97
rect 23 96 24 97
rect 22 96 23 97
rect 21 96 22 97
rect 20 96 21 97
rect 19 96 20 97
rect 18 96 19 97
rect 17 96 18 97
rect 16 96 17 97
rect 15 96 16 97
rect 14 96 15 97
rect 137 97 138 98
rect 136 97 137 98
rect 135 97 136 98
rect 134 97 135 98
rect 133 97 134 98
rect 132 97 133 98
rect 131 97 132 98
rect 130 97 131 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 50 97 51 98
rect 49 97 50 98
rect 48 97 49 98
rect 47 97 48 98
rect 46 97 47 98
rect 45 97 46 98
rect 27 97 28 98
rect 26 97 27 98
rect 25 97 26 98
rect 24 97 25 98
rect 23 97 24 98
rect 22 97 23 98
rect 21 97 22 98
rect 20 97 21 98
rect 19 97 20 98
rect 18 97 19 98
rect 17 97 18 98
rect 16 97 17 98
rect 15 97 16 98
rect 14 97 15 98
rect 137 98 138 99
rect 136 98 137 99
rect 135 98 136 99
rect 134 98 135 99
rect 133 98 134 99
rect 132 98 133 99
rect 131 98 132 99
rect 130 98 131 99
rect 129 98 130 99
rect 128 98 129 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 51 98 52 99
rect 50 98 51 99
rect 49 98 50 99
rect 48 98 49 99
rect 47 98 48 99
rect 46 98 47 99
rect 45 98 46 99
rect 27 98 28 99
rect 26 98 27 99
rect 25 98 26 99
rect 24 98 25 99
rect 23 98 24 99
rect 22 98 23 99
rect 21 98 22 99
rect 20 98 21 99
rect 19 98 20 99
rect 18 98 19 99
rect 17 98 18 99
rect 16 98 17 99
rect 15 98 16 99
rect 14 98 15 99
rect 137 99 138 100
rect 136 99 137 100
rect 135 99 136 100
rect 134 99 135 100
rect 133 99 134 100
rect 132 99 133 100
rect 131 99 132 100
rect 130 99 131 100
rect 129 99 130 100
rect 128 99 129 100
rect 127 99 128 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 51 99 52 100
rect 50 99 51 100
rect 49 99 50 100
rect 48 99 49 100
rect 47 99 48 100
rect 46 99 47 100
rect 45 99 46 100
rect 27 99 28 100
rect 26 99 27 100
rect 25 99 26 100
rect 24 99 25 100
rect 23 99 24 100
rect 22 99 23 100
rect 21 99 22 100
rect 20 99 21 100
rect 19 99 20 100
rect 18 99 19 100
rect 17 99 18 100
rect 16 99 17 100
rect 15 99 16 100
rect 14 99 15 100
rect 137 100 138 101
rect 136 100 137 101
rect 135 100 136 101
rect 134 100 135 101
rect 131 100 132 101
rect 130 100 131 101
rect 129 100 130 101
rect 128 100 129 101
rect 127 100 128 101
rect 126 100 127 101
rect 125 100 126 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 51 100 52 101
rect 50 100 51 101
rect 49 100 50 101
rect 48 100 49 101
rect 47 100 48 101
rect 46 100 47 101
rect 45 100 46 101
rect 27 100 28 101
rect 26 100 27 101
rect 25 100 26 101
rect 24 100 25 101
rect 23 100 24 101
rect 22 100 23 101
rect 21 100 22 101
rect 20 100 21 101
rect 19 100 20 101
rect 18 100 19 101
rect 17 100 18 101
rect 16 100 17 101
rect 15 100 16 101
rect 14 100 15 101
rect 137 101 138 102
rect 136 101 137 102
rect 135 101 136 102
rect 134 101 135 102
rect 130 101 131 102
rect 129 101 130 102
rect 128 101 129 102
rect 127 101 128 102
rect 126 101 127 102
rect 125 101 126 102
rect 124 101 125 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 51 101 52 102
rect 50 101 51 102
rect 49 101 50 102
rect 48 101 49 102
rect 47 101 48 102
rect 46 101 47 102
rect 45 101 46 102
rect 27 101 28 102
rect 26 101 27 102
rect 25 101 26 102
rect 24 101 25 102
rect 23 101 24 102
rect 22 101 23 102
rect 21 101 22 102
rect 20 101 21 102
rect 19 101 20 102
rect 18 101 19 102
rect 17 101 18 102
rect 16 101 17 102
rect 15 101 16 102
rect 14 101 15 102
rect 137 102 138 103
rect 136 102 137 103
rect 135 102 136 103
rect 134 102 135 103
rect 128 102 129 103
rect 127 102 128 103
rect 126 102 127 103
rect 125 102 126 103
rect 124 102 125 103
rect 123 102 124 103
rect 122 102 123 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 51 102 52 103
rect 50 102 51 103
rect 49 102 50 103
rect 48 102 49 103
rect 47 102 48 103
rect 46 102 47 103
rect 45 102 46 103
rect 27 102 28 103
rect 26 102 27 103
rect 25 102 26 103
rect 24 102 25 103
rect 23 102 24 103
rect 22 102 23 103
rect 21 102 22 103
rect 20 102 21 103
rect 19 102 20 103
rect 18 102 19 103
rect 17 102 18 103
rect 16 102 17 103
rect 15 102 16 103
rect 14 102 15 103
rect 137 103 138 104
rect 136 103 137 104
rect 135 103 136 104
rect 134 103 135 104
rect 127 103 128 104
rect 126 103 127 104
rect 125 103 126 104
rect 124 103 125 104
rect 123 103 124 104
rect 122 103 123 104
rect 121 103 122 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 50 103 51 104
rect 49 103 50 104
rect 48 103 49 104
rect 47 103 48 104
rect 46 103 47 104
rect 45 103 46 104
rect 27 103 28 104
rect 26 103 27 104
rect 25 103 26 104
rect 24 103 25 104
rect 23 103 24 104
rect 22 103 23 104
rect 21 103 22 104
rect 20 103 21 104
rect 19 103 20 104
rect 18 103 19 104
rect 17 103 18 104
rect 16 103 17 104
rect 15 103 16 104
rect 14 103 15 104
rect 137 104 138 105
rect 136 104 137 105
rect 135 104 136 105
rect 134 104 135 105
rect 125 104 126 105
rect 124 104 125 105
rect 123 104 124 105
rect 122 104 123 105
rect 121 104 122 105
rect 120 104 121 105
rect 119 104 120 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 51 104 52 105
rect 50 104 51 105
rect 49 104 50 105
rect 48 104 49 105
rect 47 104 48 105
rect 46 104 47 105
rect 45 104 46 105
rect 28 104 29 105
rect 27 104 28 105
rect 26 104 27 105
rect 25 104 26 105
rect 24 104 25 105
rect 23 104 24 105
rect 22 104 23 105
rect 21 104 22 105
rect 20 104 21 105
rect 19 104 20 105
rect 18 104 19 105
rect 17 104 18 105
rect 16 104 17 105
rect 15 104 16 105
rect 14 104 15 105
rect 137 105 138 106
rect 136 105 137 106
rect 135 105 136 106
rect 134 105 135 106
rect 133 105 134 106
rect 124 105 125 106
rect 123 105 124 106
rect 122 105 123 106
rect 121 105 122 106
rect 120 105 121 106
rect 119 105 120 106
rect 118 105 119 106
rect 117 105 118 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 51 105 52 106
rect 50 105 51 106
rect 49 105 50 106
rect 48 105 49 106
rect 47 105 48 106
rect 46 105 47 106
rect 45 105 46 106
rect 44 105 45 106
rect 28 105 29 106
rect 27 105 28 106
rect 26 105 27 106
rect 25 105 26 106
rect 24 105 25 106
rect 23 105 24 106
rect 22 105 23 106
rect 21 105 22 106
rect 20 105 21 106
rect 19 105 20 106
rect 18 105 19 106
rect 17 105 18 106
rect 16 105 17 106
rect 15 105 16 106
rect 14 105 15 106
rect 142 106 143 107
rect 141 106 142 107
rect 140 106 141 107
rect 139 106 140 107
rect 138 106 139 107
rect 137 106 138 107
rect 136 106 137 107
rect 135 106 136 107
rect 134 106 135 107
rect 133 106 134 107
rect 132 106 133 107
rect 131 106 132 107
rect 130 106 131 107
rect 129 106 130 107
rect 128 106 129 107
rect 127 106 128 107
rect 126 106 127 107
rect 125 106 126 107
rect 124 106 125 107
rect 123 106 124 107
rect 122 106 123 107
rect 121 106 122 107
rect 120 106 121 107
rect 119 106 120 107
rect 118 106 119 107
rect 117 106 118 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 51 106 52 107
rect 50 106 51 107
rect 49 106 50 107
rect 48 106 49 107
rect 47 106 48 107
rect 46 106 47 107
rect 45 106 46 107
rect 44 106 45 107
rect 29 106 30 107
rect 28 106 29 107
rect 27 106 28 107
rect 26 106 27 107
rect 25 106 26 107
rect 24 106 25 107
rect 23 106 24 107
rect 22 106 23 107
rect 21 106 22 107
rect 20 106 21 107
rect 19 106 20 107
rect 18 106 19 107
rect 17 106 18 107
rect 16 106 17 107
rect 15 106 16 107
rect 14 106 15 107
rect 142 107 143 108
rect 141 107 142 108
rect 140 107 141 108
rect 139 107 140 108
rect 138 107 139 108
rect 137 107 138 108
rect 136 107 137 108
rect 135 107 136 108
rect 134 107 135 108
rect 133 107 134 108
rect 132 107 133 108
rect 131 107 132 108
rect 130 107 131 108
rect 129 107 130 108
rect 128 107 129 108
rect 127 107 128 108
rect 126 107 127 108
rect 125 107 126 108
rect 124 107 125 108
rect 123 107 124 108
rect 122 107 123 108
rect 121 107 122 108
rect 120 107 121 108
rect 119 107 120 108
rect 118 107 119 108
rect 117 107 118 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 51 107 52 108
rect 50 107 51 108
rect 49 107 50 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 45 107 46 108
rect 44 107 45 108
rect 43 107 44 108
rect 29 107 30 108
rect 28 107 29 108
rect 27 107 28 108
rect 26 107 27 108
rect 25 107 26 108
rect 24 107 25 108
rect 23 107 24 108
rect 22 107 23 108
rect 21 107 22 108
rect 20 107 21 108
rect 19 107 20 108
rect 18 107 19 108
rect 17 107 18 108
rect 16 107 17 108
rect 15 107 16 108
rect 14 107 15 108
rect 142 108 143 109
rect 141 108 142 109
rect 140 108 141 109
rect 139 108 140 109
rect 138 108 139 109
rect 137 108 138 109
rect 136 108 137 109
rect 135 108 136 109
rect 134 108 135 109
rect 133 108 134 109
rect 132 108 133 109
rect 131 108 132 109
rect 130 108 131 109
rect 129 108 130 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 125 108 126 109
rect 124 108 125 109
rect 123 108 124 109
rect 122 108 123 109
rect 121 108 122 109
rect 120 108 121 109
rect 119 108 120 109
rect 118 108 119 109
rect 117 108 118 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 51 108 52 109
rect 50 108 51 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 45 108 46 109
rect 44 108 45 109
rect 43 108 44 109
rect 42 108 43 109
rect 31 108 32 109
rect 30 108 31 109
rect 29 108 30 109
rect 28 108 29 109
rect 27 108 28 109
rect 26 108 27 109
rect 25 108 26 109
rect 24 108 25 109
rect 23 108 24 109
rect 22 108 23 109
rect 21 108 22 109
rect 20 108 21 109
rect 19 108 20 109
rect 18 108 19 109
rect 17 108 18 109
rect 16 108 17 109
rect 15 108 16 109
rect 14 108 15 109
rect 142 109 143 110
rect 141 109 142 110
rect 140 109 141 110
rect 139 109 140 110
rect 138 109 139 110
rect 137 109 138 110
rect 136 109 137 110
rect 135 109 136 110
rect 134 109 135 110
rect 133 109 134 110
rect 132 109 133 110
rect 131 109 132 110
rect 130 109 131 110
rect 129 109 130 110
rect 128 109 129 110
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 124 109 125 110
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 120 109 121 110
rect 119 109 120 110
rect 118 109 119 110
rect 117 109 118 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 52 109 53 110
rect 51 109 52 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 44 109 45 110
rect 43 109 44 110
rect 42 109 43 110
rect 41 109 42 110
rect 40 109 41 110
rect 39 109 40 110
rect 33 109 34 110
rect 32 109 33 110
rect 31 109 32 110
rect 30 109 31 110
rect 29 109 30 110
rect 28 109 29 110
rect 27 109 28 110
rect 26 109 27 110
rect 25 109 26 110
rect 24 109 25 110
rect 23 109 24 110
rect 22 109 23 110
rect 21 109 22 110
rect 20 109 21 110
rect 19 109 20 110
rect 18 109 19 110
rect 17 109 18 110
rect 16 109 17 110
rect 15 109 16 110
rect 14 109 15 110
rect 142 110 143 111
rect 141 110 142 111
rect 140 110 141 111
rect 139 110 140 111
rect 138 110 139 111
rect 137 110 138 111
rect 136 110 137 111
rect 135 110 136 111
rect 134 110 135 111
rect 133 110 134 111
rect 132 110 133 111
rect 131 110 132 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 127 110 128 111
rect 126 110 127 111
rect 125 110 126 111
rect 124 110 125 111
rect 123 110 124 111
rect 122 110 123 111
rect 121 110 122 111
rect 120 110 121 111
rect 119 110 120 111
rect 118 110 119 111
rect 117 110 118 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 52 110 53 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 43 110 44 111
rect 42 110 43 111
rect 41 110 42 111
rect 40 110 41 111
rect 39 110 40 111
rect 38 110 39 111
rect 37 110 38 111
rect 36 110 37 111
rect 35 110 36 111
rect 34 110 35 111
rect 33 110 34 111
rect 32 110 33 111
rect 31 110 32 111
rect 30 110 31 111
rect 29 110 30 111
rect 28 110 29 111
rect 27 110 28 111
rect 26 110 27 111
rect 25 110 26 111
rect 24 110 25 111
rect 23 110 24 111
rect 22 110 23 111
rect 21 110 22 111
rect 20 110 21 111
rect 19 110 20 111
rect 18 110 19 111
rect 17 110 18 111
rect 16 110 17 111
rect 15 110 16 111
rect 14 110 15 111
rect 137 111 138 112
rect 136 111 137 112
rect 135 111 136 112
rect 134 111 135 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 52 111 53 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 40 111 41 112
rect 39 111 40 112
rect 38 111 39 112
rect 37 111 38 112
rect 36 111 37 112
rect 35 111 36 112
rect 34 111 35 112
rect 33 111 34 112
rect 32 111 33 112
rect 31 111 32 112
rect 30 111 31 112
rect 29 111 30 112
rect 28 111 29 112
rect 27 111 28 112
rect 26 111 27 112
rect 25 111 26 112
rect 24 111 25 112
rect 23 111 24 112
rect 22 111 23 112
rect 21 111 22 112
rect 20 111 21 112
rect 19 111 20 112
rect 18 111 19 112
rect 17 111 18 112
rect 16 111 17 112
rect 15 111 16 112
rect 137 112 138 113
rect 136 112 137 113
rect 135 112 136 113
rect 134 112 135 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 53 112 54 113
rect 52 112 53 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 35 112 36 113
rect 34 112 35 113
rect 33 112 34 113
rect 32 112 33 113
rect 31 112 32 113
rect 30 112 31 113
rect 29 112 30 113
rect 28 112 29 113
rect 27 112 28 113
rect 26 112 27 113
rect 25 112 26 113
rect 24 112 25 113
rect 23 112 24 113
rect 22 112 23 113
rect 21 112 22 113
rect 20 112 21 113
rect 19 112 20 113
rect 18 112 19 113
rect 17 112 18 113
rect 16 112 17 113
rect 15 112 16 113
rect 137 113 138 114
rect 136 113 137 114
rect 135 113 136 114
rect 134 113 135 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 53 113 54 114
rect 52 113 53 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 35 113 36 114
rect 34 113 35 114
rect 33 113 34 114
rect 32 113 33 114
rect 31 113 32 114
rect 30 113 31 114
rect 29 113 30 114
rect 28 113 29 114
rect 27 113 28 114
rect 26 113 27 114
rect 25 113 26 114
rect 24 113 25 114
rect 23 113 24 114
rect 22 113 23 114
rect 21 113 22 114
rect 20 113 21 114
rect 19 113 20 114
rect 18 113 19 114
rect 17 113 18 114
rect 16 113 17 114
rect 15 113 16 114
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 53 114 54 115
rect 52 114 53 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 35 114 36 115
rect 34 114 35 115
rect 33 114 34 115
rect 32 114 33 115
rect 31 114 32 115
rect 30 114 31 115
rect 29 114 30 115
rect 28 114 29 115
rect 27 114 28 115
rect 26 114 27 115
rect 25 114 26 115
rect 24 114 25 115
rect 23 114 24 115
rect 22 114 23 115
rect 21 114 22 115
rect 20 114 21 115
rect 19 114 20 115
rect 18 114 19 115
rect 17 114 18 115
rect 16 114 17 115
rect 15 114 16 115
rect 56 115 57 116
rect 55 115 56 116
rect 54 115 55 116
rect 53 115 54 116
rect 52 115 53 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 35 115 36 116
rect 34 115 35 116
rect 33 115 34 116
rect 32 115 33 116
rect 31 115 32 116
rect 30 115 31 116
rect 29 115 30 116
rect 28 115 29 116
rect 27 115 28 116
rect 26 115 27 116
rect 25 115 26 116
rect 24 115 25 116
rect 23 115 24 116
rect 22 115 23 116
rect 21 115 22 116
rect 20 115 21 116
rect 19 115 20 116
rect 18 115 19 116
rect 17 115 18 116
rect 16 115 17 116
rect 15 115 16 116
rect 147 116 148 117
rect 146 116 147 117
rect 145 116 146 117
rect 144 116 145 117
rect 56 116 57 117
rect 55 116 56 117
rect 54 116 55 117
rect 53 116 54 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 34 116 35 117
rect 33 116 34 117
rect 32 116 33 117
rect 31 116 32 117
rect 30 116 31 117
rect 29 116 30 117
rect 28 116 29 117
rect 27 116 28 117
rect 26 116 27 117
rect 25 116 26 117
rect 24 116 25 117
rect 23 116 24 117
rect 22 116 23 117
rect 21 116 22 117
rect 20 116 21 117
rect 19 116 20 117
rect 18 116 19 117
rect 17 116 18 117
rect 16 116 17 117
rect 15 116 16 117
rect 147 117 148 118
rect 146 117 147 118
rect 145 117 146 118
rect 144 117 145 118
rect 143 117 144 118
rect 142 117 143 118
rect 141 117 142 118
rect 140 117 141 118
rect 139 117 140 118
rect 55 117 56 118
rect 54 117 55 118
rect 53 117 54 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 35 117 36 118
rect 34 117 35 118
rect 33 117 34 118
rect 32 117 33 118
rect 31 117 32 118
rect 30 117 31 118
rect 29 117 30 118
rect 28 117 29 118
rect 27 117 28 118
rect 26 117 27 118
rect 25 117 26 118
rect 24 117 25 118
rect 23 117 24 118
rect 22 117 23 118
rect 21 117 22 118
rect 20 117 21 118
rect 19 117 20 118
rect 18 117 19 118
rect 17 117 18 118
rect 16 117 17 118
rect 147 118 148 119
rect 146 118 147 119
rect 145 118 146 119
rect 144 118 145 119
rect 143 118 144 119
rect 142 118 143 119
rect 141 118 142 119
rect 140 118 141 119
rect 139 118 140 119
rect 55 118 56 119
rect 54 118 55 119
rect 53 118 54 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 35 118 36 119
rect 34 118 35 119
rect 33 118 34 119
rect 32 118 33 119
rect 31 118 32 119
rect 30 118 31 119
rect 29 118 30 119
rect 28 118 29 119
rect 27 118 28 119
rect 26 118 27 119
rect 25 118 26 119
rect 24 118 25 119
rect 23 118 24 119
rect 22 118 23 119
rect 21 118 22 119
rect 20 118 21 119
rect 19 118 20 119
rect 18 118 19 119
rect 17 118 18 119
rect 16 118 17 119
rect 147 119 148 120
rect 146 119 147 120
rect 145 119 146 120
rect 144 119 145 120
rect 143 119 144 120
rect 142 119 143 120
rect 141 119 142 120
rect 140 119 141 120
rect 139 119 140 120
rect 54 119 55 120
rect 53 119 54 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 35 119 36 120
rect 34 119 35 120
rect 33 119 34 120
rect 32 119 33 120
rect 31 119 32 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 27 119 28 120
rect 26 119 27 120
rect 25 119 26 120
rect 24 119 25 120
rect 23 119 24 120
rect 22 119 23 120
rect 21 119 22 120
rect 20 119 21 120
rect 19 119 20 120
rect 18 119 19 120
rect 17 119 18 120
rect 16 119 17 120
rect 145 120 146 121
rect 144 120 145 121
rect 143 120 144 121
rect 142 120 143 121
rect 141 120 142 121
rect 140 120 141 121
rect 139 120 140 121
rect 54 120 55 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 35 120 36 121
rect 34 120 35 121
rect 33 120 34 121
rect 32 120 33 121
rect 31 120 32 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 26 120 27 121
rect 25 120 26 121
rect 24 120 25 121
rect 23 120 24 121
rect 22 120 23 121
rect 21 120 22 121
rect 20 120 21 121
rect 19 120 20 121
rect 18 120 19 121
rect 17 120 18 121
rect 142 121 143 122
rect 141 121 142 122
rect 140 121 141 122
rect 139 121 140 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 36 121 37 122
rect 35 121 36 122
rect 34 121 35 122
rect 33 121 34 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 26 121 27 122
rect 25 121 26 122
rect 24 121 25 122
rect 23 121 24 122
rect 22 121 23 122
rect 21 121 22 122
rect 20 121 21 122
rect 19 121 20 122
rect 18 121 19 122
rect 17 121 18 122
rect 139 122 140 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 36 122 37 123
rect 35 122 36 123
rect 34 122 35 123
rect 33 122 34 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 26 122 27 123
rect 25 122 26 123
rect 24 122 25 123
rect 23 122 24 123
rect 22 122 23 123
rect 21 122 22 123
rect 20 122 21 123
rect 19 122 20 123
rect 18 122 19 123
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 36 123 37 124
rect 35 123 36 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 26 123 27 124
rect 25 123 26 124
rect 24 123 25 124
rect 23 123 24 124
rect 22 123 23 124
rect 21 123 22 124
rect 20 123 21 124
rect 19 123 20 124
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 36 124 37 125
rect 35 124 36 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 26 124 27 125
rect 25 124 26 125
rect 24 124 25 125
rect 23 124 24 125
rect 22 124 23 125
rect 21 124 22 125
rect 20 124 21 125
rect 19 124 20 125
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 37 125 38 126
rect 36 125 37 126
rect 35 125 36 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 27 125 28 126
rect 26 125 27 126
rect 25 125 26 126
rect 24 125 25 126
rect 23 125 24 126
rect 22 125 23 126
rect 21 125 22 126
rect 20 125 21 126
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 37 126 38 127
rect 36 126 37 127
rect 35 126 36 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 27 126 28 127
rect 26 126 27 127
rect 25 126 26 127
rect 24 126 25 127
rect 23 126 24 127
rect 22 126 23 127
rect 21 126 22 127
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 38 127 39 128
rect 37 127 38 128
rect 36 127 37 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 27 127 28 128
rect 26 127 27 128
rect 25 127 26 128
rect 24 127 25 128
rect 23 127 24 128
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 38 128 39 129
rect 37 128 38 129
rect 36 128 37 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 28 128 29 129
rect 27 128 28 129
rect 26 128 27 129
rect 25 128 26 129
rect 24 128 25 129
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 39 129 40 130
rect 38 129 39 130
rect 37 129 38 130
rect 36 129 37 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 28 129 29 130
rect 27 129 28 130
rect 26 129 27 130
rect 40 130 41 131
rect 39 130 40 131
rect 38 130 39 131
rect 37 130 38 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 142 136 143 137
rect 141 136 142 137
rect 140 136 141 137
rect 139 136 140 137
rect 138 136 139 137
rect 137 136 138 137
rect 142 137 143 138
rect 141 137 142 138
rect 140 137 141 138
rect 139 137 140 138
rect 138 137 139 138
rect 142 138 143 139
rect 141 138 142 139
rect 140 138 141 139
rect 139 138 140 139
rect 138 138 139 139
rect 50 138 51 139
rect 49 138 50 139
rect 48 138 49 139
rect 47 138 48 139
rect 46 138 47 139
rect 45 138 46 139
rect 44 138 45 139
rect 43 138 44 139
rect 42 138 43 139
rect 41 138 42 139
rect 40 138 41 139
rect 39 138 40 139
rect 38 138 39 139
rect 37 138 38 139
rect 36 138 37 139
rect 35 138 36 139
rect 34 138 35 139
rect 33 138 34 139
rect 32 138 33 139
rect 31 138 32 139
rect 30 138 31 139
rect 29 138 30 139
rect 28 138 29 139
rect 27 138 28 139
rect 26 138 27 139
rect 25 138 26 139
rect 24 138 25 139
rect 23 138 24 139
rect 22 138 23 139
rect 21 138 22 139
rect 20 138 21 139
rect 19 138 20 139
rect 18 138 19 139
rect 17 138 18 139
rect 16 138 17 139
rect 15 138 16 139
rect 14 138 15 139
rect 142 139 143 140
rect 141 139 142 140
rect 140 139 141 140
rect 139 139 140 140
rect 138 139 139 140
rect 61 139 62 140
rect 60 139 61 140
rect 59 139 60 140
rect 58 139 59 140
rect 57 139 58 140
rect 56 139 57 140
rect 55 139 56 140
rect 54 139 55 140
rect 53 139 54 140
rect 52 139 53 140
rect 51 139 52 140
rect 50 139 51 140
rect 49 139 50 140
rect 48 139 49 140
rect 47 139 48 140
rect 46 139 47 140
rect 45 139 46 140
rect 44 139 45 140
rect 43 139 44 140
rect 42 139 43 140
rect 41 139 42 140
rect 40 139 41 140
rect 39 139 40 140
rect 38 139 39 140
rect 37 139 38 140
rect 36 139 37 140
rect 35 139 36 140
rect 34 139 35 140
rect 33 139 34 140
rect 32 139 33 140
rect 31 139 32 140
rect 30 139 31 140
rect 29 139 30 140
rect 28 139 29 140
rect 27 139 28 140
rect 26 139 27 140
rect 25 139 26 140
rect 24 139 25 140
rect 23 139 24 140
rect 22 139 23 140
rect 21 139 22 140
rect 20 139 21 140
rect 19 139 20 140
rect 18 139 19 140
rect 17 139 18 140
rect 16 139 17 140
rect 15 139 16 140
rect 14 139 15 140
rect 142 140 143 141
rect 141 140 142 141
rect 140 140 141 141
rect 139 140 140 141
rect 138 140 139 141
rect 64 140 65 141
rect 63 140 64 141
rect 62 140 63 141
rect 61 140 62 141
rect 60 140 61 141
rect 59 140 60 141
rect 58 140 59 141
rect 57 140 58 141
rect 56 140 57 141
rect 55 140 56 141
rect 54 140 55 141
rect 53 140 54 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 48 140 49 141
rect 47 140 48 141
rect 46 140 47 141
rect 45 140 46 141
rect 44 140 45 141
rect 43 140 44 141
rect 42 140 43 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 37 140 38 141
rect 36 140 37 141
rect 35 140 36 141
rect 34 140 35 141
rect 33 140 34 141
rect 32 140 33 141
rect 31 140 32 141
rect 30 140 31 141
rect 29 140 30 141
rect 28 140 29 141
rect 27 140 28 141
rect 26 140 27 141
rect 25 140 26 141
rect 24 140 25 141
rect 23 140 24 141
rect 22 140 23 141
rect 21 140 22 141
rect 20 140 21 141
rect 19 140 20 141
rect 18 140 19 141
rect 17 140 18 141
rect 16 140 17 141
rect 15 140 16 141
rect 14 140 15 141
rect 142 141 143 142
rect 141 141 142 142
rect 140 141 141 142
rect 139 141 140 142
rect 138 141 139 142
rect 137 141 138 142
rect 67 141 68 142
rect 66 141 67 142
rect 65 141 66 142
rect 64 141 65 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 49 141 50 142
rect 48 141 49 142
rect 47 141 48 142
rect 46 141 47 142
rect 45 141 46 142
rect 44 141 45 142
rect 43 141 44 142
rect 42 141 43 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 38 141 39 142
rect 37 141 38 142
rect 36 141 37 142
rect 35 141 36 142
rect 34 141 35 142
rect 33 141 34 142
rect 32 141 33 142
rect 31 141 32 142
rect 30 141 31 142
rect 29 141 30 142
rect 28 141 29 142
rect 27 141 28 142
rect 26 141 27 142
rect 25 141 26 142
rect 24 141 25 142
rect 23 141 24 142
rect 22 141 23 142
rect 21 141 22 142
rect 20 141 21 142
rect 19 141 20 142
rect 18 141 19 142
rect 17 141 18 142
rect 16 141 17 142
rect 15 141 16 142
rect 14 141 15 142
rect 142 142 143 143
rect 141 142 142 143
rect 140 142 141 143
rect 139 142 140 143
rect 138 142 139 143
rect 137 142 138 143
rect 136 142 137 143
rect 69 142 70 143
rect 68 142 69 143
rect 67 142 68 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 50 142 51 143
rect 49 142 50 143
rect 48 142 49 143
rect 47 142 48 143
rect 46 142 47 143
rect 45 142 46 143
rect 44 142 45 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 37 142 38 143
rect 36 142 37 143
rect 35 142 36 143
rect 34 142 35 143
rect 33 142 34 143
rect 32 142 33 143
rect 31 142 32 143
rect 30 142 31 143
rect 29 142 30 143
rect 28 142 29 143
rect 27 142 28 143
rect 26 142 27 143
rect 25 142 26 143
rect 24 142 25 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 19 142 20 143
rect 18 142 19 143
rect 17 142 18 143
rect 16 142 17 143
rect 15 142 16 143
rect 14 142 15 143
rect 141 143 142 144
rect 140 143 141 144
rect 139 143 140 144
rect 138 143 139 144
rect 137 143 138 144
rect 136 143 137 144
rect 135 143 136 144
rect 134 143 135 144
rect 133 143 134 144
rect 132 143 133 144
rect 131 143 132 144
rect 130 143 131 144
rect 129 143 130 144
rect 128 143 129 144
rect 127 143 128 144
rect 126 143 127 144
rect 125 143 126 144
rect 124 143 125 144
rect 123 143 124 144
rect 122 143 123 144
rect 121 143 122 144
rect 120 143 121 144
rect 119 143 120 144
rect 118 143 119 144
rect 117 143 118 144
rect 70 143 71 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 51 143 52 144
rect 50 143 51 144
rect 49 143 50 144
rect 48 143 49 144
rect 47 143 48 144
rect 46 143 47 144
rect 45 143 46 144
rect 44 143 45 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 37 143 38 144
rect 36 143 37 144
rect 35 143 36 144
rect 34 143 35 144
rect 33 143 34 144
rect 32 143 33 144
rect 31 143 32 144
rect 30 143 31 144
rect 29 143 30 144
rect 28 143 29 144
rect 27 143 28 144
rect 26 143 27 144
rect 25 143 26 144
rect 24 143 25 144
rect 23 143 24 144
rect 22 143 23 144
rect 21 143 22 144
rect 20 143 21 144
rect 19 143 20 144
rect 18 143 19 144
rect 17 143 18 144
rect 16 143 17 144
rect 15 143 16 144
rect 14 143 15 144
rect 141 144 142 145
rect 140 144 141 145
rect 139 144 140 145
rect 138 144 139 145
rect 137 144 138 145
rect 136 144 137 145
rect 135 144 136 145
rect 134 144 135 145
rect 133 144 134 145
rect 132 144 133 145
rect 131 144 132 145
rect 130 144 131 145
rect 129 144 130 145
rect 128 144 129 145
rect 127 144 128 145
rect 126 144 127 145
rect 125 144 126 145
rect 124 144 125 145
rect 123 144 124 145
rect 122 144 123 145
rect 121 144 122 145
rect 120 144 121 145
rect 119 144 120 145
rect 118 144 119 145
rect 117 144 118 145
rect 72 144 73 145
rect 71 144 72 145
rect 70 144 71 145
rect 69 144 70 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 52 144 53 145
rect 51 144 52 145
rect 50 144 51 145
rect 49 144 50 145
rect 48 144 49 145
rect 47 144 48 145
rect 46 144 47 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 37 144 38 145
rect 36 144 37 145
rect 35 144 36 145
rect 34 144 35 145
rect 33 144 34 145
rect 32 144 33 145
rect 31 144 32 145
rect 30 144 31 145
rect 29 144 30 145
rect 28 144 29 145
rect 27 144 28 145
rect 26 144 27 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 21 144 22 145
rect 20 144 21 145
rect 19 144 20 145
rect 18 144 19 145
rect 17 144 18 145
rect 16 144 17 145
rect 15 144 16 145
rect 14 144 15 145
rect 140 145 141 146
rect 139 145 140 146
rect 138 145 139 146
rect 137 145 138 146
rect 136 145 137 146
rect 135 145 136 146
rect 134 145 135 146
rect 133 145 134 146
rect 132 145 133 146
rect 131 145 132 146
rect 130 145 131 146
rect 129 145 130 146
rect 128 145 129 146
rect 127 145 128 146
rect 126 145 127 146
rect 125 145 126 146
rect 124 145 125 146
rect 123 145 124 146
rect 122 145 123 146
rect 121 145 122 146
rect 120 145 121 146
rect 119 145 120 146
rect 118 145 119 146
rect 117 145 118 146
rect 73 145 74 146
rect 72 145 73 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 54 145 55 146
rect 53 145 54 146
rect 52 145 53 146
rect 51 145 52 146
rect 50 145 51 146
rect 49 145 50 146
rect 48 145 49 146
rect 47 145 48 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 37 145 38 146
rect 36 145 37 146
rect 35 145 36 146
rect 34 145 35 146
rect 33 145 34 146
rect 32 145 33 146
rect 31 145 32 146
rect 30 145 31 146
rect 29 145 30 146
rect 28 145 29 146
rect 27 145 28 146
rect 26 145 27 146
rect 25 145 26 146
rect 24 145 25 146
rect 23 145 24 146
rect 22 145 23 146
rect 21 145 22 146
rect 20 145 21 146
rect 19 145 20 146
rect 18 145 19 146
rect 17 145 18 146
rect 16 145 17 146
rect 15 145 16 146
rect 14 145 15 146
rect 139 146 140 147
rect 138 146 139 147
rect 137 146 138 147
rect 136 146 137 147
rect 135 146 136 147
rect 134 146 135 147
rect 133 146 134 147
rect 132 146 133 147
rect 131 146 132 147
rect 130 146 131 147
rect 129 146 130 147
rect 128 146 129 147
rect 127 146 128 147
rect 126 146 127 147
rect 125 146 126 147
rect 124 146 125 147
rect 123 146 124 147
rect 122 146 123 147
rect 121 146 122 147
rect 120 146 121 147
rect 119 146 120 147
rect 118 146 119 147
rect 117 146 118 147
rect 74 146 75 147
rect 73 146 74 147
rect 72 146 73 147
rect 71 146 72 147
rect 70 146 71 147
rect 69 146 70 147
rect 68 146 69 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 57 146 58 147
rect 56 146 57 147
rect 55 146 56 147
rect 54 146 55 147
rect 53 146 54 147
rect 52 146 53 147
rect 51 146 52 147
rect 50 146 51 147
rect 49 146 50 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 37 146 38 147
rect 36 146 37 147
rect 35 146 36 147
rect 34 146 35 147
rect 33 146 34 147
rect 32 146 33 147
rect 31 146 32 147
rect 30 146 31 147
rect 29 146 30 147
rect 28 146 29 147
rect 27 146 28 147
rect 26 146 27 147
rect 25 146 26 147
rect 24 146 25 147
rect 23 146 24 147
rect 22 146 23 147
rect 21 146 22 147
rect 20 146 21 147
rect 19 146 20 147
rect 18 146 19 147
rect 17 146 18 147
rect 16 146 17 147
rect 15 146 16 147
rect 14 146 15 147
rect 138 147 139 148
rect 137 147 138 148
rect 136 147 137 148
rect 135 147 136 148
rect 134 147 135 148
rect 133 147 134 148
rect 132 147 133 148
rect 131 147 132 148
rect 130 147 131 148
rect 129 147 130 148
rect 128 147 129 148
rect 127 147 128 148
rect 126 147 127 148
rect 125 147 126 148
rect 124 147 125 148
rect 123 147 124 148
rect 122 147 123 148
rect 121 147 122 148
rect 120 147 121 148
rect 119 147 120 148
rect 118 147 119 148
rect 117 147 118 148
rect 75 147 76 148
rect 74 147 75 148
rect 73 147 74 148
rect 72 147 73 148
rect 71 147 72 148
rect 70 147 71 148
rect 69 147 70 148
rect 68 147 69 148
rect 67 147 68 148
rect 66 147 67 148
rect 65 147 66 148
rect 64 147 65 148
rect 63 147 64 148
rect 62 147 63 148
rect 61 147 62 148
rect 60 147 61 148
rect 59 147 60 148
rect 58 147 59 148
rect 57 147 58 148
rect 56 147 57 148
rect 55 147 56 148
rect 54 147 55 148
rect 53 147 54 148
rect 52 147 53 148
rect 51 147 52 148
rect 50 147 51 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 36 147 37 148
rect 35 147 36 148
rect 34 147 35 148
rect 33 147 34 148
rect 32 147 33 148
rect 31 147 32 148
rect 30 147 31 148
rect 29 147 30 148
rect 28 147 29 148
rect 27 147 28 148
rect 26 147 27 148
rect 25 147 26 148
rect 24 147 25 148
rect 23 147 24 148
rect 22 147 23 148
rect 21 147 22 148
rect 20 147 21 148
rect 19 147 20 148
rect 18 147 19 148
rect 17 147 18 148
rect 16 147 17 148
rect 15 147 16 148
rect 14 147 15 148
rect 135 148 136 149
rect 134 148 135 149
rect 133 148 134 149
rect 132 148 133 149
rect 131 148 132 149
rect 130 148 131 149
rect 129 148 130 149
rect 128 148 129 149
rect 127 148 128 149
rect 126 148 127 149
rect 125 148 126 149
rect 124 148 125 149
rect 123 148 124 149
rect 122 148 123 149
rect 121 148 122 149
rect 120 148 121 149
rect 119 148 120 149
rect 118 148 119 149
rect 117 148 118 149
rect 76 148 77 149
rect 75 148 76 149
rect 74 148 75 149
rect 73 148 74 149
rect 72 148 73 149
rect 71 148 72 149
rect 70 148 71 149
rect 69 148 70 149
rect 68 148 69 149
rect 67 148 68 149
rect 66 148 67 149
rect 65 148 66 149
rect 64 148 65 149
rect 63 148 64 149
rect 62 148 63 149
rect 61 148 62 149
rect 60 148 61 149
rect 59 148 60 149
rect 58 148 59 149
rect 57 148 58 149
rect 56 148 57 149
rect 55 148 56 149
rect 54 148 55 149
rect 53 148 54 149
rect 52 148 53 149
rect 51 148 52 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 36 148 37 149
rect 35 148 36 149
rect 34 148 35 149
rect 33 148 34 149
rect 32 148 33 149
rect 31 148 32 149
rect 30 148 31 149
rect 29 148 30 149
rect 28 148 29 149
rect 27 148 28 149
rect 26 148 27 149
rect 25 148 26 149
rect 24 148 25 149
rect 23 148 24 149
rect 22 148 23 149
rect 21 148 22 149
rect 20 148 21 149
rect 19 148 20 149
rect 18 148 19 149
rect 17 148 18 149
rect 16 148 17 149
rect 15 148 16 149
rect 14 148 15 149
rect 76 149 77 150
rect 75 149 76 150
rect 74 149 75 150
rect 73 149 74 150
rect 72 149 73 150
rect 71 149 72 150
rect 70 149 71 150
rect 69 149 70 150
rect 68 149 69 150
rect 67 149 68 150
rect 66 149 67 150
rect 65 149 66 150
rect 64 149 65 150
rect 63 149 64 150
rect 62 149 63 150
rect 61 149 62 150
rect 60 149 61 150
rect 59 149 60 150
rect 58 149 59 150
rect 57 149 58 150
rect 56 149 57 150
rect 55 149 56 150
rect 54 149 55 150
rect 53 149 54 150
rect 52 149 53 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 38 149 39 150
rect 37 149 38 150
rect 36 149 37 150
rect 35 149 36 150
rect 34 149 35 150
rect 33 149 34 150
rect 32 149 33 150
rect 31 149 32 150
rect 30 149 31 150
rect 29 149 30 150
rect 28 149 29 150
rect 27 149 28 150
rect 26 149 27 150
rect 25 149 26 150
rect 24 149 25 150
rect 23 149 24 150
rect 22 149 23 150
rect 21 149 22 150
rect 20 149 21 150
rect 19 149 20 150
rect 18 149 19 150
rect 17 149 18 150
rect 16 149 17 150
rect 15 149 16 150
rect 14 149 15 150
rect 77 150 78 151
rect 76 150 77 151
rect 75 150 76 151
rect 74 150 75 151
rect 73 150 74 151
rect 72 150 73 151
rect 71 150 72 151
rect 70 150 71 151
rect 69 150 70 151
rect 68 150 69 151
rect 67 150 68 151
rect 66 150 67 151
rect 65 150 66 151
rect 64 150 65 151
rect 63 150 64 151
rect 62 150 63 151
rect 61 150 62 151
rect 60 150 61 151
rect 59 150 60 151
rect 58 150 59 151
rect 57 150 58 151
rect 56 150 57 151
rect 55 150 56 151
rect 54 150 55 151
rect 53 150 54 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 38 150 39 151
rect 37 150 38 151
rect 36 150 37 151
rect 35 150 36 151
rect 34 150 35 151
rect 33 150 34 151
rect 32 150 33 151
rect 31 150 32 151
rect 30 150 31 151
rect 29 150 30 151
rect 28 150 29 151
rect 27 150 28 151
rect 26 150 27 151
rect 25 150 26 151
rect 24 150 25 151
rect 23 150 24 151
rect 22 150 23 151
rect 21 150 22 151
rect 20 150 21 151
rect 19 150 20 151
rect 18 150 19 151
rect 17 150 18 151
rect 16 150 17 151
rect 15 150 16 151
rect 14 150 15 151
rect 77 151 78 152
rect 76 151 77 152
rect 75 151 76 152
rect 74 151 75 152
rect 73 151 74 152
rect 72 151 73 152
rect 71 151 72 152
rect 70 151 71 152
rect 69 151 70 152
rect 68 151 69 152
rect 67 151 68 152
rect 66 151 67 152
rect 65 151 66 152
rect 64 151 65 152
rect 63 151 64 152
rect 62 151 63 152
rect 61 151 62 152
rect 60 151 61 152
rect 59 151 60 152
rect 58 151 59 152
rect 57 151 58 152
rect 56 151 57 152
rect 55 151 56 152
rect 54 151 55 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 40 151 41 152
rect 39 151 40 152
rect 38 151 39 152
rect 37 151 38 152
rect 36 151 37 152
rect 35 151 36 152
rect 34 151 35 152
rect 33 151 34 152
rect 32 151 33 152
rect 31 151 32 152
rect 30 151 31 152
rect 29 151 30 152
rect 28 151 29 152
rect 27 151 28 152
rect 26 151 27 152
rect 25 151 26 152
rect 24 151 25 152
rect 23 151 24 152
rect 22 151 23 152
rect 21 151 22 152
rect 20 151 21 152
rect 19 151 20 152
rect 18 151 19 152
rect 17 151 18 152
rect 16 151 17 152
rect 15 151 16 152
rect 14 151 15 152
rect 78 152 79 153
rect 77 152 78 153
rect 76 152 77 153
rect 75 152 76 153
rect 74 152 75 153
rect 73 152 74 153
rect 72 152 73 153
rect 71 152 72 153
rect 70 152 71 153
rect 69 152 70 153
rect 68 152 69 153
rect 67 152 68 153
rect 66 152 67 153
rect 65 152 66 153
rect 64 152 65 153
rect 63 152 64 153
rect 62 152 63 153
rect 61 152 62 153
rect 60 152 61 153
rect 59 152 60 153
rect 58 152 59 153
rect 57 152 58 153
rect 56 152 57 153
rect 55 152 56 153
rect 54 152 55 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 40 152 41 153
rect 39 152 40 153
rect 38 152 39 153
rect 37 152 38 153
rect 36 152 37 153
rect 35 152 36 153
rect 34 152 35 153
rect 33 152 34 153
rect 32 152 33 153
rect 31 152 32 153
rect 30 152 31 153
rect 29 152 30 153
rect 28 152 29 153
rect 27 152 28 153
rect 26 152 27 153
rect 25 152 26 153
rect 24 152 25 153
rect 23 152 24 153
rect 22 152 23 153
rect 21 152 22 153
rect 20 152 21 153
rect 19 152 20 153
rect 18 152 19 153
rect 17 152 18 153
rect 16 152 17 153
rect 15 152 16 153
rect 14 152 15 153
rect 139 153 140 154
rect 138 153 139 154
rect 137 153 138 154
rect 136 153 137 154
rect 135 153 136 154
rect 78 153 79 154
rect 77 153 78 154
rect 76 153 77 154
rect 75 153 76 154
rect 74 153 75 154
rect 73 153 74 154
rect 72 153 73 154
rect 71 153 72 154
rect 70 153 71 154
rect 69 153 70 154
rect 68 153 69 154
rect 67 153 68 154
rect 66 153 67 154
rect 65 153 66 154
rect 64 153 65 154
rect 63 153 64 154
rect 62 153 63 154
rect 61 153 62 154
rect 60 153 61 154
rect 59 153 60 154
rect 58 153 59 154
rect 57 153 58 154
rect 56 153 57 154
rect 55 153 56 154
rect 54 153 55 154
rect 53 153 54 154
rect 52 153 53 154
rect 51 153 52 154
rect 50 153 51 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 43 153 44 154
rect 42 153 43 154
rect 41 153 42 154
rect 40 153 41 154
rect 39 153 40 154
rect 38 153 39 154
rect 37 153 38 154
rect 36 153 37 154
rect 35 153 36 154
rect 34 153 35 154
rect 33 153 34 154
rect 32 153 33 154
rect 31 153 32 154
rect 30 153 31 154
rect 29 153 30 154
rect 28 153 29 154
rect 27 153 28 154
rect 26 153 27 154
rect 25 153 26 154
rect 24 153 25 154
rect 23 153 24 154
rect 22 153 23 154
rect 21 153 22 154
rect 20 153 21 154
rect 19 153 20 154
rect 18 153 19 154
rect 17 153 18 154
rect 16 153 17 154
rect 15 153 16 154
rect 14 153 15 154
rect 140 154 141 155
rect 139 154 140 155
rect 138 154 139 155
rect 137 154 138 155
rect 136 154 137 155
rect 135 154 136 155
rect 134 154 135 155
rect 79 154 80 155
rect 78 154 79 155
rect 77 154 78 155
rect 76 154 77 155
rect 75 154 76 155
rect 74 154 75 155
rect 73 154 74 155
rect 72 154 73 155
rect 71 154 72 155
rect 70 154 71 155
rect 69 154 70 155
rect 68 154 69 155
rect 67 154 68 155
rect 66 154 67 155
rect 65 154 66 155
rect 64 154 65 155
rect 63 154 64 155
rect 62 154 63 155
rect 61 154 62 155
rect 60 154 61 155
rect 59 154 60 155
rect 58 154 59 155
rect 57 154 58 155
rect 56 154 57 155
rect 55 154 56 155
rect 54 154 55 155
rect 53 154 54 155
rect 52 154 53 155
rect 51 154 52 155
rect 50 154 51 155
rect 49 154 50 155
rect 48 154 49 155
rect 47 154 48 155
rect 46 154 47 155
rect 45 154 46 155
rect 44 154 45 155
rect 43 154 44 155
rect 42 154 43 155
rect 41 154 42 155
rect 40 154 41 155
rect 39 154 40 155
rect 38 154 39 155
rect 37 154 38 155
rect 36 154 37 155
rect 35 154 36 155
rect 34 154 35 155
rect 33 154 34 155
rect 32 154 33 155
rect 31 154 32 155
rect 30 154 31 155
rect 29 154 30 155
rect 28 154 29 155
rect 27 154 28 155
rect 26 154 27 155
rect 25 154 26 155
rect 24 154 25 155
rect 23 154 24 155
rect 22 154 23 155
rect 21 154 22 155
rect 20 154 21 155
rect 19 154 20 155
rect 18 154 19 155
rect 17 154 18 155
rect 16 154 17 155
rect 15 154 16 155
rect 14 154 15 155
rect 141 155 142 156
rect 140 155 141 156
rect 139 155 140 156
rect 138 155 139 156
rect 137 155 138 156
rect 136 155 137 156
rect 135 155 136 156
rect 134 155 135 156
rect 133 155 134 156
rect 129 155 130 156
rect 128 155 129 156
rect 127 155 128 156
rect 126 155 127 156
rect 125 155 126 156
rect 79 155 80 156
rect 78 155 79 156
rect 77 155 78 156
rect 76 155 77 156
rect 75 155 76 156
rect 74 155 75 156
rect 73 155 74 156
rect 72 155 73 156
rect 71 155 72 156
rect 70 155 71 156
rect 69 155 70 156
rect 68 155 69 156
rect 67 155 68 156
rect 66 155 67 156
rect 65 155 66 156
rect 64 155 65 156
rect 63 155 64 156
rect 62 155 63 156
rect 61 155 62 156
rect 60 155 61 156
rect 59 155 60 156
rect 58 155 59 156
rect 57 155 58 156
rect 56 155 57 156
rect 55 155 56 156
rect 54 155 55 156
rect 53 155 54 156
rect 52 155 53 156
rect 51 155 52 156
rect 50 155 51 156
rect 49 155 50 156
rect 48 155 49 156
rect 47 155 48 156
rect 46 155 47 156
rect 45 155 46 156
rect 44 155 45 156
rect 43 155 44 156
rect 42 155 43 156
rect 41 155 42 156
rect 40 155 41 156
rect 39 155 40 156
rect 38 155 39 156
rect 37 155 38 156
rect 36 155 37 156
rect 35 155 36 156
rect 34 155 35 156
rect 33 155 34 156
rect 32 155 33 156
rect 31 155 32 156
rect 30 155 31 156
rect 29 155 30 156
rect 28 155 29 156
rect 27 155 28 156
rect 26 155 27 156
rect 25 155 26 156
rect 24 155 25 156
rect 23 155 24 156
rect 22 155 23 156
rect 21 155 22 156
rect 20 155 21 156
rect 19 155 20 156
rect 18 155 19 156
rect 17 155 18 156
rect 16 155 17 156
rect 15 155 16 156
rect 14 155 15 156
rect 142 156 143 157
rect 141 156 142 157
rect 140 156 141 157
rect 139 156 140 157
rect 138 156 139 157
rect 137 156 138 157
rect 136 156 137 157
rect 135 156 136 157
rect 134 156 135 157
rect 133 156 134 157
rect 132 156 133 157
rect 128 156 129 157
rect 127 156 128 157
rect 126 156 127 157
rect 125 156 126 157
rect 80 156 81 157
rect 79 156 80 157
rect 78 156 79 157
rect 77 156 78 157
rect 76 156 77 157
rect 75 156 76 157
rect 74 156 75 157
rect 73 156 74 157
rect 72 156 73 157
rect 71 156 72 157
rect 70 156 71 157
rect 69 156 70 157
rect 68 156 69 157
rect 67 156 68 157
rect 66 156 67 157
rect 65 156 66 157
rect 64 156 65 157
rect 63 156 64 157
rect 62 156 63 157
rect 61 156 62 157
rect 60 156 61 157
rect 59 156 60 157
rect 58 156 59 157
rect 57 156 58 157
rect 56 156 57 157
rect 55 156 56 157
rect 54 156 55 157
rect 53 156 54 157
rect 52 156 53 157
rect 51 156 52 157
rect 50 156 51 157
rect 49 156 50 157
rect 48 156 49 157
rect 47 156 48 157
rect 46 156 47 157
rect 45 156 46 157
rect 44 156 45 157
rect 43 156 44 157
rect 42 156 43 157
rect 41 156 42 157
rect 40 156 41 157
rect 39 156 40 157
rect 38 156 39 157
rect 37 156 38 157
rect 36 156 37 157
rect 35 156 36 157
rect 34 156 35 157
rect 33 156 34 157
rect 32 156 33 157
rect 31 156 32 157
rect 30 156 31 157
rect 29 156 30 157
rect 28 156 29 157
rect 27 156 28 157
rect 26 156 27 157
rect 25 156 26 157
rect 24 156 25 157
rect 23 156 24 157
rect 22 156 23 157
rect 21 156 22 157
rect 20 156 21 157
rect 19 156 20 157
rect 18 156 19 157
rect 17 156 18 157
rect 16 156 17 157
rect 15 156 16 157
rect 14 156 15 157
rect 142 157 143 158
rect 141 157 142 158
rect 140 157 141 158
rect 139 157 140 158
rect 138 157 139 158
rect 137 157 138 158
rect 136 157 137 158
rect 135 157 136 158
rect 134 157 135 158
rect 133 157 134 158
rect 132 157 133 158
rect 128 157 129 158
rect 127 157 128 158
rect 126 157 127 158
rect 125 157 126 158
rect 80 157 81 158
rect 79 157 80 158
rect 78 157 79 158
rect 77 157 78 158
rect 76 157 77 158
rect 75 157 76 158
rect 74 157 75 158
rect 73 157 74 158
rect 72 157 73 158
rect 71 157 72 158
rect 70 157 71 158
rect 69 157 70 158
rect 68 157 69 158
rect 67 157 68 158
rect 66 157 67 158
rect 65 157 66 158
rect 64 157 65 158
rect 63 157 64 158
rect 62 157 63 158
rect 61 157 62 158
rect 60 157 61 158
rect 59 157 60 158
rect 58 157 59 158
rect 57 157 58 158
rect 56 157 57 158
rect 55 157 56 158
rect 54 157 55 158
rect 53 157 54 158
rect 52 157 53 158
rect 51 157 52 158
rect 50 157 51 158
rect 49 157 50 158
rect 48 157 49 158
rect 47 157 48 158
rect 46 157 47 158
rect 45 157 46 158
rect 44 157 45 158
rect 43 157 44 158
rect 42 157 43 158
rect 41 157 42 158
rect 40 157 41 158
rect 39 157 40 158
rect 38 157 39 158
rect 37 157 38 158
rect 36 157 37 158
rect 35 157 36 158
rect 34 157 35 158
rect 33 157 34 158
rect 32 157 33 158
rect 31 157 32 158
rect 30 157 31 158
rect 29 157 30 158
rect 28 157 29 158
rect 27 157 28 158
rect 26 157 27 158
rect 25 157 26 158
rect 24 157 25 158
rect 23 157 24 158
rect 22 157 23 158
rect 21 157 22 158
rect 20 157 21 158
rect 19 157 20 158
rect 18 157 19 158
rect 17 157 18 158
rect 16 157 17 158
rect 15 157 16 158
rect 14 157 15 158
rect 142 158 143 159
rect 141 158 142 159
rect 140 158 141 159
rect 139 158 140 159
rect 138 158 139 159
rect 135 158 136 159
rect 134 158 135 159
rect 133 158 134 159
rect 132 158 133 159
rect 127 158 128 159
rect 126 158 127 159
rect 125 158 126 159
rect 124 158 125 159
rect 80 158 81 159
rect 79 158 80 159
rect 78 158 79 159
rect 77 158 78 159
rect 76 158 77 159
rect 75 158 76 159
rect 74 158 75 159
rect 73 158 74 159
rect 72 158 73 159
rect 71 158 72 159
rect 70 158 71 159
rect 69 158 70 159
rect 68 158 69 159
rect 67 158 68 159
rect 66 158 67 159
rect 65 158 66 159
rect 64 158 65 159
rect 63 158 64 159
rect 62 158 63 159
rect 61 158 62 159
rect 60 158 61 159
rect 59 158 60 159
rect 58 158 59 159
rect 57 158 58 159
rect 56 158 57 159
rect 55 158 56 159
rect 54 158 55 159
rect 53 158 54 159
rect 52 158 53 159
rect 51 158 52 159
rect 50 158 51 159
rect 49 158 50 159
rect 48 158 49 159
rect 47 158 48 159
rect 46 158 47 159
rect 45 158 46 159
rect 44 158 45 159
rect 43 158 44 159
rect 42 158 43 159
rect 41 158 42 159
rect 40 158 41 159
rect 39 158 40 159
rect 38 158 39 159
rect 37 158 38 159
rect 36 158 37 159
rect 35 158 36 159
rect 34 158 35 159
rect 33 158 34 159
rect 32 158 33 159
rect 31 158 32 159
rect 30 158 31 159
rect 29 158 30 159
rect 28 158 29 159
rect 27 158 28 159
rect 26 158 27 159
rect 25 158 26 159
rect 24 158 25 159
rect 23 158 24 159
rect 22 158 23 159
rect 21 158 22 159
rect 20 158 21 159
rect 19 158 20 159
rect 18 158 19 159
rect 17 158 18 159
rect 16 158 17 159
rect 15 158 16 159
rect 14 158 15 159
rect 142 159 143 160
rect 141 159 142 160
rect 140 159 141 160
rect 139 159 140 160
rect 134 159 135 160
rect 133 159 134 160
rect 132 159 133 160
rect 131 159 132 160
rect 127 159 128 160
rect 126 159 127 160
rect 125 159 126 160
rect 124 159 125 160
rect 80 159 81 160
rect 79 159 80 160
rect 78 159 79 160
rect 77 159 78 160
rect 76 159 77 160
rect 75 159 76 160
rect 74 159 75 160
rect 73 159 74 160
rect 72 159 73 160
rect 71 159 72 160
rect 70 159 71 160
rect 69 159 70 160
rect 68 159 69 160
rect 67 159 68 160
rect 66 159 67 160
rect 65 159 66 160
rect 64 159 65 160
rect 63 159 64 160
rect 62 159 63 160
rect 61 159 62 160
rect 60 159 61 160
rect 59 159 60 160
rect 58 159 59 160
rect 142 160 143 161
rect 141 160 142 161
rect 140 160 141 161
rect 139 160 140 161
rect 133 160 134 161
rect 132 160 133 161
rect 131 160 132 161
rect 127 160 128 161
rect 126 160 127 161
rect 125 160 126 161
rect 124 160 125 161
rect 80 160 81 161
rect 79 160 80 161
rect 78 160 79 161
rect 77 160 78 161
rect 76 160 77 161
rect 75 160 76 161
rect 74 160 75 161
rect 73 160 74 161
rect 72 160 73 161
rect 71 160 72 161
rect 70 160 71 161
rect 69 160 70 161
rect 68 160 69 161
rect 67 160 68 161
rect 66 160 67 161
rect 65 160 66 161
rect 64 160 65 161
rect 63 160 64 161
rect 62 160 63 161
rect 61 160 62 161
rect 141 161 142 162
rect 140 161 141 162
rect 139 161 140 162
rect 133 161 134 162
rect 132 161 133 162
rect 131 161 132 162
rect 127 161 128 162
rect 126 161 127 162
rect 125 161 126 162
rect 124 161 125 162
rect 81 161 82 162
rect 80 161 81 162
rect 79 161 80 162
rect 78 161 79 162
rect 77 161 78 162
rect 76 161 77 162
rect 75 161 76 162
rect 74 161 75 162
rect 73 161 74 162
rect 72 161 73 162
rect 71 161 72 162
rect 70 161 71 162
rect 69 161 70 162
rect 68 161 69 162
rect 67 161 68 162
rect 66 161 67 162
rect 65 161 66 162
rect 64 161 65 162
rect 63 161 64 162
rect 62 161 63 162
rect 141 162 142 163
rect 140 162 141 163
rect 139 162 140 163
rect 133 162 134 163
rect 132 162 133 163
rect 131 162 132 163
rect 127 162 128 163
rect 126 162 127 163
rect 125 162 126 163
rect 124 162 125 163
rect 81 162 82 163
rect 80 162 81 163
rect 79 162 80 163
rect 78 162 79 163
rect 77 162 78 163
rect 76 162 77 163
rect 75 162 76 163
rect 74 162 75 163
rect 73 162 74 163
rect 72 162 73 163
rect 71 162 72 163
rect 70 162 71 163
rect 69 162 70 163
rect 68 162 69 163
rect 67 162 68 163
rect 66 162 67 163
rect 65 162 66 163
rect 64 162 65 163
rect 63 162 64 163
rect 140 163 141 164
rect 139 163 140 164
rect 138 163 139 164
rect 133 163 134 164
rect 132 163 133 164
rect 131 163 132 164
rect 127 163 128 164
rect 126 163 127 164
rect 125 163 126 164
rect 124 163 125 164
rect 81 163 82 164
rect 80 163 81 164
rect 79 163 80 164
rect 78 163 79 164
rect 77 163 78 164
rect 76 163 77 164
rect 75 163 76 164
rect 74 163 75 164
rect 73 163 74 164
rect 72 163 73 164
rect 71 163 72 164
rect 70 163 71 164
rect 69 163 70 164
rect 68 163 69 164
rect 67 163 68 164
rect 66 163 67 164
rect 65 163 66 164
rect 64 163 65 164
rect 140 164 141 165
rect 139 164 140 165
rect 138 164 139 165
rect 137 164 138 165
rect 136 164 137 165
rect 133 164 134 165
rect 132 164 133 165
rect 131 164 132 165
rect 130 164 131 165
rect 129 164 130 165
rect 128 164 129 165
rect 127 164 128 165
rect 126 164 127 165
rect 125 164 126 165
rect 124 164 125 165
rect 81 164 82 165
rect 80 164 81 165
rect 79 164 80 165
rect 78 164 79 165
rect 77 164 78 165
rect 76 164 77 165
rect 75 164 76 165
rect 74 164 75 165
rect 73 164 74 165
rect 72 164 73 165
rect 71 164 72 165
rect 70 164 71 165
rect 69 164 70 165
rect 68 164 69 165
rect 67 164 68 165
rect 66 164 67 165
rect 65 164 66 165
rect 64 164 65 165
rect 142 165 143 166
rect 141 165 142 166
rect 140 165 141 166
rect 139 165 140 166
rect 138 165 139 166
rect 137 165 138 166
rect 136 165 137 166
rect 135 165 136 166
rect 134 165 135 166
rect 133 165 134 166
rect 132 165 133 166
rect 131 165 132 166
rect 130 165 131 166
rect 129 165 130 166
rect 128 165 129 166
rect 127 165 128 166
rect 126 165 127 166
rect 125 165 126 166
rect 81 165 82 166
rect 80 165 81 166
rect 79 165 80 166
rect 78 165 79 166
rect 77 165 78 166
rect 76 165 77 166
rect 75 165 76 166
rect 74 165 75 166
rect 73 165 74 166
rect 72 165 73 166
rect 71 165 72 166
rect 70 165 71 166
rect 69 165 70 166
rect 68 165 69 166
rect 67 165 68 166
rect 66 165 67 166
rect 65 165 66 166
rect 142 166 143 167
rect 141 166 142 167
rect 140 166 141 167
rect 139 166 140 167
rect 138 166 139 167
rect 137 166 138 167
rect 136 166 137 167
rect 135 166 136 167
rect 134 166 135 167
rect 133 166 134 167
rect 132 166 133 167
rect 131 166 132 167
rect 130 166 131 167
rect 129 166 130 167
rect 128 166 129 167
rect 127 166 128 167
rect 126 166 127 167
rect 125 166 126 167
rect 81 166 82 167
rect 80 166 81 167
rect 79 166 80 167
rect 78 166 79 167
rect 77 166 78 167
rect 76 166 77 167
rect 75 166 76 167
rect 74 166 75 167
rect 73 166 74 167
rect 72 166 73 167
rect 71 166 72 167
rect 70 166 71 167
rect 69 166 70 167
rect 68 166 69 167
rect 67 166 68 167
rect 66 166 67 167
rect 65 166 66 167
rect 142 167 143 168
rect 141 167 142 168
rect 140 167 141 168
rect 139 167 140 168
rect 138 167 139 168
rect 137 167 138 168
rect 136 167 137 168
rect 135 167 136 168
rect 134 167 135 168
rect 133 167 134 168
rect 132 167 133 168
rect 131 167 132 168
rect 130 167 131 168
rect 129 167 130 168
rect 128 167 129 168
rect 127 167 128 168
rect 126 167 127 168
rect 81 167 82 168
rect 80 167 81 168
rect 79 167 80 168
rect 78 167 79 168
rect 77 167 78 168
rect 76 167 77 168
rect 75 167 76 168
rect 74 167 75 168
rect 73 167 74 168
rect 72 167 73 168
rect 71 167 72 168
rect 70 167 71 168
rect 69 167 70 168
rect 68 167 69 168
rect 67 167 68 168
rect 66 167 67 168
rect 65 167 66 168
rect 142 168 143 169
rect 141 168 142 169
rect 140 168 141 169
rect 139 168 140 169
rect 138 168 139 169
rect 137 168 138 169
rect 136 168 137 169
rect 135 168 136 169
rect 134 168 135 169
rect 133 168 134 169
rect 132 168 133 169
rect 131 168 132 169
rect 130 168 131 169
rect 129 168 130 169
rect 128 168 129 169
rect 127 168 128 169
rect 81 168 82 169
rect 80 168 81 169
rect 79 168 80 169
rect 78 168 79 169
rect 77 168 78 169
rect 76 168 77 169
rect 75 168 76 169
rect 74 168 75 169
rect 73 168 74 169
rect 72 168 73 169
rect 71 168 72 169
rect 70 168 71 169
rect 69 168 70 169
rect 68 168 69 169
rect 67 168 68 169
rect 66 168 67 169
rect 65 168 66 169
rect 142 169 143 170
rect 141 169 142 170
rect 140 169 141 170
rect 139 169 140 170
rect 138 169 139 170
rect 137 169 138 170
rect 136 169 137 170
rect 135 169 136 170
rect 134 169 135 170
rect 133 169 134 170
rect 132 169 133 170
rect 131 169 132 170
rect 130 169 131 170
rect 129 169 130 170
rect 81 169 82 170
rect 80 169 81 170
rect 79 169 80 170
rect 78 169 79 170
rect 77 169 78 170
rect 76 169 77 170
rect 75 169 76 170
rect 74 169 75 170
rect 73 169 74 170
rect 72 169 73 170
rect 71 169 72 170
rect 70 169 71 170
rect 69 169 70 170
rect 68 169 69 170
rect 67 169 68 170
rect 66 169 67 170
rect 65 169 66 170
rect 81 170 82 171
rect 80 170 81 171
rect 79 170 80 171
rect 78 170 79 171
rect 77 170 78 171
rect 76 170 77 171
rect 75 170 76 171
rect 74 170 75 171
rect 73 170 74 171
rect 72 170 73 171
rect 71 170 72 171
rect 70 170 71 171
rect 69 170 70 171
rect 68 170 69 171
rect 67 170 68 171
rect 66 170 67 171
rect 65 170 66 171
rect 81 171 82 172
rect 80 171 81 172
rect 79 171 80 172
rect 78 171 79 172
rect 77 171 78 172
rect 76 171 77 172
rect 75 171 76 172
rect 74 171 75 172
rect 73 171 74 172
rect 72 171 73 172
rect 71 171 72 172
rect 70 171 71 172
rect 69 171 70 172
rect 68 171 69 172
rect 67 171 68 172
rect 66 171 67 172
rect 65 171 66 172
rect 64 171 65 172
rect 81 172 82 173
rect 80 172 81 173
rect 79 172 80 173
rect 78 172 79 173
rect 77 172 78 173
rect 76 172 77 173
rect 75 172 76 173
rect 74 172 75 173
rect 73 172 74 173
rect 72 172 73 173
rect 71 172 72 173
rect 70 172 71 173
rect 69 172 70 173
rect 68 172 69 173
rect 67 172 68 173
rect 66 172 67 173
rect 65 172 66 173
rect 64 172 65 173
rect 81 173 82 174
rect 80 173 81 174
rect 79 173 80 174
rect 78 173 79 174
rect 77 173 78 174
rect 76 173 77 174
rect 75 173 76 174
rect 74 173 75 174
rect 73 173 74 174
rect 72 173 73 174
rect 71 173 72 174
rect 70 173 71 174
rect 69 173 70 174
rect 68 173 69 174
rect 67 173 68 174
rect 66 173 67 174
rect 65 173 66 174
rect 64 173 65 174
rect 63 173 64 174
rect 80 174 81 175
rect 79 174 80 175
rect 78 174 79 175
rect 77 174 78 175
rect 76 174 77 175
rect 75 174 76 175
rect 74 174 75 175
rect 73 174 74 175
rect 72 174 73 175
rect 71 174 72 175
rect 70 174 71 175
rect 69 174 70 175
rect 68 174 69 175
rect 67 174 68 175
rect 66 174 67 175
rect 65 174 66 175
rect 64 174 65 175
rect 63 174 64 175
rect 62 174 63 175
rect 142 175 143 176
rect 141 175 142 176
rect 140 175 141 176
rect 139 175 140 176
rect 138 175 139 176
rect 137 175 138 176
rect 136 175 137 176
rect 135 175 136 176
rect 134 175 135 176
rect 133 175 134 176
rect 132 175 133 176
rect 131 175 132 176
rect 130 175 131 176
rect 129 175 130 176
rect 128 175 129 176
rect 127 175 128 176
rect 126 175 127 176
rect 125 175 126 176
rect 124 175 125 176
rect 80 175 81 176
rect 79 175 80 176
rect 78 175 79 176
rect 77 175 78 176
rect 76 175 77 176
rect 75 175 76 176
rect 74 175 75 176
rect 73 175 74 176
rect 72 175 73 176
rect 71 175 72 176
rect 70 175 71 176
rect 69 175 70 176
rect 68 175 69 176
rect 67 175 68 176
rect 66 175 67 176
rect 65 175 66 176
rect 64 175 65 176
rect 63 175 64 176
rect 62 175 63 176
rect 61 175 62 176
rect 142 176 143 177
rect 141 176 142 177
rect 140 176 141 177
rect 139 176 140 177
rect 138 176 139 177
rect 137 176 138 177
rect 136 176 137 177
rect 135 176 136 177
rect 134 176 135 177
rect 133 176 134 177
rect 132 176 133 177
rect 131 176 132 177
rect 130 176 131 177
rect 129 176 130 177
rect 128 176 129 177
rect 127 176 128 177
rect 126 176 127 177
rect 125 176 126 177
rect 124 176 125 177
rect 80 176 81 177
rect 79 176 80 177
rect 78 176 79 177
rect 77 176 78 177
rect 76 176 77 177
rect 75 176 76 177
rect 74 176 75 177
rect 73 176 74 177
rect 72 176 73 177
rect 71 176 72 177
rect 70 176 71 177
rect 69 176 70 177
rect 68 176 69 177
rect 67 176 68 177
rect 66 176 67 177
rect 65 176 66 177
rect 64 176 65 177
rect 63 176 64 177
rect 62 176 63 177
rect 61 176 62 177
rect 60 176 61 177
rect 59 176 60 177
rect 58 176 59 177
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 126 177 127 178
rect 125 177 126 178
rect 124 177 125 178
rect 80 177 81 178
rect 79 177 80 178
rect 78 177 79 178
rect 77 177 78 178
rect 76 177 77 178
rect 75 177 76 178
rect 74 177 75 178
rect 73 177 74 178
rect 72 177 73 178
rect 71 177 72 178
rect 70 177 71 178
rect 69 177 70 178
rect 68 177 69 178
rect 67 177 68 178
rect 66 177 67 178
rect 65 177 66 178
rect 64 177 65 178
rect 63 177 64 178
rect 62 177 63 178
rect 61 177 62 178
rect 60 177 61 178
rect 59 177 60 178
rect 58 177 59 178
rect 57 177 58 178
rect 56 177 57 178
rect 55 177 56 178
rect 54 177 55 178
rect 53 177 54 178
rect 52 177 53 178
rect 51 177 52 178
rect 50 177 51 178
rect 49 177 50 178
rect 48 177 49 178
rect 47 177 48 178
rect 46 177 47 178
rect 45 177 46 178
rect 44 177 45 178
rect 43 177 44 178
rect 42 177 43 178
rect 41 177 42 178
rect 40 177 41 178
rect 39 177 40 178
rect 38 177 39 178
rect 37 177 38 178
rect 36 177 37 178
rect 35 177 36 178
rect 34 177 35 178
rect 33 177 34 178
rect 32 177 33 178
rect 31 177 32 178
rect 30 177 31 178
rect 29 177 30 178
rect 28 177 29 178
rect 27 177 28 178
rect 26 177 27 178
rect 25 177 26 178
rect 24 177 25 178
rect 23 177 24 178
rect 22 177 23 178
rect 21 177 22 178
rect 20 177 21 178
rect 19 177 20 178
rect 18 177 19 178
rect 17 177 18 178
rect 16 177 17 178
rect 15 177 16 178
rect 14 177 15 178
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 125 178 126 179
rect 124 178 125 179
rect 80 178 81 179
rect 79 178 80 179
rect 78 178 79 179
rect 77 178 78 179
rect 76 178 77 179
rect 75 178 76 179
rect 74 178 75 179
rect 73 178 74 179
rect 72 178 73 179
rect 71 178 72 179
rect 70 178 71 179
rect 69 178 70 179
rect 68 178 69 179
rect 67 178 68 179
rect 66 178 67 179
rect 65 178 66 179
rect 64 178 65 179
rect 63 178 64 179
rect 62 178 63 179
rect 61 178 62 179
rect 60 178 61 179
rect 59 178 60 179
rect 58 178 59 179
rect 57 178 58 179
rect 56 178 57 179
rect 55 178 56 179
rect 54 178 55 179
rect 53 178 54 179
rect 52 178 53 179
rect 51 178 52 179
rect 50 178 51 179
rect 49 178 50 179
rect 48 178 49 179
rect 47 178 48 179
rect 46 178 47 179
rect 45 178 46 179
rect 44 178 45 179
rect 43 178 44 179
rect 42 178 43 179
rect 41 178 42 179
rect 40 178 41 179
rect 39 178 40 179
rect 38 178 39 179
rect 37 178 38 179
rect 36 178 37 179
rect 35 178 36 179
rect 34 178 35 179
rect 33 178 34 179
rect 32 178 33 179
rect 31 178 32 179
rect 30 178 31 179
rect 29 178 30 179
rect 28 178 29 179
rect 27 178 28 179
rect 26 178 27 179
rect 25 178 26 179
rect 24 178 25 179
rect 23 178 24 179
rect 22 178 23 179
rect 21 178 22 179
rect 20 178 21 179
rect 19 178 20 179
rect 18 178 19 179
rect 17 178 18 179
rect 16 178 17 179
rect 15 178 16 179
rect 14 178 15 179
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 125 179 126 180
rect 124 179 125 180
rect 79 179 80 180
rect 78 179 79 180
rect 77 179 78 180
rect 76 179 77 180
rect 75 179 76 180
rect 74 179 75 180
rect 73 179 74 180
rect 72 179 73 180
rect 71 179 72 180
rect 70 179 71 180
rect 69 179 70 180
rect 68 179 69 180
rect 67 179 68 180
rect 66 179 67 180
rect 65 179 66 180
rect 64 179 65 180
rect 63 179 64 180
rect 62 179 63 180
rect 61 179 62 180
rect 60 179 61 180
rect 59 179 60 180
rect 58 179 59 180
rect 57 179 58 180
rect 56 179 57 180
rect 55 179 56 180
rect 54 179 55 180
rect 53 179 54 180
rect 52 179 53 180
rect 51 179 52 180
rect 50 179 51 180
rect 49 179 50 180
rect 48 179 49 180
rect 47 179 48 180
rect 46 179 47 180
rect 45 179 46 180
rect 44 179 45 180
rect 43 179 44 180
rect 42 179 43 180
rect 41 179 42 180
rect 40 179 41 180
rect 39 179 40 180
rect 38 179 39 180
rect 37 179 38 180
rect 36 179 37 180
rect 35 179 36 180
rect 34 179 35 180
rect 33 179 34 180
rect 32 179 33 180
rect 31 179 32 180
rect 30 179 31 180
rect 29 179 30 180
rect 28 179 29 180
rect 27 179 28 180
rect 26 179 27 180
rect 25 179 26 180
rect 24 179 25 180
rect 23 179 24 180
rect 22 179 23 180
rect 21 179 22 180
rect 20 179 21 180
rect 19 179 20 180
rect 18 179 19 180
rect 17 179 18 180
rect 16 179 17 180
rect 15 179 16 180
rect 14 179 15 180
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 79 180 80 181
rect 78 180 79 181
rect 77 180 78 181
rect 76 180 77 181
rect 75 180 76 181
rect 74 180 75 181
rect 73 180 74 181
rect 72 180 73 181
rect 71 180 72 181
rect 70 180 71 181
rect 69 180 70 181
rect 68 180 69 181
rect 67 180 68 181
rect 66 180 67 181
rect 65 180 66 181
rect 64 180 65 181
rect 63 180 64 181
rect 62 180 63 181
rect 61 180 62 181
rect 60 180 61 181
rect 59 180 60 181
rect 58 180 59 181
rect 57 180 58 181
rect 56 180 57 181
rect 55 180 56 181
rect 54 180 55 181
rect 53 180 54 181
rect 52 180 53 181
rect 51 180 52 181
rect 50 180 51 181
rect 49 180 50 181
rect 48 180 49 181
rect 47 180 48 181
rect 46 180 47 181
rect 45 180 46 181
rect 44 180 45 181
rect 43 180 44 181
rect 42 180 43 181
rect 41 180 42 181
rect 40 180 41 181
rect 39 180 40 181
rect 38 180 39 181
rect 37 180 38 181
rect 36 180 37 181
rect 35 180 36 181
rect 34 180 35 181
rect 33 180 34 181
rect 32 180 33 181
rect 31 180 32 181
rect 30 180 31 181
rect 29 180 30 181
rect 28 180 29 181
rect 27 180 28 181
rect 26 180 27 181
rect 25 180 26 181
rect 24 180 25 181
rect 23 180 24 181
rect 22 180 23 181
rect 21 180 22 181
rect 20 180 21 181
rect 19 180 20 181
rect 18 180 19 181
rect 17 180 18 181
rect 16 180 17 181
rect 15 180 16 181
rect 14 180 15 181
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 79 181 80 182
rect 78 181 79 182
rect 77 181 78 182
rect 76 181 77 182
rect 75 181 76 182
rect 74 181 75 182
rect 73 181 74 182
rect 72 181 73 182
rect 71 181 72 182
rect 70 181 71 182
rect 69 181 70 182
rect 68 181 69 182
rect 67 181 68 182
rect 66 181 67 182
rect 65 181 66 182
rect 64 181 65 182
rect 63 181 64 182
rect 62 181 63 182
rect 61 181 62 182
rect 60 181 61 182
rect 59 181 60 182
rect 58 181 59 182
rect 57 181 58 182
rect 56 181 57 182
rect 55 181 56 182
rect 54 181 55 182
rect 53 181 54 182
rect 52 181 53 182
rect 51 181 52 182
rect 50 181 51 182
rect 49 181 50 182
rect 48 181 49 182
rect 47 181 48 182
rect 46 181 47 182
rect 45 181 46 182
rect 44 181 45 182
rect 43 181 44 182
rect 42 181 43 182
rect 41 181 42 182
rect 40 181 41 182
rect 39 181 40 182
rect 38 181 39 182
rect 37 181 38 182
rect 36 181 37 182
rect 35 181 36 182
rect 34 181 35 182
rect 33 181 34 182
rect 32 181 33 182
rect 31 181 32 182
rect 30 181 31 182
rect 29 181 30 182
rect 28 181 29 182
rect 27 181 28 182
rect 26 181 27 182
rect 25 181 26 182
rect 24 181 25 182
rect 23 181 24 182
rect 22 181 23 182
rect 21 181 22 182
rect 20 181 21 182
rect 19 181 20 182
rect 18 181 19 182
rect 17 181 18 182
rect 16 181 17 182
rect 15 181 16 182
rect 14 181 15 182
rect 128 182 129 183
rect 127 182 128 183
rect 126 182 127 183
rect 125 182 126 183
rect 78 182 79 183
rect 77 182 78 183
rect 76 182 77 183
rect 75 182 76 183
rect 74 182 75 183
rect 73 182 74 183
rect 72 182 73 183
rect 71 182 72 183
rect 70 182 71 183
rect 69 182 70 183
rect 68 182 69 183
rect 67 182 68 183
rect 66 182 67 183
rect 65 182 66 183
rect 64 182 65 183
rect 63 182 64 183
rect 62 182 63 183
rect 61 182 62 183
rect 60 182 61 183
rect 59 182 60 183
rect 58 182 59 183
rect 57 182 58 183
rect 56 182 57 183
rect 55 182 56 183
rect 54 182 55 183
rect 53 182 54 183
rect 52 182 53 183
rect 51 182 52 183
rect 50 182 51 183
rect 49 182 50 183
rect 48 182 49 183
rect 47 182 48 183
rect 46 182 47 183
rect 45 182 46 183
rect 44 182 45 183
rect 43 182 44 183
rect 42 182 43 183
rect 41 182 42 183
rect 40 182 41 183
rect 39 182 40 183
rect 38 182 39 183
rect 37 182 38 183
rect 36 182 37 183
rect 35 182 36 183
rect 34 182 35 183
rect 33 182 34 183
rect 32 182 33 183
rect 31 182 32 183
rect 30 182 31 183
rect 29 182 30 183
rect 28 182 29 183
rect 27 182 28 183
rect 26 182 27 183
rect 25 182 26 183
rect 24 182 25 183
rect 23 182 24 183
rect 22 182 23 183
rect 21 182 22 183
rect 20 182 21 183
rect 19 182 20 183
rect 18 182 19 183
rect 17 182 18 183
rect 16 182 17 183
rect 15 182 16 183
rect 14 182 15 183
rect 127 183 128 184
rect 126 183 127 184
rect 125 183 126 184
rect 78 183 79 184
rect 77 183 78 184
rect 76 183 77 184
rect 75 183 76 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 70 183 71 184
rect 69 183 70 184
rect 68 183 69 184
rect 67 183 68 184
rect 66 183 67 184
rect 65 183 66 184
rect 64 183 65 184
rect 63 183 64 184
rect 62 183 63 184
rect 61 183 62 184
rect 60 183 61 184
rect 59 183 60 184
rect 58 183 59 184
rect 57 183 58 184
rect 56 183 57 184
rect 55 183 56 184
rect 54 183 55 184
rect 53 183 54 184
rect 52 183 53 184
rect 51 183 52 184
rect 50 183 51 184
rect 49 183 50 184
rect 48 183 49 184
rect 47 183 48 184
rect 46 183 47 184
rect 45 183 46 184
rect 44 183 45 184
rect 43 183 44 184
rect 42 183 43 184
rect 41 183 42 184
rect 40 183 41 184
rect 39 183 40 184
rect 38 183 39 184
rect 37 183 38 184
rect 36 183 37 184
rect 35 183 36 184
rect 34 183 35 184
rect 33 183 34 184
rect 32 183 33 184
rect 31 183 32 184
rect 30 183 31 184
rect 29 183 30 184
rect 28 183 29 184
rect 27 183 28 184
rect 26 183 27 184
rect 25 183 26 184
rect 24 183 25 184
rect 23 183 24 184
rect 22 183 23 184
rect 21 183 22 184
rect 20 183 21 184
rect 19 183 20 184
rect 18 183 19 184
rect 17 183 18 184
rect 16 183 17 184
rect 15 183 16 184
rect 14 183 15 184
rect 128 184 129 185
rect 127 184 128 185
rect 126 184 127 185
rect 125 184 126 185
rect 124 184 125 185
rect 77 184 78 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 70 184 71 185
rect 69 184 70 185
rect 68 184 69 185
rect 67 184 68 185
rect 66 184 67 185
rect 65 184 66 185
rect 64 184 65 185
rect 63 184 64 185
rect 62 184 63 185
rect 61 184 62 185
rect 60 184 61 185
rect 59 184 60 185
rect 58 184 59 185
rect 57 184 58 185
rect 56 184 57 185
rect 55 184 56 185
rect 54 184 55 185
rect 53 184 54 185
rect 52 184 53 185
rect 51 184 52 185
rect 50 184 51 185
rect 49 184 50 185
rect 48 184 49 185
rect 47 184 48 185
rect 46 184 47 185
rect 45 184 46 185
rect 44 184 45 185
rect 43 184 44 185
rect 42 184 43 185
rect 41 184 42 185
rect 40 184 41 185
rect 39 184 40 185
rect 38 184 39 185
rect 37 184 38 185
rect 36 184 37 185
rect 35 184 36 185
rect 34 184 35 185
rect 33 184 34 185
rect 32 184 33 185
rect 31 184 32 185
rect 30 184 31 185
rect 29 184 30 185
rect 28 184 29 185
rect 27 184 28 185
rect 26 184 27 185
rect 25 184 26 185
rect 24 184 25 185
rect 23 184 24 185
rect 22 184 23 185
rect 21 184 22 185
rect 20 184 21 185
rect 19 184 20 185
rect 18 184 19 185
rect 17 184 18 185
rect 16 184 17 185
rect 15 184 16 185
rect 14 184 15 185
rect 128 185 129 186
rect 127 185 128 186
rect 126 185 127 186
rect 125 185 126 186
rect 124 185 125 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 69 185 70 186
rect 68 185 69 186
rect 67 185 68 186
rect 66 185 67 186
rect 65 185 66 186
rect 64 185 65 186
rect 63 185 64 186
rect 62 185 63 186
rect 61 185 62 186
rect 60 185 61 186
rect 59 185 60 186
rect 58 185 59 186
rect 57 185 58 186
rect 56 185 57 186
rect 55 185 56 186
rect 54 185 55 186
rect 53 185 54 186
rect 52 185 53 186
rect 51 185 52 186
rect 50 185 51 186
rect 49 185 50 186
rect 48 185 49 186
rect 47 185 48 186
rect 46 185 47 186
rect 45 185 46 186
rect 44 185 45 186
rect 43 185 44 186
rect 42 185 43 186
rect 41 185 42 186
rect 40 185 41 186
rect 39 185 40 186
rect 38 185 39 186
rect 37 185 38 186
rect 36 185 37 186
rect 35 185 36 186
rect 34 185 35 186
rect 33 185 34 186
rect 32 185 33 186
rect 31 185 32 186
rect 30 185 31 186
rect 29 185 30 186
rect 28 185 29 186
rect 27 185 28 186
rect 26 185 27 186
rect 25 185 26 186
rect 24 185 25 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 20 185 21 186
rect 19 185 20 186
rect 18 185 19 186
rect 17 185 18 186
rect 16 185 17 186
rect 15 185 16 186
rect 14 185 15 186
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 125 186 126 187
rect 124 186 125 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 69 186 70 187
rect 68 186 69 187
rect 67 186 68 187
rect 66 186 67 187
rect 65 186 66 187
rect 64 186 65 187
rect 63 186 64 187
rect 62 186 63 187
rect 61 186 62 187
rect 60 186 61 187
rect 59 186 60 187
rect 58 186 59 187
rect 57 186 58 187
rect 56 186 57 187
rect 55 186 56 187
rect 54 186 55 187
rect 53 186 54 187
rect 52 186 53 187
rect 51 186 52 187
rect 50 186 51 187
rect 49 186 50 187
rect 48 186 49 187
rect 47 186 48 187
rect 46 186 47 187
rect 45 186 46 187
rect 44 186 45 187
rect 43 186 44 187
rect 42 186 43 187
rect 41 186 42 187
rect 40 186 41 187
rect 39 186 40 187
rect 38 186 39 187
rect 37 186 38 187
rect 36 186 37 187
rect 35 186 36 187
rect 34 186 35 187
rect 33 186 34 187
rect 32 186 33 187
rect 31 186 32 187
rect 30 186 31 187
rect 29 186 30 187
rect 28 186 29 187
rect 27 186 28 187
rect 26 186 27 187
rect 25 186 26 187
rect 24 186 25 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 19 186 20 187
rect 18 186 19 187
rect 17 186 18 187
rect 16 186 17 187
rect 15 186 16 187
rect 14 186 15 187
rect 142 187 143 188
rect 141 187 142 188
rect 140 187 141 188
rect 139 187 140 188
rect 138 187 139 188
rect 137 187 138 188
rect 136 187 137 188
rect 135 187 136 188
rect 134 187 135 188
rect 133 187 134 188
rect 132 187 133 188
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 125 187 126 188
rect 124 187 125 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 67 187 68 188
rect 66 187 67 188
rect 65 187 66 188
rect 64 187 65 188
rect 63 187 64 188
rect 62 187 63 188
rect 61 187 62 188
rect 60 187 61 188
rect 59 187 60 188
rect 58 187 59 188
rect 57 187 58 188
rect 56 187 57 188
rect 55 187 56 188
rect 54 187 55 188
rect 53 187 54 188
rect 52 187 53 188
rect 51 187 52 188
rect 50 187 51 188
rect 49 187 50 188
rect 48 187 49 188
rect 47 187 48 188
rect 46 187 47 188
rect 45 187 46 188
rect 44 187 45 188
rect 43 187 44 188
rect 42 187 43 188
rect 41 187 42 188
rect 40 187 41 188
rect 39 187 40 188
rect 38 187 39 188
rect 37 187 38 188
rect 36 187 37 188
rect 35 187 36 188
rect 34 187 35 188
rect 33 187 34 188
rect 32 187 33 188
rect 31 187 32 188
rect 30 187 31 188
rect 29 187 30 188
rect 28 187 29 188
rect 27 187 28 188
rect 26 187 27 188
rect 25 187 26 188
rect 24 187 25 188
rect 23 187 24 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 18 187 19 188
rect 17 187 18 188
rect 16 187 17 188
rect 15 187 16 188
rect 14 187 15 188
rect 142 188 143 189
rect 141 188 142 189
rect 140 188 141 189
rect 139 188 140 189
rect 138 188 139 189
rect 137 188 138 189
rect 136 188 137 189
rect 135 188 136 189
rect 134 188 135 189
rect 133 188 134 189
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 125 188 126 189
rect 124 188 125 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 66 188 67 189
rect 65 188 66 189
rect 64 188 65 189
rect 63 188 64 189
rect 62 188 63 189
rect 61 188 62 189
rect 60 188 61 189
rect 59 188 60 189
rect 58 188 59 189
rect 57 188 58 189
rect 56 188 57 189
rect 55 188 56 189
rect 54 188 55 189
rect 53 188 54 189
rect 52 188 53 189
rect 51 188 52 189
rect 50 188 51 189
rect 49 188 50 189
rect 48 188 49 189
rect 47 188 48 189
rect 46 188 47 189
rect 45 188 46 189
rect 44 188 45 189
rect 43 188 44 189
rect 42 188 43 189
rect 41 188 42 189
rect 40 188 41 189
rect 39 188 40 189
rect 38 188 39 189
rect 37 188 38 189
rect 36 188 37 189
rect 35 188 36 189
rect 34 188 35 189
rect 33 188 34 189
rect 32 188 33 189
rect 31 188 32 189
rect 30 188 31 189
rect 29 188 30 189
rect 28 188 29 189
rect 27 188 28 189
rect 26 188 27 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 17 188 18 189
rect 16 188 17 189
rect 15 188 16 189
rect 14 188 15 189
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 125 189 126 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 69 189 70 190
rect 68 189 69 190
rect 67 189 68 190
rect 66 189 67 190
rect 65 189 66 190
rect 64 189 65 190
rect 63 189 64 190
rect 62 189 63 190
rect 61 189 62 190
rect 60 189 61 190
rect 59 189 60 190
rect 58 189 59 190
rect 57 189 58 190
rect 56 189 57 190
rect 55 189 56 190
rect 54 189 55 190
rect 53 189 54 190
rect 52 189 53 190
rect 51 189 52 190
rect 50 189 51 190
rect 49 189 50 190
rect 48 189 49 190
rect 47 189 48 190
rect 46 189 47 190
rect 45 189 46 190
rect 44 189 45 190
rect 43 189 44 190
rect 42 189 43 190
rect 41 189 42 190
rect 40 189 41 190
rect 39 189 40 190
rect 38 189 39 190
rect 37 189 38 190
rect 36 189 37 190
rect 35 189 36 190
rect 34 189 35 190
rect 33 189 34 190
rect 32 189 33 190
rect 31 189 32 190
rect 30 189 31 190
rect 29 189 30 190
rect 28 189 29 190
rect 27 189 28 190
rect 26 189 27 190
rect 25 189 26 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 16 189 17 190
rect 15 189 16 190
rect 14 189 15 190
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 68 190 69 191
rect 67 190 68 191
rect 66 190 67 191
rect 65 190 66 191
rect 64 190 65 191
rect 63 190 64 191
rect 62 190 63 191
rect 61 190 62 191
rect 60 190 61 191
rect 59 190 60 191
rect 58 190 59 191
rect 57 190 58 191
rect 56 190 57 191
rect 55 190 56 191
rect 54 190 55 191
rect 53 190 54 191
rect 52 190 53 191
rect 51 190 52 191
rect 50 190 51 191
rect 49 190 50 191
rect 48 190 49 191
rect 47 190 48 191
rect 46 190 47 191
rect 45 190 46 191
rect 44 190 45 191
rect 43 190 44 191
rect 42 190 43 191
rect 41 190 42 191
rect 40 190 41 191
rect 39 190 40 191
rect 38 190 39 191
rect 37 190 38 191
rect 36 190 37 191
rect 35 190 36 191
rect 34 190 35 191
rect 33 190 34 191
rect 32 190 33 191
rect 31 190 32 191
rect 30 190 31 191
rect 29 190 30 191
rect 28 190 29 191
rect 27 190 28 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 16 190 17 191
rect 15 190 16 191
rect 14 190 15 191
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 72 191 73 192
rect 71 191 72 192
rect 70 191 71 192
rect 69 191 70 192
rect 68 191 69 192
rect 67 191 68 192
rect 66 191 67 192
rect 65 191 66 192
rect 64 191 65 192
rect 63 191 64 192
rect 62 191 63 192
rect 61 191 62 192
rect 60 191 61 192
rect 59 191 60 192
rect 58 191 59 192
rect 57 191 58 192
rect 56 191 57 192
rect 55 191 56 192
rect 54 191 55 192
rect 53 191 54 192
rect 52 191 53 192
rect 51 191 52 192
rect 50 191 51 192
rect 49 191 50 192
rect 48 191 49 192
rect 47 191 48 192
rect 46 191 47 192
rect 45 191 46 192
rect 44 191 45 192
rect 43 191 44 192
rect 42 191 43 192
rect 41 191 42 192
rect 40 191 41 192
rect 39 191 40 192
rect 38 191 39 192
rect 37 191 38 192
rect 36 191 37 192
rect 35 191 36 192
rect 34 191 35 192
rect 33 191 34 192
rect 32 191 33 192
rect 31 191 32 192
rect 30 191 31 192
rect 29 191 30 192
rect 28 191 29 192
rect 27 191 28 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 15 191 16 192
rect 14 191 15 192
rect 70 192 71 193
rect 69 192 70 193
rect 68 192 69 193
rect 67 192 68 193
rect 66 192 67 193
rect 65 192 66 193
rect 64 192 65 193
rect 63 192 64 193
rect 62 192 63 193
rect 61 192 62 193
rect 60 192 61 193
rect 59 192 60 193
rect 58 192 59 193
rect 57 192 58 193
rect 56 192 57 193
rect 55 192 56 193
rect 54 192 55 193
rect 53 192 54 193
rect 52 192 53 193
rect 51 192 52 193
rect 50 192 51 193
rect 49 192 50 193
rect 48 192 49 193
rect 47 192 48 193
rect 46 192 47 193
rect 45 192 46 193
rect 44 192 45 193
rect 43 192 44 193
rect 42 192 43 193
rect 41 192 42 193
rect 40 192 41 193
rect 39 192 40 193
rect 38 192 39 193
rect 37 192 38 193
rect 36 192 37 193
rect 35 192 36 193
rect 34 192 35 193
rect 33 192 34 193
rect 32 192 33 193
rect 31 192 32 193
rect 30 192 31 193
rect 29 192 30 193
rect 28 192 29 193
rect 27 192 28 193
rect 26 192 27 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 16 192 17 193
rect 15 192 16 193
rect 14 192 15 193
rect 69 193 70 194
rect 68 193 69 194
rect 67 193 68 194
rect 66 193 67 194
rect 65 193 66 194
rect 64 193 65 194
rect 63 193 64 194
rect 62 193 63 194
rect 61 193 62 194
rect 60 193 61 194
rect 59 193 60 194
rect 58 193 59 194
rect 57 193 58 194
rect 56 193 57 194
rect 55 193 56 194
rect 54 193 55 194
rect 53 193 54 194
rect 52 193 53 194
rect 51 193 52 194
rect 50 193 51 194
rect 49 193 50 194
rect 48 193 49 194
rect 47 193 48 194
rect 46 193 47 194
rect 45 193 46 194
rect 44 193 45 194
rect 43 193 44 194
rect 42 193 43 194
rect 41 193 42 194
rect 40 193 41 194
rect 39 193 40 194
rect 38 193 39 194
rect 37 193 38 194
rect 36 193 37 194
rect 35 193 36 194
rect 34 193 35 194
rect 33 193 34 194
rect 32 193 33 194
rect 31 193 32 194
rect 30 193 31 194
rect 29 193 30 194
rect 28 193 29 194
rect 27 193 28 194
rect 26 193 27 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 16 193 17 194
rect 15 193 16 194
rect 14 193 15 194
rect 67 194 68 195
rect 66 194 67 195
rect 65 194 66 195
rect 64 194 65 195
rect 63 194 64 195
rect 62 194 63 195
rect 61 194 62 195
rect 60 194 61 195
rect 59 194 60 195
rect 58 194 59 195
rect 57 194 58 195
rect 56 194 57 195
rect 55 194 56 195
rect 54 194 55 195
rect 53 194 54 195
rect 52 194 53 195
rect 51 194 52 195
rect 50 194 51 195
rect 49 194 50 195
rect 48 194 49 195
rect 47 194 48 195
rect 46 194 47 195
rect 45 194 46 195
rect 44 194 45 195
rect 43 194 44 195
rect 42 194 43 195
rect 41 194 42 195
rect 40 194 41 195
rect 39 194 40 195
rect 38 194 39 195
rect 37 194 38 195
rect 36 194 37 195
rect 35 194 36 195
rect 34 194 35 195
rect 33 194 34 195
rect 32 194 33 195
rect 31 194 32 195
rect 30 194 31 195
rect 29 194 30 195
rect 28 194 29 195
rect 27 194 28 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 17 194 18 195
rect 16 194 17 195
rect 15 194 16 195
rect 14 194 15 195
rect 64 195 65 196
rect 63 195 64 196
rect 62 195 63 196
rect 61 195 62 196
rect 60 195 61 196
rect 59 195 60 196
rect 58 195 59 196
rect 57 195 58 196
rect 56 195 57 196
rect 55 195 56 196
rect 54 195 55 196
rect 53 195 54 196
rect 52 195 53 196
rect 51 195 52 196
rect 50 195 51 196
rect 49 195 50 196
rect 48 195 49 196
rect 47 195 48 196
rect 46 195 47 196
rect 45 195 46 196
rect 44 195 45 196
rect 43 195 44 196
rect 42 195 43 196
rect 41 195 42 196
rect 40 195 41 196
rect 39 195 40 196
rect 38 195 39 196
rect 37 195 38 196
rect 36 195 37 196
rect 35 195 36 196
rect 34 195 35 196
rect 33 195 34 196
rect 32 195 33 196
rect 31 195 32 196
rect 30 195 31 196
rect 29 195 30 196
rect 28 195 29 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 17 195 18 196
rect 16 195 17 196
rect 15 195 16 196
rect 14 195 15 196
rect 140 196 141 197
rect 139 196 140 197
rect 61 196 62 197
rect 60 196 61 197
rect 59 196 60 197
rect 58 196 59 197
rect 57 196 58 197
rect 56 196 57 197
rect 55 196 56 197
rect 54 196 55 197
rect 53 196 54 197
rect 52 196 53 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 48 196 49 197
rect 47 196 48 197
rect 46 196 47 197
rect 45 196 46 197
rect 44 196 45 197
rect 43 196 44 197
rect 42 196 43 197
rect 41 196 42 197
rect 40 196 41 197
rect 39 196 40 197
rect 38 196 39 197
rect 37 196 38 197
rect 36 196 37 197
rect 35 196 36 197
rect 34 196 35 197
rect 33 196 34 197
rect 32 196 33 197
rect 31 196 32 197
rect 30 196 31 197
rect 29 196 30 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 17 196 18 197
rect 16 196 17 197
rect 15 196 16 197
rect 14 196 15 197
rect 141 197 142 198
rect 140 197 141 198
rect 139 197 140 198
rect 138 197 139 198
rect 53 197 54 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 48 197 49 198
rect 47 197 48 198
rect 46 197 47 198
rect 45 197 46 198
rect 44 197 45 198
rect 43 197 44 198
rect 42 197 43 198
rect 41 197 42 198
rect 40 197 41 198
rect 39 197 40 198
rect 38 197 39 198
rect 37 197 38 198
rect 36 197 37 198
rect 35 197 36 198
rect 34 197 35 198
rect 33 197 34 198
rect 32 197 33 198
rect 31 197 32 198
rect 30 197 31 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 17 197 18 198
rect 16 197 17 198
rect 15 197 16 198
rect 14 197 15 198
rect 142 198 143 199
rect 141 198 142 199
rect 140 198 141 199
rect 139 198 140 199
rect 138 198 139 199
rect 137 198 138 199
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 139 199 140 200
rect 138 199 139 200
rect 137 199 138 200
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 138 200 139 201
rect 137 200 138 201
rect 141 201 142 202
rect 140 201 141 202
rect 139 201 140 202
rect 138 201 139 202
rect 140 202 141 203
rect 139 202 140 203
rect 138 218 139 219
rect 137 218 138 219
rect 136 218 137 219
rect 135 218 136 219
rect 134 218 135 219
rect 133 218 134 219
rect 132 218 133 219
rect 131 218 132 219
rect 130 218 131 219
rect 129 218 130 219
rect 128 218 129 219
rect 141 219 142 220
rect 140 219 141 220
rect 139 219 140 220
rect 138 219 139 220
rect 137 219 138 220
rect 136 219 137 220
rect 135 219 136 220
rect 134 219 135 220
rect 133 219 134 220
rect 132 219 133 220
rect 131 219 132 220
rect 130 219 131 220
rect 129 219 130 220
rect 128 219 129 220
rect 127 219 128 220
rect 126 219 127 220
rect 125 219 126 220
rect 124 219 125 220
rect 143 220 144 221
rect 142 220 143 221
rect 141 220 142 221
rect 140 220 141 221
rect 139 220 140 221
rect 138 220 139 221
rect 137 220 138 221
rect 136 220 137 221
rect 135 220 136 221
rect 134 220 135 221
rect 133 220 134 221
rect 132 220 133 221
rect 131 220 132 221
rect 130 220 131 221
rect 129 220 130 221
rect 128 220 129 221
rect 127 220 128 221
rect 126 220 127 221
rect 125 220 126 221
rect 124 220 125 221
rect 123 220 124 221
rect 122 220 123 221
rect 145 221 146 222
rect 144 221 145 222
rect 143 221 144 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 139 221 140 222
rect 138 221 139 222
rect 137 221 138 222
rect 136 221 137 222
rect 135 221 136 222
rect 134 221 135 222
rect 133 221 134 222
rect 132 221 133 222
rect 131 221 132 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 125 221 126 222
rect 124 221 125 222
rect 123 221 124 222
rect 122 221 123 222
rect 121 221 122 222
rect 120 221 121 222
rect 147 222 148 223
rect 146 222 147 223
rect 145 222 146 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 137 222 138 223
rect 136 222 137 223
rect 135 222 136 223
rect 134 222 135 223
rect 133 222 134 223
rect 132 222 133 223
rect 131 222 132 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 123 222 124 223
rect 122 222 123 223
rect 121 222 122 223
rect 120 222 121 223
rect 119 222 120 223
rect 148 223 149 224
rect 147 223 148 224
rect 146 223 147 224
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 121 223 122 224
rect 120 223 121 224
rect 119 223 120 224
rect 118 223 119 224
rect 117 223 118 224
rect 148 224 149 225
rect 147 224 148 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 120 224 121 225
rect 119 224 120 225
rect 118 224 119 225
rect 117 224 118 225
rect 148 225 149 226
rect 147 225 148 226
rect 146 225 147 226
rect 145 225 146 226
rect 121 225 122 226
rect 120 225 121 226
rect 119 225 120 226
rect 118 225 119 226
rect 117 225 118 226
rect 148 226 149 227
rect 147 226 148 227
rect 146 226 147 227
rect 119 226 120 227
rect 118 226 119 227
rect 117 226 118 227
rect 148 227 149 228
rect 117 227 118 228
rect 136 230 137 231
rect 135 230 136 231
rect 134 230 135 231
rect 133 230 134 231
rect 132 230 133 231
rect 131 230 132 231
rect 138 231 139 232
rect 137 231 138 232
rect 136 231 137 232
rect 135 231 136 232
rect 134 231 135 232
rect 133 231 134 232
rect 132 231 133 232
rect 131 231 132 232
rect 130 231 131 232
rect 129 231 130 232
rect 128 231 129 232
rect 139 232 140 233
rect 138 232 139 233
rect 137 232 138 233
rect 136 232 137 233
rect 135 232 136 233
rect 134 232 135 233
rect 133 232 134 233
rect 132 232 133 233
rect 131 232 132 233
rect 130 232 131 233
rect 129 232 130 233
rect 128 232 129 233
rect 127 232 128 233
rect 140 233 141 234
rect 139 233 140 234
rect 138 233 139 234
rect 137 233 138 234
rect 136 233 137 234
rect 135 233 136 234
rect 134 233 135 234
rect 133 233 134 234
rect 132 233 133 234
rect 131 233 132 234
rect 130 233 131 234
rect 129 233 130 234
rect 128 233 129 234
rect 127 233 128 234
rect 126 233 127 234
rect 141 234 142 235
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 137 234 138 235
rect 136 234 137 235
rect 135 234 136 235
rect 134 234 135 235
rect 133 234 134 235
rect 132 234 133 235
rect 131 234 132 235
rect 130 234 131 235
rect 129 234 130 235
rect 128 234 129 235
rect 127 234 128 235
rect 126 234 127 235
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 137 235 138 236
rect 136 235 137 236
rect 135 235 136 236
rect 134 235 135 236
rect 133 235 134 236
rect 132 235 133 236
rect 131 235 132 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 127 235 128 236
rect 126 235 127 236
rect 125 235 126 236
rect 59 235 60 236
rect 58 235 59 236
rect 57 235 58 236
rect 56 235 57 236
rect 55 235 56 236
rect 54 235 55 236
rect 53 235 54 236
rect 52 235 53 236
rect 51 235 52 236
rect 50 235 51 236
rect 49 235 50 236
rect 48 235 49 236
rect 47 235 48 236
rect 46 235 47 236
rect 45 235 46 236
rect 44 235 45 236
rect 43 235 44 236
rect 42 235 43 236
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 137 236 138 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 127 236 128 237
rect 126 236 127 237
rect 125 236 126 237
rect 63 236 64 237
rect 62 236 63 237
rect 61 236 62 237
rect 60 236 61 237
rect 59 236 60 237
rect 58 236 59 237
rect 57 236 58 237
rect 56 236 57 237
rect 55 236 56 237
rect 54 236 55 237
rect 53 236 54 237
rect 52 236 53 237
rect 51 236 52 237
rect 50 236 51 237
rect 49 236 50 237
rect 48 236 49 237
rect 47 236 48 237
rect 46 236 47 237
rect 45 236 46 237
rect 44 236 45 237
rect 43 236 44 237
rect 42 236 43 237
rect 41 236 42 237
rect 40 236 41 237
rect 39 236 40 237
rect 38 236 39 237
rect 37 236 38 237
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 128 237 129 238
rect 127 237 128 238
rect 126 237 127 238
rect 125 237 126 238
rect 124 237 125 238
rect 66 237 67 238
rect 65 237 66 238
rect 64 237 65 238
rect 63 237 64 238
rect 62 237 63 238
rect 61 237 62 238
rect 60 237 61 238
rect 59 237 60 238
rect 58 237 59 238
rect 57 237 58 238
rect 56 237 57 238
rect 55 237 56 238
rect 54 237 55 238
rect 53 237 54 238
rect 52 237 53 238
rect 51 237 52 238
rect 50 237 51 238
rect 49 237 50 238
rect 48 237 49 238
rect 47 237 48 238
rect 46 237 47 238
rect 45 237 46 238
rect 44 237 45 238
rect 43 237 44 238
rect 42 237 43 238
rect 41 237 42 238
rect 40 237 41 238
rect 39 237 40 238
rect 38 237 39 238
rect 37 237 38 238
rect 36 237 37 238
rect 35 237 36 238
rect 34 237 35 238
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 138 238 139 239
rect 128 238 129 239
rect 127 238 128 239
rect 126 238 127 239
rect 125 238 126 239
rect 124 238 125 239
rect 68 238 69 239
rect 67 238 68 239
rect 66 238 67 239
rect 65 238 66 239
rect 64 238 65 239
rect 63 238 64 239
rect 62 238 63 239
rect 61 238 62 239
rect 60 238 61 239
rect 59 238 60 239
rect 58 238 59 239
rect 57 238 58 239
rect 56 238 57 239
rect 55 238 56 239
rect 54 238 55 239
rect 53 238 54 239
rect 52 238 53 239
rect 51 238 52 239
rect 50 238 51 239
rect 49 238 50 239
rect 48 238 49 239
rect 47 238 48 239
rect 46 238 47 239
rect 45 238 46 239
rect 44 238 45 239
rect 43 238 44 239
rect 42 238 43 239
rect 41 238 42 239
rect 40 238 41 239
rect 39 238 40 239
rect 38 238 39 239
rect 37 238 38 239
rect 36 238 37 239
rect 35 238 36 239
rect 34 238 35 239
rect 33 238 34 239
rect 32 238 33 239
rect 31 238 32 239
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 139 239 140 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 125 239 126 240
rect 124 239 125 240
rect 70 239 71 240
rect 69 239 70 240
rect 68 239 69 240
rect 67 239 68 240
rect 66 239 67 240
rect 65 239 66 240
rect 64 239 65 240
rect 63 239 64 240
rect 62 239 63 240
rect 61 239 62 240
rect 60 239 61 240
rect 59 239 60 240
rect 58 239 59 240
rect 57 239 58 240
rect 56 239 57 240
rect 55 239 56 240
rect 54 239 55 240
rect 53 239 54 240
rect 52 239 53 240
rect 51 239 52 240
rect 50 239 51 240
rect 49 239 50 240
rect 48 239 49 240
rect 47 239 48 240
rect 46 239 47 240
rect 45 239 46 240
rect 44 239 45 240
rect 43 239 44 240
rect 42 239 43 240
rect 41 239 42 240
rect 40 239 41 240
rect 39 239 40 240
rect 38 239 39 240
rect 37 239 38 240
rect 36 239 37 240
rect 35 239 36 240
rect 34 239 35 240
rect 33 239 34 240
rect 32 239 33 240
rect 31 239 32 240
rect 30 239 31 240
rect 29 239 30 240
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 139 240 140 241
rect 127 240 128 241
rect 126 240 127 241
rect 125 240 126 241
rect 124 240 125 241
rect 72 240 73 241
rect 71 240 72 241
rect 70 240 71 241
rect 69 240 70 241
rect 68 240 69 241
rect 67 240 68 241
rect 66 240 67 241
rect 65 240 66 241
rect 64 240 65 241
rect 63 240 64 241
rect 62 240 63 241
rect 61 240 62 241
rect 60 240 61 241
rect 59 240 60 241
rect 58 240 59 241
rect 57 240 58 241
rect 56 240 57 241
rect 55 240 56 241
rect 54 240 55 241
rect 53 240 54 241
rect 52 240 53 241
rect 51 240 52 241
rect 50 240 51 241
rect 49 240 50 241
rect 48 240 49 241
rect 47 240 48 241
rect 46 240 47 241
rect 45 240 46 241
rect 44 240 45 241
rect 43 240 44 241
rect 42 240 43 241
rect 41 240 42 241
rect 40 240 41 241
rect 39 240 40 241
rect 38 240 39 241
rect 37 240 38 241
rect 36 240 37 241
rect 35 240 36 241
rect 34 240 35 241
rect 33 240 34 241
rect 32 240 33 241
rect 31 240 32 241
rect 30 240 31 241
rect 29 240 30 241
rect 28 240 29 241
rect 142 241 143 242
rect 141 241 142 242
rect 140 241 141 242
rect 139 241 140 242
rect 127 241 128 242
rect 126 241 127 242
rect 125 241 126 242
rect 124 241 125 242
rect 73 241 74 242
rect 72 241 73 242
rect 71 241 72 242
rect 70 241 71 242
rect 69 241 70 242
rect 68 241 69 242
rect 67 241 68 242
rect 66 241 67 242
rect 65 241 66 242
rect 64 241 65 242
rect 63 241 64 242
rect 62 241 63 242
rect 61 241 62 242
rect 60 241 61 242
rect 59 241 60 242
rect 58 241 59 242
rect 57 241 58 242
rect 56 241 57 242
rect 55 241 56 242
rect 54 241 55 242
rect 53 241 54 242
rect 52 241 53 242
rect 51 241 52 242
rect 50 241 51 242
rect 49 241 50 242
rect 48 241 49 242
rect 47 241 48 242
rect 46 241 47 242
rect 45 241 46 242
rect 44 241 45 242
rect 43 241 44 242
rect 42 241 43 242
rect 41 241 42 242
rect 40 241 41 242
rect 39 241 40 242
rect 38 241 39 242
rect 37 241 38 242
rect 36 241 37 242
rect 35 241 36 242
rect 34 241 35 242
rect 33 241 34 242
rect 32 241 33 242
rect 31 241 32 242
rect 30 241 31 242
rect 29 241 30 242
rect 28 241 29 242
rect 27 241 28 242
rect 26 241 27 242
rect 142 242 143 243
rect 141 242 142 243
rect 140 242 141 243
rect 139 242 140 243
rect 138 242 139 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 125 242 126 243
rect 124 242 125 243
rect 74 242 75 243
rect 73 242 74 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 56 242 57 243
rect 55 242 56 243
rect 54 242 55 243
rect 53 242 54 243
rect 52 242 53 243
rect 51 242 52 243
rect 50 242 51 243
rect 49 242 50 243
rect 48 242 49 243
rect 47 242 48 243
rect 46 242 47 243
rect 45 242 46 243
rect 44 242 45 243
rect 43 242 44 243
rect 42 242 43 243
rect 41 242 42 243
rect 40 242 41 243
rect 39 242 40 243
rect 38 242 39 243
rect 37 242 38 243
rect 36 242 37 243
rect 35 242 36 243
rect 34 242 35 243
rect 33 242 34 243
rect 32 242 33 243
rect 31 242 32 243
rect 30 242 31 243
rect 29 242 30 243
rect 28 242 29 243
rect 27 242 28 243
rect 26 242 27 243
rect 25 242 26 243
rect 142 243 143 244
rect 141 243 142 244
rect 140 243 141 244
rect 139 243 140 244
rect 138 243 139 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 125 243 126 244
rect 124 243 125 244
rect 75 243 76 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 56 243 57 244
rect 55 243 56 244
rect 54 243 55 244
rect 53 243 54 244
rect 52 243 53 244
rect 51 243 52 244
rect 50 243 51 244
rect 49 243 50 244
rect 48 243 49 244
rect 47 243 48 244
rect 46 243 47 244
rect 45 243 46 244
rect 44 243 45 244
rect 43 243 44 244
rect 42 243 43 244
rect 41 243 42 244
rect 40 243 41 244
rect 39 243 40 244
rect 38 243 39 244
rect 37 243 38 244
rect 36 243 37 244
rect 35 243 36 244
rect 34 243 35 244
rect 33 243 34 244
rect 32 243 33 244
rect 31 243 32 244
rect 30 243 31 244
rect 29 243 30 244
rect 28 243 29 244
rect 27 243 28 244
rect 26 243 27 244
rect 25 243 26 244
rect 24 243 25 244
rect 23 243 24 244
rect 141 244 142 245
rect 140 244 141 245
rect 139 244 140 245
rect 138 244 139 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 125 244 126 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 56 244 57 245
rect 55 244 56 245
rect 54 244 55 245
rect 53 244 54 245
rect 52 244 53 245
rect 51 244 52 245
rect 50 244 51 245
rect 49 244 50 245
rect 48 244 49 245
rect 47 244 48 245
rect 46 244 47 245
rect 45 244 46 245
rect 44 244 45 245
rect 43 244 44 245
rect 42 244 43 245
rect 41 244 42 245
rect 40 244 41 245
rect 39 244 40 245
rect 38 244 39 245
rect 37 244 38 245
rect 36 244 37 245
rect 35 244 36 245
rect 34 244 35 245
rect 33 244 34 245
rect 32 244 33 245
rect 31 244 32 245
rect 30 244 31 245
rect 29 244 30 245
rect 28 244 29 245
rect 27 244 28 245
rect 26 244 27 245
rect 25 244 26 245
rect 24 244 25 245
rect 23 244 24 245
rect 22 244 23 245
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 56 245 57 246
rect 55 245 56 246
rect 54 245 55 246
rect 53 245 54 246
rect 52 245 53 246
rect 51 245 52 246
rect 50 245 51 246
rect 49 245 50 246
rect 48 245 49 246
rect 47 245 48 246
rect 46 245 47 246
rect 45 245 46 246
rect 44 245 45 246
rect 43 245 44 246
rect 42 245 43 246
rect 41 245 42 246
rect 40 245 41 246
rect 39 245 40 246
rect 38 245 39 246
rect 37 245 38 246
rect 36 245 37 246
rect 35 245 36 246
rect 34 245 35 246
rect 33 245 34 246
rect 32 245 33 246
rect 31 245 32 246
rect 30 245 31 246
rect 29 245 30 246
rect 28 245 29 246
rect 27 245 28 246
rect 26 245 27 246
rect 25 245 26 246
rect 24 245 25 246
rect 23 245 24 246
rect 22 245 23 246
rect 21 245 22 246
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 56 246 57 247
rect 55 246 56 247
rect 54 246 55 247
rect 53 246 54 247
rect 52 246 53 247
rect 51 246 52 247
rect 50 246 51 247
rect 49 246 50 247
rect 48 246 49 247
rect 47 246 48 247
rect 46 246 47 247
rect 45 246 46 247
rect 44 246 45 247
rect 43 246 44 247
rect 42 246 43 247
rect 41 246 42 247
rect 40 246 41 247
rect 39 246 40 247
rect 38 246 39 247
rect 37 246 38 247
rect 36 246 37 247
rect 35 246 36 247
rect 34 246 35 247
rect 33 246 34 247
rect 32 246 33 247
rect 31 246 32 247
rect 30 246 31 247
rect 29 246 30 247
rect 28 246 29 247
rect 27 246 28 247
rect 26 246 27 247
rect 25 246 26 247
rect 24 246 25 247
rect 23 246 24 247
rect 22 246 23 247
rect 21 246 22 247
rect 20 246 21 247
rect 148 247 149 248
rect 117 247 118 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 58 247 59 248
rect 57 247 58 248
rect 56 247 57 248
rect 55 247 56 248
rect 54 247 55 248
rect 53 247 54 248
rect 52 247 53 248
rect 51 247 52 248
rect 50 247 51 248
rect 49 247 50 248
rect 48 247 49 248
rect 47 247 48 248
rect 46 247 47 248
rect 45 247 46 248
rect 44 247 45 248
rect 43 247 44 248
rect 42 247 43 248
rect 41 247 42 248
rect 40 247 41 248
rect 39 247 40 248
rect 38 247 39 248
rect 37 247 38 248
rect 36 247 37 248
rect 35 247 36 248
rect 34 247 35 248
rect 33 247 34 248
rect 32 247 33 248
rect 31 247 32 248
rect 30 247 31 248
rect 29 247 30 248
rect 28 247 29 248
rect 27 247 28 248
rect 26 247 27 248
rect 25 247 26 248
rect 24 247 25 248
rect 23 247 24 248
rect 22 247 23 248
rect 21 247 22 248
rect 20 247 21 248
rect 19 247 20 248
rect 148 248 149 249
rect 147 248 148 249
rect 118 248 119 249
rect 117 248 118 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 57 248 58 249
rect 56 248 57 249
rect 55 248 56 249
rect 54 248 55 249
rect 53 248 54 249
rect 52 248 53 249
rect 51 248 52 249
rect 50 248 51 249
rect 49 248 50 249
rect 48 248 49 249
rect 47 248 48 249
rect 46 248 47 249
rect 45 248 46 249
rect 44 248 45 249
rect 43 248 44 249
rect 42 248 43 249
rect 41 248 42 249
rect 40 248 41 249
rect 39 248 40 249
rect 38 248 39 249
rect 37 248 38 249
rect 36 248 37 249
rect 35 248 36 249
rect 34 248 35 249
rect 33 248 34 249
rect 32 248 33 249
rect 31 248 32 249
rect 30 248 31 249
rect 29 248 30 249
rect 28 248 29 249
rect 27 248 28 249
rect 26 248 27 249
rect 25 248 26 249
rect 24 248 25 249
rect 23 248 24 249
rect 22 248 23 249
rect 21 248 22 249
rect 20 248 21 249
rect 19 248 20 249
rect 148 249 149 250
rect 147 249 148 250
rect 146 249 147 250
rect 145 249 146 250
rect 120 249 121 250
rect 119 249 120 250
rect 118 249 119 250
rect 117 249 118 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 56 249 57 250
rect 55 249 56 250
rect 54 249 55 250
rect 53 249 54 250
rect 52 249 53 250
rect 51 249 52 250
rect 50 249 51 250
rect 49 249 50 250
rect 48 249 49 250
rect 47 249 48 250
rect 46 249 47 250
rect 45 249 46 250
rect 44 249 45 250
rect 43 249 44 250
rect 42 249 43 250
rect 41 249 42 250
rect 40 249 41 250
rect 39 249 40 250
rect 38 249 39 250
rect 37 249 38 250
rect 36 249 37 250
rect 35 249 36 250
rect 34 249 35 250
rect 33 249 34 250
rect 32 249 33 250
rect 31 249 32 250
rect 30 249 31 250
rect 29 249 30 250
rect 28 249 29 250
rect 27 249 28 250
rect 26 249 27 250
rect 25 249 26 250
rect 24 249 25 250
rect 23 249 24 250
rect 22 249 23 250
rect 21 249 22 250
rect 20 249 21 250
rect 19 249 20 250
rect 18 249 19 250
rect 148 250 149 251
rect 147 250 148 251
rect 146 250 147 251
rect 145 250 146 251
rect 144 250 145 251
rect 143 250 144 251
rect 122 250 123 251
rect 121 250 122 251
rect 120 250 121 251
rect 119 250 120 251
rect 118 250 119 251
rect 117 250 118 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 56 250 57 251
rect 55 250 56 251
rect 54 250 55 251
rect 53 250 54 251
rect 52 250 53 251
rect 51 250 52 251
rect 50 250 51 251
rect 49 250 50 251
rect 48 250 49 251
rect 47 250 48 251
rect 46 250 47 251
rect 45 250 46 251
rect 44 250 45 251
rect 43 250 44 251
rect 42 250 43 251
rect 41 250 42 251
rect 40 250 41 251
rect 39 250 40 251
rect 38 250 39 251
rect 37 250 38 251
rect 36 250 37 251
rect 35 250 36 251
rect 34 250 35 251
rect 33 250 34 251
rect 32 250 33 251
rect 31 250 32 251
rect 30 250 31 251
rect 29 250 30 251
rect 28 250 29 251
rect 27 250 28 251
rect 26 250 27 251
rect 25 250 26 251
rect 24 250 25 251
rect 23 250 24 251
rect 22 250 23 251
rect 21 250 22 251
rect 20 250 21 251
rect 19 250 20 251
rect 18 250 19 251
rect 17 250 18 251
rect 148 251 149 252
rect 147 251 148 252
rect 146 251 147 252
rect 145 251 146 252
rect 144 251 145 252
rect 143 251 144 252
rect 142 251 143 252
rect 141 251 142 252
rect 124 251 125 252
rect 123 251 124 252
rect 122 251 123 252
rect 121 251 122 252
rect 120 251 121 252
rect 119 251 120 252
rect 118 251 119 252
rect 117 251 118 252
rect 80 251 81 252
rect 79 251 80 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 71 251 72 252
rect 70 251 71 252
rect 69 251 70 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 56 251 57 252
rect 55 251 56 252
rect 54 251 55 252
rect 53 251 54 252
rect 52 251 53 252
rect 51 251 52 252
rect 50 251 51 252
rect 49 251 50 252
rect 48 251 49 252
rect 47 251 48 252
rect 46 251 47 252
rect 45 251 46 252
rect 44 251 45 252
rect 43 251 44 252
rect 42 251 43 252
rect 41 251 42 252
rect 40 251 41 252
rect 39 251 40 252
rect 38 251 39 252
rect 37 251 38 252
rect 36 251 37 252
rect 35 251 36 252
rect 34 251 35 252
rect 33 251 34 252
rect 32 251 33 252
rect 31 251 32 252
rect 30 251 31 252
rect 29 251 30 252
rect 28 251 29 252
rect 27 251 28 252
rect 26 251 27 252
rect 25 251 26 252
rect 24 251 25 252
rect 23 251 24 252
rect 22 251 23 252
rect 21 251 22 252
rect 20 251 21 252
rect 19 251 20 252
rect 18 251 19 252
rect 17 251 18 252
rect 147 252 148 253
rect 146 252 147 253
rect 145 252 146 253
rect 144 252 145 253
rect 143 252 144 253
rect 142 252 143 253
rect 141 252 142 253
rect 140 252 141 253
rect 139 252 140 253
rect 138 252 139 253
rect 137 252 138 253
rect 136 252 137 253
rect 129 252 130 253
rect 128 252 129 253
rect 127 252 128 253
rect 126 252 127 253
rect 125 252 126 253
rect 124 252 125 253
rect 123 252 124 253
rect 122 252 123 253
rect 121 252 122 253
rect 120 252 121 253
rect 119 252 120 253
rect 118 252 119 253
rect 80 252 81 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 72 252 73 253
rect 71 252 72 253
rect 70 252 71 253
rect 69 252 70 253
rect 68 252 69 253
rect 67 252 68 253
rect 66 252 67 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 55 252 56 253
rect 54 252 55 253
rect 53 252 54 253
rect 52 252 53 253
rect 51 252 52 253
rect 50 252 51 253
rect 49 252 50 253
rect 48 252 49 253
rect 47 252 48 253
rect 46 252 47 253
rect 45 252 46 253
rect 44 252 45 253
rect 43 252 44 253
rect 42 252 43 253
rect 41 252 42 253
rect 40 252 41 253
rect 39 252 40 253
rect 38 252 39 253
rect 37 252 38 253
rect 36 252 37 253
rect 35 252 36 253
rect 34 252 35 253
rect 33 252 34 253
rect 32 252 33 253
rect 31 252 32 253
rect 30 252 31 253
rect 29 252 30 253
rect 28 252 29 253
rect 27 252 28 253
rect 26 252 27 253
rect 25 252 26 253
rect 24 252 25 253
rect 23 252 24 253
rect 22 252 23 253
rect 21 252 22 253
rect 20 252 21 253
rect 19 252 20 253
rect 18 252 19 253
rect 17 252 18 253
rect 16 252 17 253
rect 146 253 147 254
rect 145 253 146 254
rect 144 253 145 254
rect 143 253 144 254
rect 142 253 143 254
rect 141 253 142 254
rect 140 253 141 254
rect 139 253 140 254
rect 138 253 139 254
rect 137 253 138 254
rect 136 253 137 254
rect 135 253 136 254
rect 134 253 135 254
rect 133 253 134 254
rect 132 253 133 254
rect 131 253 132 254
rect 130 253 131 254
rect 129 253 130 254
rect 128 253 129 254
rect 127 253 128 254
rect 126 253 127 254
rect 125 253 126 254
rect 124 253 125 254
rect 123 253 124 254
rect 122 253 123 254
rect 121 253 122 254
rect 120 253 121 254
rect 119 253 120 254
rect 80 253 81 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 72 253 73 254
rect 71 253 72 254
rect 70 253 71 254
rect 69 253 70 254
rect 68 253 69 254
rect 67 253 68 254
rect 66 253 67 254
rect 65 253 66 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 60 253 61 254
rect 59 253 60 254
rect 58 253 59 254
rect 57 253 58 254
rect 56 253 57 254
rect 55 253 56 254
rect 54 253 55 254
rect 53 253 54 254
rect 52 253 53 254
rect 51 253 52 254
rect 50 253 51 254
rect 49 253 50 254
rect 48 253 49 254
rect 47 253 48 254
rect 46 253 47 254
rect 45 253 46 254
rect 44 253 45 254
rect 43 253 44 254
rect 42 253 43 254
rect 41 253 42 254
rect 40 253 41 254
rect 39 253 40 254
rect 38 253 39 254
rect 37 253 38 254
rect 36 253 37 254
rect 35 253 36 254
rect 34 253 35 254
rect 33 253 34 254
rect 32 253 33 254
rect 31 253 32 254
rect 30 253 31 254
rect 29 253 30 254
rect 28 253 29 254
rect 27 253 28 254
rect 26 253 27 254
rect 25 253 26 254
rect 24 253 25 254
rect 23 253 24 254
rect 22 253 23 254
rect 21 253 22 254
rect 20 253 21 254
rect 19 253 20 254
rect 18 253 19 254
rect 17 253 18 254
rect 16 253 17 254
rect 144 254 145 255
rect 143 254 144 255
rect 142 254 143 255
rect 141 254 142 255
rect 140 254 141 255
rect 139 254 140 255
rect 138 254 139 255
rect 137 254 138 255
rect 136 254 137 255
rect 135 254 136 255
rect 134 254 135 255
rect 133 254 134 255
rect 132 254 133 255
rect 131 254 132 255
rect 130 254 131 255
rect 129 254 130 255
rect 128 254 129 255
rect 127 254 128 255
rect 126 254 127 255
rect 125 254 126 255
rect 124 254 125 255
rect 123 254 124 255
rect 122 254 123 255
rect 121 254 122 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 71 254 72 255
rect 70 254 71 255
rect 69 254 70 255
rect 68 254 69 255
rect 67 254 68 255
rect 66 254 67 255
rect 65 254 66 255
rect 64 254 65 255
rect 63 254 64 255
rect 62 254 63 255
rect 61 254 62 255
rect 60 254 61 255
rect 57 254 58 255
rect 56 254 57 255
rect 55 254 56 255
rect 54 254 55 255
rect 53 254 54 255
rect 52 254 53 255
rect 51 254 52 255
rect 50 254 51 255
rect 49 254 50 255
rect 48 254 49 255
rect 47 254 48 255
rect 46 254 47 255
rect 45 254 46 255
rect 44 254 45 255
rect 43 254 44 255
rect 38 254 39 255
rect 37 254 38 255
rect 36 254 37 255
rect 35 254 36 255
rect 34 254 35 255
rect 33 254 34 255
rect 32 254 33 255
rect 31 254 32 255
rect 30 254 31 255
rect 29 254 30 255
rect 28 254 29 255
rect 27 254 28 255
rect 26 254 27 255
rect 25 254 26 255
rect 24 254 25 255
rect 23 254 24 255
rect 22 254 23 255
rect 21 254 22 255
rect 20 254 21 255
rect 19 254 20 255
rect 18 254 19 255
rect 17 254 18 255
rect 16 254 17 255
rect 15 254 16 255
rect 142 255 143 256
rect 141 255 142 256
rect 140 255 141 256
rect 139 255 140 256
rect 138 255 139 256
rect 137 255 138 256
rect 136 255 137 256
rect 135 255 136 256
rect 134 255 135 256
rect 133 255 134 256
rect 132 255 133 256
rect 131 255 132 256
rect 130 255 131 256
rect 129 255 130 256
rect 128 255 129 256
rect 127 255 128 256
rect 126 255 127 256
rect 125 255 126 256
rect 124 255 125 256
rect 123 255 124 256
rect 81 255 82 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 69 255 70 256
rect 68 255 69 256
rect 67 255 68 256
rect 66 255 67 256
rect 65 255 66 256
rect 64 255 65 256
rect 53 255 54 256
rect 52 255 53 256
rect 51 255 52 256
rect 50 255 51 256
rect 49 255 50 256
rect 48 255 49 256
rect 47 255 48 256
rect 46 255 47 256
rect 45 255 46 256
rect 44 255 45 256
rect 43 255 44 256
rect 42 255 43 256
rect 35 255 36 256
rect 34 255 35 256
rect 33 255 34 256
rect 32 255 33 256
rect 31 255 32 256
rect 30 255 31 256
rect 29 255 30 256
rect 28 255 29 256
rect 27 255 28 256
rect 26 255 27 256
rect 25 255 26 256
rect 24 255 25 256
rect 23 255 24 256
rect 22 255 23 256
rect 21 255 22 256
rect 20 255 21 256
rect 19 255 20 256
rect 18 255 19 256
rect 17 255 18 256
rect 16 255 17 256
rect 15 255 16 256
rect 140 256 141 257
rect 139 256 140 257
rect 138 256 139 257
rect 137 256 138 257
rect 136 256 137 257
rect 135 256 136 257
rect 134 256 135 257
rect 133 256 134 257
rect 132 256 133 257
rect 131 256 132 257
rect 130 256 131 257
rect 129 256 130 257
rect 128 256 129 257
rect 127 256 128 257
rect 126 256 127 257
rect 81 256 82 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 65 256 66 257
rect 52 256 53 257
rect 51 256 52 257
rect 50 256 51 257
rect 49 256 50 257
rect 48 256 49 257
rect 47 256 48 257
rect 46 256 47 257
rect 45 256 46 257
rect 44 256 45 257
rect 43 256 44 257
rect 42 256 43 257
rect 41 256 42 257
rect 34 256 35 257
rect 33 256 34 257
rect 32 256 33 257
rect 31 256 32 257
rect 30 256 31 257
rect 29 256 30 257
rect 28 256 29 257
rect 27 256 28 257
rect 26 256 27 257
rect 25 256 26 257
rect 24 256 25 257
rect 23 256 24 257
rect 22 256 23 257
rect 21 256 22 257
rect 20 256 21 257
rect 19 256 20 257
rect 18 256 19 257
rect 17 256 18 257
rect 16 256 17 257
rect 15 256 16 257
rect 81 257 82 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 66 257 67 258
rect 51 257 52 258
rect 50 257 51 258
rect 49 257 50 258
rect 48 257 49 258
rect 47 257 48 258
rect 46 257 47 258
rect 45 257 46 258
rect 44 257 45 258
rect 43 257 44 258
rect 42 257 43 258
rect 41 257 42 258
rect 40 257 41 258
rect 32 257 33 258
rect 31 257 32 258
rect 30 257 31 258
rect 29 257 30 258
rect 28 257 29 258
rect 27 257 28 258
rect 26 257 27 258
rect 25 257 26 258
rect 24 257 25 258
rect 23 257 24 258
rect 22 257 23 258
rect 21 257 22 258
rect 20 257 21 258
rect 19 257 20 258
rect 18 257 19 258
rect 17 257 18 258
rect 16 257 17 258
rect 15 257 16 258
rect 14 257 15 258
rect 81 258 82 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 67 258 68 259
rect 50 258 51 259
rect 49 258 50 259
rect 48 258 49 259
rect 47 258 48 259
rect 46 258 47 259
rect 45 258 46 259
rect 44 258 45 259
rect 43 258 44 259
rect 42 258 43 259
rect 41 258 42 259
rect 40 258 41 259
rect 39 258 40 259
rect 31 258 32 259
rect 30 258 31 259
rect 29 258 30 259
rect 28 258 29 259
rect 27 258 28 259
rect 26 258 27 259
rect 25 258 26 259
rect 24 258 25 259
rect 23 258 24 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 16 258 17 259
rect 15 258 16 259
rect 14 258 15 259
rect 81 259 82 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 68 259 69 260
rect 67 259 68 260
rect 50 259 51 260
rect 49 259 50 260
rect 48 259 49 260
rect 47 259 48 260
rect 46 259 47 260
rect 45 259 46 260
rect 44 259 45 260
rect 43 259 44 260
rect 42 259 43 260
rect 41 259 42 260
rect 40 259 41 260
rect 39 259 40 260
rect 30 259 31 260
rect 29 259 30 260
rect 28 259 29 260
rect 27 259 28 260
rect 26 259 27 260
rect 25 259 26 260
rect 24 259 25 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 15 259 16 260
rect 14 259 15 260
rect 81 260 82 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 69 260 70 261
rect 68 260 69 261
rect 67 260 68 261
rect 50 260 51 261
rect 49 260 50 261
rect 48 260 49 261
rect 47 260 48 261
rect 46 260 47 261
rect 45 260 46 261
rect 44 260 45 261
rect 43 260 44 261
rect 42 260 43 261
rect 41 260 42 261
rect 40 260 41 261
rect 39 260 40 261
rect 38 260 39 261
rect 29 260 30 261
rect 28 260 29 261
rect 27 260 28 261
rect 26 260 27 261
rect 25 260 26 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 15 260 16 261
rect 14 260 15 261
rect 81 261 82 262
rect 80 261 81 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 70 261 71 262
rect 69 261 70 262
rect 68 261 69 262
rect 67 261 68 262
rect 50 261 51 262
rect 49 261 50 262
rect 48 261 49 262
rect 47 261 48 262
rect 46 261 47 262
rect 45 261 46 262
rect 44 261 45 262
rect 43 261 44 262
rect 42 261 43 262
rect 41 261 42 262
rect 40 261 41 262
rect 39 261 40 262
rect 38 261 39 262
rect 29 261 30 262
rect 28 261 29 262
rect 27 261 28 262
rect 26 261 27 262
rect 25 261 26 262
rect 24 261 25 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 15 261 16 262
rect 14 261 15 262
rect 134 262 135 263
rect 133 262 134 263
rect 132 262 133 263
rect 131 262 132 263
rect 130 262 131 263
rect 129 262 130 263
rect 128 262 129 263
rect 127 262 128 263
rect 126 262 127 263
rect 81 262 82 263
rect 80 262 81 263
rect 79 262 80 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 71 262 72 263
rect 70 262 71 263
rect 69 262 70 263
rect 68 262 69 263
rect 67 262 68 263
rect 50 262 51 263
rect 49 262 50 263
rect 48 262 49 263
rect 47 262 48 263
rect 46 262 47 263
rect 45 262 46 263
rect 44 262 45 263
rect 43 262 44 263
rect 42 262 43 263
rect 41 262 42 263
rect 40 262 41 263
rect 39 262 40 263
rect 38 262 39 263
rect 28 262 29 263
rect 27 262 28 263
rect 26 262 27 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 15 262 16 263
rect 14 262 15 263
rect 13 262 14 263
rect 136 263 137 264
rect 135 263 136 264
rect 134 263 135 264
rect 133 263 134 264
rect 132 263 133 264
rect 131 263 132 264
rect 130 263 131 264
rect 129 263 130 264
rect 128 263 129 264
rect 127 263 128 264
rect 126 263 127 264
rect 125 263 126 264
rect 124 263 125 264
rect 81 263 82 264
rect 80 263 81 264
rect 79 263 80 264
rect 78 263 79 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 72 263 73 264
rect 71 263 72 264
rect 70 263 71 264
rect 69 263 70 264
rect 68 263 69 264
rect 67 263 68 264
rect 66 263 67 264
rect 51 263 52 264
rect 50 263 51 264
rect 49 263 50 264
rect 48 263 49 264
rect 47 263 48 264
rect 46 263 47 264
rect 45 263 46 264
rect 44 263 45 264
rect 43 263 44 264
rect 42 263 43 264
rect 41 263 42 264
rect 40 263 41 264
rect 39 263 40 264
rect 38 263 39 264
rect 37 263 38 264
rect 28 263 29 264
rect 27 263 28 264
rect 26 263 27 264
rect 25 263 26 264
rect 24 263 25 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 16 263 17 264
rect 15 263 16 264
rect 14 263 15 264
rect 13 263 14 264
rect 138 264 139 265
rect 137 264 138 265
rect 136 264 137 265
rect 135 264 136 265
rect 134 264 135 265
rect 133 264 134 265
rect 132 264 133 265
rect 131 264 132 265
rect 130 264 131 265
rect 129 264 130 265
rect 128 264 129 265
rect 127 264 128 265
rect 126 264 127 265
rect 125 264 126 265
rect 124 264 125 265
rect 123 264 124 265
rect 122 264 123 265
rect 81 264 82 265
rect 80 264 81 265
rect 79 264 80 265
rect 78 264 79 265
rect 77 264 78 265
rect 76 264 77 265
rect 75 264 76 265
rect 74 264 75 265
rect 73 264 74 265
rect 72 264 73 265
rect 71 264 72 265
rect 70 264 71 265
rect 69 264 70 265
rect 68 264 69 265
rect 67 264 68 265
rect 66 264 67 265
rect 65 264 66 265
rect 52 264 53 265
rect 51 264 52 265
rect 50 264 51 265
rect 49 264 50 265
rect 48 264 49 265
rect 47 264 48 265
rect 46 264 47 265
rect 45 264 46 265
rect 44 264 45 265
rect 43 264 44 265
rect 42 264 43 265
rect 41 264 42 265
rect 40 264 41 265
rect 39 264 40 265
rect 38 264 39 265
rect 37 264 38 265
rect 28 264 29 265
rect 27 264 28 265
rect 26 264 27 265
rect 25 264 26 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 16 264 17 265
rect 15 264 16 265
rect 14 264 15 265
rect 13 264 14 265
rect 139 265 140 266
rect 138 265 139 266
rect 137 265 138 266
rect 136 265 137 266
rect 135 265 136 266
rect 134 265 135 266
rect 133 265 134 266
rect 132 265 133 266
rect 131 265 132 266
rect 130 265 131 266
rect 129 265 130 266
rect 128 265 129 266
rect 127 265 128 266
rect 126 265 127 266
rect 125 265 126 266
rect 124 265 125 266
rect 123 265 124 266
rect 122 265 123 266
rect 121 265 122 266
rect 80 265 81 266
rect 79 265 80 266
rect 78 265 79 266
rect 77 265 78 266
rect 76 265 77 266
rect 75 265 76 266
rect 74 265 75 266
rect 73 265 74 266
rect 72 265 73 266
rect 71 265 72 266
rect 70 265 71 266
rect 69 265 70 266
rect 68 265 69 266
rect 67 265 68 266
rect 66 265 67 266
rect 65 265 66 266
rect 64 265 65 266
rect 63 265 64 266
rect 54 265 55 266
rect 53 265 54 266
rect 52 265 53 266
rect 51 265 52 266
rect 50 265 51 266
rect 49 265 50 266
rect 48 265 49 266
rect 47 265 48 266
rect 46 265 47 266
rect 45 265 46 266
rect 44 265 45 266
rect 43 265 44 266
rect 42 265 43 266
rect 41 265 42 266
rect 40 265 41 266
rect 39 265 40 266
rect 38 265 39 266
rect 37 265 38 266
rect 27 265 28 266
rect 26 265 27 266
rect 25 265 26 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 18 265 19 266
rect 17 265 18 266
rect 16 265 17 266
rect 15 265 16 266
rect 14 265 15 266
rect 13 265 14 266
rect 139 266 140 267
rect 138 266 139 267
rect 137 266 138 267
rect 136 266 137 267
rect 135 266 136 267
rect 134 266 135 267
rect 133 266 134 267
rect 132 266 133 267
rect 131 266 132 267
rect 130 266 131 267
rect 129 266 130 267
rect 128 266 129 267
rect 127 266 128 267
rect 126 266 127 267
rect 125 266 126 267
rect 124 266 125 267
rect 123 266 124 267
rect 122 266 123 267
rect 121 266 122 267
rect 120 266 121 267
rect 80 266 81 267
rect 79 266 80 267
rect 78 266 79 267
rect 77 266 78 267
rect 76 266 77 267
rect 75 266 76 267
rect 74 266 75 267
rect 73 266 74 267
rect 72 266 73 267
rect 71 266 72 267
rect 70 266 71 267
rect 69 266 70 267
rect 68 266 69 267
rect 67 266 68 267
rect 66 266 67 267
rect 65 266 66 267
rect 64 266 65 267
rect 63 266 64 267
rect 62 266 63 267
rect 61 266 62 267
rect 60 266 61 267
rect 59 266 60 267
rect 58 266 59 267
rect 57 266 58 267
rect 56 266 57 267
rect 55 266 56 267
rect 54 266 55 267
rect 53 266 54 267
rect 52 266 53 267
rect 51 266 52 267
rect 50 266 51 267
rect 49 266 50 267
rect 48 266 49 267
rect 47 266 48 267
rect 46 266 47 267
rect 45 266 46 267
rect 44 266 45 267
rect 43 266 44 267
rect 42 266 43 267
rect 41 266 42 267
rect 40 266 41 267
rect 39 266 40 267
rect 38 266 39 267
rect 37 266 38 267
rect 27 266 28 267
rect 26 266 27 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 16 266 17 267
rect 15 266 16 267
rect 14 266 15 267
rect 13 266 14 267
rect 140 267 141 268
rect 139 267 140 268
rect 138 267 139 268
rect 137 267 138 268
rect 136 267 137 268
rect 135 267 136 268
rect 134 267 135 268
rect 133 267 134 268
rect 132 267 133 268
rect 131 267 132 268
rect 130 267 131 268
rect 129 267 130 268
rect 128 267 129 268
rect 127 267 128 268
rect 126 267 127 268
rect 125 267 126 268
rect 124 267 125 268
rect 123 267 124 268
rect 122 267 123 268
rect 121 267 122 268
rect 120 267 121 268
rect 119 267 120 268
rect 80 267 81 268
rect 79 267 80 268
rect 78 267 79 268
rect 77 267 78 268
rect 76 267 77 268
rect 75 267 76 268
rect 74 267 75 268
rect 73 267 74 268
rect 72 267 73 268
rect 71 267 72 268
rect 70 267 71 268
rect 69 267 70 268
rect 68 267 69 268
rect 67 267 68 268
rect 66 267 67 268
rect 65 267 66 268
rect 64 267 65 268
rect 63 267 64 268
rect 62 267 63 268
rect 61 267 62 268
rect 60 267 61 268
rect 59 267 60 268
rect 58 267 59 268
rect 57 267 58 268
rect 56 267 57 268
rect 55 267 56 268
rect 54 267 55 268
rect 53 267 54 268
rect 52 267 53 268
rect 51 267 52 268
rect 50 267 51 268
rect 49 267 50 268
rect 48 267 49 268
rect 47 267 48 268
rect 46 267 47 268
rect 45 267 46 268
rect 44 267 45 268
rect 43 267 44 268
rect 42 267 43 268
rect 41 267 42 268
rect 40 267 41 268
rect 39 267 40 268
rect 38 267 39 268
rect 37 267 38 268
rect 27 267 28 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 14 267 15 268
rect 13 267 14 268
rect 141 268 142 269
rect 140 268 141 269
rect 139 268 140 269
rect 138 268 139 269
rect 137 268 138 269
rect 136 268 137 269
rect 135 268 136 269
rect 134 268 135 269
rect 133 268 134 269
rect 126 268 127 269
rect 125 268 126 269
rect 124 268 125 269
rect 123 268 124 269
rect 122 268 123 269
rect 121 268 122 269
rect 120 268 121 269
rect 119 268 120 269
rect 80 268 81 269
rect 79 268 80 269
rect 78 268 79 269
rect 77 268 78 269
rect 76 268 77 269
rect 75 268 76 269
rect 74 268 75 269
rect 73 268 74 269
rect 72 268 73 269
rect 71 268 72 269
rect 70 268 71 269
rect 69 268 70 269
rect 68 268 69 269
rect 67 268 68 269
rect 66 268 67 269
rect 65 268 66 269
rect 64 268 65 269
rect 63 268 64 269
rect 62 268 63 269
rect 61 268 62 269
rect 60 268 61 269
rect 59 268 60 269
rect 58 268 59 269
rect 57 268 58 269
rect 56 268 57 269
rect 55 268 56 269
rect 54 268 55 269
rect 53 268 54 269
rect 52 268 53 269
rect 51 268 52 269
rect 50 268 51 269
rect 49 268 50 269
rect 48 268 49 269
rect 47 268 48 269
rect 46 268 47 269
rect 45 268 46 269
rect 44 268 45 269
rect 43 268 44 269
rect 42 268 43 269
rect 41 268 42 269
rect 40 268 41 269
rect 39 268 40 269
rect 38 268 39 269
rect 37 268 38 269
rect 27 268 28 269
rect 26 268 27 269
rect 25 268 26 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 14 268 15 269
rect 13 268 14 269
rect 141 269 142 270
rect 140 269 141 270
rect 139 269 140 270
rect 138 269 139 270
rect 137 269 138 270
rect 136 269 137 270
rect 135 269 136 270
rect 124 269 125 270
rect 123 269 124 270
rect 122 269 123 270
rect 121 269 122 270
rect 120 269 121 270
rect 119 269 120 270
rect 118 269 119 270
rect 79 269 80 270
rect 78 269 79 270
rect 77 269 78 270
rect 76 269 77 270
rect 75 269 76 270
rect 74 269 75 270
rect 73 269 74 270
rect 72 269 73 270
rect 71 269 72 270
rect 70 269 71 270
rect 69 269 70 270
rect 68 269 69 270
rect 67 269 68 270
rect 66 269 67 270
rect 65 269 66 270
rect 64 269 65 270
rect 63 269 64 270
rect 62 269 63 270
rect 61 269 62 270
rect 60 269 61 270
rect 59 269 60 270
rect 58 269 59 270
rect 57 269 58 270
rect 56 269 57 270
rect 55 269 56 270
rect 54 269 55 270
rect 53 269 54 270
rect 52 269 53 270
rect 51 269 52 270
rect 50 269 51 270
rect 49 269 50 270
rect 48 269 49 270
rect 47 269 48 270
rect 46 269 47 270
rect 45 269 46 270
rect 44 269 45 270
rect 43 269 44 270
rect 42 269 43 270
rect 41 269 42 270
rect 40 269 41 270
rect 39 269 40 270
rect 38 269 39 270
rect 37 269 38 270
rect 27 269 28 270
rect 26 269 27 270
rect 25 269 26 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 16 269 17 270
rect 15 269 16 270
rect 14 269 15 270
rect 13 269 14 270
rect 141 270 142 271
rect 140 270 141 271
rect 139 270 140 271
rect 138 270 139 271
rect 137 270 138 271
rect 136 270 137 271
rect 123 270 124 271
rect 122 270 123 271
rect 121 270 122 271
rect 120 270 121 271
rect 119 270 120 271
rect 118 270 119 271
rect 79 270 80 271
rect 78 270 79 271
rect 77 270 78 271
rect 76 270 77 271
rect 75 270 76 271
rect 74 270 75 271
rect 73 270 74 271
rect 72 270 73 271
rect 71 270 72 271
rect 70 270 71 271
rect 69 270 70 271
rect 68 270 69 271
rect 67 270 68 271
rect 66 270 67 271
rect 65 270 66 271
rect 64 270 65 271
rect 63 270 64 271
rect 62 270 63 271
rect 61 270 62 271
rect 60 270 61 271
rect 59 270 60 271
rect 58 270 59 271
rect 57 270 58 271
rect 56 270 57 271
rect 55 270 56 271
rect 54 270 55 271
rect 53 270 54 271
rect 52 270 53 271
rect 51 270 52 271
rect 50 270 51 271
rect 49 270 50 271
rect 48 270 49 271
rect 47 270 48 271
rect 46 270 47 271
rect 45 270 46 271
rect 44 270 45 271
rect 43 270 44 271
rect 42 270 43 271
rect 41 270 42 271
rect 40 270 41 271
rect 39 270 40 271
rect 38 270 39 271
rect 37 270 38 271
rect 27 270 28 271
rect 26 270 27 271
rect 25 270 26 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 15 270 16 271
rect 14 270 15 271
rect 13 270 14 271
rect 142 271 143 272
rect 141 271 142 272
rect 140 271 141 272
rect 139 271 140 272
rect 138 271 139 272
rect 137 271 138 272
rect 122 271 123 272
rect 121 271 122 272
rect 120 271 121 272
rect 119 271 120 272
rect 118 271 119 272
rect 79 271 80 272
rect 78 271 79 272
rect 77 271 78 272
rect 76 271 77 272
rect 75 271 76 272
rect 74 271 75 272
rect 73 271 74 272
rect 72 271 73 272
rect 71 271 72 272
rect 70 271 71 272
rect 69 271 70 272
rect 68 271 69 272
rect 67 271 68 272
rect 66 271 67 272
rect 65 271 66 272
rect 64 271 65 272
rect 63 271 64 272
rect 62 271 63 272
rect 61 271 62 272
rect 60 271 61 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 55 271 56 272
rect 54 271 55 272
rect 53 271 54 272
rect 52 271 53 272
rect 51 271 52 272
rect 50 271 51 272
rect 49 271 50 272
rect 48 271 49 272
rect 47 271 48 272
rect 46 271 47 272
rect 45 271 46 272
rect 44 271 45 272
rect 43 271 44 272
rect 42 271 43 272
rect 41 271 42 272
rect 40 271 41 272
rect 39 271 40 272
rect 38 271 39 272
rect 37 271 38 272
rect 27 271 28 272
rect 26 271 27 272
rect 25 271 26 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 15 271 16 272
rect 14 271 15 272
rect 13 271 14 272
rect 142 272 143 273
rect 141 272 142 273
rect 140 272 141 273
rect 139 272 140 273
rect 138 272 139 273
rect 122 272 123 273
rect 121 272 122 273
rect 120 272 121 273
rect 119 272 120 273
rect 118 272 119 273
rect 117 272 118 273
rect 78 272 79 273
rect 77 272 78 273
rect 76 272 77 273
rect 75 272 76 273
rect 74 272 75 273
rect 73 272 74 273
rect 72 272 73 273
rect 71 272 72 273
rect 70 272 71 273
rect 69 272 70 273
rect 68 272 69 273
rect 67 272 68 273
rect 66 272 67 273
rect 65 272 66 273
rect 64 272 65 273
rect 63 272 64 273
rect 62 272 63 273
rect 61 272 62 273
rect 60 272 61 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 55 272 56 273
rect 54 272 55 273
rect 53 272 54 273
rect 52 272 53 273
rect 51 272 52 273
rect 50 272 51 273
rect 49 272 50 273
rect 48 272 49 273
rect 47 272 48 273
rect 46 272 47 273
rect 45 272 46 273
rect 44 272 45 273
rect 43 272 44 273
rect 42 272 43 273
rect 41 272 42 273
rect 40 272 41 273
rect 39 272 40 273
rect 38 272 39 273
rect 27 272 28 273
rect 26 272 27 273
rect 25 272 26 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 15 272 16 273
rect 14 272 15 273
rect 13 272 14 273
rect 142 273 143 274
rect 141 273 142 274
rect 140 273 141 274
rect 139 273 140 274
rect 138 273 139 274
rect 121 273 122 274
rect 120 273 121 274
rect 119 273 120 274
rect 118 273 119 274
rect 117 273 118 274
rect 78 273 79 274
rect 77 273 78 274
rect 76 273 77 274
rect 75 273 76 274
rect 74 273 75 274
rect 73 273 74 274
rect 72 273 73 274
rect 71 273 72 274
rect 70 273 71 274
rect 69 273 70 274
rect 68 273 69 274
rect 67 273 68 274
rect 66 273 67 274
rect 65 273 66 274
rect 64 273 65 274
rect 63 273 64 274
rect 62 273 63 274
rect 61 273 62 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 55 273 56 274
rect 54 273 55 274
rect 53 273 54 274
rect 52 273 53 274
rect 51 273 52 274
rect 50 273 51 274
rect 49 273 50 274
rect 48 273 49 274
rect 47 273 48 274
rect 46 273 47 274
rect 45 273 46 274
rect 44 273 45 274
rect 43 273 44 274
rect 42 273 43 274
rect 41 273 42 274
rect 40 273 41 274
rect 39 273 40 274
rect 38 273 39 274
rect 27 273 28 274
rect 26 273 27 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 15 273 16 274
rect 14 273 15 274
rect 13 273 14 274
rect 142 274 143 275
rect 141 274 142 275
rect 140 274 141 275
rect 139 274 140 275
rect 138 274 139 275
rect 132 274 133 275
rect 131 274 132 275
rect 130 274 131 275
rect 129 274 130 275
rect 128 274 129 275
rect 121 274 122 275
rect 120 274 121 275
rect 119 274 120 275
rect 118 274 119 275
rect 117 274 118 275
rect 77 274 78 275
rect 76 274 77 275
rect 75 274 76 275
rect 74 274 75 275
rect 73 274 74 275
rect 72 274 73 275
rect 71 274 72 275
rect 70 274 71 275
rect 69 274 70 275
rect 68 274 69 275
rect 67 274 68 275
rect 66 274 67 275
rect 65 274 66 275
rect 64 274 65 275
rect 63 274 64 275
rect 62 274 63 275
rect 61 274 62 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 55 274 56 275
rect 54 274 55 275
rect 53 274 54 275
rect 52 274 53 275
rect 51 274 52 275
rect 50 274 51 275
rect 49 274 50 275
rect 48 274 49 275
rect 47 274 48 275
rect 46 274 47 275
rect 45 274 46 275
rect 44 274 45 275
rect 43 274 44 275
rect 42 274 43 275
rect 41 274 42 275
rect 40 274 41 275
rect 39 274 40 275
rect 38 274 39 275
rect 27 274 28 275
rect 26 274 27 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 16 274 17 275
rect 15 274 16 275
rect 14 274 15 275
rect 13 274 14 275
rect 142 275 143 276
rect 141 275 142 276
rect 140 275 141 276
rect 139 275 140 276
rect 138 275 139 276
rect 132 275 133 276
rect 131 275 132 276
rect 130 275 131 276
rect 129 275 130 276
rect 128 275 129 276
rect 121 275 122 276
rect 120 275 121 276
rect 119 275 120 276
rect 118 275 119 276
rect 117 275 118 276
rect 76 275 77 276
rect 75 275 76 276
rect 74 275 75 276
rect 73 275 74 276
rect 72 275 73 276
rect 71 275 72 276
rect 70 275 71 276
rect 69 275 70 276
rect 68 275 69 276
rect 67 275 68 276
rect 66 275 67 276
rect 65 275 66 276
rect 64 275 65 276
rect 63 275 64 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 56 275 57 276
rect 55 275 56 276
rect 54 275 55 276
rect 53 275 54 276
rect 52 275 53 276
rect 51 275 52 276
rect 50 275 51 276
rect 49 275 50 276
rect 48 275 49 276
rect 47 275 48 276
rect 46 275 47 276
rect 45 275 46 276
rect 44 275 45 276
rect 43 275 44 276
rect 42 275 43 276
rect 41 275 42 276
rect 40 275 41 276
rect 39 275 40 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 17 275 18 276
rect 16 275 17 276
rect 15 275 16 276
rect 14 275 15 276
rect 142 276 143 277
rect 141 276 142 277
rect 140 276 141 277
rect 139 276 140 277
rect 138 276 139 277
rect 132 276 133 277
rect 131 276 132 277
rect 130 276 131 277
rect 129 276 130 277
rect 128 276 129 277
rect 121 276 122 277
rect 120 276 121 277
rect 119 276 120 277
rect 118 276 119 277
rect 117 276 118 277
rect 76 276 77 277
rect 75 276 76 277
rect 74 276 75 277
rect 73 276 74 277
rect 72 276 73 277
rect 71 276 72 277
rect 70 276 71 277
rect 69 276 70 277
rect 68 276 69 277
rect 67 276 68 277
rect 66 276 67 277
rect 65 276 66 277
rect 64 276 65 277
rect 63 276 64 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 56 276 57 277
rect 55 276 56 277
rect 54 276 55 277
rect 53 276 54 277
rect 52 276 53 277
rect 51 276 52 277
rect 50 276 51 277
rect 49 276 50 277
rect 48 276 49 277
rect 47 276 48 277
rect 46 276 47 277
rect 45 276 46 277
rect 44 276 45 277
rect 43 276 44 277
rect 42 276 43 277
rect 41 276 42 277
rect 40 276 41 277
rect 39 276 40 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 18 276 19 277
rect 17 276 18 277
rect 16 276 17 277
rect 15 276 16 277
rect 14 276 15 277
rect 142 277 143 278
rect 141 277 142 278
rect 140 277 141 278
rect 139 277 140 278
rect 138 277 139 278
rect 132 277 133 278
rect 131 277 132 278
rect 130 277 131 278
rect 129 277 130 278
rect 128 277 129 278
rect 121 277 122 278
rect 120 277 121 278
rect 119 277 120 278
rect 118 277 119 278
rect 117 277 118 278
rect 75 277 76 278
rect 74 277 75 278
rect 73 277 74 278
rect 72 277 73 278
rect 71 277 72 278
rect 70 277 71 278
rect 69 277 70 278
rect 68 277 69 278
rect 67 277 68 278
rect 66 277 67 278
rect 65 277 66 278
rect 64 277 65 278
rect 63 277 64 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 56 277 57 278
rect 55 277 56 278
rect 54 277 55 278
rect 53 277 54 278
rect 52 277 53 278
rect 51 277 52 278
rect 50 277 51 278
rect 49 277 50 278
rect 48 277 49 278
rect 47 277 48 278
rect 46 277 47 278
rect 45 277 46 278
rect 44 277 45 278
rect 43 277 44 278
rect 42 277 43 278
rect 41 277 42 278
rect 40 277 41 278
rect 28 277 29 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 19 277 20 278
rect 18 277 19 278
rect 17 277 18 278
rect 16 277 17 278
rect 15 277 16 278
rect 14 277 15 278
rect 142 278 143 279
rect 141 278 142 279
rect 140 278 141 279
rect 139 278 140 279
rect 138 278 139 279
rect 132 278 133 279
rect 131 278 132 279
rect 130 278 131 279
rect 129 278 130 279
rect 128 278 129 279
rect 121 278 122 279
rect 120 278 121 279
rect 119 278 120 279
rect 118 278 119 279
rect 117 278 118 279
rect 74 278 75 279
rect 73 278 74 279
rect 72 278 73 279
rect 71 278 72 279
rect 70 278 71 279
rect 69 278 70 279
rect 68 278 69 279
rect 67 278 68 279
rect 66 278 67 279
rect 65 278 66 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 57 278 58 279
rect 56 278 57 279
rect 55 278 56 279
rect 54 278 55 279
rect 53 278 54 279
rect 52 278 53 279
rect 51 278 52 279
rect 50 278 51 279
rect 49 278 50 279
rect 48 278 49 279
rect 47 278 48 279
rect 46 278 47 279
rect 45 278 46 279
rect 44 278 45 279
rect 43 278 44 279
rect 42 278 43 279
rect 41 278 42 279
rect 28 278 29 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 17 278 18 279
rect 16 278 17 279
rect 15 278 16 279
rect 14 278 15 279
rect 142 279 143 280
rect 141 279 142 280
rect 140 279 141 280
rect 139 279 140 280
rect 138 279 139 280
rect 137 279 138 280
rect 136 279 137 280
rect 135 279 136 280
rect 134 279 135 280
rect 133 279 134 280
rect 132 279 133 280
rect 131 279 132 280
rect 130 279 131 280
rect 129 279 130 280
rect 128 279 129 280
rect 121 279 122 280
rect 120 279 121 280
rect 119 279 120 280
rect 118 279 119 280
rect 117 279 118 280
rect 73 279 74 280
rect 72 279 73 280
rect 71 279 72 280
rect 70 279 71 280
rect 69 279 70 280
rect 68 279 69 280
rect 67 279 68 280
rect 66 279 67 280
rect 65 279 66 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 58 279 59 280
rect 57 279 58 280
rect 56 279 57 280
rect 55 279 56 280
rect 54 279 55 280
rect 53 279 54 280
rect 52 279 53 280
rect 51 279 52 280
rect 50 279 51 280
rect 49 279 50 280
rect 48 279 49 280
rect 47 279 48 280
rect 46 279 47 280
rect 45 279 46 280
rect 44 279 45 280
rect 43 279 44 280
rect 42 279 43 280
rect 28 279 29 280
rect 27 279 28 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 17 279 18 280
rect 16 279 17 280
rect 15 279 16 280
rect 141 280 142 281
rect 140 280 141 281
rect 139 280 140 281
rect 138 280 139 281
rect 137 280 138 281
rect 136 280 137 281
rect 135 280 136 281
rect 134 280 135 281
rect 133 280 134 281
rect 132 280 133 281
rect 131 280 132 281
rect 130 280 131 281
rect 129 280 130 281
rect 128 280 129 281
rect 121 280 122 281
rect 120 280 121 281
rect 119 280 120 281
rect 118 280 119 281
rect 117 280 118 281
rect 71 280 72 281
rect 70 280 71 281
rect 69 280 70 281
rect 68 280 69 281
rect 67 280 68 281
rect 66 280 67 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 59 280 60 281
rect 58 280 59 281
rect 57 280 58 281
rect 56 280 57 281
rect 55 280 56 281
rect 54 280 55 281
rect 53 280 54 281
rect 52 280 53 281
rect 51 280 52 281
rect 50 280 51 281
rect 49 280 50 281
rect 48 280 49 281
rect 47 280 48 281
rect 46 280 47 281
rect 45 280 46 281
rect 44 280 45 281
rect 43 280 44 281
rect 141 281 142 282
rect 140 281 141 282
rect 139 281 140 282
rect 138 281 139 282
rect 137 281 138 282
rect 136 281 137 282
rect 135 281 136 282
rect 134 281 135 282
rect 133 281 134 282
rect 132 281 133 282
rect 131 281 132 282
rect 130 281 131 282
rect 129 281 130 282
rect 128 281 129 282
rect 122 281 123 282
rect 121 281 122 282
rect 120 281 121 282
rect 119 281 120 282
rect 118 281 119 282
rect 70 281 71 282
rect 69 281 70 282
rect 68 281 69 282
rect 67 281 68 282
rect 66 281 67 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 60 281 61 282
rect 59 281 60 282
rect 58 281 59 282
rect 57 281 58 282
rect 56 281 57 282
rect 55 281 56 282
rect 54 281 55 282
rect 53 281 54 282
rect 52 281 53 282
rect 51 281 52 282
rect 50 281 51 282
rect 49 281 50 282
rect 48 281 49 282
rect 47 281 48 282
rect 46 281 47 282
rect 45 281 46 282
rect 44 281 45 282
rect 141 282 142 283
rect 140 282 141 283
rect 139 282 140 283
rect 138 282 139 283
rect 137 282 138 283
rect 136 282 137 283
rect 135 282 136 283
rect 134 282 135 283
rect 133 282 134 283
rect 132 282 133 283
rect 131 282 132 283
rect 130 282 131 283
rect 129 282 130 283
rect 128 282 129 283
rect 122 282 123 283
rect 121 282 122 283
rect 120 282 121 283
rect 119 282 120 283
rect 118 282 119 283
rect 68 282 69 283
rect 67 282 68 283
rect 66 282 67 283
rect 65 282 66 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 61 282 62 283
rect 60 282 61 283
rect 59 282 60 283
rect 58 282 59 283
rect 57 282 58 283
rect 56 282 57 283
rect 55 282 56 283
rect 54 282 55 283
rect 53 282 54 283
rect 52 282 53 283
rect 51 282 52 283
rect 50 282 51 283
rect 49 282 50 283
rect 48 282 49 283
rect 47 282 48 283
rect 46 282 47 283
rect 140 283 141 284
rect 139 283 140 284
rect 138 283 139 284
rect 137 283 138 284
rect 136 283 137 284
rect 135 283 136 284
rect 134 283 135 284
rect 133 283 134 284
rect 132 283 133 284
rect 131 283 132 284
rect 130 283 131 284
rect 129 283 130 284
rect 128 283 129 284
rect 66 283 67 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 62 283 63 284
rect 61 283 62 284
rect 60 283 61 284
rect 59 283 60 284
rect 58 283 59 284
rect 57 283 58 284
rect 56 283 57 284
rect 55 283 56 284
rect 54 283 55 284
rect 53 283 54 284
rect 52 283 53 284
rect 51 283 52 284
rect 50 283 51 284
rect 49 283 50 284
rect 48 283 49 284
rect 140 284 141 285
rect 139 284 140 285
rect 138 284 139 285
rect 137 284 138 285
rect 136 284 137 285
rect 135 284 136 285
rect 134 284 135 285
rect 133 284 134 285
rect 132 284 133 285
rect 131 284 132 285
rect 130 284 131 285
rect 129 284 130 285
rect 128 284 129 285
rect 62 284 63 285
rect 61 284 62 285
rect 60 284 61 285
rect 59 284 60 285
rect 58 284 59 285
rect 57 284 58 285
rect 56 284 57 285
rect 55 284 56 285
rect 54 284 55 285
rect 53 284 54 285
rect 52 284 53 285
rect 134 288 135 289
rect 133 288 134 289
rect 132 288 133 289
rect 137 289 138 290
rect 136 289 137 290
rect 135 289 136 290
rect 134 289 135 290
rect 133 289 134 290
rect 132 289 133 290
rect 131 289 132 290
rect 130 289 131 290
rect 129 289 130 290
rect 139 290 140 291
rect 138 290 139 291
rect 137 290 138 291
rect 136 290 137 291
rect 135 290 136 291
rect 134 290 135 291
rect 133 290 134 291
rect 132 290 133 291
rect 131 290 132 291
rect 130 290 131 291
rect 129 290 130 291
rect 128 290 129 291
rect 127 290 128 291
rect 140 291 141 292
rect 139 291 140 292
rect 138 291 139 292
rect 137 291 138 292
rect 136 291 137 292
rect 135 291 136 292
rect 134 291 135 292
rect 133 291 134 292
rect 132 291 133 292
rect 131 291 132 292
rect 130 291 131 292
rect 129 291 130 292
rect 128 291 129 292
rect 127 291 128 292
rect 126 291 127 292
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 135 292 136 293
rect 134 292 135 293
rect 133 292 134 293
rect 132 292 133 293
rect 131 292 132 293
rect 130 292 131 293
rect 129 292 130 293
rect 128 292 129 293
rect 127 292 128 293
rect 126 292 127 293
rect 125 292 126 293
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 136 293 137 294
rect 135 293 136 294
rect 134 293 135 294
rect 133 293 134 294
rect 132 293 133 294
rect 131 293 132 294
rect 130 293 131 294
rect 129 293 130 294
rect 128 293 129 294
rect 127 293 128 294
rect 126 293 127 294
rect 125 293 126 294
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 137 294 138 295
rect 136 294 137 295
rect 130 294 131 295
rect 129 294 130 295
rect 128 294 129 295
rect 127 294 128 295
rect 126 294 127 295
rect 125 294 126 295
rect 79 294 80 295
rect 78 294 79 295
rect 77 294 78 295
rect 76 294 77 295
rect 75 294 76 295
rect 74 294 75 295
rect 73 294 74 295
rect 72 294 73 295
rect 71 294 72 295
rect 70 294 71 295
rect 69 294 70 295
rect 68 294 69 295
rect 67 294 68 295
rect 66 294 67 295
rect 65 294 66 295
rect 64 294 65 295
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 138 295 139 296
rect 128 295 129 296
rect 127 295 128 296
rect 126 295 127 296
rect 125 295 126 296
rect 124 295 125 296
rect 79 295 80 296
rect 78 295 79 296
rect 77 295 78 296
rect 76 295 77 296
rect 75 295 76 296
rect 74 295 75 296
rect 73 295 74 296
rect 72 295 73 296
rect 71 295 72 296
rect 70 295 71 296
rect 69 295 70 296
rect 68 295 69 296
rect 67 295 68 296
rect 66 295 67 296
rect 65 295 66 296
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 139 296 140 297
rect 138 296 139 297
rect 128 296 129 297
rect 127 296 128 297
rect 126 296 127 297
rect 125 296 126 297
rect 124 296 125 297
rect 79 296 80 297
rect 78 296 79 297
rect 77 296 78 297
rect 76 296 77 297
rect 75 296 76 297
rect 74 296 75 297
rect 73 296 74 297
rect 72 296 73 297
rect 71 296 72 297
rect 70 296 71 297
rect 69 296 70 297
rect 68 296 69 297
rect 67 296 68 297
rect 66 296 67 297
rect 65 296 66 297
rect 53 296 54 297
rect 52 296 53 297
rect 51 296 52 297
rect 50 296 51 297
rect 49 296 50 297
rect 48 296 49 297
rect 47 296 48 297
rect 46 296 47 297
rect 45 296 46 297
rect 44 296 45 297
rect 43 296 44 297
rect 42 296 43 297
rect 41 296 42 297
rect 40 296 41 297
rect 39 296 40 297
rect 38 296 39 297
rect 142 297 143 298
rect 141 297 142 298
rect 140 297 141 298
rect 139 297 140 298
rect 127 297 128 298
rect 126 297 127 298
rect 125 297 126 298
rect 124 297 125 298
rect 79 297 80 298
rect 78 297 79 298
rect 77 297 78 298
rect 76 297 77 298
rect 75 297 76 298
rect 74 297 75 298
rect 73 297 74 298
rect 72 297 73 298
rect 71 297 72 298
rect 70 297 71 298
rect 69 297 70 298
rect 68 297 69 298
rect 67 297 68 298
rect 66 297 67 298
rect 65 297 66 298
rect 53 297 54 298
rect 52 297 53 298
rect 51 297 52 298
rect 50 297 51 298
rect 49 297 50 298
rect 48 297 49 298
rect 47 297 48 298
rect 46 297 47 298
rect 45 297 46 298
rect 44 297 45 298
rect 43 297 44 298
rect 42 297 43 298
rect 41 297 42 298
rect 40 297 41 298
rect 39 297 40 298
rect 38 297 39 298
rect 37 297 38 298
rect 36 297 37 298
rect 35 297 36 298
rect 34 297 35 298
rect 33 297 34 298
rect 32 297 33 298
rect 31 297 32 298
rect 30 297 31 298
rect 29 297 30 298
rect 28 297 29 298
rect 27 297 28 298
rect 26 297 27 298
rect 25 297 26 298
rect 24 297 25 298
rect 23 297 24 298
rect 22 297 23 298
rect 142 298 143 299
rect 141 298 142 299
rect 140 298 141 299
rect 139 298 140 299
rect 127 298 128 299
rect 126 298 127 299
rect 125 298 126 299
rect 124 298 125 299
rect 80 298 81 299
rect 79 298 80 299
rect 78 298 79 299
rect 77 298 78 299
rect 76 298 77 299
rect 75 298 76 299
rect 74 298 75 299
rect 73 298 74 299
rect 72 298 73 299
rect 71 298 72 299
rect 70 298 71 299
rect 69 298 70 299
rect 68 298 69 299
rect 67 298 68 299
rect 66 298 67 299
rect 52 298 53 299
rect 51 298 52 299
rect 50 298 51 299
rect 49 298 50 299
rect 48 298 49 299
rect 47 298 48 299
rect 46 298 47 299
rect 45 298 46 299
rect 44 298 45 299
rect 43 298 44 299
rect 42 298 43 299
rect 41 298 42 299
rect 40 298 41 299
rect 39 298 40 299
rect 38 298 39 299
rect 37 298 38 299
rect 36 298 37 299
rect 35 298 36 299
rect 34 298 35 299
rect 33 298 34 299
rect 32 298 33 299
rect 31 298 32 299
rect 30 298 31 299
rect 29 298 30 299
rect 28 298 29 299
rect 27 298 28 299
rect 26 298 27 299
rect 25 298 26 299
rect 24 298 25 299
rect 23 298 24 299
rect 22 298 23 299
rect 21 298 22 299
rect 20 298 21 299
rect 19 298 20 299
rect 18 298 19 299
rect 17 298 18 299
rect 16 298 17 299
rect 15 298 16 299
rect 14 298 15 299
rect 142 299 143 300
rect 141 299 142 300
rect 140 299 141 300
rect 139 299 140 300
rect 127 299 128 300
rect 126 299 127 300
rect 125 299 126 300
rect 124 299 125 300
rect 80 299 81 300
rect 79 299 80 300
rect 78 299 79 300
rect 77 299 78 300
rect 76 299 77 300
rect 75 299 76 300
rect 74 299 75 300
rect 73 299 74 300
rect 72 299 73 300
rect 71 299 72 300
rect 70 299 71 300
rect 69 299 70 300
rect 68 299 69 300
rect 67 299 68 300
rect 66 299 67 300
rect 52 299 53 300
rect 51 299 52 300
rect 50 299 51 300
rect 49 299 50 300
rect 48 299 49 300
rect 47 299 48 300
rect 46 299 47 300
rect 45 299 46 300
rect 44 299 45 300
rect 43 299 44 300
rect 42 299 43 300
rect 41 299 42 300
rect 40 299 41 300
rect 39 299 40 300
rect 38 299 39 300
rect 37 299 38 300
rect 36 299 37 300
rect 35 299 36 300
rect 34 299 35 300
rect 33 299 34 300
rect 32 299 33 300
rect 31 299 32 300
rect 30 299 31 300
rect 29 299 30 300
rect 28 299 29 300
rect 27 299 28 300
rect 26 299 27 300
rect 25 299 26 300
rect 24 299 25 300
rect 23 299 24 300
rect 22 299 23 300
rect 21 299 22 300
rect 20 299 21 300
rect 19 299 20 300
rect 18 299 19 300
rect 17 299 18 300
rect 16 299 17 300
rect 15 299 16 300
rect 14 299 15 300
rect 142 300 143 301
rect 141 300 142 301
rect 140 300 141 301
rect 139 300 140 301
rect 138 300 139 301
rect 128 300 129 301
rect 127 300 128 301
rect 126 300 127 301
rect 125 300 126 301
rect 124 300 125 301
rect 80 300 81 301
rect 79 300 80 301
rect 78 300 79 301
rect 77 300 78 301
rect 76 300 77 301
rect 75 300 76 301
rect 74 300 75 301
rect 73 300 74 301
rect 72 300 73 301
rect 71 300 72 301
rect 70 300 71 301
rect 69 300 70 301
rect 68 300 69 301
rect 67 300 68 301
rect 66 300 67 301
rect 52 300 53 301
rect 51 300 52 301
rect 50 300 51 301
rect 49 300 50 301
rect 48 300 49 301
rect 47 300 48 301
rect 46 300 47 301
rect 45 300 46 301
rect 44 300 45 301
rect 43 300 44 301
rect 42 300 43 301
rect 41 300 42 301
rect 40 300 41 301
rect 39 300 40 301
rect 38 300 39 301
rect 37 300 38 301
rect 36 300 37 301
rect 35 300 36 301
rect 34 300 35 301
rect 33 300 34 301
rect 32 300 33 301
rect 31 300 32 301
rect 30 300 31 301
rect 29 300 30 301
rect 28 300 29 301
rect 27 300 28 301
rect 26 300 27 301
rect 25 300 26 301
rect 24 300 25 301
rect 23 300 24 301
rect 22 300 23 301
rect 21 300 22 301
rect 20 300 21 301
rect 19 300 20 301
rect 18 300 19 301
rect 17 300 18 301
rect 16 300 17 301
rect 15 300 16 301
rect 14 300 15 301
rect 142 301 143 302
rect 141 301 142 302
rect 140 301 141 302
rect 139 301 140 302
rect 138 301 139 302
rect 137 301 138 302
rect 129 301 130 302
rect 128 301 129 302
rect 127 301 128 302
rect 126 301 127 302
rect 125 301 126 302
rect 124 301 125 302
rect 80 301 81 302
rect 79 301 80 302
rect 78 301 79 302
rect 77 301 78 302
rect 76 301 77 302
rect 75 301 76 302
rect 74 301 75 302
rect 73 301 74 302
rect 72 301 73 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 68 301 69 302
rect 67 301 68 302
rect 66 301 67 302
rect 52 301 53 302
rect 51 301 52 302
rect 50 301 51 302
rect 49 301 50 302
rect 48 301 49 302
rect 47 301 48 302
rect 46 301 47 302
rect 45 301 46 302
rect 44 301 45 302
rect 43 301 44 302
rect 42 301 43 302
rect 41 301 42 302
rect 40 301 41 302
rect 39 301 40 302
rect 38 301 39 302
rect 37 301 38 302
rect 36 301 37 302
rect 35 301 36 302
rect 34 301 35 302
rect 33 301 34 302
rect 32 301 33 302
rect 31 301 32 302
rect 30 301 31 302
rect 29 301 30 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 25 301 26 302
rect 24 301 25 302
rect 23 301 24 302
rect 22 301 23 302
rect 21 301 22 302
rect 20 301 21 302
rect 19 301 20 302
rect 18 301 19 302
rect 17 301 18 302
rect 16 301 17 302
rect 15 301 16 302
rect 14 301 15 302
rect 141 302 142 303
rect 140 302 141 303
rect 139 302 140 303
rect 138 302 139 303
rect 137 302 138 303
rect 136 302 137 303
rect 135 302 136 303
rect 131 302 132 303
rect 130 302 131 303
rect 129 302 130 303
rect 128 302 129 303
rect 127 302 128 303
rect 126 302 127 303
rect 125 302 126 303
rect 80 302 81 303
rect 79 302 80 303
rect 78 302 79 303
rect 77 302 78 303
rect 76 302 77 303
rect 75 302 76 303
rect 74 302 75 303
rect 73 302 74 303
rect 72 302 73 303
rect 71 302 72 303
rect 70 302 71 303
rect 69 302 70 303
rect 68 302 69 303
rect 67 302 68 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 48 302 49 303
rect 47 302 48 303
rect 46 302 47 303
rect 45 302 46 303
rect 44 302 45 303
rect 43 302 44 303
rect 42 302 43 303
rect 41 302 42 303
rect 40 302 41 303
rect 39 302 40 303
rect 38 302 39 303
rect 37 302 38 303
rect 36 302 37 303
rect 35 302 36 303
rect 34 302 35 303
rect 33 302 34 303
rect 32 302 33 303
rect 31 302 32 303
rect 30 302 31 303
rect 29 302 30 303
rect 28 302 29 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 24 302 25 303
rect 23 302 24 303
rect 22 302 23 303
rect 21 302 22 303
rect 20 302 21 303
rect 19 302 20 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 15 302 16 303
rect 14 302 15 303
rect 141 303 142 304
rect 140 303 141 304
rect 139 303 140 304
rect 138 303 139 304
rect 137 303 138 304
rect 136 303 137 304
rect 135 303 136 304
rect 134 303 135 304
rect 133 303 134 304
rect 132 303 133 304
rect 131 303 132 304
rect 130 303 131 304
rect 129 303 130 304
rect 128 303 129 304
rect 127 303 128 304
rect 126 303 127 304
rect 125 303 126 304
rect 80 303 81 304
rect 79 303 80 304
rect 78 303 79 304
rect 77 303 78 304
rect 76 303 77 304
rect 75 303 76 304
rect 74 303 75 304
rect 73 303 74 304
rect 72 303 73 304
rect 71 303 72 304
rect 70 303 71 304
rect 69 303 70 304
rect 68 303 69 304
rect 67 303 68 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 48 303 49 304
rect 47 303 48 304
rect 46 303 47 304
rect 45 303 46 304
rect 44 303 45 304
rect 43 303 44 304
rect 42 303 43 304
rect 41 303 42 304
rect 40 303 41 304
rect 39 303 40 304
rect 38 303 39 304
rect 37 303 38 304
rect 36 303 37 304
rect 35 303 36 304
rect 34 303 35 304
rect 33 303 34 304
rect 32 303 33 304
rect 31 303 32 304
rect 30 303 31 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 26 303 27 304
rect 25 303 26 304
rect 24 303 25 304
rect 23 303 24 304
rect 22 303 23 304
rect 21 303 22 304
rect 20 303 21 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 15 303 16 304
rect 14 303 15 304
rect 140 304 141 305
rect 139 304 140 305
rect 138 304 139 305
rect 137 304 138 305
rect 136 304 137 305
rect 135 304 136 305
rect 134 304 135 305
rect 133 304 134 305
rect 132 304 133 305
rect 131 304 132 305
rect 130 304 131 305
rect 129 304 130 305
rect 128 304 129 305
rect 127 304 128 305
rect 126 304 127 305
rect 80 304 81 305
rect 79 304 80 305
rect 78 304 79 305
rect 77 304 78 305
rect 76 304 77 305
rect 75 304 76 305
rect 74 304 75 305
rect 73 304 74 305
rect 72 304 73 305
rect 71 304 72 305
rect 70 304 71 305
rect 69 304 70 305
rect 68 304 69 305
rect 67 304 68 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 48 304 49 305
rect 47 304 48 305
rect 46 304 47 305
rect 45 304 46 305
rect 44 304 45 305
rect 43 304 44 305
rect 42 304 43 305
rect 41 304 42 305
rect 40 304 41 305
rect 39 304 40 305
rect 38 304 39 305
rect 37 304 38 305
rect 36 304 37 305
rect 35 304 36 305
rect 34 304 35 305
rect 33 304 34 305
rect 32 304 33 305
rect 31 304 32 305
rect 30 304 31 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 22 304 23 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 17 304 18 305
rect 16 304 17 305
rect 15 304 16 305
rect 14 304 15 305
rect 139 305 140 306
rect 138 305 139 306
rect 137 305 138 306
rect 136 305 137 306
rect 135 305 136 306
rect 134 305 135 306
rect 133 305 134 306
rect 132 305 133 306
rect 131 305 132 306
rect 130 305 131 306
rect 129 305 130 306
rect 128 305 129 306
rect 127 305 128 306
rect 126 305 127 306
rect 81 305 82 306
rect 80 305 81 306
rect 79 305 80 306
rect 78 305 79 306
rect 77 305 78 306
rect 76 305 77 306
rect 75 305 76 306
rect 74 305 75 306
rect 73 305 74 306
rect 72 305 73 306
rect 71 305 72 306
rect 70 305 71 306
rect 69 305 70 306
rect 68 305 69 306
rect 67 305 68 306
rect 52 305 53 306
rect 51 305 52 306
rect 50 305 51 306
rect 49 305 50 306
rect 48 305 49 306
rect 47 305 48 306
rect 46 305 47 306
rect 45 305 46 306
rect 44 305 45 306
rect 43 305 44 306
rect 42 305 43 306
rect 41 305 42 306
rect 40 305 41 306
rect 39 305 40 306
rect 38 305 39 306
rect 37 305 38 306
rect 36 305 37 306
rect 35 305 36 306
rect 34 305 35 306
rect 33 305 34 306
rect 32 305 33 306
rect 31 305 32 306
rect 30 305 31 306
rect 29 305 30 306
rect 28 305 29 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 17 305 18 306
rect 16 305 17 306
rect 15 305 16 306
rect 14 305 15 306
rect 138 306 139 307
rect 137 306 138 307
rect 136 306 137 307
rect 135 306 136 307
rect 134 306 135 307
rect 133 306 134 307
rect 132 306 133 307
rect 131 306 132 307
rect 130 306 131 307
rect 129 306 130 307
rect 128 306 129 307
rect 81 306 82 307
rect 80 306 81 307
rect 79 306 80 307
rect 78 306 79 307
rect 77 306 78 307
rect 76 306 77 307
rect 75 306 76 307
rect 74 306 75 307
rect 73 306 74 307
rect 72 306 73 307
rect 71 306 72 307
rect 70 306 71 307
rect 69 306 70 307
rect 68 306 69 307
rect 67 306 68 307
rect 52 306 53 307
rect 51 306 52 307
rect 50 306 51 307
rect 49 306 50 307
rect 48 306 49 307
rect 47 306 48 307
rect 46 306 47 307
rect 45 306 46 307
rect 44 306 45 307
rect 43 306 44 307
rect 42 306 43 307
rect 41 306 42 307
rect 40 306 41 307
rect 39 306 40 307
rect 38 306 39 307
rect 37 306 38 307
rect 36 306 37 307
rect 35 306 36 307
rect 34 306 35 307
rect 33 306 34 307
rect 32 306 33 307
rect 31 306 32 307
rect 30 306 31 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 17 306 18 307
rect 16 306 17 307
rect 15 306 16 307
rect 14 306 15 307
rect 136 307 137 308
rect 135 307 136 308
rect 134 307 135 308
rect 133 307 134 308
rect 132 307 133 308
rect 131 307 132 308
rect 130 307 131 308
rect 129 307 130 308
rect 81 307 82 308
rect 80 307 81 308
rect 79 307 80 308
rect 78 307 79 308
rect 77 307 78 308
rect 76 307 77 308
rect 75 307 76 308
rect 74 307 75 308
rect 73 307 74 308
rect 72 307 73 308
rect 71 307 72 308
rect 70 307 71 308
rect 69 307 70 308
rect 68 307 69 308
rect 67 307 68 308
rect 52 307 53 308
rect 51 307 52 308
rect 50 307 51 308
rect 49 307 50 308
rect 48 307 49 308
rect 47 307 48 308
rect 46 307 47 308
rect 45 307 46 308
rect 44 307 45 308
rect 43 307 44 308
rect 42 307 43 308
rect 41 307 42 308
rect 40 307 41 308
rect 39 307 40 308
rect 38 307 39 308
rect 37 307 38 308
rect 36 307 37 308
rect 35 307 36 308
rect 34 307 35 308
rect 33 307 34 308
rect 32 307 33 308
rect 31 307 32 308
rect 30 307 31 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 17 307 18 308
rect 16 307 17 308
rect 15 307 16 308
rect 14 307 15 308
rect 81 308 82 309
rect 80 308 81 309
rect 79 308 80 309
rect 78 308 79 309
rect 77 308 78 309
rect 76 308 77 309
rect 75 308 76 309
rect 74 308 75 309
rect 73 308 74 309
rect 72 308 73 309
rect 71 308 72 309
rect 70 308 71 309
rect 69 308 70 309
rect 68 308 69 309
rect 67 308 68 309
rect 52 308 53 309
rect 51 308 52 309
rect 50 308 51 309
rect 49 308 50 309
rect 48 308 49 309
rect 47 308 48 309
rect 46 308 47 309
rect 45 308 46 309
rect 44 308 45 309
rect 43 308 44 309
rect 42 308 43 309
rect 41 308 42 309
rect 40 308 41 309
rect 39 308 40 309
rect 38 308 39 309
rect 37 308 38 309
rect 36 308 37 309
rect 35 308 36 309
rect 34 308 35 309
rect 33 308 34 309
rect 32 308 33 309
rect 31 308 32 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 15 308 16 309
rect 14 308 15 309
rect 81 309 82 310
rect 80 309 81 310
rect 79 309 80 310
rect 78 309 79 310
rect 77 309 78 310
rect 76 309 77 310
rect 75 309 76 310
rect 74 309 75 310
rect 73 309 74 310
rect 72 309 73 310
rect 71 309 72 310
rect 70 309 71 310
rect 69 309 70 310
rect 68 309 69 310
rect 67 309 68 310
rect 52 309 53 310
rect 51 309 52 310
rect 50 309 51 310
rect 49 309 50 310
rect 48 309 49 310
rect 47 309 48 310
rect 46 309 47 310
rect 45 309 46 310
rect 44 309 45 310
rect 43 309 44 310
rect 42 309 43 310
rect 41 309 42 310
rect 40 309 41 310
rect 39 309 40 310
rect 38 309 39 310
rect 37 309 38 310
rect 36 309 37 310
rect 35 309 36 310
rect 34 309 35 310
rect 33 309 34 310
rect 32 309 33 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 17 309 18 310
rect 16 309 17 310
rect 15 309 16 310
rect 14 309 15 310
rect 81 310 82 311
rect 80 310 81 311
rect 79 310 80 311
rect 78 310 79 311
rect 77 310 78 311
rect 76 310 77 311
rect 75 310 76 311
rect 74 310 75 311
rect 73 310 74 311
rect 72 310 73 311
rect 71 310 72 311
rect 70 310 71 311
rect 69 310 70 311
rect 68 310 69 311
rect 67 310 68 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 48 310 49 311
rect 47 310 48 311
rect 46 310 47 311
rect 45 310 46 311
rect 44 310 45 311
rect 43 310 44 311
rect 42 310 43 311
rect 41 310 42 311
rect 40 310 41 311
rect 39 310 40 311
rect 38 310 39 311
rect 37 310 38 311
rect 36 310 37 311
rect 35 310 36 311
rect 34 310 35 311
rect 33 310 34 311
rect 32 310 33 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 16 310 17 311
rect 15 310 16 311
rect 14 310 15 311
rect 136 311 137 312
rect 135 311 136 312
rect 134 311 135 312
rect 133 311 134 312
rect 132 311 133 312
rect 131 311 132 312
rect 130 311 131 312
rect 81 311 82 312
rect 80 311 81 312
rect 79 311 80 312
rect 78 311 79 312
rect 77 311 78 312
rect 76 311 77 312
rect 75 311 76 312
rect 74 311 75 312
rect 73 311 74 312
rect 72 311 73 312
rect 71 311 72 312
rect 70 311 71 312
rect 69 311 70 312
rect 68 311 69 312
rect 67 311 68 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 48 311 49 312
rect 47 311 48 312
rect 46 311 47 312
rect 45 311 46 312
rect 44 311 45 312
rect 43 311 44 312
rect 42 311 43 312
rect 41 311 42 312
rect 40 311 41 312
rect 39 311 40 312
rect 38 311 39 312
rect 37 311 38 312
rect 36 311 37 312
rect 35 311 36 312
rect 34 311 35 312
rect 33 311 34 312
rect 32 311 33 312
rect 31 311 32 312
rect 30 311 31 312
rect 29 311 30 312
rect 28 311 29 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 15 311 16 312
rect 14 311 15 312
rect 138 312 139 313
rect 137 312 138 313
rect 136 312 137 313
rect 135 312 136 313
rect 134 312 135 313
rect 133 312 134 313
rect 132 312 133 313
rect 131 312 132 313
rect 130 312 131 313
rect 129 312 130 313
rect 128 312 129 313
rect 81 312 82 313
rect 80 312 81 313
rect 79 312 80 313
rect 78 312 79 313
rect 77 312 78 313
rect 76 312 77 313
rect 75 312 76 313
rect 74 312 75 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 68 312 69 313
rect 67 312 68 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 48 312 49 313
rect 47 312 48 313
rect 46 312 47 313
rect 45 312 46 313
rect 44 312 45 313
rect 43 312 44 313
rect 42 312 43 313
rect 41 312 42 313
rect 40 312 41 313
rect 39 312 40 313
rect 38 312 39 313
rect 37 312 38 313
rect 36 312 37 313
rect 35 312 36 313
rect 34 312 35 313
rect 33 312 34 313
rect 32 312 33 313
rect 31 312 32 313
rect 30 312 31 313
rect 29 312 30 313
rect 28 312 29 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 15 312 16 313
rect 14 312 15 313
rect 139 313 140 314
rect 138 313 139 314
rect 137 313 138 314
rect 136 313 137 314
rect 135 313 136 314
rect 134 313 135 314
rect 133 313 134 314
rect 132 313 133 314
rect 131 313 132 314
rect 130 313 131 314
rect 129 313 130 314
rect 128 313 129 314
rect 127 313 128 314
rect 81 313 82 314
rect 80 313 81 314
rect 79 313 80 314
rect 78 313 79 314
rect 77 313 78 314
rect 76 313 77 314
rect 75 313 76 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 68 313 69 314
rect 67 313 68 314
rect 66 313 67 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 48 313 49 314
rect 47 313 48 314
rect 46 313 47 314
rect 45 313 46 314
rect 44 313 45 314
rect 43 313 44 314
rect 42 313 43 314
rect 41 313 42 314
rect 40 313 41 314
rect 39 313 40 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 17 313 18 314
rect 16 313 17 314
rect 15 313 16 314
rect 14 313 15 314
rect 140 314 141 315
rect 139 314 140 315
rect 138 314 139 315
rect 137 314 138 315
rect 136 314 137 315
rect 135 314 136 315
rect 134 314 135 315
rect 133 314 134 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 129 314 130 315
rect 128 314 129 315
rect 127 314 128 315
rect 126 314 127 315
rect 81 314 82 315
rect 80 314 81 315
rect 79 314 80 315
rect 78 314 79 315
rect 77 314 78 315
rect 76 314 77 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 68 314 69 315
rect 67 314 68 315
rect 66 314 67 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 48 314 49 315
rect 47 314 48 315
rect 46 314 47 315
rect 45 314 46 315
rect 44 314 45 315
rect 43 314 44 315
rect 42 314 43 315
rect 41 314 42 315
rect 40 314 41 315
rect 39 314 40 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 17 314 18 315
rect 16 314 17 315
rect 15 314 16 315
rect 14 314 15 315
rect 141 315 142 316
rect 140 315 141 316
rect 139 315 140 316
rect 138 315 139 316
rect 137 315 138 316
rect 136 315 137 316
rect 135 315 136 316
rect 134 315 135 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 128 315 129 316
rect 127 315 128 316
rect 126 315 127 316
rect 125 315 126 316
rect 81 315 82 316
rect 80 315 81 316
rect 79 315 80 316
rect 78 315 79 316
rect 77 315 78 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 67 315 68 316
rect 66 315 67 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 48 315 49 316
rect 47 315 48 316
rect 46 315 47 316
rect 45 315 46 316
rect 44 315 45 316
rect 43 315 44 316
rect 42 315 43 316
rect 41 315 42 316
rect 40 315 41 316
rect 39 315 40 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 17 315 18 316
rect 16 315 17 316
rect 15 315 16 316
rect 14 315 15 316
rect 141 316 142 317
rect 140 316 141 317
rect 139 316 140 317
rect 138 316 139 317
rect 137 316 138 317
rect 136 316 137 317
rect 135 316 136 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 131 316 132 317
rect 130 316 131 317
rect 129 316 130 317
rect 128 316 129 317
rect 127 316 128 317
rect 126 316 127 317
rect 125 316 126 317
rect 81 316 82 317
rect 80 316 81 317
rect 79 316 80 317
rect 78 316 79 317
rect 77 316 78 317
rect 76 316 77 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 67 316 68 317
rect 66 316 67 317
rect 65 316 66 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 48 316 49 317
rect 47 316 48 317
rect 46 316 47 317
rect 45 316 46 317
rect 44 316 45 317
rect 43 316 44 317
rect 42 316 43 317
rect 41 316 42 317
rect 40 316 41 317
rect 39 316 40 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 18 316 19 317
rect 17 316 18 317
rect 16 316 17 317
rect 15 316 16 317
rect 14 316 15 317
rect 142 317 143 318
rect 141 317 142 318
rect 140 317 141 318
rect 139 317 140 318
rect 138 317 139 318
rect 137 317 138 318
rect 129 317 130 318
rect 128 317 129 318
rect 127 317 128 318
rect 126 317 127 318
rect 125 317 126 318
rect 124 317 125 318
rect 81 317 82 318
rect 80 317 81 318
rect 79 317 80 318
rect 78 317 79 318
rect 77 317 78 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 67 317 68 318
rect 66 317 67 318
rect 65 317 66 318
rect 64 317 65 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 48 317 49 318
rect 47 317 48 318
rect 46 317 47 318
rect 45 317 46 318
rect 44 317 45 318
rect 43 317 44 318
rect 42 317 43 318
rect 41 317 42 318
rect 40 317 41 318
rect 39 317 40 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 19 317 20 318
rect 18 317 19 318
rect 17 317 18 318
rect 16 317 17 318
rect 15 317 16 318
rect 14 317 15 318
rect 142 318 143 319
rect 141 318 142 319
rect 140 318 141 319
rect 139 318 140 319
rect 138 318 139 319
rect 128 318 129 319
rect 127 318 128 319
rect 126 318 127 319
rect 125 318 126 319
rect 124 318 125 319
rect 80 318 81 319
rect 79 318 80 319
rect 78 318 79 319
rect 77 318 78 319
rect 76 318 77 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 69 318 70 319
rect 68 318 69 319
rect 67 318 68 319
rect 66 318 67 319
rect 65 318 66 319
rect 64 318 65 319
rect 63 318 64 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 48 318 49 319
rect 47 318 48 319
rect 46 318 47 319
rect 45 318 46 319
rect 44 318 45 319
rect 43 318 44 319
rect 42 318 43 319
rect 41 318 42 319
rect 40 318 41 319
rect 39 318 40 319
rect 29 318 30 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 17 318 18 319
rect 16 318 17 319
rect 15 318 16 319
rect 14 318 15 319
rect 142 319 143 320
rect 141 319 142 320
rect 140 319 141 320
rect 139 319 140 320
rect 138 319 139 320
rect 128 319 129 320
rect 127 319 128 320
rect 126 319 127 320
rect 125 319 126 320
rect 124 319 125 320
rect 80 319 81 320
rect 79 319 80 320
rect 78 319 79 320
rect 77 319 78 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 69 319 70 320
rect 68 319 69 320
rect 67 319 68 320
rect 66 319 67 320
rect 65 319 66 320
rect 64 319 65 320
rect 63 319 64 320
rect 62 319 63 320
rect 61 319 62 320
rect 60 319 61 320
rect 59 319 60 320
rect 58 319 59 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 48 319 49 320
rect 47 319 48 320
rect 46 319 47 320
rect 45 319 46 320
rect 44 319 45 320
rect 43 319 44 320
rect 42 319 43 320
rect 41 319 42 320
rect 40 319 41 320
rect 39 319 40 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 17 319 18 320
rect 16 319 17 320
rect 15 319 16 320
rect 14 319 15 320
rect 142 320 143 321
rect 141 320 142 321
rect 140 320 141 321
rect 139 320 140 321
rect 127 320 128 321
rect 126 320 127 321
rect 125 320 126 321
rect 124 320 125 321
rect 80 320 81 321
rect 79 320 80 321
rect 78 320 79 321
rect 77 320 78 321
rect 76 320 77 321
rect 75 320 76 321
rect 74 320 75 321
rect 73 320 74 321
rect 72 320 73 321
rect 71 320 72 321
rect 70 320 71 321
rect 69 320 70 321
rect 68 320 69 321
rect 67 320 68 321
rect 66 320 67 321
rect 65 320 66 321
rect 64 320 65 321
rect 63 320 64 321
rect 62 320 63 321
rect 61 320 62 321
rect 60 320 61 321
rect 59 320 60 321
rect 58 320 59 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 48 320 49 321
rect 47 320 48 321
rect 46 320 47 321
rect 45 320 46 321
rect 44 320 45 321
rect 43 320 44 321
rect 42 320 43 321
rect 41 320 42 321
rect 40 320 41 321
rect 39 320 40 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 17 320 18 321
rect 16 320 17 321
rect 15 320 16 321
rect 14 320 15 321
rect 142 321 143 322
rect 141 321 142 322
rect 140 321 141 322
rect 139 321 140 322
rect 127 321 128 322
rect 126 321 127 322
rect 125 321 126 322
rect 124 321 125 322
rect 80 321 81 322
rect 79 321 80 322
rect 78 321 79 322
rect 77 321 78 322
rect 76 321 77 322
rect 75 321 76 322
rect 74 321 75 322
rect 73 321 74 322
rect 72 321 73 322
rect 71 321 72 322
rect 70 321 71 322
rect 69 321 70 322
rect 68 321 69 322
rect 67 321 68 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 61 321 62 322
rect 60 321 61 322
rect 59 321 60 322
rect 58 321 59 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 48 321 49 322
rect 47 321 48 322
rect 46 321 47 322
rect 45 321 46 322
rect 44 321 45 322
rect 43 321 44 322
rect 42 321 43 322
rect 41 321 42 322
rect 40 321 41 322
rect 39 321 40 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 18 321 19 322
rect 17 321 18 322
rect 16 321 17 322
rect 15 321 16 322
rect 14 321 15 322
rect 142 322 143 323
rect 141 322 142 323
rect 140 322 141 323
rect 139 322 140 323
rect 138 322 139 323
rect 128 322 129 323
rect 127 322 128 323
rect 126 322 127 323
rect 125 322 126 323
rect 124 322 125 323
rect 79 322 80 323
rect 78 322 79 323
rect 77 322 78 323
rect 76 322 77 323
rect 75 322 76 323
rect 74 322 75 323
rect 73 322 74 323
rect 72 322 73 323
rect 71 322 72 323
rect 70 322 71 323
rect 69 322 70 323
rect 68 322 69 323
rect 67 322 68 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 61 322 62 323
rect 60 322 61 323
rect 59 322 60 323
rect 58 322 59 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 48 322 49 323
rect 47 322 48 323
rect 46 322 47 323
rect 45 322 46 323
rect 44 322 45 323
rect 43 322 44 323
rect 42 322 43 323
rect 41 322 42 323
rect 40 322 41 323
rect 39 322 40 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 18 322 19 323
rect 17 322 18 323
rect 16 322 17 323
rect 15 322 16 323
rect 14 322 15 323
rect 142 323 143 324
rect 141 323 142 324
rect 140 323 141 324
rect 139 323 140 324
rect 138 323 139 324
rect 128 323 129 324
rect 127 323 128 324
rect 126 323 127 324
rect 125 323 126 324
rect 124 323 125 324
rect 79 323 80 324
rect 78 323 79 324
rect 77 323 78 324
rect 76 323 77 324
rect 75 323 76 324
rect 74 323 75 324
rect 73 323 74 324
rect 72 323 73 324
rect 71 323 72 324
rect 70 323 71 324
rect 69 323 70 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 59 323 60 324
rect 58 323 59 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 48 323 49 324
rect 47 323 48 324
rect 46 323 47 324
rect 45 323 46 324
rect 44 323 45 324
rect 43 323 44 324
rect 42 323 43 324
rect 41 323 42 324
rect 40 323 41 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 20 323 21 324
rect 19 323 20 324
rect 18 323 19 324
rect 17 323 18 324
rect 16 323 17 324
rect 15 323 16 324
rect 14 323 15 324
rect 142 324 143 325
rect 141 324 142 325
rect 140 324 141 325
rect 139 324 140 325
rect 138 324 139 325
rect 137 324 138 325
rect 129 324 130 325
rect 128 324 129 325
rect 127 324 128 325
rect 126 324 127 325
rect 125 324 126 325
rect 124 324 125 325
rect 79 324 80 325
rect 78 324 79 325
rect 77 324 78 325
rect 76 324 77 325
rect 75 324 76 325
rect 74 324 75 325
rect 73 324 74 325
rect 72 324 73 325
rect 71 324 72 325
rect 70 324 71 325
rect 69 324 70 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 59 324 60 325
rect 58 324 59 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 49 324 50 325
rect 48 324 49 325
rect 47 324 48 325
rect 46 324 47 325
rect 45 324 46 325
rect 44 324 45 325
rect 43 324 44 325
rect 42 324 43 325
rect 41 324 42 325
rect 40 324 41 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 19 324 20 325
rect 18 324 19 325
rect 17 324 18 325
rect 16 324 17 325
rect 15 324 16 325
rect 14 324 15 325
rect 141 325 142 326
rect 140 325 141 326
rect 139 325 140 326
rect 138 325 139 326
rect 137 325 138 326
rect 136 325 137 326
rect 135 325 136 326
rect 134 325 135 326
rect 133 325 134 326
rect 132 325 133 326
rect 131 325 132 326
rect 130 325 131 326
rect 129 325 130 326
rect 128 325 129 326
rect 127 325 128 326
rect 126 325 127 326
rect 125 325 126 326
rect 78 325 79 326
rect 77 325 78 326
rect 76 325 77 326
rect 75 325 76 326
rect 74 325 75 326
rect 73 325 74 326
rect 72 325 73 326
rect 71 325 72 326
rect 70 325 71 326
rect 69 325 70 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 59 325 60 326
rect 58 325 59 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 49 325 50 326
rect 48 325 49 326
rect 47 325 48 326
rect 46 325 47 326
rect 45 325 46 326
rect 44 325 45 326
rect 43 325 44 326
rect 42 325 43 326
rect 41 325 42 326
rect 40 325 41 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 20 325 21 326
rect 19 325 20 326
rect 18 325 19 326
rect 17 325 18 326
rect 16 325 17 326
rect 15 325 16 326
rect 14 325 15 326
rect 141 326 142 327
rect 140 326 141 327
rect 139 326 140 327
rect 138 326 139 327
rect 137 326 138 327
rect 136 326 137 327
rect 135 326 136 327
rect 134 326 135 327
rect 133 326 134 327
rect 132 326 133 327
rect 131 326 132 327
rect 130 326 131 327
rect 129 326 130 327
rect 128 326 129 327
rect 127 326 128 327
rect 126 326 127 327
rect 125 326 126 327
rect 78 326 79 327
rect 77 326 78 327
rect 76 326 77 327
rect 75 326 76 327
rect 74 326 75 327
rect 73 326 74 327
rect 72 326 73 327
rect 71 326 72 327
rect 70 326 71 327
rect 69 326 70 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 59 326 60 327
rect 58 326 59 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 49 326 50 327
rect 48 326 49 327
rect 47 326 48 327
rect 46 326 47 327
rect 45 326 46 327
rect 44 326 45 327
rect 43 326 44 327
rect 42 326 43 327
rect 41 326 42 327
rect 40 326 41 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 21 326 22 327
rect 20 326 21 327
rect 19 326 20 327
rect 18 326 19 327
rect 17 326 18 327
rect 16 326 17 327
rect 15 326 16 327
rect 14 326 15 327
rect 140 327 141 328
rect 139 327 140 328
rect 138 327 139 328
rect 137 327 138 328
rect 136 327 137 328
rect 135 327 136 328
rect 134 327 135 328
rect 133 327 134 328
rect 132 327 133 328
rect 131 327 132 328
rect 130 327 131 328
rect 129 327 130 328
rect 128 327 129 328
rect 127 327 128 328
rect 126 327 127 328
rect 77 327 78 328
rect 76 327 77 328
rect 75 327 76 328
rect 74 327 75 328
rect 73 327 74 328
rect 72 327 73 328
rect 71 327 72 328
rect 70 327 71 328
rect 69 327 70 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 61 327 62 328
rect 60 327 61 328
rect 59 327 60 328
rect 58 327 59 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 50 327 51 328
rect 49 327 50 328
rect 48 327 49 328
rect 47 327 48 328
rect 46 327 47 328
rect 45 327 46 328
rect 44 327 45 328
rect 43 327 44 328
rect 42 327 43 328
rect 41 327 42 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 22 327 23 328
rect 21 327 22 328
rect 20 327 21 328
rect 19 327 20 328
rect 18 327 19 328
rect 17 327 18 328
rect 16 327 17 328
rect 15 327 16 328
rect 14 327 15 328
rect 139 328 140 329
rect 138 328 139 329
rect 137 328 138 329
rect 136 328 137 329
rect 135 328 136 329
rect 134 328 135 329
rect 133 328 134 329
rect 132 328 133 329
rect 131 328 132 329
rect 130 328 131 329
rect 129 328 130 329
rect 128 328 129 329
rect 127 328 128 329
rect 77 328 78 329
rect 76 328 77 329
rect 75 328 76 329
rect 74 328 75 329
rect 73 328 74 329
rect 72 328 73 329
rect 71 328 72 329
rect 70 328 71 329
rect 69 328 70 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 61 328 62 329
rect 60 328 61 329
rect 59 328 60 329
rect 58 328 59 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 50 328 51 329
rect 49 328 50 329
rect 48 328 49 329
rect 47 328 48 329
rect 46 328 47 329
rect 45 328 46 329
rect 44 328 45 329
rect 43 328 44 329
rect 42 328 43 329
rect 41 328 42 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 22 328 23 329
rect 21 328 22 329
rect 20 328 21 329
rect 19 328 20 329
rect 18 328 19 329
rect 17 328 18 329
rect 16 328 17 329
rect 15 328 16 329
rect 14 328 15 329
rect 138 329 139 330
rect 137 329 138 330
rect 136 329 137 330
rect 135 329 136 330
rect 134 329 135 330
rect 133 329 134 330
rect 132 329 133 330
rect 131 329 132 330
rect 130 329 131 330
rect 129 329 130 330
rect 128 329 129 330
rect 76 329 77 330
rect 75 329 76 330
rect 74 329 75 330
rect 73 329 74 330
rect 72 329 73 330
rect 71 329 72 330
rect 70 329 71 330
rect 69 329 70 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 63 329 64 330
rect 62 329 63 330
rect 61 329 62 330
rect 60 329 61 330
rect 59 329 60 330
rect 58 329 59 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 51 329 52 330
rect 50 329 51 330
rect 49 329 50 330
rect 48 329 49 330
rect 47 329 48 330
rect 46 329 47 330
rect 45 329 46 330
rect 44 329 45 330
rect 43 329 44 330
rect 42 329 43 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 23 329 24 330
rect 22 329 23 330
rect 21 329 22 330
rect 20 329 21 330
rect 19 329 20 330
rect 18 329 19 330
rect 17 329 18 330
rect 16 329 17 330
rect 15 329 16 330
rect 14 329 15 330
rect 135 330 136 331
rect 134 330 135 331
rect 133 330 134 331
rect 132 330 133 331
rect 131 330 132 331
rect 130 330 131 331
rect 75 330 76 331
rect 74 330 75 331
rect 73 330 74 331
rect 72 330 73 331
rect 71 330 72 331
rect 70 330 71 331
rect 69 330 70 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 63 330 64 331
rect 62 330 63 331
rect 61 330 62 331
rect 60 330 61 331
rect 59 330 60 331
rect 58 330 59 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 51 330 52 331
rect 50 330 51 331
rect 49 330 50 331
rect 48 330 49 331
rect 47 330 48 331
rect 46 330 47 331
rect 45 330 46 331
rect 44 330 45 331
rect 43 330 44 331
rect 42 330 43 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 24 330 25 331
rect 23 330 24 331
rect 22 330 23 331
rect 21 330 22 331
rect 20 330 21 331
rect 19 330 20 331
rect 18 330 19 331
rect 17 330 18 331
rect 16 330 17 331
rect 15 330 16 331
rect 14 330 15 331
rect 75 331 76 332
rect 74 331 75 332
rect 73 331 74 332
rect 72 331 73 332
rect 71 331 72 332
rect 70 331 71 332
rect 69 331 70 332
rect 68 331 69 332
rect 67 331 68 332
rect 66 331 67 332
rect 65 331 66 332
rect 64 331 65 332
rect 63 331 64 332
rect 62 331 63 332
rect 61 331 62 332
rect 60 331 61 332
rect 59 331 60 332
rect 58 331 59 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 52 331 53 332
rect 51 331 52 332
rect 50 331 51 332
rect 49 331 50 332
rect 48 331 49 332
rect 47 331 48 332
rect 46 331 47 332
rect 45 331 46 332
rect 44 331 45 332
rect 43 331 44 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 26 331 27 332
rect 25 331 26 332
rect 24 331 25 332
rect 23 331 24 332
rect 22 331 23 332
rect 21 331 22 332
rect 20 331 21 332
rect 19 331 20 332
rect 18 331 19 332
rect 17 331 18 332
rect 16 331 17 332
rect 15 331 16 332
rect 14 331 15 332
rect 74 332 75 333
rect 73 332 74 333
rect 72 332 73 333
rect 71 332 72 333
rect 70 332 71 333
rect 69 332 70 333
rect 68 332 69 333
rect 67 332 68 333
rect 66 332 67 333
rect 65 332 66 333
rect 64 332 65 333
rect 63 332 64 333
rect 62 332 63 333
rect 61 332 62 333
rect 60 332 61 333
rect 59 332 60 333
rect 58 332 59 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 52 332 53 333
rect 51 332 52 333
rect 50 332 51 333
rect 49 332 50 333
rect 48 332 49 333
rect 47 332 48 333
rect 46 332 47 333
rect 45 332 46 333
rect 44 332 45 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 26 332 27 333
rect 25 332 26 333
rect 24 332 25 333
rect 23 332 24 333
rect 22 332 23 333
rect 21 332 22 333
rect 20 332 21 333
rect 19 332 20 333
rect 18 332 19 333
rect 17 332 18 333
rect 16 332 17 333
rect 15 332 16 333
rect 14 332 15 333
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 52 333 53 334
rect 51 333 52 334
rect 50 333 51 334
rect 49 333 50 334
rect 48 333 49 334
rect 47 333 48 334
rect 46 333 47 334
rect 45 333 46 334
rect 44 333 45 334
rect 29 333 30 334
rect 28 333 29 334
rect 27 333 28 334
rect 26 333 27 334
rect 25 333 26 334
rect 24 333 25 334
rect 23 333 24 334
rect 22 333 23 334
rect 21 333 22 334
rect 20 333 21 334
rect 19 333 20 334
rect 18 333 19 334
rect 17 333 18 334
rect 16 333 17 334
rect 15 333 16 334
rect 14 333 15 334
rect 136 334 137 335
rect 135 334 136 335
rect 134 334 135 335
rect 133 334 134 335
rect 132 334 133 335
rect 131 334 132 335
rect 130 334 131 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 52 334 53 335
rect 51 334 52 335
rect 50 334 51 335
rect 49 334 50 335
rect 48 334 49 335
rect 47 334 48 335
rect 46 334 47 335
rect 29 334 30 335
rect 28 334 29 335
rect 27 334 28 335
rect 26 334 27 335
rect 25 334 26 335
rect 24 334 25 335
rect 23 334 24 335
rect 22 334 23 335
rect 21 334 22 335
rect 20 334 21 335
rect 19 334 20 335
rect 18 334 19 335
rect 17 334 18 335
rect 16 334 17 335
rect 15 334 16 335
rect 14 334 15 335
rect 139 335 140 336
rect 138 335 139 336
rect 137 335 138 336
rect 136 335 137 336
rect 135 335 136 336
rect 134 335 135 336
rect 133 335 134 336
rect 132 335 133 336
rect 131 335 132 336
rect 130 335 131 336
rect 129 335 130 336
rect 128 335 129 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 52 335 53 336
rect 51 335 52 336
rect 50 335 51 336
rect 49 335 50 336
rect 48 335 49 336
rect 47 335 48 336
rect 29 335 30 336
rect 28 335 29 336
rect 27 335 28 336
rect 26 335 27 336
rect 25 335 26 336
rect 24 335 25 336
rect 23 335 24 336
rect 22 335 23 336
rect 21 335 22 336
rect 20 335 21 336
rect 19 335 20 336
rect 18 335 19 336
rect 17 335 18 336
rect 16 335 17 336
rect 15 335 16 336
rect 14 335 15 336
rect 140 336 141 337
rect 139 336 140 337
rect 138 336 139 337
rect 137 336 138 337
rect 136 336 137 337
rect 135 336 136 337
rect 134 336 135 337
rect 133 336 134 337
rect 132 336 133 337
rect 131 336 132 337
rect 130 336 131 337
rect 129 336 130 337
rect 128 336 129 337
rect 127 336 128 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 52 336 53 337
rect 51 336 52 337
rect 50 336 51 337
rect 49 336 50 337
rect 48 336 49 337
rect 141 337 142 338
rect 140 337 141 338
rect 139 337 140 338
rect 138 337 139 338
rect 137 337 138 338
rect 136 337 137 338
rect 135 337 136 338
rect 134 337 135 338
rect 133 337 134 338
rect 132 337 133 338
rect 131 337 132 338
rect 130 337 131 338
rect 129 337 130 338
rect 128 337 129 338
rect 127 337 128 338
rect 126 337 127 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 52 337 53 338
rect 51 337 52 338
rect 141 338 142 339
rect 140 338 141 339
rect 139 338 140 339
rect 138 338 139 339
rect 137 338 138 339
rect 136 338 137 339
rect 135 338 136 339
rect 134 338 135 339
rect 133 338 134 339
rect 132 338 133 339
rect 131 338 132 339
rect 130 338 131 339
rect 129 338 130 339
rect 128 338 129 339
rect 127 338 128 339
rect 126 338 127 339
rect 125 338 126 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 142 339 143 340
rect 141 339 142 340
rect 140 339 141 340
rect 139 339 140 340
rect 138 339 139 340
rect 137 339 138 340
rect 136 339 137 340
rect 135 339 136 340
rect 134 339 135 340
rect 133 339 134 340
rect 132 339 133 340
rect 131 339 132 340
rect 130 339 131 340
rect 129 339 130 340
rect 128 339 129 340
rect 127 339 128 340
rect 126 339 127 340
rect 125 339 126 340
rect 142 340 143 341
rect 141 340 142 341
rect 140 340 141 341
rect 139 340 140 341
rect 138 340 139 341
rect 137 340 138 341
rect 129 340 130 341
rect 128 340 129 341
rect 127 340 128 341
rect 126 340 127 341
rect 125 340 126 341
rect 124 340 125 341
rect 142 341 143 342
rect 141 341 142 342
rect 140 341 141 342
rect 139 341 140 342
rect 138 341 139 342
rect 128 341 129 342
rect 127 341 128 342
rect 126 341 127 342
rect 125 341 126 342
rect 124 341 125 342
rect 142 342 143 343
rect 141 342 142 343
rect 140 342 141 343
rect 139 342 140 343
rect 138 342 139 343
rect 128 342 129 343
rect 127 342 128 343
rect 126 342 127 343
rect 125 342 126 343
rect 124 342 125 343
rect 142 343 143 344
rect 141 343 142 344
rect 140 343 141 344
rect 139 343 140 344
rect 127 343 128 344
rect 126 343 127 344
rect 125 343 126 344
rect 124 343 125 344
rect 141 344 142 345
rect 140 344 141 345
rect 139 344 140 345
rect 127 344 128 345
rect 126 344 127 345
rect 125 344 126 345
rect 124 344 125 345
rect 141 345 142 346
rect 140 345 141 346
rect 139 345 140 346
rect 138 345 139 346
rect 128 345 129 346
rect 127 345 128 346
rect 126 345 127 346
rect 125 345 126 346
rect 140 346 141 347
rect 139 346 140 347
rect 138 346 139 347
rect 137 346 138 347
rect 128 346 129 347
rect 127 346 128 347
rect 126 346 127 347
rect 125 346 126 347
rect 140 347 141 348
rect 139 347 140 348
rect 138 347 139 348
rect 137 347 138 348
rect 136 347 137 348
rect 135 347 136 348
rect 130 347 131 348
rect 129 347 130 348
rect 128 347 129 348
rect 127 347 128 348
rect 126 347 127 348
rect 142 348 143 349
rect 141 348 142 349
rect 140 348 141 349
rect 139 348 140 349
rect 138 348 139 349
rect 137 348 138 349
rect 136 348 137 349
rect 135 348 136 349
rect 134 348 135 349
rect 133 348 134 349
rect 132 348 133 349
rect 131 348 132 349
rect 130 348 131 349
rect 129 348 130 349
rect 128 348 129 349
rect 127 348 128 349
rect 126 348 127 349
rect 125 348 126 349
rect 124 348 125 349
rect 123 348 124 349
rect 122 348 123 349
rect 121 348 122 349
rect 120 348 121 349
rect 119 348 120 349
rect 118 348 119 349
rect 117 348 118 349
rect 116 348 117 349
rect 115 348 116 349
rect 53 348 54 349
rect 52 348 53 349
rect 51 348 52 349
rect 50 348 51 349
rect 49 348 50 349
rect 48 348 49 349
rect 47 348 48 349
rect 46 348 47 349
rect 45 348 46 349
rect 44 348 45 349
rect 43 348 44 349
rect 42 348 43 349
rect 142 349 143 350
rect 141 349 142 350
rect 140 349 141 350
rect 139 349 140 350
rect 138 349 139 350
rect 137 349 138 350
rect 136 349 137 350
rect 135 349 136 350
rect 134 349 135 350
rect 133 349 134 350
rect 132 349 133 350
rect 131 349 132 350
rect 130 349 131 350
rect 129 349 130 350
rect 128 349 129 350
rect 127 349 128 350
rect 126 349 127 350
rect 125 349 126 350
rect 124 349 125 350
rect 123 349 124 350
rect 122 349 123 350
rect 121 349 122 350
rect 120 349 121 350
rect 119 349 120 350
rect 118 349 119 350
rect 117 349 118 350
rect 116 349 117 350
rect 115 349 116 350
rect 61 349 62 350
rect 60 349 61 350
rect 59 349 60 350
rect 58 349 59 350
rect 57 349 58 350
rect 56 349 57 350
rect 55 349 56 350
rect 54 349 55 350
rect 53 349 54 350
rect 52 349 53 350
rect 51 349 52 350
rect 50 349 51 350
rect 49 349 50 350
rect 48 349 49 350
rect 47 349 48 350
rect 46 349 47 350
rect 45 349 46 350
rect 44 349 45 350
rect 43 349 44 350
rect 42 349 43 350
rect 41 349 42 350
rect 40 349 41 350
rect 39 349 40 350
rect 38 349 39 350
rect 37 349 38 350
rect 36 349 37 350
rect 35 349 36 350
rect 142 350 143 351
rect 141 350 142 351
rect 140 350 141 351
rect 139 350 140 351
rect 138 350 139 351
rect 137 350 138 351
rect 136 350 137 351
rect 135 350 136 351
rect 134 350 135 351
rect 133 350 134 351
rect 132 350 133 351
rect 131 350 132 351
rect 130 350 131 351
rect 129 350 130 351
rect 128 350 129 351
rect 127 350 128 351
rect 126 350 127 351
rect 125 350 126 351
rect 124 350 125 351
rect 123 350 124 351
rect 122 350 123 351
rect 121 350 122 351
rect 120 350 121 351
rect 119 350 120 351
rect 118 350 119 351
rect 117 350 118 351
rect 116 350 117 351
rect 115 350 116 351
rect 65 350 66 351
rect 64 350 65 351
rect 63 350 64 351
rect 62 350 63 351
rect 61 350 62 351
rect 60 350 61 351
rect 59 350 60 351
rect 58 350 59 351
rect 57 350 58 351
rect 56 350 57 351
rect 55 350 56 351
rect 54 350 55 351
rect 53 350 54 351
rect 52 350 53 351
rect 51 350 52 351
rect 50 350 51 351
rect 49 350 50 351
rect 48 350 49 351
rect 47 350 48 351
rect 46 350 47 351
rect 45 350 46 351
rect 44 350 45 351
rect 43 350 44 351
rect 42 350 43 351
rect 41 350 42 351
rect 40 350 41 351
rect 39 350 40 351
rect 38 350 39 351
rect 37 350 38 351
rect 36 350 37 351
rect 35 350 36 351
rect 34 350 35 351
rect 33 350 34 351
rect 32 350 33 351
rect 31 350 32 351
rect 142 351 143 352
rect 141 351 142 352
rect 140 351 141 352
rect 139 351 140 352
rect 138 351 139 352
rect 137 351 138 352
rect 136 351 137 352
rect 135 351 136 352
rect 134 351 135 352
rect 133 351 134 352
rect 132 351 133 352
rect 131 351 132 352
rect 130 351 131 352
rect 129 351 130 352
rect 128 351 129 352
rect 127 351 128 352
rect 126 351 127 352
rect 125 351 126 352
rect 124 351 125 352
rect 123 351 124 352
rect 122 351 123 352
rect 121 351 122 352
rect 120 351 121 352
rect 119 351 120 352
rect 118 351 119 352
rect 117 351 118 352
rect 116 351 117 352
rect 115 351 116 352
rect 67 351 68 352
rect 66 351 67 352
rect 65 351 66 352
rect 64 351 65 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 59 351 60 352
rect 58 351 59 352
rect 57 351 58 352
rect 56 351 57 352
rect 55 351 56 352
rect 54 351 55 352
rect 53 351 54 352
rect 52 351 53 352
rect 51 351 52 352
rect 50 351 51 352
rect 49 351 50 352
rect 48 351 49 352
rect 47 351 48 352
rect 46 351 47 352
rect 45 351 46 352
rect 44 351 45 352
rect 43 351 44 352
rect 42 351 43 352
rect 41 351 42 352
rect 40 351 41 352
rect 39 351 40 352
rect 38 351 39 352
rect 37 351 38 352
rect 36 351 37 352
rect 35 351 36 352
rect 34 351 35 352
rect 33 351 34 352
rect 32 351 33 352
rect 31 351 32 352
rect 30 351 31 352
rect 29 351 30 352
rect 28 351 29 352
rect 142 352 143 353
rect 141 352 142 353
rect 140 352 141 353
rect 139 352 140 353
rect 138 352 139 353
rect 137 352 138 353
rect 136 352 137 353
rect 135 352 136 353
rect 134 352 135 353
rect 133 352 134 353
rect 132 352 133 353
rect 131 352 132 353
rect 130 352 131 353
rect 129 352 130 353
rect 128 352 129 353
rect 127 352 128 353
rect 126 352 127 353
rect 125 352 126 353
rect 124 352 125 353
rect 123 352 124 353
rect 122 352 123 353
rect 121 352 122 353
rect 120 352 121 353
rect 119 352 120 353
rect 118 352 119 353
rect 117 352 118 353
rect 116 352 117 353
rect 115 352 116 353
rect 69 352 70 353
rect 68 352 69 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 60 352 61 353
rect 59 352 60 353
rect 58 352 59 353
rect 57 352 58 353
rect 56 352 57 353
rect 55 352 56 353
rect 54 352 55 353
rect 53 352 54 353
rect 52 352 53 353
rect 51 352 52 353
rect 50 352 51 353
rect 49 352 50 353
rect 48 352 49 353
rect 47 352 48 353
rect 46 352 47 353
rect 45 352 46 353
rect 44 352 45 353
rect 43 352 44 353
rect 42 352 43 353
rect 41 352 42 353
rect 40 352 41 353
rect 39 352 40 353
rect 38 352 39 353
rect 37 352 38 353
rect 36 352 37 353
rect 35 352 36 353
rect 34 352 35 353
rect 33 352 34 353
rect 32 352 33 353
rect 31 352 32 353
rect 30 352 31 353
rect 29 352 30 353
rect 28 352 29 353
rect 27 352 28 353
rect 26 352 27 353
rect 71 353 72 354
rect 70 353 71 354
rect 69 353 70 354
rect 68 353 69 354
rect 67 353 68 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 61 353 62 354
rect 60 353 61 354
rect 59 353 60 354
rect 58 353 59 354
rect 57 353 58 354
rect 56 353 57 354
rect 55 353 56 354
rect 54 353 55 354
rect 53 353 54 354
rect 52 353 53 354
rect 51 353 52 354
rect 50 353 51 354
rect 49 353 50 354
rect 48 353 49 354
rect 47 353 48 354
rect 46 353 47 354
rect 45 353 46 354
rect 44 353 45 354
rect 43 353 44 354
rect 42 353 43 354
rect 41 353 42 354
rect 40 353 41 354
rect 39 353 40 354
rect 38 353 39 354
rect 37 353 38 354
rect 36 353 37 354
rect 35 353 36 354
rect 34 353 35 354
rect 33 353 34 354
rect 32 353 33 354
rect 31 353 32 354
rect 30 353 31 354
rect 29 353 30 354
rect 28 353 29 354
rect 27 353 28 354
rect 26 353 27 354
rect 25 353 26 354
rect 24 353 25 354
rect 73 354 74 355
rect 72 354 73 355
rect 71 354 72 355
rect 70 354 71 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 62 354 63 355
rect 61 354 62 355
rect 60 354 61 355
rect 59 354 60 355
rect 58 354 59 355
rect 57 354 58 355
rect 56 354 57 355
rect 55 354 56 355
rect 54 354 55 355
rect 53 354 54 355
rect 52 354 53 355
rect 51 354 52 355
rect 50 354 51 355
rect 49 354 50 355
rect 48 354 49 355
rect 47 354 48 355
rect 46 354 47 355
rect 45 354 46 355
rect 44 354 45 355
rect 43 354 44 355
rect 42 354 43 355
rect 41 354 42 355
rect 40 354 41 355
rect 39 354 40 355
rect 38 354 39 355
rect 37 354 38 355
rect 36 354 37 355
rect 35 354 36 355
rect 34 354 35 355
rect 33 354 34 355
rect 32 354 33 355
rect 31 354 32 355
rect 30 354 31 355
rect 29 354 30 355
rect 28 354 29 355
rect 27 354 28 355
rect 26 354 27 355
rect 25 354 26 355
rect 24 354 25 355
rect 23 354 24 355
rect 74 355 75 356
rect 73 355 74 356
rect 72 355 73 356
rect 71 355 72 356
rect 70 355 71 356
rect 69 355 70 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 63 355 64 356
rect 62 355 63 356
rect 61 355 62 356
rect 60 355 61 356
rect 59 355 60 356
rect 58 355 59 356
rect 57 355 58 356
rect 56 355 57 356
rect 55 355 56 356
rect 54 355 55 356
rect 53 355 54 356
rect 52 355 53 356
rect 51 355 52 356
rect 50 355 51 356
rect 49 355 50 356
rect 48 355 49 356
rect 47 355 48 356
rect 46 355 47 356
rect 45 355 46 356
rect 44 355 45 356
rect 43 355 44 356
rect 42 355 43 356
rect 41 355 42 356
rect 40 355 41 356
rect 39 355 40 356
rect 38 355 39 356
rect 37 355 38 356
rect 36 355 37 356
rect 35 355 36 356
rect 34 355 35 356
rect 33 355 34 356
rect 32 355 33 356
rect 31 355 32 356
rect 30 355 31 356
rect 29 355 30 356
rect 28 355 29 356
rect 27 355 28 356
rect 26 355 27 356
rect 25 355 26 356
rect 24 355 25 356
rect 23 355 24 356
rect 22 355 23 356
rect 75 356 76 357
rect 74 356 75 357
rect 73 356 74 357
rect 72 356 73 357
rect 71 356 72 357
rect 70 356 71 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 64 356 65 357
rect 63 356 64 357
rect 62 356 63 357
rect 61 356 62 357
rect 60 356 61 357
rect 59 356 60 357
rect 58 356 59 357
rect 57 356 58 357
rect 56 356 57 357
rect 55 356 56 357
rect 54 356 55 357
rect 53 356 54 357
rect 52 356 53 357
rect 51 356 52 357
rect 50 356 51 357
rect 49 356 50 357
rect 48 356 49 357
rect 47 356 48 357
rect 46 356 47 357
rect 45 356 46 357
rect 44 356 45 357
rect 43 356 44 357
rect 42 356 43 357
rect 41 356 42 357
rect 40 356 41 357
rect 39 356 40 357
rect 38 356 39 357
rect 37 356 38 357
rect 36 356 37 357
rect 35 356 36 357
rect 34 356 35 357
rect 33 356 34 357
rect 32 356 33 357
rect 31 356 32 357
rect 30 356 31 357
rect 29 356 30 357
rect 28 356 29 357
rect 27 356 28 357
rect 26 356 27 357
rect 25 356 26 357
rect 24 356 25 357
rect 23 356 24 357
rect 22 356 23 357
rect 21 356 22 357
rect 20 356 21 357
rect 76 357 77 358
rect 75 357 76 358
rect 74 357 75 358
rect 73 357 74 358
rect 72 357 73 358
rect 71 357 72 358
rect 70 357 71 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 65 357 66 358
rect 64 357 65 358
rect 63 357 64 358
rect 62 357 63 358
rect 61 357 62 358
rect 60 357 61 358
rect 59 357 60 358
rect 58 357 59 358
rect 57 357 58 358
rect 56 357 57 358
rect 55 357 56 358
rect 54 357 55 358
rect 53 357 54 358
rect 52 357 53 358
rect 51 357 52 358
rect 50 357 51 358
rect 49 357 50 358
rect 48 357 49 358
rect 47 357 48 358
rect 46 357 47 358
rect 45 357 46 358
rect 44 357 45 358
rect 43 357 44 358
rect 42 357 43 358
rect 41 357 42 358
rect 40 357 41 358
rect 39 357 40 358
rect 38 357 39 358
rect 37 357 38 358
rect 36 357 37 358
rect 35 357 36 358
rect 34 357 35 358
rect 33 357 34 358
rect 32 357 33 358
rect 31 357 32 358
rect 30 357 31 358
rect 29 357 30 358
rect 28 357 29 358
rect 27 357 28 358
rect 26 357 27 358
rect 25 357 26 358
rect 24 357 25 358
rect 23 357 24 358
rect 22 357 23 358
rect 21 357 22 358
rect 20 357 21 358
rect 19 357 20 358
rect 77 358 78 359
rect 76 358 77 359
rect 75 358 76 359
rect 74 358 75 359
rect 73 358 74 359
rect 72 358 73 359
rect 71 358 72 359
rect 70 358 71 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 66 358 67 359
rect 65 358 66 359
rect 64 358 65 359
rect 63 358 64 359
rect 62 358 63 359
rect 61 358 62 359
rect 60 358 61 359
rect 59 358 60 359
rect 58 358 59 359
rect 57 358 58 359
rect 56 358 57 359
rect 55 358 56 359
rect 54 358 55 359
rect 53 358 54 359
rect 52 358 53 359
rect 51 358 52 359
rect 50 358 51 359
rect 49 358 50 359
rect 48 358 49 359
rect 47 358 48 359
rect 46 358 47 359
rect 45 358 46 359
rect 44 358 45 359
rect 43 358 44 359
rect 42 358 43 359
rect 41 358 42 359
rect 40 358 41 359
rect 39 358 40 359
rect 38 358 39 359
rect 37 358 38 359
rect 36 358 37 359
rect 35 358 36 359
rect 34 358 35 359
rect 33 358 34 359
rect 32 358 33 359
rect 31 358 32 359
rect 30 358 31 359
rect 29 358 30 359
rect 28 358 29 359
rect 27 358 28 359
rect 26 358 27 359
rect 25 358 26 359
rect 24 358 25 359
rect 23 358 24 359
rect 22 358 23 359
rect 21 358 22 359
rect 20 358 21 359
rect 19 358 20 359
rect 18 358 19 359
rect 142 359 143 360
rect 141 359 142 360
rect 140 359 141 360
rect 139 359 140 360
rect 138 359 139 360
rect 137 359 138 360
rect 136 359 137 360
rect 135 359 136 360
rect 134 359 135 360
rect 133 359 134 360
rect 132 359 133 360
rect 131 359 132 360
rect 130 359 131 360
rect 129 359 130 360
rect 128 359 129 360
rect 127 359 128 360
rect 126 359 127 360
rect 125 359 126 360
rect 124 359 125 360
rect 123 359 124 360
rect 122 359 123 360
rect 121 359 122 360
rect 120 359 121 360
rect 119 359 120 360
rect 118 359 119 360
rect 117 359 118 360
rect 77 359 78 360
rect 76 359 77 360
rect 75 359 76 360
rect 74 359 75 360
rect 73 359 74 360
rect 72 359 73 360
rect 71 359 72 360
rect 70 359 71 360
rect 69 359 70 360
rect 68 359 69 360
rect 67 359 68 360
rect 66 359 67 360
rect 65 359 66 360
rect 64 359 65 360
rect 63 359 64 360
rect 62 359 63 360
rect 61 359 62 360
rect 60 359 61 360
rect 59 359 60 360
rect 58 359 59 360
rect 57 359 58 360
rect 56 359 57 360
rect 55 359 56 360
rect 54 359 55 360
rect 53 359 54 360
rect 52 359 53 360
rect 51 359 52 360
rect 50 359 51 360
rect 49 359 50 360
rect 48 359 49 360
rect 47 359 48 360
rect 46 359 47 360
rect 45 359 46 360
rect 44 359 45 360
rect 43 359 44 360
rect 42 359 43 360
rect 41 359 42 360
rect 40 359 41 360
rect 39 359 40 360
rect 38 359 39 360
rect 37 359 38 360
rect 36 359 37 360
rect 35 359 36 360
rect 34 359 35 360
rect 33 359 34 360
rect 32 359 33 360
rect 31 359 32 360
rect 30 359 31 360
rect 29 359 30 360
rect 28 359 29 360
rect 27 359 28 360
rect 26 359 27 360
rect 25 359 26 360
rect 24 359 25 360
rect 23 359 24 360
rect 22 359 23 360
rect 21 359 22 360
rect 20 359 21 360
rect 19 359 20 360
rect 18 359 19 360
rect 142 360 143 361
rect 141 360 142 361
rect 140 360 141 361
rect 139 360 140 361
rect 138 360 139 361
rect 137 360 138 361
rect 136 360 137 361
rect 135 360 136 361
rect 134 360 135 361
rect 133 360 134 361
rect 132 360 133 361
rect 131 360 132 361
rect 130 360 131 361
rect 129 360 130 361
rect 128 360 129 361
rect 127 360 128 361
rect 126 360 127 361
rect 125 360 126 361
rect 124 360 125 361
rect 123 360 124 361
rect 122 360 123 361
rect 121 360 122 361
rect 120 360 121 361
rect 119 360 120 361
rect 118 360 119 361
rect 117 360 118 361
rect 78 360 79 361
rect 77 360 78 361
rect 76 360 77 361
rect 75 360 76 361
rect 74 360 75 361
rect 73 360 74 361
rect 72 360 73 361
rect 71 360 72 361
rect 70 360 71 361
rect 69 360 70 361
rect 68 360 69 361
rect 67 360 68 361
rect 66 360 67 361
rect 65 360 66 361
rect 64 360 65 361
rect 63 360 64 361
rect 62 360 63 361
rect 61 360 62 361
rect 60 360 61 361
rect 59 360 60 361
rect 58 360 59 361
rect 57 360 58 361
rect 56 360 57 361
rect 55 360 56 361
rect 54 360 55 361
rect 53 360 54 361
rect 52 360 53 361
rect 51 360 52 361
rect 50 360 51 361
rect 49 360 50 361
rect 48 360 49 361
rect 47 360 48 361
rect 46 360 47 361
rect 45 360 46 361
rect 44 360 45 361
rect 43 360 44 361
rect 42 360 43 361
rect 41 360 42 361
rect 40 360 41 361
rect 39 360 40 361
rect 38 360 39 361
rect 37 360 38 361
rect 36 360 37 361
rect 35 360 36 361
rect 34 360 35 361
rect 33 360 34 361
rect 32 360 33 361
rect 31 360 32 361
rect 30 360 31 361
rect 29 360 30 361
rect 28 360 29 361
rect 27 360 28 361
rect 26 360 27 361
rect 25 360 26 361
rect 24 360 25 361
rect 23 360 24 361
rect 22 360 23 361
rect 21 360 22 361
rect 20 360 21 361
rect 19 360 20 361
rect 18 360 19 361
rect 17 360 18 361
rect 142 361 143 362
rect 141 361 142 362
rect 140 361 141 362
rect 139 361 140 362
rect 138 361 139 362
rect 137 361 138 362
rect 136 361 137 362
rect 135 361 136 362
rect 134 361 135 362
rect 133 361 134 362
rect 132 361 133 362
rect 131 361 132 362
rect 130 361 131 362
rect 129 361 130 362
rect 128 361 129 362
rect 127 361 128 362
rect 126 361 127 362
rect 125 361 126 362
rect 124 361 125 362
rect 123 361 124 362
rect 122 361 123 362
rect 121 361 122 362
rect 120 361 121 362
rect 119 361 120 362
rect 118 361 119 362
rect 117 361 118 362
rect 78 361 79 362
rect 77 361 78 362
rect 76 361 77 362
rect 75 361 76 362
rect 74 361 75 362
rect 73 361 74 362
rect 72 361 73 362
rect 71 361 72 362
rect 70 361 71 362
rect 69 361 70 362
rect 68 361 69 362
rect 67 361 68 362
rect 66 361 67 362
rect 65 361 66 362
rect 64 361 65 362
rect 63 361 64 362
rect 62 361 63 362
rect 61 361 62 362
rect 60 361 61 362
rect 59 361 60 362
rect 58 361 59 362
rect 57 361 58 362
rect 56 361 57 362
rect 55 361 56 362
rect 54 361 55 362
rect 53 361 54 362
rect 52 361 53 362
rect 51 361 52 362
rect 50 361 51 362
rect 49 361 50 362
rect 48 361 49 362
rect 47 361 48 362
rect 46 361 47 362
rect 45 361 46 362
rect 44 361 45 362
rect 43 361 44 362
rect 42 361 43 362
rect 41 361 42 362
rect 40 361 41 362
rect 39 361 40 362
rect 38 361 39 362
rect 37 361 38 362
rect 36 361 37 362
rect 35 361 36 362
rect 34 361 35 362
rect 33 361 34 362
rect 32 361 33 362
rect 31 361 32 362
rect 30 361 31 362
rect 29 361 30 362
rect 28 361 29 362
rect 27 361 28 362
rect 26 361 27 362
rect 25 361 26 362
rect 24 361 25 362
rect 23 361 24 362
rect 22 361 23 362
rect 21 361 22 362
rect 20 361 21 362
rect 19 361 20 362
rect 18 361 19 362
rect 17 361 18 362
rect 16 361 17 362
rect 142 362 143 363
rect 141 362 142 363
rect 140 362 141 363
rect 139 362 140 363
rect 138 362 139 363
rect 137 362 138 363
rect 136 362 137 363
rect 135 362 136 363
rect 134 362 135 363
rect 133 362 134 363
rect 132 362 133 363
rect 131 362 132 363
rect 130 362 131 363
rect 129 362 130 363
rect 128 362 129 363
rect 127 362 128 363
rect 126 362 127 363
rect 125 362 126 363
rect 124 362 125 363
rect 123 362 124 363
rect 122 362 123 363
rect 121 362 122 363
rect 120 362 121 363
rect 119 362 120 363
rect 118 362 119 363
rect 117 362 118 363
rect 79 362 80 363
rect 78 362 79 363
rect 77 362 78 363
rect 76 362 77 363
rect 75 362 76 363
rect 74 362 75 363
rect 73 362 74 363
rect 72 362 73 363
rect 71 362 72 363
rect 70 362 71 363
rect 69 362 70 363
rect 68 362 69 363
rect 67 362 68 363
rect 66 362 67 363
rect 65 362 66 363
rect 64 362 65 363
rect 63 362 64 363
rect 62 362 63 363
rect 61 362 62 363
rect 60 362 61 363
rect 59 362 60 363
rect 58 362 59 363
rect 57 362 58 363
rect 56 362 57 363
rect 55 362 56 363
rect 54 362 55 363
rect 53 362 54 363
rect 52 362 53 363
rect 51 362 52 363
rect 50 362 51 363
rect 49 362 50 363
rect 48 362 49 363
rect 47 362 48 363
rect 46 362 47 363
rect 45 362 46 363
rect 44 362 45 363
rect 43 362 44 363
rect 42 362 43 363
rect 41 362 42 363
rect 40 362 41 363
rect 39 362 40 363
rect 38 362 39 363
rect 37 362 38 363
rect 36 362 37 363
rect 35 362 36 363
rect 34 362 35 363
rect 33 362 34 363
rect 32 362 33 363
rect 31 362 32 363
rect 30 362 31 363
rect 29 362 30 363
rect 28 362 29 363
rect 27 362 28 363
rect 26 362 27 363
rect 25 362 26 363
rect 24 362 25 363
rect 23 362 24 363
rect 22 362 23 363
rect 21 362 22 363
rect 20 362 21 363
rect 19 362 20 363
rect 18 362 19 363
rect 17 362 18 363
rect 16 362 17 363
rect 142 363 143 364
rect 141 363 142 364
rect 140 363 141 364
rect 139 363 140 364
rect 138 363 139 364
rect 137 363 138 364
rect 136 363 137 364
rect 135 363 136 364
rect 134 363 135 364
rect 133 363 134 364
rect 132 363 133 364
rect 131 363 132 364
rect 130 363 131 364
rect 129 363 130 364
rect 128 363 129 364
rect 127 363 128 364
rect 126 363 127 364
rect 125 363 126 364
rect 124 363 125 364
rect 123 363 124 364
rect 122 363 123 364
rect 121 363 122 364
rect 120 363 121 364
rect 119 363 120 364
rect 118 363 119 364
rect 117 363 118 364
rect 79 363 80 364
rect 78 363 79 364
rect 77 363 78 364
rect 76 363 77 364
rect 75 363 76 364
rect 74 363 75 364
rect 73 363 74 364
rect 72 363 73 364
rect 71 363 72 364
rect 70 363 71 364
rect 69 363 70 364
rect 68 363 69 364
rect 67 363 68 364
rect 66 363 67 364
rect 65 363 66 364
rect 64 363 65 364
rect 63 363 64 364
rect 62 363 63 364
rect 61 363 62 364
rect 60 363 61 364
rect 59 363 60 364
rect 58 363 59 364
rect 57 363 58 364
rect 56 363 57 364
rect 55 363 56 364
rect 54 363 55 364
rect 53 363 54 364
rect 52 363 53 364
rect 51 363 52 364
rect 50 363 51 364
rect 49 363 50 364
rect 48 363 49 364
rect 47 363 48 364
rect 46 363 47 364
rect 45 363 46 364
rect 44 363 45 364
rect 43 363 44 364
rect 42 363 43 364
rect 41 363 42 364
rect 40 363 41 364
rect 39 363 40 364
rect 38 363 39 364
rect 37 363 38 364
rect 36 363 37 364
rect 35 363 36 364
rect 34 363 35 364
rect 33 363 34 364
rect 32 363 33 364
rect 31 363 32 364
rect 30 363 31 364
rect 29 363 30 364
rect 28 363 29 364
rect 27 363 28 364
rect 26 363 27 364
rect 25 363 26 364
rect 24 363 25 364
rect 23 363 24 364
rect 22 363 23 364
rect 21 363 22 364
rect 20 363 21 364
rect 19 363 20 364
rect 18 363 19 364
rect 17 363 18 364
rect 16 363 17 364
rect 15 363 16 364
rect 130 364 131 365
rect 129 364 130 365
rect 128 364 129 365
rect 80 364 81 365
rect 79 364 80 365
rect 78 364 79 365
rect 77 364 78 365
rect 76 364 77 365
rect 75 364 76 365
rect 74 364 75 365
rect 73 364 74 365
rect 72 364 73 365
rect 71 364 72 365
rect 70 364 71 365
rect 69 364 70 365
rect 68 364 69 365
rect 67 364 68 365
rect 66 364 67 365
rect 65 364 66 365
rect 64 364 65 365
rect 63 364 64 365
rect 62 364 63 365
rect 61 364 62 365
rect 60 364 61 365
rect 59 364 60 365
rect 58 364 59 365
rect 57 364 58 365
rect 56 364 57 365
rect 55 364 56 365
rect 54 364 55 365
rect 53 364 54 365
rect 52 364 53 365
rect 51 364 52 365
rect 50 364 51 365
rect 49 364 50 365
rect 48 364 49 365
rect 47 364 48 365
rect 46 364 47 365
rect 45 364 46 365
rect 44 364 45 365
rect 43 364 44 365
rect 42 364 43 365
rect 41 364 42 365
rect 40 364 41 365
rect 39 364 40 365
rect 38 364 39 365
rect 37 364 38 365
rect 36 364 37 365
rect 35 364 36 365
rect 34 364 35 365
rect 33 364 34 365
rect 32 364 33 365
rect 31 364 32 365
rect 30 364 31 365
rect 29 364 30 365
rect 28 364 29 365
rect 27 364 28 365
rect 26 364 27 365
rect 25 364 26 365
rect 24 364 25 365
rect 23 364 24 365
rect 22 364 23 365
rect 21 364 22 365
rect 20 364 21 365
rect 19 364 20 365
rect 18 364 19 365
rect 17 364 18 365
rect 16 364 17 365
rect 15 364 16 365
rect 131 365 132 366
rect 130 365 131 366
rect 129 365 130 366
rect 128 365 129 366
rect 80 365 81 366
rect 79 365 80 366
rect 78 365 79 366
rect 77 365 78 366
rect 76 365 77 366
rect 75 365 76 366
rect 74 365 75 366
rect 73 365 74 366
rect 72 365 73 366
rect 71 365 72 366
rect 70 365 71 366
rect 69 365 70 366
rect 68 365 69 366
rect 67 365 68 366
rect 66 365 67 366
rect 65 365 66 366
rect 64 365 65 366
rect 63 365 64 366
rect 62 365 63 366
rect 61 365 62 366
rect 60 365 61 366
rect 59 365 60 366
rect 58 365 59 366
rect 57 365 58 366
rect 56 365 57 366
rect 55 365 56 366
rect 54 365 55 366
rect 53 365 54 366
rect 52 365 53 366
rect 51 365 52 366
rect 50 365 51 366
rect 49 365 50 366
rect 48 365 49 366
rect 47 365 48 366
rect 46 365 47 366
rect 45 365 46 366
rect 44 365 45 366
rect 43 365 44 366
rect 42 365 43 366
rect 41 365 42 366
rect 40 365 41 366
rect 39 365 40 366
rect 38 365 39 366
rect 37 365 38 366
rect 36 365 37 366
rect 35 365 36 366
rect 34 365 35 366
rect 33 365 34 366
rect 32 365 33 366
rect 31 365 32 366
rect 30 365 31 366
rect 29 365 30 366
rect 28 365 29 366
rect 27 365 28 366
rect 26 365 27 366
rect 25 365 26 366
rect 24 365 25 366
rect 23 365 24 366
rect 22 365 23 366
rect 21 365 22 366
rect 20 365 21 366
rect 19 365 20 366
rect 18 365 19 366
rect 17 365 18 366
rect 16 365 17 366
rect 15 365 16 366
rect 132 366 133 367
rect 131 366 132 367
rect 130 366 131 367
rect 129 366 130 367
rect 128 366 129 367
rect 127 366 128 367
rect 126 366 127 367
rect 80 366 81 367
rect 79 366 80 367
rect 78 366 79 367
rect 77 366 78 367
rect 76 366 77 367
rect 75 366 76 367
rect 74 366 75 367
rect 73 366 74 367
rect 72 366 73 367
rect 71 366 72 367
rect 70 366 71 367
rect 69 366 70 367
rect 68 366 69 367
rect 67 366 68 367
rect 66 366 67 367
rect 65 366 66 367
rect 64 366 65 367
rect 63 366 64 367
rect 62 366 63 367
rect 61 366 62 367
rect 60 366 61 367
rect 59 366 60 367
rect 58 366 59 367
rect 57 366 58 367
rect 56 366 57 367
rect 55 366 56 367
rect 54 366 55 367
rect 53 366 54 367
rect 52 366 53 367
rect 51 366 52 367
rect 50 366 51 367
rect 49 366 50 367
rect 48 366 49 367
rect 47 366 48 367
rect 46 366 47 367
rect 45 366 46 367
rect 44 366 45 367
rect 43 366 44 367
rect 42 366 43 367
rect 41 366 42 367
rect 40 366 41 367
rect 39 366 40 367
rect 38 366 39 367
rect 37 366 38 367
rect 36 366 37 367
rect 35 366 36 367
rect 34 366 35 367
rect 33 366 34 367
rect 32 366 33 367
rect 31 366 32 367
rect 30 366 31 367
rect 29 366 30 367
rect 28 366 29 367
rect 27 366 28 367
rect 26 366 27 367
rect 25 366 26 367
rect 24 366 25 367
rect 23 366 24 367
rect 22 366 23 367
rect 21 366 22 367
rect 20 366 21 367
rect 19 366 20 367
rect 18 366 19 367
rect 17 366 18 367
rect 16 366 17 367
rect 15 366 16 367
rect 14 366 15 367
rect 134 367 135 368
rect 133 367 134 368
rect 132 367 133 368
rect 131 367 132 368
rect 130 367 131 368
rect 129 367 130 368
rect 128 367 129 368
rect 127 367 128 368
rect 126 367 127 368
rect 125 367 126 368
rect 80 367 81 368
rect 79 367 80 368
rect 78 367 79 368
rect 77 367 78 368
rect 76 367 77 368
rect 75 367 76 368
rect 74 367 75 368
rect 73 367 74 368
rect 72 367 73 368
rect 71 367 72 368
rect 70 367 71 368
rect 69 367 70 368
rect 68 367 69 368
rect 67 367 68 368
rect 66 367 67 368
rect 65 367 66 368
rect 64 367 65 368
rect 63 367 64 368
rect 62 367 63 368
rect 61 367 62 368
rect 60 367 61 368
rect 59 367 60 368
rect 58 367 59 368
rect 57 367 58 368
rect 56 367 57 368
rect 55 367 56 368
rect 54 367 55 368
rect 53 367 54 368
rect 52 367 53 368
rect 51 367 52 368
rect 50 367 51 368
rect 49 367 50 368
rect 48 367 49 368
rect 47 367 48 368
rect 46 367 47 368
rect 45 367 46 368
rect 44 367 45 368
rect 43 367 44 368
rect 42 367 43 368
rect 41 367 42 368
rect 40 367 41 368
rect 39 367 40 368
rect 38 367 39 368
rect 37 367 38 368
rect 36 367 37 368
rect 35 367 36 368
rect 34 367 35 368
rect 33 367 34 368
rect 32 367 33 368
rect 31 367 32 368
rect 30 367 31 368
rect 29 367 30 368
rect 28 367 29 368
rect 27 367 28 368
rect 26 367 27 368
rect 25 367 26 368
rect 24 367 25 368
rect 23 367 24 368
rect 22 367 23 368
rect 21 367 22 368
rect 20 367 21 368
rect 19 367 20 368
rect 18 367 19 368
rect 17 367 18 368
rect 16 367 17 368
rect 15 367 16 368
rect 14 367 15 368
rect 135 368 136 369
rect 134 368 135 369
rect 133 368 134 369
rect 132 368 133 369
rect 131 368 132 369
rect 130 368 131 369
rect 129 368 130 369
rect 128 368 129 369
rect 127 368 128 369
rect 126 368 127 369
rect 125 368 126 369
rect 124 368 125 369
rect 123 368 124 369
rect 81 368 82 369
rect 80 368 81 369
rect 79 368 80 369
rect 78 368 79 369
rect 77 368 78 369
rect 76 368 77 369
rect 75 368 76 369
rect 74 368 75 369
rect 73 368 74 369
rect 72 368 73 369
rect 71 368 72 369
rect 70 368 71 369
rect 69 368 70 369
rect 68 368 69 369
rect 67 368 68 369
rect 66 368 67 369
rect 65 368 66 369
rect 64 368 65 369
rect 63 368 64 369
rect 62 368 63 369
rect 61 368 62 369
rect 60 368 61 369
rect 59 368 60 369
rect 58 368 59 369
rect 37 368 38 369
rect 36 368 37 369
rect 35 368 36 369
rect 34 368 35 369
rect 33 368 34 369
rect 32 368 33 369
rect 31 368 32 369
rect 30 368 31 369
rect 29 368 30 369
rect 28 368 29 369
rect 27 368 28 369
rect 26 368 27 369
rect 25 368 26 369
rect 24 368 25 369
rect 23 368 24 369
rect 22 368 23 369
rect 21 368 22 369
rect 20 368 21 369
rect 19 368 20 369
rect 18 368 19 369
rect 17 368 18 369
rect 16 368 17 369
rect 15 368 16 369
rect 14 368 15 369
rect 137 369 138 370
rect 136 369 137 370
rect 135 369 136 370
rect 134 369 135 370
rect 133 369 134 370
rect 132 369 133 370
rect 131 369 132 370
rect 130 369 131 370
rect 129 369 130 370
rect 128 369 129 370
rect 127 369 128 370
rect 126 369 127 370
rect 125 369 126 370
rect 124 369 125 370
rect 123 369 124 370
rect 122 369 123 370
rect 81 369 82 370
rect 80 369 81 370
rect 79 369 80 370
rect 78 369 79 370
rect 77 369 78 370
rect 76 369 77 370
rect 75 369 76 370
rect 74 369 75 370
rect 73 369 74 370
rect 72 369 73 370
rect 71 369 72 370
rect 70 369 71 370
rect 69 369 70 370
rect 68 369 69 370
rect 67 369 68 370
rect 66 369 67 370
rect 65 369 66 370
rect 64 369 65 370
rect 63 369 64 370
rect 32 369 33 370
rect 31 369 32 370
rect 30 369 31 370
rect 29 369 30 370
rect 28 369 29 370
rect 27 369 28 370
rect 26 369 27 370
rect 25 369 26 370
rect 24 369 25 370
rect 23 369 24 370
rect 22 369 23 370
rect 21 369 22 370
rect 20 369 21 370
rect 19 369 20 370
rect 18 369 19 370
rect 17 369 18 370
rect 16 369 17 370
rect 15 369 16 370
rect 14 369 15 370
rect 138 370 139 371
rect 137 370 138 371
rect 136 370 137 371
rect 135 370 136 371
rect 134 370 135 371
rect 133 370 134 371
rect 132 370 133 371
rect 131 370 132 371
rect 130 370 131 371
rect 129 370 130 371
rect 128 370 129 371
rect 127 370 128 371
rect 126 370 127 371
rect 125 370 126 371
rect 124 370 125 371
rect 123 370 124 371
rect 122 370 123 371
rect 121 370 122 371
rect 120 370 121 371
rect 81 370 82 371
rect 80 370 81 371
rect 79 370 80 371
rect 78 370 79 371
rect 77 370 78 371
rect 76 370 77 371
rect 75 370 76 371
rect 74 370 75 371
rect 73 370 74 371
rect 72 370 73 371
rect 71 370 72 371
rect 70 370 71 371
rect 69 370 70 371
rect 68 370 69 371
rect 67 370 68 371
rect 66 370 67 371
rect 65 370 66 371
rect 29 370 30 371
rect 28 370 29 371
rect 27 370 28 371
rect 26 370 27 371
rect 25 370 26 371
rect 24 370 25 371
rect 23 370 24 371
rect 22 370 23 371
rect 21 370 22 371
rect 20 370 21 371
rect 19 370 20 371
rect 18 370 19 371
rect 17 370 18 371
rect 16 370 17 371
rect 15 370 16 371
rect 14 370 15 371
rect 13 370 14 371
rect 140 371 141 372
rect 139 371 140 372
rect 138 371 139 372
rect 137 371 138 372
rect 136 371 137 372
rect 135 371 136 372
rect 134 371 135 372
rect 133 371 134 372
rect 132 371 133 372
rect 131 371 132 372
rect 127 371 128 372
rect 126 371 127 372
rect 125 371 126 372
rect 124 371 125 372
rect 123 371 124 372
rect 122 371 123 372
rect 121 371 122 372
rect 120 371 121 372
rect 119 371 120 372
rect 81 371 82 372
rect 80 371 81 372
rect 79 371 80 372
rect 78 371 79 372
rect 77 371 78 372
rect 76 371 77 372
rect 75 371 76 372
rect 74 371 75 372
rect 73 371 74 372
rect 72 371 73 372
rect 71 371 72 372
rect 70 371 71 372
rect 69 371 70 372
rect 68 371 69 372
rect 67 371 68 372
rect 66 371 67 372
rect 28 371 29 372
rect 27 371 28 372
rect 26 371 27 372
rect 25 371 26 372
rect 24 371 25 372
rect 23 371 24 372
rect 22 371 23 372
rect 21 371 22 372
rect 20 371 21 372
rect 19 371 20 372
rect 18 371 19 372
rect 17 371 18 372
rect 16 371 17 372
rect 15 371 16 372
rect 14 371 15 372
rect 13 371 14 372
rect 141 372 142 373
rect 140 372 141 373
rect 139 372 140 373
rect 138 372 139 373
rect 137 372 138 373
rect 136 372 137 373
rect 135 372 136 373
rect 134 372 135 373
rect 133 372 134 373
rect 132 372 133 373
rect 126 372 127 373
rect 125 372 126 373
rect 124 372 125 373
rect 123 372 124 373
rect 122 372 123 373
rect 121 372 122 373
rect 120 372 121 373
rect 119 372 120 373
rect 118 372 119 373
rect 117 372 118 373
rect 81 372 82 373
rect 80 372 81 373
rect 79 372 80 373
rect 78 372 79 373
rect 77 372 78 373
rect 76 372 77 373
rect 75 372 76 373
rect 74 372 75 373
rect 73 372 74 373
rect 72 372 73 373
rect 71 372 72 373
rect 70 372 71 373
rect 69 372 70 373
rect 68 372 69 373
rect 67 372 68 373
rect 27 372 28 373
rect 26 372 27 373
rect 25 372 26 373
rect 24 372 25 373
rect 23 372 24 373
rect 22 372 23 373
rect 21 372 22 373
rect 20 372 21 373
rect 19 372 20 373
rect 18 372 19 373
rect 17 372 18 373
rect 16 372 17 373
rect 15 372 16 373
rect 14 372 15 373
rect 13 372 14 373
rect 142 373 143 374
rect 141 373 142 374
rect 140 373 141 374
rect 139 373 140 374
rect 138 373 139 374
rect 137 373 138 374
rect 136 373 137 374
rect 135 373 136 374
rect 134 373 135 374
rect 124 373 125 374
rect 123 373 124 374
rect 122 373 123 374
rect 121 373 122 374
rect 120 373 121 374
rect 119 373 120 374
rect 118 373 119 374
rect 117 373 118 374
rect 81 373 82 374
rect 80 373 81 374
rect 79 373 80 374
rect 78 373 79 374
rect 77 373 78 374
rect 76 373 77 374
rect 75 373 76 374
rect 74 373 75 374
rect 73 373 74 374
rect 72 373 73 374
rect 71 373 72 374
rect 70 373 71 374
rect 69 373 70 374
rect 68 373 69 374
rect 67 373 68 374
rect 27 373 28 374
rect 26 373 27 374
rect 25 373 26 374
rect 24 373 25 374
rect 23 373 24 374
rect 22 373 23 374
rect 21 373 22 374
rect 20 373 21 374
rect 19 373 20 374
rect 18 373 19 374
rect 17 373 18 374
rect 16 373 17 374
rect 15 373 16 374
rect 14 373 15 374
rect 13 373 14 374
rect 142 374 143 375
rect 141 374 142 375
rect 140 374 141 375
rect 139 374 140 375
rect 138 374 139 375
rect 137 374 138 375
rect 136 374 137 375
rect 135 374 136 375
rect 123 374 124 375
rect 122 374 123 375
rect 121 374 122 375
rect 120 374 121 375
rect 119 374 120 375
rect 118 374 119 375
rect 117 374 118 375
rect 81 374 82 375
rect 80 374 81 375
rect 79 374 80 375
rect 78 374 79 375
rect 77 374 78 375
rect 76 374 77 375
rect 75 374 76 375
rect 74 374 75 375
rect 73 374 74 375
rect 72 374 73 375
rect 71 374 72 375
rect 70 374 71 375
rect 69 374 70 375
rect 68 374 69 375
rect 67 374 68 375
rect 27 374 28 375
rect 26 374 27 375
rect 25 374 26 375
rect 24 374 25 375
rect 23 374 24 375
rect 22 374 23 375
rect 21 374 22 375
rect 20 374 21 375
rect 19 374 20 375
rect 18 374 19 375
rect 17 374 18 375
rect 16 374 17 375
rect 15 374 16 375
rect 14 374 15 375
rect 13 374 14 375
rect 142 375 143 376
rect 141 375 142 376
rect 140 375 141 376
rect 139 375 140 376
rect 138 375 139 376
rect 137 375 138 376
rect 136 375 137 376
rect 121 375 122 376
rect 120 375 121 376
rect 119 375 120 376
rect 118 375 119 376
rect 117 375 118 376
rect 81 375 82 376
rect 80 375 81 376
rect 79 375 80 376
rect 78 375 79 376
rect 77 375 78 376
rect 76 375 77 376
rect 75 375 76 376
rect 74 375 75 376
rect 73 375 74 376
rect 72 375 73 376
rect 71 375 72 376
rect 70 375 71 376
rect 69 375 70 376
rect 68 375 69 376
rect 67 375 68 376
rect 27 375 28 376
rect 26 375 27 376
rect 25 375 26 376
rect 24 375 25 376
rect 23 375 24 376
rect 22 375 23 376
rect 21 375 22 376
rect 20 375 21 376
rect 19 375 20 376
rect 18 375 19 376
rect 17 375 18 376
rect 16 375 17 376
rect 15 375 16 376
rect 14 375 15 376
rect 13 375 14 376
rect 142 376 143 377
rect 141 376 142 377
rect 140 376 141 377
rect 139 376 140 377
rect 138 376 139 377
rect 120 376 121 377
rect 119 376 120 377
rect 118 376 119 377
rect 117 376 118 377
rect 81 376 82 377
rect 80 376 81 377
rect 79 376 80 377
rect 78 376 79 377
rect 77 376 78 377
rect 76 376 77 377
rect 75 376 76 377
rect 74 376 75 377
rect 73 376 74 377
rect 72 376 73 377
rect 71 376 72 377
rect 70 376 71 377
rect 69 376 70 377
rect 68 376 69 377
rect 67 376 68 377
rect 66 376 67 377
rect 28 376 29 377
rect 27 376 28 377
rect 26 376 27 377
rect 25 376 26 377
rect 24 376 25 377
rect 23 376 24 377
rect 22 376 23 377
rect 21 376 22 377
rect 20 376 21 377
rect 19 376 20 377
rect 18 376 19 377
rect 17 376 18 377
rect 16 376 17 377
rect 15 376 16 377
rect 14 376 15 377
rect 13 376 14 377
rect 142 377 143 378
rect 141 377 142 378
rect 140 377 141 378
rect 139 377 140 378
rect 119 377 120 378
rect 118 377 119 378
rect 117 377 118 378
rect 81 377 82 378
rect 80 377 81 378
rect 79 377 80 378
rect 78 377 79 378
rect 77 377 78 378
rect 76 377 77 378
rect 75 377 76 378
rect 74 377 75 378
rect 73 377 74 378
rect 72 377 73 378
rect 71 377 72 378
rect 70 377 71 378
rect 69 377 70 378
rect 68 377 69 378
rect 67 377 68 378
rect 66 377 67 378
rect 65 377 66 378
rect 29 377 30 378
rect 28 377 29 378
rect 27 377 28 378
rect 26 377 27 378
rect 25 377 26 378
rect 24 377 25 378
rect 23 377 24 378
rect 22 377 23 378
rect 21 377 22 378
rect 20 377 21 378
rect 19 377 20 378
rect 18 377 19 378
rect 17 377 18 378
rect 16 377 17 378
rect 15 377 16 378
rect 14 377 15 378
rect 13 377 14 378
rect 142 378 143 379
rect 141 378 142 379
rect 117 378 118 379
rect 81 378 82 379
rect 80 378 81 379
rect 79 378 80 379
rect 78 378 79 379
rect 77 378 78 379
rect 76 378 77 379
rect 75 378 76 379
rect 74 378 75 379
rect 73 378 74 379
rect 72 378 73 379
rect 71 378 72 379
rect 70 378 71 379
rect 69 378 70 379
rect 68 378 69 379
rect 67 378 68 379
rect 66 378 67 379
rect 65 378 66 379
rect 64 378 65 379
rect 63 378 64 379
rect 62 378 63 379
rect 31 378 32 379
rect 30 378 31 379
rect 29 378 30 379
rect 28 378 29 379
rect 27 378 28 379
rect 26 378 27 379
rect 25 378 26 379
rect 24 378 25 379
rect 23 378 24 379
rect 22 378 23 379
rect 21 378 22 379
rect 20 378 21 379
rect 19 378 20 379
rect 18 378 19 379
rect 17 378 18 379
rect 16 378 17 379
rect 15 378 16 379
rect 14 378 15 379
rect 13 378 14 379
rect 142 379 143 380
rect 80 379 81 380
rect 79 379 80 380
rect 78 379 79 380
rect 77 379 78 380
rect 76 379 77 380
rect 75 379 76 380
rect 74 379 75 380
rect 73 379 74 380
rect 72 379 73 380
rect 71 379 72 380
rect 70 379 71 380
rect 69 379 70 380
rect 68 379 69 380
rect 67 379 68 380
rect 66 379 67 380
rect 65 379 66 380
rect 64 379 65 380
rect 63 379 64 380
rect 62 379 63 380
rect 61 379 62 380
rect 60 379 61 380
rect 59 379 60 380
rect 58 379 59 380
rect 35 379 36 380
rect 34 379 35 380
rect 33 379 34 380
rect 32 379 33 380
rect 31 379 32 380
rect 30 379 31 380
rect 29 379 30 380
rect 28 379 29 380
rect 27 379 28 380
rect 26 379 27 380
rect 25 379 26 380
rect 24 379 25 380
rect 23 379 24 380
rect 22 379 23 380
rect 21 379 22 380
rect 20 379 21 380
rect 19 379 20 380
rect 18 379 19 380
rect 17 379 18 380
rect 16 379 17 380
rect 15 379 16 380
rect 14 379 15 380
rect 13 379 14 380
rect 80 380 81 381
rect 79 380 80 381
rect 78 380 79 381
rect 77 380 78 381
rect 76 380 77 381
rect 75 380 76 381
rect 74 380 75 381
rect 73 380 74 381
rect 72 380 73 381
rect 71 380 72 381
rect 70 380 71 381
rect 69 380 70 381
rect 68 380 69 381
rect 67 380 68 381
rect 66 380 67 381
rect 65 380 66 381
rect 64 380 65 381
rect 63 380 64 381
rect 62 380 63 381
rect 61 380 62 381
rect 60 380 61 381
rect 59 380 60 381
rect 58 380 59 381
rect 57 380 58 381
rect 56 380 57 381
rect 55 380 56 381
rect 54 380 55 381
rect 53 380 54 381
rect 52 380 53 381
rect 51 380 52 381
rect 50 380 51 381
rect 49 380 50 381
rect 48 380 49 381
rect 47 380 48 381
rect 46 380 47 381
rect 45 380 46 381
rect 44 380 45 381
rect 43 380 44 381
rect 42 380 43 381
rect 41 380 42 381
rect 40 380 41 381
rect 39 380 40 381
rect 38 380 39 381
rect 37 380 38 381
rect 36 380 37 381
rect 35 380 36 381
rect 34 380 35 381
rect 33 380 34 381
rect 32 380 33 381
rect 31 380 32 381
rect 30 380 31 381
rect 29 380 30 381
rect 28 380 29 381
rect 27 380 28 381
rect 26 380 27 381
rect 25 380 26 381
rect 24 380 25 381
rect 23 380 24 381
rect 22 380 23 381
rect 21 380 22 381
rect 20 380 21 381
rect 19 380 20 381
rect 18 380 19 381
rect 17 380 18 381
rect 16 380 17 381
rect 15 380 16 381
rect 14 380 15 381
rect 134 381 135 382
rect 133 381 134 382
rect 132 381 133 382
rect 80 381 81 382
rect 79 381 80 382
rect 78 381 79 382
rect 77 381 78 382
rect 76 381 77 382
rect 75 381 76 382
rect 74 381 75 382
rect 73 381 74 382
rect 72 381 73 382
rect 71 381 72 382
rect 70 381 71 382
rect 69 381 70 382
rect 68 381 69 382
rect 67 381 68 382
rect 66 381 67 382
rect 65 381 66 382
rect 64 381 65 382
rect 63 381 64 382
rect 62 381 63 382
rect 61 381 62 382
rect 60 381 61 382
rect 59 381 60 382
rect 58 381 59 382
rect 57 381 58 382
rect 56 381 57 382
rect 55 381 56 382
rect 54 381 55 382
rect 53 381 54 382
rect 52 381 53 382
rect 51 381 52 382
rect 50 381 51 382
rect 49 381 50 382
rect 48 381 49 382
rect 47 381 48 382
rect 46 381 47 382
rect 45 381 46 382
rect 44 381 45 382
rect 43 381 44 382
rect 42 381 43 382
rect 41 381 42 382
rect 40 381 41 382
rect 39 381 40 382
rect 38 381 39 382
rect 37 381 38 382
rect 36 381 37 382
rect 35 381 36 382
rect 34 381 35 382
rect 33 381 34 382
rect 32 381 33 382
rect 31 381 32 382
rect 30 381 31 382
rect 29 381 30 382
rect 28 381 29 382
rect 27 381 28 382
rect 26 381 27 382
rect 25 381 26 382
rect 24 381 25 382
rect 23 381 24 382
rect 22 381 23 382
rect 21 381 22 382
rect 20 381 21 382
rect 19 381 20 382
rect 18 381 19 382
rect 17 381 18 382
rect 16 381 17 382
rect 15 381 16 382
rect 14 381 15 382
rect 137 382 138 383
rect 136 382 137 383
rect 135 382 136 383
rect 134 382 135 383
rect 133 382 134 383
rect 132 382 133 383
rect 131 382 132 383
rect 130 382 131 383
rect 129 382 130 383
rect 80 382 81 383
rect 79 382 80 383
rect 78 382 79 383
rect 77 382 78 383
rect 76 382 77 383
rect 75 382 76 383
rect 74 382 75 383
rect 73 382 74 383
rect 72 382 73 383
rect 71 382 72 383
rect 70 382 71 383
rect 69 382 70 383
rect 68 382 69 383
rect 67 382 68 383
rect 66 382 67 383
rect 65 382 66 383
rect 64 382 65 383
rect 63 382 64 383
rect 62 382 63 383
rect 61 382 62 383
rect 60 382 61 383
rect 59 382 60 383
rect 58 382 59 383
rect 57 382 58 383
rect 56 382 57 383
rect 55 382 56 383
rect 54 382 55 383
rect 53 382 54 383
rect 52 382 53 383
rect 51 382 52 383
rect 50 382 51 383
rect 49 382 50 383
rect 48 382 49 383
rect 47 382 48 383
rect 46 382 47 383
rect 45 382 46 383
rect 44 382 45 383
rect 43 382 44 383
rect 42 382 43 383
rect 41 382 42 383
rect 40 382 41 383
rect 39 382 40 383
rect 38 382 39 383
rect 37 382 38 383
rect 36 382 37 383
rect 35 382 36 383
rect 34 382 35 383
rect 33 382 34 383
rect 32 382 33 383
rect 31 382 32 383
rect 30 382 31 383
rect 29 382 30 383
rect 28 382 29 383
rect 27 382 28 383
rect 26 382 27 383
rect 25 382 26 383
rect 24 382 25 383
rect 23 382 24 383
rect 22 382 23 383
rect 21 382 22 383
rect 20 382 21 383
rect 19 382 20 383
rect 18 382 19 383
rect 17 382 18 383
rect 16 382 17 383
rect 15 382 16 383
rect 14 382 15 383
rect 139 383 140 384
rect 138 383 139 384
rect 137 383 138 384
rect 136 383 137 384
rect 135 383 136 384
rect 134 383 135 384
rect 133 383 134 384
rect 132 383 133 384
rect 131 383 132 384
rect 130 383 131 384
rect 129 383 130 384
rect 128 383 129 384
rect 127 383 128 384
rect 79 383 80 384
rect 78 383 79 384
rect 77 383 78 384
rect 76 383 77 384
rect 75 383 76 384
rect 74 383 75 384
rect 73 383 74 384
rect 72 383 73 384
rect 71 383 72 384
rect 70 383 71 384
rect 69 383 70 384
rect 68 383 69 384
rect 67 383 68 384
rect 66 383 67 384
rect 65 383 66 384
rect 64 383 65 384
rect 63 383 64 384
rect 62 383 63 384
rect 61 383 62 384
rect 60 383 61 384
rect 59 383 60 384
rect 58 383 59 384
rect 57 383 58 384
rect 56 383 57 384
rect 55 383 56 384
rect 54 383 55 384
rect 53 383 54 384
rect 52 383 53 384
rect 51 383 52 384
rect 50 383 51 384
rect 49 383 50 384
rect 48 383 49 384
rect 47 383 48 384
rect 46 383 47 384
rect 45 383 46 384
rect 44 383 45 384
rect 43 383 44 384
rect 42 383 43 384
rect 41 383 42 384
rect 40 383 41 384
rect 39 383 40 384
rect 38 383 39 384
rect 37 383 38 384
rect 36 383 37 384
rect 35 383 36 384
rect 34 383 35 384
rect 33 383 34 384
rect 32 383 33 384
rect 31 383 32 384
rect 30 383 31 384
rect 29 383 30 384
rect 28 383 29 384
rect 27 383 28 384
rect 26 383 27 384
rect 25 383 26 384
rect 24 383 25 384
rect 23 383 24 384
rect 22 383 23 384
rect 21 383 22 384
rect 20 383 21 384
rect 19 383 20 384
rect 18 383 19 384
rect 17 383 18 384
rect 16 383 17 384
rect 15 383 16 384
rect 14 383 15 384
rect 140 384 141 385
rect 139 384 140 385
rect 138 384 139 385
rect 137 384 138 385
rect 136 384 137 385
rect 135 384 136 385
rect 134 384 135 385
rect 133 384 134 385
rect 132 384 133 385
rect 131 384 132 385
rect 130 384 131 385
rect 129 384 130 385
rect 128 384 129 385
rect 127 384 128 385
rect 126 384 127 385
rect 79 384 80 385
rect 78 384 79 385
rect 77 384 78 385
rect 76 384 77 385
rect 75 384 76 385
rect 74 384 75 385
rect 73 384 74 385
rect 72 384 73 385
rect 71 384 72 385
rect 70 384 71 385
rect 69 384 70 385
rect 68 384 69 385
rect 67 384 68 385
rect 66 384 67 385
rect 65 384 66 385
rect 64 384 65 385
rect 63 384 64 385
rect 62 384 63 385
rect 61 384 62 385
rect 60 384 61 385
rect 59 384 60 385
rect 58 384 59 385
rect 57 384 58 385
rect 56 384 57 385
rect 55 384 56 385
rect 54 384 55 385
rect 53 384 54 385
rect 52 384 53 385
rect 51 384 52 385
rect 50 384 51 385
rect 49 384 50 385
rect 48 384 49 385
rect 47 384 48 385
rect 46 384 47 385
rect 45 384 46 385
rect 44 384 45 385
rect 43 384 44 385
rect 42 384 43 385
rect 41 384 42 385
rect 40 384 41 385
rect 39 384 40 385
rect 38 384 39 385
rect 37 384 38 385
rect 36 384 37 385
rect 35 384 36 385
rect 34 384 35 385
rect 33 384 34 385
rect 32 384 33 385
rect 31 384 32 385
rect 30 384 31 385
rect 29 384 30 385
rect 28 384 29 385
rect 27 384 28 385
rect 26 384 27 385
rect 25 384 26 385
rect 24 384 25 385
rect 23 384 24 385
rect 22 384 23 385
rect 21 384 22 385
rect 20 384 21 385
rect 19 384 20 385
rect 18 384 19 385
rect 17 384 18 385
rect 16 384 17 385
rect 15 384 16 385
rect 141 385 142 386
rect 140 385 141 386
rect 139 385 140 386
rect 138 385 139 386
rect 137 385 138 386
rect 136 385 137 386
rect 135 385 136 386
rect 134 385 135 386
rect 133 385 134 386
rect 132 385 133 386
rect 131 385 132 386
rect 130 385 131 386
rect 129 385 130 386
rect 128 385 129 386
rect 127 385 128 386
rect 126 385 127 386
rect 125 385 126 386
rect 79 385 80 386
rect 78 385 79 386
rect 77 385 78 386
rect 76 385 77 386
rect 75 385 76 386
rect 74 385 75 386
rect 73 385 74 386
rect 72 385 73 386
rect 71 385 72 386
rect 70 385 71 386
rect 69 385 70 386
rect 68 385 69 386
rect 67 385 68 386
rect 66 385 67 386
rect 65 385 66 386
rect 64 385 65 386
rect 63 385 64 386
rect 62 385 63 386
rect 61 385 62 386
rect 60 385 61 386
rect 59 385 60 386
rect 58 385 59 386
rect 57 385 58 386
rect 56 385 57 386
rect 55 385 56 386
rect 54 385 55 386
rect 53 385 54 386
rect 52 385 53 386
rect 51 385 52 386
rect 50 385 51 386
rect 49 385 50 386
rect 48 385 49 386
rect 47 385 48 386
rect 46 385 47 386
rect 45 385 46 386
rect 44 385 45 386
rect 43 385 44 386
rect 42 385 43 386
rect 41 385 42 386
rect 40 385 41 386
rect 39 385 40 386
rect 38 385 39 386
rect 37 385 38 386
rect 36 385 37 386
rect 35 385 36 386
rect 34 385 35 386
rect 33 385 34 386
rect 32 385 33 386
rect 31 385 32 386
rect 30 385 31 386
rect 29 385 30 386
rect 28 385 29 386
rect 27 385 28 386
rect 26 385 27 386
rect 25 385 26 386
rect 24 385 25 386
rect 23 385 24 386
rect 22 385 23 386
rect 21 385 22 386
rect 20 385 21 386
rect 19 385 20 386
rect 18 385 19 386
rect 17 385 18 386
rect 16 385 17 386
rect 15 385 16 386
rect 141 386 142 387
rect 140 386 141 387
rect 139 386 140 387
rect 138 386 139 387
rect 137 386 138 387
rect 136 386 137 387
rect 135 386 136 387
rect 134 386 135 387
rect 133 386 134 387
rect 132 386 133 387
rect 131 386 132 387
rect 130 386 131 387
rect 129 386 130 387
rect 128 386 129 387
rect 127 386 128 387
rect 126 386 127 387
rect 125 386 126 387
rect 78 386 79 387
rect 77 386 78 387
rect 76 386 77 387
rect 75 386 76 387
rect 74 386 75 387
rect 73 386 74 387
rect 72 386 73 387
rect 71 386 72 387
rect 70 386 71 387
rect 69 386 70 387
rect 68 386 69 387
rect 67 386 68 387
rect 66 386 67 387
rect 65 386 66 387
rect 64 386 65 387
rect 63 386 64 387
rect 62 386 63 387
rect 61 386 62 387
rect 60 386 61 387
rect 59 386 60 387
rect 58 386 59 387
rect 57 386 58 387
rect 56 386 57 387
rect 55 386 56 387
rect 54 386 55 387
rect 53 386 54 387
rect 52 386 53 387
rect 51 386 52 387
rect 50 386 51 387
rect 49 386 50 387
rect 48 386 49 387
rect 47 386 48 387
rect 46 386 47 387
rect 45 386 46 387
rect 44 386 45 387
rect 43 386 44 387
rect 42 386 43 387
rect 41 386 42 387
rect 40 386 41 387
rect 39 386 40 387
rect 38 386 39 387
rect 37 386 38 387
rect 36 386 37 387
rect 35 386 36 387
rect 34 386 35 387
rect 33 386 34 387
rect 32 386 33 387
rect 31 386 32 387
rect 30 386 31 387
rect 29 386 30 387
rect 28 386 29 387
rect 27 386 28 387
rect 26 386 27 387
rect 25 386 26 387
rect 24 386 25 387
rect 23 386 24 387
rect 22 386 23 387
rect 21 386 22 387
rect 20 386 21 387
rect 19 386 20 387
rect 18 386 19 387
rect 17 386 18 387
rect 16 386 17 387
rect 15 386 16 387
rect 141 387 142 388
rect 140 387 141 388
rect 139 387 140 388
rect 138 387 139 388
rect 137 387 138 388
rect 136 387 137 388
rect 130 387 131 388
rect 129 387 130 388
rect 128 387 129 388
rect 127 387 128 388
rect 126 387 127 388
rect 125 387 126 388
rect 77 387 78 388
rect 76 387 77 388
rect 75 387 76 388
rect 74 387 75 388
rect 73 387 74 388
rect 72 387 73 388
rect 71 387 72 388
rect 70 387 71 388
rect 69 387 70 388
rect 68 387 69 388
rect 67 387 68 388
rect 66 387 67 388
rect 65 387 66 388
rect 64 387 65 388
rect 63 387 64 388
rect 62 387 63 388
rect 61 387 62 388
rect 60 387 61 388
rect 59 387 60 388
rect 58 387 59 388
rect 57 387 58 388
rect 56 387 57 388
rect 55 387 56 388
rect 54 387 55 388
rect 53 387 54 388
rect 52 387 53 388
rect 51 387 52 388
rect 50 387 51 388
rect 49 387 50 388
rect 48 387 49 388
rect 47 387 48 388
rect 46 387 47 388
rect 45 387 46 388
rect 44 387 45 388
rect 43 387 44 388
rect 42 387 43 388
rect 41 387 42 388
rect 40 387 41 388
rect 39 387 40 388
rect 38 387 39 388
rect 37 387 38 388
rect 36 387 37 388
rect 35 387 36 388
rect 34 387 35 388
rect 33 387 34 388
rect 32 387 33 388
rect 31 387 32 388
rect 30 387 31 388
rect 29 387 30 388
rect 28 387 29 388
rect 27 387 28 388
rect 26 387 27 388
rect 25 387 26 388
rect 24 387 25 388
rect 23 387 24 388
rect 22 387 23 388
rect 21 387 22 388
rect 20 387 21 388
rect 19 387 20 388
rect 18 387 19 388
rect 17 387 18 388
rect 16 387 17 388
rect 142 388 143 389
rect 141 388 142 389
rect 140 388 141 389
rect 139 388 140 389
rect 138 388 139 389
rect 128 388 129 389
rect 127 388 128 389
rect 126 388 127 389
rect 125 388 126 389
rect 124 388 125 389
rect 77 388 78 389
rect 76 388 77 389
rect 75 388 76 389
rect 74 388 75 389
rect 73 388 74 389
rect 72 388 73 389
rect 71 388 72 389
rect 70 388 71 389
rect 69 388 70 389
rect 68 388 69 389
rect 67 388 68 389
rect 66 388 67 389
rect 65 388 66 389
rect 64 388 65 389
rect 63 388 64 389
rect 62 388 63 389
rect 61 388 62 389
rect 60 388 61 389
rect 59 388 60 389
rect 58 388 59 389
rect 57 388 58 389
rect 56 388 57 389
rect 55 388 56 389
rect 54 388 55 389
rect 53 388 54 389
rect 52 388 53 389
rect 51 388 52 389
rect 50 388 51 389
rect 49 388 50 389
rect 48 388 49 389
rect 47 388 48 389
rect 46 388 47 389
rect 45 388 46 389
rect 44 388 45 389
rect 43 388 44 389
rect 42 388 43 389
rect 41 388 42 389
rect 40 388 41 389
rect 39 388 40 389
rect 38 388 39 389
rect 37 388 38 389
rect 36 388 37 389
rect 35 388 36 389
rect 34 388 35 389
rect 33 388 34 389
rect 32 388 33 389
rect 31 388 32 389
rect 30 388 31 389
rect 29 388 30 389
rect 28 388 29 389
rect 27 388 28 389
rect 26 388 27 389
rect 25 388 26 389
rect 24 388 25 389
rect 23 388 24 389
rect 22 388 23 389
rect 21 388 22 389
rect 20 388 21 389
rect 19 388 20 389
rect 18 388 19 389
rect 17 388 18 389
rect 142 389 143 390
rect 141 389 142 390
rect 140 389 141 390
rect 139 389 140 390
rect 138 389 139 390
rect 128 389 129 390
rect 127 389 128 390
rect 126 389 127 390
rect 125 389 126 390
rect 124 389 125 390
rect 76 389 77 390
rect 75 389 76 390
rect 74 389 75 390
rect 73 389 74 390
rect 72 389 73 390
rect 71 389 72 390
rect 70 389 71 390
rect 69 389 70 390
rect 68 389 69 390
rect 67 389 68 390
rect 66 389 67 390
rect 65 389 66 390
rect 64 389 65 390
rect 63 389 64 390
rect 62 389 63 390
rect 61 389 62 390
rect 60 389 61 390
rect 59 389 60 390
rect 58 389 59 390
rect 57 389 58 390
rect 56 389 57 390
rect 55 389 56 390
rect 54 389 55 390
rect 53 389 54 390
rect 52 389 53 390
rect 51 389 52 390
rect 50 389 51 390
rect 49 389 50 390
rect 48 389 49 390
rect 47 389 48 390
rect 46 389 47 390
rect 45 389 46 390
rect 44 389 45 390
rect 43 389 44 390
rect 42 389 43 390
rect 41 389 42 390
rect 40 389 41 390
rect 39 389 40 390
rect 38 389 39 390
rect 37 389 38 390
rect 36 389 37 390
rect 35 389 36 390
rect 34 389 35 390
rect 33 389 34 390
rect 32 389 33 390
rect 31 389 32 390
rect 30 389 31 390
rect 29 389 30 390
rect 28 389 29 390
rect 27 389 28 390
rect 26 389 27 390
rect 25 389 26 390
rect 24 389 25 390
rect 23 389 24 390
rect 22 389 23 390
rect 21 389 22 390
rect 20 389 21 390
rect 19 389 20 390
rect 18 389 19 390
rect 17 389 18 390
rect 142 390 143 391
rect 141 390 142 391
rect 140 390 141 391
rect 139 390 140 391
rect 127 390 128 391
rect 126 390 127 391
rect 125 390 126 391
rect 124 390 125 391
rect 75 390 76 391
rect 74 390 75 391
rect 73 390 74 391
rect 72 390 73 391
rect 71 390 72 391
rect 70 390 71 391
rect 69 390 70 391
rect 68 390 69 391
rect 67 390 68 391
rect 66 390 67 391
rect 65 390 66 391
rect 64 390 65 391
rect 63 390 64 391
rect 62 390 63 391
rect 61 390 62 391
rect 60 390 61 391
rect 59 390 60 391
rect 58 390 59 391
rect 57 390 58 391
rect 56 390 57 391
rect 55 390 56 391
rect 54 390 55 391
rect 53 390 54 391
rect 52 390 53 391
rect 51 390 52 391
rect 50 390 51 391
rect 49 390 50 391
rect 48 390 49 391
rect 47 390 48 391
rect 46 390 47 391
rect 45 390 46 391
rect 44 390 45 391
rect 43 390 44 391
rect 42 390 43 391
rect 41 390 42 391
rect 40 390 41 391
rect 39 390 40 391
rect 38 390 39 391
rect 37 390 38 391
rect 36 390 37 391
rect 35 390 36 391
rect 34 390 35 391
rect 33 390 34 391
rect 32 390 33 391
rect 31 390 32 391
rect 30 390 31 391
rect 29 390 30 391
rect 28 390 29 391
rect 27 390 28 391
rect 26 390 27 391
rect 25 390 26 391
rect 24 390 25 391
rect 23 390 24 391
rect 22 390 23 391
rect 21 390 22 391
rect 20 390 21 391
rect 19 390 20 391
rect 18 390 19 391
rect 142 391 143 392
rect 141 391 142 392
rect 140 391 141 392
rect 139 391 140 392
rect 127 391 128 392
rect 126 391 127 392
rect 125 391 126 392
rect 124 391 125 392
rect 74 391 75 392
rect 73 391 74 392
rect 72 391 73 392
rect 71 391 72 392
rect 70 391 71 392
rect 69 391 70 392
rect 68 391 69 392
rect 67 391 68 392
rect 66 391 67 392
rect 65 391 66 392
rect 64 391 65 392
rect 63 391 64 392
rect 62 391 63 392
rect 61 391 62 392
rect 60 391 61 392
rect 59 391 60 392
rect 58 391 59 392
rect 57 391 58 392
rect 56 391 57 392
rect 55 391 56 392
rect 54 391 55 392
rect 53 391 54 392
rect 52 391 53 392
rect 51 391 52 392
rect 50 391 51 392
rect 49 391 50 392
rect 48 391 49 392
rect 47 391 48 392
rect 46 391 47 392
rect 45 391 46 392
rect 44 391 45 392
rect 43 391 44 392
rect 42 391 43 392
rect 41 391 42 392
rect 40 391 41 392
rect 39 391 40 392
rect 38 391 39 392
rect 37 391 38 392
rect 36 391 37 392
rect 35 391 36 392
rect 34 391 35 392
rect 33 391 34 392
rect 32 391 33 392
rect 31 391 32 392
rect 30 391 31 392
rect 29 391 30 392
rect 28 391 29 392
rect 27 391 28 392
rect 26 391 27 392
rect 25 391 26 392
rect 24 391 25 392
rect 23 391 24 392
rect 22 391 23 392
rect 21 391 22 392
rect 20 391 21 392
rect 19 391 20 392
rect 142 392 143 393
rect 141 392 142 393
rect 140 392 141 393
rect 139 392 140 393
rect 127 392 128 393
rect 126 392 127 393
rect 125 392 126 393
rect 124 392 125 393
rect 73 392 74 393
rect 72 392 73 393
rect 71 392 72 393
rect 70 392 71 393
rect 69 392 70 393
rect 68 392 69 393
rect 67 392 68 393
rect 66 392 67 393
rect 65 392 66 393
rect 64 392 65 393
rect 63 392 64 393
rect 62 392 63 393
rect 61 392 62 393
rect 60 392 61 393
rect 59 392 60 393
rect 58 392 59 393
rect 57 392 58 393
rect 56 392 57 393
rect 55 392 56 393
rect 54 392 55 393
rect 53 392 54 393
rect 52 392 53 393
rect 51 392 52 393
rect 50 392 51 393
rect 49 392 50 393
rect 48 392 49 393
rect 47 392 48 393
rect 46 392 47 393
rect 45 392 46 393
rect 44 392 45 393
rect 43 392 44 393
rect 42 392 43 393
rect 41 392 42 393
rect 40 392 41 393
rect 39 392 40 393
rect 38 392 39 393
rect 37 392 38 393
rect 36 392 37 393
rect 35 392 36 393
rect 34 392 35 393
rect 33 392 34 393
rect 32 392 33 393
rect 31 392 32 393
rect 30 392 31 393
rect 29 392 30 393
rect 28 392 29 393
rect 27 392 28 393
rect 26 392 27 393
rect 25 392 26 393
rect 24 392 25 393
rect 23 392 24 393
rect 22 392 23 393
rect 21 392 22 393
rect 20 392 21 393
rect 142 393 143 394
rect 141 393 142 394
rect 140 393 141 394
rect 139 393 140 394
rect 138 393 139 394
rect 128 393 129 394
rect 127 393 128 394
rect 126 393 127 394
rect 125 393 126 394
rect 124 393 125 394
rect 72 393 73 394
rect 71 393 72 394
rect 70 393 71 394
rect 69 393 70 394
rect 68 393 69 394
rect 67 393 68 394
rect 66 393 67 394
rect 65 393 66 394
rect 64 393 65 394
rect 63 393 64 394
rect 62 393 63 394
rect 61 393 62 394
rect 60 393 61 394
rect 59 393 60 394
rect 58 393 59 394
rect 57 393 58 394
rect 56 393 57 394
rect 55 393 56 394
rect 54 393 55 394
rect 53 393 54 394
rect 52 393 53 394
rect 51 393 52 394
rect 50 393 51 394
rect 49 393 50 394
rect 48 393 49 394
rect 47 393 48 394
rect 46 393 47 394
rect 45 393 46 394
rect 44 393 45 394
rect 43 393 44 394
rect 42 393 43 394
rect 41 393 42 394
rect 40 393 41 394
rect 39 393 40 394
rect 38 393 39 394
rect 37 393 38 394
rect 36 393 37 394
rect 35 393 36 394
rect 34 393 35 394
rect 33 393 34 394
rect 32 393 33 394
rect 31 393 32 394
rect 30 393 31 394
rect 29 393 30 394
rect 28 393 29 394
rect 27 393 28 394
rect 26 393 27 394
rect 25 393 26 394
rect 24 393 25 394
rect 23 393 24 394
rect 22 393 23 394
rect 21 393 22 394
rect 142 394 143 395
rect 141 394 142 395
rect 140 394 141 395
rect 139 394 140 395
rect 138 394 139 395
rect 137 394 138 395
rect 129 394 130 395
rect 128 394 129 395
rect 127 394 128 395
rect 126 394 127 395
rect 125 394 126 395
rect 124 394 125 395
rect 70 394 71 395
rect 69 394 70 395
rect 68 394 69 395
rect 67 394 68 395
rect 66 394 67 395
rect 65 394 66 395
rect 64 394 65 395
rect 63 394 64 395
rect 62 394 63 395
rect 61 394 62 395
rect 60 394 61 395
rect 59 394 60 395
rect 58 394 59 395
rect 57 394 58 395
rect 56 394 57 395
rect 55 394 56 395
rect 54 394 55 395
rect 53 394 54 395
rect 52 394 53 395
rect 51 394 52 395
rect 50 394 51 395
rect 49 394 50 395
rect 48 394 49 395
rect 47 394 48 395
rect 46 394 47 395
rect 45 394 46 395
rect 44 394 45 395
rect 43 394 44 395
rect 42 394 43 395
rect 41 394 42 395
rect 40 394 41 395
rect 39 394 40 395
rect 38 394 39 395
rect 37 394 38 395
rect 36 394 37 395
rect 35 394 36 395
rect 34 394 35 395
rect 33 394 34 395
rect 32 394 33 395
rect 31 394 32 395
rect 30 394 31 395
rect 29 394 30 395
rect 28 394 29 395
rect 27 394 28 395
rect 26 394 27 395
rect 25 394 26 395
rect 24 394 25 395
rect 23 394 24 395
rect 141 395 142 396
rect 140 395 141 396
rect 139 395 140 396
rect 138 395 139 396
rect 137 395 138 396
rect 136 395 137 396
rect 135 395 136 396
rect 131 395 132 396
rect 130 395 131 396
rect 129 395 130 396
rect 128 395 129 396
rect 127 395 128 396
rect 126 395 127 396
rect 125 395 126 396
rect 68 395 69 396
rect 67 395 68 396
rect 66 395 67 396
rect 65 395 66 396
rect 64 395 65 396
rect 63 395 64 396
rect 62 395 63 396
rect 61 395 62 396
rect 60 395 61 396
rect 59 395 60 396
rect 58 395 59 396
rect 57 395 58 396
rect 56 395 57 396
rect 55 395 56 396
rect 54 395 55 396
rect 53 395 54 396
rect 52 395 53 396
rect 51 395 52 396
rect 50 395 51 396
rect 49 395 50 396
rect 48 395 49 396
rect 47 395 48 396
rect 46 395 47 396
rect 45 395 46 396
rect 44 395 45 396
rect 43 395 44 396
rect 42 395 43 396
rect 41 395 42 396
rect 40 395 41 396
rect 39 395 40 396
rect 38 395 39 396
rect 37 395 38 396
rect 36 395 37 396
rect 35 395 36 396
rect 34 395 35 396
rect 33 395 34 396
rect 32 395 33 396
rect 31 395 32 396
rect 30 395 31 396
rect 29 395 30 396
rect 28 395 29 396
rect 27 395 28 396
rect 26 395 27 396
rect 25 395 26 396
rect 141 396 142 397
rect 140 396 141 397
rect 139 396 140 397
rect 138 396 139 397
rect 137 396 138 397
rect 136 396 137 397
rect 135 396 136 397
rect 134 396 135 397
rect 133 396 134 397
rect 132 396 133 397
rect 131 396 132 397
rect 130 396 131 397
rect 129 396 130 397
rect 128 396 129 397
rect 127 396 128 397
rect 126 396 127 397
rect 125 396 126 397
rect 66 396 67 397
rect 65 396 66 397
rect 64 396 65 397
rect 63 396 64 397
rect 62 396 63 397
rect 61 396 62 397
rect 60 396 61 397
rect 59 396 60 397
rect 58 396 59 397
rect 57 396 58 397
rect 56 396 57 397
rect 55 396 56 397
rect 54 396 55 397
rect 53 396 54 397
rect 52 396 53 397
rect 51 396 52 397
rect 50 396 51 397
rect 49 396 50 397
rect 48 396 49 397
rect 47 396 48 397
rect 46 396 47 397
rect 45 396 46 397
rect 44 396 45 397
rect 43 396 44 397
rect 42 396 43 397
rect 41 396 42 397
rect 40 396 41 397
rect 39 396 40 397
rect 38 396 39 397
rect 37 396 38 397
rect 36 396 37 397
rect 35 396 36 397
rect 34 396 35 397
rect 33 396 34 397
rect 32 396 33 397
rect 31 396 32 397
rect 30 396 31 397
rect 29 396 30 397
rect 28 396 29 397
rect 27 396 28 397
rect 140 397 141 398
rect 139 397 140 398
rect 138 397 139 398
rect 137 397 138 398
rect 136 397 137 398
rect 135 397 136 398
rect 134 397 135 398
rect 133 397 134 398
rect 132 397 133 398
rect 131 397 132 398
rect 130 397 131 398
rect 129 397 130 398
rect 128 397 129 398
rect 127 397 128 398
rect 126 397 127 398
rect 64 397 65 398
rect 63 397 64 398
rect 62 397 63 398
rect 61 397 62 398
rect 60 397 61 398
rect 59 397 60 398
rect 58 397 59 398
rect 57 397 58 398
rect 56 397 57 398
rect 55 397 56 398
rect 54 397 55 398
rect 53 397 54 398
rect 52 397 53 398
rect 51 397 52 398
rect 50 397 51 398
rect 49 397 50 398
rect 48 397 49 398
rect 47 397 48 398
rect 46 397 47 398
rect 45 397 46 398
rect 44 397 45 398
rect 43 397 44 398
rect 42 397 43 398
rect 41 397 42 398
rect 40 397 41 398
rect 39 397 40 398
rect 38 397 39 398
rect 37 397 38 398
rect 36 397 37 398
rect 35 397 36 398
rect 34 397 35 398
rect 33 397 34 398
rect 32 397 33 398
rect 31 397 32 398
rect 30 397 31 398
rect 29 397 30 398
rect 139 398 140 399
rect 138 398 139 399
rect 137 398 138 399
rect 136 398 137 399
rect 135 398 136 399
rect 134 398 135 399
rect 133 398 134 399
rect 132 398 133 399
rect 131 398 132 399
rect 130 398 131 399
rect 129 398 130 399
rect 128 398 129 399
rect 127 398 128 399
rect 126 398 127 399
rect 60 398 61 399
rect 59 398 60 399
rect 58 398 59 399
rect 57 398 58 399
rect 56 398 57 399
rect 55 398 56 399
rect 54 398 55 399
rect 53 398 54 399
rect 52 398 53 399
rect 51 398 52 399
rect 50 398 51 399
rect 49 398 50 399
rect 48 398 49 399
rect 47 398 48 399
rect 46 398 47 399
rect 45 398 46 399
rect 44 398 45 399
rect 43 398 44 399
rect 42 398 43 399
rect 41 398 42 399
rect 40 398 41 399
rect 39 398 40 399
rect 38 398 39 399
rect 37 398 38 399
rect 36 398 37 399
rect 35 398 36 399
rect 34 398 35 399
rect 33 398 34 399
rect 138 399 139 400
rect 137 399 138 400
rect 136 399 137 400
rect 135 399 136 400
rect 134 399 135 400
rect 133 399 134 400
rect 132 399 133 400
rect 131 399 132 400
rect 130 399 131 400
rect 129 399 130 400
rect 128 399 129 400
rect 53 399 54 400
rect 52 399 53 400
rect 51 399 52 400
rect 50 399 51 400
rect 49 399 50 400
rect 48 399 49 400
rect 47 399 48 400
rect 46 399 47 400
rect 45 399 46 400
rect 44 399 45 400
rect 43 399 44 400
rect 42 399 43 400
rect 41 399 42 400
rect 40 399 41 400
rect 136 400 137 401
rect 135 400 136 401
rect 134 400 135 401
rect 133 400 134 401
rect 132 400 133 401
rect 131 400 132 401
rect 130 400 131 401
rect 129 400 130 401
rect 136 404 137 405
rect 135 404 136 405
rect 134 404 135 405
rect 133 404 134 405
rect 132 404 133 405
rect 131 404 132 405
rect 130 404 131 405
rect 138 405 139 406
rect 137 405 138 406
rect 136 405 137 406
rect 135 405 136 406
rect 134 405 135 406
rect 133 405 134 406
rect 132 405 133 406
rect 131 405 132 406
rect 130 405 131 406
rect 129 405 130 406
rect 128 405 129 406
rect 139 406 140 407
rect 138 406 139 407
rect 137 406 138 407
rect 136 406 137 407
rect 135 406 136 407
rect 134 406 135 407
rect 133 406 134 407
rect 132 406 133 407
rect 131 406 132 407
rect 130 406 131 407
rect 129 406 130 407
rect 128 406 129 407
rect 127 406 128 407
rect 140 407 141 408
rect 139 407 140 408
rect 138 407 139 408
rect 137 407 138 408
rect 136 407 137 408
rect 135 407 136 408
rect 134 407 135 408
rect 133 407 134 408
rect 132 407 133 408
rect 131 407 132 408
rect 130 407 131 408
rect 129 407 130 408
rect 128 407 129 408
rect 127 407 128 408
rect 126 407 127 408
rect 80 407 81 408
rect 79 407 80 408
rect 78 407 79 408
rect 77 407 78 408
rect 76 407 77 408
rect 75 407 76 408
rect 74 407 75 408
rect 73 407 74 408
rect 72 407 73 408
rect 71 407 72 408
rect 70 407 71 408
rect 141 408 142 409
rect 140 408 141 409
rect 139 408 140 409
rect 138 408 139 409
rect 137 408 138 409
rect 136 408 137 409
rect 135 408 136 409
rect 134 408 135 409
rect 133 408 134 409
rect 132 408 133 409
rect 131 408 132 409
rect 130 408 131 409
rect 129 408 130 409
rect 128 408 129 409
rect 127 408 128 409
rect 126 408 127 409
rect 125 408 126 409
rect 80 408 81 409
rect 79 408 80 409
rect 78 408 79 409
rect 77 408 78 409
rect 76 408 77 409
rect 75 408 76 409
rect 74 408 75 409
rect 73 408 74 409
rect 72 408 73 409
rect 71 408 72 409
rect 70 408 71 409
rect 69 408 70 409
rect 68 408 69 409
rect 67 408 68 409
rect 66 408 67 409
rect 141 409 142 410
rect 140 409 141 410
rect 139 409 140 410
rect 138 409 139 410
rect 137 409 138 410
rect 136 409 137 410
rect 135 409 136 410
rect 134 409 135 410
rect 133 409 134 410
rect 132 409 133 410
rect 131 409 132 410
rect 130 409 131 410
rect 129 409 130 410
rect 128 409 129 410
rect 127 409 128 410
rect 126 409 127 410
rect 125 409 126 410
rect 80 409 81 410
rect 79 409 80 410
rect 78 409 79 410
rect 77 409 78 410
rect 76 409 77 410
rect 75 409 76 410
rect 74 409 75 410
rect 73 409 74 410
rect 72 409 73 410
rect 71 409 72 410
rect 70 409 71 410
rect 69 409 70 410
rect 68 409 69 410
rect 67 409 68 410
rect 66 409 67 410
rect 65 409 66 410
rect 64 409 65 410
rect 63 409 64 410
rect 142 410 143 411
rect 141 410 142 411
rect 140 410 141 411
rect 139 410 140 411
rect 138 410 139 411
rect 137 410 138 411
rect 129 410 130 411
rect 128 410 129 411
rect 127 410 128 411
rect 126 410 127 411
rect 125 410 126 411
rect 124 410 125 411
rect 80 410 81 411
rect 79 410 80 411
rect 78 410 79 411
rect 77 410 78 411
rect 76 410 77 411
rect 75 410 76 411
rect 74 410 75 411
rect 73 410 74 411
rect 72 410 73 411
rect 71 410 72 411
rect 70 410 71 411
rect 69 410 70 411
rect 68 410 69 411
rect 67 410 68 411
rect 66 410 67 411
rect 65 410 66 411
rect 64 410 65 411
rect 63 410 64 411
rect 62 410 63 411
rect 33 410 34 411
rect 32 410 33 411
rect 31 410 32 411
rect 30 410 31 411
rect 29 410 30 411
rect 28 410 29 411
rect 27 410 28 411
rect 26 410 27 411
rect 25 410 26 411
rect 24 410 25 411
rect 23 410 24 411
rect 22 410 23 411
rect 21 410 22 411
rect 20 410 21 411
rect 19 410 20 411
rect 18 410 19 411
rect 142 411 143 412
rect 141 411 142 412
rect 140 411 141 412
rect 139 411 140 412
rect 138 411 139 412
rect 128 411 129 412
rect 127 411 128 412
rect 126 411 127 412
rect 125 411 126 412
rect 124 411 125 412
rect 80 411 81 412
rect 79 411 80 412
rect 78 411 79 412
rect 77 411 78 412
rect 76 411 77 412
rect 75 411 76 412
rect 74 411 75 412
rect 73 411 74 412
rect 72 411 73 412
rect 71 411 72 412
rect 70 411 71 412
rect 69 411 70 412
rect 68 411 69 412
rect 67 411 68 412
rect 66 411 67 412
rect 65 411 66 412
rect 64 411 65 412
rect 63 411 64 412
rect 62 411 63 412
rect 61 411 62 412
rect 60 411 61 412
rect 32 411 33 412
rect 31 411 32 412
rect 30 411 31 412
rect 29 411 30 412
rect 28 411 29 412
rect 27 411 28 412
rect 26 411 27 412
rect 25 411 26 412
rect 24 411 25 412
rect 23 411 24 412
rect 22 411 23 412
rect 21 411 22 412
rect 20 411 21 412
rect 19 411 20 412
rect 18 411 19 412
rect 17 411 18 412
rect 142 412 143 413
rect 141 412 142 413
rect 140 412 141 413
rect 139 412 140 413
rect 138 412 139 413
rect 128 412 129 413
rect 127 412 128 413
rect 126 412 127 413
rect 125 412 126 413
rect 124 412 125 413
rect 80 412 81 413
rect 79 412 80 413
rect 78 412 79 413
rect 77 412 78 413
rect 76 412 77 413
rect 75 412 76 413
rect 74 412 75 413
rect 73 412 74 413
rect 72 412 73 413
rect 71 412 72 413
rect 70 412 71 413
rect 69 412 70 413
rect 68 412 69 413
rect 67 412 68 413
rect 66 412 67 413
rect 65 412 66 413
rect 64 412 65 413
rect 63 412 64 413
rect 62 412 63 413
rect 61 412 62 413
rect 60 412 61 413
rect 59 412 60 413
rect 32 412 33 413
rect 31 412 32 413
rect 30 412 31 413
rect 29 412 30 413
rect 28 412 29 413
rect 27 412 28 413
rect 26 412 27 413
rect 25 412 26 413
rect 24 412 25 413
rect 23 412 24 413
rect 22 412 23 413
rect 21 412 22 413
rect 20 412 21 413
rect 19 412 20 413
rect 18 412 19 413
rect 17 412 18 413
rect 142 413 143 414
rect 141 413 142 414
rect 140 413 141 414
rect 139 413 140 414
rect 127 413 128 414
rect 126 413 127 414
rect 125 413 126 414
rect 124 413 125 414
rect 80 413 81 414
rect 79 413 80 414
rect 78 413 79 414
rect 77 413 78 414
rect 76 413 77 414
rect 75 413 76 414
rect 74 413 75 414
rect 73 413 74 414
rect 72 413 73 414
rect 71 413 72 414
rect 70 413 71 414
rect 69 413 70 414
rect 68 413 69 414
rect 67 413 68 414
rect 66 413 67 414
rect 65 413 66 414
rect 64 413 65 414
rect 63 413 64 414
rect 62 413 63 414
rect 61 413 62 414
rect 60 413 61 414
rect 59 413 60 414
rect 58 413 59 414
rect 57 413 58 414
rect 31 413 32 414
rect 30 413 31 414
rect 29 413 30 414
rect 28 413 29 414
rect 27 413 28 414
rect 26 413 27 414
rect 25 413 26 414
rect 24 413 25 414
rect 23 413 24 414
rect 22 413 23 414
rect 21 413 22 414
rect 20 413 21 414
rect 19 413 20 414
rect 18 413 19 414
rect 17 413 18 414
rect 142 414 143 415
rect 141 414 142 415
rect 140 414 141 415
rect 139 414 140 415
rect 127 414 128 415
rect 126 414 127 415
rect 125 414 126 415
rect 124 414 125 415
rect 80 414 81 415
rect 79 414 80 415
rect 78 414 79 415
rect 77 414 78 415
rect 76 414 77 415
rect 75 414 76 415
rect 74 414 75 415
rect 73 414 74 415
rect 72 414 73 415
rect 71 414 72 415
rect 70 414 71 415
rect 69 414 70 415
rect 68 414 69 415
rect 67 414 68 415
rect 66 414 67 415
rect 65 414 66 415
rect 64 414 65 415
rect 63 414 64 415
rect 62 414 63 415
rect 61 414 62 415
rect 60 414 61 415
rect 59 414 60 415
rect 58 414 59 415
rect 57 414 58 415
rect 56 414 57 415
rect 31 414 32 415
rect 30 414 31 415
rect 29 414 30 415
rect 28 414 29 415
rect 27 414 28 415
rect 26 414 27 415
rect 25 414 26 415
rect 24 414 25 415
rect 23 414 24 415
rect 22 414 23 415
rect 21 414 22 415
rect 20 414 21 415
rect 19 414 20 415
rect 18 414 19 415
rect 17 414 18 415
rect 16 414 17 415
rect 142 415 143 416
rect 141 415 142 416
rect 140 415 141 416
rect 139 415 140 416
rect 138 415 139 416
rect 128 415 129 416
rect 127 415 128 416
rect 126 415 127 416
rect 125 415 126 416
rect 124 415 125 416
rect 80 415 81 416
rect 79 415 80 416
rect 78 415 79 416
rect 77 415 78 416
rect 76 415 77 416
rect 75 415 76 416
rect 74 415 75 416
rect 73 415 74 416
rect 72 415 73 416
rect 71 415 72 416
rect 70 415 71 416
rect 69 415 70 416
rect 68 415 69 416
rect 67 415 68 416
rect 66 415 67 416
rect 65 415 66 416
rect 64 415 65 416
rect 63 415 64 416
rect 62 415 63 416
rect 61 415 62 416
rect 60 415 61 416
rect 59 415 60 416
rect 58 415 59 416
rect 57 415 58 416
rect 56 415 57 416
rect 55 415 56 416
rect 30 415 31 416
rect 29 415 30 416
rect 28 415 29 416
rect 27 415 28 416
rect 26 415 27 416
rect 25 415 26 416
rect 24 415 25 416
rect 23 415 24 416
rect 22 415 23 416
rect 21 415 22 416
rect 20 415 21 416
rect 19 415 20 416
rect 18 415 19 416
rect 17 415 18 416
rect 16 415 17 416
rect 142 416 143 417
rect 141 416 142 417
rect 140 416 141 417
rect 139 416 140 417
rect 138 416 139 417
rect 128 416 129 417
rect 127 416 128 417
rect 126 416 127 417
rect 125 416 126 417
rect 124 416 125 417
rect 80 416 81 417
rect 79 416 80 417
rect 78 416 79 417
rect 77 416 78 417
rect 76 416 77 417
rect 75 416 76 417
rect 74 416 75 417
rect 73 416 74 417
rect 72 416 73 417
rect 71 416 72 417
rect 70 416 71 417
rect 69 416 70 417
rect 68 416 69 417
rect 67 416 68 417
rect 66 416 67 417
rect 65 416 66 417
rect 64 416 65 417
rect 63 416 64 417
rect 62 416 63 417
rect 61 416 62 417
rect 60 416 61 417
rect 59 416 60 417
rect 58 416 59 417
rect 57 416 58 417
rect 56 416 57 417
rect 55 416 56 417
rect 54 416 55 417
rect 30 416 31 417
rect 29 416 30 417
rect 28 416 29 417
rect 27 416 28 417
rect 26 416 27 417
rect 25 416 26 417
rect 24 416 25 417
rect 23 416 24 417
rect 22 416 23 417
rect 21 416 22 417
rect 20 416 21 417
rect 19 416 20 417
rect 18 416 19 417
rect 17 416 18 417
rect 16 416 17 417
rect 15 416 16 417
rect 142 417 143 418
rect 141 417 142 418
rect 140 417 141 418
rect 139 417 140 418
rect 138 417 139 418
rect 137 417 138 418
rect 129 417 130 418
rect 128 417 129 418
rect 127 417 128 418
rect 126 417 127 418
rect 125 417 126 418
rect 124 417 125 418
rect 80 417 81 418
rect 79 417 80 418
rect 78 417 79 418
rect 77 417 78 418
rect 76 417 77 418
rect 75 417 76 418
rect 74 417 75 418
rect 73 417 74 418
rect 72 417 73 418
rect 71 417 72 418
rect 70 417 71 418
rect 69 417 70 418
rect 68 417 69 418
rect 67 417 68 418
rect 66 417 67 418
rect 65 417 66 418
rect 64 417 65 418
rect 63 417 64 418
rect 62 417 63 418
rect 61 417 62 418
rect 60 417 61 418
rect 59 417 60 418
rect 58 417 59 418
rect 57 417 58 418
rect 56 417 57 418
rect 55 417 56 418
rect 54 417 55 418
rect 29 417 30 418
rect 28 417 29 418
rect 27 417 28 418
rect 26 417 27 418
rect 25 417 26 418
rect 24 417 25 418
rect 23 417 24 418
rect 22 417 23 418
rect 21 417 22 418
rect 20 417 21 418
rect 19 417 20 418
rect 18 417 19 418
rect 17 417 18 418
rect 16 417 17 418
rect 15 417 16 418
rect 141 418 142 419
rect 140 418 141 419
rect 139 418 140 419
rect 138 418 139 419
rect 137 418 138 419
rect 136 418 137 419
rect 135 418 136 419
rect 134 418 135 419
rect 133 418 134 419
rect 132 418 133 419
rect 131 418 132 419
rect 130 418 131 419
rect 129 418 130 419
rect 128 418 129 419
rect 127 418 128 419
rect 126 418 127 419
rect 125 418 126 419
rect 80 418 81 419
rect 79 418 80 419
rect 78 418 79 419
rect 77 418 78 419
rect 76 418 77 419
rect 75 418 76 419
rect 74 418 75 419
rect 73 418 74 419
rect 72 418 73 419
rect 71 418 72 419
rect 70 418 71 419
rect 69 418 70 419
rect 68 418 69 419
rect 67 418 68 419
rect 66 418 67 419
rect 65 418 66 419
rect 64 418 65 419
rect 63 418 64 419
rect 62 418 63 419
rect 61 418 62 419
rect 60 418 61 419
rect 59 418 60 419
rect 58 418 59 419
rect 57 418 58 419
rect 56 418 57 419
rect 55 418 56 419
rect 54 418 55 419
rect 53 418 54 419
rect 29 418 30 419
rect 28 418 29 419
rect 27 418 28 419
rect 26 418 27 419
rect 25 418 26 419
rect 24 418 25 419
rect 23 418 24 419
rect 22 418 23 419
rect 21 418 22 419
rect 20 418 21 419
rect 19 418 20 419
rect 18 418 19 419
rect 17 418 18 419
rect 16 418 17 419
rect 15 418 16 419
rect 141 419 142 420
rect 140 419 141 420
rect 139 419 140 420
rect 138 419 139 420
rect 137 419 138 420
rect 136 419 137 420
rect 135 419 136 420
rect 134 419 135 420
rect 133 419 134 420
rect 132 419 133 420
rect 131 419 132 420
rect 130 419 131 420
rect 129 419 130 420
rect 128 419 129 420
rect 127 419 128 420
rect 126 419 127 420
rect 125 419 126 420
rect 80 419 81 420
rect 79 419 80 420
rect 78 419 79 420
rect 77 419 78 420
rect 76 419 77 420
rect 75 419 76 420
rect 74 419 75 420
rect 73 419 74 420
rect 72 419 73 420
rect 71 419 72 420
rect 70 419 71 420
rect 69 419 70 420
rect 68 419 69 420
rect 67 419 68 420
rect 66 419 67 420
rect 65 419 66 420
rect 64 419 65 420
rect 63 419 64 420
rect 62 419 63 420
rect 61 419 62 420
rect 60 419 61 420
rect 59 419 60 420
rect 58 419 59 420
rect 57 419 58 420
rect 56 419 57 420
rect 55 419 56 420
rect 54 419 55 420
rect 53 419 54 420
rect 52 419 53 420
rect 29 419 30 420
rect 28 419 29 420
rect 27 419 28 420
rect 26 419 27 420
rect 25 419 26 420
rect 24 419 25 420
rect 23 419 24 420
rect 22 419 23 420
rect 21 419 22 420
rect 20 419 21 420
rect 19 419 20 420
rect 18 419 19 420
rect 17 419 18 420
rect 16 419 17 420
rect 15 419 16 420
rect 14 419 15 420
rect 140 420 141 421
rect 139 420 140 421
rect 138 420 139 421
rect 137 420 138 421
rect 136 420 137 421
rect 135 420 136 421
rect 134 420 135 421
rect 133 420 134 421
rect 132 420 133 421
rect 131 420 132 421
rect 130 420 131 421
rect 129 420 130 421
rect 128 420 129 421
rect 127 420 128 421
rect 126 420 127 421
rect 80 420 81 421
rect 79 420 80 421
rect 78 420 79 421
rect 77 420 78 421
rect 76 420 77 421
rect 75 420 76 421
rect 74 420 75 421
rect 73 420 74 421
rect 72 420 73 421
rect 71 420 72 421
rect 70 420 71 421
rect 69 420 70 421
rect 68 420 69 421
rect 67 420 68 421
rect 66 420 67 421
rect 65 420 66 421
rect 64 420 65 421
rect 63 420 64 421
rect 62 420 63 421
rect 61 420 62 421
rect 60 420 61 421
rect 59 420 60 421
rect 58 420 59 421
rect 57 420 58 421
rect 56 420 57 421
rect 55 420 56 421
rect 54 420 55 421
rect 53 420 54 421
rect 52 420 53 421
rect 51 420 52 421
rect 29 420 30 421
rect 28 420 29 421
rect 27 420 28 421
rect 26 420 27 421
rect 25 420 26 421
rect 24 420 25 421
rect 23 420 24 421
rect 22 420 23 421
rect 21 420 22 421
rect 20 420 21 421
rect 19 420 20 421
rect 18 420 19 421
rect 17 420 18 421
rect 16 420 17 421
rect 15 420 16 421
rect 14 420 15 421
rect 139 421 140 422
rect 138 421 139 422
rect 137 421 138 422
rect 136 421 137 422
rect 135 421 136 422
rect 134 421 135 422
rect 133 421 134 422
rect 132 421 133 422
rect 131 421 132 422
rect 130 421 131 422
rect 129 421 130 422
rect 128 421 129 422
rect 127 421 128 422
rect 80 421 81 422
rect 79 421 80 422
rect 78 421 79 422
rect 77 421 78 422
rect 76 421 77 422
rect 75 421 76 422
rect 74 421 75 422
rect 73 421 74 422
rect 72 421 73 422
rect 71 421 72 422
rect 70 421 71 422
rect 69 421 70 422
rect 68 421 69 422
rect 67 421 68 422
rect 66 421 67 422
rect 65 421 66 422
rect 64 421 65 422
rect 63 421 64 422
rect 62 421 63 422
rect 61 421 62 422
rect 60 421 61 422
rect 59 421 60 422
rect 58 421 59 422
rect 57 421 58 422
rect 56 421 57 422
rect 55 421 56 422
rect 54 421 55 422
rect 53 421 54 422
rect 52 421 53 422
rect 51 421 52 422
rect 50 421 51 422
rect 28 421 29 422
rect 27 421 28 422
rect 26 421 27 422
rect 25 421 26 422
rect 24 421 25 422
rect 23 421 24 422
rect 22 421 23 422
rect 21 421 22 422
rect 20 421 21 422
rect 19 421 20 422
rect 18 421 19 422
rect 17 421 18 422
rect 16 421 17 422
rect 15 421 16 422
rect 14 421 15 422
rect 138 422 139 423
rect 137 422 138 423
rect 136 422 137 423
rect 135 422 136 423
rect 134 422 135 423
rect 133 422 134 423
rect 132 422 133 423
rect 131 422 132 423
rect 130 422 131 423
rect 129 422 130 423
rect 128 422 129 423
rect 80 422 81 423
rect 79 422 80 423
rect 78 422 79 423
rect 77 422 78 423
rect 76 422 77 423
rect 75 422 76 423
rect 74 422 75 423
rect 73 422 74 423
rect 72 422 73 423
rect 71 422 72 423
rect 70 422 71 423
rect 69 422 70 423
rect 68 422 69 423
rect 67 422 68 423
rect 66 422 67 423
rect 65 422 66 423
rect 64 422 65 423
rect 63 422 64 423
rect 62 422 63 423
rect 61 422 62 423
rect 60 422 61 423
rect 59 422 60 423
rect 58 422 59 423
rect 57 422 58 423
rect 56 422 57 423
rect 55 422 56 423
rect 54 422 55 423
rect 53 422 54 423
rect 52 422 53 423
rect 51 422 52 423
rect 50 422 51 423
rect 49 422 50 423
rect 28 422 29 423
rect 27 422 28 423
rect 26 422 27 423
rect 25 422 26 423
rect 24 422 25 423
rect 23 422 24 423
rect 22 422 23 423
rect 21 422 22 423
rect 20 422 21 423
rect 19 422 20 423
rect 18 422 19 423
rect 17 422 18 423
rect 16 422 17 423
rect 15 422 16 423
rect 14 422 15 423
rect 135 423 136 424
rect 134 423 135 424
rect 133 423 134 424
rect 132 423 133 424
rect 131 423 132 424
rect 130 423 131 424
rect 80 423 81 424
rect 79 423 80 424
rect 78 423 79 424
rect 77 423 78 424
rect 76 423 77 424
rect 75 423 76 424
rect 74 423 75 424
rect 73 423 74 424
rect 72 423 73 424
rect 71 423 72 424
rect 70 423 71 424
rect 69 423 70 424
rect 68 423 69 424
rect 67 423 68 424
rect 66 423 67 424
rect 65 423 66 424
rect 64 423 65 424
rect 63 423 64 424
rect 62 423 63 424
rect 61 423 62 424
rect 60 423 61 424
rect 59 423 60 424
rect 58 423 59 424
rect 57 423 58 424
rect 56 423 57 424
rect 55 423 56 424
rect 54 423 55 424
rect 53 423 54 424
rect 52 423 53 424
rect 51 423 52 424
rect 50 423 51 424
rect 49 423 50 424
rect 28 423 29 424
rect 27 423 28 424
rect 26 423 27 424
rect 25 423 26 424
rect 24 423 25 424
rect 23 423 24 424
rect 22 423 23 424
rect 21 423 22 424
rect 20 423 21 424
rect 19 423 20 424
rect 18 423 19 424
rect 17 423 18 424
rect 16 423 17 424
rect 15 423 16 424
rect 14 423 15 424
rect 80 424 81 425
rect 79 424 80 425
rect 78 424 79 425
rect 77 424 78 425
rect 76 424 77 425
rect 75 424 76 425
rect 74 424 75 425
rect 73 424 74 425
rect 72 424 73 425
rect 71 424 72 425
rect 70 424 71 425
rect 69 424 70 425
rect 68 424 69 425
rect 67 424 68 425
rect 66 424 67 425
rect 65 424 66 425
rect 64 424 65 425
rect 63 424 64 425
rect 62 424 63 425
rect 61 424 62 425
rect 60 424 61 425
rect 59 424 60 425
rect 58 424 59 425
rect 57 424 58 425
rect 56 424 57 425
rect 55 424 56 425
rect 54 424 55 425
rect 53 424 54 425
rect 52 424 53 425
rect 51 424 52 425
rect 50 424 51 425
rect 49 424 50 425
rect 48 424 49 425
rect 28 424 29 425
rect 27 424 28 425
rect 26 424 27 425
rect 25 424 26 425
rect 24 424 25 425
rect 23 424 24 425
rect 22 424 23 425
rect 21 424 22 425
rect 20 424 21 425
rect 19 424 20 425
rect 18 424 19 425
rect 17 424 18 425
rect 16 424 17 425
rect 15 424 16 425
rect 14 424 15 425
rect 80 425 81 426
rect 79 425 80 426
rect 78 425 79 426
rect 77 425 78 426
rect 76 425 77 426
rect 75 425 76 426
rect 74 425 75 426
rect 73 425 74 426
rect 72 425 73 426
rect 71 425 72 426
rect 70 425 71 426
rect 69 425 70 426
rect 68 425 69 426
rect 67 425 68 426
rect 66 425 67 426
rect 65 425 66 426
rect 64 425 65 426
rect 63 425 64 426
rect 62 425 63 426
rect 61 425 62 426
rect 60 425 61 426
rect 59 425 60 426
rect 58 425 59 426
rect 57 425 58 426
rect 56 425 57 426
rect 55 425 56 426
rect 54 425 55 426
rect 53 425 54 426
rect 52 425 53 426
rect 51 425 52 426
rect 50 425 51 426
rect 49 425 50 426
rect 48 425 49 426
rect 47 425 48 426
rect 28 425 29 426
rect 27 425 28 426
rect 26 425 27 426
rect 25 425 26 426
rect 24 425 25 426
rect 23 425 24 426
rect 22 425 23 426
rect 21 425 22 426
rect 20 425 21 426
rect 19 425 20 426
rect 18 425 19 426
rect 17 425 18 426
rect 16 425 17 426
rect 15 425 16 426
rect 14 425 15 426
rect 13 425 14 426
rect 80 426 81 427
rect 79 426 80 427
rect 78 426 79 427
rect 77 426 78 427
rect 76 426 77 427
rect 75 426 76 427
rect 74 426 75 427
rect 73 426 74 427
rect 72 426 73 427
rect 71 426 72 427
rect 70 426 71 427
rect 69 426 70 427
rect 68 426 69 427
rect 67 426 68 427
rect 66 426 67 427
rect 65 426 66 427
rect 64 426 65 427
rect 63 426 64 427
rect 62 426 63 427
rect 61 426 62 427
rect 60 426 61 427
rect 59 426 60 427
rect 58 426 59 427
rect 57 426 58 427
rect 56 426 57 427
rect 55 426 56 427
rect 54 426 55 427
rect 53 426 54 427
rect 52 426 53 427
rect 51 426 52 427
rect 50 426 51 427
rect 49 426 50 427
rect 48 426 49 427
rect 47 426 48 427
rect 46 426 47 427
rect 28 426 29 427
rect 27 426 28 427
rect 26 426 27 427
rect 25 426 26 427
rect 24 426 25 427
rect 23 426 24 427
rect 22 426 23 427
rect 21 426 22 427
rect 20 426 21 427
rect 19 426 20 427
rect 18 426 19 427
rect 17 426 18 427
rect 16 426 17 427
rect 15 426 16 427
rect 14 426 15 427
rect 13 426 14 427
rect 80 427 81 428
rect 79 427 80 428
rect 78 427 79 428
rect 77 427 78 428
rect 76 427 77 428
rect 75 427 76 428
rect 74 427 75 428
rect 73 427 74 428
rect 72 427 73 428
rect 71 427 72 428
rect 70 427 71 428
rect 69 427 70 428
rect 68 427 69 428
rect 67 427 68 428
rect 66 427 67 428
rect 65 427 66 428
rect 64 427 65 428
rect 63 427 64 428
rect 62 427 63 428
rect 61 427 62 428
rect 60 427 61 428
rect 59 427 60 428
rect 58 427 59 428
rect 57 427 58 428
rect 56 427 57 428
rect 55 427 56 428
rect 54 427 55 428
rect 53 427 54 428
rect 52 427 53 428
rect 51 427 52 428
rect 50 427 51 428
rect 49 427 50 428
rect 48 427 49 428
rect 47 427 48 428
rect 46 427 47 428
rect 45 427 46 428
rect 28 427 29 428
rect 27 427 28 428
rect 26 427 27 428
rect 25 427 26 428
rect 24 427 25 428
rect 23 427 24 428
rect 22 427 23 428
rect 21 427 22 428
rect 20 427 21 428
rect 19 427 20 428
rect 18 427 19 428
rect 17 427 18 428
rect 16 427 17 428
rect 15 427 16 428
rect 14 427 15 428
rect 13 427 14 428
rect 142 428 143 429
rect 141 428 142 429
rect 140 428 141 429
rect 139 428 140 429
rect 138 428 139 429
rect 137 428 138 429
rect 136 428 137 429
rect 135 428 136 429
rect 134 428 135 429
rect 133 428 134 429
rect 132 428 133 429
rect 131 428 132 429
rect 130 428 131 429
rect 129 428 130 429
rect 128 428 129 429
rect 127 428 128 429
rect 126 428 127 429
rect 125 428 126 429
rect 124 428 125 429
rect 123 428 124 429
rect 122 428 123 429
rect 121 428 122 429
rect 120 428 121 429
rect 119 428 120 429
rect 118 428 119 429
rect 117 428 118 429
rect 116 428 117 429
rect 115 428 116 429
rect 80 428 81 429
rect 79 428 80 429
rect 78 428 79 429
rect 77 428 78 429
rect 76 428 77 429
rect 75 428 76 429
rect 74 428 75 429
rect 73 428 74 429
rect 72 428 73 429
rect 71 428 72 429
rect 70 428 71 429
rect 69 428 70 429
rect 68 428 69 429
rect 67 428 68 429
rect 66 428 67 429
rect 65 428 66 429
rect 63 428 64 429
rect 62 428 63 429
rect 61 428 62 429
rect 60 428 61 429
rect 59 428 60 429
rect 58 428 59 429
rect 57 428 58 429
rect 56 428 57 429
rect 55 428 56 429
rect 54 428 55 429
rect 53 428 54 429
rect 52 428 53 429
rect 51 428 52 429
rect 50 428 51 429
rect 49 428 50 429
rect 48 428 49 429
rect 47 428 48 429
rect 46 428 47 429
rect 45 428 46 429
rect 28 428 29 429
rect 27 428 28 429
rect 26 428 27 429
rect 25 428 26 429
rect 24 428 25 429
rect 23 428 24 429
rect 22 428 23 429
rect 21 428 22 429
rect 20 428 21 429
rect 19 428 20 429
rect 18 428 19 429
rect 17 428 18 429
rect 16 428 17 429
rect 15 428 16 429
rect 14 428 15 429
rect 13 428 14 429
rect 142 429 143 430
rect 141 429 142 430
rect 140 429 141 430
rect 139 429 140 430
rect 138 429 139 430
rect 137 429 138 430
rect 136 429 137 430
rect 135 429 136 430
rect 134 429 135 430
rect 133 429 134 430
rect 132 429 133 430
rect 131 429 132 430
rect 130 429 131 430
rect 129 429 130 430
rect 128 429 129 430
rect 127 429 128 430
rect 126 429 127 430
rect 125 429 126 430
rect 124 429 125 430
rect 123 429 124 430
rect 122 429 123 430
rect 121 429 122 430
rect 120 429 121 430
rect 119 429 120 430
rect 118 429 119 430
rect 117 429 118 430
rect 116 429 117 430
rect 115 429 116 430
rect 80 429 81 430
rect 79 429 80 430
rect 78 429 79 430
rect 77 429 78 430
rect 76 429 77 430
rect 75 429 76 430
rect 74 429 75 430
rect 73 429 74 430
rect 72 429 73 430
rect 71 429 72 430
rect 70 429 71 430
rect 69 429 70 430
rect 68 429 69 430
rect 67 429 68 430
rect 66 429 67 430
rect 65 429 66 430
rect 62 429 63 430
rect 61 429 62 430
rect 60 429 61 430
rect 59 429 60 430
rect 58 429 59 430
rect 57 429 58 430
rect 56 429 57 430
rect 55 429 56 430
rect 54 429 55 430
rect 53 429 54 430
rect 52 429 53 430
rect 51 429 52 430
rect 50 429 51 430
rect 49 429 50 430
rect 48 429 49 430
rect 47 429 48 430
rect 46 429 47 430
rect 45 429 46 430
rect 44 429 45 430
rect 28 429 29 430
rect 27 429 28 430
rect 26 429 27 430
rect 25 429 26 430
rect 24 429 25 430
rect 23 429 24 430
rect 22 429 23 430
rect 21 429 22 430
rect 20 429 21 430
rect 19 429 20 430
rect 18 429 19 430
rect 17 429 18 430
rect 16 429 17 430
rect 15 429 16 430
rect 14 429 15 430
rect 13 429 14 430
rect 142 430 143 431
rect 141 430 142 431
rect 140 430 141 431
rect 139 430 140 431
rect 138 430 139 431
rect 137 430 138 431
rect 136 430 137 431
rect 135 430 136 431
rect 134 430 135 431
rect 133 430 134 431
rect 132 430 133 431
rect 131 430 132 431
rect 130 430 131 431
rect 129 430 130 431
rect 128 430 129 431
rect 127 430 128 431
rect 126 430 127 431
rect 125 430 126 431
rect 124 430 125 431
rect 123 430 124 431
rect 122 430 123 431
rect 121 430 122 431
rect 120 430 121 431
rect 119 430 120 431
rect 118 430 119 431
rect 117 430 118 431
rect 116 430 117 431
rect 115 430 116 431
rect 80 430 81 431
rect 79 430 80 431
rect 78 430 79 431
rect 77 430 78 431
rect 76 430 77 431
rect 75 430 76 431
rect 74 430 75 431
rect 73 430 74 431
rect 72 430 73 431
rect 71 430 72 431
rect 70 430 71 431
rect 69 430 70 431
rect 68 430 69 431
rect 67 430 68 431
rect 66 430 67 431
rect 65 430 66 431
rect 61 430 62 431
rect 60 430 61 431
rect 59 430 60 431
rect 58 430 59 431
rect 57 430 58 431
rect 56 430 57 431
rect 55 430 56 431
rect 54 430 55 431
rect 53 430 54 431
rect 52 430 53 431
rect 51 430 52 431
rect 50 430 51 431
rect 49 430 50 431
rect 48 430 49 431
rect 47 430 48 431
rect 46 430 47 431
rect 45 430 46 431
rect 44 430 45 431
rect 43 430 44 431
rect 29 430 30 431
rect 28 430 29 431
rect 27 430 28 431
rect 26 430 27 431
rect 25 430 26 431
rect 24 430 25 431
rect 23 430 24 431
rect 22 430 23 431
rect 21 430 22 431
rect 20 430 21 431
rect 19 430 20 431
rect 18 430 19 431
rect 17 430 18 431
rect 16 430 17 431
rect 15 430 16 431
rect 14 430 15 431
rect 13 430 14 431
rect 142 431 143 432
rect 141 431 142 432
rect 140 431 141 432
rect 139 431 140 432
rect 138 431 139 432
rect 137 431 138 432
rect 136 431 137 432
rect 135 431 136 432
rect 134 431 135 432
rect 133 431 134 432
rect 132 431 133 432
rect 131 431 132 432
rect 130 431 131 432
rect 129 431 130 432
rect 128 431 129 432
rect 127 431 128 432
rect 126 431 127 432
rect 125 431 126 432
rect 124 431 125 432
rect 123 431 124 432
rect 122 431 123 432
rect 121 431 122 432
rect 120 431 121 432
rect 119 431 120 432
rect 118 431 119 432
rect 117 431 118 432
rect 116 431 117 432
rect 115 431 116 432
rect 80 431 81 432
rect 79 431 80 432
rect 78 431 79 432
rect 77 431 78 432
rect 76 431 77 432
rect 75 431 76 432
rect 74 431 75 432
rect 73 431 74 432
rect 72 431 73 432
rect 71 431 72 432
rect 70 431 71 432
rect 69 431 70 432
rect 68 431 69 432
rect 67 431 68 432
rect 66 431 67 432
rect 65 431 66 432
rect 60 431 61 432
rect 59 431 60 432
rect 58 431 59 432
rect 57 431 58 432
rect 56 431 57 432
rect 55 431 56 432
rect 54 431 55 432
rect 53 431 54 432
rect 52 431 53 432
rect 51 431 52 432
rect 50 431 51 432
rect 49 431 50 432
rect 48 431 49 432
rect 47 431 48 432
rect 46 431 47 432
rect 45 431 46 432
rect 44 431 45 432
rect 43 431 44 432
rect 42 431 43 432
rect 29 431 30 432
rect 28 431 29 432
rect 27 431 28 432
rect 26 431 27 432
rect 25 431 26 432
rect 24 431 25 432
rect 23 431 24 432
rect 22 431 23 432
rect 21 431 22 432
rect 20 431 21 432
rect 19 431 20 432
rect 18 431 19 432
rect 17 431 18 432
rect 16 431 17 432
rect 15 431 16 432
rect 14 431 15 432
rect 13 431 14 432
rect 142 432 143 433
rect 141 432 142 433
rect 140 432 141 433
rect 139 432 140 433
rect 138 432 139 433
rect 137 432 138 433
rect 136 432 137 433
rect 135 432 136 433
rect 134 432 135 433
rect 133 432 134 433
rect 132 432 133 433
rect 131 432 132 433
rect 130 432 131 433
rect 129 432 130 433
rect 128 432 129 433
rect 127 432 128 433
rect 126 432 127 433
rect 125 432 126 433
rect 124 432 125 433
rect 123 432 124 433
rect 122 432 123 433
rect 121 432 122 433
rect 120 432 121 433
rect 119 432 120 433
rect 118 432 119 433
rect 117 432 118 433
rect 116 432 117 433
rect 115 432 116 433
rect 80 432 81 433
rect 79 432 80 433
rect 78 432 79 433
rect 77 432 78 433
rect 76 432 77 433
rect 75 432 76 433
rect 74 432 75 433
rect 73 432 74 433
rect 72 432 73 433
rect 71 432 72 433
rect 70 432 71 433
rect 69 432 70 433
rect 68 432 69 433
rect 67 432 68 433
rect 66 432 67 433
rect 65 432 66 433
rect 59 432 60 433
rect 58 432 59 433
rect 57 432 58 433
rect 56 432 57 433
rect 55 432 56 433
rect 54 432 55 433
rect 53 432 54 433
rect 52 432 53 433
rect 51 432 52 433
rect 50 432 51 433
rect 49 432 50 433
rect 48 432 49 433
rect 47 432 48 433
rect 46 432 47 433
rect 45 432 46 433
rect 44 432 45 433
rect 43 432 44 433
rect 42 432 43 433
rect 41 432 42 433
rect 40 432 41 433
rect 30 432 31 433
rect 29 432 30 433
rect 28 432 29 433
rect 27 432 28 433
rect 26 432 27 433
rect 25 432 26 433
rect 24 432 25 433
rect 23 432 24 433
rect 22 432 23 433
rect 21 432 22 433
rect 20 432 21 433
rect 19 432 20 433
rect 18 432 19 433
rect 17 432 18 433
rect 16 432 17 433
rect 15 432 16 433
rect 14 432 15 433
rect 13 432 14 433
rect 142 433 143 434
rect 141 433 142 434
rect 140 433 141 434
rect 139 433 140 434
rect 138 433 139 434
rect 137 433 138 434
rect 136 433 137 434
rect 135 433 136 434
rect 134 433 135 434
rect 133 433 134 434
rect 132 433 133 434
rect 131 433 132 434
rect 130 433 131 434
rect 129 433 130 434
rect 128 433 129 434
rect 127 433 128 434
rect 126 433 127 434
rect 125 433 126 434
rect 124 433 125 434
rect 123 433 124 434
rect 122 433 123 434
rect 121 433 122 434
rect 120 433 121 434
rect 119 433 120 434
rect 118 433 119 434
rect 117 433 118 434
rect 116 433 117 434
rect 115 433 116 434
rect 80 433 81 434
rect 79 433 80 434
rect 78 433 79 434
rect 77 433 78 434
rect 76 433 77 434
rect 75 433 76 434
rect 74 433 75 434
rect 73 433 74 434
rect 72 433 73 434
rect 71 433 72 434
rect 70 433 71 434
rect 69 433 70 434
rect 68 433 69 434
rect 67 433 68 434
rect 66 433 67 434
rect 65 433 66 434
rect 58 433 59 434
rect 57 433 58 434
rect 56 433 57 434
rect 55 433 56 434
rect 54 433 55 434
rect 53 433 54 434
rect 52 433 53 434
rect 51 433 52 434
rect 50 433 51 434
rect 49 433 50 434
rect 48 433 49 434
rect 47 433 48 434
rect 46 433 47 434
rect 45 433 46 434
rect 44 433 45 434
rect 43 433 44 434
rect 42 433 43 434
rect 41 433 42 434
rect 40 433 41 434
rect 39 433 40 434
rect 38 433 39 434
rect 32 433 33 434
rect 31 433 32 434
rect 30 433 31 434
rect 29 433 30 434
rect 28 433 29 434
rect 27 433 28 434
rect 26 433 27 434
rect 25 433 26 434
rect 24 433 25 434
rect 23 433 24 434
rect 22 433 23 434
rect 21 433 22 434
rect 20 433 21 434
rect 19 433 20 434
rect 18 433 19 434
rect 17 433 18 434
rect 16 433 17 434
rect 15 433 16 434
rect 14 433 15 434
rect 13 433 14 434
rect 134 434 135 435
rect 133 434 134 435
rect 132 434 133 435
rect 80 434 81 435
rect 79 434 80 435
rect 78 434 79 435
rect 77 434 78 435
rect 76 434 77 435
rect 75 434 76 435
rect 74 434 75 435
rect 73 434 74 435
rect 72 434 73 435
rect 71 434 72 435
rect 70 434 71 435
rect 69 434 70 435
rect 68 434 69 435
rect 67 434 68 435
rect 66 434 67 435
rect 65 434 66 435
rect 58 434 59 435
rect 57 434 58 435
rect 56 434 57 435
rect 55 434 56 435
rect 54 434 55 435
rect 53 434 54 435
rect 52 434 53 435
rect 51 434 52 435
rect 50 434 51 435
rect 49 434 50 435
rect 48 434 49 435
rect 47 434 48 435
rect 46 434 47 435
rect 45 434 46 435
rect 44 434 45 435
rect 43 434 44 435
rect 42 434 43 435
rect 41 434 42 435
rect 40 434 41 435
rect 39 434 40 435
rect 38 434 39 435
rect 37 434 38 435
rect 36 434 37 435
rect 35 434 36 435
rect 34 434 35 435
rect 33 434 34 435
rect 32 434 33 435
rect 31 434 32 435
rect 30 434 31 435
rect 29 434 30 435
rect 28 434 29 435
rect 27 434 28 435
rect 26 434 27 435
rect 25 434 26 435
rect 24 434 25 435
rect 23 434 24 435
rect 22 434 23 435
rect 21 434 22 435
rect 20 434 21 435
rect 19 434 20 435
rect 18 434 19 435
rect 17 434 18 435
rect 16 434 17 435
rect 15 434 16 435
rect 14 434 15 435
rect 13 434 14 435
rect 135 435 136 436
rect 134 435 135 436
rect 133 435 134 436
rect 132 435 133 436
rect 131 435 132 436
rect 130 435 131 436
rect 80 435 81 436
rect 79 435 80 436
rect 78 435 79 436
rect 77 435 78 436
rect 76 435 77 436
rect 75 435 76 436
rect 74 435 75 436
rect 73 435 74 436
rect 72 435 73 436
rect 71 435 72 436
rect 70 435 71 436
rect 69 435 70 436
rect 68 435 69 436
rect 67 435 68 436
rect 66 435 67 436
rect 65 435 66 436
rect 57 435 58 436
rect 56 435 57 436
rect 55 435 56 436
rect 54 435 55 436
rect 53 435 54 436
rect 52 435 53 436
rect 51 435 52 436
rect 50 435 51 436
rect 49 435 50 436
rect 48 435 49 436
rect 47 435 48 436
rect 46 435 47 436
rect 45 435 46 436
rect 44 435 45 436
rect 43 435 44 436
rect 42 435 43 436
rect 41 435 42 436
rect 40 435 41 436
rect 39 435 40 436
rect 38 435 39 436
rect 37 435 38 436
rect 36 435 37 436
rect 35 435 36 436
rect 34 435 35 436
rect 33 435 34 436
rect 32 435 33 436
rect 31 435 32 436
rect 30 435 31 436
rect 29 435 30 436
rect 28 435 29 436
rect 27 435 28 436
rect 26 435 27 436
rect 25 435 26 436
rect 24 435 25 436
rect 23 435 24 436
rect 22 435 23 436
rect 21 435 22 436
rect 20 435 21 436
rect 19 435 20 436
rect 18 435 19 436
rect 17 435 18 436
rect 16 435 17 436
rect 15 435 16 436
rect 14 435 15 436
rect 13 435 14 436
rect 137 436 138 437
rect 136 436 137 437
rect 135 436 136 437
rect 134 436 135 437
rect 133 436 134 437
rect 132 436 133 437
rect 131 436 132 437
rect 130 436 131 437
rect 129 436 130 437
rect 80 436 81 437
rect 79 436 80 437
rect 78 436 79 437
rect 77 436 78 437
rect 76 436 77 437
rect 75 436 76 437
rect 74 436 75 437
rect 73 436 74 437
rect 72 436 73 437
rect 71 436 72 437
rect 70 436 71 437
rect 69 436 70 437
rect 68 436 69 437
rect 67 436 68 437
rect 66 436 67 437
rect 65 436 66 437
rect 56 436 57 437
rect 55 436 56 437
rect 54 436 55 437
rect 53 436 54 437
rect 52 436 53 437
rect 51 436 52 437
rect 50 436 51 437
rect 49 436 50 437
rect 48 436 49 437
rect 47 436 48 437
rect 46 436 47 437
rect 45 436 46 437
rect 44 436 45 437
rect 43 436 44 437
rect 42 436 43 437
rect 41 436 42 437
rect 40 436 41 437
rect 39 436 40 437
rect 38 436 39 437
rect 37 436 38 437
rect 36 436 37 437
rect 35 436 36 437
rect 34 436 35 437
rect 33 436 34 437
rect 32 436 33 437
rect 31 436 32 437
rect 30 436 31 437
rect 29 436 30 437
rect 28 436 29 437
rect 27 436 28 437
rect 26 436 27 437
rect 25 436 26 437
rect 24 436 25 437
rect 23 436 24 437
rect 22 436 23 437
rect 21 436 22 437
rect 20 436 21 437
rect 19 436 20 437
rect 18 436 19 437
rect 17 436 18 437
rect 16 436 17 437
rect 15 436 16 437
rect 14 436 15 437
rect 13 436 14 437
rect 138 437 139 438
rect 137 437 138 438
rect 136 437 137 438
rect 135 437 136 438
rect 134 437 135 438
rect 133 437 134 438
rect 132 437 133 438
rect 131 437 132 438
rect 130 437 131 438
rect 129 437 130 438
rect 128 437 129 438
rect 127 437 128 438
rect 80 437 81 438
rect 79 437 80 438
rect 78 437 79 438
rect 77 437 78 438
rect 76 437 77 438
rect 75 437 76 438
rect 74 437 75 438
rect 73 437 74 438
rect 72 437 73 438
rect 71 437 72 438
rect 70 437 71 438
rect 69 437 70 438
rect 68 437 69 438
rect 67 437 68 438
rect 66 437 67 438
rect 65 437 66 438
rect 55 437 56 438
rect 54 437 55 438
rect 53 437 54 438
rect 52 437 53 438
rect 51 437 52 438
rect 50 437 51 438
rect 49 437 50 438
rect 48 437 49 438
rect 47 437 48 438
rect 46 437 47 438
rect 45 437 46 438
rect 44 437 45 438
rect 43 437 44 438
rect 42 437 43 438
rect 41 437 42 438
rect 40 437 41 438
rect 39 437 40 438
rect 38 437 39 438
rect 37 437 38 438
rect 36 437 37 438
rect 35 437 36 438
rect 34 437 35 438
rect 33 437 34 438
rect 32 437 33 438
rect 31 437 32 438
rect 30 437 31 438
rect 29 437 30 438
rect 28 437 29 438
rect 27 437 28 438
rect 26 437 27 438
rect 25 437 26 438
rect 24 437 25 438
rect 23 437 24 438
rect 22 437 23 438
rect 21 437 22 438
rect 20 437 21 438
rect 19 437 20 438
rect 18 437 19 438
rect 17 437 18 438
rect 16 437 17 438
rect 15 437 16 438
rect 14 437 15 438
rect 140 438 141 439
rect 139 438 140 439
rect 138 438 139 439
rect 137 438 138 439
rect 136 438 137 439
rect 135 438 136 439
rect 134 438 135 439
rect 133 438 134 439
rect 132 438 133 439
rect 131 438 132 439
rect 130 438 131 439
rect 129 438 130 439
rect 128 438 129 439
rect 127 438 128 439
rect 126 438 127 439
rect 80 438 81 439
rect 79 438 80 439
rect 78 438 79 439
rect 77 438 78 439
rect 76 438 77 439
rect 75 438 76 439
rect 74 438 75 439
rect 73 438 74 439
rect 72 438 73 439
rect 71 438 72 439
rect 70 438 71 439
rect 69 438 70 439
rect 68 438 69 439
rect 67 438 68 439
rect 66 438 67 439
rect 65 438 66 439
rect 55 438 56 439
rect 54 438 55 439
rect 53 438 54 439
rect 52 438 53 439
rect 51 438 52 439
rect 50 438 51 439
rect 49 438 50 439
rect 48 438 49 439
rect 47 438 48 439
rect 46 438 47 439
rect 45 438 46 439
rect 44 438 45 439
rect 43 438 44 439
rect 42 438 43 439
rect 41 438 42 439
rect 40 438 41 439
rect 39 438 40 439
rect 38 438 39 439
rect 37 438 38 439
rect 36 438 37 439
rect 35 438 36 439
rect 34 438 35 439
rect 33 438 34 439
rect 32 438 33 439
rect 31 438 32 439
rect 30 438 31 439
rect 29 438 30 439
rect 28 438 29 439
rect 27 438 28 439
rect 26 438 27 439
rect 25 438 26 439
rect 24 438 25 439
rect 23 438 24 439
rect 22 438 23 439
rect 21 438 22 439
rect 20 438 21 439
rect 19 438 20 439
rect 18 438 19 439
rect 17 438 18 439
rect 16 438 17 439
rect 15 438 16 439
rect 14 438 15 439
rect 141 439 142 440
rect 140 439 141 440
rect 139 439 140 440
rect 138 439 139 440
rect 137 439 138 440
rect 136 439 137 440
rect 135 439 136 440
rect 134 439 135 440
rect 133 439 134 440
rect 132 439 133 440
rect 131 439 132 440
rect 130 439 131 440
rect 129 439 130 440
rect 128 439 129 440
rect 127 439 128 440
rect 126 439 127 440
rect 125 439 126 440
rect 124 439 125 440
rect 80 439 81 440
rect 79 439 80 440
rect 78 439 79 440
rect 77 439 78 440
rect 76 439 77 440
rect 75 439 76 440
rect 74 439 75 440
rect 73 439 74 440
rect 72 439 73 440
rect 71 439 72 440
rect 70 439 71 440
rect 69 439 70 440
rect 68 439 69 440
rect 67 439 68 440
rect 66 439 67 440
rect 65 439 66 440
rect 54 439 55 440
rect 53 439 54 440
rect 52 439 53 440
rect 51 439 52 440
rect 50 439 51 440
rect 49 439 50 440
rect 48 439 49 440
rect 47 439 48 440
rect 46 439 47 440
rect 45 439 46 440
rect 44 439 45 440
rect 43 439 44 440
rect 42 439 43 440
rect 41 439 42 440
rect 40 439 41 440
rect 39 439 40 440
rect 38 439 39 440
rect 37 439 38 440
rect 36 439 37 440
rect 35 439 36 440
rect 34 439 35 440
rect 33 439 34 440
rect 32 439 33 440
rect 31 439 32 440
rect 30 439 31 440
rect 29 439 30 440
rect 28 439 29 440
rect 27 439 28 440
rect 26 439 27 440
rect 25 439 26 440
rect 24 439 25 440
rect 23 439 24 440
rect 22 439 23 440
rect 21 439 22 440
rect 20 439 21 440
rect 19 439 20 440
rect 18 439 19 440
rect 17 439 18 440
rect 16 439 17 440
rect 15 439 16 440
rect 14 439 15 440
rect 142 440 143 441
rect 141 440 142 441
rect 140 440 141 441
rect 139 440 140 441
rect 138 440 139 441
rect 137 440 138 441
rect 136 440 137 441
rect 135 440 136 441
rect 134 440 135 441
rect 131 440 132 441
rect 130 440 131 441
rect 129 440 130 441
rect 128 440 129 441
rect 127 440 128 441
rect 126 440 127 441
rect 125 440 126 441
rect 124 440 125 441
rect 80 440 81 441
rect 79 440 80 441
rect 78 440 79 441
rect 77 440 78 441
rect 76 440 77 441
rect 75 440 76 441
rect 74 440 75 441
rect 73 440 74 441
rect 72 440 73 441
rect 71 440 72 441
rect 70 440 71 441
rect 69 440 70 441
rect 68 440 69 441
rect 67 440 68 441
rect 66 440 67 441
rect 65 440 66 441
rect 54 440 55 441
rect 53 440 54 441
rect 52 440 53 441
rect 51 440 52 441
rect 50 440 51 441
rect 49 440 50 441
rect 48 440 49 441
rect 47 440 48 441
rect 46 440 47 441
rect 45 440 46 441
rect 44 440 45 441
rect 43 440 44 441
rect 42 440 43 441
rect 41 440 42 441
rect 40 440 41 441
rect 39 440 40 441
rect 38 440 39 441
rect 37 440 38 441
rect 36 440 37 441
rect 35 440 36 441
rect 34 440 35 441
rect 33 440 34 441
rect 32 440 33 441
rect 31 440 32 441
rect 30 440 31 441
rect 29 440 30 441
rect 28 440 29 441
rect 27 440 28 441
rect 26 440 27 441
rect 25 440 26 441
rect 24 440 25 441
rect 23 440 24 441
rect 22 440 23 441
rect 21 440 22 441
rect 20 440 21 441
rect 19 440 20 441
rect 18 440 19 441
rect 17 440 18 441
rect 16 440 17 441
rect 15 440 16 441
rect 14 440 15 441
rect 142 441 143 442
rect 141 441 142 442
rect 140 441 141 442
rect 139 441 140 442
rect 138 441 139 442
rect 137 441 138 442
rect 136 441 137 442
rect 129 441 130 442
rect 128 441 129 442
rect 127 441 128 442
rect 126 441 127 442
rect 125 441 126 442
rect 124 441 125 442
rect 80 441 81 442
rect 79 441 80 442
rect 78 441 79 442
rect 77 441 78 442
rect 76 441 77 442
rect 75 441 76 442
rect 74 441 75 442
rect 73 441 74 442
rect 72 441 73 442
rect 71 441 72 442
rect 70 441 71 442
rect 69 441 70 442
rect 68 441 69 442
rect 67 441 68 442
rect 66 441 67 442
rect 65 441 66 442
rect 53 441 54 442
rect 52 441 53 442
rect 51 441 52 442
rect 50 441 51 442
rect 49 441 50 442
rect 48 441 49 442
rect 47 441 48 442
rect 46 441 47 442
rect 45 441 46 442
rect 44 441 45 442
rect 43 441 44 442
rect 42 441 43 442
rect 41 441 42 442
rect 40 441 41 442
rect 39 441 40 442
rect 38 441 39 442
rect 37 441 38 442
rect 36 441 37 442
rect 35 441 36 442
rect 34 441 35 442
rect 33 441 34 442
rect 32 441 33 442
rect 31 441 32 442
rect 30 441 31 442
rect 29 441 30 442
rect 28 441 29 442
rect 27 441 28 442
rect 26 441 27 442
rect 25 441 26 442
rect 24 441 25 442
rect 23 441 24 442
rect 22 441 23 442
rect 21 441 22 442
rect 20 441 21 442
rect 19 441 20 442
rect 18 441 19 442
rect 17 441 18 442
rect 16 441 17 442
rect 15 441 16 442
rect 142 442 143 443
rect 141 442 142 443
rect 140 442 141 443
rect 139 442 140 443
rect 138 442 139 443
rect 137 442 138 443
rect 128 442 129 443
rect 127 442 128 443
rect 126 442 127 443
rect 125 442 126 443
rect 124 442 125 443
rect 80 442 81 443
rect 79 442 80 443
rect 78 442 79 443
rect 77 442 78 443
rect 76 442 77 443
rect 75 442 76 443
rect 74 442 75 443
rect 73 442 74 443
rect 72 442 73 443
rect 71 442 72 443
rect 70 442 71 443
rect 69 442 70 443
rect 68 442 69 443
rect 67 442 68 443
rect 66 442 67 443
rect 65 442 66 443
rect 52 442 53 443
rect 51 442 52 443
rect 50 442 51 443
rect 49 442 50 443
rect 48 442 49 443
rect 47 442 48 443
rect 46 442 47 443
rect 45 442 46 443
rect 44 442 45 443
rect 43 442 44 443
rect 42 442 43 443
rect 41 442 42 443
rect 40 442 41 443
rect 39 442 40 443
rect 38 442 39 443
rect 37 442 38 443
rect 36 442 37 443
rect 35 442 36 443
rect 34 442 35 443
rect 33 442 34 443
rect 32 442 33 443
rect 31 442 32 443
rect 30 442 31 443
rect 29 442 30 443
rect 28 442 29 443
rect 27 442 28 443
rect 26 442 27 443
rect 25 442 26 443
rect 24 442 25 443
rect 23 442 24 443
rect 22 442 23 443
rect 21 442 22 443
rect 20 442 21 443
rect 19 442 20 443
rect 18 442 19 443
rect 17 442 18 443
rect 16 442 17 443
rect 15 442 16 443
rect 142 443 143 444
rect 141 443 142 444
rect 140 443 141 444
rect 139 443 140 444
rect 138 443 139 444
rect 127 443 128 444
rect 126 443 127 444
rect 125 443 126 444
rect 124 443 125 444
rect 80 443 81 444
rect 79 443 80 444
rect 78 443 79 444
rect 77 443 78 444
rect 76 443 77 444
rect 75 443 76 444
rect 74 443 75 444
rect 73 443 74 444
rect 72 443 73 444
rect 71 443 72 444
rect 70 443 71 444
rect 69 443 70 444
rect 68 443 69 444
rect 67 443 68 444
rect 66 443 67 444
rect 65 443 66 444
rect 51 443 52 444
rect 50 443 51 444
rect 49 443 50 444
rect 48 443 49 444
rect 47 443 48 444
rect 46 443 47 444
rect 45 443 46 444
rect 44 443 45 444
rect 43 443 44 444
rect 42 443 43 444
rect 41 443 42 444
rect 40 443 41 444
rect 39 443 40 444
rect 38 443 39 444
rect 37 443 38 444
rect 36 443 37 444
rect 35 443 36 444
rect 34 443 35 444
rect 33 443 34 444
rect 32 443 33 444
rect 31 443 32 444
rect 30 443 31 444
rect 29 443 30 444
rect 28 443 29 444
rect 27 443 28 444
rect 26 443 27 444
rect 25 443 26 444
rect 24 443 25 444
rect 23 443 24 444
rect 22 443 23 444
rect 21 443 22 444
rect 20 443 21 444
rect 19 443 20 444
rect 18 443 19 444
rect 17 443 18 444
rect 16 443 17 444
rect 142 444 143 445
rect 141 444 142 445
rect 140 444 141 445
rect 125 444 126 445
rect 124 444 125 445
rect 80 444 81 445
rect 79 444 80 445
rect 78 444 79 445
rect 77 444 78 445
rect 76 444 77 445
rect 75 444 76 445
rect 74 444 75 445
rect 73 444 74 445
rect 72 444 73 445
rect 71 444 72 445
rect 70 444 71 445
rect 69 444 70 445
rect 68 444 69 445
rect 67 444 68 445
rect 66 444 67 445
rect 65 444 66 445
rect 51 444 52 445
rect 50 444 51 445
rect 49 444 50 445
rect 48 444 49 445
rect 47 444 48 445
rect 46 444 47 445
rect 45 444 46 445
rect 44 444 45 445
rect 43 444 44 445
rect 42 444 43 445
rect 41 444 42 445
rect 40 444 41 445
rect 39 444 40 445
rect 38 444 39 445
rect 37 444 38 445
rect 36 444 37 445
rect 35 444 36 445
rect 34 444 35 445
rect 33 444 34 445
rect 32 444 33 445
rect 31 444 32 445
rect 30 444 31 445
rect 29 444 30 445
rect 28 444 29 445
rect 27 444 28 445
rect 26 444 27 445
rect 25 444 26 445
rect 24 444 25 445
rect 23 444 24 445
rect 22 444 23 445
rect 21 444 22 445
rect 20 444 21 445
rect 19 444 20 445
rect 18 444 19 445
rect 17 444 18 445
rect 16 444 17 445
rect 142 445 143 446
rect 141 445 142 446
rect 124 445 125 446
rect 80 445 81 446
rect 79 445 80 446
rect 78 445 79 446
rect 77 445 78 446
rect 76 445 77 446
rect 75 445 76 446
rect 74 445 75 446
rect 73 445 74 446
rect 72 445 73 446
rect 71 445 72 446
rect 70 445 71 446
rect 69 445 70 446
rect 68 445 69 446
rect 67 445 68 446
rect 66 445 67 446
rect 65 445 66 446
rect 50 445 51 446
rect 49 445 50 446
rect 48 445 49 446
rect 47 445 48 446
rect 46 445 47 446
rect 45 445 46 446
rect 44 445 45 446
rect 43 445 44 446
rect 42 445 43 446
rect 41 445 42 446
rect 40 445 41 446
rect 39 445 40 446
rect 38 445 39 446
rect 37 445 38 446
rect 36 445 37 446
rect 35 445 36 446
rect 34 445 35 446
rect 33 445 34 446
rect 32 445 33 446
rect 31 445 32 446
rect 30 445 31 446
rect 29 445 30 446
rect 28 445 29 446
rect 27 445 28 446
rect 26 445 27 446
rect 25 445 26 446
rect 24 445 25 446
rect 23 445 24 446
rect 22 445 23 446
rect 21 445 22 446
rect 20 445 21 446
rect 19 445 20 446
rect 18 445 19 446
rect 17 445 18 446
rect 80 446 81 447
rect 79 446 80 447
rect 78 446 79 447
rect 77 446 78 447
rect 76 446 77 447
rect 75 446 76 447
rect 74 446 75 447
rect 73 446 74 447
rect 72 446 73 447
rect 71 446 72 447
rect 70 446 71 447
rect 69 446 70 447
rect 68 446 69 447
rect 67 446 68 447
rect 66 446 67 447
rect 65 446 66 447
rect 49 446 50 447
rect 48 446 49 447
rect 47 446 48 447
rect 46 446 47 447
rect 45 446 46 447
rect 44 446 45 447
rect 43 446 44 447
rect 42 446 43 447
rect 41 446 42 447
rect 40 446 41 447
rect 39 446 40 447
rect 38 446 39 447
rect 37 446 38 447
rect 36 446 37 447
rect 35 446 36 447
rect 34 446 35 447
rect 33 446 34 447
rect 32 446 33 447
rect 31 446 32 447
rect 30 446 31 447
rect 29 446 30 447
rect 28 446 29 447
rect 27 446 28 447
rect 26 446 27 447
rect 25 446 26 447
rect 24 446 25 447
rect 23 446 24 447
rect 22 446 23 447
rect 21 446 22 447
rect 20 446 21 447
rect 19 446 20 447
rect 18 446 19 447
rect 17 446 18 447
rect 80 447 81 448
rect 79 447 80 448
rect 78 447 79 448
rect 77 447 78 448
rect 76 447 77 448
rect 75 447 76 448
rect 74 447 75 448
rect 73 447 74 448
rect 72 447 73 448
rect 71 447 72 448
rect 70 447 71 448
rect 69 447 70 448
rect 68 447 69 448
rect 67 447 68 448
rect 66 447 67 448
rect 65 447 66 448
rect 48 447 49 448
rect 47 447 48 448
rect 46 447 47 448
rect 45 447 46 448
rect 44 447 45 448
rect 43 447 44 448
rect 42 447 43 448
rect 41 447 42 448
rect 40 447 41 448
rect 39 447 40 448
rect 38 447 39 448
rect 37 447 38 448
rect 36 447 37 448
rect 35 447 36 448
rect 34 447 35 448
rect 33 447 34 448
rect 32 447 33 448
rect 31 447 32 448
rect 30 447 31 448
rect 29 447 30 448
rect 28 447 29 448
rect 27 447 28 448
rect 26 447 27 448
rect 25 447 26 448
rect 24 447 25 448
rect 23 447 24 448
rect 22 447 23 448
rect 21 447 22 448
rect 20 447 21 448
rect 19 447 20 448
rect 18 447 19 448
rect 80 448 81 449
rect 79 448 80 449
rect 78 448 79 449
rect 77 448 78 449
rect 76 448 77 449
rect 75 448 76 449
rect 74 448 75 449
rect 73 448 74 449
rect 72 448 73 449
rect 71 448 72 449
rect 70 448 71 449
rect 69 448 70 449
rect 68 448 69 449
rect 67 448 68 449
rect 66 448 67 449
rect 65 448 66 449
rect 47 448 48 449
rect 46 448 47 449
rect 45 448 46 449
rect 44 448 45 449
rect 43 448 44 449
rect 42 448 43 449
rect 41 448 42 449
rect 40 448 41 449
rect 39 448 40 449
rect 38 448 39 449
rect 37 448 38 449
rect 36 448 37 449
rect 35 448 36 449
rect 34 448 35 449
rect 33 448 34 449
rect 32 448 33 449
rect 31 448 32 449
rect 30 448 31 449
rect 29 448 30 449
rect 28 448 29 449
rect 27 448 28 449
rect 26 448 27 449
rect 25 448 26 449
rect 24 448 25 449
rect 23 448 24 449
rect 22 448 23 449
rect 21 448 22 449
rect 20 448 21 449
rect 19 448 20 449
rect 80 449 81 450
rect 79 449 80 450
rect 78 449 79 450
rect 77 449 78 450
rect 76 449 77 450
rect 75 449 76 450
rect 74 449 75 450
rect 73 449 74 450
rect 72 449 73 450
rect 71 449 72 450
rect 70 449 71 450
rect 69 449 70 450
rect 68 449 69 450
rect 67 449 68 450
rect 66 449 67 450
rect 65 449 66 450
rect 46 449 47 450
rect 45 449 46 450
rect 44 449 45 450
rect 43 449 44 450
rect 42 449 43 450
rect 41 449 42 450
rect 40 449 41 450
rect 39 449 40 450
rect 38 449 39 450
rect 37 449 38 450
rect 36 449 37 450
rect 35 449 36 450
rect 34 449 35 450
rect 33 449 34 450
rect 32 449 33 450
rect 31 449 32 450
rect 30 449 31 450
rect 29 449 30 450
rect 28 449 29 450
rect 27 449 28 450
rect 26 449 27 450
rect 25 449 26 450
rect 24 449 25 450
rect 23 449 24 450
rect 22 449 23 450
rect 21 449 22 450
rect 20 449 21 450
rect 80 450 81 451
rect 79 450 80 451
rect 78 450 79 451
rect 77 450 78 451
rect 76 450 77 451
rect 75 450 76 451
rect 74 450 75 451
rect 73 450 74 451
rect 72 450 73 451
rect 71 450 72 451
rect 70 450 71 451
rect 69 450 70 451
rect 68 450 69 451
rect 67 450 68 451
rect 66 450 67 451
rect 65 450 66 451
rect 44 450 45 451
rect 43 450 44 451
rect 42 450 43 451
rect 41 450 42 451
rect 40 450 41 451
rect 39 450 40 451
rect 38 450 39 451
rect 37 450 38 451
rect 36 450 37 451
rect 35 450 36 451
rect 34 450 35 451
rect 33 450 34 451
rect 32 450 33 451
rect 31 450 32 451
rect 30 450 31 451
rect 29 450 30 451
rect 28 450 29 451
rect 27 450 28 451
rect 26 450 27 451
rect 25 450 26 451
rect 24 450 25 451
rect 23 450 24 451
rect 22 450 23 451
rect 21 450 22 451
rect 80 451 81 452
rect 79 451 80 452
rect 78 451 79 452
rect 77 451 78 452
rect 76 451 77 452
rect 75 451 76 452
rect 74 451 75 452
rect 73 451 74 452
rect 72 451 73 452
rect 71 451 72 452
rect 70 451 71 452
rect 69 451 70 452
rect 68 451 69 452
rect 67 451 68 452
rect 66 451 67 452
rect 65 451 66 452
rect 42 451 43 452
rect 41 451 42 452
rect 40 451 41 452
rect 39 451 40 452
rect 38 451 39 452
rect 37 451 38 452
rect 36 451 37 452
rect 35 451 36 452
rect 34 451 35 452
rect 33 451 34 452
rect 32 451 33 452
rect 31 451 32 452
rect 30 451 31 452
rect 29 451 30 452
rect 28 451 29 452
rect 27 451 28 452
rect 26 451 27 452
rect 25 451 26 452
rect 24 451 25 452
rect 23 451 24 452
rect 80 452 81 453
rect 79 452 80 453
rect 78 452 79 453
rect 77 452 78 453
rect 76 452 77 453
rect 75 452 76 453
rect 74 452 75 453
rect 73 452 74 453
rect 72 452 73 453
rect 71 452 72 453
rect 70 452 71 453
rect 69 452 70 453
rect 68 452 69 453
rect 67 452 68 453
rect 66 452 67 453
rect 65 452 66 453
rect 40 452 41 453
rect 39 452 40 453
rect 38 452 39 453
rect 37 452 38 453
rect 36 452 37 453
rect 35 452 36 453
rect 34 452 35 453
rect 33 452 34 453
rect 32 452 33 453
rect 31 452 32 453
rect 30 452 31 453
rect 29 452 30 453
rect 28 452 29 453
rect 27 452 28 453
rect 26 452 27 453
rect 25 452 26 453
rect 80 453 81 454
rect 79 453 80 454
rect 78 453 79 454
rect 77 453 78 454
rect 76 453 77 454
rect 75 453 76 454
rect 74 453 75 454
rect 73 453 74 454
rect 72 453 73 454
rect 71 453 72 454
rect 70 453 71 454
rect 69 453 70 454
rect 68 453 69 454
rect 67 453 68 454
rect 66 453 67 454
rect 65 453 66 454
rect 35 453 36 454
rect 34 453 35 454
rect 33 453 34 454
rect 32 453 33 454
rect 31 453 32 454
rect 30 453 31 454
<< metal2 >>
rect 57 14 58 15
rect 56 14 57 15
rect 55 14 56 15
rect 54 14 55 15
rect 53 14 54 15
rect 52 14 53 15
rect 51 14 52 15
rect 50 14 51 15
rect 49 14 50 15
rect 48 14 49 15
rect 47 14 48 15
rect 46 14 47 15
rect 45 14 46 15
rect 44 14 45 15
rect 61 15 62 16
rect 60 15 61 16
rect 59 15 60 16
rect 58 15 59 16
rect 57 15 58 16
rect 56 15 57 16
rect 55 15 56 16
rect 54 15 55 16
rect 53 15 54 16
rect 52 15 53 16
rect 51 15 52 16
rect 50 15 51 16
rect 49 15 50 16
rect 48 15 49 16
rect 47 15 48 16
rect 46 15 47 16
rect 45 15 46 16
rect 44 15 45 16
rect 43 15 44 16
rect 42 15 43 16
rect 41 15 42 16
rect 40 15 41 16
rect 39 15 40 16
rect 64 16 65 17
rect 63 16 64 17
rect 62 16 63 17
rect 61 16 62 17
rect 60 16 61 17
rect 59 16 60 17
rect 58 16 59 17
rect 57 16 58 17
rect 56 16 57 17
rect 55 16 56 17
rect 54 16 55 17
rect 53 16 54 17
rect 52 16 53 17
rect 51 16 52 17
rect 50 16 51 17
rect 49 16 50 17
rect 48 16 49 17
rect 47 16 48 17
rect 46 16 47 17
rect 45 16 46 17
rect 44 16 45 17
rect 43 16 44 17
rect 42 16 43 17
rect 41 16 42 17
rect 40 16 41 17
rect 39 16 40 17
rect 38 16 39 17
rect 37 16 38 17
rect 36 16 37 17
rect 66 17 67 18
rect 65 17 66 18
rect 64 17 65 18
rect 63 17 64 18
rect 62 17 63 18
rect 61 17 62 18
rect 60 17 61 18
rect 59 17 60 18
rect 58 17 59 18
rect 57 17 58 18
rect 56 17 57 18
rect 55 17 56 18
rect 54 17 55 18
rect 53 17 54 18
rect 52 17 53 18
rect 51 17 52 18
rect 50 17 51 18
rect 49 17 50 18
rect 48 17 49 18
rect 47 17 48 18
rect 46 17 47 18
rect 45 17 46 18
rect 44 17 45 18
rect 43 17 44 18
rect 42 17 43 18
rect 41 17 42 18
rect 40 17 41 18
rect 39 17 40 18
rect 38 17 39 18
rect 37 17 38 18
rect 36 17 37 18
rect 35 17 36 18
rect 34 17 35 18
rect 68 18 69 19
rect 67 18 68 19
rect 66 18 67 19
rect 65 18 66 19
rect 64 18 65 19
rect 63 18 64 19
rect 62 18 63 19
rect 61 18 62 19
rect 60 18 61 19
rect 59 18 60 19
rect 58 18 59 19
rect 57 18 58 19
rect 56 18 57 19
rect 55 18 56 19
rect 54 18 55 19
rect 53 18 54 19
rect 52 18 53 19
rect 51 18 52 19
rect 50 18 51 19
rect 49 18 50 19
rect 48 18 49 19
rect 47 18 48 19
rect 46 18 47 19
rect 45 18 46 19
rect 44 18 45 19
rect 43 18 44 19
rect 42 18 43 19
rect 41 18 42 19
rect 40 18 41 19
rect 39 18 40 19
rect 38 18 39 19
rect 37 18 38 19
rect 36 18 37 19
rect 35 18 36 19
rect 34 18 35 19
rect 33 18 34 19
rect 32 18 33 19
rect 70 19 71 20
rect 69 19 70 20
rect 68 19 69 20
rect 67 19 68 20
rect 66 19 67 20
rect 65 19 66 20
rect 64 19 65 20
rect 63 19 64 20
rect 62 19 63 20
rect 61 19 62 20
rect 60 19 61 20
rect 59 19 60 20
rect 58 19 59 20
rect 57 19 58 20
rect 56 19 57 20
rect 55 19 56 20
rect 54 19 55 20
rect 53 19 54 20
rect 52 19 53 20
rect 51 19 52 20
rect 50 19 51 20
rect 49 19 50 20
rect 48 19 49 20
rect 47 19 48 20
rect 46 19 47 20
rect 45 19 46 20
rect 44 19 45 20
rect 43 19 44 20
rect 42 19 43 20
rect 41 19 42 20
rect 40 19 41 20
rect 39 19 40 20
rect 38 19 39 20
rect 37 19 38 20
rect 36 19 37 20
rect 35 19 36 20
rect 34 19 35 20
rect 33 19 34 20
rect 32 19 33 20
rect 31 19 32 20
rect 71 20 72 21
rect 70 20 71 21
rect 69 20 70 21
rect 68 20 69 21
rect 67 20 68 21
rect 66 20 67 21
rect 65 20 66 21
rect 64 20 65 21
rect 63 20 64 21
rect 62 20 63 21
rect 61 20 62 21
rect 60 20 61 21
rect 59 20 60 21
rect 58 20 59 21
rect 57 20 58 21
rect 56 20 57 21
rect 55 20 56 21
rect 54 20 55 21
rect 53 20 54 21
rect 52 20 53 21
rect 51 20 52 21
rect 50 20 51 21
rect 49 20 50 21
rect 48 20 49 21
rect 47 20 48 21
rect 46 20 47 21
rect 45 20 46 21
rect 44 20 45 21
rect 43 20 44 21
rect 42 20 43 21
rect 41 20 42 21
rect 40 20 41 21
rect 39 20 40 21
rect 38 20 39 21
rect 37 20 38 21
rect 36 20 37 21
rect 35 20 36 21
rect 34 20 35 21
rect 33 20 34 21
rect 32 20 33 21
rect 31 20 32 21
rect 30 20 31 21
rect 29 20 30 21
rect 72 21 73 22
rect 71 21 72 22
rect 70 21 71 22
rect 69 21 70 22
rect 68 21 69 22
rect 67 21 68 22
rect 66 21 67 22
rect 65 21 66 22
rect 64 21 65 22
rect 63 21 64 22
rect 62 21 63 22
rect 61 21 62 22
rect 60 21 61 22
rect 59 21 60 22
rect 58 21 59 22
rect 57 21 58 22
rect 56 21 57 22
rect 55 21 56 22
rect 54 21 55 22
rect 53 21 54 22
rect 52 21 53 22
rect 51 21 52 22
rect 50 21 51 22
rect 49 21 50 22
rect 48 21 49 22
rect 47 21 48 22
rect 46 21 47 22
rect 45 21 46 22
rect 44 21 45 22
rect 43 21 44 22
rect 42 21 43 22
rect 41 21 42 22
rect 40 21 41 22
rect 39 21 40 22
rect 38 21 39 22
rect 37 21 38 22
rect 36 21 37 22
rect 35 21 36 22
rect 34 21 35 22
rect 33 21 34 22
rect 32 21 33 22
rect 31 21 32 22
rect 30 21 31 22
rect 29 21 30 22
rect 28 21 29 22
rect 73 22 74 23
rect 72 22 73 23
rect 71 22 72 23
rect 70 22 71 23
rect 69 22 70 23
rect 68 22 69 23
rect 67 22 68 23
rect 66 22 67 23
rect 65 22 66 23
rect 64 22 65 23
rect 63 22 64 23
rect 62 22 63 23
rect 61 22 62 23
rect 60 22 61 23
rect 59 22 60 23
rect 58 22 59 23
rect 57 22 58 23
rect 56 22 57 23
rect 55 22 56 23
rect 54 22 55 23
rect 53 22 54 23
rect 52 22 53 23
rect 51 22 52 23
rect 50 22 51 23
rect 49 22 50 23
rect 48 22 49 23
rect 47 22 48 23
rect 46 22 47 23
rect 45 22 46 23
rect 44 22 45 23
rect 43 22 44 23
rect 42 22 43 23
rect 41 22 42 23
rect 40 22 41 23
rect 39 22 40 23
rect 38 22 39 23
rect 37 22 38 23
rect 36 22 37 23
rect 35 22 36 23
rect 34 22 35 23
rect 33 22 34 23
rect 32 22 33 23
rect 31 22 32 23
rect 30 22 31 23
rect 29 22 30 23
rect 28 22 29 23
rect 27 22 28 23
rect 74 23 75 24
rect 73 23 74 24
rect 72 23 73 24
rect 71 23 72 24
rect 70 23 71 24
rect 69 23 70 24
rect 68 23 69 24
rect 67 23 68 24
rect 66 23 67 24
rect 65 23 66 24
rect 64 23 65 24
rect 63 23 64 24
rect 62 23 63 24
rect 61 23 62 24
rect 60 23 61 24
rect 59 23 60 24
rect 58 23 59 24
rect 57 23 58 24
rect 56 23 57 24
rect 55 23 56 24
rect 54 23 55 24
rect 53 23 54 24
rect 52 23 53 24
rect 51 23 52 24
rect 50 23 51 24
rect 49 23 50 24
rect 48 23 49 24
rect 47 23 48 24
rect 46 23 47 24
rect 45 23 46 24
rect 44 23 45 24
rect 43 23 44 24
rect 42 23 43 24
rect 41 23 42 24
rect 40 23 41 24
rect 39 23 40 24
rect 38 23 39 24
rect 37 23 38 24
rect 36 23 37 24
rect 35 23 36 24
rect 34 23 35 24
rect 33 23 34 24
rect 32 23 33 24
rect 31 23 32 24
rect 30 23 31 24
rect 29 23 30 24
rect 28 23 29 24
rect 27 23 28 24
rect 26 23 27 24
rect 25 23 26 24
rect 75 24 76 25
rect 74 24 75 25
rect 73 24 74 25
rect 72 24 73 25
rect 71 24 72 25
rect 70 24 71 25
rect 69 24 70 25
rect 68 24 69 25
rect 67 24 68 25
rect 66 24 67 25
rect 65 24 66 25
rect 64 24 65 25
rect 63 24 64 25
rect 62 24 63 25
rect 61 24 62 25
rect 60 24 61 25
rect 59 24 60 25
rect 58 24 59 25
rect 57 24 58 25
rect 56 24 57 25
rect 55 24 56 25
rect 54 24 55 25
rect 53 24 54 25
rect 52 24 53 25
rect 51 24 52 25
rect 50 24 51 25
rect 49 24 50 25
rect 48 24 49 25
rect 47 24 48 25
rect 46 24 47 25
rect 45 24 46 25
rect 44 24 45 25
rect 43 24 44 25
rect 42 24 43 25
rect 41 24 42 25
rect 40 24 41 25
rect 39 24 40 25
rect 38 24 39 25
rect 37 24 38 25
rect 36 24 37 25
rect 35 24 36 25
rect 34 24 35 25
rect 33 24 34 25
rect 32 24 33 25
rect 31 24 32 25
rect 30 24 31 25
rect 29 24 30 25
rect 28 24 29 25
rect 27 24 28 25
rect 26 24 27 25
rect 25 24 26 25
rect 24 24 25 25
rect 76 25 77 26
rect 75 25 76 26
rect 74 25 75 26
rect 73 25 74 26
rect 72 25 73 26
rect 71 25 72 26
rect 70 25 71 26
rect 69 25 70 26
rect 68 25 69 26
rect 67 25 68 26
rect 66 25 67 26
rect 65 25 66 26
rect 64 25 65 26
rect 63 25 64 26
rect 62 25 63 26
rect 61 25 62 26
rect 60 25 61 26
rect 59 25 60 26
rect 58 25 59 26
rect 57 25 58 26
rect 56 25 57 26
rect 55 25 56 26
rect 54 25 55 26
rect 53 25 54 26
rect 52 25 53 26
rect 51 25 52 26
rect 50 25 51 26
rect 49 25 50 26
rect 48 25 49 26
rect 47 25 48 26
rect 46 25 47 26
rect 45 25 46 26
rect 44 25 45 26
rect 43 25 44 26
rect 42 25 43 26
rect 41 25 42 26
rect 40 25 41 26
rect 39 25 40 26
rect 38 25 39 26
rect 37 25 38 26
rect 36 25 37 26
rect 35 25 36 26
rect 34 25 35 26
rect 33 25 34 26
rect 32 25 33 26
rect 31 25 32 26
rect 30 25 31 26
rect 29 25 30 26
rect 28 25 29 26
rect 27 25 28 26
rect 26 25 27 26
rect 25 25 26 26
rect 24 25 25 26
rect 77 26 78 27
rect 76 26 77 27
rect 75 26 76 27
rect 74 26 75 27
rect 73 26 74 27
rect 72 26 73 27
rect 71 26 72 27
rect 70 26 71 27
rect 69 26 70 27
rect 68 26 69 27
rect 67 26 68 27
rect 66 26 67 27
rect 65 26 66 27
rect 64 26 65 27
rect 63 26 64 27
rect 62 26 63 27
rect 61 26 62 27
rect 60 26 61 27
rect 59 26 60 27
rect 58 26 59 27
rect 57 26 58 27
rect 56 26 57 27
rect 55 26 56 27
rect 54 26 55 27
rect 53 26 54 27
rect 52 26 53 27
rect 51 26 52 27
rect 50 26 51 27
rect 49 26 50 27
rect 48 26 49 27
rect 47 26 48 27
rect 46 26 47 27
rect 45 26 46 27
rect 44 26 45 27
rect 43 26 44 27
rect 42 26 43 27
rect 41 26 42 27
rect 40 26 41 27
rect 39 26 40 27
rect 38 26 39 27
rect 37 26 38 27
rect 36 26 37 27
rect 35 26 36 27
rect 34 26 35 27
rect 33 26 34 27
rect 32 26 33 27
rect 31 26 32 27
rect 30 26 31 27
rect 29 26 30 27
rect 28 26 29 27
rect 27 26 28 27
rect 26 26 27 27
rect 25 26 26 27
rect 24 26 25 27
rect 23 26 24 27
rect 78 27 79 28
rect 77 27 78 28
rect 76 27 77 28
rect 75 27 76 28
rect 74 27 75 28
rect 73 27 74 28
rect 72 27 73 28
rect 71 27 72 28
rect 70 27 71 28
rect 69 27 70 28
rect 68 27 69 28
rect 67 27 68 28
rect 66 27 67 28
rect 65 27 66 28
rect 64 27 65 28
rect 63 27 64 28
rect 62 27 63 28
rect 61 27 62 28
rect 60 27 61 28
rect 59 27 60 28
rect 58 27 59 28
rect 57 27 58 28
rect 56 27 57 28
rect 55 27 56 28
rect 54 27 55 28
rect 53 27 54 28
rect 52 27 53 28
rect 51 27 52 28
rect 50 27 51 28
rect 49 27 50 28
rect 48 27 49 28
rect 47 27 48 28
rect 46 27 47 28
rect 45 27 46 28
rect 44 27 45 28
rect 43 27 44 28
rect 42 27 43 28
rect 41 27 42 28
rect 40 27 41 28
rect 39 27 40 28
rect 38 27 39 28
rect 37 27 38 28
rect 36 27 37 28
rect 35 27 36 28
rect 34 27 35 28
rect 33 27 34 28
rect 32 27 33 28
rect 31 27 32 28
rect 30 27 31 28
rect 29 27 30 28
rect 28 27 29 28
rect 27 27 28 28
rect 26 27 27 28
rect 25 27 26 28
rect 24 27 25 28
rect 23 27 24 28
rect 22 27 23 28
rect 78 28 79 29
rect 77 28 78 29
rect 76 28 77 29
rect 75 28 76 29
rect 74 28 75 29
rect 73 28 74 29
rect 72 28 73 29
rect 71 28 72 29
rect 70 28 71 29
rect 69 28 70 29
rect 68 28 69 29
rect 67 28 68 29
rect 66 28 67 29
rect 65 28 66 29
rect 64 28 65 29
rect 63 28 64 29
rect 62 28 63 29
rect 61 28 62 29
rect 60 28 61 29
rect 59 28 60 29
rect 58 28 59 29
rect 57 28 58 29
rect 56 28 57 29
rect 55 28 56 29
rect 54 28 55 29
rect 53 28 54 29
rect 52 28 53 29
rect 51 28 52 29
rect 50 28 51 29
rect 49 28 50 29
rect 48 28 49 29
rect 47 28 48 29
rect 46 28 47 29
rect 45 28 46 29
rect 44 28 45 29
rect 43 28 44 29
rect 42 28 43 29
rect 41 28 42 29
rect 40 28 41 29
rect 39 28 40 29
rect 38 28 39 29
rect 37 28 38 29
rect 36 28 37 29
rect 35 28 36 29
rect 34 28 35 29
rect 33 28 34 29
rect 32 28 33 29
rect 31 28 32 29
rect 30 28 31 29
rect 29 28 30 29
rect 28 28 29 29
rect 27 28 28 29
rect 26 28 27 29
rect 25 28 26 29
rect 24 28 25 29
rect 23 28 24 29
rect 22 28 23 29
rect 21 28 22 29
rect 79 29 80 30
rect 78 29 79 30
rect 77 29 78 30
rect 76 29 77 30
rect 75 29 76 30
rect 74 29 75 30
rect 73 29 74 30
rect 72 29 73 30
rect 71 29 72 30
rect 70 29 71 30
rect 69 29 70 30
rect 68 29 69 30
rect 67 29 68 30
rect 66 29 67 30
rect 65 29 66 30
rect 64 29 65 30
rect 63 29 64 30
rect 62 29 63 30
rect 61 29 62 30
rect 60 29 61 30
rect 59 29 60 30
rect 58 29 59 30
rect 57 29 58 30
rect 56 29 57 30
rect 55 29 56 30
rect 54 29 55 30
rect 53 29 54 30
rect 52 29 53 30
rect 51 29 52 30
rect 50 29 51 30
rect 49 29 50 30
rect 48 29 49 30
rect 47 29 48 30
rect 46 29 47 30
rect 45 29 46 30
rect 44 29 45 30
rect 43 29 44 30
rect 42 29 43 30
rect 41 29 42 30
rect 40 29 41 30
rect 39 29 40 30
rect 38 29 39 30
rect 37 29 38 30
rect 36 29 37 30
rect 35 29 36 30
rect 34 29 35 30
rect 33 29 34 30
rect 32 29 33 30
rect 31 29 32 30
rect 30 29 31 30
rect 29 29 30 30
rect 28 29 29 30
rect 27 29 28 30
rect 26 29 27 30
rect 25 29 26 30
rect 24 29 25 30
rect 23 29 24 30
rect 22 29 23 30
rect 21 29 22 30
rect 79 30 80 31
rect 78 30 79 31
rect 77 30 78 31
rect 76 30 77 31
rect 75 30 76 31
rect 74 30 75 31
rect 73 30 74 31
rect 72 30 73 31
rect 71 30 72 31
rect 70 30 71 31
rect 69 30 70 31
rect 68 30 69 31
rect 67 30 68 31
rect 66 30 67 31
rect 65 30 66 31
rect 64 30 65 31
rect 63 30 64 31
rect 62 30 63 31
rect 61 30 62 31
rect 60 30 61 31
rect 59 30 60 31
rect 58 30 59 31
rect 57 30 58 31
rect 56 30 57 31
rect 55 30 56 31
rect 54 30 55 31
rect 53 30 54 31
rect 52 30 53 31
rect 51 30 52 31
rect 50 30 51 31
rect 49 30 50 31
rect 48 30 49 31
rect 47 30 48 31
rect 46 30 47 31
rect 45 30 46 31
rect 44 30 45 31
rect 43 30 44 31
rect 42 30 43 31
rect 41 30 42 31
rect 40 30 41 31
rect 39 30 40 31
rect 38 30 39 31
rect 37 30 38 31
rect 36 30 37 31
rect 35 30 36 31
rect 34 30 35 31
rect 33 30 34 31
rect 32 30 33 31
rect 31 30 32 31
rect 30 30 31 31
rect 29 30 30 31
rect 28 30 29 31
rect 27 30 28 31
rect 26 30 27 31
rect 25 30 26 31
rect 24 30 25 31
rect 23 30 24 31
rect 22 30 23 31
rect 21 30 22 31
rect 20 30 21 31
rect 80 31 81 32
rect 79 31 80 32
rect 78 31 79 32
rect 77 31 78 32
rect 76 31 77 32
rect 75 31 76 32
rect 74 31 75 32
rect 73 31 74 32
rect 72 31 73 32
rect 71 31 72 32
rect 70 31 71 32
rect 69 31 70 32
rect 68 31 69 32
rect 67 31 68 32
rect 66 31 67 32
rect 65 31 66 32
rect 64 31 65 32
rect 63 31 64 32
rect 62 31 63 32
rect 61 31 62 32
rect 60 31 61 32
rect 59 31 60 32
rect 58 31 59 32
rect 57 31 58 32
rect 56 31 57 32
rect 55 31 56 32
rect 54 31 55 32
rect 53 31 54 32
rect 52 31 53 32
rect 51 31 52 32
rect 50 31 51 32
rect 49 31 50 32
rect 48 31 49 32
rect 47 31 48 32
rect 46 31 47 32
rect 45 31 46 32
rect 44 31 45 32
rect 43 31 44 32
rect 42 31 43 32
rect 41 31 42 32
rect 40 31 41 32
rect 39 31 40 32
rect 38 31 39 32
rect 37 31 38 32
rect 36 31 37 32
rect 35 31 36 32
rect 34 31 35 32
rect 33 31 34 32
rect 32 31 33 32
rect 31 31 32 32
rect 30 31 31 32
rect 29 31 30 32
rect 28 31 29 32
rect 27 31 28 32
rect 26 31 27 32
rect 25 31 26 32
rect 24 31 25 32
rect 23 31 24 32
rect 22 31 23 32
rect 21 31 22 32
rect 20 31 21 32
rect 80 32 81 33
rect 79 32 80 33
rect 78 32 79 33
rect 77 32 78 33
rect 76 32 77 33
rect 75 32 76 33
rect 74 32 75 33
rect 73 32 74 33
rect 72 32 73 33
rect 71 32 72 33
rect 70 32 71 33
rect 69 32 70 33
rect 68 32 69 33
rect 67 32 68 33
rect 66 32 67 33
rect 65 32 66 33
rect 64 32 65 33
rect 63 32 64 33
rect 62 32 63 33
rect 61 32 62 33
rect 60 32 61 33
rect 59 32 60 33
rect 58 32 59 33
rect 57 32 58 33
rect 56 32 57 33
rect 55 32 56 33
rect 54 32 55 33
rect 53 32 54 33
rect 52 32 53 33
rect 51 32 52 33
rect 50 32 51 33
rect 49 32 50 33
rect 48 32 49 33
rect 47 32 48 33
rect 46 32 47 33
rect 45 32 46 33
rect 44 32 45 33
rect 43 32 44 33
rect 42 32 43 33
rect 41 32 42 33
rect 40 32 41 33
rect 39 32 40 33
rect 38 32 39 33
rect 37 32 38 33
rect 36 32 37 33
rect 35 32 36 33
rect 34 32 35 33
rect 33 32 34 33
rect 32 32 33 33
rect 31 32 32 33
rect 30 32 31 33
rect 29 32 30 33
rect 28 32 29 33
rect 27 32 28 33
rect 26 32 27 33
rect 25 32 26 33
rect 24 32 25 33
rect 23 32 24 33
rect 22 32 23 33
rect 21 32 22 33
rect 20 32 21 33
rect 19 32 20 33
rect 144 33 145 34
rect 143 33 144 34
rect 142 33 143 34
rect 141 33 142 34
rect 140 33 141 34
rect 139 33 140 34
rect 81 33 82 34
rect 80 33 81 34
rect 79 33 80 34
rect 78 33 79 34
rect 77 33 78 34
rect 76 33 77 34
rect 75 33 76 34
rect 74 33 75 34
rect 73 33 74 34
rect 72 33 73 34
rect 71 33 72 34
rect 70 33 71 34
rect 69 33 70 34
rect 68 33 69 34
rect 67 33 68 34
rect 66 33 67 34
rect 65 33 66 34
rect 64 33 65 34
rect 63 33 64 34
rect 62 33 63 34
rect 61 33 62 34
rect 60 33 61 34
rect 59 33 60 34
rect 58 33 59 34
rect 57 33 58 34
rect 56 33 57 34
rect 55 33 56 34
rect 54 33 55 34
rect 53 33 54 34
rect 52 33 53 34
rect 51 33 52 34
rect 50 33 51 34
rect 49 33 50 34
rect 48 33 49 34
rect 47 33 48 34
rect 46 33 47 34
rect 45 33 46 34
rect 44 33 45 34
rect 43 33 44 34
rect 42 33 43 34
rect 41 33 42 34
rect 40 33 41 34
rect 39 33 40 34
rect 38 33 39 34
rect 37 33 38 34
rect 36 33 37 34
rect 35 33 36 34
rect 34 33 35 34
rect 33 33 34 34
rect 32 33 33 34
rect 31 33 32 34
rect 30 33 31 34
rect 29 33 30 34
rect 28 33 29 34
rect 27 33 28 34
rect 26 33 27 34
rect 25 33 26 34
rect 24 33 25 34
rect 23 33 24 34
rect 22 33 23 34
rect 21 33 22 34
rect 20 33 21 34
rect 19 33 20 34
rect 144 34 145 35
rect 143 34 144 35
rect 142 34 143 35
rect 141 34 142 35
rect 140 34 141 35
rect 139 34 140 35
rect 138 34 139 35
rect 137 34 138 35
rect 124 34 125 35
rect 123 34 124 35
rect 122 34 123 35
rect 121 34 122 35
rect 81 34 82 35
rect 80 34 81 35
rect 79 34 80 35
rect 78 34 79 35
rect 77 34 78 35
rect 76 34 77 35
rect 75 34 76 35
rect 74 34 75 35
rect 73 34 74 35
rect 72 34 73 35
rect 71 34 72 35
rect 70 34 71 35
rect 69 34 70 35
rect 68 34 69 35
rect 67 34 68 35
rect 66 34 67 35
rect 65 34 66 35
rect 64 34 65 35
rect 63 34 64 35
rect 62 34 63 35
rect 61 34 62 35
rect 60 34 61 35
rect 59 34 60 35
rect 58 34 59 35
rect 57 34 58 35
rect 56 34 57 35
rect 55 34 56 35
rect 54 34 55 35
rect 53 34 54 35
rect 52 34 53 35
rect 51 34 52 35
rect 50 34 51 35
rect 49 34 50 35
rect 48 34 49 35
rect 47 34 48 35
rect 46 34 47 35
rect 45 34 46 35
rect 44 34 45 35
rect 43 34 44 35
rect 42 34 43 35
rect 41 34 42 35
rect 40 34 41 35
rect 39 34 40 35
rect 38 34 39 35
rect 37 34 38 35
rect 36 34 37 35
rect 35 34 36 35
rect 34 34 35 35
rect 33 34 34 35
rect 32 34 33 35
rect 31 34 32 35
rect 30 34 31 35
rect 29 34 30 35
rect 28 34 29 35
rect 27 34 28 35
rect 26 34 27 35
rect 25 34 26 35
rect 24 34 25 35
rect 23 34 24 35
rect 22 34 23 35
rect 21 34 22 35
rect 20 34 21 35
rect 19 34 20 35
rect 18 34 19 35
rect 144 35 145 36
rect 143 35 144 36
rect 142 35 143 36
rect 141 35 142 36
rect 140 35 141 36
rect 139 35 140 36
rect 138 35 139 36
rect 137 35 138 36
rect 136 35 137 36
rect 124 35 125 36
rect 123 35 124 36
rect 122 35 123 36
rect 121 35 122 36
rect 120 35 121 36
rect 81 35 82 36
rect 80 35 81 36
rect 79 35 80 36
rect 78 35 79 36
rect 77 35 78 36
rect 76 35 77 36
rect 75 35 76 36
rect 74 35 75 36
rect 73 35 74 36
rect 72 35 73 36
rect 71 35 72 36
rect 70 35 71 36
rect 69 35 70 36
rect 68 35 69 36
rect 67 35 68 36
rect 66 35 67 36
rect 65 35 66 36
rect 64 35 65 36
rect 63 35 64 36
rect 62 35 63 36
rect 61 35 62 36
rect 60 35 61 36
rect 59 35 60 36
rect 58 35 59 36
rect 57 35 58 36
rect 56 35 57 36
rect 55 35 56 36
rect 54 35 55 36
rect 53 35 54 36
rect 45 35 46 36
rect 44 35 45 36
rect 43 35 44 36
rect 42 35 43 36
rect 41 35 42 36
rect 40 35 41 36
rect 39 35 40 36
rect 38 35 39 36
rect 37 35 38 36
rect 36 35 37 36
rect 35 35 36 36
rect 34 35 35 36
rect 33 35 34 36
rect 32 35 33 36
rect 31 35 32 36
rect 30 35 31 36
rect 29 35 30 36
rect 28 35 29 36
rect 27 35 28 36
rect 26 35 27 36
rect 25 35 26 36
rect 24 35 25 36
rect 23 35 24 36
rect 22 35 23 36
rect 21 35 22 36
rect 20 35 21 36
rect 19 35 20 36
rect 18 35 19 36
rect 144 36 145 37
rect 143 36 144 37
rect 142 36 143 37
rect 141 36 142 37
rect 140 36 141 37
rect 139 36 140 37
rect 138 36 139 37
rect 137 36 138 37
rect 136 36 137 37
rect 135 36 136 37
rect 123 36 124 37
rect 122 36 123 37
rect 121 36 122 37
rect 120 36 121 37
rect 81 36 82 37
rect 80 36 81 37
rect 79 36 80 37
rect 78 36 79 37
rect 77 36 78 37
rect 76 36 77 37
rect 75 36 76 37
rect 74 36 75 37
rect 73 36 74 37
rect 72 36 73 37
rect 71 36 72 37
rect 70 36 71 37
rect 69 36 70 37
rect 68 36 69 37
rect 67 36 68 37
rect 66 36 67 37
rect 65 36 66 37
rect 64 36 65 37
rect 63 36 64 37
rect 62 36 63 37
rect 61 36 62 37
rect 60 36 61 37
rect 59 36 60 37
rect 58 36 59 37
rect 57 36 58 37
rect 41 36 42 37
rect 40 36 41 37
rect 39 36 40 37
rect 38 36 39 37
rect 37 36 38 37
rect 36 36 37 37
rect 35 36 36 37
rect 34 36 35 37
rect 33 36 34 37
rect 32 36 33 37
rect 31 36 32 37
rect 30 36 31 37
rect 29 36 30 37
rect 28 36 29 37
rect 27 36 28 37
rect 26 36 27 37
rect 25 36 26 37
rect 24 36 25 37
rect 23 36 24 37
rect 22 36 23 37
rect 21 36 22 37
rect 20 36 21 37
rect 19 36 20 37
rect 18 36 19 37
rect 17 36 18 37
rect 144 37 145 38
rect 143 37 144 38
rect 142 37 143 38
rect 141 37 142 38
rect 140 37 141 38
rect 139 37 140 38
rect 138 37 139 38
rect 137 37 138 38
rect 136 37 137 38
rect 135 37 136 38
rect 134 37 135 38
rect 123 37 124 38
rect 122 37 123 38
rect 121 37 122 38
rect 120 37 121 38
rect 82 37 83 38
rect 81 37 82 38
rect 80 37 81 38
rect 79 37 80 38
rect 78 37 79 38
rect 77 37 78 38
rect 76 37 77 38
rect 75 37 76 38
rect 74 37 75 38
rect 73 37 74 38
rect 72 37 73 38
rect 71 37 72 38
rect 70 37 71 38
rect 69 37 70 38
rect 68 37 69 38
rect 67 37 68 38
rect 66 37 67 38
rect 65 37 66 38
rect 64 37 65 38
rect 63 37 64 38
rect 62 37 63 38
rect 61 37 62 38
rect 60 37 61 38
rect 59 37 60 38
rect 39 37 40 38
rect 38 37 39 38
rect 37 37 38 38
rect 36 37 37 38
rect 35 37 36 38
rect 34 37 35 38
rect 33 37 34 38
rect 32 37 33 38
rect 31 37 32 38
rect 30 37 31 38
rect 29 37 30 38
rect 28 37 29 38
rect 27 37 28 38
rect 26 37 27 38
rect 25 37 26 38
rect 24 37 25 38
rect 23 37 24 38
rect 22 37 23 38
rect 21 37 22 38
rect 20 37 21 38
rect 19 37 20 38
rect 18 37 19 38
rect 17 37 18 38
rect 144 38 145 39
rect 143 38 144 39
rect 142 38 143 39
rect 141 38 142 39
rect 140 38 141 39
rect 139 38 140 39
rect 138 38 139 39
rect 137 38 138 39
rect 136 38 137 39
rect 135 38 136 39
rect 134 38 135 39
rect 123 38 124 39
rect 122 38 123 39
rect 121 38 122 39
rect 120 38 121 39
rect 119 38 120 39
rect 82 38 83 39
rect 81 38 82 39
rect 80 38 81 39
rect 79 38 80 39
rect 78 38 79 39
rect 77 38 78 39
rect 76 38 77 39
rect 75 38 76 39
rect 74 38 75 39
rect 73 38 74 39
rect 72 38 73 39
rect 71 38 72 39
rect 70 38 71 39
rect 69 38 70 39
rect 68 38 69 39
rect 67 38 68 39
rect 66 38 67 39
rect 65 38 66 39
rect 64 38 65 39
rect 63 38 64 39
rect 62 38 63 39
rect 61 38 62 39
rect 60 38 61 39
rect 38 38 39 39
rect 37 38 38 39
rect 36 38 37 39
rect 35 38 36 39
rect 34 38 35 39
rect 33 38 34 39
rect 32 38 33 39
rect 31 38 32 39
rect 30 38 31 39
rect 29 38 30 39
rect 28 38 29 39
rect 27 38 28 39
rect 26 38 27 39
rect 25 38 26 39
rect 24 38 25 39
rect 23 38 24 39
rect 22 38 23 39
rect 21 38 22 39
rect 20 38 21 39
rect 19 38 20 39
rect 18 38 19 39
rect 17 38 18 39
rect 144 39 145 40
rect 143 39 144 40
rect 142 39 143 40
rect 141 39 142 40
rect 140 39 141 40
rect 138 39 139 40
rect 137 39 138 40
rect 136 39 137 40
rect 135 39 136 40
rect 134 39 135 40
rect 133 39 134 40
rect 122 39 123 40
rect 121 39 122 40
rect 120 39 121 40
rect 119 39 120 40
rect 82 39 83 40
rect 81 39 82 40
rect 80 39 81 40
rect 79 39 80 40
rect 78 39 79 40
rect 77 39 78 40
rect 76 39 77 40
rect 75 39 76 40
rect 74 39 75 40
rect 73 39 74 40
rect 72 39 73 40
rect 71 39 72 40
rect 70 39 71 40
rect 69 39 70 40
rect 68 39 69 40
rect 67 39 68 40
rect 66 39 67 40
rect 65 39 66 40
rect 64 39 65 40
rect 63 39 64 40
rect 62 39 63 40
rect 36 39 37 40
rect 35 39 36 40
rect 34 39 35 40
rect 33 39 34 40
rect 32 39 33 40
rect 31 39 32 40
rect 30 39 31 40
rect 29 39 30 40
rect 28 39 29 40
rect 27 39 28 40
rect 26 39 27 40
rect 25 39 26 40
rect 24 39 25 40
rect 23 39 24 40
rect 22 39 23 40
rect 21 39 22 40
rect 20 39 21 40
rect 19 39 20 40
rect 18 39 19 40
rect 17 39 18 40
rect 16 39 17 40
rect 144 40 145 41
rect 143 40 144 41
rect 142 40 143 41
rect 141 40 142 41
rect 140 40 141 41
rect 137 40 138 41
rect 136 40 137 41
rect 135 40 136 41
rect 134 40 135 41
rect 133 40 134 41
rect 132 40 133 41
rect 122 40 123 41
rect 121 40 122 41
rect 120 40 121 41
rect 119 40 120 41
rect 82 40 83 41
rect 81 40 82 41
rect 80 40 81 41
rect 79 40 80 41
rect 78 40 79 41
rect 77 40 78 41
rect 76 40 77 41
rect 75 40 76 41
rect 74 40 75 41
rect 73 40 74 41
rect 72 40 73 41
rect 71 40 72 41
rect 70 40 71 41
rect 69 40 70 41
rect 68 40 69 41
rect 67 40 68 41
rect 66 40 67 41
rect 65 40 66 41
rect 64 40 65 41
rect 63 40 64 41
rect 35 40 36 41
rect 34 40 35 41
rect 33 40 34 41
rect 32 40 33 41
rect 31 40 32 41
rect 30 40 31 41
rect 29 40 30 41
rect 28 40 29 41
rect 27 40 28 41
rect 26 40 27 41
rect 25 40 26 41
rect 24 40 25 41
rect 23 40 24 41
rect 22 40 23 41
rect 21 40 22 41
rect 20 40 21 41
rect 19 40 20 41
rect 18 40 19 41
rect 17 40 18 41
rect 16 40 17 41
rect 144 41 145 42
rect 143 41 144 42
rect 142 41 143 42
rect 141 41 142 42
rect 140 41 141 42
rect 136 41 137 42
rect 135 41 136 42
rect 134 41 135 42
rect 133 41 134 42
rect 132 41 133 42
rect 131 41 132 42
rect 123 41 124 42
rect 122 41 123 42
rect 121 41 122 42
rect 120 41 121 42
rect 119 41 120 42
rect 82 41 83 42
rect 81 41 82 42
rect 80 41 81 42
rect 79 41 80 42
rect 78 41 79 42
rect 77 41 78 42
rect 76 41 77 42
rect 75 41 76 42
rect 74 41 75 42
rect 73 41 74 42
rect 72 41 73 42
rect 71 41 72 42
rect 70 41 71 42
rect 69 41 70 42
rect 68 41 69 42
rect 67 41 68 42
rect 66 41 67 42
rect 65 41 66 42
rect 64 41 65 42
rect 34 41 35 42
rect 33 41 34 42
rect 32 41 33 42
rect 31 41 32 42
rect 30 41 31 42
rect 29 41 30 42
rect 28 41 29 42
rect 27 41 28 42
rect 26 41 27 42
rect 25 41 26 42
rect 24 41 25 42
rect 23 41 24 42
rect 22 41 23 42
rect 21 41 22 42
rect 20 41 21 42
rect 19 41 20 42
rect 18 41 19 42
rect 17 41 18 42
rect 16 41 17 42
rect 144 42 145 43
rect 143 42 144 43
rect 142 42 143 43
rect 141 42 142 43
rect 140 42 141 43
rect 135 42 136 43
rect 134 42 135 43
rect 133 42 134 43
rect 132 42 133 43
rect 131 42 132 43
rect 130 42 131 43
rect 123 42 124 43
rect 122 42 123 43
rect 121 42 122 43
rect 120 42 121 43
rect 119 42 120 43
rect 83 42 84 43
rect 82 42 83 43
rect 81 42 82 43
rect 80 42 81 43
rect 79 42 80 43
rect 78 42 79 43
rect 77 42 78 43
rect 76 42 77 43
rect 75 42 76 43
rect 74 42 75 43
rect 73 42 74 43
rect 72 42 73 43
rect 71 42 72 43
rect 70 42 71 43
rect 69 42 70 43
rect 68 42 69 43
rect 67 42 68 43
rect 66 42 67 43
rect 65 42 66 43
rect 64 42 65 43
rect 34 42 35 43
rect 33 42 34 43
rect 32 42 33 43
rect 31 42 32 43
rect 30 42 31 43
rect 29 42 30 43
rect 28 42 29 43
rect 27 42 28 43
rect 26 42 27 43
rect 25 42 26 43
rect 24 42 25 43
rect 23 42 24 43
rect 22 42 23 43
rect 21 42 22 43
rect 20 42 21 43
rect 19 42 20 43
rect 18 42 19 43
rect 17 42 18 43
rect 16 42 17 43
rect 144 43 145 44
rect 143 43 144 44
rect 142 43 143 44
rect 141 43 142 44
rect 140 43 141 44
rect 135 43 136 44
rect 134 43 135 44
rect 133 43 134 44
rect 132 43 133 44
rect 131 43 132 44
rect 130 43 131 44
rect 129 43 130 44
rect 124 43 125 44
rect 123 43 124 44
rect 122 43 123 44
rect 121 43 122 44
rect 120 43 121 44
rect 119 43 120 44
rect 83 43 84 44
rect 82 43 83 44
rect 81 43 82 44
rect 80 43 81 44
rect 79 43 80 44
rect 78 43 79 44
rect 77 43 78 44
rect 76 43 77 44
rect 75 43 76 44
rect 74 43 75 44
rect 73 43 74 44
rect 72 43 73 44
rect 71 43 72 44
rect 70 43 71 44
rect 69 43 70 44
rect 68 43 69 44
rect 67 43 68 44
rect 66 43 67 44
rect 65 43 66 44
rect 33 43 34 44
rect 32 43 33 44
rect 31 43 32 44
rect 30 43 31 44
rect 29 43 30 44
rect 28 43 29 44
rect 27 43 28 44
rect 26 43 27 44
rect 25 43 26 44
rect 24 43 25 44
rect 23 43 24 44
rect 22 43 23 44
rect 21 43 22 44
rect 20 43 21 44
rect 19 43 20 44
rect 18 43 19 44
rect 17 43 18 44
rect 16 43 17 44
rect 144 44 145 45
rect 143 44 144 45
rect 142 44 143 45
rect 141 44 142 45
rect 140 44 141 45
rect 134 44 135 45
rect 133 44 134 45
rect 132 44 133 45
rect 131 44 132 45
rect 130 44 131 45
rect 129 44 130 45
rect 128 44 129 45
rect 127 44 128 45
rect 126 44 127 45
rect 125 44 126 45
rect 124 44 125 45
rect 123 44 124 45
rect 122 44 123 45
rect 121 44 122 45
rect 120 44 121 45
rect 119 44 120 45
rect 83 44 84 45
rect 82 44 83 45
rect 81 44 82 45
rect 80 44 81 45
rect 79 44 80 45
rect 78 44 79 45
rect 77 44 78 45
rect 76 44 77 45
rect 75 44 76 45
rect 74 44 75 45
rect 73 44 74 45
rect 72 44 73 45
rect 71 44 72 45
rect 70 44 71 45
rect 69 44 70 45
rect 68 44 69 45
rect 67 44 68 45
rect 66 44 67 45
rect 65 44 66 45
rect 33 44 34 45
rect 32 44 33 45
rect 31 44 32 45
rect 30 44 31 45
rect 29 44 30 45
rect 28 44 29 45
rect 27 44 28 45
rect 26 44 27 45
rect 25 44 26 45
rect 24 44 25 45
rect 23 44 24 45
rect 22 44 23 45
rect 21 44 22 45
rect 20 44 21 45
rect 19 44 20 45
rect 18 44 19 45
rect 17 44 18 45
rect 16 44 17 45
rect 15 44 16 45
rect 144 45 145 46
rect 143 45 144 46
rect 142 45 143 46
rect 141 45 142 46
rect 140 45 141 46
rect 133 45 134 46
rect 132 45 133 46
rect 131 45 132 46
rect 130 45 131 46
rect 129 45 130 46
rect 128 45 129 46
rect 127 45 128 46
rect 126 45 127 46
rect 125 45 126 46
rect 124 45 125 46
rect 123 45 124 46
rect 122 45 123 46
rect 121 45 122 46
rect 120 45 121 46
rect 83 45 84 46
rect 82 45 83 46
rect 81 45 82 46
rect 80 45 81 46
rect 79 45 80 46
rect 78 45 79 46
rect 77 45 78 46
rect 76 45 77 46
rect 75 45 76 46
rect 74 45 75 46
rect 73 45 74 46
rect 72 45 73 46
rect 71 45 72 46
rect 70 45 71 46
rect 69 45 70 46
rect 68 45 69 46
rect 67 45 68 46
rect 66 45 67 46
rect 32 45 33 46
rect 31 45 32 46
rect 30 45 31 46
rect 29 45 30 46
rect 28 45 29 46
rect 27 45 28 46
rect 26 45 27 46
rect 25 45 26 46
rect 24 45 25 46
rect 23 45 24 46
rect 22 45 23 46
rect 21 45 22 46
rect 20 45 21 46
rect 19 45 20 46
rect 18 45 19 46
rect 17 45 18 46
rect 16 45 17 46
rect 15 45 16 46
rect 144 46 145 47
rect 143 46 144 47
rect 142 46 143 47
rect 141 46 142 47
rect 140 46 141 47
rect 132 46 133 47
rect 131 46 132 47
rect 130 46 131 47
rect 129 46 130 47
rect 128 46 129 47
rect 127 46 128 47
rect 126 46 127 47
rect 125 46 126 47
rect 124 46 125 47
rect 123 46 124 47
rect 122 46 123 47
rect 121 46 122 47
rect 120 46 121 47
rect 83 46 84 47
rect 82 46 83 47
rect 81 46 82 47
rect 80 46 81 47
rect 79 46 80 47
rect 78 46 79 47
rect 77 46 78 47
rect 76 46 77 47
rect 75 46 76 47
rect 74 46 75 47
rect 73 46 74 47
rect 72 46 73 47
rect 71 46 72 47
rect 70 46 71 47
rect 69 46 70 47
rect 68 46 69 47
rect 67 46 68 47
rect 66 46 67 47
rect 32 46 33 47
rect 31 46 32 47
rect 30 46 31 47
rect 29 46 30 47
rect 28 46 29 47
rect 27 46 28 47
rect 26 46 27 47
rect 25 46 26 47
rect 24 46 25 47
rect 23 46 24 47
rect 22 46 23 47
rect 21 46 22 47
rect 20 46 21 47
rect 19 46 20 47
rect 18 46 19 47
rect 17 46 18 47
rect 16 46 17 47
rect 15 46 16 47
rect 144 47 145 48
rect 143 47 144 48
rect 142 47 143 48
rect 141 47 142 48
rect 140 47 141 48
rect 131 47 132 48
rect 130 47 131 48
rect 129 47 130 48
rect 128 47 129 48
rect 127 47 128 48
rect 126 47 127 48
rect 125 47 126 48
rect 124 47 125 48
rect 123 47 124 48
rect 122 47 123 48
rect 121 47 122 48
rect 83 47 84 48
rect 82 47 83 48
rect 81 47 82 48
rect 80 47 81 48
rect 79 47 80 48
rect 78 47 79 48
rect 77 47 78 48
rect 76 47 77 48
rect 75 47 76 48
rect 74 47 75 48
rect 73 47 74 48
rect 72 47 73 48
rect 71 47 72 48
rect 70 47 71 48
rect 69 47 70 48
rect 68 47 69 48
rect 67 47 68 48
rect 66 47 67 48
rect 32 47 33 48
rect 31 47 32 48
rect 30 47 31 48
rect 29 47 30 48
rect 28 47 29 48
rect 27 47 28 48
rect 26 47 27 48
rect 25 47 26 48
rect 24 47 25 48
rect 23 47 24 48
rect 22 47 23 48
rect 21 47 22 48
rect 20 47 21 48
rect 19 47 20 48
rect 18 47 19 48
rect 17 47 18 48
rect 16 47 17 48
rect 15 47 16 48
rect 144 48 145 49
rect 143 48 144 49
rect 142 48 143 49
rect 141 48 142 49
rect 140 48 141 49
rect 130 48 131 49
rect 129 48 130 49
rect 128 48 129 49
rect 127 48 128 49
rect 126 48 127 49
rect 125 48 126 49
rect 124 48 125 49
rect 123 48 124 49
rect 122 48 123 49
rect 83 48 84 49
rect 82 48 83 49
rect 81 48 82 49
rect 80 48 81 49
rect 79 48 80 49
rect 78 48 79 49
rect 77 48 78 49
rect 76 48 77 49
rect 75 48 76 49
rect 74 48 75 49
rect 73 48 74 49
rect 72 48 73 49
rect 71 48 72 49
rect 70 48 71 49
rect 69 48 70 49
rect 68 48 69 49
rect 67 48 68 49
rect 31 48 32 49
rect 30 48 31 49
rect 29 48 30 49
rect 28 48 29 49
rect 27 48 28 49
rect 26 48 27 49
rect 25 48 26 49
rect 24 48 25 49
rect 23 48 24 49
rect 22 48 23 49
rect 21 48 22 49
rect 20 48 21 49
rect 19 48 20 49
rect 18 48 19 49
rect 17 48 18 49
rect 16 48 17 49
rect 15 48 16 49
rect 144 49 145 50
rect 143 49 144 50
rect 142 49 143 50
rect 141 49 142 50
rect 140 49 141 50
rect 127 49 128 50
rect 126 49 127 50
rect 125 49 126 50
rect 83 49 84 50
rect 82 49 83 50
rect 81 49 82 50
rect 80 49 81 50
rect 79 49 80 50
rect 78 49 79 50
rect 77 49 78 50
rect 76 49 77 50
rect 75 49 76 50
rect 74 49 75 50
rect 73 49 74 50
rect 72 49 73 50
rect 71 49 72 50
rect 70 49 71 50
rect 69 49 70 50
rect 68 49 69 50
rect 67 49 68 50
rect 31 49 32 50
rect 30 49 31 50
rect 29 49 30 50
rect 28 49 29 50
rect 27 49 28 50
rect 26 49 27 50
rect 25 49 26 50
rect 24 49 25 50
rect 23 49 24 50
rect 22 49 23 50
rect 21 49 22 50
rect 20 49 21 50
rect 19 49 20 50
rect 18 49 19 50
rect 17 49 18 50
rect 16 49 17 50
rect 15 49 16 50
rect 83 50 84 51
rect 82 50 83 51
rect 81 50 82 51
rect 80 50 81 51
rect 79 50 80 51
rect 78 50 79 51
rect 77 50 78 51
rect 76 50 77 51
rect 75 50 76 51
rect 74 50 75 51
rect 73 50 74 51
rect 72 50 73 51
rect 71 50 72 51
rect 70 50 71 51
rect 69 50 70 51
rect 68 50 69 51
rect 67 50 68 51
rect 31 50 32 51
rect 30 50 31 51
rect 29 50 30 51
rect 28 50 29 51
rect 27 50 28 51
rect 26 50 27 51
rect 25 50 26 51
rect 24 50 25 51
rect 23 50 24 51
rect 22 50 23 51
rect 21 50 22 51
rect 20 50 21 51
rect 19 50 20 51
rect 18 50 19 51
rect 17 50 18 51
rect 16 50 17 51
rect 15 50 16 51
rect 83 51 84 52
rect 82 51 83 52
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 78 51 79 52
rect 77 51 78 52
rect 76 51 77 52
rect 75 51 76 52
rect 74 51 75 52
rect 73 51 74 52
rect 72 51 73 52
rect 71 51 72 52
rect 70 51 71 52
rect 69 51 70 52
rect 68 51 69 52
rect 67 51 68 52
rect 31 51 32 52
rect 30 51 31 52
rect 29 51 30 52
rect 28 51 29 52
rect 27 51 28 52
rect 26 51 27 52
rect 25 51 26 52
rect 24 51 25 52
rect 23 51 24 52
rect 22 51 23 52
rect 21 51 22 52
rect 20 51 21 52
rect 19 51 20 52
rect 18 51 19 52
rect 17 51 18 52
rect 16 51 17 52
rect 15 51 16 52
rect 83 52 84 53
rect 82 52 83 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 77 52 78 53
rect 76 52 77 53
rect 75 52 76 53
rect 74 52 75 53
rect 73 52 74 53
rect 72 52 73 53
rect 71 52 72 53
rect 70 52 71 53
rect 69 52 70 53
rect 68 52 69 53
rect 67 52 68 53
rect 31 52 32 53
rect 30 52 31 53
rect 29 52 30 53
rect 28 52 29 53
rect 27 52 28 53
rect 26 52 27 53
rect 25 52 26 53
rect 24 52 25 53
rect 23 52 24 53
rect 22 52 23 53
rect 21 52 22 53
rect 20 52 21 53
rect 19 52 20 53
rect 18 52 19 53
rect 17 52 18 53
rect 16 52 17 53
rect 15 52 16 53
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 76 53 77 54
rect 75 53 76 54
rect 74 53 75 54
rect 73 53 74 54
rect 72 53 73 54
rect 71 53 72 54
rect 70 53 71 54
rect 69 53 70 54
rect 68 53 69 54
rect 67 53 68 54
rect 31 53 32 54
rect 30 53 31 54
rect 29 53 30 54
rect 28 53 29 54
rect 27 53 28 54
rect 26 53 27 54
rect 25 53 26 54
rect 24 53 25 54
rect 23 53 24 54
rect 22 53 23 54
rect 21 53 22 54
rect 20 53 21 54
rect 19 53 20 54
rect 18 53 19 54
rect 17 53 18 54
rect 16 53 17 54
rect 15 53 16 54
rect 137 54 138 55
rect 136 54 137 55
rect 135 54 136 55
rect 134 54 135 55
rect 133 54 134 55
rect 132 54 133 55
rect 131 54 132 55
rect 130 54 131 55
rect 129 54 130 55
rect 128 54 129 55
rect 127 54 128 55
rect 126 54 127 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 75 54 76 55
rect 74 54 75 55
rect 73 54 74 55
rect 72 54 73 55
rect 71 54 72 55
rect 70 54 71 55
rect 69 54 70 55
rect 68 54 69 55
rect 67 54 68 55
rect 31 54 32 55
rect 30 54 31 55
rect 29 54 30 55
rect 28 54 29 55
rect 27 54 28 55
rect 26 54 27 55
rect 25 54 26 55
rect 24 54 25 55
rect 23 54 24 55
rect 22 54 23 55
rect 21 54 22 55
rect 20 54 21 55
rect 19 54 20 55
rect 18 54 19 55
rect 17 54 18 55
rect 16 54 17 55
rect 15 54 16 55
rect 140 55 141 56
rect 139 55 140 56
rect 138 55 139 56
rect 137 55 138 56
rect 136 55 137 56
rect 135 55 136 56
rect 134 55 135 56
rect 133 55 134 56
rect 132 55 133 56
rect 131 55 132 56
rect 130 55 131 56
rect 129 55 130 56
rect 128 55 129 56
rect 127 55 128 56
rect 126 55 127 56
rect 125 55 126 56
rect 124 55 125 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 75 55 76 56
rect 74 55 75 56
rect 73 55 74 56
rect 72 55 73 56
rect 71 55 72 56
rect 70 55 71 56
rect 69 55 70 56
rect 68 55 69 56
rect 67 55 68 56
rect 31 55 32 56
rect 30 55 31 56
rect 29 55 30 56
rect 28 55 29 56
rect 27 55 28 56
rect 26 55 27 56
rect 25 55 26 56
rect 24 55 25 56
rect 23 55 24 56
rect 22 55 23 56
rect 21 55 22 56
rect 20 55 21 56
rect 19 55 20 56
rect 18 55 19 56
rect 17 55 18 56
rect 16 55 17 56
rect 15 55 16 56
rect 141 56 142 57
rect 140 56 141 57
rect 139 56 140 57
rect 138 56 139 57
rect 137 56 138 57
rect 136 56 137 57
rect 135 56 136 57
rect 134 56 135 57
rect 133 56 134 57
rect 132 56 133 57
rect 131 56 132 57
rect 130 56 131 57
rect 129 56 130 57
rect 128 56 129 57
rect 127 56 128 57
rect 126 56 127 57
rect 125 56 126 57
rect 124 56 125 57
rect 123 56 124 57
rect 122 56 123 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 74 56 75 57
rect 73 56 74 57
rect 72 56 73 57
rect 71 56 72 57
rect 70 56 71 57
rect 69 56 70 57
rect 68 56 69 57
rect 67 56 68 57
rect 31 56 32 57
rect 30 56 31 57
rect 29 56 30 57
rect 28 56 29 57
rect 27 56 28 57
rect 26 56 27 57
rect 25 56 26 57
rect 24 56 25 57
rect 23 56 24 57
rect 22 56 23 57
rect 21 56 22 57
rect 20 56 21 57
rect 19 56 20 57
rect 18 56 19 57
rect 17 56 18 57
rect 16 56 17 57
rect 15 56 16 57
rect 142 57 143 58
rect 141 57 142 58
rect 140 57 141 58
rect 139 57 140 58
rect 138 57 139 58
rect 137 57 138 58
rect 136 57 137 58
rect 135 57 136 58
rect 134 57 135 58
rect 133 57 134 58
rect 132 57 133 58
rect 131 57 132 58
rect 130 57 131 58
rect 129 57 130 58
rect 128 57 129 58
rect 127 57 128 58
rect 126 57 127 58
rect 125 57 126 58
rect 124 57 125 58
rect 123 57 124 58
rect 122 57 123 58
rect 121 57 122 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 73 57 74 58
rect 72 57 73 58
rect 71 57 72 58
rect 70 57 71 58
rect 69 57 70 58
rect 68 57 69 58
rect 67 57 68 58
rect 31 57 32 58
rect 30 57 31 58
rect 29 57 30 58
rect 28 57 29 58
rect 27 57 28 58
rect 26 57 27 58
rect 25 57 26 58
rect 24 57 25 58
rect 23 57 24 58
rect 22 57 23 58
rect 21 57 22 58
rect 20 57 21 58
rect 19 57 20 58
rect 18 57 19 58
rect 17 57 18 58
rect 16 57 17 58
rect 15 57 16 58
rect 143 58 144 59
rect 142 58 143 59
rect 141 58 142 59
rect 140 58 141 59
rect 139 58 140 59
rect 138 58 139 59
rect 137 58 138 59
rect 136 58 137 59
rect 135 58 136 59
rect 134 58 135 59
rect 133 58 134 59
rect 132 58 133 59
rect 131 58 132 59
rect 130 58 131 59
rect 129 58 130 59
rect 128 58 129 59
rect 127 58 128 59
rect 126 58 127 59
rect 125 58 126 59
rect 124 58 125 59
rect 123 58 124 59
rect 122 58 123 59
rect 121 58 122 59
rect 120 58 121 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 73 58 74 59
rect 72 58 73 59
rect 71 58 72 59
rect 70 58 71 59
rect 69 58 70 59
rect 68 58 69 59
rect 67 58 68 59
rect 66 58 67 59
rect 31 58 32 59
rect 30 58 31 59
rect 29 58 30 59
rect 28 58 29 59
rect 27 58 28 59
rect 26 58 27 59
rect 25 58 26 59
rect 24 58 25 59
rect 23 58 24 59
rect 22 58 23 59
rect 21 58 22 59
rect 20 58 21 59
rect 19 58 20 59
rect 18 58 19 59
rect 17 58 18 59
rect 16 58 17 59
rect 143 59 144 60
rect 142 59 143 60
rect 141 59 142 60
rect 140 59 141 60
rect 139 59 140 60
rect 138 59 139 60
rect 137 59 138 60
rect 136 59 137 60
rect 135 59 136 60
rect 128 59 129 60
rect 127 59 128 60
rect 126 59 127 60
rect 125 59 126 60
rect 124 59 125 60
rect 123 59 124 60
rect 122 59 123 60
rect 121 59 122 60
rect 120 59 121 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 72 59 73 60
rect 71 59 72 60
rect 70 59 71 60
rect 69 59 70 60
rect 68 59 69 60
rect 67 59 68 60
rect 66 59 67 60
rect 32 59 33 60
rect 31 59 32 60
rect 30 59 31 60
rect 29 59 30 60
rect 28 59 29 60
rect 27 59 28 60
rect 26 59 27 60
rect 25 59 26 60
rect 24 59 25 60
rect 23 59 24 60
rect 22 59 23 60
rect 21 59 22 60
rect 20 59 21 60
rect 19 59 20 60
rect 18 59 19 60
rect 17 59 18 60
rect 16 59 17 60
rect 144 60 145 61
rect 143 60 144 61
rect 142 60 143 61
rect 141 60 142 61
rect 140 60 141 61
rect 139 60 140 61
rect 124 60 125 61
rect 123 60 124 61
rect 122 60 123 61
rect 121 60 122 61
rect 120 60 121 61
rect 119 60 120 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 72 60 73 61
rect 71 60 72 61
rect 70 60 71 61
rect 69 60 70 61
rect 68 60 69 61
rect 67 60 68 61
rect 66 60 67 61
rect 32 60 33 61
rect 31 60 32 61
rect 30 60 31 61
rect 29 60 30 61
rect 28 60 29 61
rect 27 60 28 61
rect 26 60 27 61
rect 25 60 26 61
rect 24 60 25 61
rect 23 60 24 61
rect 22 60 23 61
rect 21 60 22 61
rect 20 60 21 61
rect 19 60 20 61
rect 18 60 19 61
rect 17 60 18 61
rect 16 60 17 61
rect 144 61 145 62
rect 143 61 144 62
rect 142 61 143 62
rect 141 61 142 62
rect 140 61 141 62
rect 123 61 124 62
rect 122 61 123 62
rect 121 61 122 62
rect 120 61 121 62
rect 119 61 120 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 71 61 72 62
rect 70 61 71 62
rect 69 61 70 62
rect 68 61 69 62
rect 67 61 68 62
rect 66 61 67 62
rect 32 61 33 62
rect 31 61 32 62
rect 30 61 31 62
rect 29 61 30 62
rect 28 61 29 62
rect 27 61 28 62
rect 26 61 27 62
rect 25 61 26 62
rect 24 61 25 62
rect 23 61 24 62
rect 22 61 23 62
rect 21 61 22 62
rect 20 61 21 62
rect 19 61 20 62
rect 18 61 19 62
rect 17 61 18 62
rect 16 61 17 62
rect 144 62 145 63
rect 143 62 144 63
rect 142 62 143 63
rect 141 62 142 63
rect 122 62 123 63
rect 121 62 122 63
rect 120 62 121 63
rect 119 62 120 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 71 62 72 63
rect 70 62 71 63
rect 69 62 70 63
rect 68 62 69 63
rect 67 62 68 63
rect 66 62 67 63
rect 65 62 66 63
rect 33 62 34 63
rect 32 62 33 63
rect 31 62 32 63
rect 30 62 31 63
rect 29 62 30 63
rect 28 62 29 63
rect 27 62 28 63
rect 26 62 27 63
rect 25 62 26 63
rect 24 62 25 63
rect 23 62 24 63
rect 22 62 23 63
rect 21 62 22 63
rect 20 62 21 63
rect 19 62 20 63
rect 18 62 19 63
rect 17 62 18 63
rect 16 62 17 63
rect 144 63 145 64
rect 143 63 144 64
rect 142 63 143 64
rect 141 63 142 64
rect 122 63 123 64
rect 121 63 122 64
rect 120 63 121 64
rect 119 63 120 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 70 63 71 64
rect 69 63 70 64
rect 68 63 69 64
rect 67 63 68 64
rect 66 63 67 64
rect 65 63 66 64
rect 33 63 34 64
rect 32 63 33 64
rect 31 63 32 64
rect 30 63 31 64
rect 29 63 30 64
rect 28 63 29 64
rect 27 63 28 64
rect 26 63 27 64
rect 25 63 26 64
rect 24 63 25 64
rect 23 63 24 64
rect 22 63 23 64
rect 21 63 22 64
rect 20 63 21 64
rect 19 63 20 64
rect 18 63 19 64
rect 17 63 18 64
rect 16 63 17 64
rect 144 64 145 65
rect 143 64 144 65
rect 142 64 143 65
rect 141 64 142 65
rect 140 64 141 65
rect 123 64 124 65
rect 122 64 123 65
rect 121 64 122 65
rect 120 64 121 65
rect 119 64 120 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 70 64 71 65
rect 69 64 70 65
rect 68 64 69 65
rect 67 64 68 65
rect 66 64 67 65
rect 65 64 66 65
rect 33 64 34 65
rect 32 64 33 65
rect 31 64 32 65
rect 30 64 31 65
rect 29 64 30 65
rect 28 64 29 65
rect 27 64 28 65
rect 26 64 27 65
rect 25 64 26 65
rect 24 64 25 65
rect 23 64 24 65
rect 22 64 23 65
rect 21 64 22 65
rect 20 64 21 65
rect 19 64 20 65
rect 18 64 19 65
rect 17 64 18 65
rect 16 64 17 65
rect 144 65 145 66
rect 143 65 144 66
rect 142 65 143 66
rect 141 65 142 66
rect 140 65 141 66
rect 139 65 140 66
rect 124 65 125 66
rect 123 65 124 66
rect 122 65 123 66
rect 121 65 122 66
rect 120 65 121 66
rect 119 65 120 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 69 65 70 66
rect 68 65 69 66
rect 67 65 68 66
rect 66 65 67 66
rect 65 65 66 66
rect 64 65 65 66
rect 34 65 35 66
rect 33 65 34 66
rect 32 65 33 66
rect 31 65 32 66
rect 30 65 31 66
rect 29 65 30 66
rect 28 65 29 66
rect 27 65 28 66
rect 26 65 27 66
rect 25 65 26 66
rect 24 65 25 66
rect 23 65 24 66
rect 22 65 23 66
rect 21 65 22 66
rect 20 65 21 66
rect 19 65 20 66
rect 18 65 19 66
rect 17 65 18 66
rect 143 66 144 67
rect 142 66 143 67
rect 141 66 142 67
rect 140 66 141 67
rect 139 66 140 67
rect 138 66 139 67
rect 137 66 138 67
rect 136 66 137 67
rect 127 66 128 67
rect 126 66 127 67
rect 125 66 126 67
rect 124 66 125 67
rect 123 66 124 67
rect 122 66 123 67
rect 121 66 122 67
rect 120 66 121 67
rect 119 66 120 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 71 66 72 67
rect 70 66 71 67
rect 69 66 70 67
rect 68 66 69 67
rect 67 66 68 67
rect 66 66 67 67
rect 65 66 66 67
rect 64 66 65 67
rect 34 66 35 67
rect 33 66 34 67
rect 32 66 33 67
rect 31 66 32 67
rect 30 66 31 67
rect 29 66 30 67
rect 28 66 29 67
rect 27 66 28 67
rect 26 66 27 67
rect 25 66 26 67
rect 24 66 25 67
rect 23 66 24 67
rect 22 66 23 67
rect 21 66 22 67
rect 20 66 21 67
rect 19 66 20 67
rect 18 66 19 67
rect 17 66 18 67
rect 143 67 144 68
rect 142 67 143 68
rect 141 67 142 68
rect 140 67 141 68
rect 139 67 140 68
rect 138 67 139 68
rect 137 67 138 68
rect 136 67 137 68
rect 135 67 136 68
rect 134 67 135 68
rect 133 67 134 68
rect 132 67 133 68
rect 131 67 132 68
rect 130 67 131 68
rect 129 67 130 68
rect 128 67 129 68
rect 127 67 128 68
rect 126 67 127 68
rect 125 67 126 68
rect 124 67 125 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 120 67 121 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 71 67 72 68
rect 70 67 71 68
rect 69 67 70 68
rect 68 67 69 68
rect 67 67 68 68
rect 66 67 67 68
rect 65 67 66 68
rect 64 67 65 68
rect 63 67 64 68
rect 35 67 36 68
rect 34 67 35 68
rect 33 67 34 68
rect 32 67 33 68
rect 31 67 32 68
rect 30 67 31 68
rect 29 67 30 68
rect 28 67 29 68
rect 27 67 28 68
rect 26 67 27 68
rect 25 67 26 68
rect 24 67 25 68
rect 23 67 24 68
rect 22 67 23 68
rect 21 67 22 68
rect 20 67 21 68
rect 19 67 20 68
rect 18 67 19 68
rect 17 67 18 68
rect 142 68 143 69
rect 141 68 142 69
rect 140 68 141 69
rect 139 68 140 69
rect 138 68 139 69
rect 137 68 138 69
rect 136 68 137 69
rect 135 68 136 69
rect 134 68 135 69
rect 133 68 134 69
rect 132 68 133 69
rect 131 68 132 69
rect 130 68 131 69
rect 129 68 130 69
rect 128 68 129 69
rect 127 68 128 69
rect 126 68 127 69
rect 125 68 126 69
rect 124 68 125 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 120 68 121 69
rect 141 69 142 70
rect 140 69 141 70
rect 139 69 140 70
rect 138 69 139 70
rect 137 69 138 70
rect 136 69 137 70
rect 135 69 136 70
rect 134 69 135 70
rect 133 69 134 70
rect 132 69 133 70
rect 131 69 132 70
rect 130 69 131 70
rect 129 69 130 70
rect 128 69 129 70
rect 127 69 128 70
rect 126 69 127 70
rect 125 69 126 70
rect 124 69 125 70
rect 123 69 124 70
rect 122 69 123 70
rect 121 69 122 70
rect 140 70 141 71
rect 139 70 140 71
rect 138 70 139 71
rect 137 70 138 71
rect 136 70 137 71
rect 135 70 136 71
rect 134 70 135 71
rect 133 70 134 71
rect 132 70 133 71
rect 131 70 132 71
rect 130 70 131 71
rect 129 70 130 71
rect 128 70 129 71
rect 127 70 128 71
rect 126 70 127 71
rect 125 70 126 71
rect 124 70 125 71
rect 123 70 124 71
rect 138 71 139 72
rect 137 71 138 72
rect 136 71 137 72
rect 135 71 136 72
rect 134 71 135 72
rect 133 71 134 72
rect 132 71 133 72
rect 131 71 132 72
rect 130 71 131 72
rect 129 71 130 72
rect 128 71 129 72
rect 127 71 128 72
rect 126 71 127 72
rect 125 71 126 72
rect 144 76 145 77
rect 143 76 144 77
rect 142 76 143 77
rect 141 76 142 77
rect 140 76 141 77
rect 139 76 140 77
rect 144 77 145 78
rect 143 77 144 78
rect 142 77 143 78
rect 141 77 142 78
rect 140 77 141 78
rect 139 77 140 78
rect 138 77 139 78
rect 137 77 138 78
rect 124 77 125 78
rect 123 77 124 78
rect 122 77 123 78
rect 121 77 122 78
rect 144 78 145 79
rect 143 78 144 79
rect 142 78 143 79
rect 141 78 142 79
rect 140 78 141 79
rect 139 78 140 79
rect 138 78 139 79
rect 137 78 138 79
rect 136 78 137 79
rect 124 78 125 79
rect 123 78 124 79
rect 122 78 123 79
rect 121 78 122 79
rect 120 78 121 79
rect 82 78 83 79
rect 81 78 82 79
rect 80 78 81 79
rect 79 78 80 79
rect 78 78 79 79
rect 77 78 78 79
rect 76 78 77 79
rect 75 78 76 79
rect 74 78 75 79
rect 73 78 74 79
rect 72 78 73 79
rect 71 78 72 79
rect 70 78 71 79
rect 69 78 70 79
rect 68 78 69 79
rect 67 78 68 79
rect 66 78 67 79
rect 65 78 66 79
rect 64 78 65 79
rect 63 78 64 79
rect 62 78 63 79
rect 61 78 62 79
rect 60 78 61 79
rect 59 78 60 79
rect 58 78 59 79
rect 57 78 58 79
rect 56 78 57 79
rect 55 78 56 79
rect 54 78 55 79
rect 53 78 54 79
rect 52 78 53 79
rect 51 78 52 79
rect 50 78 51 79
rect 49 78 50 79
rect 48 78 49 79
rect 47 78 48 79
rect 46 78 47 79
rect 45 78 46 79
rect 44 78 45 79
rect 43 78 44 79
rect 42 78 43 79
rect 41 78 42 79
rect 40 78 41 79
rect 39 78 40 79
rect 38 78 39 79
rect 37 78 38 79
rect 36 78 37 79
rect 35 78 36 79
rect 34 78 35 79
rect 33 78 34 79
rect 32 78 33 79
rect 31 78 32 79
rect 30 78 31 79
rect 29 78 30 79
rect 28 78 29 79
rect 27 78 28 79
rect 26 78 27 79
rect 25 78 26 79
rect 24 78 25 79
rect 23 78 24 79
rect 22 78 23 79
rect 21 78 22 79
rect 20 78 21 79
rect 19 78 20 79
rect 18 78 19 79
rect 17 78 18 79
rect 16 78 17 79
rect 144 79 145 80
rect 143 79 144 80
rect 142 79 143 80
rect 141 79 142 80
rect 140 79 141 80
rect 139 79 140 80
rect 138 79 139 80
rect 137 79 138 80
rect 136 79 137 80
rect 135 79 136 80
rect 123 79 124 80
rect 122 79 123 80
rect 121 79 122 80
rect 120 79 121 80
rect 82 79 83 80
rect 81 79 82 80
rect 80 79 81 80
rect 79 79 80 80
rect 78 79 79 80
rect 77 79 78 80
rect 76 79 77 80
rect 75 79 76 80
rect 74 79 75 80
rect 73 79 74 80
rect 72 79 73 80
rect 71 79 72 80
rect 70 79 71 80
rect 69 79 70 80
rect 68 79 69 80
rect 67 79 68 80
rect 66 79 67 80
rect 65 79 66 80
rect 64 79 65 80
rect 63 79 64 80
rect 62 79 63 80
rect 61 79 62 80
rect 60 79 61 80
rect 59 79 60 80
rect 58 79 59 80
rect 57 79 58 80
rect 56 79 57 80
rect 55 79 56 80
rect 54 79 55 80
rect 53 79 54 80
rect 52 79 53 80
rect 51 79 52 80
rect 50 79 51 80
rect 49 79 50 80
rect 48 79 49 80
rect 47 79 48 80
rect 46 79 47 80
rect 45 79 46 80
rect 44 79 45 80
rect 43 79 44 80
rect 42 79 43 80
rect 41 79 42 80
rect 40 79 41 80
rect 39 79 40 80
rect 38 79 39 80
rect 37 79 38 80
rect 36 79 37 80
rect 35 79 36 80
rect 34 79 35 80
rect 33 79 34 80
rect 32 79 33 80
rect 31 79 32 80
rect 30 79 31 80
rect 29 79 30 80
rect 28 79 29 80
rect 27 79 28 80
rect 26 79 27 80
rect 25 79 26 80
rect 24 79 25 80
rect 23 79 24 80
rect 22 79 23 80
rect 21 79 22 80
rect 20 79 21 80
rect 19 79 20 80
rect 18 79 19 80
rect 17 79 18 80
rect 16 79 17 80
rect 144 80 145 81
rect 143 80 144 81
rect 142 80 143 81
rect 141 80 142 81
rect 140 80 141 81
rect 139 80 140 81
rect 138 80 139 81
rect 137 80 138 81
rect 136 80 137 81
rect 135 80 136 81
rect 134 80 135 81
rect 123 80 124 81
rect 122 80 123 81
rect 121 80 122 81
rect 120 80 121 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 61 80 62 81
rect 60 80 61 81
rect 59 80 60 81
rect 58 80 59 81
rect 57 80 58 81
rect 56 80 57 81
rect 55 80 56 81
rect 54 80 55 81
rect 53 80 54 81
rect 52 80 53 81
rect 51 80 52 81
rect 50 80 51 81
rect 49 80 50 81
rect 48 80 49 81
rect 47 80 48 81
rect 46 80 47 81
rect 45 80 46 81
rect 44 80 45 81
rect 43 80 44 81
rect 42 80 43 81
rect 41 80 42 81
rect 40 80 41 81
rect 39 80 40 81
rect 38 80 39 81
rect 37 80 38 81
rect 36 80 37 81
rect 35 80 36 81
rect 34 80 35 81
rect 33 80 34 81
rect 32 80 33 81
rect 31 80 32 81
rect 30 80 31 81
rect 29 80 30 81
rect 28 80 29 81
rect 27 80 28 81
rect 26 80 27 81
rect 25 80 26 81
rect 24 80 25 81
rect 23 80 24 81
rect 22 80 23 81
rect 21 80 22 81
rect 20 80 21 81
rect 19 80 20 81
rect 18 80 19 81
rect 17 80 18 81
rect 16 80 17 81
rect 144 81 145 82
rect 143 81 144 82
rect 142 81 143 82
rect 141 81 142 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 136 81 137 82
rect 135 81 136 82
rect 134 81 135 82
rect 123 81 124 82
rect 122 81 123 82
rect 121 81 122 82
rect 120 81 121 82
rect 119 81 120 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 61 81 62 82
rect 60 81 61 82
rect 59 81 60 82
rect 58 81 59 82
rect 57 81 58 82
rect 56 81 57 82
rect 55 81 56 82
rect 54 81 55 82
rect 53 81 54 82
rect 52 81 53 82
rect 51 81 52 82
rect 50 81 51 82
rect 49 81 50 82
rect 48 81 49 82
rect 47 81 48 82
rect 46 81 47 82
rect 45 81 46 82
rect 44 81 45 82
rect 43 81 44 82
rect 42 81 43 82
rect 41 81 42 82
rect 40 81 41 82
rect 39 81 40 82
rect 38 81 39 82
rect 37 81 38 82
rect 36 81 37 82
rect 35 81 36 82
rect 34 81 35 82
rect 33 81 34 82
rect 32 81 33 82
rect 31 81 32 82
rect 30 81 31 82
rect 29 81 30 82
rect 28 81 29 82
rect 27 81 28 82
rect 26 81 27 82
rect 25 81 26 82
rect 24 81 25 82
rect 23 81 24 82
rect 22 81 23 82
rect 21 81 22 82
rect 20 81 21 82
rect 19 81 20 82
rect 18 81 19 82
rect 17 81 18 82
rect 16 81 17 82
rect 144 82 145 83
rect 143 82 144 83
rect 142 82 143 83
rect 141 82 142 83
rect 140 82 141 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 135 82 136 83
rect 134 82 135 83
rect 133 82 134 83
rect 122 82 123 83
rect 121 82 122 83
rect 120 82 121 83
rect 119 82 120 83
rect 82 82 83 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 60 82 61 83
rect 59 82 60 83
rect 58 82 59 83
rect 57 82 58 83
rect 56 82 57 83
rect 55 82 56 83
rect 54 82 55 83
rect 53 82 54 83
rect 52 82 53 83
rect 51 82 52 83
rect 50 82 51 83
rect 49 82 50 83
rect 48 82 49 83
rect 47 82 48 83
rect 46 82 47 83
rect 45 82 46 83
rect 44 82 45 83
rect 43 82 44 83
rect 42 82 43 83
rect 41 82 42 83
rect 40 82 41 83
rect 39 82 40 83
rect 38 82 39 83
rect 37 82 38 83
rect 36 82 37 83
rect 35 82 36 83
rect 34 82 35 83
rect 33 82 34 83
rect 32 82 33 83
rect 31 82 32 83
rect 30 82 31 83
rect 29 82 30 83
rect 28 82 29 83
rect 27 82 28 83
rect 26 82 27 83
rect 25 82 26 83
rect 24 82 25 83
rect 23 82 24 83
rect 22 82 23 83
rect 21 82 22 83
rect 20 82 21 83
rect 19 82 20 83
rect 18 82 19 83
rect 17 82 18 83
rect 16 82 17 83
rect 144 83 145 84
rect 143 83 144 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 137 83 138 84
rect 136 83 137 84
rect 135 83 136 84
rect 134 83 135 84
rect 133 83 134 84
rect 132 83 133 84
rect 122 83 123 84
rect 121 83 122 84
rect 120 83 121 84
rect 119 83 120 84
rect 82 83 83 84
rect 81 83 82 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 59 83 60 84
rect 58 83 59 84
rect 57 83 58 84
rect 56 83 57 84
rect 55 83 56 84
rect 54 83 55 84
rect 53 83 54 84
rect 52 83 53 84
rect 51 83 52 84
rect 50 83 51 84
rect 49 83 50 84
rect 48 83 49 84
rect 47 83 48 84
rect 46 83 47 84
rect 45 83 46 84
rect 44 83 45 84
rect 43 83 44 84
rect 42 83 43 84
rect 41 83 42 84
rect 40 83 41 84
rect 39 83 40 84
rect 38 83 39 84
rect 37 83 38 84
rect 36 83 37 84
rect 35 83 36 84
rect 34 83 35 84
rect 33 83 34 84
rect 32 83 33 84
rect 31 83 32 84
rect 30 83 31 84
rect 29 83 30 84
rect 28 83 29 84
rect 27 83 28 84
rect 26 83 27 84
rect 25 83 26 84
rect 24 83 25 84
rect 23 83 24 84
rect 22 83 23 84
rect 21 83 22 84
rect 20 83 21 84
rect 19 83 20 84
rect 18 83 19 84
rect 17 83 18 84
rect 16 83 17 84
rect 144 84 145 85
rect 143 84 144 85
rect 142 84 143 85
rect 141 84 142 85
rect 140 84 141 85
rect 136 84 137 85
rect 135 84 136 85
rect 134 84 135 85
rect 133 84 134 85
rect 132 84 133 85
rect 131 84 132 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 120 84 121 85
rect 119 84 120 85
rect 82 84 83 85
rect 81 84 82 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 59 84 60 85
rect 58 84 59 85
rect 57 84 58 85
rect 56 84 57 85
rect 55 84 56 85
rect 54 84 55 85
rect 53 84 54 85
rect 52 84 53 85
rect 51 84 52 85
rect 50 84 51 85
rect 49 84 50 85
rect 48 84 49 85
rect 47 84 48 85
rect 46 84 47 85
rect 45 84 46 85
rect 44 84 45 85
rect 43 84 44 85
rect 42 84 43 85
rect 41 84 42 85
rect 40 84 41 85
rect 39 84 40 85
rect 38 84 39 85
rect 37 84 38 85
rect 36 84 37 85
rect 35 84 36 85
rect 34 84 35 85
rect 33 84 34 85
rect 32 84 33 85
rect 31 84 32 85
rect 30 84 31 85
rect 29 84 30 85
rect 28 84 29 85
rect 27 84 28 85
rect 26 84 27 85
rect 25 84 26 85
rect 24 84 25 85
rect 23 84 24 85
rect 22 84 23 85
rect 21 84 22 85
rect 20 84 21 85
rect 19 84 20 85
rect 18 84 19 85
rect 17 84 18 85
rect 16 84 17 85
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 141 85 142 86
rect 140 85 141 86
rect 135 85 136 86
rect 134 85 135 86
rect 133 85 134 86
rect 132 85 133 86
rect 131 85 132 86
rect 130 85 131 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 120 85 121 86
rect 119 85 120 86
rect 82 85 83 86
rect 81 85 82 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 58 85 59 86
rect 57 85 58 86
rect 56 85 57 86
rect 55 85 56 86
rect 54 85 55 86
rect 53 85 54 86
rect 52 85 53 86
rect 51 85 52 86
rect 50 85 51 86
rect 49 85 50 86
rect 48 85 49 86
rect 47 85 48 86
rect 46 85 47 86
rect 45 85 46 86
rect 44 85 45 86
rect 43 85 44 86
rect 42 85 43 86
rect 41 85 42 86
rect 40 85 41 86
rect 39 85 40 86
rect 38 85 39 86
rect 37 85 38 86
rect 36 85 37 86
rect 35 85 36 86
rect 34 85 35 86
rect 33 85 34 86
rect 32 85 33 86
rect 31 85 32 86
rect 30 85 31 86
rect 29 85 30 86
rect 28 85 29 86
rect 27 85 28 86
rect 26 85 27 86
rect 25 85 26 86
rect 24 85 25 86
rect 23 85 24 86
rect 22 85 23 86
rect 21 85 22 86
rect 20 85 21 86
rect 19 85 20 86
rect 18 85 19 86
rect 17 85 18 86
rect 16 85 17 86
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 141 86 142 87
rect 140 86 141 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 132 86 133 87
rect 131 86 132 87
rect 130 86 131 87
rect 129 86 130 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 120 86 121 87
rect 119 86 120 87
rect 82 86 83 87
rect 81 86 82 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 57 86 58 87
rect 56 86 57 87
rect 55 86 56 87
rect 54 86 55 87
rect 53 86 54 87
rect 52 86 53 87
rect 51 86 52 87
rect 50 86 51 87
rect 49 86 50 87
rect 48 86 49 87
rect 47 86 48 87
rect 46 86 47 87
rect 45 86 46 87
rect 44 86 45 87
rect 43 86 44 87
rect 42 86 43 87
rect 41 86 42 87
rect 40 86 41 87
rect 39 86 40 87
rect 38 86 39 87
rect 37 86 38 87
rect 36 86 37 87
rect 35 86 36 87
rect 34 86 35 87
rect 33 86 34 87
rect 32 86 33 87
rect 31 86 32 87
rect 30 86 31 87
rect 29 86 30 87
rect 28 86 29 87
rect 27 86 28 87
rect 26 86 27 87
rect 25 86 26 87
rect 24 86 25 87
rect 23 86 24 87
rect 22 86 23 87
rect 21 86 22 87
rect 20 86 21 87
rect 19 86 20 87
rect 18 86 19 87
rect 17 86 18 87
rect 16 86 17 87
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 141 87 142 88
rect 140 87 141 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 131 87 132 88
rect 130 87 131 88
rect 129 87 130 88
rect 128 87 129 88
rect 127 87 128 88
rect 126 87 127 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 120 87 121 88
rect 119 87 120 88
rect 82 87 83 88
rect 81 87 82 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 57 87 58 88
rect 56 87 57 88
rect 55 87 56 88
rect 54 87 55 88
rect 53 87 54 88
rect 52 87 53 88
rect 51 87 52 88
rect 50 87 51 88
rect 49 87 50 88
rect 48 87 49 88
rect 47 87 48 88
rect 46 87 47 88
rect 45 87 46 88
rect 44 87 45 88
rect 43 87 44 88
rect 42 87 43 88
rect 41 87 42 88
rect 40 87 41 88
rect 39 87 40 88
rect 38 87 39 88
rect 37 87 38 88
rect 36 87 37 88
rect 35 87 36 88
rect 34 87 35 88
rect 33 87 34 88
rect 32 87 33 88
rect 31 87 32 88
rect 30 87 31 88
rect 29 87 30 88
rect 28 87 29 88
rect 27 87 28 88
rect 26 87 27 88
rect 25 87 26 88
rect 24 87 25 88
rect 23 87 24 88
rect 22 87 23 88
rect 21 87 22 88
rect 20 87 21 88
rect 19 87 20 88
rect 18 87 19 88
rect 17 87 18 88
rect 16 87 17 88
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 141 88 142 89
rect 140 88 141 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 130 88 131 89
rect 129 88 130 89
rect 128 88 129 89
rect 127 88 128 89
rect 126 88 127 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 120 88 121 89
rect 82 88 83 89
rect 81 88 82 89
rect 80 88 81 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 56 88 57 89
rect 55 88 56 89
rect 54 88 55 89
rect 53 88 54 89
rect 52 88 53 89
rect 51 88 52 89
rect 50 88 51 89
rect 49 88 50 89
rect 48 88 49 89
rect 47 88 48 89
rect 46 88 47 89
rect 45 88 46 89
rect 44 88 45 89
rect 43 88 44 89
rect 42 88 43 89
rect 41 88 42 89
rect 40 88 41 89
rect 39 88 40 89
rect 38 88 39 89
rect 37 88 38 89
rect 36 88 37 89
rect 35 88 36 89
rect 34 88 35 89
rect 33 88 34 89
rect 32 88 33 89
rect 31 88 32 89
rect 30 88 31 89
rect 29 88 30 89
rect 28 88 29 89
rect 27 88 28 89
rect 26 88 27 89
rect 25 88 26 89
rect 24 88 25 89
rect 23 88 24 89
rect 22 88 23 89
rect 21 88 22 89
rect 20 88 21 89
rect 19 88 20 89
rect 18 88 19 89
rect 17 88 18 89
rect 16 88 17 89
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 141 89 142 90
rect 140 89 141 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 129 89 130 90
rect 128 89 129 90
rect 127 89 128 90
rect 126 89 127 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 120 89 121 90
rect 82 89 83 90
rect 81 89 82 90
rect 80 89 81 90
rect 79 89 80 90
rect 78 89 79 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 55 89 56 90
rect 54 89 55 90
rect 53 89 54 90
rect 52 89 53 90
rect 51 89 52 90
rect 50 89 51 90
rect 49 89 50 90
rect 48 89 49 90
rect 47 89 48 90
rect 46 89 47 90
rect 45 89 46 90
rect 44 89 45 90
rect 43 89 44 90
rect 42 89 43 90
rect 41 89 42 90
rect 40 89 41 90
rect 39 89 40 90
rect 38 89 39 90
rect 37 89 38 90
rect 36 89 37 90
rect 35 89 36 90
rect 34 89 35 90
rect 33 89 34 90
rect 32 89 33 90
rect 31 89 32 90
rect 30 89 31 90
rect 29 89 30 90
rect 28 89 29 90
rect 27 89 28 90
rect 26 89 27 90
rect 25 89 26 90
rect 24 89 25 90
rect 23 89 24 90
rect 22 89 23 90
rect 21 89 22 90
rect 20 89 21 90
rect 19 89 20 90
rect 18 89 19 90
rect 17 89 18 90
rect 16 89 17 90
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 141 90 142 91
rect 140 90 141 91
rect 131 90 132 91
rect 130 90 131 91
rect 129 90 130 91
rect 128 90 129 91
rect 127 90 128 91
rect 126 90 127 91
rect 125 90 126 91
rect 124 90 125 91
rect 123 90 124 91
rect 122 90 123 91
rect 121 90 122 91
rect 82 90 83 91
rect 81 90 82 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 77 90 78 91
rect 76 90 77 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 55 90 56 91
rect 54 90 55 91
rect 53 90 54 91
rect 52 90 53 91
rect 51 90 52 91
rect 50 90 51 91
rect 49 90 50 91
rect 48 90 49 91
rect 47 90 48 91
rect 46 90 47 91
rect 45 90 46 91
rect 44 90 45 91
rect 43 90 44 91
rect 42 90 43 91
rect 41 90 42 91
rect 40 90 41 91
rect 39 90 40 91
rect 38 90 39 91
rect 37 90 38 91
rect 36 90 37 91
rect 35 90 36 91
rect 34 90 35 91
rect 33 90 34 91
rect 32 90 33 91
rect 31 90 32 91
rect 30 90 31 91
rect 29 90 30 91
rect 28 90 29 91
rect 27 90 28 91
rect 26 90 27 91
rect 25 90 26 91
rect 24 90 25 91
rect 23 90 24 91
rect 22 90 23 91
rect 21 90 22 91
rect 20 90 21 91
rect 19 90 20 91
rect 18 90 19 91
rect 17 90 18 91
rect 16 90 17 91
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 141 91 142 92
rect 140 91 141 92
rect 130 91 131 92
rect 129 91 130 92
rect 128 91 129 92
rect 127 91 128 92
rect 126 91 127 92
rect 125 91 126 92
rect 124 91 125 92
rect 123 91 124 92
rect 122 91 123 92
rect 82 91 83 92
rect 81 91 82 92
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 74 91 75 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 54 91 55 92
rect 53 91 54 92
rect 52 91 53 92
rect 51 91 52 92
rect 50 91 51 92
rect 49 91 50 92
rect 48 91 49 92
rect 47 91 48 92
rect 46 91 47 92
rect 45 91 46 92
rect 44 91 45 92
rect 43 91 44 92
rect 42 91 43 92
rect 41 91 42 92
rect 40 91 41 92
rect 39 91 40 92
rect 38 91 39 92
rect 37 91 38 92
rect 36 91 37 92
rect 35 91 36 92
rect 34 91 35 92
rect 33 91 34 92
rect 32 91 33 92
rect 31 91 32 92
rect 30 91 31 92
rect 29 91 30 92
rect 28 91 29 92
rect 27 91 28 92
rect 26 91 27 92
rect 25 91 26 92
rect 24 91 25 92
rect 23 91 24 92
rect 22 91 23 92
rect 21 91 22 92
rect 20 91 21 92
rect 19 91 20 92
rect 18 91 19 92
rect 17 91 18 92
rect 16 91 17 92
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 141 92 142 93
rect 140 92 141 93
rect 127 92 128 93
rect 126 92 127 93
rect 125 92 126 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 72 92 73 93
rect 71 92 72 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 53 92 54 93
rect 52 92 53 93
rect 51 92 52 93
rect 50 92 51 93
rect 49 92 50 93
rect 48 92 49 93
rect 47 92 48 93
rect 46 92 47 93
rect 45 92 46 93
rect 44 92 45 93
rect 43 92 44 93
rect 42 92 43 93
rect 41 92 42 93
rect 40 92 41 93
rect 39 92 40 93
rect 38 92 39 93
rect 37 92 38 93
rect 36 92 37 93
rect 35 92 36 93
rect 34 92 35 93
rect 33 92 34 93
rect 32 92 33 93
rect 31 92 32 93
rect 30 92 31 93
rect 29 92 30 93
rect 28 92 29 93
rect 27 92 28 93
rect 26 92 27 93
rect 25 92 26 93
rect 24 92 25 93
rect 23 92 24 93
rect 22 92 23 93
rect 21 92 22 93
rect 20 92 21 93
rect 19 92 20 93
rect 18 92 19 93
rect 17 92 18 93
rect 16 92 17 93
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 70 93 71 94
rect 69 93 70 94
rect 68 93 69 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 52 93 53 94
rect 51 93 52 94
rect 50 93 51 94
rect 49 93 50 94
rect 48 93 49 94
rect 47 93 48 94
rect 46 93 47 94
rect 45 93 46 94
rect 44 93 45 94
rect 43 93 44 94
rect 42 93 43 94
rect 41 93 42 94
rect 40 93 41 94
rect 39 93 40 94
rect 38 93 39 94
rect 37 93 38 94
rect 36 93 37 94
rect 35 93 36 94
rect 34 93 35 94
rect 33 93 34 94
rect 32 93 33 94
rect 31 93 32 94
rect 30 93 31 94
rect 29 93 30 94
rect 28 93 29 94
rect 27 93 28 94
rect 26 93 27 94
rect 25 93 26 94
rect 24 93 25 94
rect 23 93 24 94
rect 22 93 23 94
rect 21 93 22 94
rect 20 93 21 94
rect 19 93 20 94
rect 18 93 19 94
rect 17 93 18 94
rect 16 93 17 94
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 68 94 69 95
rect 67 94 68 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 51 94 52 95
rect 50 94 51 95
rect 49 94 50 95
rect 48 94 49 95
rect 47 94 48 95
rect 46 94 47 95
rect 45 94 46 95
rect 44 94 45 95
rect 43 94 44 95
rect 42 94 43 95
rect 41 94 42 95
rect 40 94 41 95
rect 39 94 40 95
rect 38 94 39 95
rect 37 94 38 95
rect 36 94 37 95
rect 35 94 36 95
rect 34 94 35 95
rect 33 94 34 95
rect 32 94 33 95
rect 31 94 32 95
rect 30 94 31 95
rect 29 94 30 95
rect 28 94 29 95
rect 27 94 28 95
rect 26 94 27 95
rect 25 94 26 95
rect 24 94 25 95
rect 23 94 24 95
rect 22 94 23 95
rect 21 94 22 95
rect 20 94 21 95
rect 19 94 20 95
rect 18 94 19 95
rect 17 94 18 95
rect 16 94 17 95
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 72 95 73 96
rect 71 95 72 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 67 95 68 96
rect 66 95 67 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 50 95 51 96
rect 49 95 50 96
rect 48 95 49 96
rect 47 95 48 96
rect 46 95 47 96
rect 45 95 46 96
rect 44 95 45 96
rect 43 95 44 96
rect 42 95 43 96
rect 41 95 42 96
rect 40 95 41 96
rect 39 95 40 96
rect 38 95 39 96
rect 37 95 38 96
rect 36 95 37 96
rect 35 95 36 96
rect 34 95 35 96
rect 33 95 34 96
rect 32 95 33 96
rect 31 95 32 96
rect 30 95 31 96
rect 29 95 30 96
rect 28 95 29 96
rect 27 95 28 96
rect 26 95 27 96
rect 25 95 26 96
rect 24 95 25 96
rect 23 95 24 96
rect 22 95 23 96
rect 21 95 22 96
rect 20 95 21 96
rect 19 95 20 96
rect 18 95 19 96
rect 17 95 18 96
rect 16 95 17 96
rect 139 96 140 97
rect 138 96 139 97
rect 137 96 138 97
rect 136 96 137 97
rect 135 96 136 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 72 96 73 97
rect 71 96 72 97
rect 70 96 71 97
rect 69 96 70 97
rect 68 96 69 97
rect 67 96 68 97
rect 66 96 67 97
rect 65 96 66 97
rect 64 96 65 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 49 96 50 97
rect 48 96 49 97
rect 47 96 48 97
rect 46 96 47 97
rect 45 96 46 97
rect 44 96 45 97
rect 43 96 44 97
rect 42 96 43 97
rect 41 96 42 97
rect 40 96 41 97
rect 39 96 40 97
rect 38 96 39 97
rect 37 96 38 97
rect 36 96 37 97
rect 35 96 36 97
rect 34 96 35 97
rect 33 96 34 97
rect 32 96 33 97
rect 31 96 32 97
rect 30 96 31 97
rect 29 96 30 97
rect 28 96 29 97
rect 27 96 28 97
rect 26 96 27 97
rect 25 96 26 97
rect 24 96 25 97
rect 23 96 24 97
rect 22 96 23 97
rect 21 96 22 97
rect 20 96 21 97
rect 19 96 20 97
rect 18 96 19 97
rect 17 96 18 97
rect 16 96 17 97
rect 139 97 140 98
rect 138 97 139 98
rect 137 97 138 98
rect 136 97 137 98
rect 135 97 136 98
rect 134 97 135 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 74 97 75 98
rect 73 97 74 98
rect 72 97 73 98
rect 71 97 72 98
rect 70 97 71 98
rect 69 97 70 98
rect 68 97 69 98
rect 67 97 68 98
rect 66 97 67 98
rect 65 97 66 98
rect 64 97 65 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 50 97 51 98
rect 49 97 50 98
rect 48 97 49 98
rect 47 97 48 98
rect 46 97 47 98
rect 45 97 46 98
rect 44 97 45 98
rect 43 97 44 98
rect 42 97 43 98
rect 41 97 42 98
rect 40 97 41 98
rect 39 97 40 98
rect 38 97 39 98
rect 37 97 38 98
rect 36 97 37 98
rect 35 97 36 98
rect 34 97 35 98
rect 33 97 34 98
rect 32 97 33 98
rect 31 97 32 98
rect 30 97 31 98
rect 29 97 30 98
rect 28 97 29 98
rect 27 97 28 98
rect 26 97 27 98
rect 25 97 26 98
rect 24 97 25 98
rect 23 97 24 98
rect 22 97 23 98
rect 21 97 22 98
rect 20 97 21 98
rect 19 97 20 98
rect 18 97 19 98
rect 17 97 18 98
rect 16 97 17 98
rect 139 98 140 99
rect 138 98 139 99
rect 137 98 138 99
rect 136 98 137 99
rect 135 98 136 99
rect 134 98 135 99
rect 133 98 134 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 51 98 52 99
rect 50 98 51 99
rect 49 98 50 99
rect 48 98 49 99
rect 47 98 48 99
rect 29 98 30 99
rect 28 98 29 99
rect 27 98 28 99
rect 26 98 27 99
rect 25 98 26 99
rect 24 98 25 99
rect 23 98 24 99
rect 22 98 23 99
rect 21 98 22 99
rect 20 98 21 99
rect 19 98 20 99
rect 18 98 19 99
rect 17 98 18 99
rect 16 98 17 99
rect 139 99 140 100
rect 138 99 139 100
rect 137 99 138 100
rect 136 99 137 100
rect 135 99 136 100
rect 134 99 135 100
rect 133 99 134 100
rect 132 99 133 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 51 99 52 100
rect 50 99 51 100
rect 49 99 50 100
rect 48 99 49 100
rect 47 99 48 100
rect 29 99 30 100
rect 28 99 29 100
rect 27 99 28 100
rect 26 99 27 100
rect 25 99 26 100
rect 24 99 25 100
rect 23 99 24 100
rect 22 99 23 100
rect 21 99 22 100
rect 20 99 21 100
rect 19 99 20 100
rect 18 99 19 100
rect 17 99 18 100
rect 16 99 17 100
rect 139 100 140 101
rect 138 100 139 101
rect 137 100 138 101
rect 136 100 137 101
rect 135 100 136 101
rect 134 100 135 101
rect 133 100 134 101
rect 132 100 133 101
rect 131 100 132 101
rect 130 100 131 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 51 100 52 101
rect 50 100 51 101
rect 49 100 50 101
rect 48 100 49 101
rect 47 100 48 101
rect 29 100 30 101
rect 28 100 29 101
rect 27 100 28 101
rect 26 100 27 101
rect 25 100 26 101
rect 24 100 25 101
rect 23 100 24 101
rect 22 100 23 101
rect 21 100 22 101
rect 20 100 21 101
rect 19 100 20 101
rect 18 100 19 101
rect 17 100 18 101
rect 16 100 17 101
rect 139 101 140 102
rect 138 101 139 102
rect 137 101 138 102
rect 136 101 137 102
rect 135 101 136 102
rect 134 101 135 102
rect 133 101 134 102
rect 132 101 133 102
rect 131 101 132 102
rect 130 101 131 102
rect 129 101 130 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 51 101 52 102
rect 50 101 51 102
rect 49 101 50 102
rect 48 101 49 102
rect 47 101 48 102
rect 29 101 30 102
rect 28 101 29 102
rect 27 101 28 102
rect 26 101 27 102
rect 25 101 26 102
rect 24 101 25 102
rect 23 101 24 102
rect 22 101 23 102
rect 21 101 22 102
rect 20 101 21 102
rect 19 101 20 102
rect 18 101 19 102
rect 17 101 18 102
rect 16 101 17 102
rect 139 102 140 103
rect 138 102 139 103
rect 137 102 138 103
rect 136 102 137 103
rect 133 102 134 103
rect 132 102 133 103
rect 131 102 132 103
rect 130 102 131 103
rect 129 102 130 103
rect 128 102 129 103
rect 127 102 128 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 51 102 52 103
rect 50 102 51 103
rect 49 102 50 103
rect 48 102 49 103
rect 47 102 48 103
rect 29 102 30 103
rect 28 102 29 103
rect 27 102 28 103
rect 26 102 27 103
rect 25 102 26 103
rect 24 102 25 103
rect 23 102 24 103
rect 22 102 23 103
rect 21 102 22 103
rect 20 102 21 103
rect 19 102 20 103
rect 18 102 19 103
rect 17 102 18 103
rect 16 102 17 103
rect 139 103 140 104
rect 138 103 139 104
rect 137 103 138 104
rect 136 103 137 104
rect 132 103 133 104
rect 131 103 132 104
rect 130 103 131 104
rect 129 103 130 104
rect 128 103 129 104
rect 127 103 128 104
rect 126 103 127 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 50 103 51 104
rect 49 103 50 104
rect 48 103 49 104
rect 47 103 48 104
rect 29 103 30 104
rect 28 103 29 104
rect 27 103 28 104
rect 26 103 27 104
rect 25 103 26 104
rect 24 103 25 104
rect 23 103 24 104
rect 22 103 23 104
rect 21 103 22 104
rect 20 103 21 104
rect 19 103 20 104
rect 18 103 19 104
rect 17 103 18 104
rect 16 103 17 104
rect 139 104 140 105
rect 138 104 139 105
rect 137 104 138 105
rect 136 104 137 105
rect 130 104 131 105
rect 129 104 130 105
rect 128 104 129 105
rect 127 104 128 105
rect 126 104 127 105
rect 125 104 126 105
rect 124 104 125 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 51 104 52 105
rect 50 104 51 105
rect 49 104 50 105
rect 48 104 49 105
rect 47 104 48 105
rect 29 104 30 105
rect 28 104 29 105
rect 27 104 28 105
rect 26 104 27 105
rect 25 104 26 105
rect 24 104 25 105
rect 23 104 24 105
rect 22 104 23 105
rect 21 104 22 105
rect 20 104 21 105
rect 19 104 20 105
rect 18 104 19 105
rect 17 104 18 105
rect 16 104 17 105
rect 139 105 140 106
rect 138 105 139 106
rect 137 105 138 106
rect 136 105 137 106
rect 129 105 130 106
rect 128 105 129 106
rect 127 105 128 106
rect 126 105 127 106
rect 125 105 126 106
rect 124 105 125 106
rect 123 105 124 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 51 105 52 106
rect 50 105 51 106
rect 49 105 50 106
rect 48 105 49 106
rect 47 105 48 106
rect 29 105 30 106
rect 28 105 29 106
rect 27 105 28 106
rect 26 105 27 106
rect 25 105 26 106
rect 24 105 25 106
rect 23 105 24 106
rect 22 105 23 106
rect 21 105 22 106
rect 20 105 21 106
rect 19 105 20 106
rect 18 105 19 106
rect 17 105 18 106
rect 16 105 17 106
rect 139 106 140 107
rect 138 106 139 107
rect 137 106 138 107
rect 136 106 137 107
rect 127 106 128 107
rect 126 106 127 107
rect 125 106 126 107
rect 124 106 125 107
rect 123 106 124 107
rect 122 106 123 107
rect 121 106 122 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 51 106 52 107
rect 50 106 51 107
rect 49 106 50 107
rect 48 106 49 107
rect 47 106 48 107
rect 30 106 31 107
rect 29 106 30 107
rect 28 106 29 107
rect 27 106 28 107
rect 26 106 27 107
rect 25 106 26 107
rect 24 106 25 107
rect 23 106 24 107
rect 22 106 23 107
rect 21 106 22 107
rect 20 106 21 107
rect 19 106 20 107
rect 18 106 19 107
rect 17 106 18 107
rect 16 106 17 107
rect 139 107 140 108
rect 138 107 139 108
rect 137 107 138 108
rect 136 107 137 108
rect 135 107 136 108
rect 126 107 127 108
rect 125 107 126 108
rect 124 107 125 108
rect 123 107 124 108
rect 122 107 123 108
rect 121 107 122 108
rect 120 107 121 108
rect 119 107 120 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 51 107 52 108
rect 50 107 51 108
rect 49 107 50 108
rect 48 107 49 108
rect 47 107 48 108
rect 46 107 47 108
rect 30 107 31 108
rect 29 107 30 108
rect 28 107 29 108
rect 27 107 28 108
rect 26 107 27 108
rect 25 107 26 108
rect 24 107 25 108
rect 23 107 24 108
rect 22 107 23 108
rect 21 107 22 108
rect 20 107 21 108
rect 19 107 20 108
rect 18 107 19 108
rect 17 107 18 108
rect 16 107 17 108
rect 144 108 145 109
rect 143 108 144 109
rect 142 108 143 109
rect 141 108 142 109
rect 140 108 141 109
rect 139 108 140 109
rect 138 108 139 109
rect 137 108 138 109
rect 136 108 137 109
rect 135 108 136 109
rect 134 108 135 109
rect 133 108 134 109
rect 132 108 133 109
rect 131 108 132 109
rect 130 108 131 109
rect 129 108 130 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 125 108 126 109
rect 124 108 125 109
rect 123 108 124 109
rect 122 108 123 109
rect 121 108 122 109
rect 120 108 121 109
rect 119 108 120 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 51 108 52 109
rect 50 108 51 109
rect 49 108 50 109
rect 48 108 49 109
rect 47 108 48 109
rect 46 108 47 109
rect 31 108 32 109
rect 30 108 31 109
rect 29 108 30 109
rect 28 108 29 109
rect 27 108 28 109
rect 26 108 27 109
rect 25 108 26 109
rect 24 108 25 109
rect 23 108 24 109
rect 22 108 23 109
rect 21 108 22 109
rect 20 108 21 109
rect 19 108 20 109
rect 18 108 19 109
rect 17 108 18 109
rect 16 108 17 109
rect 144 109 145 110
rect 143 109 144 110
rect 142 109 143 110
rect 141 109 142 110
rect 140 109 141 110
rect 139 109 140 110
rect 138 109 139 110
rect 137 109 138 110
rect 136 109 137 110
rect 135 109 136 110
rect 134 109 135 110
rect 133 109 134 110
rect 132 109 133 110
rect 131 109 132 110
rect 130 109 131 110
rect 129 109 130 110
rect 128 109 129 110
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 124 109 125 110
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 120 109 121 110
rect 119 109 120 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 52 109 53 110
rect 51 109 52 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 47 109 48 110
rect 46 109 47 110
rect 45 109 46 110
rect 31 109 32 110
rect 30 109 31 110
rect 29 109 30 110
rect 28 109 29 110
rect 27 109 28 110
rect 26 109 27 110
rect 25 109 26 110
rect 24 109 25 110
rect 23 109 24 110
rect 22 109 23 110
rect 21 109 22 110
rect 20 109 21 110
rect 19 109 20 110
rect 18 109 19 110
rect 17 109 18 110
rect 16 109 17 110
rect 144 110 145 111
rect 143 110 144 111
rect 142 110 143 111
rect 141 110 142 111
rect 140 110 141 111
rect 139 110 140 111
rect 138 110 139 111
rect 137 110 138 111
rect 136 110 137 111
rect 135 110 136 111
rect 134 110 135 111
rect 133 110 134 111
rect 132 110 133 111
rect 131 110 132 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 127 110 128 111
rect 126 110 127 111
rect 125 110 126 111
rect 124 110 125 111
rect 123 110 124 111
rect 122 110 123 111
rect 121 110 122 111
rect 120 110 121 111
rect 119 110 120 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 52 110 53 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 47 110 48 111
rect 46 110 47 111
rect 45 110 46 111
rect 44 110 45 111
rect 33 110 34 111
rect 32 110 33 111
rect 31 110 32 111
rect 30 110 31 111
rect 29 110 30 111
rect 28 110 29 111
rect 27 110 28 111
rect 26 110 27 111
rect 25 110 26 111
rect 24 110 25 111
rect 23 110 24 111
rect 22 110 23 111
rect 21 110 22 111
rect 20 110 21 111
rect 19 110 20 111
rect 18 110 19 111
rect 17 110 18 111
rect 16 110 17 111
rect 144 111 145 112
rect 143 111 144 112
rect 142 111 143 112
rect 141 111 142 112
rect 140 111 141 112
rect 139 111 140 112
rect 138 111 139 112
rect 137 111 138 112
rect 136 111 137 112
rect 135 111 136 112
rect 134 111 135 112
rect 133 111 134 112
rect 132 111 133 112
rect 131 111 132 112
rect 130 111 131 112
rect 129 111 130 112
rect 128 111 129 112
rect 127 111 128 112
rect 126 111 127 112
rect 125 111 126 112
rect 124 111 125 112
rect 123 111 124 112
rect 122 111 123 112
rect 121 111 122 112
rect 120 111 121 112
rect 119 111 120 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 52 111 53 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 46 111 47 112
rect 45 111 46 112
rect 44 111 45 112
rect 43 111 44 112
rect 42 111 43 112
rect 41 111 42 112
rect 35 111 36 112
rect 34 111 35 112
rect 33 111 34 112
rect 32 111 33 112
rect 31 111 32 112
rect 30 111 31 112
rect 29 111 30 112
rect 28 111 29 112
rect 27 111 28 112
rect 26 111 27 112
rect 25 111 26 112
rect 24 111 25 112
rect 23 111 24 112
rect 22 111 23 112
rect 21 111 22 112
rect 20 111 21 112
rect 19 111 20 112
rect 18 111 19 112
rect 17 111 18 112
rect 16 111 17 112
rect 144 112 145 113
rect 143 112 144 113
rect 142 112 143 113
rect 141 112 142 113
rect 140 112 141 113
rect 139 112 140 113
rect 138 112 139 113
rect 137 112 138 113
rect 136 112 137 113
rect 135 112 136 113
rect 134 112 135 113
rect 133 112 134 113
rect 132 112 133 113
rect 131 112 132 113
rect 130 112 131 113
rect 129 112 130 113
rect 128 112 129 113
rect 127 112 128 113
rect 126 112 127 113
rect 125 112 126 113
rect 124 112 125 113
rect 123 112 124 113
rect 122 112 123 113
rect 121 112 122 113
rect 120 112 121 113
rect 119 112 120 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 53 112 54 113
rect 52 112 53 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 45 112 46 113
rect 44 112 45 113
rect 43 112 44 113
rect 42 112 43 113
rect 41 112 42 113
rect 40 112 41 113
rect 39 112 40 113
rect 38 112 39 113
rect 37 112 38 113
rect 36 112 37 113
rect 35 112 36 113
rect 34 112 35 113
rect 33 112 34 113
rect 32 112 33 113
rect 31 112 32 113
rect 30 112 31 113
rect 29 112 30 113
rect 28 112 29 113
rect 27 112 28 113
rect 26 112 27 113
rect 25 112 26 113
rect 24 112 25 113
rect 23 112 24 113
rect 22 112 23 113
rect 21 112 22 113
rect 20 112 21 113
rect 19 112 20 113
rect 18 112 19 113
rect 17 112 18 113
rect 16 112 17 113
rect 139 113 140 114
rect 138 113 139 114
rect 137 113 138 114
rect 136 113 137 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 53 113 54 114
rect 52 113 53 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 42 113 43 114
rect 41 113 42 114
rect 40 113 41 114
rect 39 113 40 114
rect 38 113 39 114
rect 37 113 38 114
rect 36 113 37 114
rect 35 113 36 114
rect 34 113 35 114
rect 33 113 34 114
rect 32 113 33 114
rect 31 113 32 114
rect 30 113 31 114
rect 29 113 30 114
rect 28 113 29 114
rect 27 113 28 114
rect 26 113 27 114
rect 25 113 26 114
rect 24 113 25 114
rect 23 113 24 114
rect 22 113 23 114
rect 21 113 22 114
rect 20 113 21 114
rect 19 113 20 114
rect 18 113 19 114
rect 17 113 18 114
rect 139 114 140 115
rect 138 114 139 115
rect 137 114 138 115
rect 136 114 137 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 53 114 54 115
rect 52 114 53 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 35 114 36 115
rect 34 114 35 115
rect 33 114 34 115
rect 32 114 33 115
rect 31 114 32 115
rect 30 114 31 115
rect 29 114 30 115
rect 28 114 29 115
rect 27 114 28 115
rect 26 114 27 115
rect 25 114 26 115
rect 24 114 25 115
rect 23 114 24 115
rect 22 114 23 115
rect 21 114 22 115
rect 20 114 21 115
rect 19 114 20 115
rect 18 114 19 115
rect 17 114 18 115
rect 139 115 140 116
rect 138 115 139 116
rect 137 115 138 116
rect 136 115 137 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 55 115 56 116
rect 54 115 55 116
rect 53 115 54 116
rect 52 115 53 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 35 115 36 116
rect 34 115 35 116
rect 33 115 34 116
rect 32 115 33 116
rect 31 115 32 116
rect 30 115 31 116
rect 29 115 30 116
rect 28 115 29 116
rect 27 115 28 116
rect 26 115 27 116
rect 25 115 26 116
rect 24 115 25 116
rect 23 115 24 116
rect 22 115 23 116
rect 21 115 22 116
rect 20 115 21 116
rect 19 115 20 116
rect 18 115 19 116
rect 17 115 18 116
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 55 116 56 117
rect 54 116 55 117
rect 53 116 54 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 34 116 35 117
rect 33 116 34 117
rect 32 116 33 117
rect 31 116 32 117
rect 30 116 31 117
rect 29 116 30 117
rect 28 116 29 117
rect 27 116 28 117
rect 26 116 27 117
rect 25 116 26 117
rect 24 116 25 117
rect 23 116 24 117
rect 22 116 23 117
rect 21 116 22 117
rect 20 116 21 117
rect 19 116 20 117
rect 18 116 19 117
rect 17 116 18 117
rect 58 117 59 118
rect 57 117 58 118
rect 56 117 57 118
rect 55 117 56 118
rect 54 117 55 118
rect 53 117 54 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 35 117 36 118
rect 34 117 35 118
rect 33 117 34 118
rect 32 117 33 118
rect 31 117 32 118
rect 30 117 31 118
rect 29 117 30 118
rect 28 117 29 118
rect 27 117 28 118
rect 26 117 27 118
rect 25 117 26 118
rect 24 117 25 118
rect 23 117 24 118
rect 22 117 23 118
rect 21 117 22 118
rect 20 117 21 118
rect 19 117 20 118
rect 18 117 19 118
rect 17 117 18 118
rect 149 118 150 119
rect 148 118 149 119
rect 147 118 148 119
rect 146 118 147 119
rect 58 118 59 119
rect 57 118 58 119
rect 56 118 57 119
rect 55 118 56 119
rect 54 118 55 119
rect 53 118 54 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 35 118 36 119
rect 34 118 35 119
rect 33 118 34 119
rect 32 118 33 119
rect 31 118 32 119
rect 30 118 31 119
rect 29 118 30 119
rect 28 118 29 119
rect 27 118 28 119
rect 26 118 27 119
rect 25 118 26 119
rect 24 118 25 119
rect 23 118 24 119
rect 22 118 23 119
rect 21 118 22 119
rect 20 118 21 119
rect 19 118 20 119
rect 18 118 19 119
rect 17 118 18 119
rect 149 119 150 120
rect 148 119 149 120
rect 147 119 148 120
rect 146 119 147 120
rect 145 119 146 120
rect 144 119 145 120
rect 143 119 144 120
rect 142 119 143 120
rect 141 119 142 120
rect 57 119 58 120
rect 56 119 57 120
rect 55 119 56 120
rect 54 119 55 120
rect 53 119 54 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 35 119 36 120
rect 34 119 35 120
rect 33 119 34 120
rect 32 119 33 120
rect 31 119 32 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 27 119 28 120
rect 26 119 27 120
rect 25 119 26 120
rect 24 119 25 120
rect 23 119 24 120
rect 22 119 23 120
rect 21 119 22 120
rect 20 119 21 120
rect 19 119 20 120
rect 18 119 19 120
rect 149 120 150 121
rect 148 120 149 121
rect 147 120 148 121
rect 146 120 147 121
rect 145 120 146 121
rect 144 120 145 121
rect 143 120 144 121
rect 142 120 143 121
rect 141 120 142 121
rect 57 120 58 121
rect 56 120 57 121
rect 55 120 56 121
rect 54 120 55 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 35 120 36 121
rect 34 120 35 121
rect 33 120 34 121
rect 32 120 33 121
rect 31 120 32 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 26 120 27 121
rect 25 120 26 121
rect 24 120 25 121
rect 23 120 24 121
rect 22 120 23 121
rect 21 120 22 121
rect 20 120 21 121
rect 19 120 20 121
rect 18 120 19 121
rect 149 121 150 122
rect 148 121 149 122
rect 147 121 148 122
rect 146 121 147 122
rect 145 121 146 122
rect 144 121 145 122
rect 143 121 144 122
rect 142 121 143 122
rect 141 121 142 122
rect 56 121 57 122
rect 55 121 56 122
rect 54 121 55 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 36 121 37 122
rect 35 121 36 122
rect 34 121 35 122
rect 33 121 34 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 26 121 27 122
rect 25 121 26 122
rect 24 121 25 122
rect 23 121 24 122
rect 22 121 23 122
rect 21 121 22 122
rect 20 121 21 122
rect 19 121 20 122
rect 18 121 19 122
rect 147 122 148 123
rect 146 122 147 123
rect 145 122 146 123
rect 144 122 145 123
rect 143 122 144 123
rect 142 122 143 123
rect 141 122 142 123
rect 56 122 57 123
rect 55 122 56 123
rect 54 122 55 123
rect 53 122 54 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 36 122 37 123
rect 35 122 36 123
rect 34 122 35 123
rect 33 122 34 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 26 122 27 123
rect 25 122 26 123
rect 24 122 25 123
rect 23 122 24 123
rect 22 122 23 123
rect 21 122 22 123
rect 20 122 21 123
rect 19 122 20 123
rect 144 123 145 124
rect 143 123 144 124
rect 142 123 143 124
rect 141 123 142 124
rect 55 123 56 124
rect 54 123 55 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 36 123 37 124
rect 35 123 36 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 26 123 27 124
rect 25 123 26 124
rect 24 123 25 124
rect 23 123 24 124
rect 22 123 23 124
rect 21 123 22 124
rect 20 123 21 124
rect 19 123 20 124
rect 141 124 142 125
rect 54 124 55 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 36 124 37 125
rect 35 124 36 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 26 124 27 125
rect 25 124 26 125
rect 24 124 25 125
rect 23 124 24 125
rect 22 124 23 125
rect 21 124 22 125
rect 20 124 21 125
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 37 125 38 126
rect 36 125 37 126
rect 35 125 36 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 27 125 28 126
rect 26 125 27 126
rect 25 125 26 126
rect 24 125 25 126
rect 23 125 24 126
rect 22 125 23 126
rect 21 125 22 126
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 37 126 38 127
rect 36 126 37 127
rect 35 126 36 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 27 126 28 127
rect 26 126 27 127
rect 25 126 26 127
rect 24 126 25 127
rect 23 126 24 127
rect 22 126 23 127
rect 21 126 22 127
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 38 127 39 128
rect 37 127 38 128
rect 36 127 37 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 27 127 28 128
rect 26 127 27 128
rect 25 127 26 128
rect 24 127 25 128
rect 23 127 24 128
rect 22 127 23 128
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 38 128 39 129
rect 37 128 38 129
rect 36 128 37 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 28 128 29 129
rect 27 128 28 129
rect 26 128 27 129
rect 25 128 26 129
rect 24 128 25 129
rect 23 128 24 129
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 39 129 40 130
rect 38 129 39 130
rect 37 129 38 130
rect 36 129 37 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 28 129 29 130
rect 27 129 28 130
rect 26 129 27 130
rect 25 129 26 130
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 40 130 41 131
rect 39 130 40 131
rect 38 130 39 131
rect 37 130 38 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 29 130 30 131
rect 28 130 29 131
rect 27 130 28 131
rect 26 130 27 131
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 41 131 42 132
rect 40 131 41 132
rect 39 131 40 132
rect 38 131 39 132
rect 37 131 38 132
rect 36 131 37 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 30 131 31 132
rect 29 131 30 132
rect 28 131 29 132
rect 42 132 43 133
rect 41 132 42 133
rect 40 132 41 133
rect 39 132 40 133
rect 38 132 39 133
rect 37 132 38 133
rect 36 132 37 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 144 138 145 139
rect 143 138 144 139
rect 142 138 143 139
rect 141 138 142 139
rect 140 138 141 139
rect 139 138 140 139
rect 144 139 145 140
rect 143 139 144 140
rect 142 139 143 140
rect 141 139 142 140
rect 140 139 141 140
rect 144 140 145 141
rect 143 140 144 141
rect 142 140 143 141
rect 141 140 142 141
rect 140 140 141 141
rect 52 140 53 141
rect 51 140 52 141
rect 50 140 51 141
rect 49 140 50 141
rect 48 140 49 141
rect 47 140 48 141
rect 46 140 47 141
rect 45 140 46 141
rect 44 140 45 141
rect 43 140 44 141
rect 42 140 43 141
rect 41 140 42 141
rect 40 140 41 141
rect 39 140 40 141
rect 38 140 39 141
rect 37 140 38 141
rect 36 140 37 141
rect 35 140 36 141
rect 34 140 35 141
rect 33 140 34 141
rect 32 140 33 141
rect 31 140 32 141
rect 30 140 31 141
rect 29 140 30 141
rect 28 140 29 141
rect 27 140 28 141
rect 26 140 27 141
rect 25 140 26 141
rect 24 140 25 141
rect 23 140 24 141
rect 22 140 23 141
rect 21 140 22 141
rect 20 140 21 141
rect 19 140 20 141
rect 18 140 19 141
rect 17 140 18 141
rect 16 140 17 141
rect 144 141 145 142
rect 143 141 144 142
rect 142 141 143 142
rect 141 141 142 142
rect 140 141 141 142
rect 63 141 64 142
rect 62 141 63 142
rect 61 141 62 142
rect 60 141 61 142
rect 59 141 60 142
rect 58 141 59 142
rect 57 141 58 142
rect 56 141 57 142
rect 55 141 56 142
rect 54 141 55 142
rect 53 141 54 142
rect 52 141 53 142
rect 51 141 52 142
rect 50 141 51 142
rect 49 141 50 142
rect 48 141 49 142
rect 47 141 48 142
rect 46 141 47 142
rect 45 141 46 142
rect 44 141 45 142
rect 43 141 44 142
rect 42 141 43 142
rect 41 141 42 142
rect 40 141 41 142
rect 39 141 40 142
rect 38 141 39 142
rect 37 141 38 142
rect 36 141 37 142
rect 35 141 36 142
rect 34 141 35 142
rect 33 141 34 142
rect 32 141 33 142
rect 31 141 32 142
rect 30 141 31 142
rect 29 141 30 142
rect 28 141 29 142
rect 27 141 28 142
rect 26 141 27 142
rect 25 141 26 142
rect 24 141 25 142
rect 23 141 24 142
rect 22 141 23 142
rect 21 141 22 142
rect 20 141 21 142
rect 19 141 20 142
rect 18 141 19 142
rect 17 141 18 142
rect 16 141 17 142
rect 144 142 145 143
rect 143 142 144 143
rect 142 142 143 143
rect 141 142 142 143
rect 140 142 141 143
rect 66 142 67 143
rect 65 142 66 143
rect 64 142 65 143
rect 63 142 64 143
rect 62 142 63 143
rect 61 142 62 143
rect 60 142 61 143
rect 59 142 60 143
rect 58 142 59 143
rect 57 142 58 143
rect 56 142 57 143
rect 55 142 56 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 50 142 51 143
rect 49 142 50 143
rect 48 142 49 143
rect 47 142 48 143
rect 46 142 47 143
rect 45 142 46 143
rect 44 142 45 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 37 142 38 143
rect 36 142 37 143
rect 35 142 36 143
rect 34 142 35 143
rect 33 142 34 143
rect 32 142 33 143
rect 31 142 32 143
rect 30 142 31 143
rect 29 142 30 143
rect 28 142 29 143
rect 27 142 28 143
rect 26 142 27 143
rect 25 142 26 143
rect 24 142 25 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 19 142 20 143
rect 18 142 19 143
rect 17 142 18 143
rect 16 142 17 143
rect 144 143 145 144
rect 143 143 144 144
rect 142 143 143 144
rect 141 143 142 144
rect 140 143 141 144
rect 139 143 140 144
rect 69 143 70 144
rect 68 143 69 144
rect 67 143 68 144
rect 66 143 67 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 51 143 52 144
rect 50 143 51 144
rect 49 143 50 144
rect 48 143 49 144
rect 47 143 48 144
rect 46 143 47 144
rect 45 143 46 144
rect 44 143 45 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 37 143 38 144
rect 36 143 37 144
rect 35 143 36 144
rect 34 143 35 144
rect 33 143 34 144
rect 32 143 33 144
rect 31 143 32 144
rect 30 143 31 144
rect 29 143 30 144
rect 28 143 29 144
rect 27 143 28 144
rect 26 143 27 144
rect 25 143 26 144
rect 24 143 25 144
rect 23 143 24 144
rect 22 143 23 144
rect 21 143 22 144
rect 20 143 21 144
rect 19 143 20 144
rect 18 143 19 144
rect 17 143 18 144
rect 16 143 17 144
rect 144 144 145 145
rect 143 144 144 145
rect 142 144 143 145
rect 141 144 142 145
rect 140 144 141 145
rect 139 144 140 145
rect 138 144 139 145
rect 71 144 72 145
rect 70 144 71 145
rect 69 144 70 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 52 144 53 145
rect 51 144 52 145
rect 50 144 51 145
rect 49 144 50 145
rect 48 144 49 145
rect 47 144 48 145
rect 46 144 47 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 37 144 38 145
rect 36 144 37 145
rect 35 144 36 145
rect 34 144 35 145
rect 33 144 34 145
rect 32 144 33 145
rect 31 144 32 145
rect 30 144 31 145
rect 29 144 30 145
rect 28 144 29 145
rect 27 144 28 145
rect 26 144 27 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 21 144 22 145
rect 20 144 21 145
rect 19 144 20 145
rect 18 144 19 145
rect 17 144 18 145
rect 16 144 17 145
rect 143 145 144 146
rect 142 145 143 146
rect 141 145 142 146
rect 140 145 141 146
rect 139 145 140 146
rect 138 145 139 146
rect 137 145 138 146
rect 136 145 137 146
rect 135 145 136 146
rect 134 145 135 146
rect 133 145 134 146
rect 132 145 133 146
rect 131 145 132 146
rect 130 145 131 146
rect 129 145 130 146
rect 128 145 129 146
rect 127 145 128 146
rect 126 145 127 146
rect 125 145 126 146
rect 124 145 125 146
rect 123 145 124 146
rect 122 145 123 146
rect 121 145 122 146
rect 120 145 121 146
rect 119 145 120 146
rect 72 145 73 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 54 145 55 146
rect 53 145 54 146
rect 52 145 53 146
rect 51 145 52 146
rect 50 145 51 146
rect 49 145 50 146
rect 48 145 49 146
rect 47 145 48 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 37 145 38 146
rect 36 145 37 146
rect 35 145 36 146
rect 34 145 35 146
rect 33 145 34 146
rect 32 145 33 146
rect 31 145 32 146
rect 30 145 31 146
rect 29 145 30 146
rect 28 145 29 146
rect 27 145 28 146
rect 26 145 27 146
rect 25 145 26 146
rect 24 145 25 146
rect 23 145 24 146
rect 22 145 23 146
rect 21 145 22 146
rect 20 145 21 146
rect 19 145 20 146
rect 18 145 19 146
rect 17 145 18 146
rect 16 145 17 146
rect 143 146 144 147
rect 142 146 143 147
rect 141 146 142 147
rect 140 146 141 147
rect 139 146 140 147
rect 138 146 139 147
rect 137 146 138 147
rect 136 146 137 147
rect 135 146 136 147
rect 134 146 135 147
rect 133 146 134 147
rect 132 146 133 147
rect 131 146 132 147
rect 130 146 131 147
rect 129 146 130 147
rect 128 146 129 147
rect 127 146 128 147
rect 126 146 127 147
rect 125 146 126 147
rect 124 146 125 147
rect 123 146 124 147
rect 122 146 123 147
rect 121 146 122 147
rect 120 146 121 147
rect 119 146 120 147
rect 74 146 75 147
rect 73 146 74 147
rect 72 146 73 147
rect 71 146 72 147
rect 70 146 71 147
rect 69 146 70 147
rect 68 146 69 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 57 146 58 147
rect 56 146 57 147
rect 55 146 56 147
rect 54 146 55 147
rect 53 146 54 147
rect 52 146 53 147
rect 51 146 52 147
rect 50 146 51 147
rect 49 146 50 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 37 146 38 147
rect 36 146 37 147
rect 35 146 36 147
rect 34 146 35 147
rect 33 146 34 147
rect 32 146 33 147
rect 31 146 32 147
rect 30 146 31 147
rect 29 146 30 147
rect 28 146 29 147
rect 27 146 28 147
rect 26 146 27 147
rect 25 146 26 147
rect 24 146 25 147
rect 23 146 24 147
rect 22 146 23 147
rect 21 146 22 147
rect 20 146 21 147
rect 19 146 20 147
rect 18 146 19 147
rect 17 146 18 147
rect 16 146 17 147
rect 142 147 143 148
rect 141 147 142 148
rect 140 147 141 148
rect 139 147 140 148
rect 138 147 139 148
rect 137 147 138 148
rect 136 147 137 148
rect 135 147 136 148
rect 134 147 135 148
rect 133 147 134 148
rect 132 147 133 148
rect 131 147 132 148
rect 130 147 131 148
rect 129 147 130 148
rect 128 147 129 148
rect 127 147 128 148
rect 126 147 127 148
rect 125 147 126 148
rect 124 147 125 148
rect 123 147 124 148
rect 122 147 123 148
rect 121 147 122 148
rect 120 147 121 148
rect 119 147 120 148
rect 75 147 76 148
rect 74 147 75 148
rect 73 147 74 148
rect 72 147 73 148
rect 71 147 72 148
rect 70 147 71 148
rect 69 147 70 148
rect 68 147 69 148
rect 67 147 68 148
rect 66 147 67 148
rect 65 147 66 148
rect 64 147 65 148
rect 63 147 64 148
rect 62 147 63 148
rect 61 147 62 148
rect 60 147 61 148
rect 59 147 60 148
rect 58 147 59 148
rect 57 147 58 148
rect 56 147 57 148
rect 55 147 56 148
rect 54 147 55 148
rect 53 147 54 148
rect 52 147 53 148
rect 51 147 52 148
rect 50 147 51 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 36 147 37 148
rect 35 147 36 148
rect 34 147 35 148
rect 33 147 34 148
rect 32 147 33 148
rect 31 147 32 148
rect 30 147 31 148
rect 29 147 30 148
rect 28 147 29 148
rect 27 147 28 148
rect 26 147 27 148
rect 25 147 26 148
rect 24 147 25 148
rect 23 147 24 148
rect 22 147 23 148
rect 21 147 22 148
rect 20 147 21 148
rect 19 147 20 148
rect 18 147 19 148
rect 17 147 18 148
rect 16 147 17 148
rect 141 148 142 149
rect 140 148 141 149
rect 139 148 140 149
rect 138 148 139 149
rect 137 148 138 149
rect 136 148 137 149
rect 135 148 136 149
rect 134 148 135 149
rect 133 148 134 149
rect 132 148 133 149
rect 131 148 132 149
rect 130 148 131 149
rect 129 148 130 149
rect 128 148 129 149
rect 127 148 128 149
rect 126 148 127 149
rect 125 148 126 149
rect 124 148 125 149
rect 123 148 124 149
rect 122 148 123 149
rect 121 148 122 149
rect 120 148 121 149
rect 119 148 120 149
rect 76 148 77 149
rect 75 148 76 149
rect 74 148 75 149
rect 73 148 74 149
rect 72 148 73 149
rect 71 148 72 149
rect 70 148 71 149
rect 69 148 70 149
rect 68 148 69 149
rect 67 148 68 149
rect 66 148 67 149
rect 65 148 66 149
rect 64 148 65 149
rect 63 148 64 149
rect 62 148 63 149
rect 61 148 62 149
rect 60 148 61 149
rect 59 148 60 149
rect 58 148 59 149
rect 57 148 58 149
rect 56 148 57 149
rect 55 148 56 149
rect 54 148 55 149
rect 53 148 54 149
rect 52 148 53 149
rect 51 148 52 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 36 148 37 149
rect 35 148 36 149
rect 34 148 35 149
rect 33 148 34 149
rect 32 148 33 149
rect 31 148 32 149
rect 30 148 31 149
rect 29 148 30 149
rect 28 148 29 149
rect 27 148 28 149
rect 26 148 27 149
rect 25 148 26 149
rect 24 148 25 149
rect 23 148 24 149
rect 22 148 23 149
rect 21 148 22 149
rect 20 148 21 149
rect 19 148 20 149
rect 18 148 19 149
rect 17 148 18 149
rect 16 148 17 149
rect 140 149 141 150
rect 139 149 140 150
rect 138 149 139 150
rect 137 149 138 150
rect 136 149 137 150
rect 135 149 136 150
rect 134 149 135 150
rect 133 149 134 150
rect 132 149 133 150
rect 131 149 132 150
rect 130 149 131 150
rect 129 149 130 150
rect 128 149 129 150
rect 127 149 128 150
rect 126 149 127 150
rect 125 149 126 150
rect 124 149 125 150
rect 123 149 124 150
rect 122 149 123 150
rect 121 149 122 150
rect 120 149 121 150
rect 119 149 120 150
rect 77 149 78 150
rect 76 149 77 150
rect 75 149 76 150
rect 74 149 75 150
rect 73 149 74 150
rect 72 149 73 150
rect 71 149 72 150
rect 70 149 71 150
rect 69 149 70 150
rect 68 149 69 150
rect 67 149 68 150
rect 66 149 67 150
rect 65 149 66 150
rect 64 149 65 150
rect 63 149 64 150
rect 62 149 63 150
rect 61 149 62 150
rect 60 149 61 150
rect 59 149 60 150
rect 58 149 59 150
rect 57 149 58 150
rect 56 149 57 150
rect 55 149 56 150
rect 54 149 55 150
rect 53 149 54 150
rect 52 149 53 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 38 149 39 150
rect 37 149 38 150
rect 36 149 37 150
rect 35 149 36 150
rect 34 149 35 150
rect 33 149 34 150
rect 32 149 33 150
rect 31 149 32 150
rect 30 149 31 150
rect 29 149 30 150
rect 28 149 29 150
rect 27 149 28 150
rect 26 149 27 150
rect 25 149 26 150
rect 24 149 25 150
rect 23 149 24 150
rect 22 149 23 150
rect 21 149 22 150
rect 20 149 21 150
rect 19 149 20 150
rect 18 149 19 150
rect 17 149 18 150
rect 16 149 17 150
rect 137 150 138 151
rect 136 150 137 151
rect 135 150 136 151
rect 134 150 135 151
rect 133 150 134 151
rect 132 150 133 151
rect 131 150 132 151
rect 130 150 131 151
rect 129 150 130 151
rect 128 150 129 151
rect 127 150 128 151
rect 126 150 127 151
rect 125 150 126 151
rect 124 150 125 151
rect 123 150 124 151
rect 122 150 123 151
rect 121 150 122 151
rect 120 150 121 151
rect 119 150 120 151
rect 78 150 79 151
rect 77 150 78 151
rect 76 150 77 151
rect 75 150 76 151
rect 74 150 75 151
rect 73 150 74 151
rect 72 150 73 151
rect 71 150 72 151
rect 70 150 71 151
rect 69 150 70 151
rect 68 150 69 151
rect 67 150 68 151
rect 66 150 67 151
rect 65 150 66 151
rect 64 150 65 151
rect 63 150 64 151
rect 62 150 63 151
rect 61 150 62 151
rect 60 150 61 151
rect 59 150 60 151
rect 58 150 59 151
rect 57 150 58 151
rect 56 150 57 151
rect 55 150 56 151
rect 54 150 55 151
rect 53 150 54 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 38 150 39 151
rect 37 150 38 151
rect 36 150 37 151
rect 35 150 36 151
rect 34 150 35 151
rect 33 150 34 151
rect 32 150 33 151
rect 31 150 32 151
rect 30 150 31 151
rect 29 150 30 151
rect 28 150 29 151
rect 27 150 28 151
rect 26 150 27 151
rect 25 150 26 151
rect 24 150 25 151
rect 23 150 24 151
rect 22 150 23 151
rect 21 150 22 151
rect 20 150 21 151
rect 19 150 20 151
rect 18 150 19 151
rect 17 150 18 151
rect 16 150 17 151
rect 78 151 79 152
rect 77 151 78 152
rect 76 151 77 152
rect 75 151 76 152
rect 74 151 75 152
rect 73 151 74 152
rect 72 151 73 152
rect 71 151 72 152
rect 70 151 71 152
rect 69 151 70 152
rect 68 151 69 152
rect 67 151 68 152
rect 66 151 67 152
rect 65 151 66 152
rect 64 151 65 152
rect 63 151 64 152
rect 62 151 63 152
rect 61 151 62 152
rect 60 151 61 152
rect 59 151 60 152
rect 58 151 59 152
rect 57 151 58 152
rect 56 151 57 152
rect 55 151 56 152
rect 54 151 55 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 40 151 41 152
rect 39 151 40 152
rect 38 151 39 152
rect 37 151 38 152
rect 36 151 37 152
rect 35 151 36 152
rect 34 151 35 152
rect 33 151 34 152
rect 32 151 33 152
rect 31 151 32 152
rect 30 151 31 152
rect 29 151 30 152
rect 28 151 29 152
rect 27 151 28 152
rect 26 151 27 152
rect 25 151 26 152
rect 24 151 25 152
rect 23 151 24 152
rect 22 151 23 152
rect 21 151 22 152
rect 20 151 21 152
rect 19 151 20 152
rect 18 151 19 152
rect 17 151 18 152
rect 16 151 17 152
rect 79 152 80 153
rect 78 152 79 153
rect 77 152 78 153
rect 76 152 77 153
rect 75 152 76 153
rect 74 152 75 153
rect 73 152 74 153
rect 72 152 73 153
rect 71 152 72 153
rect 70 152 71 153
rect 69 152 70 153
rect 68 152 69 153
rect 67 152 68 153
rect 66 152 67 153
rect 65 152 66 153
rect 64 152 65 153
rect 63 152 64 153
rect 62 152 63 153
rect 61 152 62 153
rect 60 152 61 153
rect 59 152 60 153
rect 58 152 59 153
rect 57 152 58 153
rect 56 152 57 153
rect 55 152 56 153
rect 54 152 55 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 40 152 41 153
rect 39 152 40 153
rect 38 152 39 153
rect 37 152 38 153
rect 36 152 37 153
rect 35 152 36 153
rect 34 152 35 153
rect 33 152 34 153
rect 32 152 33 153
rect 31 152 32 153
rect 30 152 31 153
rect 29 152 30 153
rect 28 152 29 153
rect 27 152 28 153
rect 26 152 27 153
rect 25 152 26 153
rect 24 152 25 153
rect 23 152 24 153
rect 22 152 23 153
rect 21 152 22 153
rect 20 152 21 153
rect 19 152 20 153
rect 18 152 19 153
rect 17 152 18 153
rect 16 152 17 153
rect 79 153 80 154
rect 78 153 79 154
rect 77 153 78 154
rect 76 153 77 154
rect 75 153 76 154
rect 74 153 75 154
rect 73 153 74 154
rect 72 153 73 154
rect 71 153 72 154
rect 70 153 71 154
rect 69 153 70 154
rect 68 153 69 154
rect 67 153 68 154
rect 66 153 67 154
rect 65 153 66 154
rect 64 153 65 154
rect 63 153 64 154
rect 62 153 63 154
rect 61 153 62 154
rect 60 153 61 154
rect 59 153 60 154
rect 58 153 59 154
rect 57 153 58 154
rect 56 153 57 154
rect 55 153 56 154
rect 54 153 55 154
rect 53 153 54 154
rect 52 153 53 154
rect 51 153 52 154
rect 50 153 51 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 43 153 44 154
rect 42 153 43 154
rect 41 153 42 154
rect 40 153 41 154
rect 39 153 40 154
rect 38 153 39 154
rect 37 153 38 154
rect 36 153 37 154
rect 35 153 36 154
rect 34 153 35 154
rect 33 153 34 154
rect 32 153 33 154
rect 31 153 32 154
rect 30 153 31 154
rect 29 153 30 154
rect 28 153 29 154
rect 27 153 28 154
rect 26 153 27 154
rect 25 153 26 154
rect 24 153 25 154
rect 23 153 24 154
rect 22 153 23 154
rect 21 153 22 154
rect 20 153 21 154
rect 19 153 20 154
rect 18 153 19 154
rect 17 153 18 154
rect 16 153 17 154
rect 80 154 81 155
rect 79 154 80 155
rect 78 154 79 155
rect 77 154 78 155
rect 76 154 77 155
rect 75 154 76 155
rect 74 154 75 155
rect 73 154 74 155
rect 72 154 73 155
rect 71 154 72 155
rect 70 154 71 155
rect 69 154 70 155
rect 68 154 69 155
rect 67 154 68 155
rect 66 154 67 155
rect 65 154 66 155
rect 64 154 65 155
rect 63 154 64 155
rect 62 154 63 155
rect 61 154 62 155
rect 60 154 61 155
rect 59 154 60 155
rect 58 154 59 155
rect 57 154 58 155
rect 56 154 57 155
rect 55 154 56 155
rect 54 154 55 155
rect 53 154 54 155
rect 52 154 53 155
rect 51 154 52 155
rect 50 154 51 155
rect 49 154 50 155
rect 48 154 49 155
rect 47 154 48 155
rect 46 154 47 155
rect 45 154 46 155
rect 44 154 45 155
rect 43 154 44 155
rect 42 154 43 155
rect 41 154 42 155
rect 40 154 41 155
rect 39 154 40 155
rect 38 154 39 155
rect 37 154 38 155
rect 36 154 37 155
rect 35 154 36 155
rect 34 154 35 155
rect 33 154 34 155
rect 32 154 33 155
rect 31 154 32 155
rect 30 154 31 155
rect 29 154 30 155
rect 28 154 29 155
rect 27 154 28 155
rect 26 154 27 155
rect 25 154 26 155
rect 24 154 25 155
rect 23 154 24 155
rect 22 154 23 155
rect 21 154 22 155
rect 20 154 21 155
rect 19 154 20 155
rect 18 154 19 155
rect 17 154 18 155
rect 16 154 17 155
rect 141 155 142 156
rect 140 155 141 156
rect 139 155 140 156
rect 138 155 139 156
rect 137 155 138 156
rect 80 155 81 156
rect 79 155 80 156
rect 78 155 79 156
rect 77 155 78 156
rect 76 155 77 156
rect 75 155 76 156
rect 74 155 75 156
rect 73 155 74 156
rect 72 155 73 156
rect 71 155 72 156
rect 70 155 71 156
rect 69 155 70 156
rect 68 155 69 156
rect 67 155 68 156
rect 66 155 67 156
rect 65 155 66 156
rect 64 155 65 156
rect 63 155 64 156
rect 62 155 63 156
rect 61 155 62 156
rect 60 155 61 156
rect 59 155 60 156
rect 58 155 59 156
rect 57 155 58 156
rect 56 155 57 156
rect 55 155 56 156
rect 54 155 55 156
rect 53 155 54 156
rect 52 155 53 156
rect 51 155 52 156
rect 50 155 51 156
rect 49 155 50 156
rect 48 155 49 156
rect 47 155 48 156
rect 46 155 47 156
rect 45 155 46 156
rect 44 155 45 156
rect 43 155 44 156
rect 42 155 43 156
rect 41 155 42 156
rect 40 155 41 156
rect 39 155 40 156
rect 38 155 39 156
rect 37 155 38 156
rect 36 155 37 156
rect 35 155 36 156
rect 34 155 35 156
rect 33 155 34 156
rect 32 155 33 156
rect 31 155 32 156
rect 30 155 31 156
rect 29 155 30 156
rect 28 155 29 156
rect 27 155 28 156
rect 26 155 27 156
rect 25 155 26 156
rect 24 155 25 156
rect 23 155 24 156
rect 22 155 23 156
rect 21 155 22 156
rect 20 155 21 156
rect 19 155 20 156
rect 18 155 19 156
rect 17 155 18 156
rect 16 155 17 156
rect 142 156 143 157
rect 141 156 142 157
rect 140 156 141 157
rect 139 156 140 157
rect 138 156 139 157
rect 137 156 138 157
rect 136 156 137 157
rect 81 156 82 157
rect 80 156 81 157
rect 79 156 80 157
rect 78 156 79 157
rect 77 156 78 157
rect 76 156 77 157
rect 75 156 76 157
rect 74 156 75 157
rect 73 156 74 157
rect 72 156 73 157
rect 71 156 72 157
rect 70 156 71 157
rect 69 156 70 157
rect 68 156 69 157
rect 67 156 68 157
rect 66 156 67 157
rect 65 156 66 157
rect 64 156 65 157
rect 63 156 64 157
rect 62 156 63 157
rect 61 156 62 157
rect 60 156 61 157
rect 59 156 60 157
rect 58 156 59 157
rect 57 156 58 157
rect 56 156 57 157
rect 55 156 56 157
rect 54 156 55 157
rect 53 156 54 157
rect 52 156 53 157
rect 51 156 52 157
rect 50 156 51 157
rect 49 156 50 157
rect 48 156 49 157
rect 47 156 48 157
rect 46 156 47 157
rect 45 156 46 157
rect 44 156 45 157
rect 43 156 44 157
rect 42 156 43 157
rect 41 156 42 157
rect 40 156 41 157
rect 39 156 40 157
rect 38 156 39 157
rect 37 156 38 157
rect 36 156 37 157
rect 35 156 36 157
rect 34 156 35 157
rect 33 156 34 157
rect 32 156 33 157
rect 31 156 32 157
rect 30 156 31 157
rect 29 156 30 157
rect 28 156 29 157
rect 27 156 28 157
rect 26 156 27 157
rect 25 156 26 157
rect 24 156 25 157
rect 23 156 24 157
rect 22 156 23 157
rect 21 156 22 157
rect 20 156 21 157
rect 19 156 20 157
rect 18 156 19 157
rect 17 156 18 157
rect 16 156 17 157
rect 143 157 144 158
rect 142 157 143 158
rect 141 157 142 158
rect 140 157 141 158
rect 139 157 140 158
rect 138 157 139 158
rect 137 157 138 158
rect 136 157 137 158
rect 135 157 136 158
rect 131 157 132 158
rect 130 157 131 158
rect 129 157 130 158
rect 128 157 129 158
rect 127 157 128 158
rect 81 157 82 158
rect 80 157 81 158
rect 79 157 80 158
rect 78 157 79 158
rect 77 157 78 158
rect 76 157 77 158
rect 75 157 76 158
rect 74 157 75 158
rect 73 157 74 158
rect 72 157 73 158
rect 71 157 72 158
rect 70 157 71 158
rect 69 157 70 158
rect 68 157 69 158
rect 67 157 68 158
rect 66 157 67 158
rect 65 157 66 158
rect 64 157 65 158
rect 63 157 64 158
rect 62 157 63 158
rect 61 157 62 158
rect 60 157 61 158
rect 59 157 60 158
rect 58 157 59 158
rect 57 157 58 158
rect 56 157 57 158
rect 55 157 56 158
rect 54 157 55 158
rect 53 157 54 158
rect 52 157 53 158
rect 51 157 52 158
rect 50 157 51 158
rect 49 157 50 158
rect 48 157 49 158
rect 47 157 48 158
rect 46 157 47 158
rect 45 157 46 158
rect 44 157 45 158
rect 43 157 44 158
rect 42 157 43 158
rect 41 157 42 158
rect 40 157 41 158
rect 39 157 40 158
rect 38 157 39 158
rect 37 157 38 158
rect 36 157 37 158
rect 35 157 36 158
rect 34 157 35 158
rect 33 157 34 158
rect 32 157 33 158
rect 31 157 32 158
rect 30 157 31 158
rect 29 157 30 158
rect 28 157 29 158
rect 27 157 28 158
rect 26 157 27 158
rect 25 157 26 158
rect 24 157 25 158
rect 23 157 24 158
rect 22 157 23 158
rect 21 157 22 158
rect 20 157 21 158
rect 19 157 20 158
rect 18 157 19 158
rect 17 157 18 158
rect 16 157 17 158
rect 144 158 145 159
rect 143 158 144 159
rect 142 158 143 159
rect 141 158 142 159
rect 140 158 141 159
rect 139 158 140 159
rect 138 158 139 159
rect 137 158 138 159
rect 136 158 137 159
rect 135 158 136 159
rect 134 158 135 159
rect 130 158 131 159
rect 129 158 130 159
rect 128 158 129 159
rect 127 158 128 159
rect 82 158 83 159
rect 81 158 82 159
rect 80 158 81 159
rect 79 158 80 159
rect 78 158 79 159
rect 77 158 78 159
rect 76 158 77 159
rect 75 158 76 159
rect 74 158 75 159
rect 73 158 74 159
rect 72 158 73 159
rect 71 158 72 159
rect 70 158 71 159
rect 69 158 70 159
rect 68 158 69 159
rect 67 158 68 159
rect 66 158 67 159
rect 65 158 66 159
rect 64 158 65 159
rect 63 158 64 159
rect 62 158 63 159
rect 61 158 62 159
rect 60 158 61 159
rect 59 158 60 159
rect 58 158 59 159
rect 57 158 58 159
rect 56 158 57 159
rect 55 158 56 159
rect 54 158 55 159
rect 53 158 54 159
rect 52 158 53 159
rect 51 158 52 159
rect 50 158 51 159
rect 49 158 50 159
rect 48 158 49 159
rect 47 158 48 159
rect 46 158 47 159
rect 45 158 46 159
rect 44 158 45 159
rect 43 158 44 159
rect 42 158 43 159
rect 41 158 42 159
rect 40 158 41 159
rect 39 158 40 159
rect 38 158 39 159
rect 37 158 38 159
rect 36 158 37 159
rect 35 158 36 159
rect 34 158 35 159
rect 33 158 34 159
rect 32 158 33 159
rect 31 158 32 159
rect 30 158 31 159
rect 29 158 30 159
rect 28 158 29 159
rect 27 158 28 159
rect 26 158 27 159
rect 25 158 26 159
rect 24 158 25 159
rect 23 158 24 159
rect 22 158 23 159
rect 21 158 22 159
rect 20 158 21 159
rect 19 158 20 159
rect 18 158 19 159
rect 17 158 18 159
rect 16 158 17 159
rect 144 159 145 160
rect 143 159 144 160
rect 142 159 143 160
rect 141 159 142 160
rect 140 159 141 160
rect 139 159 140 160
rect 138 159 139 160
rect 137 159 138 160
rect 136 159 137 160
rect 135 159 136 160
rect 134 159 135 160
rect 130 159 131 160
rect 129 159 130 160
rect 128 159 129 160
rect 127 159 128 160
rect 82 159 83 160
rect 81 159 82 160
rect 80 159 81 160
rect 79 159 80 160
rect 78 159 79 160
rect 77 159 78 160
rect 76 159 77 160
rect 75 159 76 160
rect 74 159 75 160
rect 73 159 74 160
rect 72 159 73 160
rect 71 159 72 160
rect 70 159 71 160
rect 69 159 70 160
rect 68 159 69 160
rect 67 159 68 160
rect 66 159 67 160
rect 65 159 66 160
rect 64 159 65 160
rect 63 159 64 160
rect 62 159 63 160
rect 61 159 62 160
rect 60 159 61 160
rect 59 159 60 160
rect 58 159 59 160
rect 57 159 58 160
rect 56 159 57 160
rect 55 159 56 160
rect 54 159 55 160
rect 53 159 54 160
rect 52 159 53 160
rect 51 159 52 160
rect 50 159 51 160
rect 49 159 50 160
rect 48 159 49 160
rect 47 159 48 160
rect 46 159 47 160
rect 45 159 46 160
rect 44 159 45 160
rect 43 159 44 160
rect 42 159 43 160
rect 41 159 42 160
rect 40 159 41 160
rect 39 159 40 160
rect 38 159 39 160
rect 37 159 38 160
rect 36 159 37 160
rect 35 159 36 160
rect 34 159 35 160
rect 33 159 34 160
rect 32 159 33 160
rect 31 159 32 160
rect 30 159 31 160
rect 29 159 30 160
rect 28 159 29 160
rect 27 159 28 160
rect 26 159 27 160
rect 25 159 26 160
rect 24 159 25 160
rect 23 159 24 160
rect 22 159 23 160
rect 21 159 22 160
rect 20 159 21 160
rect 19 159 20 160
rect 18 159 19 160
rect 17 159 18 160
rect 16 159 17 160
rect 144 160 145 161
rect 143 160 144 161
rect 142 160 143 161
rect 141 160 142 161
rect 140 160 141 161
rect 137 160 138 161
rect 136 160 137 161
rect 135 160 136 161
rect 134 160 135 161
rect 129 160 130 161
rect 128 160 129 161
rect 127 160 128 161
rect 126 160 127 161
rect 82 160 83 161
rect 81 160 82 161
rect 80 160 81 161
rect 79 160 80 161
rect 78 160 79 161
rect 77 160 78 161
rect 76 160 77 161
rect 75 160 76 161
rect 74 160 75 161
rect 73 160 74 161
rect 72 160 73 161
rect 71 160 72 161
rect 70 160 71 161
rect 69 160 70 161
rect 68 160 69 161
rect 67 160 68 161
rect 66 160 67 161
rect 65 160 66 161
rect 64 160 65 161
rect 63 160 64 161
rect 62 160 63 161
rect 61 160 62 161
rect 60 160 61 161
rect 59 160 60 161
rect 58 160 59 161
rect 57 160 58 161
rect 56 160 57 161
rect 55 160 56 161
rect 54 160 55 161
rect 53 160 54 161
rect 52 160 53 161
rect 51 160 52 161
rect 50 160 51 161
rect 49 160 50 161
rect 48 160 49 161
rect 47 160 48 161
rect 46 160 47 161
rect 45 160 46 161
rect 44 160 45 161
rect 43 160 44 161
rect 42 160 43 161
rect 41 160 42 161
rect 40 160 41 161
rect 39 160 40 161
rect 38 160 39 161
rect 37 160 38 161
rect 36 160 37 161
rect 35 160 36 161
rect 34 160 35 161
rect 33 160 34 161
rect 32 160 33 161
rect 31 160 32 161
rect 30 160 31 161
rect 29 160 30 161
rect 28 160 29 161
rect 27 160 28 161
rect 26 160 27 161
rect 25 160 26 161
rect 24 160 25 161
rect 23 160 24 161
rect 22 160 23 161
rect 21 160 22 161
rect 20 160 21 161
rect 19 160 20 161
rect 18 160 19 161
rect 17 160 18 161
rect 16 160 17 161
rect 144 161 145 162
rect 143 161 144 162
rect 142 161 143 162
rect 141 161 142 162
rect 136 161 137 162
rect 135 161 136 162
rect 134 161 135 162
rect 133 161 134 162
rect 129 161 130 162
rect 128 161 129 162
rect 127 161 128 162
rect 126 161 127 162
rect 82 161 83 162
rect 81 161 82 162
rect 80 161 81 162
rect 79 161 80 162
rect 78 161 79 162
rect 77 161 78 162
rect 76 161 77 162
rect 75 161 76 162
rect 74 161 75 162
rect 73 161 74 162
rect 72 161 73 162
rect 71 161 72 162
rect 70 161 71 162
rect 69 161 70 162
rect 68 161 69 162
rect 67 161 68 162
rect 66 161 67 162
rect 65 161 66 162
rect 64 161 65 162
rect 63 161 64 162
rect 62 161 63 162
rect 61 161 62 162
rect 60 161 61 162
rect 144 162 145 163
rect 143 162 144 163
rect 142 162 143 163
rect 141 162 142 163
rect 135 162 136 163
rect 134 162 135 163
rect 133 162 134 163
rect 129 162 130 163
rect 128 162 129 163
rect 127 162 128 163
rect 126 162 127 163
rect 82 162 83 163
rect 81 162 82 163
rect 80 162 81 163
rect 79 162 80 163
rect 78 162 79 163
rect 77 162 78 163
rect 76 162 77 163
rect 75 162 76 163
rect 74 162 75 163
rect 73 162 74 163
rect 72 162 73 163
rect 71 162 72 163
rect 70 162 71 163
rect 69 162 70 163
rect 68 162 69 163
rect 67 162 68 163
rect 66 162 67 163
rect 65 162 66 163
rect 64 162 65 163
rect 63 162 64 163
rect 143 163 144 164
rect 142 163 143 164
rect 141 163 142 164
rect 135 163 136 164
rect 134 163 135 164
rect 133 163 134 164
rect 129 163 130 164
rect 128 163 129 164
rect 127 163 128 164
rect 126 163 127 164
rect 83 163 84 164
rect 82 163 83 164
rect 81 163 82 164
rect 80 163 81 164
rect 79 163 80 164
rect 78 163 79 164
rect 77 163 78 164
rect 76 163 77 164
rect 75 163 76 164
rect 74 163 75 164
rect 73 163 74 164
rect 72 163 73 164
rect 71 163 72 164
rect 70 163 71 164
rect 69 163 70 164
rect 68 163 69 164
rect 67 163 68 164
rect 66 163 67 164
rect 65 163 66 164
rect 64 163 65 164
rect 143 164 144 165
rect 142 164 143 165
rect 141 164 142 165
rect 135 164 136 165
rect 134 164 135 165
rect 133 164 134 165
rect 129 164 130 165
rect 128 164 129 165
rect 127 164 128 165
rect 126 164 127 165
rect 83 164 84 165
rect 82 164 83 165
rect 81 164 82 165
rect 80 164 81 165
rect 79 164 80 165
rect 78 164 79 165
rect 77 164 78 165
rect 76 164 77 165
rect 75 164 76 165
rect 74 164 75 165
rect 73 164 74 165
rect 72 164 73 165
rect 71 164 72 165
rect 70 164 71 165
rect 69 164 70 165
rect 68 164 69 165
rect 67 164 68 165
rect 66 164 67 165
rect 65 164 66 165
rect 142 165 143 166
rect 141 165 142 166
rect 140 165 141 166
rect 135 165 136 166
rect 134 165 135 166
rect 133 165 134 166
rect 129 165 130 166
rect 128 165 129 166
rect 127 165 128 166
rect 126 165 127 166
rect 83 165 84 166
rect 82 165 83 166
rect 81 165 82 166
rect 80 165 81 166
rect 79 165 80 166
rect 78 165 79 166
rect 77 165 78 166
rect 76 165 77 166
rect 75 165 76 166
rect 74 165 75 166
rect 73 165 74 166
rect 72 165 73 166
rect 71 165 72 166
rect 70 165 71 166
rect 69 165 70 166
rect 68 165 69 166
rect 67 165 68 166
rect 66 165 67 166
rect 142 166 143 167
rect 141 166 142 167
rect 140 166 141 167
rect 139 166 140 167
rect 138 166 139 167
rect 135 166 136 167
rect 134 166 135 167
rect 133 166 134 167
rect 132 166 133 167
rect 131 166 132 167
rect 130 166 131 167
rect 129 166 130 167
rect 128 166 129 167
rect 127 166 128 167
rect 126 166 127 167
rect 83 166 84 167
rect 82 166 83 167
rect 81 166 82 167
rect 80 166 81 167
rect 79 166 80 167
rect 78 166 79 167
rect 77 166 78 167
rect 76 166 77 167
rect 75 166 76 167
rect 74 166 75 167
rect 73 166 74 167
rect 72 166 73 167
rect 71 166 72 167
rect 70 166 71 167
rect 69 166 70 167
rect 68 166 69 167
rect 67 166 68 167
rect 66 166 67 167
rect 144 167 145 168
rect 143 167 144 168
rect 142 167 143 168
rect 141 167 142 168
rect 140 167 141 168
rect 139 167 140 168
rect 138 167 139 168
rect 137 167 138 168
rect 136 167 137 168
rect 135 167 136 168
rect 134 167 135 168
rect 133 167 134 168
rect 132 167 133 168
rect 131 167 132 168
rect 130 167 131 168
rect 129 167 130 168
rect 128 167 129 168
rect 127 167 128 168
rect 83 167 84 168
rect 82 167 83 168
rect 81 167 82 168
rect 80 167 81 168
rect 79 167 80 168
rect 78 167 79 168
rect 77 167 78 168
rect 76 167 77 168
rect 75 167 76 168
rect 74 167 75 168
rect 73 167 74 168
rect 72 167 73 168
rect 71 167 72 168
rect 70 167 71 168
rect 69 167 70 168
rect 68 167 69 168
rect 67 167 68 168
rect 144 168 145 169
rect 143 168 144 169
rect 142 168 143 169
rect 141 168 142 169
rect 140 168 141 169
rect 139 168 140 169
rect 138 168 139 169
rect 137 168 138 169
rect 136 168 137 169
rect 135 168 136 169
rect 134 168 135 169
rect 133 168 134 169
rect 132 168 133 169
rect 131 168 132 169
rect 130 168 131 169
rect 129 168 130 169
rect 128 168 129 169
rect 127 168 128 169
rect 83 168 84 169
rect 82 168 83 169
rect 81 168 82 169
rect 80 168 81 169
rect 79 168 80 169
rect 78 168 79 169
rect 77 168 78 169
rect 76 168 77 169
rect 75 168 76 169
rect 74 168 75 169
rect 73 168 74 169
rect 72 168 73 169
rect 71 168 72 169
rect 70 168 71 169
rect 69 168 70 169
rect 68 168 69 169
rect 67 168 68 169
rect 144 169 145 170
rect 143 169 144 170
rect 142 169 143 170
rect 141 169 142 170
rect 140 169 141 170
rect 139 169 140 170
rect 138 169 139 170
rect 137 169 138 170
rect 136 169 137 170
rect 135 169 136 170
rect 134 169 135 170
rect 133 169 134 170
rect 132 169 133 170
rect 131 169 132 170
rect 130 169 131 170
rect 129 169 130 170
rect 128 169 129 170
rect 83 169 84 170
rect 82 169 83 170
rect 81 169 82 170
rect 80 169 81 170
rect 79 169 80 170
rect 78 169 79 170
rect 77 169 78 170
rect 76 169 77 170
rect 75 169 76 170
rect 74 169 75 170
rect 73 169 74 170
rect 72 169 73 170
rect 71 169 72 170
rect 70 169 71 170
rect 69 169 70 170
rect 68 169 69 170
rect 67 169 68 170
rect 144 170 145 171
rect 143 170 144 171
rect 142 170 143 171
rect 141 170 142 171
rect 140 170 141 171
rect 139 170 140 171
rect 138 170 139 171
rect 137 170 138 171
rect 136 170 137 171
rect 135 170 136 171
rect 134 170 135 171
rect 133 170 134 171
rect 132 170 133 171
rect 131 170 132 171
rect 130 170 131 171
rect 129 170 130 171
rect 83 170 84 171
rect 82 170 83 171
rect 81 170 82 171
rect 80 170 81 171
rect 79 170 80 171
rect 78 170 79 171
rect 77 170 78 171
rect 76 170 77 171
rect 75 170 76 171
rect 74 170 75 171
rect 73 170 74 171
rect 72 170 73 171
rect 71 170 72 171
rect 70 170 71 171
rect 69 170 70 171
rect 68 170 69 171
rect 67 170 68 171
rect 144 171 145 172
rect 143 171 144 172
rect 142 171 143 172
rect 141 171 142 172
rect 140 171 141 172
rect 139 171 140 172
rect 138 171 139 172
rect 137 171 138 172
rect 136 171 137 172
rect 135 171 136 172
rect 134 171 135 172
rect 133 171 134 172
rect 132 171 133 172
rect 131 171 132 172
rect 83 171 84 172
rect 82 171 83 172
rect 81 171 82 172
rect 80 171 81 172
rect 79 171 80 172
rect 78 171 79 172
rect 77 171 78 172
rect 76 171 77 172
rect 75 171 76 172
rect 74 171 75 172
rect 73 171 74 172
rect 72 171 73 172
rect 71 171 72 172
rect 70 171 71 172
rect 69 171 70 172
rect 68 171 69 172
rect 67 171 68 172
rect 83 172 84 173
rect 82 172 83 173
rect 81 172 82 173
rect 80 172 81 173
rect 79 172 80 173
rect 78 172 79 173
rect 77 172 78 173
rect 76 172 77 173
rect 75 172 76 173
rect 74 172 75 173
rect 73 172 74 173
rect 72 172 73 173
rect 71 172 72 173
rect 70 172 71 173
rect 69 172 70 173
rect 68 172 69 173
rect 67 172 68 173
rect 83 173 84 174
rect 82 173 83 174
rect 81 173 82 174
rect 80 173 81 174
rect 79 173 80 174
rect 78 173 79 174
rect 77 173 78 174
rect 76 173 77 174
rect 75 173 76 174
rect 74 173 75 174
rect 73 173 74 174
rect 72 173 73 174
rect 71 173 72 174
rect 70 173 71 174
rect 69 173 70 174
rect 68 173 69 174
rect 67 173 68 174
rect 66 173 67 174
rect 83 174 84 175
rect 82 174 83 175
rect 81 174 82 175
rect 80 174 81 175
rect 79 174 80 175
rect 78 174 79 175
rect 77 174 78 175
rect 76 174 77 175
rect 75 174 76 175
rect 74 174 75 175
rect 73 174 74 175
rect 72 174 73 175
rect 71 174 72 175
rect 70 174 71 175
rect 69 174 70 175
rect 68 174 69 175
rect 67 174 68 175
rect 66 174 67 175
rect 83 175 84 176
rect 82 175 83 176
rect 81 175 82 176
rect 80 175 81 176
rect 79 175 80 176
rect 78 175 79 176
rect 77 175 78 176
rect 76 175 77 176
rect 75 175 76 176
rect 74 175 75 176
rect 73 175 74 176
rect 72 175 73 176
rect 71 175 72 176
rect 70 175 71 176
rect 69 175 70 176
rect 68 175 69 176
rect 67 175 68 176
rect 66 175 67 176
rect 65 175 66 176
rect 82 176 83 177
rect 81 176 82 177
rect 80 176 81 177
rect 79 176 80 177
rect 78 176 79 177
rect 77 176 78 177
rect 76 176 77 177
rect 75 176 76 177
rect 74 176 75 177
rect 73 176 74 177
rect 72 176 73 177
rect 71 176 72 177
rect 70 176 71 177
rect 69 176 70 177
rect 68 176 69 177
rect 67 176 68 177
rect 66 176 67 177
rect 65 176 66 177
rect 64 176 65 177
rect 144 177 145 178
rect 143 177 144 178
rect 142 177 143 178
rect 141 177 142 178
rect 140 177 141 178
rect 139 177 140 178
rect 138 177 139 178
rect 137 177 138 178
rect 136 177 137 178
rect 135 177 136 178
rect 134 177 135 178
rect 133 177 134 178
rect 132 177 133 178
rect 131 177 132 178
rect 130 177 131 178
rect 129 177 130 178
rect 128 177 129 178
rect 127 177 128 178
rect 126 177 127 178
rect 82 177 83 178
rect 81 177 82 178
rect 80 177 81 178
rect 79 177 80 178
rect 78 177 79 178
rect 77 177 78 178
rect 76 177 77 178
rect 75 177 76 178
rect 74 177 75 178
rect 73 177 74 178
rect 72 177 73 178
rect 71 177 72 178
rect 70 177 71 178
rect 69 177 70 178
rect 68 177 69 178
rect 67 177 68 178
rect 66 177 67 178
rect 65 177 66 178
rect 64 177 65 178
rect 63 177 64 178
rect 144 178 145 179
rect 143 178 144 179
rect 142 178 143 179
rect 141 178 142 179
rect 140 178 141 179
rect 139 178 140 179
rect 138 178 139 179
rect 137 178 138 179
rect 136 178 137 179
rect 135 178 136 179
rect 134 178 135 179
rect 133 178 134 179
rect 132 178 133 179
rect 131 178 132 179
rect 130 178 131 179
rect 129 178 130 179
rect 128 178 129 179
rect 127 178 128 179
rect 126 178 127 179
rect 82 178 83 179
rect 81 178 82 179
rect 80 178 81 179
rect 79 178 80 179
rect 78 178 79 179
rect 77 178 78 179
rect 76 178 77 179
rect 75 178 76 179
rect 74 178 75 179
rect 73 178 74 179
rect 72 178 73 179
rect 71 178 72 179
rect 70 178 71 179
rect 69 178 70 179
rect 68 178 69 179
rect 67 178 68 179
rect 66 178 67 179
rect 65 178 66 179
rect 64 178 65 179
rect 63 178 64 179
rect 62 178 63 179
rect 61 178 62 179
rect 60 178 61 179
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 127 179 128 180
rect 126 179 127 180
rect 82 179 83 180
rect 81 179 82 180
rect 80 179 81 180
rect 79 179 80 180
rect 78 179 79 180
rect 77 179 78 180
rect 76 179 77 180
rect 75 179 76 180
rect 74 179 75 180
rect 73 179 74 180
rect 72 179 73 180
rect 71 179 72 180
rect 70 179 71 180
rect 69 179 70 180
rect 68 179 69 180
rect 67 179 68 180
rect 66 179 67 180
rect 65 179 66 180
rect 64 179 65 180
rect 63 179 64 180
rect 62 179 63 180
rect 61 179 62 180
rect 60 179 61 180
rect 59 179 60 180
rect 58 179 59 180
rect 57 179 58 180
rect 56 179 57 180
rect 55 179 56 180
rect 54 179 55 180
rect 53 179 54 180
rect 52 179 53 180
rect 51 179 52 180
rect 50 179 51 180
rect 49 179 50 180
rect 48 179 49 180
rect 47 179 48 180
rect 46 179 47 180
rect 45 179 46 180
rect 44 179 45 180
rect 43 179 44 180
rect 42 179 43 180
rect 41 179 42 180
rect 40 179 41 180
rect 39 179 40 180
rect 38 179 39 180
rect 37 179 38 180
rect 36 179 37 180
rect 35 179 36 180
rect 34 179 35 180
rect 33 179 34 180
rect 32 179 33 180
rect 31 179 32 180
rect 30 179 31 180
rect 29 179 30 180
rect 28 179 29 180
rect 27 179 28 180
rect 26 179 27 180
rect 25 179 26 180
rect 24 179 25 180
rect 23 179 24 180
rect 22 179 23 180
rect 21 179 22 180
rect 20 179 21 180
rect 19 179 20 180
rect 18 179 19 180
rect 17 179 18 180
rect 16 179 17 180
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 127 180 128 181
rect 126 180 127 181
rect 82 180 83 181
rect 81 180 82 181
rect 80 180 81 181
rect 79 180 80 181
rect 78 180 79 181
rect 77 180 78 181
rect 76 180 77 181
rect 75 180 76 181
rect 74 180 75 181
rect 73 180 74 181
rect 72 180 73 181
rect 71 180 72 181
rect 70 180 71 181
rect 69 180 70 181
rect 68 180 69 181
rect 67 180 68 181
rect 66 180 67 181
rect 65 180 66 181
rect 64 180 65 181
rect 63 180 64 181
rect 62 180 63 181
rect 61 180 62 181
rect 60 180 61 181
rect 59 180 60 181
rect 58 180 59 181
rect 57 180 58 181
rect 56 180 57 181
rect 55 180 56 181
rect 54 180 55 181
rect 53 180 54 181
rect 52 180 53 181
rect 51 180 52 181
rect 50 180 51 181
rect 49 180 50 181
rect 48 180 49 181
rect 47 180 48 181
rect 46 180 47 181
rect 45 180 46 181
rect 44 180 45 181
rect 43 180 44 181
rect 42 180 43 181
rect 41 180 42 181
rect 40 180 41 181
rect 39 180 40 181
rect 38 180 39 181
rect 37 180 38 181
rect 36 180 37 181
rect 35 180 36 181
rect 34 180 35 181
rect 33 180 34 181
rect 32 180 33 181
rect 31 180 32 181
rect 30 180 31 181
rect 29 180 30 181
rect 28 180 29 181
rect 27 180 28 181
rect 26 180 27 181
rect 25 180 26 181
rect 24 180 25 181
rect 23 180 24 181
rect 22 180 23 181
rect 21 180 22 181
rect 20 180 21 181
rect 19 180 20 181
rect 18 180 19 181
rect 17 180 18 181
rect 16 180 17 181
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 127 181 128 182
rect 126 181 127 182
rect 81 181 82 182
rect 80 181 81 182
rect 79 181 80 182
rect 78 181 79 182
rect 77 181 78 182
rect 76 181 77 182
rect 75 181 76 182
rect 74 181 75 182
rect 73 181 74 182
rect 72 181 73 182
rect 71 181 72 182
rect 70 181 71 182
rect 69 181 70 182
rect 68 181 69 182
rect 67 181 68 182
rect 66 181 67 182
rect 65 181 66 182
rect 64 181 65 182
rect 63 181 64 182
rect 62 181 63 182
rect 61 181 62 182
rect 60 181 61 182
rect 59 181 60 182
rect 58 181 59 182
rect 57 181 58 182
rect 56 181 57 182
rect 55 181 56 182
rect 54 181 55 182
rect 53 181 54 182
rect 52 181 53 182
rect 51 181 52 182
rect 50 181 51 182
rect 49 181 50 182
rect 48 181 49 182
rect 47 181 48 182
rect 46 181 47 182
rect 45 181 46 182
rect 44 181 45 182
rect 43 181 44 182
rect 42 181 43 182
rect 41 181 42 182
rect 40 181 41 182
rect 39 181 40 182
rect 38 181 39 182
rect 37 181 38 182
rect 36 181 37 182
rect 35 181 36 182
rect 34 181 35 182
rect 33 181 34 182
rect 32 181 33 182
rect 31 181 32 182
rect 30 181 31 182
rect 29 181 30 182
rect 28 181 29 182
rect 27 181 28 182
rect 26 181 27 182
rect 25 181 26 182
rect 24 181 25 182
rect 23 181 24 182
rect 22 181 23 182
rect 21 181 22 182
rect 20 181 21 182
rect 19 181 20 182
rect 18 181 19 182
rect 17 181 18 182
rect 16 181 17 182
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 81 182 82 183
rect 80 182 81 183
rect 79 182 80 183
rect 78 182 79 183
rect 77 182 78 183
rect 76 182 77 183
rect 75 182 76 183
rect 74 182 75 183
rect 73 182 74 183
rect 72 182 73 183
rect 71 182 72 183
rect 70 182 71 183
rect 69 182 70 183
rect 68 182 69 183
rect 67 182 68 183
rect 66 182 67 183
rect 65 182 66 183
rect 64 182 65 183
rect 63 182 64 183
rect 62 182 63 183
rect 61 182 62 183
rect 60 182 61 183
rect 59 182 60 183
rect 58 182 59 183
rect 57 182 58 183
rect 56 182 57 183
rect 55 182 56 183
rect 54 182 55 183
rect 53 182 54 183
rect 52 182 53 183
rect 51 182 52 183
rect 50 182 51 183
rect 49 182 50 183
rect 48 182 49 183
rect 47 182 48 183
rect 46 182 47 183
rect 45 182 46 183
rect 44 182 45 183
rect 43 182 44 183
rect 42 182 43 183
rect 41 182 42 183
rect 40 182 41 183
rect 39 182 40 183
rect 38 182 39 183
rect 37 182 38 183
rect 36 182 37 183
rect 35 182 36 183
rect 34 182 35 183
rect 33 182 34 183
rect 32 182 33 183
rect 31 182 32 183
rect 30 182 31 183
rect 29 182 30 183
rect 28 182 29 183
rect 27 182 28 183
rect 26 182 27 183
rect 25 182 26 183
rect 24 182 25 183
rect 23 182 24 183
rect 22 182 23 183
rect 21 182 22 183
rect 20 182 21 183
rect 19 182 20 183
rect 18 182 19 183
rect 17 182 18 183
rect 16 182 17 183
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 81 183 82 184
rect 80 183 81 184
rect 79 183 80 184
rect 78 183 79 184
rect 77 183 78 184
rect 76 183 77 184
rect 75 183 76 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 70 183 71 184
rect 69 183 70 184
rect 68 183 69 184
rect 67 183 68 184
rect 66 183 67 184
rect 65 183 66 184
rect 64 183 65 184
rect 63 183 64 184
rect 62 183 63 184
rect 61 183 62 184
rect 60 183 61 184
rect 59 183 60 184
rect 58 183 59 184
rect 57 183 58 184
rect 56 183 57 184
rect 55 183 56 184
rect 54 183 55 184
rect 53 183 54 184
rect 52 183 53 184
rect 51 183 52 184
rect 50 183 51 184
rect 49 183 50 184
rect 48 183 49 184
rect 47 183 48 184
rect 46 183 47 184
rect 45 183 46 184
rect 44 183 45 184
rect 43 183 44 184
rect 42 183 43 184
rect 41 183 42 184
rect 40 183 41 184
rect 39 183 40 184
rect 38 183 39 184
rect 37 183 38 184
rect 36 183 37 184
rect 35 183 36 184
rect 34 183 35 184
rect 33 183 34 184
rect 32 183 33 184
rect 31 183 32 184
rect 30 183 31 184
rect 29 183 30 184
rect 28 183 29 184
rect 27 183 28 184
rect 26 183 27 184
rect 25 183 26 184
rect 24 183 25 184
rect 23 183 24 184
rect 22 183 23 184
rect 21 183 22 184
rect 20 183 21 184
rect 19 183 20 184
rect 18 183 19 184
rect 17 183 18 184
rect 16 183 17 184
rect 130 184 131 185
rect 129 184 130 185
rect 128 184 129 185
rect 127 184 128 185
rect 80 184 81 185
rect 79 184 80 185
rect 78 184 79 185
rect 77 184 78 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 70 184 71 185
rect 69 184 70 185
rect 68 184 69 185
rect 67 184 68 185
rect 66 184 67 185
rect 65 184 66 185
rect 64 184 65 185
rect 63 184 64 185
rect 62 184 63 185
rect 61 184 62 185
rect 60 184 61 185
rect 59 184 60 185
rect 58 184 59 185
rect 57 184 58 185
rect 56 184 57 185
rect 55 184 56 185
rect 54 184 55 185
rect 53 184 54 185
rect 52 184 53 185
rect 51 184 52 185
rect 50 184 51 185
rect 49 184 50 185
rect 48 184 49 185
rect 47 184 48 185
rect 46 184 47 185
rect 45 184 46 185
rect 44 184 45 185
rect 43 184 44 185
rect 42 184 43 185
rect 41 184 42 185
rect 40 184 41 185
rect 39 184 40 185
rect 38 184 39 185
rect 37 184 38 185
rect 36 184 37 185
rect 35 184 36 185
rect 34 184 35 185
rect 33 184 34 185
rect 32 184 33 185
rect 31 184 32 185
rect 30 184 31 185
rect 29 184 30 185
rect 28 184 29 185
rect 27 184 28 185
rect 26 184 27 185
rect 25 184 26 185
rect 24 184 25 185
rect 23 184 24 185
rect 22 184 23 185
rect 21 184 22 185
rect 20 184 21 185
rect 19 184 20 185
rect 18 184 19 185
rect 17 184 18 185
rect 16 184 17 185
rect 129 185 130 186
rect 128 185 129 186
rect 127 185 128 186
rect 80 185 81 186
rect 79 185 80 186
rect 78 185 79 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 69 185 70 186
rect 68 185 69 186
rect 67 185 68 186
rect 66 185 67 186
rect 65 185 66 186
rect 64 185 65 186
rect 63 185 64 186
rect 62 185 63 186
rect 61 185 62 186
rect 60 185 61 186
rect 59 185 60 186
rect 58 185 59 186
rect 57 185 58 186
rect 56 185 57 186
rect 55 185 56 186
rect 54 185 55 186
rect 53 185 54 186
rect 52 185 53 186
rect 51 185 52 186
rect 50 185 51 186
rect 49 185 50 186
rect 48 185 49 186
rect 47 185 48 186
rect 46 185 47 186
rect 45 185 46 186
rect 44 185 45 186
rect 43 185 44 186
rect 42 185 43 186
rect 41 185 42 186
rect 40 185 41 186
rect 39 185 40 186
rect 38 185 39 186
rect 37 185 38 186
rect 36 185 37 186
rect 35 185 36 186
rect 34 185 35 186
rect 33 185 34 186
rect 32 185 33 186
rect 31 185 32 186
rect 30 185 31 186
rect 29 185 30 186
rect 28 185 29 186
rect 27 185 28 186
rect 26 185 27 186
rect 25 185 26 186
rect 24 185 25 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 20 185 21 186
rect 19 185 20 186
rect 18 185 19 186
rect 17 185 18 186
rect 16 185 17 186
rect 130 186 131 187
rect 129 186 130 187
rect 128 186 129 187
rect 127 186 128 187
rect 126 186 127 187
rect 79 186 80 187
rect 78 186 79 187
rect 77 186 78 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 69 186 70 187
rect 68 186 69 187
rect 67 186 68 187
rect 66 186 67 187
rect 65 186 66 187
rect 64 186 65 187
rect 63 186 64 187
rect 62 186 63 187
rect 61 186 62 187
rect 60 186 61 187
rect 59 186 60 187
rect 58 186 59 187
rect 57 186 58 187
rect 56 186 57 187
rect 55 186 56 187
rect 54 186 55 187
rect 53 186 54 187
rect 52 186 53 187
rect 51 186 52 187
rect 50 186 51 187
rect 49 186 50 187
rect 48 186 49 187
rect 47 186 48 187
rect 46 186 47 187
rect 45 186 46 187
rect 44 186 45 187
rect 43 186 44 187
rect 42 186 43 187
rect 41 186 42 187
rect 40 186 41 187
rect 39 186 40 187
rect 38 186 39 187
rect 37 186 38 187
rect 36 186 37 187
rect 35 186 36 187
rect 34 186 35 187
rect 33 186 34 187
rect 32 186 33 187
rect 31 186 32 187
rect 30 186 31 187
rect 29 186 30 187
rect 28 186 29 187
rect 27 186 28 187
rect 26 186 27 187
rect 25 186 26 187
rect 24 186 25 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 19 186 20 187
rect 18 186 19 187
rect 17 186 18 187
rect 16 186 17 187
rect 130 187 131 188
rect 129 187 130 188
rect 128 187 129 188
rect 127 187 128 188
rect 126 187 127 188
rect 79 187 80 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 67 187 68 188
rect 66 187 67 188
rect 65 187 66 188
rect 64 187 65 188
rect 63 187 64 188
rect 62 187 63 188
rect 61 187 62 188
rect 60 187 61 188
rect 59 187 60 188
rect 58 187 59 188
rect 57 187 58 188
rect 56 187 57 188
rect 55 187 56 188
rect 54 187 55 188
rect 53 187 54 188
rect 52 187 53 188
rect 51 187 52 188
rect 50 187 51 188
rect 49 187 50 188
rect 48 187 49 188
rect 47 187 48 188
rect 46 187 47 188
rect 45 187 46 188
rect 44 187 45 188
rect 43 187 44 188
rect 42 187 43 188
rect 41 187 42 188
rect 40 187 41 188
rect 39 187 40 188
rect 38 187 39 188
rect 37 187 38 188
rect 36 187 37 188
rect 35 187 36 188
rect 34 187 35 188
rect 33 187 34 188
rect 32 187 33 188
rect 31 187 32 188
rect 30 187 31 188
rect 29 187 30 188
rect 28 187 29 188
rect 27 187 28 188
rect 26 187 27 188
rect 25 187 26 188
rect 24 187 25 188
rect 23 187 24 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 18 187 19 188
rect 17 187 18 188
rect 16 187 17 188
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 127 188 128 189
rect 126 188 127 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 66 188 67 189
rect 65 188 66 189
rect 64 188 65 189
rect 63 188 64 189
rect 62 188 63 189
rect 61 188 62 189
rect 60 188 61 189
rect 59 188 60 189
rect 58 188 59 189
rect 57 188 58 189
rect 56 188 57 189
rect 55 188 56 189
rect 54 188 55 189
rect 53 188 54 189
rect 52 188 53 189
rect 51 188 52 189
rect 50 188 51 189
rect 49 188 50 189
rect 48 188 49 189
rect 47 188 48 189
rect 46 188 47 189
rect 45 188 46 189
rect 44 188 45 189
rect 43 188 44 189
rect 42 188 43 189
rect 41 188 42 189
rect 40 188 41 189
rect 39 188 40 189
rect 38 188 39 189
rect 37 188 38 189
rect 36 188 37 189
rect 35 188 36 189
rect 34 188 35 189
rect 33 188 34 189
rect 32 188 33 189
rect 31 188 32 189
rect 30 188 31 189
rect 29 188 30 189
rect 28 188 29 189
rect 27 188 28 189
rect 26 188 27 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 17 188 18 189
rect 16 188 17 189
rect 144 189 145 190
rect 143 189 144 190
rect 142 189 143 190
rect 141 189 142 190
rect 140 189 141 190
rect 139 189 140 190
rect 138 189 139 190
rect 137 189 138 190
rect 136 189 137 190
rect 135 189 136 190
rect 134 189 135 190
rect 133 189 134 190
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 127 189 128 190
rect 126 189 127 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 69 189 70 190
rect 68 189 69 190
rect 67 189 68 190
rect 66 189 67 190
rect 65 189 66 190
rect 64 189 65 190
rect 63 189 64 190
rect 62 189 63 190
rect 61 189 62 190
rect 60 189 61 190
rect 59 189 60 190
rect 58 189 59 190
rect 57 189 58 190
rect 56 189 57 190
rect 55 189 56 190
rect 54 189 55 190
rect 53 189 54 190
rect 52 189 53 190
rect 51 189 52 190
rect 50 189 51 190
rect 49 189 50 190
rect 48 189 49 190
rect 47 189 48 190
rect 46 189 47 190
rect 45 189 46 190
rect 44 189 45 190
rect 43 189 44 190
rect 42 189 43 190
rect 41 189 42 190
rect 40 189 41 190
rect 39 189 40 190
rect 38 189 39 190
rect 37 189 38 190
rect 36 189 37 190
rect 35 189 36 190
rect 34 189 35 190
rect 33 189 34 190
rect 32 189 33 190
rect 31 189 32 190
rect 30 189 31 190
rect 29 189 30 190
rect 28 189 29 190
rect 27 189 28 190
rect 26 189 27 190
rect 25 189 26 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 17 189 18 190
rect 16 189 17 190
rect 144 190 145 191
rect 143 190 144 191
rect 142 190 143 191
rect 141 190 142 191
rect 140 190 141 191
rect 139 190 140 191
rect 138 190 139 191
rect 137 190 138 191
rect 136 190 137 191
rect 135 190 136 191
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 127 190 128 191
rect 126 190 127 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 68 190 69 191
rect 67 190 68 191
rect 66 190 67 191
rect 65 190 66 191
rect 64 190 65 191
rect 63 190 64 191
rect 62 190 63 191
rect 61 190 62 191
rect 60 190 61 191
rect 59 190 60 191
rect 58 190 59 191
rect 57 190 58 191
rect 56 190 57 191
rect 55 190 56 191
rect 54 190 55 191
rect 53 190 54 191
rect 52 190 53 191
rect 51 190 52 191
rect 50 190 51 191
rect 49 190 50 191
rect 48 190 49 191
rect 47 190 48 191
rect 46 190 47 191
rect 45 190 46 191
rect 44 190 45 191
rect 43 190 44 191
rect 42 190 43 191
rect 41 190 42 191
rect 40 190 41 191
rect 39 190 40 191
rect 38 190 39 191
rect 37 190 38 191
rect 36 190 37 191
rect 35 190 36 191
rect 34 190 35 191
rect 33 190 34 191
rect 32 190 33 191
rect 31 190 32 191
rect 30 190 31 191
rect 29 190 30 191
rect 28 190 29 191
rect 27 190 28 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 19 190 20 191
rect 18 190 19 191
rect 17 190 18 191
rect 16 190 17 191
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 127 191 128 192
rect 76 191 77 192
rect 75 191 76 192
rect 74 191 75 192
rect 73 191 74 192
rect 72 191 73 192
rect 71 191 72 192
rect 70 191 71 192
rect 69 191 70 192
rect 68 191 69 192
rect 67 191 68 192
rect 66 191 67 192
rect 65 191 66 192
rect 64 191 65 192
rect 63 191 64 192
rect 62 191 63 192
rect 61 191 62 192
rect 60 191 61 192
rect 59 191 60 192
rect 58 191 59 192
rect 57 191 58 192
rect 56 191 57 192
rect 55 191 56 192
rect 54 191 55 192
rect 53 191 54 192
rect 52 191 53 192
rect 51 191 52 192
rect 50 191 51 192
rect 49 191 50 192
rect 48 191 49 192
rect 47 191 48 192
rect 46 191 47 192
rect 45 191 46 192
rect 44 191 45 192
rect 43 191 44 192
rect 42 191 43 192
rect 41 191 42 192
rect 40 191 41 192
rect 39 191 40 192
rect 38 191 39 192
rect 37 191 38 192
rect 36 191 37 192
rect 35 191 36 192
rect 34 191 35 192
rect 33 191 34 192
rect 32 191 33 192
rect 31 191 32 192
rect 30 191 31 192
rect 29 191 30 192
rect 28 191 29 192
rect 27 191 28 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 17 191 18 192
rect 16 191 17 192
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 75 192 76 193
rect 74 192 75 193
rect 73 192 74 193
rect 72 192 73 193
rect 71 192 72 193
rect 70 192 71 193
rect 69 192 70 193
rect 68 192 69 193
rect 67 192 68 193
rect 66 192 67 193
rect 65 192 66 193
rect 64 192 65 193
rect 63 192 64 193
rect 62 192 63 193
rect 61 192 62 193
rect 60 192 61 193
rect 59 192 60 193
rect 58 192 59 193
rect 57 192 58 193
rect 56 192 57 193
rect 55 192 56 193
rect 54 192 55 193
rect 53 192 54 193
rect 52 192 53 193
rect 51 192 52 193
rect 50 192 51 193
rect 49 192 50 193
rect 48 192 49 193
rect 47 192 48 193
rect 46 192 47 193
rect 45 192 46 193
rect 44 192 45 193
rect 43 192 44 193
rect 42 192 43 193
rect 41 192 42 193
rect 40 192 41 193
rect 39 192 40 193
rect 38 192 39 193
rect 37 192 38 193
rect 36 192 37 193
rect 35 192 36 193
rect 34 192 35 193
rect 33 192 34 193
rect 32 192 33 193
rect 31 192 32 193
rect 30 192 31 193
rect 29 192 30 193
rect 28 192 29 193
rect 27 192 28 193
rect 26 192 27 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 17 192 18 193
rect 16 192 17 193
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 74 193 75 194
rect 73 193 74 194
rect 72 193 73 194
rect 71 193 72 194
rect 70 193 71 194
rect 69 193 70 194
rect 68 193 69 194
rect 67 193 68 194
rect 66 193 67 194
rect 65 193 66 194
rect 64 193 65 194
rect 63 193 64 194
rect 62 193 63 194
rect 61 193 62 194
rect 60 193 61 194
rect 59 193 60 194
rect 58 193 59 194
rect 57 193 58 194
rect 56 193 57 194
rect 55 193 56 194
rect 54 193 55 194
rect 53 193 54 194
rect 52 193 53 194
rect 51 193 52 194
rect 50 193 51 194
rect 49 193 50 194
rect 48 193 49 194
rect 47 193 48 194
rect 46 193 47 194
rect 45 193 46 194
rect 44 193 45 194
rect 43 193 44 194
rect 42 193 43 194
rect 41 193 42 194
rect 40 193 41 194
rect 39 193 40 194
rect 38 193 39 194
rect 37 193 38 194
rect 36 193 37 194
rect 35 193 36 194
rect 34 193 35 194
rect 33 193 34 194
rect 32 193 33 194
rect 31 193 32 194
rect 30 193 31 194
rect 29 193 30 194
rect 28 193 29 194
rect 27 193 28 194
rect 26 193 27 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 17 193 18 194
rect 16 193 17 194
rect 72 194 73 195
rect 71 194 72 195
rect 70 194 71 195
rect 69 194 70 195
rect 68 194 69 195
rect 67 194 68 195
rect 66 194 67 195
rect 65 194 66 195
rect 64 194 65 195
rect 63 194 64 195
rect 62 194 63 195
rect 61 194 62 195
rect 60 194 61 195
rect 59 194 60 195
rect 58 194 59 195
rect 57 194 58 195
rect 56 194 57 195
rect 55 194 56 195
rect 54 194 55 195
rect 53 194 54 195
rect 52 194 53 195
rect 51 194 52 195
rect 50 194 51 195
rect 49 194 50 195
rect 48 194 49 195
rect 47 194 48 195
rect 46 194 47 195
rect 45 194 46 195
rect 44 194 45 195
rect 43 194 44 195
rect 42 194 43 195
rect 41 194 42 195
rect 40 194 41 195
rect 39 194 40 195
rect 38 194 39 195
rect 37 194 38 195
rect 36 194 37 195
rect 35 194 36 195
rect 34 194 35 195
rect 33 194 34 195
rect 32 194 33 195
rect 31 194 32 195
rect 30 194 31 195
rect 29 194 30 195
rect 28 194 29 195
rect 27 194 28 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 17 194 18 195
rect 16 194 17 195
rect 71 195 72 196
rect 70 195 71 196
rect 69 195 70 196
rect 68 195 69 196
rect 67 195 68 196
rect 66 195 67 196
rect 65 195 66 196
rect 64 195 65 196
rect 63 195 64 196
rect 62 195 63 196
rect 61 195 62 196
rect 60 195 61 196
rect 59 195 60 196
rect 58 195 59 196
rect 57 195 58 196
rect 56 195 57 196
rect 55 195 56 196
rect 54 195 55 196
rect 53 195 54 196
rect 52 195 53 196
rect 51 195 52 196
rect 50 195 51 196
rect 49 195 50 196
rect 48 195 49 196
rect 47 195 48 196
rect 46 195 47 196
rect 45 195 46 196
rect 44 195 45 196
rect 43 195 44 196
rect 42 195 43 196
rect 41 195 42 196
rect 40 195 41 196
rect 39 195 40 196
rect 38 195 39 196
rect 37 195 38 196
rect 36 195 37 196
rect 35 195 36 196
rect 34 195 35 196
rect 33 195 34 196
rect 32 195 33 196
rect 31 195 32 196
rect 30 195 31 196
rect 29 195 30 196
rect 28 195 29 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 17 195 18 196
rect 16 195 17 196
rect 69 196 70 197
rect 68 196 69 197
rect 67 196 68 197
rect 66 196 67 197
rect 65 196 66 197
rect 64 196 65 197
rect 63 196 64 197
rect 62 196 63 197
rect 61 196 62 197
rect 60 196 61 197
rect 59 196 60 197
rect 58 196 59 197
rect 57 196 58 197
rect 56 196 57 197
rect 55 196 56 197
rect 54 196 55 197
rect 53 196 54 197
rect 52 196 53 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 48 196 49 197
rect 47 196 48 197
rect 46 196 47 197
rect 45 196 46 197
rect 44 196 45 197
rect 43 196 44 197
rect 42 196 43 197
rect 41 196 42 197
rect 40 196 41 197
rect 39 196 40 197
rect 38 196 39 197
rect 37 196 38 197
rect 36 196 37 197
rect 35 196 36 197
rect 34 196 35 197
rect 33 196 34 197
rect 32 196 33 197
rect 31 196 32 197
rect 30 196 31 197
rect 29 196 30 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 17 196 18 197
rect 16 196 17 197
rect 66 197 67 198
rect 65 197 66 198
rect 64 197 65 198
rect 63 197 64 198
rect 62 197 63 198
rect 61 197 62 198
rect 60 197 61 198
rect 59 197 60 198
rect 58 197 59 198
rect 57 197 58 198
rect 56 197 57 198
rect 55 197 56 198
rect 54 197 55 198
rect 53 197 54 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 48 197 49 198
rect 47 197 48 198
rect 46 197 47 198
rect 45 197 46 198
rect 44 197 45 198
rect 43 197 44 198
rect 42 197 43 198
rect 41 197 42 198
rect 40 197 41 198
rect 39 197 40 198
rect 38 197 39 198
rect 37 197 38 198
rect 36 197 37 198
rect 35 197 36 198
rect 34 197 35 198
rect 33 197 34 198
rect 32 197 33 198
rect 31 197 32 198
rect 30 197 31 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 17 197 18 198
rect 16 197 17 198
rect 142 198 143 199
rect 141 198 142 199
rect 63 198 64 199
rect 62 198 63 199
rect 61 198 62 199
rect 60 198 61 199
rect 59 198 60 199
rect 58 198 59 199
rect 57 198 58 199
rect 56 198 57 199
rect 55 198 56 199
rect 54 198 55 199
rect 53 198 54 199
rect 52 198 53 199
rect 51 198 52 199
rect 50 198 51 199
rect 49 198 50 199
rect 48 198 49 199
rect 47 198 48 199
rect 46 198 47 199
rect 45 198 46 199
rect 44 198 45 199
rect 43 198 44 199
rect 42 198 43 199
rect 41 198 42 199
rect 40 198 41 199
rect 39 198 40 199
rect 38 198 39 199
rect 37 198 38 199
rect 36 198 37 199
rect 35 198 36 199
rect 34 198 35 199
rect 33 198 34 199
rect 32 198 33 199
rect 31 198 32 199
rect 30 198 31 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 24 198 25 199
rect 23 198 24 199
rect 22 198 23 199
rect 21 198 22 199
rect 20 198 21 199
rect 19 198 20 199
rect 18 198 19 199
rect 17 198 18 199
rect 16 198 17 199
rect 143 199 144 200
rect 142 199 143 200
rect 141 199 142 200
rect 140 199 141 200
rect 55 199 56 200
rect 54 199 55 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 50 199 51 200
rect 49 199 50 200
rect 48 199 49 200
rect 47 199 48 200
rect 46 199 47 200
rect 45 199 46 200
rect 44 199 45 200
rect 43 199 44 200
rect 42 199 43 200
rect 41 199 42 200
rect 40 199 41 200
rect 39 199 40 200
rect 38 199 39 200
rect 37 199 38 200
rect 36 199 37 200
rect 35 199 36 200
rect 34 199 35 200
rect 33 199 34 200
rect 32 199 33 200
rect 31 199 32 200
rect 30 199 31 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 22 199 23 200
rect 21 199 22 200
rect 20 199 21 200
rect 19 199 20 200
rect 18 199 19 200
rect 17 199 18 200
rect 16 199 17 200
rect 144 200 145 201
rect 143 200 144 201
rect 142 200 143 201
rect 141 200 142 201
rect 140 200 141 201
rect 139 200 140 201
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 141 201 142 202
rect 140 201 141 202
rect 139 201 140 202
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 140 202 141 203
rect 139 202 140 203
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 140 203 141 204
rect 142 204 143 205
rect 141 204 142 205
rect 140 220 141 221
rect 139 220 140 221
rect 138 220 139 221
rect 137 220 138 221
rect 136 220 137 221
rect 135 220 136 221
rect 134 220 135 221
rect 133 220 134 221
rect 132 220 133 221
rect 131 220 132 221
rect 130 220 131 221
rect 143 221 144 222
rect 142 221 143 222
rect 141 221 142 222
rect 140 221 141 222
rect 139 221 140 222
rect 138 221 139 222
rect 137 221 138 222
rect 136 221 137 222
rect 135 221 136 222
rect 134 221 135 222
rect 133 221 134 222
rect 132 221 133 222
rect 131 221 132 222
rect 130 221 131 222
rect 129 221 130 222
rect 128 221 129 222
rect 127 221 128 222
rect 126 221 127 222
rect 145 222 146 223
rect 144 222 145 223
rect 143 222 144 223
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 137 222 138 223
rect 136 222 137 223
rect 135 222 136 223
rect 134 222 135 223
rect 133 222 134 223
rect 132 222 133 223
rect 131 222 132 223
rect 130 222 131 223
rect 129 222 130 223
rect 128 222 129 223
rect 127 222 128 223
rect 126 222 127 223
rect 125 222 126 223
rect 124 222 125 223
rect 147 223 148 224
rect 146 223 147 224
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 138 223 139 224
rect 137 223 138 224
rect 136 223 137 224
rect 135 223 136 224
rect 134 223 135 224
rect 133 223 134 224
rect 132 223 133 224
rect 131 223 132 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 127 223 128 224
rect 126 223 127 224
rect 125 223 126 224
rect 124 223 125 224
rect 123 223 124 224
rect 122 223 123 224
rect 149 224 150 225
rect 148 224 149 225
rect 147 224 148 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 139 224 140 225
rect 138 224 139 225
rect 137 224 138 225
rect 136 224 137 225
rect 135 224 136 225
rect 134 224 135 225
rect 133 224 134 225
rect 132 224 133 225
rect 131 224 132 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 125 224 126 225
rect 124 224 125 225
rect 123 224 124 225
rect 122 224 123 225
rect 121 224 122 225
rect 150 225 151 226
rect 149 225 150 226
rect 148 225 149 226
rect 147 225 148 226
rect 146 225 147 226
rect 145 225 146 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 141 225 142 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 123 225 124 226
rect 122 225 123 226
rect 121 225 122 226
rect 120 225 121 226
rect 119 225 120 226
rect 150 226 151 227
rect 149 226 150 227
rect 148 226 149 227
rect 147 226 148 227
rect 146 226 147 227
rect 145 226 146 227
rect 144 226 145 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 122 226 123 227
rect 121 226 122 227
rect 120 226 121 227
rect 119 226 120 227
rect 150 227 151 228
rect 149 227 150 228
rect 148 227 149 228
rect 147 227 148 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 120 227 121 228
rect 119 227 120 228
rect 150 228 151 229
rect 149 228 150 229
rect 148 228 149 229
rect 121 228 122 229
rect 120 228 121 229
rect 119 228 120 229
rect 150 229 151 230
rect 119 229 120 230
rect 138 232 139 233
rect 137 232 138 233
rect 136 232 137 233
rect 135 232 136 233
rect 134 232 135 233
rect 133 232 134 233
rect 140 233 141 234
rect 139 233 140 234
rect 138 233 139 234
rect 137 233 138 234
rect 136 233 137 234
rect 135 233 136 234
rect 134 233 135 234
rect 133 233 134 234
rect 132 233 133 234
rect 131 233 132 234
rect 130 233 131 234
rect 141 234 142 235
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 137 234 138 235
rect 136 234 137 235
rect 135 234 136 235
rect 134 234 135 235
rect 133 234 134 235
rect 132 234 133 235
rect 131 234 132 235
rect 130 234 131 235
rect 129 234 130 235
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 137 235 138 236
rect 136 235 137 236
rect 135 235 136 236
rect 134 235 135 236
rect 133 235 134 236
rect 132 235 133 236
rect 131 235 132 236
rect 130 235 131 236
rect 129 235 130 236
rect 128 235 129 236
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 137 236 138 237
rect 136 236 137 237
rect 135 236 136 237
rect 134 236 135 237
rect 133 236 134 237
rect 132 236 133 237
rect 131 236 132 237
rect 130 236 131 237
rect 129 236 130 237
rect 128 236 129 237
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 137 237 138 238
rect 136 237 137 238
rect 135 237 136 238
rect 134 237 135 238
rect 133 237 134 238
rect 132 237 133 238
rect 131 237 132 238
rect 130 237 131 238
rect 129 237 130 238
rect 128 237 129 238
rect 127 237 128 238
rect 61 237 62 238
rect 60 237 61 238
rect 59 237 60 238
rect 58 237 59 238
rect 57 237 58 238
rect 56 237 57 238
rect 55 237 56 238
rect 54 237 55 238
rect 53 237 54 238
rect 52 237 53 238
rect 51 237 52 238
rect 50 237 51 238
rect 49 237 50 238
rect 48 237 49 238
rect 47 237 48 238
rect 46 237 47 238
rect 45 237 46 238
rect 44 237 45 238
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 132 238 133 239
rect 131 238 132 239
rect 130 238 131 239
rect 129 238 130 239
rect 128 238 129 239
rect 127 238 128 239
rect 65 238 66 239
rect 64 238 65 239
rect 63 238 64 239
rect 62 238 63 239
rect 61 238 62 239
rect 60 238 61 239
rect 59 238 60 239
rect 58 238 59 239
rect 57 238 58 239
rect 56 238 57 239
rect 55 238 56 239
rect 54 238 55 239
rect 53 238 54 239
rect 52 238 53 239
rect 51 238 52 239
rect 50 238 51 239
rect 49 238 50 239
rect 48 238 49 239
rect 47 238 48 239
rect 46 238 47 239
rect 45 238 46 239
rect 44 238 45 239
rect 43 238 44 239
rect 42 238 43 239
rect 41 238 42 239
rect 40 238 41 239
rect 39 238 40 239
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 130 239 131 240
rect 129 239 130 240
rect 128 239 129 240
rect 127 239 128 240
rect 126 239 127 240
rect 68 239 69 240
rect 67 239 68 240
rect 66 239 67 240
rect 65 239 66 240
rect 64 239 65 240
rect 63 239 64 240
rect 62 239 63 240
rect 61 239 62 240
rect 60 239 61 240
rect 59 239 60 240
rect 58 239 59 240
rect 57 239 58 240
rect 56 239 57 240
rect 55 239 56 240
rect 54 239 55 240
rect 53 239 54 240
rect 52 239 53 240
rect 51 239 52 240
rect 50 239 51 240
rect 49 239 50 240
rect 48 239 49 240
rect 47 239 48 240
rect 46 239 47 240
rect 45 239 46 240
rect 44 239 45 240
rect 43 239 44 240
rect 42 239 43 240
rect 41 239 42 240
rect 40 239 41 240
rect 39 239 40 240
rect 38 239 39 240
rect 37 239 38 240
rect 36 239 37 240
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 140 240 141 241
rect 130 240 131 241
rect 129 240 130 241
rect 128 240 129 241
rect 127 240 128 241
rect 126 240 127 241
rect 70 240 71 241
rect 69 240 70 241
rect 68 240 69 241
rect 67 240 68 241
rect 66 240 67 241
rect 65 240 66 241
rect 64 240 65 241
rect 63 240 64 241
rect 62 240 63 241
rect 61 240 62 241
rect 60 240 61 241
rect 59 240 60 241
rect 58 240 59 241
rect 57 240 58 241
rect 56 240 57 241
rect 55 240 56 241
rect 54 240 55 241
rect 53 240 54 241
rect 52 240 53 241
rect 51 240 52 241
rect 50 240 51 241
rect 49 240 50 241
rect 48 240 49 241
rect 47 240 48 241
rect 46 240 47 241
rect 45 240 46 241
rect 44 240 45 241
rect 43 240 44 241
rect 42 240 43 241
rect 41 240 42 241
rect 40 240 41 241
rect 39 240 40 241
rect 38 240 39 241
rect 37 240 38 241
rect 36 240 37 241
rect 35 240 36 241
rect 34 240 35 241
rect 33 240 34 241
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 141 241 142 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 127 241 128 242
rect 126 241 127 242
rect 72 241 73 242
rect 71 241 72 242
rect 70 241 71 242
rect 69 241 70 242
rect 68 241 69 242
rect 67 241 68 242
rect 66 241 67 242
rect 65 241 66 242
rect 64 241 65 242
rect 63 241 64 242
rect 62 241 63 242
rect 61 241 62 242
rect 60 241 61 242
rect 59 241 60 242
rect 58 241 59 242
rect 57 241 58 242
rect 56 241 57 242
rect 55 241 56 242
rect 54 241 55 242
rect 53 241 54 242
rect 52 241 53 242
rect 51 241 52 242
rect 50 241 51 242
rect 49 241 50 242
rect 48 241 49 242
rect 47 241 48 242
rect 46 241 47 242
rect 45 241 46 242
rect 44 241 45 242
rect 43 241 44 242
rect 42 241 43 242
rect 41 241 42 242
rect 40 241 41 242
rect 39 241 40 242
rect 38 241 39 242
rect 37 241 38 242
rect 36 241 37 242
rect 35 241 36 242
rect 34 241 35 242
rect 33 241 34 242
rect 32 241 33 242
rect 31 241 32 242
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 141 242 142 243
rect 129 242 130 243
rect 128 242 129 243
rect 127 242 128 243
rect 126 242 127 243
rect 74 242 75 243
rect 73 242 74 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 56 242 57 243
rect 55 242 56 243
rect 54 242 55 243
rect 53 242 54 243
rect 52 242 53 243
rect 51 242 52 243
rect 50 242 51 243
rect 49 242 50 243
rect 48 242 49 243
rect 47 242 48 243
rect 46 242 47 243
rect 45 242 46 243
rect 44 242 45 243
rect 43 242 44 243
rect 42 242 43 243
rect 41 242 42 243
rect 40 242 41 243
rect 39 242 40 243
rect 38 242 39 243
rect 37 242 38 243
rect 36 242 37 243
rect 35 242 36 243
rect 34 242 35 243
rect 33 242 34 243
rect 32 242 33 243
rect 31 242 32 243
rect 30 242 31 243
rect 144 243 145 244
rect 143 243 144 244
rect 142 243 143 244
rect 141 243 142 244
rect 129 243 130 244
rect 128 243 129 244
rect 127 243 128 244
rect 126 243 127 244
rect 75 243 76 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 56 243 57 244
rect 55 243 56 244
rect 54 243 55 244
rect 53 243 54 244
rect 52 243 53 244
rect 51 243 52 244
rect 50 243 51 244
rect 49 243 50 244
rect 48 243 49 244
rect 47 243 48 244
rect 46 243 47 244
rect 45 243 46 244
rect 44 243 45 244
rect 43 243 44 244
rect 42 243 43 244
rect 41 243 42 244
rect 40 243 41 244
rect 39 243 40 244
rect 38 243 39 244
rect 37 243 38 244
rect 36 243 37 244
rect 35 243 36 244
rect 34 243 35 244
rect 33 243 34 244
rect 32 243 33 244
rect 31 243 32 244
rect 30 243 31 244
rect 29 243 30 244
rect 28 243 29 244
rect 144 244 145 245
rect 143 244 144 245
rect 142 244 143 245
rect 141 244 142 245
rect 140 244 141 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 127 244 128 245
rect 126 244 127 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 56 244 57 245
rect 55 244 56 245
rect 54 244 55 245
rect 53 244 54 245
rect 52 244 53 245
rect 51 244 52 245
rect 50 244 51 245
rect 49 244 50 245
rect 48 244 49 245
rect 47 244 48 245
rect 46 244 47 245
rect 45 244 46 245
rect 44 244 45 245
rect 43 244 44 245
rect 42 244 43 245
rect 41 244 42 245
rect 40 244 41 245
rect 39 244 40 245
rect 38 244 39 245
rect 37 244 38 245
rect 36 244 37 245
rect 35 244 36 245
rect 34 244 35 245
rect 33 244 34 245
rect 32 244 33 245
rect 31 244 32 245
rect 30 244 31 245
rect 29 244 30 245
rect 28 244 29 245
rect 27 244 28 245
rect 144 245 145 246
rect 143 245 144 246
rect 142 245 143 246
rect 141 245 142 246
rect 140 245 141 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 127 245 128 246
rect 126 245 127 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 56 245 57 246
rect 55 245 56 246
rect 54 245 55 246
rect 53 245 54 246
rect 52 245 53 246
rect 51 245 52 246
rect 50 245 51 246
rect 49 245 50 246
rect 48 245 49 246
rect 47 245 48 246
rect 46 245 47 246
rect 45 245 46 246
rect 44 245 45 246
rect 43 245 44 246
rect 42 245 43 246
rect 41 245 42 246
rect 40 245 41 246
rect 39 245 40 246
rect 38 245 39 246
rect 37 245 38 246
rect 36 245 37 246
rect 35 245 36 246
rect 34 245 35 246
rect 33 245 34 246
rect 32 245 33 246
rect 31 245 32 246
rect 30 245 31 246
rect 29 245 30 246
rect 28 245 29 246
rect 27 245 28 246
rect 26 245 27 246
rect 25 245 26 246
rect 143 246 144 247
rect 142 246 143 247
rect 141 246 142 247
rect 140 246 141 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 127 246 128 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 56 246 57 247
rect 55 246 56 247
rect 54 246 55 247
rect 53 246 54 247
rect 52 246 53 247
rect 51 246 52 247
rect 50 246 51 247
rect 49 246 50 247
rect 48 246 49 247
rect 47 246 48 247
rect 46 246 47 247
rect 45 246 46 247
rect 44 246 45 247
rect 43 246 44 247
rect 42 246 43 247
rect 41 246 42 247
rect 40 246 41 247
rect 39 246 40 247
rect 38 246 39 247
rect 37 246 38 247
rect 36 246 37 247
rect 35 246 36 247
rect 34 246 35 247
rect 33 246 34 247
rect 32 246 33 247
rect 31 246 32 247
rect 30 246 31 247
rect 29 246 30 247
rect 28 246 29 247
rect 27 246 28 247
rect 26 246 27 247
rect 25 246 26 247
rect 24 246 25 247
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 58 247 59 248
rect 57 247 58 248
rect 56 247 57 248
rect 55 247 56 248
rect 54 247 55 248
rect 53 247 54 248
rect 52 247 53 248
rect 51 247 52 248
rect 50 247 51 248
rect 49 247 50 248
rect 48 247 49 248
rect 47 247 48 248
rect 46 247 47 248
rect 45 247 46 248
rect 44 247 45 248
rect 43 247 44 248
rect 42 247 43 248
rect 41 247 42 248
rect 40 247 41 248
rect 39 247 40 248
rect 38 247 39 248
rect 37 247 38 248
rect 36 247 37 248
rect 35 247 36 248
rect 34 247 35 248
rect 33 247 34 248
rect 32 247 33 248
rect 31 247 32 248
rect 30 247 31 248
rect 29 247 30 248
rect 28 247 29 248
rect 27 247 28 248
rect 26 247 27 248
rect 25 247 26 248
rect 24 247 25 248
rect 23 247 24 248
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 57 248 58 249
rect 56 248 57 249
rect 55 248 56 249
rect 54 248 55 249
rect 53 248 54 249
rect 52 248 53 249
rect 51 248 52 249
rect 50 248 51 249
rect 49 248 50 249
rect 48 248 49 249
rect 47 248 48 249
rect 46 248 47 249
rect 45 248 46 249
rect 44 248 45 249
rect 43 248 44 249
rect 42 248 43 249
rect 41 248 42 249
rect 40 248 41 249
rect 39 248 40 249
rect 38 248 39 249
rect 37 248 38 249
rect 36 248 37 249
rect 35 248 36 249
rect 34 248 35 249
rect 33 248 34 249
rect 32 248 33 249
rect 31 248 32 249
rect 30 248 31 249
rect 29 248 30 249
rect 28 248 29 249
rect 27 248 28 249
rect 26 248 27 249
rect 25 248 26 249
rect 24 248 25 249
rect 23 248 24 249
rect 22 248 23 249
rect 150 249 151 250
rect 119 249 120 250
rect 80 249 81 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 56 249 57 250
rect 55 249 56 250
rect 54 249 55 250
rect 53 249 54 250
rect 52 249 53 250
rect 51 249 52 250
rect 50 249 51 250
rect 49 249 50 250
rect 48 249 49 250
rect 47 249 48 250
rect 46 249 47 250
rect 45 249 46 250
rect 44 249 45 250
rect 43 249 44 250
rect 42 249 43 250
rect 41 249 42 250
rect 40 249 41 250
rect 39 249 40 250
rect 38 249 39 250
rect 37 249 38 250
rect 36 249 37 250
rect 35 249 36 250
rect 34 249 35 250
rect 33 249 34 250
rect 32 249 33 250
rect 31 249 32 250
rect 30 249 31 250
rect 29 249 30 250
rect 28 249 29 250
rect 27 249 28 250
rect 26 249 27 250
rect 25 249 26 250
rect 24 249 25 250
rect 23 249 24 250
rect 22 249 23 250
rect 21 249 22 250
rect 150 250 151 251
rect 149 250 150 251
rect 120 250 121 251
rect 119 250 120 251
rect 80 250 81 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 56 250 57 251
rect 55 250 56 251
rect 54 250 55 251
rect 53 250 54 251
rect 52 250 53 251
rect 51 250 52 251
rect 50 250 51 251
rect 49 250 50 251
rect 48 250 49 251
rect 47 250 48 251
rect 46 250 47 251
rect 45 250 46 251
rect 44 250 45 251
rect 43 250 44 251
rect 42 250 43 251
rect 41 250 42 251
rect 40 250 41 251
rect 39 250 40 251
rect 38 250 39 251
rect 37 250 38 251
rect 36 250 37 251
rect 35 250 36 251
rect 34 250 35 251
rect 33 250 34 251
rect 32 250 33 251
rect 31 250 32 251
rect 30 250 31 251
rect 29 250 30 251
rect 28 250 29 251
rect 27 250 28 251
rect 26 250 27 251
rect 25 250 26 251
rect 24 250 25 251
rect 23 250 24 251
rect 22 250 23 251
rect 21 250 22 251
rect 150 251 151 252
rect 149 251 150 252
rect 148 251 149 252
rect 147 251 148 252
rect 122 251 123 252
rect 121 251 122 252
rect 120 251 121 252
rect 119 251 120 252
rect 81 251 82 252
rect 80 251 81 252
rect 79 251 80 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 71 251 72 252
rect 70 251 71 252
rect 69 251 70 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 56 251 57 252
rect 55 251 56 252
rect 54 251 55 252
rect 53 251 54 252
rect 52 251 53 252
rect 51 251 52 252
rect 50 251 51 252
rect 49 251 50 252
rect 48 251 49 252
rect 47 251 48 252
rect 46 251 47 252
rect 45 251 46 252
rect 44 251 45 252
rect 43 251 44 252
rect 42 251 43 252
rect 41 251 42 252
rect 40 251 41 252
rect 39 251 40 252
rect 38 251 39 252
rect 37 251 38 252
rect 36 251 37 252
rect 35 251 36 252
rect 34 251 35 252
rect 33 251 34 252
rect 32 251 33 252
rect 31 251 32 252
rect 30 251 31 252
rect 29 251 30 252
rect 28 251 29 252
rect 27 251 28 252
rect 26 251 27 252
rect 25 251 26 252
rect 24 251 25 252
rect 23 251 24 252
rect 22 251 23 252
rect 21 251 22 252
rect 20 251 21 252
rect 150 252 151 253
rect 149 252 150 253
rect 148 252 149 253
rect 147 252 148 253
rect 146 252 147 253
rect 145 252 146 253
rect 124 252 125 253
rect 123 252 124 253
rect 122 252 123 253
rect 121 252 122 253
rect 120 252 121 253
rect 119 252 120 253
rect 81 252 82 253
rect 80 252 81 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 72 252 73 253
rect 71 252 72 253
rect 70 252 71 253
rect 69 252 70 253
rect 68 252 69 253
rect 67 252 68 253
rect 66 252 67 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 55 252 56 253
rect 54 252 55 253
rect 53 252 54 253
rect 52 252 53 253
rect 51 252 52 253
rect 50 252 51 253
rect 49 252 50 253
rect 48 252 49 253
rect 47 252 48 253
rect 46 252 47 253
rect 45 252 46 253
rect 44 252 45 253
rect 43 252 44 253
rect 42 252 43 253
rect 41 252 42 253
rect 40 252 41 253
rect 39 252 40 253
rect 38 252 39 253
rect 37 252 38 253
rect 36 252 37 253
rect 35 252 36 253
rect 34 252 35 253
rect 33 252 34 253
rect 32 252 33 253
rect 31 252 32 253
rect 30 252 31 253
rect 29 252 30 253
rect 28 252 29 253
rect 27 252 28 253
rect 26 252 27 253
rect 25 252 26 253
rect 24 252 25 253
rect 23 252 24 253
rect 22 252 23 253
rect 21 252 22 253
rect 20 252 21 253
rect 19 252 20 253
rect 150 253 151 254
rect 149 253 150 254
rect 148 253 149 254
rect 147 253 148 254
rect 146 253 147 254
rect 145 253 146 254
rect 144 253 145 254
rect 143 253 144 254
rect 126 253 127 254
rect 125 253 126 254
rect 124 253 125 254
rect 123 253 124 254
rect 122 253 123 254
rect 121 253 122 254
rect 120 253 121 254
rect 119 253 120 254
rect 82 253 83 254
rect 81 253 82 254
rect 80 253 81 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 72 253 73 254
rect 71 253 72 254
rect 70 253 71 254
rect 69 253 70 254
rect 68 253 69 254
rect 67 253 68 254
rect 66 253 67 254
rect 65 253 66 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 60 253 61 254
rect 59 253 60 254
rect 58 253 59 254
rect 57 253 58 254
rect 56 253 57 254
rect 55 253 56 254
rect 54 253 55 254
rect 53 253 54 254
rect 52 253 53 254
rect 51 253 52 254
rect 50 253 51 254
rect 49 253 50 254
rect 48 253 49 254
rect 47 253 48 254
rect 46 253 47 254
rect 45 253 46 254
rect 44 253 45 254
rect 43 253 44 254
rect 42 253 43 254
rect 41 253 42 254
rect 40 253 41 254
rect 39 253 40 254
rect 38 253 39 254
rect 37 253 38 254
rect 36 253 37 254
rect 35 253 36 254
rect 34 253 35 254
rect 33 253 34 254
rect 32 253 33 254
rect 31 253 32 254
rect 30 253 31 254
rect 29 253 30 254
rect 28 253 29 254
rect 27 253 28 254
rect 26 253 27 254
rect 25 253 26 254
rect 24 253 25 254
rect 23 253 24 254
rect 22 253 23 254
rect 21 253 22 254
rect 20 253 21 254
rect 19 253 20 254
rect 149 254 150 255
rect 148 254 149 255
rect 147 254 148 255
rect 146 254 147 255
rect 145 254 146 255
rect 144 254 145 255
rect 143 254 144 255
rect 142 254 143 255
rect 141 254 142 255
rect 140 254 141 255
rect 139 254 140 255
rect 138 254 139 255
rect 131 254 132 255
rect 130 254 131 255
rect 129 254 130 255
rect 128 254 129 255
rect 127 254 128 255
rect 126 254 127 255
rect 125 254 126 255
rect 124 254 125 255
rect 123 254 124 255
rect 122 254 123 255
rect 121 254 122 255
rect 120 254 121 255
rect 82 254 83 255
rect 81 254 82 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 71 254 72 255
rect 70 254 71 255
rect 69 254 70 255
rect 68 254 69 255
rect 67 254 68 255
rect 66 254 67 255
rect 65 254 66 255
rect 64 254 65 255
rect 63 254 64 255
rect 62 254 63 255
rect 61 254 62 255
rect 60 254 61 255
rect 59 254 60 255
rect 58 254 59 255
rect 57 254 58 255
rect 56 254 57 255
rect 55 254 56 255
rect 54 254 55 255
rect 53 254 54 255
rect 52 254 53 255
rect 51 254 52 255
rect 50 254 51 255
rect 49 254 50 255
rect 48 254 49 255
rect 47 254 48 255
rect 46 254 47 255
rect 45 254 46 255
rect 44 254 45 255
rect 43 254 44 255
rect 42 254 43 255
rect 41 254 42 255
rect 40 254 41 255
rect 39 254 40 255
rect 38 254 39 255
rect 37 254 38 255
rect 36 254 37 255
rect 35 254 36 255
rect 34 254 35 255
rect 33 254 34 255
rect 32 254 33 255
rect 31 254 32 255
rect 30 254 31 255
rect 29 254 30 255
rect 28 254 29 255
rect 27 254 28 255
rect 26 254 27 255
rect 25 254 26 255
rect 24 254 25 255
rect 23 254 24 255
rect 22 254 23 255
rect 21 254 22 255
rect 20 254 21 255
rect 19 254 20 255
rect 18 254 19 255
rect 148 255 149 256
rect 147 255 148 256
rect 146 255 147 256
rect 145 255 146 256
rect 144 255 145 256
rect 143 255 144 256
rect 142 255 143 256
rect 141 255 142 256
rect 140 255 141 256
rect 139 255 140 256
rect 138 255 139 256
rect 137 255 138 256
rect 136 255 137 256
rect 135 255 136 256
rect 134 255 135 256
rect 133 255 134 256
rect 132 255 133 256
rect 131 255 132 256
rect 130 255 131 256
rect 129 255 130 256
rect 128 255 129 256
rect 127 255 128 256
rect 126 255 127 256
rect 125 255 126 256
rect 124 255 125 256
rect 123 255 124 256
rect 122 255 123 256
rect 121 255 122 256
rect 82 255 83 256
rect 81 255 82 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 69 255 70 256
rect 68 255 69 256
rect 67 255 68 256
rect 66 255 67 256
rect 65 255 66 256
rect 64 255 65 256
rect 63 255 64 256
rect 62 255 63 256
rect 61 255 62 256
rect 60 255 61 256
rect 59 255 60 256
rect 58 255 59 256
rect 57 255 58 256
rect 56 255 57 256
rect 55 255 56 256
rect 54 255 55 256
rect 53 255 54 256
rect 52 255 53 256
rect 51 255 52 256
rect 50 255 51 256
rect 49 255 50 256
rect 48 255 49 256
rect 47 255 48 256
rect 46 255 47 256
rect 45 255 46 256
rect 44 255 45 256
rect 43 255 44 256
rect 42 255 43 256
rect 41 255 42 256
rect 40 255 41 256
rect 39 255 40 256
rect 38 255 39 256
rect 37 255 38 256
rect 36 255 37 256
rect 35 255 36 256
rect 34 255 35 256
rect 33 255 34 256
rect 32 255 33 256
rect 31 255 32 256
rect 30 255 31 256
rect 29 255 30 256
rect 28 255 29 256
rect 27 255 28 256
rect 26 255 27 256
rect 25 255 26 256
rect 24 255 25 256
rect 23 255 24 256
rect 22 255 23 256
rect 21 255 22 256
rect 20 255 21 256
rect 19 255 20 256
rect 18 255 19 256
rect 146 256 147 257
rect 145 256 146 257
rect 144 256 145 257
rect 143 256 144 257
rect 142 256 143 257
rect 141 256 142 257
rect 140 256 141 257
rect 139 256 140 257
rect 138 256 139 257
rect 137 256 138 257
rect 136 256 137 257
rect 135 256 136 257
rect 134 256 135 257
rect 133 256 134 257
rect 132 256 133 257
rect 131 256 132 257
rect 130 256 131 257
rect 129 256 130 257
rect 128 256 129 257
rect 127 256 128 257
rect 126 256 127 257
rect 125 256 126 257
rect 124 256 125 257
rect 123 256 124 257
rect 82 256 83 257
rect 81 256 82 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 65 256 66 257
rect 64 256 65 257
rect 63 256 64 257
rect 62 256 63 257
rect 59 256 60 257
rect 58 256 59 257
rect 57 256 58 257
rect 56 256 57 257
rect 55 256 56 257
rect 54 256 55 257
rect 53 256 54 257
rect 52 256 53 257
rect 51 256 52 257
rect 50 256 51 257
rect 49 256 50 257
rect 48 256 49 257
rect 47 256 48 257
rect 46 256 47 257
rect 45 256 46 257
rect 40 256 41 257
rect 39 256 40 257
rect 38 256 39 257
rect 37 256 38 257
rect 36 256 37 257
rect 35 256 36 257
rect 34 256 35 257
rect 33 256 34 257
rect 32 256 33 257
rect 31 256 32 257
rect 30 256 31 257
rect 29 256 30 257
rect 28 256 29 257
rect 27 256 28 257
rect 26 256 27 257
rect 25 256 26 257
rect 24 256 25 257
rect 23 256 24 257
rect 22 256 23 257
rect 21 256 22 257
rect 20 256 21 257
rect 19 256 20 257
rect 18 256 19 257
rect 17 256 18 257
rect 144 257 145 258
rect 143 257 144 258
rect 142 257 143 258
rect 141 257 142 258
rect 140 257 141 258
rect 139 257 140 258
rect 138 257 139 258
rect 137 257 138 258
rect 136 257 137 258
rect 135 257 136 258
rect 134 257 135 258
rect 133 257 134 258
rect 132 257 133 258
rect 131 257 132 258
rect 130 257 131 258
rect 129 257 130 258
rect 128 257 129 258
rect 127 257 128 258
rect 126 257 127 258
rect 125 257 126 258
rect 83 257 84 258
rect 82 257 83 258
rect 81 257 82 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 66 257 67 258
rect 55 257 56 258
rect 54 257 55 258
rect 53 257 54 258
rect 52 257 53 258
rect 51 257 52 258
rect 50 257 51 258
rect 49 257 50 258
rect 48 257 49 258
rect 47 257 48 258
rect 46 257 47 258
rect 45 257 46 258
rect 44 257 45 258
rect 37 257 38 258
rect 36 257 37 258
rect 35 257 36 258
rect 34 257 35 258
rect 33 257 34 258
rect 32 257 33 258
rect 31 257 32 258
rect 30 257 31 258
rect 29 257 30 258
rect 28 257 29 258
rect 27 257 28 258
rect 26 257 27 258
rect 25 257 26 258
rect 24 257 25 258
rect 23 257 24 258
rect 22 257 23 258
rect 21 257 22 258
rect 20 257 21 258
rect 19 257 20 258
rect 18 257 19 258
rect 17 257 18 258
rect 142 258 143 259
rect 141 258 142 259
rect 140 258 141 259
rect 139 258 140 259
rect 138 258 139 259
rect 137 258 138 259
rect 136 258 137 259
rect 135 258 136 259
rect 134 258 135 259
rect 133 258 134 259
rect 132 258 133 259
rect 131 258 132 259
rect 130 258 131 259
rect 129 258 130 259
rect 128 258 129 259
rect 83 258 84 259
rect 82 258 83 259
rect 81 258 82 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 67 258 68 259
rect 54 258 55 259
rect 53 258 54 259
rect 52 258 53 259
rect 51 258 52 259
rect 50 258 51 259
rect 49 258 50 259
rect 48 258 49 259
rect 47 258 48 259
rect 46 258 47 259
rect 45 258 46 259
rect 44 258 45 259
rect 43 258 44 259
rect 36 258 37 259
rect 35 258 36 259
rect 34 258 35 259
rect 33 258 34 259
rect 32 258 33 259
rect 31 258 32 259
rect 30 258 31 259
rect 29 258 30 259
rect 28 258 29 259
rect 27 258 28 259
rect 26 258 27 259
rect 25 258 26 259
rect 24 258 25 259
rect 23 258 24 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 18 258 19 259
rect 17 258 18 259
rect 83 259 84 260
rect 82 259 83 260
rect 81 259 82 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 68 259 69 260
rect 53 259 54 260
rect 52 259 53 260
rect 51 259 52 260
rect 50 259 51 260
rect 49 259 50 260
rect 48 259 49 260
rect 47 259 48 260
rect 46 259 47 260
rect 45 259 46 260
rect 44 259 45 260
rect 43 259 44 260
rect 42 259 43 260
rect 34 259 35 260
rect 33 259 34 260
rect 32 259 33 260
rect 31 259 32 260
rect 30 259 31 260
rect 29 259 30 260
rect 28 259 29 260
rect 27 259 28 260
rect 26 259 27 260
rect 25 259 26 260
rect 24 259 25 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 18 259 19 260
rect 17 259 18 260
rect 16 259 17 260
rect 83 260 84 261
rect 82 260 83 261
rect 81 260 82 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 69 260 70 261
rect 52 260 53 261
rect 51 260 52 261
rect 50 260 51 261
rect 49 260 50 261
rect 48 260 49 261
rect 47 260 48 261
rect 46 260 47 261
rect 45 260 46 261
rect 44 260 45 261
rect 43 260 44 261
rect 42 260 43 261
rect 41 260 42 261
rect 33 260 34 261
rect 32 260 33 261
rect 31 260 32 261
rect 30 260 31 261
rect 29 260 30 261
rect 28 260 29 261
rect 27 260 28 261
rect 26 260 27 261
rect 25 260 26 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 18 260 19 261
rect 17 260 18 261
rect 16 260 17 261
rect 83 261 84 262
rect 82 261 83 262
rect 81 261 82 262
rect 80 261 81 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 70 261 71 262
rect 69 261 70 262
rect 52 261 53 262
rect 51 261 52 262
rect 50 261 51 262
rect 49 261 50 262
rect 48 261 49 262
rect 47 261 48 262
rect 46 261 47 262
rect 45 261 46 262
rect 44 261 45 262
rect 43 261 44 262
rect 42 261 43 262
rect 41 261 42 262
rect 32 261 33 262
rect 31 261 32 262
rect 30 261 31 262
rect 29 261 30 262
rect 28 261 29 262
rect 27 261 28 262
rect 26 261 27 262
rect 25 261 26 262
rect 24 261 25 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 17 261 18 262
rect 16 261 17 262
rect 83 262 84 263
rect 82 262 83 263
rect 81 262 82 263
rect 80 262 81 263
rect 79 262 80 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 71 262 72 263
rect 70 262 71 263
rect 69 262 70 263
rect 52 262 53 263
rect 51 262 52 263
rect 50 262 51 263
rect 49 262 50 263
rect 48 262 49 263
rect 47 262 48 263
rect 46 262 47 263
rect 45 262 46 263
rect 44 262 45 263
rect 43 262 44 263
rect 42 262 43 263
rect 41 262 42 263
rect 40 262 41 263
rect 31 262 32 263
rect 30 262 31 263
rect 29 262 30 263
rect 28 262 29 263
rect 27 262 28 263
rect 26 262 27 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 17 262 18 263
rect 16 262 17 263
rect 83 263 84 264
rect 82 263 83 264
rect 81 263 82 264
rect 80 263 81 264
rect 79 263 80 264
rect 78 263 79 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 72 263 73 264
rect 71 263 72 264
rect 70 263 71 264
rect 69 263 70 264
rect 52 263 53 264
rect 51 263 52 264
rect 50 263 51 264
rect 49 263 50 264
rect 48 263 49 264
rect 47 263 48 264
rect 46 263 47 264
rect 45 263 46 264
rect 44 263 45 264
rect 43 263 44 264
rect 42 263 43 264
rect 41 263 42 264
rect 40 263 41 264
rect 31 263 32 264
rect 30 263 31 264
rect 29 263 30 264
rect 28 263 29 264
rect 27 263 28 264
rect 26 263 27 264
rect 25 263 26 264
rect 24 263 25 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 17 263 18 264
rect 16 263 17 264
rect 136 264 137 265
rect 135 264 136 265
rect 134 264 135 265
rect 133 264 134 265
rect 132 264 133 265
rect 131 264 132 265
rect 130 264 131 265
rect 129 264 130 265
rect 128 264 129 265
rect 83 264 84 265
rect 82 264 83 265
rect 81 264 82 265
rect 80 264 81 265
rect 79 264 80 265
rect 78 264 79 265
rect 77 264 78 265
rect 76 264 77 265
rect 75 264 76 265
rect 74 264 75 265
rect 73 264 74 265
rect 72 264 73 265
rect 71 264 72 265
rect 70 264 71 265
rect 69 264 70 265
rect 52 264 53 265
rect 51 264 52 265
rect 50 264 51 265
rect 49 264 50 265
rect 48 264 49 265
rect 47 264 48 265
rect 46 264 47 265
rect 45 264 46 265
rect 44 264 45 265
rect 43 264 44 265
rect 42 264 43 265
rect 41 264 42 265
rect 40 264 41 265
rect 30 264 31 265
rect 29 264 30 265
rect 28 264 29 265
rect 27 264 28 265
rect 26 264 27 265
rect 25 264 26 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 17 264 18 265
rect 16 264 17 265
rect 15 264 16 265
rect 138 265 139 266
rect 137 265 138 266
rect 136 265 137 266
rect 135 265 136 266
rect 134 265 135 266
rect 133 265 134 266
rect 132 265 133 266
rect 131 265 132 266
rect 130 265 131 266
rect 129 265 130 266
rect 128 265 129 266
rect 127 265 128 266
rect 126 265 127 266
rect 83 265 84 266
rect 82 265 83 266
rect 81 265 82 266
rect 80 265 81 266
rect 79 265 80 266
rect 78 265 79 266
rect 77 265 78 266
rect 76 265 77 266
rect 75 265 76 266
rect 74 265 75 266
rect 73 265 74 266
rect 72 265 73 266
rect 71 265 72 266
rect 70 265 71 266
rect 69 265 70 266
rect 68 265 69 266
rect 53 265 54 266
rect 52 265 53 266
rect 51 265 52 266
rect 50 265 51 266
rect 49 265 50 266
rect 48 265 49 266
rect 47 265 48 266
rect 46 265 47 266
rect 45 265 46 266
rect 44 265 45 266
rect 43 265 44 266
rect 42 265 43 266
rect 41 265 42 266
rect 40 265 41 266
rect 39 265 40 266
rect 30 265 31 266
rect 29 265 30 266
rect 28 265 29 266
rect 27 265 28 266
rect 26 265 27 266
rect 25 265 26 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 18 265 19 266
rect 17 265 18 266
rect 16 265 17 266
rect 15 265 16 266
rect 140 266 141 267
rect 139 266 140 267
rect 138 266 139 267
rect 137 266 138 267
rect 136 266 137 267
rect 135 266 136 267
rect 134 266 135 267
rect 133 266 134 267
rect 132 266 133 267
rect 131 266 132 267
rect 130 266 131 267
rect 129 266 130 267
rect 128 266 129 267
rect 127 266 128 267
rect 126 266 127 267
rect 125 266 126 267
rect 124 266 125 267
rect 83 266 84 267
rect 82 266 83 267
rect 81 266 82 267
rect 80 266 81 267
rect 79 266 80 267
rect 78 266 79 267
rect 77 266 78 267
rect 76 266 77 267
rect 75 266 76 267
rect 74 266 75 267
rect 73 266 74 267
rect 72 266 73 267
rect 71 266 72 267
rect 70 266 71 267
rect 69 266 70 267
rect 68 266 69 267
rect 67 266 68 267
rect 54 266 55 267
rect 53 266 54 267
rect 52 266 53 267
rect 51 266 52 267
rect 50 266 51 267
rect 49 266 50 267
rect 48 266 49 267
rect 47 266 48 267
rect 46 266 47 267
rect 45 266 46 267
rect 44 266 45 267
rect 43 266 44 267
rect 42 266 43 267
rect 41 266 42 267
rect 40 266 41 267
rect 39 266 40 267
rect 30 266 31 267
rect 29 266 30 267
rect 28 266 29 267
rect 27 266 28 267
rect 26 266 27 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 16 266 17 267
rect 15 266 16 267
rect 141 267 142 268
rect 140 267 141 268
rect 139 267 140 268
rect 138 267 139 268
rect 137 267 138 268
rect 136 267 137 268
rect 135 267 136 268
rect 134 267 135 268
rect 133 267 134 268
rect 132 267 133 268
rect 131 267 132 268
rect 130 267 131 268
rect 129 267 130 268
rect 128 267 129 268
rect 127 267 128 268
rect 126 267 127 268
rect 125 267 126 268
rect 124 267 125 268
rect 123 267 124 268
rect 82 267 83 268
rect 81 267 82 268
rect 80 267 81 268
rect 79 267 80 268
rect 78 267 79 268
rect 77 267 78 268
rect 76 267 77 268
rect 75 267 76 268
rect 74 267 75 268
rect 73 267 74 268
rect 72 267 73 268
rect 71 267 72 268
rect 70 267 71 268
rect 69 267 70 268
rect 68 267 69 268
rect 67 267 68 268
rect 66 267 67 268
rect 65 267 66 268
rect 56 267 57 268
rect 55 267 56 268
rect 54 267 55 268
rect 53 267 54 268
rect 52 267 53 268
rect 51 267 52 268
rect 50 267 51 268
rect 49 267 50 268
rect 48 267 49 268
rect 47 267 48 268
rect 46 267 47 268
rect 45 267 46 268
rect 44 267 45 268
rect 43 267 44 268
rect 42 267 43 268
rect 41 267 42 268
rect 40 267 41 268
rect 39 267 40 268
rect 29 267 30 268
rect 28 267 29 268
rect 27 267 28 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 16 267 17 268
rect 15 267 16 268
rect 141 268 142 269
rect 140 268 141 269
rect 139 268 140 269
rect 138 268 139 269
rect 137 268 138 269
rect 136 268 137 269
rect 135 268 136 269
rect 134 268 135 269
rect 133 268 134 269
rect 132 268 133 269
rect 131 268 132 269
rect 130 268 131 269
rect 129 268 130 269
rect 128 268 129 269
rect 127 268 128 269
rect 126 268 127 269
rect 125 268 126 269
rect 124 268 125 269
rect 123 268 124 269
rect 122 268 123 269
rect 82 268 83 269
rect 81 268 82 269
rect 80 268 81 269
rect 79 268 80 269
rect 78 268 79 269
rect 77 268 78 269
rect 76 268 77 269
rect 75 268 76 269
rect 74 268 75 269
rect 73 268 74 269
rect 72 268 73 269
rect 71 268 72 269
rect 70 268 71 269
rect 69 268 70 269
rect 68 268 69 269
rect 67 268 68 269
rect 66 268 67 269
rect 65 268 66 269
rect 64 268 65 269
rect 63 268 64 269
rect 62 268 63 269
rect 61 268 62 269
rect 60 268 61 269
rect 59 268 60 269
rect 58 268 59 269
rect 57 268 58 269
rect 56 268 57 269
rect 55 268 56 269
rect 54 268 55 269
rect 53 268 54 269
rect 52 268 53 269
rect 51 268 52 269
rect 50 268 51 269
rect 49 268 50 269
rect 48 268 49 269
rect 47 268 48 269
rect 46 268 47 269
rect 45 268 46 269
rect 44 268 45 269
rect 43 268 44 269
rect 42 268 43 269
rect 41 268 42 269
rect 40 268 41 269
rect 39 268 40 269
rect 29 268 30 269
rect 28 268 29 269
rect 27 268 28 269
rect 26 268 27 269
rect 25 268 26 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 16 268 17 269
rect 15 268 16 269
rect 142 269 143 270
rect 141 269 142 270
rect 140 269 141 270
rect 139 269 140 270
rect 138 269 139 270
rect 137 269 138 270
rect 136 269 137 270
rect 135 269 136 270
rect 134 269 135 270
rect 133 269 134 270
rect 132 269 133 270
rect 131 269 132 270
rect 130 269 131 270
rect 129 269 130 270
rect 128 269 129 270
rect 127 269 128 270
rect 126 269 127 270
rect 125 269 126 270
rect 124 269 125 270
rect 123 269 124 270
rect 122 269 123 270
rect 121 269 122 270
rect 82 269 83 270
rect 81 269 82 270
rect 80 269 81 270
rect 79 269 80 270
rect 78 269 79 270
rect 77 269 78 270
rect 76 269 77 270
rect 75 269 76 270
rect 74 269 75 270
rect 73 269 74 270
rect 72 269 73 270
rect 71 269 72 270
rect 70 269 71 270
rect 69 269 70 270
rect 68 269 69 270
rect 67 269 68 270
rect 66 269 67 270
rect 65 269 66 270
rect 64 269 65 270
rect 63 269 64 270
rect 62 269 63 270
rect 61 269 62 270
rect 60 269 61 270
rect 59 269 60 270
rect 58 269 59 270
rect 57 269 58 270
rect 56 269 57 270
rect 55 269 56 270
rect 54 269 55 270
rect 53 269 54 270
rect 52 269 53 270
rect 51 269 52 270
rect 50 269 51 270
rect 49 269 50 270
rect 48 269 49 270
rect 47 269 48 270
rect 46 269 47 270
rect 45 269 46 270
rect 44 269 45 270
rect 43 269 44 270
rect 42 269 43 270
rect 41 269 42 270
rect 40 269 41 270
rect 39 269 40 270
rect 29 269 30 270
rect 28 269 29 270
rect 27 269 28 270
rect 26 269 27 270
rect 25 269 26 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 16 269 17 270
rect 15 269 16 270
rect 143 270 144 271
rect 142 270 143 271
rect 141 270 142 271
rect 140 270 141 271
rect 139 270 140 271
rect 138 270 139 271
rect 137 270 138 271
rect 136 270 137 271
rect 135 270 136 271
rect 128 270 129 271
rect 127 270 128 271
rect 126 270 127 271
rect 125 270 126 271
rect 124 270 125 271
rect 123 270 124 271
rect 122 270 123 271
rect 121 270 122 271
rect 82 270 83 271
rect 81 270 82 271
rect 80 270 81 271
rect 79 270 80 271
rect 78 270 79 271
rect 77 270 78 271
rect 76 270 77 271
rect 75 270 76 271
rect 74 270 75 271
rect 73 270 74 271
rect 72 270 73 271
rect 71 270 72 271
rect 70 270 71 271
rect 69 270 70 271
rect 68 270 69 271
rect 67 270 68 271
rect 66 270 67 271
rect 65 270 66 271
rect 64 270 65 271
rect 63 270 64 271
rect 62 270 63 271
rect 61 270 62 271
rect 60 270 61 271
rect 59 270 60 271
rect 58 270 59 271
rect 57 270 58 271
rect 56 270 57 271
rect 55 270 56 271
rect 54 270 55 271
rect 53 270 54 271
rect 52 270 53 271
rect 51 270 52 271
rect 50 270 51 271
rect 49 270 50 271
rect 48 270 49 271
rect 47 270 48 271
rect 46 270 47 271
rect 45 270 46 271
rect 44 270 45 271
rect 43 270 44 271
rect 42 270 43 271
rect 41 270 42 271
rect 40 270 41 271
rect 39 270 40 271
rect 29 270 30 271
rect 28 270 29 271
rect 27 270 28 271
rect 26 270 27 271
rect 25 270 26 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 16 270 17 271
rect 15 270 16 271
rect 143 271 144 272
rect 142 271 143 272
rect 141 271 142 272
rect 140 271 141 272
rect 139 271 140 272
rect 138 271 139 272
rect 137 271 138 272
rect 126 271 127 272
rect 125 271 126 272
rect 124 271 125 272
rect 123 271 124 272
rect 122 271 123 272
rect 121 271 122 272
rect 120 271 121 272
rect 81 271 82 272
rect 80 271 81 272
rect 79 271 80 272
rect 78 271 79 272
rect 77 271 78 272
rect 76 271 77 272
rect 75 271 76 272
rect 74 271 75 272
rect 73 271 74 272
rect 72 271 73 272
rect 71 271 72 272
rect 70 271 71 272
rect 69 271 70 272
rect 68 271 69 272
rect 67 271 68 272
rect 66 271 67 272
rect 65 271 66 272
rect 64 271 65 272
rect 63 271 64 272
rect 62 271 63 272
rect 61 271 62 272
rect 60 271 61 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 55 271 56 272
rect 54 271 55 272
rect 53 271 54 272
rect 52 271 53 272
rect 51 271 52 272
rect 50 271 51 272
rect 49 271 50 272
rect 48 271 49 272
rect 47 271 48 272
rect 46 271 47 272
rect 45 271 46 272
rect 44 271 45 272
rect 43 271 44 272
rect 42 271 43 272
rect 41 271 42 272
rect 40 271 41 272
rect 39 271 40 272
rect 29 271 30 272
rect 28 271 29 272
rect 27 271 28 272
rect 26 271 27 272
rect 25 271 26 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 16 271 17 272
rect 15 271 16 272
rect 143 272 144 273
rect 142 272 143 273
rect 141 272 142 273
rect 140 272 141 273
rect 139 272 140 273
rect 138 272 139 273
rect 125 272 126 273
rect 124 272 125 273
rect 123 272 124 273
rect 122 272 123 273
rect 121 272 122 273
rect 120 272 121 273
rect 81 272 82 273
rect 80 272 81 273
rect 79 272 80 273
rect 78 272 79 273
rect 77 272 78 273
rect 76 272 77 273
rect 75 272 76 273
rect 74 272 75 273
rect 73 272 74 273
rect 72 272 73 273
rect 71 272 72 273
rect 70 272 71 273
rect 69 272 70 273
rect 68 272 69 273
rect 67 272 68 273
rect 66 272 67 273
rect 65 272 66 273
rect 64 272 65 273
rect 63 272 64 273
rect 62 272 63 273
rect 61 272 62 273
rect 60 272 61 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 55 272 56 273
rect 54 272 55 273
rect 53 272 54 273
rect 52 272 53 273
rect 51 272 52 273
rect 50 272 51 273
rect 49 272 50 273
rect 48 272 49 273
rect 47 272 48 273
rect 46 272 47 273
rect 45 272 46 273
rect 44 272 45 273
rect 43 272 44 273
rect 42 272 43 273
rect 41 272 42 273
rect 40 272 41 273
rect 39 272 40 273
rect 29 272 30 273
rect 28 272 29 273
rect 27 272 28 273
rect 26 272 27 273
rect 25 272 26 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 16 272 17 273
rect 15 272 16 273
rect 144 273 145 274
rect 143 273 144 274
rect 142 273 143 274
rect 141 273 142 274
rect 140 273 141 274
rect 139 273 140 274
rect 124 273 125 274
rect 123 273 124 274
rect 122 273 123 274
rect 121 273 122 274
rect 120 273 121 274
rect 81 273 82 274
rect 80 273 81 274
rect 79 273 80 274
rect 78 273 79 274
rect 77 273 78 274
rect 76 273 77 274
rect 75 273 76 274
rect 74 273 75 274
rect 73 273 74 274
rect 72 273 73 274
rect 71 273 72 274
rect 70 273 71 274
rect 69 273 70 274
rect 68 273 69 274
rect 67 273 68 274
rect 66 273 67 274
rect 65 273 66 274
rect 64 273 65 274
rect 63 273 64 274
rect 62 273 63 274
rect 61 273 62 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 55 273 56 274
rect 54 273 55 274
rect 53 273 54 274
rect 52 273 53 274
rect 51 273 52 274
rect 50 273 51 274
rect 49 273 50 274
rect 48 273 49 274
rect 47 273 48 274
rect 46 273 47 274
rect 45 273 46 274
rect 44 273 45 274
rect 43 273 44 274
rect 42 273 43 274
rect 41 273 42 274
rect 40 273 41 274
rect 39 273 40 274
rect 29 273 30 274
rect 28 273 29 274
rect 27 273 28 274
rect 26 273 27 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 16 273 17 274
rect 15 273 16 274
rect 144 274 145 275
rect 143 274 144 275
rect 142 274 143 275
rect 141 274 142 275
rect 140 274 141 275
rect 124 274 125 275
rect 123 274 124 275
rect 122 274 123 275
rect 121 274 122 275
rect 120 274 121 275
rect 119 274 120 275
rect 80 274 81 275
rect 79 274 80 275
rect 78 274 79 275
rect 77 274 78 275
rect 76 274 77 275
rect 75 274 76 275
rect 74 274 75 275
rect 73 274 74 275
rect 72 274 73 275
rect 71 274 72 275
rect 70 274 71 275
rect 69 274 70 275
rect 68 274 69 275
rect 67 274 68 275
rect 66 274 67 275
rect 65 274 66 275
rect 64 274 65 275
rect 63 274 64 275
rect 62 274 63 275
rect 61 274 62 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 55 274 56 275
rect 54 274 55 275
rect 53 274 54 275
rect 52 274 53 275
rect 51 274 52 275
rect 50 274 51 275
rect 49 274 50 275
rect 48 274 49 275
rect 47 274 48 275
rect 46 274 47 275
rect 45 274 46 275
rect 44 274 45 275
rect 43 274 44 275
rect 42 274 43 275
rect 41 274 42 275
rect 40 274 41 275
rect 29 274 30 275
rect 28 274 29 275
rect 27 274 28 275
rect 26 274 27 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 16 274 17 275
rect 15 274 16 275
rect 144 275 145 276
rect 143 275 144 276
rect 142 275 143 276
rect 141 275 142 276
rect 140 275 141 276
rect 123 275 124 276
rect 122 275 123 276
rect 121 275 122 276
rect 120 275 121 276
rect 119 275 120 276
rect 80 275 81 276
rect 79 275 80 276
rect 78 275 79 276
rect 77 275 78 276
rect 76 275 77 276
rect 75 275 76 276
rect 74 275 75 276
rect 73 275 74 276
rect 72 275 73 276
rect 71 275 72 276
rect 70 275 71 276
rect 69 275 70 276
rect 68 275 69 276
rect 67 275 68 276
rect 66 275 67 276
rect 65 275 66 276
rect 64 275 65 276
rect 63 275 64 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 56 275 57 276
rect 55 275 56 276
rect 54 275 55 276
rect 53 275 54 276
rect 52 275 53 276
rect 51 275 52 276
rect 50 275 51 276
rect 49 275 50 276
rect 48 275 49 276
rect 47 275 48 276
rect 46 275 47 276
rect 45 275 46 276
rect 44 275 45 276
rect 43 275 44 276
rect 42 275 43 276
rect 41 275 42 276
rect 40 275 41 276
rect 29 275 30 276
rect 28 275 29 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 17 275 18 276
rect 16 275 17 276
rect 15 275 16 276
rect 144 276 145 277
rect 143 276 144 277
rect 142 276 143 277
rect 141 276 142 277
rect 140 276 141 277
rect 134 276 135 277
rect 133 276 134 277
rect 132 276 133 277
rect 131 276 132 277
rect 130 276 131 277
rect 123 276 124 277
rect 122 276 123 277
rect 121 276 122 277
rect 120 276 121 277
rect 119 276 120 277
rect 79 276 80 277
rect 78 276 79 277
rect 77 276 78 277
rect 76 276 77 277
rect 75 276 76 277
rect 74 276 75 277
rect 73 276 74 277
rect 72 276 73 277
rect 71 276 72 277
rect 70 276 71 277
rect 69 276 70 277
rect 68 276 69 277
rect 67 276 68 277
rect 66 276 67 277
rect 65 276 66 277
rect 64 276 65 277
rect 63 276 64 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 56 276 57 277
rect 55 276 56 277
rect 54 276 55 277
rect 53 276 54 277
rect 52 276 53 277
rect 51 276 52 277
rect 50 276 51 277
rect 49 276 50 277
rect 48 276 49 277
rect 47 276 48 277
rect 46 276 47 277
rect 45 276 46 277
rect 44 276 45 277
rect 43 276 44 277
rect 42 276 43 277
rect 41 276 42 277
rect 40 276 41 277
rect 29 276 30 277
rect 28 276 29 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 18 276 19 277
rect 17 276 18 277
rect 16 276 17 277
rect 15 276 16 277
rect 144 277 145 278
rect 143 277 144 278
rect 142 277 143 278
rect 141 277 142 278
rect 140 277 141 278
rect 134 277 135 278
rect 133 277 134 278
rect 132 277 133 278
rect 131 277 132 278
rect 130 277 131 278
rect 123 277 124 278
rect 122 277 123 278
rect 121 277 122 278
rect 120 277 121 278
rect 119 277 120 278
rect 78 277 79 278
rect 77 277 78 278
rect 76 277 77 278
rect 75 277 76 278
rect 74 277 75 278
rect 73 277 74 278
rect 72 277 73 278
rect 71 277 72 278
rect 70 277 71 278
rect 69 277 70 278
rect 68 277 69 278
rect 67 277 68 278
rect 66 277 67 278
rect 65 277 66 278
rect 64 277 65 278
rect 63 277 64 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 56 277 57 278
rect 55 277 56 278
rect 54 277 55 278
rect 53 277 54 278
rect 52 277 53 278
rect 51 277 52 278
rect 50 277 51 278
rect 49 277 50 278
rect 48 277 49 278
rect 47 277 48 278
rect 46 277 47 278
rect 45 277 46 278
rect 44 277 45 278
rect 43 277 44 278
rect 42 277 43 278
rect 41 277 42 278
rect 29 277 30 278
rect 28 277 29 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 19 277 20 278
rect 18 277 19 278
rect 17 277 18 278
rect 16 277 17 278
rect 144 278 145 279
rect 143 278 144 279
rect 142 278 143 279
rect 141 278 142 279
rect 140 278 141 279
rect 134 278 135 279
rect 133 278 134 279
rect 132 278 133 279
rect 131 278 132 279
rect 130 278 131 279
rect 123 278 124 279
rect 122 278 123 279
rect 121 278 122 279
rect 120 278 121 279
rect 119 278 120 279
rect 78 278 79 279
rect 77 278 78 279
rect 76 278 77 279
rect 75 278 76 279
rect 74 278 75 279
rect 73 278 74 279
rect 72 278 73 279
rect 71 278 72 279
rect 70 278 71 279
rect 69 278 70 279
rect 68 278 69 279
rect 67 278 68 279
rect 66 278 67 279
rect 65 278 66 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 57 278 58 279
rect 56 278 57 279
rect 55 278 56 279
rect 54 278 55 279
rect 53 278 54 279
rect 52 278 53 279
rect 51 278 52 279
rect 50 278 51 279
rect 49 278 50 279
rect 48 278 49 279
rect 47 278 48 279
rect 46 278 47 279
rect 45 278 46 279
rect 44 278 45 279
rect 43 278 44 279
rect 42 278 43 279
rect 41 278 42 279
rect 29 278 30 279
rect 28 278 29 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 17 278 18 279
rect 16 278 17 279
rect 144 279 145 280
rect 143 279 144 280
rect 142 279 143 280
rect 141 279 142 280
rect 140 279 141 280
rect 134 279 135 280
rect 133 279 134 280
rect 132 279 133 280
rect 131 279 132 280
rect 130 279 131 280
rect 123 279 124 280
rect 122 279 123 280
rect 121 279 122 280
rect 120 279 121 280
rect 119 279 120 280
rect 77 279 78 280
rect 76 279 77 280
rect 75 279 76 280
rect 74 279 75 280
rect 73 279 74 280
rect 72 279 73 280
rect 71 279 72 280
rect 70 279 71 280
rect 69 279 70 280
rect 68 279 69 280
rect 67 279 68 280
rect 66 279 67 280
rect 65 279 66 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 58 279 59 280
rect 57 279 58 280
rect 56 279 57 280
rect 55 279 56 280
rect 54 279 55 280
rect 53 279 54 280
rect 52 279 53 280
rect 51 279 52 280
rect 50 279 51 280
rect 49 279 50 280
rect 48 279 49 280
rect 47 279 48 280
rect 46 279 47 280
rect 45 279 46 280
rect 44 279 45 280
rect 43 279 44 280
rect 42 279 43 280
rect 30 279 31 280
rect 29 279 30 280
rect 28 279 29 280
rect 27 279 28 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 17 279 18 280
rect 16 279 17 280
rect 144 280 145 281
rect 143 280 144 281
rect 142 280 143 281
rect 141 280 142 281
rect 140 280 141 281
rect 134 280 135 281
rect 133 280 134 281
rect 132 280 133 281
rect 131 280 132 281
rect 130 280 131 281
rect 123 280 124 281
rect 122 280 123 281
rect 121 280 122 281
rect 120 280 121 281
rect 119 280 120 281
rect 76 280 77 281
rect 75 280 76 281
rect 74 280 75 281
rect 73 280 74 281
rect 72 280 73 281
rect 71 280 72 281
rect 70 280 71 281
rect 69 280 70 281
rect 68 280 69 281
rect 67 280 68 281
rect 66 280 67 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 59 280 60 281
rect 58 280 59 281
rect 57 280 58 281
rect 56 280 57 281
rect 55 280 56 281
rect 54 280 55 281
rect 53 280 54 281
rect 52 280 53 281
rect 51 280 52 281
rect 50 280 51 281
rect 49 280 50 281
rect 48 280 49 281
rect 47 280 48 281
rect 46 280 47 281
rect 45 280 46 281
rect 44 280 45 281
rect 43 280 44 281
rect 30 280 31 281
rect 29 280 30 281
rect 28 280 29 281
rect 27 280 28 281
rect 26 280 27 281
rect 25 280 26 281
rect 24 280 25 281
rect 23 280 24 281
rect 22 280 23 281
rect 21 280 22 281
rect 20 280 21 281
rect 19 280 20 281
rect 18 280 19 281
rect 17 280 18 281
rect 16 280 17 281
rect 144 281 145 282
rect 143 281 144 282
rect 142 281 143 282
rect 141 281 142 282
rect 140 281 141 282
rect 139 281 140 282
rect 138 281 139 282
rect 137 281 138 282
rect 136 281 137 282
rect 135 281 136 282
rect 134 281 135 282
rect 133 281 134 282
rect 132 281 133 282
rect 131 281 132 282
rect 130 281 131 282
rect 123 281 124 282
rect 122 281 123 282
rect 121 281 122 282
rect 120 281 121 282
rect 119 281 120 282
rect 75 281 76 282
rect 74 281 75 282
rect 73 281 74 282
rect 72 281 73 282
rect 71 281 72 282
rect 70 281 71 282
rect 69 281 70 282
rect 68 281 69 282
rect 67 281 68 282
rect 66 281 67 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 60 281 61 282
rect 59 281 60 282
rect 58 281 59 282
rect 57 281 58 282
rect 56 281 57 282
rect 55 281 56 282
rect 54 281 55 282
rect 53 281 54 282
rect 52 281 53 282
rect 51 281 52 282
rect 50 281 51 282
rect 49 281 50 282
rect 48 281 49 282
rect 47 281 48 282
rect 46 281 47 282
rect 45 281 46 282
rect 44 281 45 282
rect 30 281 31 282
rect 29 281 30 282
rect 28 281 29 282
rect 27 281 28 282
rect 26 281 27 282
rect 25 281 26 282
rect 24 281 25 282
rect 23 281 24 282
rect 22 281 23 282
rect 21 281 22 282
rect 20 281 21 282
rect 19 281 20 282
rect 18 281 19 282
rect 17 281 18 282
rect 143 282 144 283
rect 142 282 143 283
rect 141 282 142 283
rect 140 282 141 283
rect 139 282 140 283
rect 138 282 139 283
rect 137 282 138 283
rect 136 282 137 283
rect 135 282 136 283
rect 134 282 135 283
rect 133 282 134 283
rect 132 282 133 283
rect 131 282 132 283
rect 130 282 131 283
rect 123 282 124 283
rect 122 282 123 283
rect 121 282 122 283
rect 120 282 121 283
rect 119 282 120 283
rect 73 282 74 283
rect 72 282 73 283
rect 71 282 72 283
rect 70 282 71 283
rect 69 282 70 283
rect 68 282 69 283
rect 67 282 68 283
rect 66 282 67 283
rect 65 282 66 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 61 282 62 283
rect 60 282 61 283
rect 59 282 60 283
rect 58 282 59 283
rect 57 282 58 283
rect 56 282 57 283
rect 55 282 56 283
rect 54 282 55 283
rect 53 282 54 283
rect 52 282 53 283
rect 51 282 52 283
rect 50 282 51 283
rect 49 282 50 283
rect 48 282 49 283
rect 47 282 48 283
rect 46 282 47 283
rect 45 282 46 283
rect 143 283 144 284
rect 142 283 143 284
rect 141 283 142 284
rect 140 283 141 284
rect 139 283 140 284
rect 138 283 139 284
rect 137 283 138 284
rect 136 283 137 284
rect 135 283 136 284
rect 134 283 135 284
rect 133 283 134 284
rect 132 283 133 284
rect 131 283 132 284
rect 130 283 131 284
rect 124 283 125 284
rect 123 283 124 284
rect 122 283 123 284
rect 121 283 122 284
rect 120 283 121 284
rect 72 283 73 284
rect 71 283 72 284
rect 70 283 71 284
rect 69 283 70 284
rect 68 283 69 284
rect 67 283 68 284
rect 66 283 67 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 62 283 63 284
rect 61 283 62 284
rect 60 283 61 284
rect 59 283 60 284
rect 58 283 59 284
rect 57 283 58 284
rect 56 283 57 284
rect 55 283 56 284
rect 54 283 55 284
rect 53 283 54 284
rect 52 283 53 284
rect 51 283 52 284
rect 50 283 51 284
rect 49 283 50 284
rect 48 283 49 284
rect 47 283 48 284
rect 46 283 47 284
rect 143 284 144 285
rect 142 284 143 285
rect 141 284 142 285
rect 140 284 141 285
rect 139 284 140 285
rect 138 284 139 285
rect 137 284 138 285
rect 136 284 137 285
rect 135 284 136 285
rect 134 284 135 285
rect 133 284 134 285
rect 132 284 133 285
rect 131 284 132 285
rect 130 284 131 285
rect 124 284 125 285
rect 123 284 124 285
rect 122 284 123 285
rect 121 284 122 285
rect 120 284 121 285
rect 70 284 71 285
rect 69 284 70 285
rect 68 284 69 285
rect 67 284 68 285
rect 66 284 67 285
rect 65 284 66 285
rect 64 284 65 285
rect 63 284 64 285
rect 62 284 63 285
rect 61 284 62 285
rect 60 284 61 285
rect 59 284 60 285
rect 58 284 59 285
rect 57 284 58 285
rect 56 284 57 285
rect 55 284 56 285
rect 54 284 55 285
rect 53 284 54 285
rect 52 284 53 285
rect 51 284 52 285
rect 50 284 51 285
rect 49 284 50 285
rect 48 284 49 285
rect 142 285 143 286
rect 141 285 142 286
rect 140 285 141 286
rect 139 285 140 286
rect 138 285 139 286
rect 137 285 138 286
rect 136 285 137 286
rect 135 285 136 286
rect 134 285 135 286
rect 133 285 134 286
rect 132 285 133 286
rect 131 285 132 286
rect 130 285 131 286
rect 68 285 69 286
rect 67 285 68 286
rect 66 285 67 286
rect 65 285 66 286
rect 64 285 65 286
rect 63 285 64 286
rect 62 285 63 286
rect 61 285 62 286
rect 60 285 61 286
rect 59 285 60 286
rect 58 285 59 286
rect 57 285 58 286
rect 56 285 57 286
rect 55 285 56 286
rect 54 285 55 286
rect 53 285 54 286
rect 52 285 53 286
rect 51 285 52 286
rect 50 285 51 286
rect 142 286 143 287
rect 141 286 142 287
rect 140 286 141 287
rect 139 286 140 287
rect 138 286 139 287
rect 137 286 138 287
rect 136 286 137 287
rect 135 286 136 287
rect 134 286 135 287
rect 133 286 134 287
rect 132 286 133 287
rect 131 286 132 287
rect 130 286 131 287
rect 64 286 65 287
rect 63 286 64 287
rect 62 286 63 287
rect 61 286 62 287
rect 60 286 61 287
rect 59 286 60 287
rect 58 286 59 287
rect 57 286 58 287
rect 56 286 57 287
rect 55 286 56 287
rect 54 286 55 287
rect 136 290 137 291
rect 135 290 136 291
rect 134 290 135 291
rect 139 291 140 292
rect 138 291 139 292
rect 137 291 138 292
rect 136 291 137 292
rect 135 291 136 292
rect 134 291 135 292
rect 133 291 134 292
rect 132 291 133 292
rect 131 291 132 292
rect 141 292 142 293
rect 140 292 141 293
rect 139 292 140 293
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 135 292 136 293
rect 134 292 135 293
rect 133 292 134 293
rect 132 292 133 293
rect 131 292 132 293
rect 130 292 131 293
rect 129 292 130 293
rect 142 293 143 294
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 136 293 137 294
rect 135 293 136 294
rect 134 293 135 294
rect 133 293 134 294
rect 132 293 133 294
rect 131 293 132 294
rect 130 293 131 294
rect 129 293 130 294
rect 128 293 129 294
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 137 294 138 295
rect 136 294 137 295
rect 135 294 136 295
rect 134 294 135 295
rect 133 294 134 295
rect 132 294 133 295
rect 131 294 132 295
rect 130 294 131 295
rect 129 294 130 295
rect 128 294 129 295
rect 127 294 128 295
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 138 295 139 296
rect 137 295 138 296
rect 136 295 137 296
rect 135 295 136 296
rect 134 295 135 296
rect 133 295 134 296
rect 132 295 133 296
rect 131 295 132 296
rect 130 295 131 296
rect 129 295 130 296
rect 128 295 129 296
rect 127 295 128 296
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 139 296 140 297
rect 138 296 139 297
rect 132 296 133 297
rect 131 296 132 297
rect 130 296 131 297
rect 129 296 130 297
rect 128 296 129 297
rect 127 296 128 297
rect 81 296 82 297
rect 80 296 81 297
rect 79 296 80 297
rect 78 296 79 297
rect 77 296 78 297
rect 76 296 77 297
rect 75 296 76 297
rect 74 296 75 297
rect 73 296 74 297
rect 72 296 73 297
rect 71 296 72 297
rect 70 296 71 297
rect 69 296 70 297
rect 68 296 69 297
rect 67 296 68 297
rect 66 296 67 297
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 140 297 141 298
rect 130 297 131 298
rect 129 297 130 298
rect 128 297 129 298
rect 127 297 128 298
rect 126 297 127 298
rect 81 297 82 298
rect 80 297 81 298
rect 79 297 80 298
rect 78 297 79 298
rect 77 297 78 298
rect 76 297 77 298
rect 75 297 76 298
rect 74 297 75 298
rect 73 297 74 298
rect 72 297 73 298
rect 71 297 72 298
rect 70 297 71 298
rect 69 297 70 298
rect 68 297 69 298
rect 67 297 68 298
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 141 298 142 299
rect 140 298 141 299
rect 130 298 131 299
rect 129 298 130 299
rect 128 298 129 299
rect 127 298 128 299
rect 126 298 127 299
rect 81 298 82 299
rect 80 298 81 299
rect 79 298 80 299
rect 78 298 79 299
rect 77 298 78 299
rect 76 298 77 299
rect 75 298 76 299
rect 74 298 75 299
rect 73 298 74 299
rect 72 298 73 299
rect 71 298 72 299
rect 70 298 71 299
rect 69 298 70 299
rect 68 298 69 299
rect 67 298 68 299
rect 55 298 56 299
rect 54 298 55 299
rect 53 298 54 299
rect 52 298 53 299
rect 51 298 52 299
rect 50 298 51 299
rect 49 298 50 299
rect 48 298 49 299
rect 47 298 48 299
rect 46 298 47 299
rect 45 298 46 299
rect 44 298 45 299
rect 43 298 44 299
rect 42 298 43 299
rect 41 298 42 299
rect 40 298 41 299
rect 144 299 145 300
rect 143 299 144 300
rect 142 299 143 300
rect 141 299 142 300
rect 129 299 130 300
rect 128 299 129 300
rect 127 299 128 300
rect 126 299 127 300
rect 81 299 82 300
rect 80 299 81 300
rect 79 299 80 300
rect 78 299 79 300
rect 77 299 78 300
rect 76 299 77 300
rect 75 299 76 300
rect 74 299 75 300
rect 73 299 74 300
rect 72 299 73 300
rect 71 299 72 300
rect 70 299 71 300
rect 69 299 70 300
rect 68 299 69 300
rect 67 299 68 300
rect 55 299 56 300
rect 54 299 55 300
rect 53 299 54 300
rect 52 299 53 300
rect 51 299 52 300
rect 50 299 51 300
rect 49 299 50 300
rect 48 299 49 300
rect 47 299 48 300
rect 46 299 47 300
rect 45 299 46 300
rect 44 299 45 300
rect 43 299 44 300
rect 42 299 43 300
rect 41 299 42 300
rect 40 299 41 300
rect 39 299 40 300
rect 38 299 39 300
rect 37 299 38 300
rect 36 299 37 300
rect 35 299 36 300
rect 34 299 35 300
rect 33 299 34 300
rect 32 299 33 300
rect 31 299 32 300
rect 30 299 31 300
rect 29 299 30 300
rect 28 299 29 300
rect 27 299 28 300
rect 26 299 27 300
rect 25 299 26 300
rect 24 299 25 300
rect 144 300 145 301
rect 143 300 144 301
rect 142 300 143 301
rect 141 300 142 301
rect 129 300 130 301
rect 128 300 129 301
rect 127 300 128 301
rect 126 300 127 301
rect 82 300 83 301
rect 81 300 82 301
rect 80 300 81 301
rect 79 300 80 301
rect 78 300 79 301
rect 77 300 78 301
rect 76 300 77 301
rect 75 300 76 301
rect 74 300 75 301
rect 73 300 74 301
rect 72 300 73 301
rect 71 300 72 301
rect 70 300 71 301
rect 69 300 70 301
rect 68 300 69 301
rect 54 300 55 301
rect 53 300 54 301
rect 52 300 53 301
rect 51 300 52 301
rect 50 300 51 301
rect 49 300 50 301
rect 48 300 49 301
rect 47 300 48 301
rect 46 300 47 301
rect 45 300 46 301
rect 44 300 45 301
rect 43 300 44 301
rect 42 300 43 301
rect 41 300 42 301
rect 40 300 41 301
rect 39 300 40 301
rect 38 300 39 301
rect 37 300 38 301
rect 36 300 37 301
rect 35 300 36 301
rect 34 300 35 301
rect 33 300 34 301
rect 32 300 33 301
rect 31 300 32 301
rect 30 300 31 301
rect 29 300 30 301
rect 28 300 29 301
rect 27 300 28 301
rect 26 300 27 301
rect 25 300 26 301
rect 24 300 25 301
rect 23 300 24 301
rect 22 300 23 301
rect 21 300 22 301
rect 20 300 21 301
rect 19 300 20 301
rect 18 300 19 301
rect 17 300 18 301
rect 16 300 17 301
rect 144 301 145 302
rect 143 301 144 302
rect 142 301 143 302
rect 141 301 142 302
rect 129 301 130 302
rect 128 301 129 302
rect 127 301 128 302
rect 126 301 127 302
rect 82 301 83 302
rect 81 301 82 302
rect 80 301 81 302
rect 79 301 80 302
rect 78 301 79 302
rect 77 301 78 302
rect 76 301 77 302
rect 75 301 76 302
rect 74 301 75 302
rect 73 301 74 302
rect 72 301 73 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 68 301 69 302
rect 54 301 55 302
rect 53 301 54 302
rect 52 301 53 302
rect 51 301 52 302
rect 50 301 51 302
rect 49 301 50 302
rect 48 301 49 302
rect 47 301 48 302
rect 46 301 47 302
rect 45 301 46 302
rect 44 301 45 302
rect 43 301 44 302
rect 42 301 43 302
rect 41 301 42 302
rect 40 301 41 302
rect 39 301 40 302
rect 38 301 39 302
rect 37 301 38 302
rect 36 301 37 302
rect 35 301 36 302
rect 34 301 35 302
rect 33 301 34 302
rect 32 301 33 302
rect 31 301 32 302
rect 30 301 31 302
rect 29 301 30 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 25 301 26 302
rect 24 301 25 302
rect 23 301 24 302
rect 22 301 23 302
rect 21 301 22 302
rect 20 301 21 302
rect 19 301 20 302
rect 18 301 19 302
rect 17 301 18 302
rect 16 301 17 302
rect 144 302 145 303
rect 143 302 144 303
rect 142 302 143 303
rect 141 302 142 303
rect 140 302 141 303
rect 130 302 131 303
rect 129 302 130 303
rect 128 302 129 303
rect 127 302 128 303
rect 126 302 127 303
rect 82 302 83 303
rect 81 302 82 303
rect 80 302 81 303
rect 79 302 80 303
rect 78 302 79 303
rect 77 302 78 303
rect 76 302 77 303
rect 75 302 76 303
rect 74 302 75 303
rect 73 302 74 303
rect 72 302 73 303
rect 71 302 72 303
rect 70 302 71 303
rect 69 302 70 303
rect 68 302 69 303
rect 54 302 55 303
rect 53 302 54 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 48 302 49 303
rect 47 302 48 303
rect 46 302 47 303
rect 45 302 46 303
rect 44 302 45 303
rect 43 302 44 303
rect 42 302 43 303
rect 41 302 42 303
rect 40 302 41 303
rect 39 302 40 303
rect 38 302 39 303
rect 37 302 38 303
rect 36 302 37 303
rect 35 302 36 303
rect 34 302 35 303
rect 33 302 34 303
rect 32 302 33 303
rect 31 302 32 303
rect 30 302 31 303
rect 29 302 30 303
rect 28 302 29 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 24 302 25 303
rect 23 302 24 303
rect 22 302 23 303
rect 21 302 22 303
rect 20 302 21 303
rect 19 302 20 303
rect 18 302 19 303
rect 17 302 18 303
rect 16 302 17 303
rect 144 303 145 304
rect 143 303 144 304
rect 142 303 143 304
rect 141 303 142 304
rect 140 303 141 304
rect 139 303 140 304
rect 131 303 132 304
rect 130 303 131 304
rect 129 303 130 304
rect 128 303 129 304
rect 127 303 128 304
rect 126 303 127 304
rect 82 303 83 304
rect 81 303 82 304
rect 80 303 81 304
rect 79 303 80 304
rect 78 303 79 304
rect 77 303 78 304
rect 76 303 77 304
rect 75 303 76 304
rect 74 303 75 304
rect 73 303 74 304
rect 72 303 73 304
rect 71 303 72 304
rect 70 303 71 304
rect 69 303 70 304
rect 68 303 69 304
rect 54 303 55 304
rect 53 303 54 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 48 303 49 304
rect 47 303 48 304
rect 46 303 47 304
rect 45 303 46 304
rect 44 303 45 304
rect 43 303 44 304
rect 42 303 43 304
rect 41 303 42 304
rect 40 303 41 304
rect 39 303 40 304
rect 38 303 39 304
rect 37 303 38 304
rect 36 303 37 304
rect 35 303 36 304
rect 34 303 35 304
rect 33 303 34 304
rect 32 303 33 304
rect 31 303 32 304
rect 30 303 31 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 26 303 27 304
rect 25 303 26 304
rect 24 303 25 304
rect 23 303 24 304
rect 22 303 23 304
rect 21 303 22 304
rect 20 303 21 304
rect 19 303 20 304
rect 18 303 19 304
rect 17 303 18 304
rect 16 303 17 304
rect 143 304 144 305
rect 142 304 143 305
rect 141 304 142 305
rect 140 304 141 305
rect 139 304 140 305
rect 138 304 139 305
rect 137 304 138 305
rect 133 304 134 305
rect 132 304 133 305
rect 131 304 132 305
rect 130 304 131 305
rect 129 304 130 305
rect 128 304 129 305
rect 127 304 128 305
rect 82 304 83 305
rect 81 304 82 305
rect 80 304 81 305
rect 79 304 80 305
rect 78 304 79 305
rect 77 304 78 305
rect 76 304 77 305
rect 75 304 76 305
rect 74 304 75 305
rect 73 304 74 305
rect 72 304 73 305
rect 71 304 72 305
rect 70 304 71 305
rect 69 304 70 305
rect 54 304 55 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 48 304 49 305
rect 47 304 48 305
rect 46 304 47 305
rect 45 304 46 305
rect 44 304 45 305
rect 43 304 44 305
rect 42 304 43 305
rect 41 304 42 305
rect 40 304 41 305
rect 39 304 40 305
rect 38 304 39 305
rect 37 304 38 305
rect 36 304 37 305
rect 35 304 36 305
rect 34 304 35 305
rect 33 304 34 305
rect 32 304 33 305
rect 31 304 32 305
rect 30 304 31 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 22 304 23 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 17 304 18 305
rect 16 304 17 305
rect 143 305 144 306
rect 142 305 143 306
rect 141 305 142 306
rect 140 305 141 306
rect 139 305 140 306
rect 138 305 139 306
rect 137 305 138 306
rect 136 305 137 306
rect 135 305 136 306
rect 134 305 135 306
rect 133 305 134 306
rect 132 305 133 306
rect 131 305 132 306
rect 130 305 131 306
rect 129 305 130 306
rect 128 305 129 306
rect 127 305 128 306
rect 82 305 83 306
rect 81 305 82 306
rect 80 305 81 306
rect 79 305 80 306
rect 78 305 79 306
rect 77 305 78 306
rect 76 305 77 306
rect 75 305 76 306
rect 74 305 75 306
rect 73 305 74 306
rect 72 305 73 306
rect 71 305 72 306
rect 70 305 71 306
rect 69 305 70 306
rect 54 305 55 306
rect 53 305 54 306
rect 52 305 53 306
rect 51 305 52 306
rect 50 305 51 306
rect 49 305 50 306
rect 48 305 49 306
rect 47 305 48 306
rect 46 305 47 306
rect 45 305 46 306
rect 44 305 45 306
rect 43 305 44 306
rect 42 305 43 306
rect 41 305 42 306
rect 40 305 41 306
rect 39 305 40 306
rect 38 305 39 306
rect 37 305 38 306
rect 36 305 37 306
rect 35 305 36 306
rect 34 305 35 306
rect 33 305 34 306
rect 32 305 33 306
rect 31 305 32 306
rect 30 305 31 306
rect 29 305 30 306
rect 28 305 29 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 17 305 18 306
rect 16 305 17 306
rect 142 306 143 307
rect 141 306 142 307
rect 140 306 141 307
rect 139 306 140 307
rect 138 306 139 307
rect 137 306 138 307
rect 136 306 137 307
rect 135 306 136 307
rect 134 306 135 307
rect 133 306 134 307
rect 132 306 133 307
rect 131 306 132 307
rect 130 306 131 307
rect 129 306 130 307
rect 128 306 129 307
rect 82 306 83 307
rect 81 306 82 307
rect 80 306 81 307
rect 79 306 80 307
rect 78 306 79 307
rect 77 306 78 307
rect 76 306 77 307
rect 75 306 76 307
rect 74 306 75 307
rect 73 306 74 307
rect 72 306 73 307
rect 71 306 72 307
rect 70 306 71 307
rect 69 306 70 307
rect 54 306 55 307
rect 53 306 54 307
rect 52 306 53 307
rect 51 306 52 307
rect 50 306 51 307
rect 49 306 50 307
rect 48 306 49 307
rect 47 306 48 307
rect 46 306 47 307
rect 45 306 46 307
rect 44 306 45 307
rect 43 306 44 307
rect 42 306 43 307
rect 41 306 42 307
rect 40 306 41 307
rect 39 306 40 307
rect 38 306 39 307
rect 37 306 38 307
rect 36 306 37 307
rect 35 306 36 307
rect 34 306 35 307
rect 33 306 34 307
rect 32 306 33 307
rect 31 306 32 307
rect 30 306 31 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 17 306 18 307
rect 16 306 17 307
rect 141 307 142 308
rect 140 307 141 308
rect 139 307 140 308
rect 138 307 139 308
rect 137 307 138 308
rect 136 307 137 308
rect 135 307 136 308
rect 134 307 135 308
rect 133 307 134 308
rect 132 307 133 308
rect 131 307 132 308
rect 130 307 131 308
rect 129 307 130 308
rect 128 307 129 308
rect 83 307 84 308
rect 82 307 83 308
rect 81 307 82 308
rect 80 307 81 308
rect 79 307 80 308
rect 78 307 79 308
rect 77 307 78 308
rect 76 307 77 308
rect 75 307 76 308
rect 74 307 75 308
rect 73 307 74 308
rect 72 307 73 308
rect 71 307 72 308
rect 70 307 71 308
rect 69 307 70 308
rect 54 307 55 308
rect 53 307 54 308
rect 52 307 53 308
rect 51 307 52 308
rect 50 307 51 308
rect 49 307 50 308
rect 48 307 49 308
rect 47 307 48 308
rect 46 307 47 308
rect 45 307 46 308
rect 44 307 45 308
rect 43 307 44 308
rect 42 307 43 308
rect 41 307 42 308
rect 40 307 41 308
rect 39 307 40 308
rect 38 307 39 308
rect 37 307 38 308
rect 36 307 37 308
rect 35 307 36 308
rect 34 307 35 308
rect 33 307 34 308
rect 32 307 33 308
rect 31 307 32 308
rect 30 307 31 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 17 307 18 308
rect 16 307 17 308
rect 140 308 141 309
rect 139 308 140 309
rect 138 308 139 309
rect 137 308 138 309
rect 136 308 137 309
rect 135 308 136 309
rect 134 308 135 309
rect 133 308 134 309
rect 132 308 133 309
rect 131 308 132 309
rect 130 308 131 309
rect 83 308 84 309
rect 82 308 83 309
rect 81 308 82 309
rect 80 308 81 309
rect 79 308 80 309
rect 78 308 79 309
rect 77 308 78 309
rect 76 308 77 309
rect 75 308 76 309
rect 74 308 75 309
rect 73 308 74 309
rect 72 308 73 309
rect 71 308 72 309
rect 70 308 71 309
rect 69 308 70 309
rect 54 308 55 309
rect 53 308 54 309
rect 52 308 53 309
rect 51 308 52 309
rect 50 308 51 309
rect 49 308 50 309
rect 48 308 49 309
rect 47 308 48 309
rect 46 308 47 309
rect 45 308 46 309
rect 44 308 45 309
rect 43 308 44 309
rect 42 308 43 309
rect 41 308 42 309
rect 40 308 41 309
rect 39 308 40 309
rect 38 308 39 309
rect 37 308 38 309
rect 36 308 37 309
rect 35 308 36 309
rect 34 308 35 309
rect 33 308 34 309
rect 32 308 33 309
rect 31 308 32 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 17 308 18 309
rect 16 308 17 309
rect 138 309 139 310
rect 137 309 138 310
rect 136 309 137 310
rect 135 309 136 310
rect 134 309 135 310
rect 133 309 134 310
rect 132 309 133 310
rect 131 309 132 310
rect 83 309 84 310
rect 82 309 83 310
rect 81 309 82 310
rect 80 309 81 310
rect 79 309 80 310
rect 78 309 79 310
rect 77 309 78 310
rect 76 309 77 310
rect 75 309 76 310
rect 74 309 75 310
rect 73 309 74 310
rect 72 309 73 310
rect 71 309 72 310
rect 70 309 71 310
rect 69 309 70 310
rect 54 309 55 310
rect 53 309 54 310
rect 52 309 53 310
rect 51 309 52 310
rect 50 309 51 310
rect 49 309 50 310
rect 48 309 49 310
rect 47 309 48 310
rect 46 309 47 310
rect 45 309 46 310
rect 44 309 45 310
rect 43 309 44 310
rect 42 309 43 310
rect 41 309 42 310
rect 40 309 41 310
rect 39 309 40 310
rect 38 309 39 310
rect 37 309 38 310
rect 36 309 37 310
rect 35 309 36 310
rect 34 309 35 310
rect 33 309 34 310
rect 32 309 33 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 17 309 18 310
rect 16 309 17 310
rect 83 310 84 311
rect 82 310 83 311
rect 81 310 82 311
rect 80 310 81 311
rect 79 310 80 311
rect 78 310 79 311
rect 77 310 78 311
rect 76 310 77 311
rect 75 310 76 311
rect 74 310 75 311
rect 73 310 74 311
rect 72 310 73 311
rect 71 310 72 311
rect 70 310 71 311
rect 69 310 70 311
rect 54 310 55 311
rect 53 310 54 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 48 310 49 311
rect 47 310 48 311
rect 46 310 47 311
rect 45 310 46 311
rect 44 310 45 311
rect 43 310 44 311
rect 42 310 43 311
rect 41 310 42 311
rect 40 310 41 311
rect 39 310 40 311
rect 38 310 39 311
rect 37 310 38 311
rect 36 310 37 311
rect 35 310 36 311
rect 34 310 35 311
rect 33 310 34 311
rect 32 310 33 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 17 310 18 311
rect 16 310 17 311
rect 83 311 84 312
rect 82 311 83 312
rect 81 311 82 312
rect 80 311 81 312
rect 79 311 80 312
rect 78 311 79 312
rect 77 311 78 312
rect 76 311 77 312
rect 75 311 76 312
rect 74 311 75 312
rect 73 311 74 312
rect 72 311 73 312
rect 71 311 72 312
rect 70 311 71 312
rect 69 311 70 312
rect 54 311 55 312
rect 53 311 54 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 48 311 49 312
rect 47 311 48 312
rect 46 311 47 312
rect 45 311 46 312
rect 44 311 45 312
rect 43 311 44 312
rect 42 311 43 312
rect 41 311 42 312
rect 40 311 41 312
rect 39 311 40 312
rect 38 311 39 312
rect 37 311 38 312
rect 36 311 37 312
rect 35 311 36 312
rect 34 311 35 312
rect 33 311 34 312
rect 32 311 33 312
rect 31 311 32 312
rect 30 311 31 312
rect 29 311 30 312
rect 28 311 29 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 17 311 18 312
rect 16 311 17 312
rect 83 312 84 313
rect 82 312 83 313
rect 81 312 82 313
rect 80 312 81 313
rect 79 312 80 313
rect 78 312 79 313
rect 77 312 78 313
rect 76 312 77 313
rect 75 312 76 313
rect 74 312 75 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 70 312 71 313
rect 69 312 70 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 48 312 49 313
rect 47 312 48 313
rect 46 312 47 313
rect 45 312 46 313
rect 44 312 45 313
rect 43 312 44 313
rect 42 312 43 313
rect 41 312 42 313
rect 40 312 41 313
rect 39 312 40 313
rect 38 312 39 313
rect 37 312 38 313
rect 36 312 37 313
rect 35 312 36 313
rect 34 312 35 313
rect 33 312 34 313
rect 32 312 33 313
rect 31 312 32 313
rect 30 312 31 313
rect 29 312 30 313
rect 28 312 29 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 17 312 18 313
rect 16 312 17 313
rect 138 313 139 314
rect 137 313 138 314
rect 136 313 137 314
rect 135 313 136 314
rect 134 313 135 314
rect 133 313 134 314
rect 132 313 133 314
rect 83 313 84 314
rect 82 313 83 314
rect 81 313 82 314
rect 80 313 81 314
rect 79 313 80 314
rect 78 313 79 314
rect 77 313 78 314
rect 76 313 77 314
rect 75 313 76 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 70 313 71 314
rect 69 313 70 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 48 313 49 314
rect 47 313 48 314
rect 46 313 47 314
rect 45 313 46 314
rect 44 313 45 314
rect 43 313 44 314
rect 42 313 43 314
rect 41 313 42 314
rect 40 313 41 314
rect 39 313 40 314
rect 38 313 39 314
rect 37 313 38 314
rect 36 313 37 314
rect 35 313 36 314
rect 34 313 35 314
rect 33 313 34 314
rect 32 313 33 314
rect 31 313 32 314
rect 30 313 31 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 17 313 18 314
rect 16 313 17 314
rect 140 314 141 315
rect 139 314 140 315
rect 138 314 139 315
rect 137 314 138 315
rect 136 314 137 315
rect 135 314 136 315
rect 134 314 135 315
rect 133 314 134 315
rect 132 314 133 315
rect 131 314 132 315
rect 130 314 131 315
rect 83 314 84 315
rect 82 314 83 315
rect 81 314 82 315
rect 80 314 81 315
rect 79 314 80 315
rect 78 314 79 315
rect 77 314 78 315
rect 76 314 77 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 70 314 71 315
rect 69 314 70 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 48 314 49 315
rect 47 314 48 315
rect 46 314 47 315
rect 45 314 46 315
rect 44 314 45 315
rect 43 314 44 315
rect 42 314 43 315
rect 41 314 42 315
rect 40 314 41 315
rect 39 314 40 315
rect 38 314 39 315
rect 37 314 38 315
rect 36 314 37 315
rect 35 314 36 315
rect 34 314 35 315
rect 33 314 34 315
rect 32 314 33 315
rect 31 314 32 315
rect 30 314 31 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 17 314 18 315
rect 16 314 17 315
rect 141 315 142 316
rect 140 315 141 316
rect 139 315 140 316
rect 138 315 139 316
rect 137 315 138 316
rect 136 315 137 316
rect 135 315 136 316
rect 134 315 135 316
rect 133 315 134 316
rect 132 315 133 316
rect 131 315 132 316
rect 130 315 131 316
rect 129 315 130 316
rect 83 315 84 316
rect 82 315 83 316
rect 81 315 82 316
rect 80 315 81 316
rect 79 315 80 316
rect 78 315 79 316
rect 77 315 78 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 70 315 71 316
rect 69 315 70 316
rect 68 315 69 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 48 315 49 316
rect 47 315 48 316
rect 46 315 47 316
rect 45 315 46 316
rect 44 315 45 316
rect 43 315 44 316
rect 42 315 43 316
rect 41 315 42 316
rect 31 315 32 316
rect 30 315 31 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 17 315 18 316
rect 16 315 17 316
rect 142 316 143 317
rect 141 316 142 317
rect 140 316 141 317
rect 139 316 140 317
rect 138 316 139 317
rect 137 316 138 317
rect 136 316 137 317
rect 135 316 136 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 131 316 132 317
rect 130 316 131 317
rect 129 316 130 317
rect 128 316 129 317
rect 83 316 84 317
rect 82 316 83 317
rect 81 316 82 317
rect 80 316 81 317
rect 79 316 80 317
rect 78 316 79 317
rect 77 316 78 317
rect 76 316 77 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 70 316 71 317
rect 69 316 70 317
rect 68 316 69 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 48 316 49 317
rect 47 316 48 317
rect 46 316 47 317
rect 45 316 46 317
rect 44 316 45 317
rect 43 316 44 317
rect 42 316 43 317
rect 41 316 42 317
rect 31 316 32 317
rect 30 316 31 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 18 316 19 317
rect 17 316 18 317
rect 16 316 17 317
rect 143 317 144 318
rect 142 317 143 318
rect 141 317 142 318
rect 140 317 141 318
rect 139 317 140 318
rect 138 317 139 318
rect 137 317 138 318
rect 136 317 137 318
rect 135 317 136 318
rect 134 317 135 318
rect 133 317 134 318
rect 132 317 133 318
rect 131 317 132 318
rect 130 317 131 318
rect 129 317 130 318
rect 128 317 129 318
rect 127 317 128 318
rect 83 317 84 318
rect 82 317 83 318
rect 81 317 82 318
rect 80 317 81 318
rect 79 317 80 318
rect 78 317 79 318
rect 77 317 78 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 69 317 70 318
rect 68 317 69 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 48 317 49 318
rect 47 317 48 318
rect 46 317 47 318
rect 45 317 46 318
rect 44 317 45 318
rect 43 317 44 318
rect 42 317 43 318
rect 41 317 42 318
rect 31 317 32 318
rect 30 317 31 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 19 317 20 318
rect 18 317 19 318
rect 17 317 18 318
rect 16 317 17 318
rect 143 318 144 319
rect 142 318 143 319
rect 141 318 142 319
rect 140 318 141 319
rect 139 318 140 319
rect 138 318 139 319
rect 137 318 138 319
rect 136 318 137 319
rect 135 318 136 319
rect 134 318 135 319
rect 133 318 134 319
rect 132 318 133 319
rect 131 318 132 319
rect 130 318 131 319
rect 129 318 130 319
rect 128 318 129 319
rect 127 318 128 319
rect 83 318 84 319
rect 82 318 83 319
rect 81 318 82 319
rect 80 318 81 319
rect 79 318 80 319
rect 78 318 79 319
rect 77 318 78 319
rect 76 318 77 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 69 318 70 319
rect 68 318 69 319
rect 67 318 68 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 48 318 49 319
rect 47 318 48 319
rect 46 318 47 319
rect 45 318 46 319
rect 44 318 45 319
rect 43 318 44 319
rect 42 318 43 319
rect 41 318 42 319
rect 31 318 32 319
rect 30 318 31 319
rect 29 318 30 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 17 318 18 319
rect 16 318 17 319
rect 144 319 145 320
rect 143 319 144 320
rect 142 319 143 320
rect 141 319 142 320
rect 140 319 141 320
rect 139 319 140 320
rect 131 319 132 320
rect 130 319 131 320
rect 129 319 130 320
rect 128 319 129 320
rect 127 319 128 320
rect 126 319 127 320
rect 83 319 84 320
rect 82 319 83 320
rect 81 319 82 320
rect 80 319 81 320
rect 79 319 80 320
rect 78 319 79 320
rect 77 319 78 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 69 319 70 320
rect 68 319 69 320
rect 67 319 68 320
rect 66 319 67 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 48 319 49 320
rect 47 319 48 320
rect 46 319 47 320
rect 45 319 46 320
rect 44 319 45 320
rect 43 319 44 320
rect 42 319 43 320
rect 41 319 42 320
rect 31 319 32 320
rect 30 319 31 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 17 319 18 320
rect 16 319 17 320
rect 144 320 145 321
rect 143 320 144 321
rect 142 320 143 321
rect 141 320 142 321
rect 140 320 141 321
rect 130 320 131 321
rect 129 320 130 321
rect 128 320 129 321
rect 127 320 128 321
rect 126 320 127 321
rect 82 320 83 321
rect 81 320 82 321
rect 80 320 81 321
rect 79 320 80 321
rect 78 320 79 321
rect 77 320 78 321
rect 76 320 77 321
rect 75 320 76 321
rect 74 320 75 321
rect 73 320 74 321
rect 72 320 73 321
rect 71 320 72 321
rect 70 320 71 321
rect 69 320 70 321
rect 68 320 69 321
rect 67 320 68 321
rect 66 320 67 321
rect 65 320 66 321
rect 58 320 59 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 48 320 49 321
rect 47 320 48 321
rect 46 320 47 321
rect 45 320 46 321
rect 44 320 45 321
rect 43 320 44 321
rect 42 320 43 321
rect 41 320 42 321
rect 31 320 32 321
rect 30 320 31 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 17 320 18 321
rect 16 320 17 321
rect 144 321 145 322
rect 143 321 144 322
rect 142 321 143 322
rect 141 321 142 322
rect 140 321 141 322
rect 130 321 131 322
rect 129 321 130 322
rect 128 321 129 322
rect 127 321 128 322
rect 126 321 127 322
rect 82 321 83 322
rect 81 321 82 322
rect 80 321 81 322
rect 79 321 80 322
rect 78 321 79 322
rect 77 321 78 322
rect 76 321 77 322
rect 75 321 76 322
rect 74 321 75 322
rect 73 321 74 322
rect 72 321 73 322
rect 71 321 72 322
rect 70 321 71 322
rect 69 321 70 322
rect 68 321 69 322
rect 67 321 68 322
rect 66 321 67 322
rect 65 321 66 322
rect 64 321 65 322
rect 63 321 64 322
rect 62 321 63 322
rect 61 321 62 322
rect 60 321 61 322
rect 59 321 60 322
rect 58 321 59 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 48 321 49 322
rect 47 321 48 322
rect 46 321 47 322
rect 45 321 46 322
rect 44 321 45 322
rect 43 321 44 322
rect 42 321 43 322
rect 41 321 42 322
rect 31 321 32 322
rect 30 321 31 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 18 321 19 322
rect 17 321 18 322
rect 16 321 17 322
rect 144 322 145 323
rect 143 322 144 323
rect 142 322 143 323
rect 141 322 142 323
rect 129 322 130 323
rect 128 322 129 323
rect 127 322 128 323
rect 126 322 127 323
rect 82 322 83 323
rect 81 322 82 323
rect 80 322 81 323
rect 79 322 80 323
rect 78 322 79 323
rect 77 322 78 323
rect 76 322 77 323
rect 75 322 76 323
rect 74 322 75 323
rect 73 322 74 323
rect 72 322 73 323
rect 71 322 72 323
rect 70 322 71 323
rect 69 322 70 323
rect 68 322 69 323
rect 67 322 68 323
rect 66 322 67 323
rect 65 322 66 323
rect 64 322 65 323
rect 63 322 64 323
rect 62 322 63 323
rect 61 322 62 323
rect 60 322 61 323
rect 59 322 60 323
rect 58 322 59 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 48 322 49 323
rect 47 322 48 323
rect 46 322 47 323
rect 45 322 46 323
rect 44 322 45 323
rect 43 322 44 323
rect 42 322 43 323
rect 41 322 42 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 18 322 19 323
rect 17 322 18 323
rect 16 322 17 323
rect 144 323 145 324
rect 143 323 144 324
rect 142 323 143 324
rect 141 323 142 324
rect 129 323 130 324
rect 128 323 129 324
rect 127 323 128 324
rect 126 323 127 324
rect 82 323 83 324
rect 81 323 82 324
rect 80 323 81 324
rect 79 323 80 324
rect 78 323 79 324
rect 77 323 78 324
rect 76 323 77 324
rect 75 323 76 324
rect 74 323 75 324
rect 73 323 74 324
rect 72 323 73 324
rect 71 323 72 324
rect 70 323 71 324
rect 69 323 70 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 59 323 60 324
rect 58 323 59 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 48 323 49 324
rect 47 323 48 324
rect 46 323 47 324
rect 45 323 46 324
rect 44 323 45 324
rect 43 323 44 324
rect 42 323 43 324
rect 41 323 42 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 20 323 21 324
rect 19 323 20 324
rect 18 323 19 324
rect 17 323 18 324
rect 16 323 17 324
rect 144 324 145 325
rect 143 324 144 325
rect 142 324 143 325
rect 141 324 142 325
rect 140 324 141 325
rect 130 324 131 325
rect 129 324 130 325
rect 128 324 129 325
rect 127 324 128 325
rect 126 324 127 325
rect 81 324 82 325
rect 80 324 81 325
rect 79 324 80 325
rect 78 324 79 325
rect 77 324 78 325
rect 76 324 77 325
rect 75 324 76 325
rect 74 324 75 325
rect 73 324 74 325
rect 72 324 73 325
rect 71 324 72 325
rect 70 324 71 325
rect 69 324 70 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 59 324 60 325
rect 58 324 59 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 49 324 50 325
rect 48 324 49 325
rect 47 324 48 325
rect 46 324 47 325
rect 45 324 46 325
rect 44 324 45 325
rect 43 324 44 325
rect 42 324 43 325
rect 41 324 42 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 19 324 20 325
rect 18 324 19 325
rect 17 324 18 325
rect 16 324 17 325
rect 144 325 145 326
rect 143 325 144 326
rect 142 325 143 326
rect 141 325 142 326
rect 140 325 141 326
rect 130 325 131 326
rect 129 325 130 326
rect 128 325 129 326
rect 127 325 128 326
rect 126 325 127 326
rect 81 325 82 326
rect 80 325 81 326
rect 79 325 80 326
rect 78 325 79 326
rect 77 325 78 326
rect 76 325 77 326
rect 75 325 76 326
rect 74 325 75 326
rect 73 325 74 326
rect 72 325 73 326
rect 71 325 72 326
rect 70 325 71 326
rect 69 325 70 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 59 325 60 326
rect 58 325 59 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 49 325 50 326
rect 48 325 49 326
rect 47 325 48 326
rect 46 325 47 326
rect 45 325 46 326
rect 44 325 45 326
rect 43 325 44 326
rect 42 325 43 326
rect 31 325 32 326
rect 30 325 31 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 20 325 21 326
rect 19 325 20 326
rect 18 325 19 326
rect 17 325 18 326
rect 16 325 17 326
rect 144 326 145 327
rect 143 326 144 327
rect 142 326 143 327
rect 141 326 142 327
rect 140 326 141 327
rect 139 326 140 327
rect 131 326 132 327
rect 130 326 131 327
rect 129 326 130 327
rect 128 326 129 327
rect 127 326 128 327
rect 126 326 127 327
rect 81 326 82 327
rect 80 326 81 327
rect 79 326 80 327
rect 78 326 79 327
rect 77 326 78 327
rect 76 326 77 327
rect 75 326 76 327
rect 74 326 75 327
rect 73 326 74 327
rect 72 326 73 327
rect 71 326 72 327
rect 70 326 71 327
rect 69 326 70 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 59 326 60 327
rect 58 326 59 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 49 326 50 327
rect 48 326 49 327
rect 47 326 48 327
rect 46 326 47 327
rect 45 326 46 327
rect 44 326 45 327
rect 43 326 44 327
rect 42 326 43 327
rect 31 326 32 327
rect 30 326 31 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 21 326 22 327
rect 20 326 21 327
rect 19 326 20 327
rect 18 326 19 327
rect 17 326 18 327
rect 16 326 17 327
rect 143 327 144 328
rect 142 327 143 328
rect 141 327 142 328
rect 140 327 141 328
rect 139 327 140 328
rect 138 327 139 328
rect 137 327 138 328
rect 136 327 137 328
rect 135 327 136 328
rect 134 327 135 328
rect 133 327 134 328
rect 132 327 133 328
rect 131 327 132 328
rect 130 327 131 328
rect 129 327 130 328
rect 128 327 129 328
rect 127 327 128 328
rect 80 327 81 328
rect 79 327 80 328
rect 78 327 79 328
rect 77 327 78 328
rect 76 327 77 328
rect 75 327 76 328
rect 74 327 75 328
rect 73 327 74 328
rect 72 327 73 328
rect 71 327 72 328
rect 70 327 71 328
rect 69 327 70 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 61 327 62 328
rect 60 327 61 328
rect 59 327 60 328
rect 58 327 59 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 50 327 51 328
rect 49 327 50 328
rect 48 327 49 328
rect 47 327 48 328
rect 46 327 47 328
rect 45 327 46 328
rect 44 327 45 328
rect 43 327 44 328
rect 42 327 43 328
rect 31 327 32 328
rect 30 327 31 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 22 327 23 328
rect 21 327 22 328
rect 20 327 21 328
rect 19 327 20 328
rect 18 327 19 328
rect 17 327 18 328
rect 16 327 17 328
rect 143 328 144 329
rect 142 328 143 329
rect 141 328 142 329
rect 140 328 141 329
rect 139 328 140 329
rect 138 328 139 329
rect 137 328 138 329
rect 136 328 137 329
rect 135 328 136 329
rect 134 328 135 329
rect 133 328 134 329
rect 132 328 133 329
rect 131 328 132 329
rect 130 328 131 329
rect 129 328 130 329
rect 128 328 129 329
rect 127 328 128 329
rect 80 328 81 329
rect 79 328 80 329
rect 78 328 79 329
rect 77 328 78 329
rect 76 328 77 329
rect 75 328 76 329
rect 74 328 75 329
rect 73 328 74 329
rect 72 328 73 329
rect 71 328 72 329
rect 70 328 71 329
rect 69 328 70 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 61 328 62 329
rect 60 328 61 329
rect 59 328 60 329
rect 58 328 59 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 50 328 51 329
rect 49 328 50 329
rect 48 328 49 329
rect 47 328 48 329
rect 46 328 47 329
rect 45 328 46 329
rect 44 328 45 329
rect 43 328 44 329
rect 42 328 43 329
rect 31 328 32 329
rect 30 328 31 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 22 328 23 329
rect 21 328 22 329
rect 20 328 21 329
rect 19 328 20 329
rect 18 328 19 329
rect 17 328 18 329
rect 16 328 17 329
rect 142 329 143 330
rect 141 329 142 330
rect 140 329 141 330
rect 139 329 140 330
rect 138 329 139 330
rect 137 329 138 330
rect 136 329 137 330
rect 135 329 136 330
rect 134 329 135 330
rect 133 329 134 330
rect 132 329 133 330
rect 131 329 132 330
rect 130 329 131 330
rect 129 329 130 330
rect 128 329 129 330
rect 79 329 80 330
rect 78 329 79 330
rect 77 329 78 330
rect 76 329 77 330
rect 75 329 76 330
rect 74 329 75 330
rect 73 329 74 330
rect 72 329 73 330
rect 71 329 72 330
rect 70 329 71 330
rect 69 329 70 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 63 329 64 330
rect 62 329 63 330
rect 61 329 62 330
rect 60 329 61 330
rect 59 329 60 330
rect 58 329 59 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 51 329 52 330
rect 50 329 51 330
rect 49 329 50 330
rect 48 329 49 330
rect 47 329 48 330
rect 46 329 47 330
rect 45 329 46 330
rect 44 329 45 330
rect 43 329 44 330
rect 31 329 32 330
rect 30 329 31 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 23 329 24 330
rect 22 329 23 330
rect 21 329 22 330
rect 20 329 21 330
rect 19 329 20 330
rect 18 329 19 330
rect 17 329 18 330
rect 16 329 17 330
rect 141 330 142 331
rect 140 330 141 331
rect 139 330 140 331
rect 138 330 139 331
rect 137 330 138 331
rect 136 330 137 331
rect 135 330 136 331
rect 134 330 135 331
rect 133 330 134 331
rect 132 330 133 331
rect 131 330 132 331
rect 130 330 131 331
rect 129 330 130 331
rect 79 330 80 331
rect 78 330 79 331
rect 77 330 78 331
rect 76 330 77 331
rect 75 330 76 331
rect 74 330 75 331
rect 73 330 74 331
rect 72 330 73 331
rect 71 330 72 331
rect 70 330 71 331
rect 69 330 70 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 63 330 64 331
rect 62 330 63 331
rect 61 330 62 331
rect 60 330 61 331
rect 59 330 60 331
rect 58 330 59 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 51 330 52 331
rect 50 330 51 331
rect 49 330 50 331
rect 48 330 49 331
rect 47 330 48 331
rect 46 330 47 331
rect 45 330 46 331
rect 44 330 45 331
rect 43 330 44 331
rect 31 330 32 331
rect 30 330 31 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 24 330 25 331
rect 23 330 24 331
rect 22 330 23 331
rect 21 330 22 331
rect 20 330 21 331
rect 19 330 20 331
rect 18 330 19 331
rect 17 330 18 331
rect 16 330 17 331
rect 140 331 141 332
rect 139 331 140 332
rect 138 331 139 332
rect 137 331 138 332
rect 136 331 137 332
rect 135 331 136 332
rect 134 331 135 332
rect 133 331 134 332
rect 132 331 133 332
rect 131 331 132 332
rect 130 331 131 332
rect 78 331 79 332
rect 77 331 78 332
rect 76 331 77 332
rect 75 331 76 332
rect 74 331 75 332
rect 73 331 74 332
rect 72 331 73 332
rect 71 331 72 332
rect 70 331 71 332
rect 69 331 70 332
rect 68 331 69 332
rect 67 331 68 332
rect 66 331 67 332
rect 65 331 66 332
rect 64 331 65 332
rect 63 331 64 332
rect 62 331 63 332
rect 61 331 62 332
rect 60 331 61 332
rect 59 331 60 332
rect 58 331 59 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 52 331 53 332
rect 51 331 52 332
rect 50 331 51 332
rect 49 331 50 332
rect 48 331 49 332
rect 47 331 48 332
rect 46 331 47 332
rect 45 331 46 332
rect 44 331 45 332
rect 31 331 32 332
rect 30 331 31 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 26 331 27 332
rect 25 331 26 332
rect 24 331 25 332
rect 23 331 24 332
rect 22 331 23 332
rect 21 331 22 332
rect 20 331 21 332
rect 19 331 20 332
rect 18 331 19 332
rect 17 331 18 332
rect 16 331 17 332
rect 137 332 138 333
rect 136 332 137 333
rect 135 332 136 333
rect 134 332 135 333
rect 133 332 134 333
rect 132 332 133 333
rect 77 332 78 333
rect 76 332 77 333
rect 75 332 76 333
rect 74 332 75 333
rect 73 332 74 333
rect 72 332 73 333
rect 71 332 72 333
rect 70 332 71 333
rect 69 332 70 333
rect 68 332 69 333
rect 67 332 68 333
rect 66 332 67 333
rect 65 332 66 333
rect 64 332 65 333
rect 63 332 64 333
rect 62 332 63 333
rect 61 332 62 333
rect 60 332 61 333
rect 59 332 60 333
rect 58 332 59 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 52 332 53 333
rect 51 332 52 333
rect 50 332 51 333
rect 49 332 50 333
rect 48 332 49 333
rect 47 332 48 333
rect 46 332 47 333
rect 45 332 46 333
rect 44 332 45 333
rect 31 332 32 333
rect 30 332 31 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 26 332 27 333
rect 25 332 26 333
rect 24 332 25 333
rect 23 332 24 333
rect 22 332 23 333
rect 21 332 22 333
rect 20 332 21 333
rect 19 332 20 333
rect 18 332 19 333
rect 17 332 18 333
rect 16 332 17 333
rect 77 333 78 334
rect 76 333 77 334
rect 75 333 76 334
rect 74 333 75 334
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 52 333 53 334
rect 51 333 52 334
rect 50 333 51 334
rect 49 333 50 334
rect 48 333 49 334
rect 47 333 48 334
rect 46 333 47 334
rect 45 333 46 334
rect 31 333 32 334
rect 30 333 31 334
rect 29 333 30 334
rect 28 333 29 334
rect 27 333 28 334
rect 26 333 27 334
rect 25 333 26 334
rect 24 333 25 334
rect 23 333 24 334
rect 22 333 23 334
rect 21 333 22 334
rect 20 333 21 334
rect 19 333 20 334
rect 18 333 19 334
rect 17 333 18 334
rect 16 333 17 334
rect 76 334 77 335
rect 75 334 76 335
rect 74 334 75 335
rect 73 334 74 335
rect 72 334 73 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 52 334 53 335
rect 51 334 52 335
rect 50 334 51 335
rect 49 334 50 335
rect 48 334 49 335
rect 47 334 48 335
rect 46 334 47 335
rect 31 334 32 335
rect 30 334 31 335
rect 29 334 30 335
rect 28 334 29 335
rect 27 334 28 335
rect 26 334 27 335
rect 25 334 26 335
rect 24 334 25 335
rect 23 334 24 335
rect 22 334 23 335
rect 21 334 22 335
rect 20 334 21 335
rect 19 334 20 335
rect 18 334 19 335
rect 17 334 18 335
rect 16 334 17 335
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 52 335 53 336
rect 51 335 52 336
rect 50 335 51 336
rect 49 335 50 336
rect 48 335 49 336
rect 47 335 48 336
rect 46 335 47 336
rect 31 335 32 336
rect 30 335 31 336
rect 29 335 30 336
rect 28 335 29 336
rect 27 335 28 336
rect 26 335 27 336
rect 25 335 26 336
rect 24 335 25 336
rect 23 335 24 336
rect 22 335 23 336
rect 21 335 22 336
rect 20 335 21 336
rect 19 335 20 336
rect 18 335 19 336
rect 17 335 18 336
rect 16 335 17 336
rect 138 336 139 337
rect 137 336 138 337
rect 136 336 137 337
rect 135 336 136 337
rect 134 336 135 337
rect 133 336 134 337
rect 132 336 133 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 52 336 53 337
rect 51 336 52 337
rect 50 336 51 337
rect 49 336 50 337
rect 48 336 49 337
rect 31 336 32 337
rect 30 336 31 337
rect 29 336 30 337
rect 28 336 29 337
rect 27 336 28 337
rect 26 336 27 337
rect 25 336 26 337
rect 24 336 25 337
rect 23 336 24 337
rect 22 336 23 337
rect 21 336 22 337
rect 20 336 21 337
rect 19 336 20 337
rect 18 336 19 337
rect 17 336 18 337
rect 16 336 17 337
rect 141 337 142 338
rect 140 337 141 338
rect 139 337 140 338
rect 138 337 139 338
rect 137 337 138 338
rect 136 337 137 338
rect 135 337 136 338
rect 134 337 135 338
rect 133 337 134 338
rect 132 337 133 338
rect 131 337 132 338
rect 130 337 131 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 52 337 53 338
rect 51 337 52 338
rect 50 337 51 338
rect 49 337 50 338
rect 31 337 32 338
rect 30 337 31 338
rect 29 337 30 338
rect 28 337 29 338
rect 27 337 28 338
rect 26 337 27 338
rect 25 337 26 338
rect 24 337 25 338
rect 23 337 24 338
rect 22 337 23 338
rect 21 337 22 338
rect 20 337 21 338
rect 19 337 20 338
rect 18 337 19 338
rect 17 337 18 338
rect 16 337 17 338
rect 142 338 143 339
rect 141 338 142 339
rect 140 338 141 339
rect 139 338 140 339
rect 138 338 139 339
rect 137 338 138 339
rect 136 338 137 339
rect 135 338 136 339
rect 134 338 135 339
rect 133 338 134 339
rect 132 338 133 339
rect 131 338 132 339
rect 130 338 131 339
rect 129 338 130 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 53 338 54 339
rect 52 338 53 339
rect 51 338 52 339
rect 50 338 51 339
rect 143 339 144 340
rect 142 339 143 340
rect 141 339 142 340
rect 140 339 141 340
rect 139 339 140 340
rect 138 339 139 340
rect 137 339 138 340
rect 136 339 137 340
rect 135 339 136 340
rect 134 339 135 340
rect 133 339 134 340
rect 132 339 133 340
rect 131 339 132 340
rect 130 339 131 340
rect 129 339 130 340
rect 128 339 129 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 54 339 55 340
rect 53 339 54 340
rect 143 340 144 341
rect 142 340 143 341
rect 141 340 142 341
rect 140 340 141 341
rect 139 340 140 341
rect 138 340 139 341
rect 137 340 138 341
rect 136 340 137 341
rect 135 340 136 341
rect 134 340 135 341
rect 133 340 134 341
rect 132 340 133 341
rect 131 340 132 341
rect 130 340 131 341
rect 129 340 130 341
rect 128 340 129 341
rect 127 340 128 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 144 341 145 342
rect 143 341 144 342
rect 142 341 143 342
rect 141 341 142 342
rect 140 341 141 342
rect 139 341 140 342
rect 138 341 139 342
rect 137 341 138 342
rect 136 341 137 342
rect 135 341 136 342
rect 134 341 135 342
rect 133 341 134 342
rect 132 341 133 342
rect 131 341 132 342
rect 130 341 131 342
rect 129 341 130 342
rect 128 341 129 342
rect 127 341 128 342
rect 144 342 145 343
rect 143 342 144 343
rect 142 342 143 343
rect 141 342 142 343
rect 140 342 141 343
rect 139 342 140 343
rect 131 342 132 343
rect 130 342 131 343
rect 129 342 130 343
rect 128 342 129 343
rect 127 342 128 343
rect 126 342 127 343
rect 144 343 145 344
rect 143 343 144 344
rect 142 343 143 344
rect 141 343 142 344
rect 140 343 141 344
rect 130 343 131 344
rect 129 343 130 344
rect 128 343 129 344
rect 127 343 128 344
rect 126 343 127 344
rect 144 344 145 345
rect 143 344 144 345
rect 142 344 143 345
rect 141 344 142 345
rect 140 344 141 345
rect 130 344 131 345
rect 129 344 130 345
rect 128 344 129 345
rect 127 344 128 345
rect 126 344 127 345
rect 144 345 145 346
rect 143 345 144 346
rect 142 345 143 346
rect 141 345 142 346
rect 129 345 130 346
rect 128 345 129 346
rect 127 345 128 346
rect 126 345 127 346
rect 143 346 144 347
rect 142 346 143 347
rect 141 346 142 347
rect 129 346 130 347
rect 128 346 129 347
rect 127 346 128 347
rect 126 346 127 347
rect 143 347 144 348
rect 142 347 143 348
rect 141 347 142 348
rect 140 347 141 348
rect 130 347 131 348
rect 129 347 130 348
rect 128 347 129 348
rect 127 347 128 348
rect 142 348 143 349
rect 141 348 142 349
rect 140 348 141 349
rect 139 348 140 349
rect 130 348 131 349
rect 129 348 130 349
rect 128 348 129 349
rect 127 348 128 349
rect 142 349 143 350
rect 141 349 142 350
rect 140 349 141 350
rect 139 349 140 350
rect 138 349 139 350
rect 137 349 138 350
rect 132 349 133 350
rect 131 349 132 350
rect 130 349 131 350
rect 129 349 130 350
rect 128 349 129 350
rect 144 350 145 351
rect 143 350 144 351
rect 142 350 143 351
rect 141 350 142 351
rect 140 350 141 351
rect 139 350 140 351
rect 138 350 139 351
rect 137 350 138 351
rect 136 350 137 351
rect 135 350 136 351
rect 134 350 135 351
rect 133 350 134 351
rect 132 350 133 351
rect 131 350 132 351
rect 130 350 131 351
rect 129 350 130 351
rect 128 350 129 351
rect 127 350 128 351
rect 126 350 127 351
rect 125 350 126 351
rect 124 350 125 351
rect 123 350 124 351
rect 122 350 123 351
rect 121 350 122 351
rect 120 350 121 351
rect 119 350 120 351
rect 118 350 119 351
rect 117 350 118 351
rect 55 350 56 351
rect 54 350 55 351
rect 53 350 54 351
rect 52 350 53 351
rect 51 350 52 351
rect 50 350 51 351
rect 49 350 50 351
rect 48 350 49 351
rect 47 350 48 351
rect 46 350 47 351
rect 45 350 46 351
rect 44 350 45 351
rect 144 351 145 352
rect 143 351 144 352
rect 142 351 143 352
rect 141 351 142 352
rect 140 351 141 352
rect 139 351 140 352
rect 138 351 139 352
rect 137 351 138 352
rect 136 351 137 352
rect 135 351 136 352
rect 134 351 135 352
rect 133 351 134 352
rect 132 351 133 352
rect 131 351 132 352
rect 130 351 131 352
rect 129 351 130 352
rect 128 351 129 352
rect 127 351 128 352
rect 126 351 127 352
rect 125 351 126 352
rect 124 351 125 352
rect 123 351 124 352
rect 122 351 123 352
rect 121 351 122 352
rect 120 351 121 352
rect 119 351 120 352
rect 118 351 119 352
rect 117 351 118 352
rect 63 351 64 352
rect 62 351 63 352
rect 61 351 62 352
rect 60 351 61 352
rect 59 351 60 352
rect 58 351 59 352
rect 57 351 58 352
rect 56 351 57 352
rect 55 351 56 352
rect 54 351 55 352
rect 53 351 54 352
rect 52 351 53 352
rect 51 351 52 352
rect 50 351 51 352
rect 49 351 50 352
rect 48 351 49 352
rect 47 351 48 352
rect 46 351 47 352
rect 45 351 46 352
rect 44 351 45 352
rect 43 351 44 352
rect 42 351 43 352
rect 41 351 42 352
rect 40 351 41 352
rect 39 351 40 352
rect 38 351 39 352
rect 37 351 38 352
rect 144 352 145 353
rect 143 352 144 353
rect 142 352 143 353
rect 141 352 142 353
rect 140 352 141 353
rect 139 352 140 353
rect 138 352 139 353
rect 137 352 138 353
rect 136 352 137 353
rect 135 352 136 353
rect 134 352 135 353
rect 133 352 134 353
rect 132 352 133 353
rect 131 352 132 353
rect 130 352 131 353
rect 129 352 130 353
rect 128 352 129 353
rect 127 352 128 353
rect 126 352 127 353
rect 125 352 126 353
rect 124 352 125 353
rect 123 352 124 353
rect 122 352 123 353
rect 121 352 122 353
rect 120 352 121 353
rect 119 352 120 353
rect 118 352 119 353
rect 117 352 118 353
rect 67 352 68 353
rect 66 352 67 353
rect 65 352 66 353
rect 64 352 65 353
rect 63 352 64 353
rect 62 352 63 353
rect 61 352 62 353
rect 60 352 61 353
rect 59 352 60 353
rect 58 352 59 353
rect 57 352 58 353
rect 56 352 57 353
rect 55 352 56 353
rect 54 352 55 353
rect 53 352 54 353
rect 52 352 53 353
rect 51 352 52 353
rect 50 352 51 353
rect 49 352 50 353
rect 48 352 49 353
rect 47 352 48 353
rect 46 352 47 353
rect 45 352 46 353
rect 44 352 45 353
rect 43 352 44 353
rect 42 352 43 353
rect 41 352 42 353
rect 40 352 41 353
rect 39 352 40 353
rect 38 352 39 353
rect 37 352 38 353
rect 36 352 37 353
rect 35 352 36 353
rect 34 352 35 353
rect 33 352 34 353
rect 144 353 145 354
rect 143 353 144 354
rect 142 353 143 354
rect 141 353 142 354
rect 140 353 141 354
rect 139 353 140 354
rect 138 353 139 354
rect 137 353 138 354
rect 136 353 137 354
rect 135 353 136 354
rect 134 353 135 354
rect 133 353 134 354
rect 132 353 133 354
rect 131 353 132 354
rect 130 353 131 354
rect 129 353 130 354
rect 128 353 129 354
rect 127 353 128 354
rect 126 353 127 354
rect 125 353 126 354
rect 124 353 125 354
rect 123 353 124 354
rect 122 353 123 354
rect 121 353 122 354
rect 120 353 121 354
rect 119 353 120 354
rect 118 353 119 354
rect 117 353 118 354
rect 69 353 70 354
rect 68 353 69 354
rect 67 353 68 354
rect 66 353 67 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 61 353 62 354
rect 60 353 61 354
rect 59 353 60 354
rect 58 353 59 354
rect 57 353 58 354
rect 56 353 57 354
rect 55 353 56 354
rect 54 353 55 354
rect 53 353 54 354
rect 52 353 53 354
rect 51 353 52 354
rect 50 353 51 354
rect 49 353 50 354
rect 48 353 49 354
rect 47 353 48 354
rect 46 353 47 354
rect 45 353 46 354
rect 44 353 45 354
rect 43 353 44 354
rect 42 353 43 354
rect 41 353 42 354
rect 40 353 41 354
rect 39 353 40 354
rect 38 353 39 354
rect 37 353 38 354
rect 36 353 37 354
rect 35 353 36 354
rect 34 353 35 354
rect 33 353 34 354
rect 32 353 33 354
rect 31 353 32 354
rect 30 353 31 354
rect 144 354 145 355
rect 143 354 144 355
rect 142 354 143 355
rect 141 354 142 355
rect 140 354 141 355
rect 139 354 140 355
rect 138 354 139 355
rect 137 354 138 355
rect 136 354 137 355
rect 135 354 136 355
rect 134 354 135 355
rect 133 354 134 355
rect 132 354 133 355
rect 131 354 132 355
rect 130 354 131 355
rect 129 354 130 355
rect 128 354 129 355
rect 127 354 128 355
rect 126 354 127 355
rect 125 354 126 355
rect 124 354 125 355
rect 123 354 124 355
rect 122 354 123 355
rect 121 354 122 355
rect 120 354 121 355
rect 119 354 120 355
rect 118 354 119 355
rect 117 354 118 355
rect 71 354 72 355
rect 70 354 71 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 62 354 63 355
rect 61 354 62 355
rect 60 354 61 355
rect 59 354 60 355
rect 58 354 59 355
rect 57 354 58 355
rect 56 354 57 355
rect 55 354 56 355
rect 54 354 55 355
rect 53 354 54 355
rect 52 354 53 355
rect 51 354 52 355
rect 50 354 51 355
rect 49 354 50 355
rect 48 354 49 355
rect 47 354 48 355
rect 46 354 47 355
rect 45 354 46 355
rect 44 354 45 355
rect 43 354 44 355
rect 42 354 43 355
rect 41 354 42 355
rect 40 354 41 355
rect 39 354 40 355
rect 38 354 39 355
rect 37 354 38 355
rect 36 354 37 355
rect 35 354 36 355
rect 34 354 35 355
rect 33 354 34 355
rect 32 354 33 355
rect 31 354 32 355
rect 30 354 31 355
rect 29 354 30 355
rect 28 354 29 355
rect 73 355 74 356
rect 72 355 73 356
rect 71 355 72 356
rect 70 355 71 356
rect 69 355 70 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 63 355 64 356
rect 62 355 63 356
rect 61 355 62 356
rect 60 355 61 356
rect 59 355 60 356
rect 58 355 59 356
rect 57 355 58 356
rect 56 355 57 356
rect 55 355 56 356
rect 54 355 55 356
rect 53 355 54 356
rect 52 355 53 356
rect 51 355 52 356
rect 50 355 51 356
rect 49 355 50 356
rect 48 355 49 356
rect 47 355 48 356
rect 46 355 47 356
rect 45 355 46 356
rect 44 355 45 356
rect 43 355 44 356
rect 42 355 43 356
rect 41 355 42 356
rect 40 355 41 356
rect 39 355 40 356
rect 38 355 39 356
rect 37 355 38 356
rect 36 355 37 356
rect 35 355 36 356
rect 34 355 35 356
rect 33 355 34 356
rect 32 355 33 356
rect 31 355 32 356
rect 30 355 31 356
rect 29 355 30 356
rect 28 355 29 356
rect 27 355 28 356
rect 26 355 27 356
rect 75 356 76 357
rect 74 356 75 357
rect 73 356 74 357
rect 72 356 73 357
rect 71 356 72 357
rect 70 356 71 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 64 356 65 357
rect 63 356 64 357
rect 62 356 63 357
rect 61 356 62 357
rect 60 356 61 357
rect 59 356 60 357
rect 58 356 59 357
rect 57 356 58 357
rect 56 356 57 357
rect 55 356 56 357
rect 54 356 55 357
rect 53 356 54 357
rect 52 356 53 357
rect 51 356 52 357
rect 50 356 51 357
rect 49 356 50 357
rect 48 356 49 357
rect 47 356 48 357
rect 46 356 47 357
rect 45 356 46 357
rect 44 356 45 357
rect 43 356 44 357
rect 42 356 43 357
rect 41 356 42 357
rect 40 356 41 357
rect 39 356 40 357
rect 38 356 39 357
rect 37 356 38 357
rect 36 356 37 357
rect 35 356 36 357
rect 34 356 35 357
rect 33 356 34 357
rect 32 356 33 357
rect 31 356 32 357
rect 30 356 31 357
rect 29 356 30 357
rect 28 356 29 357
rect 27 356 28 357
rect 26 356 27 357
rect 25 356 26 357
rect 76 357 77 358
rect 75 357 76 358
rect 74 357 75 358
rect 73 357 74 358
rect 72 357 73 358
rect 71 357 72 358
rect 70 357 71 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 65 357 66 358
rect 64 357 65 358
rect 63 357 64 358
rect 62 357 63 358
rect 61 357 62 358
rect 60 357 61 358
rect 59 357 60 358
rect 58 357 59 358
rect 57 357 58 358
rect 56 357 57 358
rect 55 357 56 358
rect 54 357 55 358
rect 53 357 54 358
rect 52 357 53 358
rect 51 357 52 358
rect 50 357 51 358
rect 49 357 50 358
rect 48 357 49 358
rect 47 357 48 358
rect 46 357 47 358
rect 45 357 46 358
rect 44 357 45 358
rect 43 357 44 358
rect 42 357 43 358
rect 41 357 42 358
rect 40 357 41 358
rect 39 357 40 358
rect 38 357 39 358
rect 37 357 38 358
rect 36 357 37 358
rect 35 357 36 358
rect 34 357 35 358
rect 33 357 34 358
rect 32 357 33 358
rect 31 357 32 358
rect 30 357 31 358
rect 29 357 30 358
rect 28 357 29 358
rect 27 357 28 358
rect 26 357 27 358
rect 25 357 26 358
rect 24 357 25 358
rect 77 358 78 359
rect 76 358 77 359
rect 75 358 76 359
rect 74 358 75 359
rect 73 358 74 359
rect 72 358 73 359
rect 71 358 72 359
rect 70 358 71 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 66 358 67 359
rect 65 358 66 359
rect 64 358 65 359
rect 63 358 64 359
rect 62 358 63 359
rect 61 358 62 359
rect 60 358 61 359
rect 59 358 60 359
rect 58 358 59 359
rect 57 358 58 359
rect 56 358 57 359
rect 55 358 56 359
rect 54 358 55 359
rect 53 358 54 359
rect 52 358 53 359
rect 51 358 52 359
rect 50 358 51 359
rect 49 358 50 359
rect 48 358 49 359
rect 47 358 48 359
rect 46 358 47 359
rect 45 358 46 359
rect 44 358 45 359
rect 43 358 44 359
rect 42 358 43 359
rect 41 358 42 359
rect 40 358 41 359
rect 39 358 40 359
rect 38 358 39 359
rect 37 358 38 359
rect 36 358 37 359
rect 35 358 36 359
rect 34 358 35 359
rect 33 358 34 359
rect 32 358 33 359
rect 31 358 32 359
rect 30 358 31 359
rect 29 358 30 359
rect 28 358 29 359
rect 27 358 28 359
rect 26 358 27 359
rect 25 358 26 359
rect 24 358 25 359
rect 23 358 24 359
rect 22 358 23 359
rect 78 359 79 360
rect 77 359 78 360
rect 76 359 77 360
rect 75 359 76 360
rect 74 359 75 360
rect 73 359 74 360
rect 72 359 73 360
rect 71 359 72 360
rect 70 359 71 360
rect 69 359 70 360
rect 68 359 69 360
rect 67 359 68 360
rect 66 359 67 360
rect 65 359 66 360
rect 64 359 65 360
rect 63 359 64 360
rect 62 359 63 360
rect 61 359 62 360
rect 60 359 61 360
rect 59 359 60 360
rect 58 359 59 360
rect 57 359 58 360
rect 56 359 57 360
rect 55 359 56 360
rect 54 359 55 360
rect 53 359 54 360
rect 52 359 53 360
rect 51 359 52 360
rect 50 359 51 360
rect 49 359 50 360
rect 48 359 49 360
rect 47 359 48 360
rect 46 359 47 360
rect 45 359 46 360
rect 44 359 45 360
rect 43 359 44 360
rect 42 359 43 360
rect 41 359 42 360
rect 40 359 41 360
rect 39 359 40 360
rect 38 359 39 360
rect 37 359 38 360
rect 36 359 37 360
rect 35 359 36 360
rect 34 359 35 360
rect 33 359 34 360
rect 32 359 33 360
rect 31 359 32 360
rect 30 359 31 360
rect 29 359 30 360
rect 28 359 29 360
rect 27 359 28 360
rect 26 359 27 360
rect 25 359 26 360
rect 24 359 25 360
rect 23 359 24 360
rect 22 359 23 360
rect 21 359 22 360
rect 79 360 80 361
rect 78 360 79 361
rect 77 360 78 361
rect 76 360 77 361
rect 75 360 76 361
rect 74 360 75 361
rect 73 360 74 361
rect 72 360 73 361
rect 71 360 72 361
rect 70 360 71 361
rect 69 360 70 361
rect 68 360 69 361
rect 67 360 68 361
rect 66 360 67 361
rect 65 360 66 361
rect 64 360 65 361
rect 63 360 64 361
rect 62 360 63 361
rect 61 360 62 361
rect 60 360 61 361
rect 59 360 60 361
rect 58 360 59 361
rect 57 360 58 361
rect 56 360 57 361
rect 55 360 56 361
rect 54 360 55 361
rect 53 360 54 361
rect 52 360 53 361
rect 51 360 52 361
rect 50 360 51 361
rect 49 360 50 361
rect 48 360 49 361
rect 47 360 48 361
rect 46 360 47 361
rect 45 360 46 361
rect 44 360 45 361
rect 43 360 44 361
rect 42 360 43 361
rect 41 360 42 361
rect 40 360 41 361
rect 39 360 40 361
rect 38 360 39 361
rect 37 360 38 361
rect 36 360 37 361
rect 35 360 36 361
rect 34 360 35 361
rect 33 360 34 361
rect 32 360 33 361
rect 31 360 32 361
rect 30 360 31 361
rect 29 360 30 361
rect 28 360 29 361
rect 27 360 28 361
rect 26 360 27 361
rect 25 360 26 361
rect 24 360 25 361
rect 23 360 24 361
rect 22 360 23 361
rect 21 360 22 361
rect 20 360 21 361
rect 144 361 145 362
rect 143 361 144 362
rect 142 361 143 362
rect 141 361 142 362
rect 140 361 141 362
rect 139 361 140 362
rect 138 361 139 362
rect 137 361 138 362
rect 136 361 137 362
rect 135 361 136 362
rect 134 361 135 362
rect 133 361 134 362
rect 132 361 133 362
rect 131 361 132 362
rect 130 361 131 362
rect 129 361 130 362
rect 128 361 129 362
rect 127 361 128 362
rect 126 361 127 362
rect 125 361 126 362
rect 124 361 125 362
rect 123 361 124 362
rect 122 361 123 362
rect 121 361 122 362
rect 120 361 121 362
rect 119 361 120 362
rect 79 361 80 362
rect 78 361 79 362
rect 77 361 78 362
rect 76 361 77 362
rect 75 361 76 362
rect 74 361 75 362
rect 73 361 74 362
rect 72 361 73 362
rect 71 361 72 362
rect 70 361 71 362
rect 69 361 70 362
rect 68 361 69 362
rect 67 361 68 362
rect 66 361 67 362
rect 65 361 66 362
rect 64 361 65 362
rect 63 361 64 362
rect 62 361 63 362
rect 61 361 62 362
rect 60 361 61 362
rect 59 361 60 362
rect 58 361 59 362
rect 57 361 58 362
rect 56 361 57 362
rect 55 361 56 362
rect 54 361 55 362
rect 53 361 54 362
rect 52 361 53 362
rect 51 361 52 362
rect 50 361 51 362
rect 49 361 50 362
rect 48 361 49 362
rect 47 361 48 362
rect 46 361 47 362
rect 45 361 46 362
rect 44 361 45 362
rect 43 361 44 362
rect 42 361 43 362
rect 41 361 42 362
rect 40 361 41 362
rect 39 361 40 362
rect 38 361 39 362
rect 37 361 38 362
rect 36 361 37 362
rect 35 361 36 362
rect 34 361 35 362
rect 33 361 34 362
rect 32 361 33 362
rect 31 361 32 362
rect 30 361 31 362
rect 29 361 30 362
rect 28 361 29 362
rect 27 361 28 362
rect 26 361 27 362
rect 25 361 26 362
rect 24 361 25 362
rect 23 361 24 362
rect 22 361 23 362
rect 21 361 22 362
rect 20 361 21 362
rect 144 362 145 363
rect 143 362 144 363
rect 142 362 143 363
rect 141 362 142 363
rect 140 362 141 363
rect 139 362 140 363
rect 138 362 139 363
rect 137 362 138 363
rect 136 362 137 363
rect 135 362 136 363
rect 134 362 135 363
rect 133 362 134 363
rect 132 362 133 363
rect 131 362 132 363
rect 130 362 131 363
rect 129 362 130 363
rect 128 362 129 363
rect 127 362 128 363
rect 126 362 127 363
rect 125 362 126 363
rect 124 362 125 363
rect 123 362 124 363
rect 122 362 123 363
rect 121 362 122 363
rect 120 362 121 363
rect 119 362 120 363
rect 80 362 81 363
rect 79 362 80 363
rect 78 362 79 363
rect 77 362 78 363
rect 76 362 77 363
rect 75 362 76 363
rect 74 362 75 363
rect 73 362 74 363
rect 72 362 73 363
rect 71 362 72 363
rect 70 362 71 363
rect 69 362 70 363
rect 68 362 69 363
rect 67 362 68 363
rect 66 362 67 363
rect 65 362 66 363
rect 64 362 65 363
rect 63 362 64 363
rect 62 362 63 363
rect 61 362 62 363
rect 60 362 61 363
rect 59 362 60 363
rect 58 362 59 363
rect 57 362 58 363
rect 56 362 57 363
rect 55 362 56 363
rect 54 362 55 363
rect 53 362 54 363
rect 52 362 53 363
rect 51 362 52 363
rect 50 362 51 363
rect 49 362 50 363
rect 48 362 49 363
rect 47 362 48 363
rect 46 362 47 363
rect 45 362 46 363
rect 44 362 45 363
rect 43 362 44 363
rect 42 362 43 363
rect 41 362 42 363
rect 40 362 41 363
rect 39 362 40 363
rect 38 362 39 363
rect 37 362 38 363
rect 36 362 37 363
rect 35 362 36 363
rect 34 362 35 363
rect 33 362 34 363
rect 32 362 33 363
rect 31 362 32 363
rect 30 362 31 363
rect 29 362 30 363
rect 28 362 29 363
rect 27 362 28 363
rect 26 362 27 363
rect 25 362 26 363
rect 24 362 25 363
rect 23 362 24 363
rect 22 362 23 363
rect 21 362 22 363
rect 20 362 21 363
rect 19 362 20 363
rect 144 363 145 364
rect 143 363 144 364
rect 142 363 143 364
rect 141 363 142 364
rect 140 363 141 364
rect 139 363 140 364
rect 138 363 139 364
rect 137 363 138 364
rect 136 363 137 364
rect 135 363 136 364
rect 134 363 135 364
rect 133 363 134 364
rect 132 363 133 364
rect 131 363 132 364
rect 130 363 131 364
rect 129 363 130 364
rect 128 363 129 364
rect 127 363 128 364
rect 126 363 127 364
rect 125 363 126 364
rect 124 363 125 364
rect 123 363 124 364
rect 122 363 123 364
rect 121 363 122 364
rect 120 363 121 364
rect 119 363 120 364
rect 80 363 81 364
rect 79 363 80 364
rect 78 363 79 364
rect 77 363 78 364
rect 76 363 77 364
rect 75 363 76 364
rect 74 363 75 364
rect 73 363 74 364
rect 72 363 73 364
rect 71 363 72 364
rect 70 363 71 364
rect 69 363 70 364
rect 68 363 69 364
rect 67 363 68 364
rect 66 363 67 364
rect 65 363 66 364
rect 64 363 65 364
rect 63 363 64 364
rect 62 363 63 364
rect 61 363 62 364
rect 60 363 61 364
rect 59 363 60 364
rect 58 363 59 364
rect 57 363 58 364
rect 56 363 57 364
rect 55 363 56 364
rect 54 363 55 364
rect 53 363 54 364
rect 52 363 53 364
rect 51 363 52 364
rect 50 363 51 364
rect 49 363 50 364
rect 48 363 49 364
rect 47 363 48 364
rect 46 363 47 364
rect 45 363 46 364
rect 44 363 45 364
rect 43 363 44 364
rect 42 363 43 364
rect 41 363 42 364
rect 40 363 41 364
rect 39 363 40 364
rect 38 363 39 364
rect 37 363 38 364
rect 36 363 37 364
rect 35 363 36 364
rect 34 363 35 364
rect 33 363 34 364
rect 32 363 33 364
rect 31 363 32 364
rect 30 363 31 364
rect 29 363 30 364
rect 28 363 29 364
rect 27 363 28 364
rect 26 363 27 364
rect 25 363 26 364
rect 24 363 25 364
rect 23 363 24 364
rect 22 363 23 364
rect 21 363 22 364
rect 20 363 21 364
rect 19 363 20 364
rect 18 363 19 364
rect 144 364 145 365
rect 143 364 144 365
rect 142 364 143 365
rect 141 364 142 365
rect 140 364 141 365
rect 139 364 140 365
rect 138 364 139 365
rect 137 364 138 365
rect 136 364 137 365
rect 135 364 136 365
rect 134 364 135 365
rect 133 364 134 365
rect 132 364 133 365
rect 131 364 132 365
rect 130 364 131 365
rect 129 364 130 365
rect 128 364 129 365
rect 127 364 128 365
rect 126 364 127 365
rect 125 364 126 365
rect 124 364 125 365
rect 123 364 124 365
rect 122 364 123 365
rect 121 364 122 365
rect 120 364 121 365
rect 119 364 120 365
rect 81 364 82 365
rect 80 364 81 365
rect 79 364 80 365
rect 78 364 79 365
rect 77 364 78 365
rect 76 364 77 365
rect 75 364 76 365
rect 74 364 75 365
rect 73 364 74 365
rect 72 364 73 365
rect 71 364 72 365
rect 70 364 71 365
rect 69 364 70 365
rect 68 364 69 365
rect 67 364 68 365
rect 66 364 67 365
rect 65 364 66 365
rect 64 364 65 365
rect 63 364 64 365
rect 62 364 63 365
rect 61 364 62 365
rect 60 364 61 365
rect 59 364 60 365
rect 58 364 59 365
rect 57 364 58 365
rect 56 364 57 365
rect 55 364 56 365
rect 54 364 55 365
rect 53 364 54 365
rect 52 364 53 365
rect 51 364 52 365
rect 50 364 51 365
rect 49 364 50 365
rect 48 364 49 365
rect 47 364 48 365
rect 46 364 47 365
rect 45 364 46 365
rect 44 364 45 365
rect 43 364 44 365
rect 42 364 43 365
rect 41 364 42 365
rect 40 364 41 365
rect 39 364 40 365
rect 38 364 39 365
rect 37 364 38 365
rect 36 364 37 365
rect 35 364 36 365
rect 34 364 35 365
rect 33 364 34 365
rect 32 364 33 365
rect 31 364 32 365
rect 30 364 31 365
rect 29 364 30 365
rect 28 364 29 365
rect 27 364 28 365
rect 26 364 27 365
rect 25 364 26 365
rect 24 364 25 365
rect 23 364 24 365
rect 22 364 23 365
rect 21 364 22 365
rect 20 364 21 365
rect 19 364 20 365
rect 18 364 19 365
rect 144 365 145 366
rect 143 365 144 366
rect 142 365 143 366
rect 141 365 142 366
rect 140 365 141 366
rect 139 365 140 366
rect 138 365 139 366
rect 137 365 138 366
rect 136 365 137 366
rect 135 365 136 366
rect 134 365 135 366
rect 133 365 134 366
rect 132 365 133 366
rect 131 365 132 366
rect 130 365 131 366
rect 129 365 130 366
rect 128 365 129 366
rect 127 365 128 366
rect 126 365 127 366
rect 125 365 126 366
rect 124 365 125 366
rect 123 365 124 366
rect 122 365 123 366
rect 121 365 122 366
rect 120 365 121 366
rect 119 365 120 366
rect 81 365 82 366
rect 80 365 81 366
rect 79 365 80 366
rect 78 365 79 366
rect 77 365 78 366
rect 76 365 77 366
rect 75 365 76 366
rect 74 365 75 366
rect 73 365 74 366
rect 72 365 73 366
rect 71 365 72 366
rect 70 365 71 366
rect 69 365 70 366
rect 68 365 69 366
rect 67 365 68 366
rect 66 365 67 366
rect 65 365 66 366
rect 64 365 65 366
rect 63 365 64 366
rect 62 365 63 366
rect 61 365 62 366
rect 60 365 61 366
rect 59 365 60 366
rect 58 365 59 366
rect 57 365 58 366
rect 56 365 57 366
rect 55 365 56 366
rect 54 365 55 366
rect 53 365 54 366
rect 52 365 53 366
rect 51 365 52 366
rect 50 365 51 366
rect 49 365 50 366
rect 48 365 49 366
rect 47 365 48 366
rect 46 365 47 366
rect 45 365 46 366
rect 44 365 45 366
rect 43 365 44 366
rect 42 365 43 366
rect 41 365 42 366
rect 40 365 41 366
rect 39 365 40 366
rect 38 365 39 366
rect 37 365 38 366
rect 36 365 37 366
rect 35 365 36 366
rect 34 365 35 366
rect 33 365 34 366
rect 32 365 33 366
rect 31 365 32 366
rect 30 365 31 366
rect 29 365 30 366
rect 28 365 29 366
rect 27 365 28 366
rect 26 365 27 366
rect 25 365 26 366
rect 24 365 25 366
rect 23 365 24 366
rect 22 365 23 366
rect 21 365 22 366
rect 20 365 21 366
rect 19 365 20 366
rect 18 365 19 366
rect 17 365 18 366
rect 132 366 133 367
rect 131 366 132 367
rect 130 366 131 367
rect 82 366 83 367
rect 81 366 82 367
rect 80 366 81 367
rect 79 366 80 367
rect 78 366 79 367
rect 77 366 78 367
rect 76 366 77 367
rect 75 366 76 367
rect 74 366 75 367
rect 73 366 74 367
rect 72 366 73 367
rect 71 366 72 367
rect 70 366 71 367
rect 69 366 70 367
rect 68 366 69 367
rect 67 366 68 367
rect 66 366 67 367
rect 65 366 66 367
rect 64 366 65 367
rect 63 366 64 367
rect 62 366 63 367
rect 61 366 62 367
rect 60 366 61 367
rect 59 366 60 367
rect 58 366 59 367
rect 57 366 58 367
rect 56 366 57 367
rect 55 366 56 367
rect 54 366 55 367
rect 53 366 54 367
rect 52 366 53 367
rect 51 366 52 367
rect 50 366 51 367
rect 49 366 50 367
rect 48 366 49 367
rect 47 366 48 367
rect 46 366 47 367
rect 45 366 46 367
rect 44 366 45 367
rect 43 366 44 367
rect 42 366 43 367
rect 41 366 42 367
rect 40 366 41 367
rect 39 366 40 367
rect 38 366 39 367
rect 37 366 38 367
rect 36 366 37 367
rect 35 366 36 367
rect 34 366 35 367
rect 33 366 34 367
rect 32 366 33 367
rect 31 366 32 367
rect 30 366 31 367
rect 29 366 30 367
rect 28 366 29 367
rect 27 366 28 367
rect 26 366 27 367
rect 25 366 26 367
rect 24 366 25 367
rect 23 366 24 367
rect 22 366 23 367
rect 21 366 22 367
rect 20 366 21 367
rect 19 366 20 367
rect 18 366 19 367
rect 17 366 18 367
rect 133 367 134 368
rect 132 367 133 368
rect 131 367 132 368
rect 130 367 131 368
rect 82 367 83 368
rect 81 367 82 368
rect 80 367 81 368
rect 79 367 80 368
rect 78 367 79 368
rect 77 367 78 368
rect 76 367 77 368
rect 75 367 76 368
rect 74 367 75 368
rect 73 367 74 368
rect 72 367 73 368
rect 71 367 72 368
rect 70 367 71 368
rect 69 367 70 368
rect 68 367 69 368
rect 67 367 68 368
rect 66 367 67 368
rect 65 367 66 368
rect 64 367 65 368
rect 63 367 64 368
rect 62 367 63 368
rect 61 367 62 368
rect 60 367 61 368
rect 59 367 60 368
rect 58 367 59 368
rect 57 367 58 368
rect 56 367 57 368
rect 55 367 56 368
rect 54 367 55 368
rect 53 367 54 368
rect 52 367 53 368
rect 51 367 52 368
rect 50 367 51 368
rect 49 367 50 368
rect 48 367 49 368
rect 47 367 48 368
rect 46 367 47 368
rect 45 367 46 368
rect 44 367 45 368
rect 43 367 44 368
rect 42 367 43 368
rect 41 367 42 368
rect 40 367 41 368
rect 39 367 40 368
rect 38 367 39 368
rect 37 367 38 368
rect 36 367 37 368
rect 35 367 36 368
rect 34 367 35 368
rect 33 367 34 368
rect 32 367 33 368
rect 31 367 32 368
rect 30 367 31 368
rect 29 367 30 368
rect 28 367 29 368
rect 27 367 28 368
rect 26 367 27 368
rect 25 367 26 368
rect 24 367 25 368
rect 23 367 24 368
rect 22 367 23 368
rect 21 367 22 368
rect 20 367 21 368
rect 19 367 20 368
rect 18 367 19 368
rect 17 367 18 368
rect 134 368 135 369
rect 133 368 134 369
rect 132 368 133 369
rect 131 368 132 369
rect 130 368 131 369
rect 129 368 130 369
rect 128 368 129 369
rect 82 368 83 369
rect 81 368 82 369
rect 80 368 81 369
rect 79 368 80 369
rect 78 368 79 369
rect 77 368 78 369
rect 76 368 77 369
rect 75 368 76 369
rect 74 368 75 369
rect 73 368 74 369
rect 72 368 73 369
rect 71 368 72 369
rect 70 368 71 369
rect 69 368 70 369
rect 68 368 69 369
rect 67 368 68 369
rect 66 368 67 369
rect 65 368 66 369
rect 64 368 65 369
rect 63 368 64 369
rect 62 368 63 369
rect 61 368 62 369
rect 60 368 61 369
rect 59 368 60 369
rect 58 368 59 369
rect 57 368 58 369
rect 56 368 57 369
rect 55 368 56 369
rect 54 368 55 369
rect 53 368 54 369
rect 52 368 53 369
rect 51 368 52 369
rect 50 368 51 369
rect 49 368 50 369
rect 48 368 49 369
rect 47 368 48 369
rect 46 368 47 369
rect 45 368 46 369
rect 44 368 45 369
rect 43 368 44 369
rect 42 368 43 369
rect 41 368 42 369
rect 40 368 41 369
rect 39 368 40 369
rect 38 368 39 369
rect 37 368 38 369
rect 36 368 37 369
rect 35 368 36 369
rect 34 368 35 369
rect 33 368 34 369
rect 32 368 33 369
rect 31 368 32 369
rect 30 368 31 369
rect 29 368 30 369
rect 28 368 29 369
rect 27 368 28 369
rect 26 368 27 369
rect 25 368 26 369
rect 24 368 25 369
rect 23 368 24 369
rect 22 368 23 369
rect 21 368 22 369
rect 20 368 21 369
rect 19 368 20 369
rect 18 368 19 369
rect 17 368 18 369
rect 16 368 17 369
rect 136 369 137 370
rect 135 369 136 370
rect 134 369 135 370
rect 133 369 134 370
rect 132 369 133 370
rect 131 369 132 370
rect 130 369 131 370
rect 129 369 130 370
rect 128 369 129 370
rect 127 369 128 370
rect 82 369 83 370
rect 81 369 82 370
rect 80 369 81 370
rect 79 369 80 370
rect 78 369 79 370
rect 77 369 78 370
rect 76 369 77 370
rect 75 369 76 370
rect 74 369 75 370
rect 73 369 74 370
rect 72 369 73 370
rect 71 369 72 370
rect 70 369 71 370
rect 69 369 70 370
rect 68 369 69 370
rect 67 369 68 370
rect 66 369 67 370
rect 65 369 66 370
rect 64 369 65 370
rect 63 369 64 370
rect 62 369 63 370
rect 61 369 62 370
rect 60 369 61 370
rect 59 369 60 370
rect 58 369 59 370
rect 57 369 58 370
rect 56 369 57 370
rect 55 369 56 370
rect 54 369 55 370
rect 53 369 54 370
rect 52 369 53 370
rect 51 369 52 370
rect 50 369 51 370
rect 49 369 50 370
rect 48 369 49 370
rect 47 369 48 370
rect 46 369 47 370
rect 45 369 46 370
rect 44 369 45 370
rect 43 369 44 370
rect 42 369 43 370
rect 41 369 42 370
rect 40 369 41 370
rect 39 369 40 370
rect 38 369 39 370
rect 37 369 38 370
rect 36 369 37 370
rect 35 369 36 370
rect 34 369 35 370
rect 33 369 34 370
rect 32 369 33 370
rect 31 369 32 370
rect 30 369 31 370
rect 29 369 30 370
rect 28 369 29 370
rect 27 369 28 370
rect 26 369 27 370
rect 25 369 26 370
rect 24 369 25 370
rect 23 369 24 370
rect 22 369 23 370
rect 21 369 22 370
rect 20 369 21 370
rect 19 369 20 370
rect 18 369 19 370
rect 17 369 18 370
rect 16 369 17 370
rect 137 370 138 371
rect 136 370 137 371
rect 135 370 136 371
rect 134 370 135 371
rect 133 370 134 371
rect 132 370 133 371
rect 131 370 132 371
rect 130 370 131 371
rect 129 370 130 371
rect 128 370 129 371
rect 127 370 128 371
rect 126 370 127 371
rect 125 370 126 371
rect 83 370 84 371
rect 82 370 83 371
rect 81 370 82 371
rect 80 370 81 371
rect 79 370 80 371
rect 78 370 79 371
rect 77 370 78 371
rect 76 370 77 371
rect 75 370 76 371
rect 74 370 75 371
rect 73 370 74 371
rect 72 370 73 371
rect 71 370 72 371
rect 70 370 71 371
rect 69 370 70 371
rect 68 370 69 371
rect 67 370 68 371
rect 66 370 67 371
rect 65 370 66 371
rect 64 370 65 371
rect 63 370 64 371
rect 62 370 63 371
rect 61 370 62 371
rect 60 370 61 371
rect 39 370 40 371
rect 38 370 39 371
rect 37 370 38 371
rect 36 370 37 371
rect 35 370 36 371
rect 34 370 35 371
rect 33 370 34 371
rect 32 370 33 371
rect 31 370 32 371
rect 30 370 31 371
rect 29 370 30 371
rect 28 370 29 371
rect 27 370 28 371
rect 26 370 27 371
rect 25 370 26 371
rect 24 370 25 371
rect 23 370 24 371
rect 22 370 23 371
rect 21 370 22 371
rect 20 370 21 371
rect 19 370 20 371
rect 18 370 19 371
rect 17 370 18 371
rect 16 370 17 371
rect 139 371 140 372
rect 138 371 139 372
rect 137 371 138 372
rect 136 371 137 372
rect 135 371 136 372
rect 134 371 135 372
rect 133 371 134 372
rect 132 371 133 372
rect 131 371 132 372
rect 130 371 131 372
rect 129 371 130 372
rect 128 371 129 372
rect 127 371 128 372
rect 126 371 127 372
rect 125 371 126 372
rect 124 371 125 372
rect 83 371 84 372
rect 82 371 83 372
rect 81 371 82 372
rect 80 371 81 372
rect 79 371 80 372
rect 78 371 79 372
rect 77 371 78 372
rect 76 371 77 372
rect 75 371 76 372
rect 74 371 75 372
rect 73 371 74 372
rect 72 371 73 372
rect 71 371 72 372
rect 70 371 71 372
rect 69 371 70 372
rect 68 371 69 372
rect 67 371 68 372
rect 66 371 67 372
rect 65 371 66 372
rect 34 371 35 372
rect 33 371 34 372
rect 32 371 33 372
rect 31 371 32 372
rect 30 371 31 372
rect 29 371 30 372
rect 28 371 29 372
rect 27 371 28 372
rect 26 371 27 372
rect 25 371 26 372
rect 24 371 25 372
rect 23 371 24 372
rect 22 371 23 372
rect 21 371 22 372
rect 20 371 21 372
rect 19 371 20 372
rect 18 371 19 372
rect 17 371 18 372
rect 16 371 17 372
rect 140 372 141 373
rect 139 372 140 373
rect 138 372 139 373
rect 137 372 138 373
rect 136 372 137 373
rect 135 372 136 373
rect 134 372 135 373
rect 133 372 134 373
rect 132 372 133 373
rect 131 372 132 373
rect 130 372 131 373
rect 129 372 130 373
rect 128 372 129 373
rect 127 372 128 373
rect 126 372 127 373
rect 125 372 126 373
rect 124 372 125 373
rect 123 372 124 373
rect 122 372 123 373
rect 83 372 84 373
rect 82 372 83 373
rect 81 372 82 373
rect 80 372 81 373
rect 79 372 80 373
rect 78 372 79 373
rect 77 372 78 373
rect 76 372 77 373
rect 75 372 76 373
rect 74 372 75 373
rect 73 372 74 373
rect 72 372 73 373
rect 71 372 72 373
rect 70 372 71 373
rect 69 372 70 373
rect 68 372 69 373
rect 67 372 68 373
rect 31 372 32 373
rect 30 372 31 373
rect 29 372 30 373
rect 28 372 29 373
rect 27 372 28 373
rect 26 372 27 373
rect 25 372 26 373
rect 24 372 25 373
rect 23 372 24 373
rect 22 372 23 373
rect 21 372 22 373
rect 20 372 21 373
rect 19 372 20 373
rect 18 372 19 373
rect 17 372 18 373
rect 16 372 17 373
rect 15 372 16 373
rect 142 373 143 374
rect 141 373 142 374
rect 140 373 141 374
rect 139 373 140 374
rect 138 373 139 374
rect 137 373 138 374
rect 136 373 137 374
rect 135 373 136 374
rect 134 373 135 374
rect 133 373 134 374
rect 129 373 130 374
rect 128 373 129 374
rect 127 373 128 374
rect 126 373 127 374
rect 125 373 126 374
rect 124 373 125 374
rect 123 373 124 374
rect 122 373 123 374
rect 121 373 122 374
rect 83 373 84 374
rect 82 373 83 374
rect 81 373 82 374
rect 80 373 81 374
rect 79 373 80 374
rect 78 373 79 374
rect 77 373 78 374
rect 76 373 77 374
rect 75 373 76 374
rect 74 373 75 374
rect 73 373 74 374
rect 72 373 73 374
rect 71 373 72 374
rect 70 373 71 374
rect 69 373 70 374
rect 68 373 69 374
rect 30 373 31 374
rect 29 373 30 374
rect 28 373 29 374
rect 27 373 28 374
rect 26 373 27 374
rect 25 373 26 374
rect 24 373 25 374
rect 23 373 24 374
rect 22 373 23 374
rect 21 373 22 374
rect 20 373 21 374
rect 19 373 20 374
rect 18 373 19 374
rect 17 373 18 374
rect 16 373 17 374
rect 15 373 16 374
rect 143 374 144 375
rect 142 374 143 375
rect 141 374 142 375
rect 140 374 141 375
rect 139 374 140 375
rect 138 374 139 375
rect 137 374 138 375
rect 136 374 137 375
rect 135 374 136 375
rect 134 374 135 375
rect 128 374 129 375
rect 127 374 128 375
rect 126 374 127 375
rect 125 374 126 375
rect 124 374 125 375
rect 123 374 124 375
rect 122 374 123 375
rect 121 374 122 375
rect 120 374 121 375
rect 119 374 120 375
rect 83 374 84 375
rect 82 374 83 375
rect 81 374 82 375
rect 80 374 81 375
rect 79 374 80 375
rect 78 374 79 375
rect 77 374 78 375
rect 76 374 77 375
rect 75 374 76 375
rect 74 374 75 375
rect 73 374 74 375
rect 72 374 73 375
rect 71 374 72 375
rect 70 374 71 375
rect 69 374 70 375
rect 29 374 30 375
rect 28 374 29 375
rect 27 374 28 375
rect 26 374 27 375
rect 25 374 26 375
rect 24 374 25 375
rect 23 374 24 375
rect 22 374 23 375
rect 21 374 22 375
rect 20 374 21 375
rect 19 374 20 375
rect 18 374 19 375
rect 17 374 18 375
rect 16 374 17 375
rect 15 374 16 375
rect 144 375 145 376
rect 143 375 144 376
rect 142 375 143 376
rect 141 375 142 376
rect 140 375 141 376
rect 139 375 140 376
rect 138 375 139 376
rect 137 375 138 376
rect 136 375 137 376
rect 126 375 127 376
rect 125 375 126 376
rect 124 375 125 376
rect 123 375 124 376
rect 122 375 123 376
rect 121 375 122 376
rect 120 375 121 376
rect 119 375 120 376
rect 83 375 84 376
rect 82 375 83 376
rect 81 375 82 376
rect 80 375 81 376
rect 79 375 80 376
rect 78 375 79 376
rect 77 375 78 376
rect 76 375 77 376
rect 75 375 76 376
rect 74 375 75 376
rect 73 375 74 376
rect 72 375 73 376
rect 71 375 72 376
rect 70 375 71 376
rect 69 375 70 376
rect 29 375 30 376
rect 28 375 29 376
rect 27 375 28 376
rect 26 375 27 376
rect 25 375 26 376
rect 24 375 25 376
rect 23 375 24 376
rect 22 375 23 376
rect 21 375 22 376
rect 20 375 21 376
rect 19 375 20 376
rect 18 375 19 376
rect 17 375 18 376
rect 16 375 17 376
rect 15 375 16 376
rect 144 376 145 377
rect 143 376 144 377
rect 142 376 143 377
rect 141 376 142 377
rect 140 376 141 377
rect 139 376 140 377
rect 138 376 139 377
rect 137 376 138 377
rect 125 376 126 377
rect 124 376 125 377
rect 123 376 124 377
rect 122 376 123 377
rect 121 376 122 377
rect 120 376 121 377
rect 119 376 120 377
rect 83 376 84 377
rect 82 376 83 377
rect 81 376 82 377
rect 80 376 81 377
rect 79 376 80 377
rect 78 376 79 377
rect 77 376 78 377
rect 76 376 77 377
rect 75 376 76 377
rect 74 376 75 377
rect 73 376 74 377
rect 72 376 73 377
rect 71 376 72 377
rect 70 376 71 377
rect 69 376 70 377
rect 29 376 30 377
rect 28 376 29 377
rect 27 376 28 377
rect 26 376 27 377
rect 25 376 26 377
rect 24 376 25 377
rect 23 376 24 377
rect 22 376 23 377
rect 21 376 22 377
rect 20 376 21 377
rect 19 376 20 377
rect 18 376 19 377
rect 17 376 18 377
rect 16 376 17 377
rect 15 376 16 377
rect 144 377 145 378
rect 143 377 144 378
rect 142 377 143 378
rect 141 377 142 378
rect 140 377 141 378
rect 139 377 140 378
rect 138 377 139 378
rect 123 377 124 378
rect 122 377 123 378
rect 121 377 122 378
rect 120 377 121 378
rect 119 377 120 378
rect 83 377 84 378
rect 82 377 83 378
rect 81 377 82 378
rect 80 377 81 378
rect 79 377 80 378
rect 78 377 79 378
rect 77 377 78 378
rect 76 377 77 378
rect 75 377 76 378
rect 74 377 75 378
rect 73 377 74 378
rect 72 377 73 378
rect 71 377 72 378
rect 70 377 71 378
rect 69 377 70 378
rect 29 377 30 378
rect 28 377 29 378
rect 27 377 28 378
rect 26 377 27 378
rect 25 377 26 378
rect 24 377 25 378
rect 23 377 24 378
rect 22 377 23 378
rect 21 377 22 378
rect 20 377 21 378
rect 19 377 20 378
rect 18 377 19 378
rect 17 377 18 378
rect 16 377 17 378
rect 15 377 16 378
rect 144 378 145 379
rect 143 378 144 379
rect 142 378 143 379
rect 141 378 142 379
rect 140 378 141 379
rect 122 378 123 379
rect 121 378 122 379
rect 120 378 121 379
rect 119 378 120 379
rect 83 378 84 379
rect 82 378 83 379
rect 81 378 82 379
rect 80 378 81 379
rect 79 378 80 379
rect 78 378 79 379
rect 77 378 78 379
rect 76 378 77 379
rect 75 378 76 379
rect 74 378 75 379
rect 73 378 74 379
rect 72 378 73 379
rect 71 378 72 379
rect 70 378 71 379
rect 69 378 70 379
rect 68 378 69 379
rect 30 378 31 379
rect 29 378 30 379
rect 28 378 29 379
rect 27 378 28 379
rect 26 378 27 379
rect 25 378 26 379
rect 24 378 25 379
rect 23 378 24 379
rect 22 378 23 379
rect 21 378 22 379
rect 20 378 21 379
rect 19 378 20 379
rect 18 378 19 379
rect 17 378 18 379
rect 16 378 17 379
rect 15 378 16 379
rect 144 379 145 380
rect 143 379 144 380
rect 142 379 143 380
rect 141 379 142 380
rect 121 379 122 380
rect 120 379 121 380
rect 119 379 120 380
rect 83 379 84 380
rect 82 379 83 380
rect 81 379 82 380
rect 80 379 81 380
rect 79 379 80 380
rect 78 379 79 380
rect 77 379 78 380
rect 76 379 77 380
rect 75 379 76 380
rect 74 379 75 380
rect 73 379 74 380
rect 72 379 73 380
rect 71 379 72 380
rect 70 379 71 380
rect 69 379 70 380
rect 68 379 69 380
rect 67 379 68 380
rect 31 379 32 380
rect 30 379 31 380
rect 29 379 30 380
rect 28 379 29 380
rect 27 379 28 380
rect 26 379 27 380
rect 25 379 26 380
rect 24 379 25 380
rect 23 379 24 380
rect 22 379 23 380
rect 21 379 22 380
rect 20 379 21 380
rect 19 379 20 380
rect 18 379 19 380
rect 17 379 18 380
rect 16 379 17 380
rect 15 379 16 380
rect 144 380 145 381
rect 143 380 144 381
rect 119 380 120 381
rect 83 380 84 381
rect 82 380 83 381
rect 81 380 82 381
rect 80 380 81 381
rect 79 380 80 381
rect 78 380 79 381
rect 77 380 78 381
rect 76 380 77 381
rect 75 380 76 381
rect 74 380 75 381
rect 73 380 74 381
rect 72 380 73 381
rect 71 380 72 381
rect 70 380 71 381
rect 69 380 70 381
rect 68 380 69 381
rect 67 380 68 381
rect 66 380 67 381
rect 65 380 66 381
rect 64 380 65 381
rect 33 380 34 381
rect 32 380 33 381
rect 31 380 32 381
rect 30 380 31 381
rect 29 380 30 381
rect 28 380 29 381
rect 27 380 28 381
rect 26 380 27 381
rect 25 380 26 381
rect 24 380 25 381
rect 23 380 24 381
rect 22 380 23 381
rect 21 380 22 381
rect 20 380 21 381
rect 19 380 20 381
rect 18 380 19 381
rect 17 380 18 381
rect 16 380 17 381
rect 15 380 16 381
rect 144 381 145 382
rect 82 381 83 382
rect 81 381 82 382
rect 80 381 81 382
rect 79 381 80 382
rect 78 381 79 382
rect 77 381 78 382
rect 76 381 77 382
rect 75 381 76 382
rect 74 381 75 382
rect 73 381 74 382
rect 72 381 73 382
rect 71 381 72 382
rect 70 381 71 382
rect 69 381 70 382
rect 68 381 69 382
rect 67 381 68 382
rect 66 381 67 382
rect 65 381 66 382
rect 64 381 65 382
rect 63 381 64 382
rect 62 381 63 382
rect 61 381 62 382
rect 60 381 61 382
rect 37 381 38 382
rect 36 381 37 382
rect 35 381 36 382
rect 34 381 35 382
rect 33 381 34 382
rect 32 381 33 382
rect 31 381 32 382
rect 30 381 31 382
rect 29 381 30 382
rect 28 381 29 382
rect 27 381 28 382
rect 26 381 27 382
rect 25 381 26 382
rect 24 381 25 382
rect 23 381 24 382
rect 22 381 23 382
rect 21 381 22 382
rect 20 381 21 382
rect 19 381 20 382
rect 18 381 19 382
rect 17 381 18 382
rect 16 381 17 382
rect 15 381 16 382
rect 82 382 83 383
rect 81 382 82 383
rect 80 382 81 383
rect 79 382 80 383
rect 78 382 79 383
rect 77 382 78 383
rect 76 382 77 383
rect 75 382 76 383
rect 74 382 75 383
rect 73 382 74 383
rect 72 382 73 383
rect 71 382 72 383
rect 70 382 71 383
rect 69 382 70 383
rect 68 382 69 383
rect 67 382 68 383
rect 66 382 67 383
rect 65 382 66 383
rect 64 382 65 383
rect 63 382 64 383
rect 62 382 63 383
rect 61 382 62 383
rect 60 382 61 383
rect 59 382 60 383
rect 58 382 59 383
rect 57 382 58 383
rect 56 382 57 383
rect 55 382 56 383
rect 54 382 55 383
rect 53 382 54 383
rect 52 382 53 383
rect 51 382 52 383
rect 50 382 51 383
rect 49 382 50 383
rect 48 382 49 383
rect 47 382 48 383
rect 46 382 47 383
rect 45 382 46 383
rect 44 382 45 383
rect 43 382 44 383
rect 42 382 43 383
rect 41 382 42 383
rect 40 382 41 383
rect 39 382 40 383
rect 38 382 39 383
rect 37 382 38 383
rect 36 382 37 383
rect 35 382 36 383
rect 34 382 35 383
rect 33 382 34 383
rect 32 382 33 383
rect 31 382 32 383
rect 30 382 31 383
rect 29 382 30 383
rect 28 382 29 383
rect 27 382 28 383
rect 26 382 27 383
rect 25 382 26 383
rect 24 382 25 383
rect 23 382 24 383
rect 22 382 23 383
rect 21 382 22 383
rect 20 382 21 383
rect 19 382 20 383
rect 18 382 19 383
rect 17 382 18 383
rect 16 382 17 383
rect 136 383 137 384
rect 135 383 136 384
rect 134 383 135 384
rect 82 383 83 384
rect 81 383 82 384
rect 80 383 81 384
rect 79 383 80 384
rect 78 383 79 384
rect 77 383 78 384
rect 76 383 77 384
rect 75 383 76 384
rect 74 383 75 384
rect 73 383 74 384
rect 72 383 73 384
rect 71 383 72 384
rect 70 383 71 384
rect 69 383 70 384
rect 68 383 69 384
rect 67 383 68 384
rect 66 383 67 384
rect 65 383 66 384
rect 64 383 65 384
rect 63 383 64 384
rect 62 383 63 384
rect 61 383 62 384
rect 60 383 61 384
rect 59 383 60 384
rect 58 383 59 384
rect 57 383 58 384
rect 56 383 57 384
rect 55 383 56 384
rect 54 383 55 384
rect 53 383 54 384
rect 52 383 53 384
rect 51 383 52 384
rect 50 383 51 384
rect 49 383 50 384
rect 48 383 49 384
rect 47 383 48 384
rect 46 383 47 384
rect 45 383 46 384
rect 44 383 45 384
rect 43 383 44 384
rect 42 383 43 384
rect 41 383 42 384
rect 40 383 41 384
rect 39 383 40 384
rect 38 383 39 384
rect 37 383 38 384
rect 36 383 37 384
rect 35 383 36 384
rect 34 383 35 384
rect 33 383 34 384
rect 32 383 33 384
rect 31 383 32 384
rect 30 383 31 384
rect 29 383 30 384
rect 28 383 29 384
rect 27 383 28 384
rect 26 383 27 384
rect 25 383 26 384
rect 24 383 25 384
rect 23 383 24 384
rect 22 383 23 384
rect 21 383 22 384
rect 20 383 21 384
rect 19 383 20 384
rect 18 383 19 384
rect 17 383 18 384
rect 16 383 17 384
rect 139 384 140 385
rect 138 384 139 385
rect 137 384 138 385
rect 136 384 137 385
rect 135 384 136 385
rect 134 384 135 385
rect 133 384 134 385
rect 132 384 133 385
rect 131 384 132 385
rect 82 384 83 385
rect 81 384 82 385
rect 80 384 81 385
rect 79 384 80 385
rect 78 384 79 385
rect 77 384 78 385
rect 76 384 77 385
rect 75 384 76 385
rect 74 384 75 385
rect 73 384 74 385
rect 72 384 73 385
rect 71 384 72 385
rect 70 384 71 385
rect 69 384 70 385
rect 68 384 69 385
rect 67 384 68 385
rect 66 384 67 385
rect 65 384 66 385
rect 64 384 65 385
rect 63 384 64 385
rect 62 384 63 385
rect 61 384 62 385
rect 60 384 61 385
rect 59 384 60 385
rect 58 384 59 385
rect 57 384 58 385
rect 56 384 57 385
rect 55 384 56 385
rect 54 384 55 385
rect 53 384 54 385
rect 52 384 53 385
rect 51 384 52 385
rect 50 384 51 385
rect 49 384 50 385
rect 48 384 49 385
rect 47 384 48 385
rect 46 384 47 385
rect 45 384 46 385
rect 44 384 45 385
rect 43 384 44 385
rect 42 384 43 385
rect 41 384 42 385
rect 40 384 41 385
rect 39 384 40 385
rect 38 384 39 385
rect 37 384 38 385
rect 36 384 37 385
rect 35 384 36 385
rect 34 384 35 385
rect 33 384 34 385
rect 32 384 33 385
rect 31 384 32 385
rect 30 384 31 385
rect 29 384 30 385
rect 28 384 29 385
rect 27 384 28 385
rect 26 384 27 385
rect 25 384 26 385
rect 24 384 25 385
rect 23 384 24 385
rect 22 384 23 385
rect 21 384 22 385
rect 20 384 21 385
rect 19 384 20 385
rect 18 384 19 385
rect 17 384 18 385
rect 16 384 17 385
rect 141 385 142 386
rect 140 385 141 386
rect 139 385 140 386
rect 138 385 139 386
rect 137 385 138 386
rect 136 385 137 386
rect 135 385 136 386
rect 134 385 135 386
rect 133 385 134 386
rect 132 385 133 386
rect 131 385 132 386
rect 130 385 131 386
rect 129 385 130 386
rect 81 385 82 386
rect 80 385 81 386
rect 79 385 80 386
rect 78 385 79 386
rect 77 385 78 386
rect 76 385 77 386
rect 75 385 76 386
rect 74 385 75 386
rect 73 385 74 386
rect 72 385 73 386
rect 71 385 72 386
rect 70 385 71 386
rect 69 385 70 386
rect 68 385 69 386
rect 67 385 68 386
rect 66 385 67 386
rect 65 385 66 386
rect 64 385 65 386
rect 63 385 64 386
rect 62 385 63 386
rect 61 385 62 386
rect 60 385 61 386
rect 59 385 60 386
rect 58 385 59 386
rect 57 385 58 386
rect 56 385 57 386
rect 55 385 56 386
rect 54 385 55 386
rect 53 385 54 386
rect 52 385 53 386
rect 51 385 52 386
rect 50 385 51 386
rect 49 385 50 386
rect 48 385 49 386
rect 47 385 48 386
rect 46 385 47 386
rect 45 385 46 386
rect 44 385 45 386
rect 43 385 44 386
rect 42 385 43 386
rect 41 385 42 386
rect 40 385 41 386
rect 39 385 40 386
rect 38 385 39 386
rect 37 385 38 386
rect 36 385 37 386
rect 35 385 36 386
rect 34 385 35 386
rect 33 385 34 386
rect 32 385 33 386
rect 31 385 32 386
rect 30 385 31 386
rect 29 385 30 386
rect 28 385 29 386
rect 27 385 28 386
rect 26 385 27 386
rect 25 385 26 386
rect 24 385 25 386
rect 23 385 24 386
rect 22 385 23 386
rect 21 385 22 386
rect 20 385 21 386
rect 19 385 20 386
rect 18 385 19 386
rect 17 385 18 386
rect 16 385 17 386
rect 142 386 143 387
rect 141 386 142 387
rect 140 386 141 387
rect 139 386 140 387
rect 138 386 139 387
rect 137 386 138 387
rect 136 386 137 387
rect 135 386 136 387
rect 134 386 135 387
rect 133 386 134 387
rect 132 386 133 387
rect 131 386 132 387
rect 130 386 131 387
rect 129 386 130 387
rect 128 386 129 387
rect 81 386 82 387
rect 80 386 81 387
rect 79 386 80 387
rect 78 386 79 387
rect 77 386 78 387
rect 76 386 77 387
rect 75 386 76 387
rect 74 386 75 387
rect 73 386 74 387
rect 72 386 73 387
rect 71 386 72 387
rect 70 386 71 387
rect 69 386 70 387
rect 68 386 69 387
rect 67 386 68 387
rect 66 386 67 387
rect 65 386 66 387
rect 64 386 65 387
rect 63 386 64 387
rect 62 386 63 387
rect 61 386 62 387
rect 60 386 61 387
rect 59 386 60 387
rect 58 386 59 387
rect 57 386 58 387
rect 56 386 57 387
rect 55 386 56 387
rect 54 386 55 387
rect 53 386 54 387
rect 52 386 53 387
rect 51 386 52 387
rect 50 386 51 387
rect 49 386 50 387
rect 48 386 49 387
rect 47 386 48 387
rect 46 386 47 387
rect 45 386 46 387
rect 44 386 45 387
rect 43 386 44 387
rect 42 386 43 387
rect 41 386 42 387
rect 40 386 41 387
rect 39 386 40 387
rect 38 386 39 387
rect 37 386 38 387
rect 36 386 37 387
rect 35 386 36 387
rect 34 386 35 387
rect 33 386 34 387
rect 32 386 33 387
rect 31 386 32 387
rect 30 386 31 387
rect 29 386 30 387
rect 28 386 29 387
rect 27 386 28 387
rect 26 386 27 387
rect 25 386 26 387
rect 24 386 25 387
rect 23 386 24 387
rect 22 386 23 387
rect 21 386 22 387
rect 20 386 21 387
rect 19 386 20 387
rect 18 386 19 387
rect 17 386 18 387
rect 143 387 144 388
rect 142 387 143 388
rect 141 387 142 388
rect 140 387 141 388
rect 139 387 140 388
rect 138 387 139 388
rect 137 387 138 388
rect 136 387 137 388
rect 135 387 136 388
rect 134 387 135 388
rect 133 387 134 388
rect 132 387 133 388
rect 131 387 132 388
rect 130 387 131 388
rect 129 387 130 388
rect 128 387 129 388
rect 127 387 128 388
rect 81 387 82 388
rect 80 387 81 388
rect 79 387 80 388
rect 78 387 79 388
rect 77 387 78 388
rect 76 387 77 388
rect 75 387 76 388
rect 74 387 75 388
rect 73 387 74 388
rect 72 387 73 388
rect 71 387 72 388
rect 70 387 71 388
rect 69 387 70 388
rect 68 387 69 388
rect 67 387 68 388
rect 66 387 67 388
rect 65 387 66 388
rect 64 387 65 388
rect 63 387 64 388
rect 62 387 63 388
rect 61 387 62 388
rect 60 387 61 388
rect 59 387 60 388
rect 58 387 59 388
rect 57 387 58 388
rect 56 387 57 388
rect 55 387 56 388
rect 54 387 55 388
rect 53 387 54 388
rect 52 387 53 388
rect 51 387 52 388
rect 50 387 51 388
rect 49 387 50 388
rect 48 387 49 388
rect 47 387 48 388
rect 46 387 47 388
rect 45 387 46 388
rect 44 387 45 388
rect 43 387 44 388
rect 42 387 43 388
rect 41 387 42 388
rect 40 387 41 388
rect 39 387 40 388
rect 38 387 39 388
rect 37 387 38 388
rect 36 387 37 388
rect 35 387 36 388
rect 34 387 35 388
rect 33 387 34 388
rect 32 387 33 388
rect 31 387 32 388
rect 30 387 31 388
rect 29 387 30 388
rect 28 387 29 388
rect 27 387 28 388
rect 26 387 27 388
rect 25 387 26 388
rect 24 387 25 388
rect 23 387 24 388
rect 22 387 23 388
rect 21 387 22 388
rect 20 387 21 388
rect 19 387 20 388
rect 18 387 19 388
rect 17 387 18 388
rect 143 388 144 389
rect 142 388 143 389
rect 141 388 142 389
rect 140 388 141 389
rect 139 388 140 389
rect 138 388 139 389
rect 137 388 138 389
rect 136 388 137 389
rect 135 388 136 389
rect 134 388 135 389
rect 133 388 134 389
rect 132 388 133 389
rect 131 388 132 389
rect 130 388 131 389
rect 129 388 130 389
rect 128 388 129 389
rect 127 388 128 389
rect 80 388 81 389
rect 79 388 80 389
rect 78 388 79 389
rect 77 388 78 389
rect 76 388 77 389
rect 75 388 76 389
rect 74 388 75 389
rect 73 388 74 389
rect 72 388 73 389
rect 71 388 72 389
rect 70 388 71 389
rect 69 388 70 389
rect 68 388 69 389
rect 67 388 68 389
rect 66 388 67 389
rect 65 388 66 389
rect 64 388 65 389
rect 63 388 64 389
rect 62 388 63 389
rect 61 388 62 389
rect 60 388 61 389
rect 59 388 60 389
rect 58 388 59 389
rect 57 388 58 389
rect 56 388 57 389
rect 55 388 56 389
rect 54 388 55 389
rect 53 388 54 389
rect 52 388 53 389
rect 51 388 52 389
rect 50 388 51 389
rect 49 388 50 389
rect 48 388 49 389
rect 47 388 48 389
rect 46 388 47 389
rect 45 388 46 389
rect 44 388 45 389
rect 43 388 44 389
rect 42 388 43 389
rect 41 388 42 389
rect 40 388 41 389
rect 39 388 40 389
rect 38 388 39 389
rect 37 388 38 389
rect 36 388 37 389
rect 35 388 36 389
rect 34 388 35 389
rect 33 388 34 389
rect 32 388 33 389
rect 31 388 32 389
rect 30 388 31 389
rect 29 388 30 389
rect 28 388 29 389
rect 27 388 28 389
rect 26 388 27 389
rect 25 388 26 389
rect 24 388 25 389
rect 23 388 24 389
rect 22 388 23 389
rect 21 388 22 389
rect 20 388 21 389
rect 19 388 20 389
rect 18 388 19 389
rect 17 388 18 389
rect 143 389 144 390
rect 142 389 143 390
rect 141 389 142 390
rect 140 389 141 390
rect 139 389 140 390
rect 138 389 139 390
rect 132 389 133 390
rect 131 389 132 390
rect 130 389 131 390
rect 129 389 130 390
rect 128 389 129 390
rect 127 389 128 390
rect 79 389 80 390
rect 78 389 79 390
rect 77 389 78 390
rect 76 389 77 390
rect 75 389 76 390
rect 74 389 75 390
rect 73 389 74 390
rect 72 389 73 390
rect 71 389 72 390
rect 70 389 71 390
rect 69 389 70 390
rect 68 389 69 390
rect 67 389 68 390
rect 66 389 67 390
rect 65 389 66 390
rect 64 389 65 390
rect 63 389 64 390
rect 62 389 63 390
rect 61 389 62 390
rect 60 389 61 390
rect 59 389 60 390
rect 58 389 59 390
rect 57 389 58 390
rect 56 389 57 390
rect 55 389 56 390
rect 54 389 55 390
rect 53 389 54 390
rect 52 389 53 390
rect 51 389 52 390
rect 50 389 51 390
rect 49 389 50 390
rect 48 389 49 390
rect 47 389 48 390
rect 46 389 47 390
rect 45 389 46 390
rect 44 389 45 390
rect 43 389 44 390
rect 42 389 43 390
rect 41 389 42 390
rect 40 389 41 390
rect 39 389 40 390
rect 38 389 39 390
rect 37 389 38 390
rect 36 389 37 390
rect 35 389 36 390
rect 34 389 35 390
rect 33 389 34 390
rect 32 389 33 390
rect 31 389 32 390
rect 30 389 31 390
rect 29 389 30 390
rect 28 389 29 390
rect 27 389 28 390
rect 26 389 27 390
rect 25 389 26 390
rect 24 389 25 390
rect 23 389 24 390
rect 22 389 23 390
rect 21 389 22 390
rect 20 389 21 390
rect 19 389 20 390
rect 18 389 19 390
rect 144 390 145 391
rect 143 390 144 391
rect 142 390 143 391
rect 141 390 142 391
rect 140 390 141 391
rect 130 390 131 391
rect 129 390 130 391
rect 128 390 129 391
rect 127 390 128 391
rect 126 390 127 391
rect 79 390 80 391
rect 78 390 79 391
rect 77 390 78 391
rect 76 390 77 391
rect 75 390 76 391
rect 74 390 75 391
rect 73 390 74 391
rect 72 390 73 391
rect 71 390 72 391
rect 70 390 71 391
rect 69 390 70 391
rect 68 390 69 391
rect 67 390 68 391
rect 66 390 67 391
rect 65 390 66 391
rect 64 390 65 391
rect 63 390 64 391
rect 62 390 63 391
rect 61 390 62 391
rect 60 390 61 391
rect 59 390 60 391
rect 58 390 59 391
rect 57 390 58 391
rect 56 390 57 391
rect 55 390 56 391
rect 54 390 55 391
rect 53 390 54 391
rect 52 390 53 391
rect 51 390 52 391
rect 50 390 51 391
rect 49 390 50 391
rect 48 390 49 391
rect 47 390 48 391
rect 46 390 47 391
rect 45 390 46 391
rect 44 390 45 391
rect 43 390 44 391
rect 42 390 43 391
rect 41 390 42 391
rect 40 390 41 391
rect 39 390 40 391
rect 38 390 39 391
rect 37 390 38 391
rect 36 390 37 391
rect 35 390 36 391
rect 34 390 35 391
rect 33 390 34 391
rect 32 390 33 391
rect 31 390 32 391
rect 30 390 31 391
rect 29 390 30 391
rect 28 390 29 391
rect 27 390 28 391
rect 26 390 27 391
rect 25 390 26 391
rect 24 390 25 391
rect 23 390 24 391
rect 22 390 23 391
rect 21 390 22 391
rect 20 390 21 391
rect 19 390 20 391
rect 144 391 145 392
rect 143 391 144 392
rect 142 391 143 392
rect 141 391 142 392
rect 140 391 141 392
rect 130 391 131 392
rect 129 391 130 392
rect 128 391 129 392
rect 127 391 128 392
rect 126 391 127 392
rect 78 391 79 392
rect 77 391 78 392
rect 76 391 77 392
rect 75 391 76 392
rect 74 391 75 392
rect 73 391 74 392
rect 72 391 73 392
rect 71 391 72 392
rect 70 391 71 392
rect 69 391 70 392
rect 68 391 69 392
rect 67 391 68 392
rect 66 391 67 392
rect 65 391 66 392
rect 64 391 65 392
rect 63 391 64 392
rect 62 391 63 392
rect 61 391 62 392
rect 60 391 61 392
rect 59 391 60 392
rect 58 391 59 392
rect 57 391 58 392
rect 56 391 57 392
rect 55 391 56 392
rect 54 391 55 392
rect 53 391 54 392
rect 52 391 53 392
rect 51 391 52 392
rect 50 391 51 392
rect 49 391 50 392
rect 48 391 49 392
rect 47 391 48 392
rect 46 391 47 392
rect 45 391 46 392
rect 44 391 45 392
rect 43 391 44 392
rect 42 391 43 392
rect 41 391 42 392
rect 40 391 41 392
rect 39 391 40 392
rect 38 391 39 392
rect 37 391 38 392
rect 36 391 37 392
rect 35 391 36 392
rect 34 391 35 392
rect 33 391 34 392
rect 32 391 33 392
rect 31 391 32 392
rect 30 391 31 392
rect 29 391 30 392
rect 28 391 29 392
rect 27 391 28 392
rect 26 391 27 392
rect 25 391 26 392
rect 24 391 25 392
rect 23 391 24 392
rect 22 391 23 392
rect 21 391 22 392
rect 20 391 21 392
rect 19 391 20 392
rect 144 392 145 393
rect 143 392 144 393
rect 142 392 143 393
rect 141 392 142 393
rect 129 392 130 393
rect 128 392 129 393
rect 127 392 128 393
rect 126 392 127 393
rect 77 392 78 393
rect 76 392 77 393
rect 75 392 76 393
rect 74 392 75 393
rect 73 392 74 393
rect 72 392 73 393
rect 71 392 72 393
rect 70 392 71 393
rect 69 392 70 393
rect 68 392 69 393
rect 67 392 68 393
rect 66 392 67 393
rect 65 392 66 393
rect 64 392 65 393
rect 63 392 64 393
rect 62 392 63 393
rect 61 392 62 393
rect 60 392 61 393
rect 59 392 60 393
rect 58 392 59 393
rect 57 392 58 393
rect 56 392 57 393
rect 55 392 56 393
rect 54 392 55 393
rect 53 392 54 393
rect 52 392 53 393
rect 51 392 52 393
rect 50 392 51 393
rect 49 392 50 393
rect 48 392 49 393
rect 47 392 48 393
rect 46 392 47 393
rect 45 392 46 393
rect 44 392 45 393
rect 43 392 44 393
rect 42 392 43 393
rect 41 392 42 393
rect 40 392 41 393
rect 39 392 40 393
rect 38 392 39 393
rect 37 392 38 393
rect 36 392 37 393
rect 35 392 36 393
rect 34 392 35 393
rect 33 392 34 393
rect 32 392 33 393
rect 31 392 32 393
rect 30 392 31 393
rect 29 392 30 393
rect 28 392 29 393
rect 27 392 28 393
rect 26 392 27 393
rect 25 392 26 393
rect 24 392 25 393
rect 23 392 24 393
rect 22 392 23 393
rect 21 392 22 393
rect 20 392 21 393
rect 144 393 145 394
rect 143 393 144 394
rect 142 393 143 394
rect 141 393 142 394
rect 129 393 130 394
rect 128 393 129 394
rect 127 393 128 394
rect 126 393 127 394
rect 76 393 77 394
rect 75 393 76 394
rect 74 393 75 394
rect 73 393 74 394
rect 72 393 73 394
rect 71 393 72 394
rect 70 393 71 394
rect 69 393 70 394
rect 68 393 69 394
rect 67 393 68 394
rect 66 393 67 394
rect 65 393 66 394
rect 64 393 65 394
rect 63 393 64 394
rect 62 393 63 394
rect 61 393 62 394
rect 60 393 61 394
rect 59 393 60 394
rect 58 393 59 394
rect 57 393 58 394
rect 56 393 57 394
rect 55 393 56 394
rect 54 393 55 394
rect 53 393 54 394
rect 52 393 53 394
rect 51 393 52 394
rect 50 393 51 394
rect 49 393 50 394
rect 48 393 49 394
rect 47 393 48 394
rect 46 393 47 394
rect 45 393 46 394
rect 44 393 45 394
rect 43 393 44 394
rect 42 393 43 394
rect 41 393 42 394
rect 40 393 41 394
rect 39 393 40 394
rect 38 393 39 394
rect 37 393 38 394
rect 36 393 37 394
rect 35 393 36 394
rect 34 393 35 394
rect 33 393 34 394
rect 32 393 33 394
rect 31 393 32 394
rect 30 393 31 394
rect 29 393 30 394
rect 28 393 29 394
rect 27 393 28 394
rect 26 393 27 394
rect 25 393 26 394
rect 24 393 25 394
rect 23 393 24 394
rect 22 393 23 394
rect 21 393 22 394
rect 144 394 145 395
rect 143 394 144 395
rect 142 394 143 395
rect 141 394 142 395
rect 129 394 130 395
rect 128 394 129 395
rect 127 394 128 395
rect 126 394 127 395
rect 75 394 76 395
rect 74 394 75 395
rect 73 394 74 395
rect 72 394 73 395
rect 71 394 72 395
rect 70 394 71 395
rect 69 394 70 395
rect 68 394 69 395
rect 67 394 68 395
rect 66 394 67 395
rect 65 394 66 395
rect 64 394 65 395
rect 63 394 64 395
rect 62 394 63 395
rect 61 394 62 395
rect 60 394 61 395
rect 59 394 60 395
rect 58 394 59 395
rect 57 394 58 395
rect 56 394 57 395
rect 55 394 56 395
rect 54 394 55 395
rect 53 394 54 395
rect 52 394 53 395
rect 51 394 52 395
rect 50 394 51 395
rect 49 394 50 395
rect 48 394 49 395
rect 47 394 48 395
rect 46 394 47 395
rect 45 394 46 395
rect 44 394 45 395
rect 43 394 44 395
rect 42 394 43 395
rect 41 394 42 395
rect 40 394 41 395
rect 39 394 40 395
rect 38 394 39 395
rect 37 394 38 395
rect 36 394 37 395
rect 35 394 36 395
rect 34 394 35 395
rect 33 394 34 395
rect 32 394 33 395
rect 31 394 32 395
rect 30 394 31 395
rect 29 394 30 395
rect 28 394 29 395
rect 27 394 28 395
rect 26 394 27 395
rect 25 394 26 395
rect 24 394 25 395
rect 23 394 24 395
rect 22 394 23 395
rect 144 395 145 396
rect 143 395 144 396
rect 142 395 143 396
rect 141 395 142 396
rect 140 395 141 396
rect 130 395 131 396
rect 129 395 130 396
rect 128 395 129 396
rect 127 395 128 396
rect 126 395 127 396
rect 74 395 75 396
rect 73 395 74 396
rect 72 395 73 396
rect 71 395 72 396
rect 70 395 71 396
rect 69 395 70 396
rect 68 395 69 396
rect 67 395 68 396
rect 66 395 67 396
rect 65 395 66 396
rect 64 395 65 396
rect 63 395 64 396
rect 62 395 63 396
rect 61 395 62 396
rect 60 395 61 396
rect 59 395 60 396
rect 58 395 59 396
rect 57 395 58 396
rect 56 395 57 396
rect 55 395 56 396
rect 54 395 55 396
rect 53 395 54 396
rect 52 395 53 396
rect 51 395 52 396
rect 50 395 51 396
rect 49 395 50 396
rect 48 395 49 396
rect 47 395 48 396
rect 46 395 47 396
rect 45 395 46 396
rect 44 395 45 396
rect 43 395 44 396
rect 42 395 43 396
rect 41 395 42 396
rect 40 395 41 396
rect 39 395 40 396
rect 38 395 39 396
rect 37 395 38 396
rect 36 395 37 396
rect 35 395 36 396
rect 34 395 35 396
rect 33 395 34 396
rect 32 395 33 396
rect 31 395 32 396
rect 30 395 31 396
rect 29 395 30 396
rect 28 395 29 396
rect 27 395 28 396
rect 26 395 27 396
rect 25 395 26 396
rect 24 395 25 396
rect 23 395 24 396
rect 144 396 145 397
rect 143 396 144 397
rect 142 396 143 397
rect 141 396 142 397
rect 140 396 141 397
rect 139 396 140 397
rect 131 396 132 397
rect 130 396 131 397
rect 129 396 130 397
rect 128 396 129 397
rect 127 396 128 397
rect 126 396 127 397
rect 72 396 73 397
rect 71 396 72 397
rect 70 396 71 397
rect 69 396 70 397
rect 68 396 69 397
rect 67 396 68 397
rect 66 396 67 397
rect 65 396 66 397
rect 64 396 65 397
rect 63 396 64 397
rect 62 396 63 397
rect 61 396 62 397
rect 60 396 61 397
rect 59 396 60 397
rect 58 396 59 397
rect 57 396 58 397
rect 56 396 57 397
rect 55 396 56 397
rect 54 396 55 397
rect 53 396 54 397
rect 52 396 53 397
rect 51 396 52 397
rect 50 396 51 397
rect 49 396 50 397
rect 48 396 49 397
rect 47 396 48 397
rect 46 396 47 397
rect 45 396 46 397
rect 44 396 45 397
rect 43 396 44 397
rect 42 396 43 397
rect 41 396 42 397
rect 40 396 41 397
rect 39 396 40 397
rect 38 396 39 397
rect 37 396 38 397
rect 36 396 37 397
rect 35 396 36 397
rect 34 396 35 397
rect 33 396 34 397
rect 32 396 33 397
rect 31 396 32 397
rect 30 396 31 397
rect 29 396 30 397
rect 28 396 29 397
rect 27 396 28 397
rect 26 396 27 397
rect 25 396 26 397
rect 143 397 144 398
rect 142 397 143 398
rect 141 397 142 398
rect 140 397 141 398
rect 139 397 140 398
rect 138 397 139 398
rect 137 397 138 398
rect 133 397 134 398
rect 132 397 133 398
rect 131 397 132 398
rect 130 397 131 398
rect 129 397 130 398
rect 128 397 129 398
rect 127 397 128 398
rect 70 397 71 398
rect 69 397 70 398
rect 68 397 69 398
rect 67 397 68 398
rect 66 397 67 398
rect 65 397 66 398
rect 64 397 65 398
rect 63 397 64 398
rect 62 397 63 398
rect 61 397 62 398
rect 60 397 61 398
rect 59 397 60 398
rect 58 397 59 398
rect 57 397 58 398
rect 56 397 57 398
rect 55 397 56 398
rect 54 397 55 398
rect 53 397 54 398
rect 52 397 53 398
rect 51 397 52 398
rect 50 397 51 398
rect 49 397 50 398
rect 48 397 49 398
rect 47 397 48 398
rect 46 397 47 398
rect 45 397 46 398
rect 44 397 45 398
rect 43 397 44 398
rect 42 397 43 398
rect 41 397 42 398
rect 40 397 41 398
rect 39 397 40 398
rect 38 397 39 398
rect 37 397 38 398
rect 36 397 37 398
rect 35 397 36 398
rect 34 397 35 398
rect 33 397 34 398
rect 32 397 33 398
rect 31 397 32 398
rect 30 397 31 398
rect 29 397 30 398
rect 28 397 29 398
rect 27 397 28 398
rect 143 398 144 399
rect 142 398 143 399
rect 141 398 142 399
rect 140 398 141 399
rect 139 398 140 399
rect 138 398 139 399
rect 137 398 138 399
rect 136 398 137 399
rect 135 398 136 399
rect 134 398 135 399
rect 133 398 134 399
rect 132 398 133 399
rect 131 398 132 399
rect 130 398 131 399
rect 129 398 130 399
rect 128 398 129 399
rect 127 398 128 399
rect 68 398 69 399
rect 67 398 68 399
rect 66 398 67 399
rect 65 398 66 399
rect 64 398 65 399
rect 63 398 64 399
rect 62 398 63 399
rect 61 398 62 399
rect 60 398 61 399
rect 59 398 60 399
rect 58 398 59 399
rect 57 398 58 399
rect 56 398 57 399
rect 55 398 56 399
rect 54 398 55 399
rect 53 398 54 399
rect 52 398 53 399
rect 51 398 52 399
rect 50 398 51 399
rect 49 398 50 399
rect 48 398 49 399
rect 47 398 48 399
rect 46 398 47 399
rect 45 398 46 399
rect 44 398 45 399
rect 43 398 44 399
rect 42 398 43 399
rect 41 398 42 399
rect 40 398 41 399
rect 39 398 40 399
rect 38 398 39 399
rect 37 398 38 399
rect 36 398 37 399
rect 35 398 36 399
rect 34 398 35 399
rect 33 398 34 399
rect 32 398 33 399
rect 31 398 32 399
rect 30 398 31 399
rect 29 398 30 399
rect 142 399 143 400
rect 141 399 142 400
rect 140 399 141 400
rect 139 399 140 400
rect 138 399 139 400
rect 137 399 138 400
rect 136 399 137 400
rect 135 399 136 400
rect 134 399 135 400
rect 133 399 134 400
rect 132 399 133 400
rect 131 399 132 400
rect 130 399 131 400
rect 129 399 130 400
rect 128 399 129 400
rect 66 399 67 400
rect 65 399 66 400
rect 64 399 65 400
rect 63 399 64 400
rect 62 399 63 400
rect 61 399 62 400
rect 60 399 61 400
rect 59 399 60 400
rect 58 399 59 400
rect 57 399 58 400
rect 56 399 57 400
rect 55 399 56 400
rect 54 399 55 400
rect 53 399 54 400
rect 52 399 53 400
rect 51 399 52 400
rect 50 399 51 400
rect 49 399 50 400
rect 48 399 49 400
rect 47 399 48 400
rect 46 399 47 400
rect 45 399 46 400
rect 44 399 45 400
rect 43 399 44 400
rect 42 399 43 400
rect 41 399 42 400
rect 40 399 41 400
rect 39 399 40 400
rect 38 399 39 400
rect 37 399 38 400
rect 36 399 37 400
rect 35 399 36 400
rect 34 399 35 400
rect 33 399 34 400
rect 32 399 33 400
rect 31 399 32 400
rect 141 400 142 401
rect 140 400 141 401
rect 139 400 140 401
rect 138 400 139 401
rect 137 400 138 401
rect 136 400 137 401
rect 135 400 136 401
rect 134 400 135 401
rect 133 400 134 401
rect 132 400 133 401
rect 131 400 132 401
rect 130 400 131 401
rect 129 400 130 401
rect 128 400 129 401
rect 62 400 63 401
rect 61 400 62 401
rect 60 400 61 401
rect 59 400 60 401
rect 58 400 59 401
rect 57 400 58 401
rect 56 400 57 401
rect 55 400 56 401
rect 54 400 55 401
rect 53 400 54 401
rect 52 400 53 401
rect 51 400 52 401
rect 50 400 51 401
rect 49 400 50 401
rect 48 400 49 401
rect 47 400 48 401
rect 46 400 47 401
rect 45 400 46 401
rect 44 400 45 401
rect 43 400 44 401
rect 42 400 43 401
rect 41 400 42 401
rect 40 400 41 401
rect 39 400 40 401
rect 38 400 39 401
rect 37 400 38 401
rect 36 400 37 401
rect 35 400 36 401
rect 140 401 141 402
rect 139 401 140 402
rect 138 401 139 402
rect 137 401 138 402
rect 136 401 137 402
rect 135 401 136 402
rect 134 401 135 402
rect 133 401 134 402
rect 132 401 133 402
rect 131 401 132 402
rect 130 401 131 402
rect 55 401 56 402
rect 54 401 55 402
rect 53 401 54 402
rect 52 401 53 402
rect 51 401 52 402
rect 50 401 51 402
rect 49 401 50 402
rect 48 401 49 402
rect 47 401 48 402
rect 46 401 47 402
rect 45 401 46 402
rect 44 401 45 402
rect 43 401 44 402
rect 42 401 43 402
rect 138 402 139 403
rect 137 402 138 403
rect 136 402 137 403
rect 135 402 136 403
rect 134 402 135 403
rect 133 402 134 403
rect 132 402 133 403
rect 131 402 132 403
rect 138 406 139 407
rect 137 406 138 407
rect 136 406 137 407
rect 135 406 136 407
rect 134 406 135 407
rect 133 406 134 407
rect 132 406 133 407
rect 140 407 141 408
rect 139 407 140 408
rect 138 407 139 408
rect 137 407 138 408
rect 136 407 137 408
rect 135 407 136 408
rect 134 407 135 408
rect 133 407 134 408
rect 132 407 133 408
rect 131 407 132 408
rect 130 407 131 408
rect 141 408 142 409
rect 140 408 141 409
rect 139 408 140 409
rect 138 408 139 409
rect 137 408 138 409
rect 136 408 137 409
rect 135 408 136 409
rect 134 408 135 409
rect 133 408 134 409
rect 132 408 133 409
rect 131 408 132 409
rect 130 408 131 409
rect 129 408 130 409
rect 142 409 143 410
rect 141 409 142 410
rect 140 409 141 410
rect 139 409 140 410
rect 138 409 139 410
rect 137 409 138 410
rect 136 409 137 410
rect 135 409 136 410
rect 134 409 135 410
rect 133 409 134 410
rect 132 409 133 410
rect 131 409 132 410
rect 130 409 131 410
rect 129 409 130 410
rect 128 409 129 410
rect 82 409 83 410
rect 81 409 82 410
rect 80 409 81 410
rect 79 409 80 410
rect 78 409 79 410
rect 77 409 78 410
rect 76 409 77 410
rect 75 409 76 410
rect 74 409 75 410
rect 73 409 74 410
rect 72 409 73 410
rect 143 410 144 411
rect 142 410 143 411
rect 141 410 142 411
rect 140 410 141 411
rect 139 410 140 411
rect 138 410 139 411
rect 137 410 138 411
rect 136 410 137 411
rect 135 410 136 411
rect 134 410 135 411
rect 133 410 134 411
rect 132 410 133 411
rect 131 410 132 411
rect 130 410 131 411
rect 129 410 130 411
rect 128 410 129 411
rect 127 410 128 411
rect 82 410 83 411
rect 81 410 82 411
rect 80 410 81 411
rect 79 410 80 411
rect 78 410 79 411
rect 77 410 78 411
rect 76 410 77 411
rect 75 410 76 411
rect 74 410 75 411
rect 73 410 74 411
rect 72 410 73 411
rect 71 410 72 411
rect 70 410 71 411
rect 69 410 70 411
rect 68 410 69 411
rect 143 411 144 412
rect 142 411 143 412
rect 141 411 142 412
rect 140 411 141 412
rect 139 411 140 412
rect 138 411 139 412
rect 137 411 138 412
rect 136 411 137 412
rect 135 411 136 412
rect 134 411 135 412
rect 133 411 134 412
rect 132 411 133 412
rect 131 411 132 412
rect 130 411 131 412
rect 129 411 130 412
rect 128 411 129 412
rect 127 411 128 412
rect 82 411 83 412
rect 81 411 82 412
rect 80 411 81 412
rect 79 411 80 412
rect 78 411 79 412
rect 77 411 78 412
rect 76 411 77 412
rect 75 411 76 412
rect 74 411 75 412
rect 73 411 74 412
rect 72 411 73 412
rect 71 411 72 412
rect 70 411 71 412
rect 69 411 70 412
rect 68 411 69 412
rect 67 411 68 412
rect 66 411 67 412
rect 65 411 66 412
rect 144 412 145 413
rect 143 412 144 413
rect 142 412 143 413
rect 141 412 142 413
rect 140 412 141 413
rect 139 412 140 413
rect 131 412 132 413
rect 130 412 131 413
rect 129 412 130 413
rect 128 412 129 413
rect 127 412 128 413
rect 126 412 127 413
rect 82 412 83 413
rect 81 412 82 413
rect 80 412 81 413
rect 79 412 80 413
rect 78 412 79 413
rect 77 412 78 413
rect 76 412 77 413
rect 75 412 76 413
rect 74 412 75 413
rect 73 412 74 413
rect 72 412 73 413
rect 71 412 72 413
rect 70 412 71 413
rect 69 412 70 413
rect 68 412 69 413
rect 67 412 68 413
rect 66 412 67 413
rect 65 412 66 413
rect 64 412 65 413
rect 35 412 36 413
rect 34 412 35 413
rect 33 412 34 413
rect 32 412 33 413
rect 31 412 32 413
rect 30 412 31 413
rect 29 412 30 413
rect 28 412 29 413
rect 27 412 28 413
rect 26 412 27 413
rect 25 412 26 413
rect 24 412 25 413
rect 23 412 24 413
rect 22 412 23 413
rect 21 412 22 413
rect 20 412 21 413
rect 144 413 145 414
rect 143 413 144 414
rect 142 413 143 414
rect 141 413 142 414
rect 140 413 141 414
rect 130 413 131 414
rect 129 413 130 414
rect 128 413 129 414
rect 127 413 128 414
rect 126 413 127 414
rect 82 413 83 414
rect 81 413 82 414
rect 80 413 81 414
rect 79 413 80 414
rect 78 413 79 414
rect 77 413 78 414
rect 76 413 77 414
rect 75 413 76 414
rect 74 413 75 414
rect 73 413 74 414
rect 72 413 73 414
rect 71 413 72 414
rect 70 413 71 414
rect 69 413 70 414
rect 68 413 69 414
rect 67 413 68 414
rect 66 413 67 414
rect 65 413 66 414
rect 64 413 65 414
rect 63 413 64 414
rect 62 413 63 414
rect 34 413 35 414
rect 33 413 34 414
rect 32 413 33 414
rect 31 413 32 414
rect 30 413 31 414
rect 29 413 30 414
rect 28 413 29 414
rect 27 413 28 414
rect 26 413 27 414
rect 25 413 26 414
rect 24 413 25 414
rect 23 413 24 414
rect 22 413 23 414
rect 21 413 22 414
rect 20 413 21 414
rect 19 413 20 414
rect 144 414 145 415
rect 143 414 144 415
rect 142 414 143 415
rect 141 414 142 415
rect 140 414 141 415
rect 130 414 131 415
rect 129 414 130 415
rect 128 414 129 415
rect 127 414 128 415
rect 126 414 127 415
rect 82 414 83 415
rect 81 414 82 415
rect 80 414 81 415
rect 79 414 80 415
rect 78 414 79 415
rect 77 414 78 415
rect 76 414 77 415
rect 75 414 76 415
rect 74 414 75 415
rect 73 414 74 415
rect 72 414 73 415
rect 71 414 72 415
rect 70 414 71 415
rect 69 414 70 415
rect 68 414 69 415
rect 67 414 68 415
rect 66 414 67 415
rect 65 414 66 415
rect 64 414 65 415
rect 63 414 64 415
rect 62 414 63 415
rect 61 414 62 415
rect 34 414 35 415
rect 33 414 34 415
rect 32 414 33 415
rect 31 414 32 415
rect 30 414 31 415
rect 29 414 30 415
rect 28 414 29 415
rect 27 414 28 415
rect 26 414 27 415
rect 25 414 26 415
rect 24 414 25 415
rect 23 414 24 415
rect 22 414 23 415
rect 21 414 22 415
rect 20 414 21 415
rect 19 414 20 415
rect 144 415 145 416
rect 143 415 144 416
rect 142 415 143 416
rect 141 415 142 416
rect 129 415 130 416
rect 128 415 129 416
rect 127 415 128 416
rect 126 415 127 416
rect 82 415 83 416
rect 81 415 82 416
rect 80 415 81 416
rect 79 415 80 416
rect 78 415 79 416
rect 77 415 78 416
rect 76 415 77 416
rect 75 415 76 416
rect 74 415 75 416
rect 73 415 74 416
rect 72 415 73 416
rect 71 415 72 416
rect 70 415 71 416
rect 69 415 70 416
rect 68 415 69 416
rect 67 415 68 416
rect 66 415 67 416
rect 65 415 66 416
rect 64 415 65 416
rect 63 415 64 416
rect 62 415 63 416
rect 61 415 62 416
rect 60 415 61 416
rect 59 415 60 416
rect 33 415 34 416
rect 32 415 33 416
rect 31 415 32 416
rect 30 415 31 416
rect 29 415 30 416
rect 28 415 29 416
rect 27 415 28 416
rect 26 415 27 416
rect 25 415 26 416
rect 24 415 25 416
rect 23 415 24 416
rect 22 415 23 416
rect 21 415 22 416
rect 20 415 21 416
rect 19 415 20 416
rect 144 416 145 417
rect 143 416 144 417
rect 142 416 143 417
rect 141 416 142 417
rect 129 416 130 417
rect 128 416 129 417
rect 127 416 128 417
rect 126 416 127 417
rect 82 416 83 417
rect 81 416 82 417
rect 80 416 81 417
rect 79 416 80 417
rect 78 416 79 417
rect 77 416 78 417
rect 76 416 77 417
rect 75 416 76 417
rect 74 416 75 417
rect 73 416 74 417
rect 72 416 73 417
rect 71 416 72 417
rect 70 416 71 417
rect 69 416 70 417
rect 68 416 69 417
rect 67 416 68 417
rect 66 416 67 417
rect 65 416 66 417
rect 64 416 65 417
rect 63 416 64 417
rect 62 416 63 417
rect 61 416 62 417
rect 60 416 61 417
rect 59 416 60 417
rect 58 416 59 417
rect 33 416 34 417
rect 32 416 33 417
rect 31 416 32 417
rect 30 416 31 417
rect 29 416 30 417
rect 28 416 29 417
rect 27 416 28 417
rect 26 416 27 417
rect 25 416 26 417
rect 24 416 25 417
rect 23 416 24 417
rect 22 416 23 417
rect 21 416 22 417
rect 20 416 21 417
rect 19 416 20 417
rect 18 416 19 417
rect 144 417 145 418
rect 143 417 144 418
rect 142 417 143 418
rect 141 417 142 418
rect 140 417 141 418
rect 130 417 131 418
rect 129 417 130 418
rect 128 417 129 418
rect 127 417 128 418
rect 126 417 127 418
rect 82 417 83 418
rect 81 417 82 418
rect 80 417 81 418
rect 79 417 80 418
rect 78 417 79 418
rect 77 417 78 418
rect 76 417 77 418
rect 75 417 76 418
rect 74 417 75 418
rect 73 417 74 418
rect 72 417 73 418
rect 71 417 72 418
rect 70 417 71 418
rect 69 417 70 418
rect 68 417 69 418
rect 67 417 68 418
rect 66 417 67 418
rect 65 417 66 418
rect 64 417 65 418
rect 63 417 64 418
rect 62 417 63 418
rect 61 417 62 418
rect 60 417 61 418
rect 59 417 60 418
rect 58 417 59 418
rect 57 417 58 418
rect 32 417 33 418
rect 31 417 32 418
rect 30 417 31 418
rect 29 417 30 418
rect 28 417 29 418
rect 27 417 28 418
rect 26 417 27 418
rect 25 417 26 418
rect 24 417 25 418
rect 23 417 24 418
rect 22 417 23 418
rect 21 417 22 418
rect 20 417 21 418
rect 19 417 20 418
rect 18 417 19 418
rect 144 418 145 419
rect 143 418 144 419
rect 142 418 143 419
rect 141 418 142 419
rect 140 418 141 419
rect 130 418 131 419
rect 129 418 130 419
rect 128 418 129 419
rect 127 418 128 419
rect 126 418 127 419
rect 82 418 83 419
rect 81 418 82 419
rect 80 418 81 419
rect 79 418 80 419
rect 78 418 79 419
rect 77 418 78 419
rect 76 418 77 419
rect 75 418 76 419
rect 74 418 75 419
rect 73 418 74 419
rect 72 418 73 419
rect 71 418 72 419
rect 70 418 71 419
rect 69 418 70 419
rect 68 418 69 419
rect 67 418 68 419
rect 66 418 67 419
rect 65 418 66 419
rect 64 418 65 419
rect 63 418 64 419
rect 62 418 63 419
rect 61 418 62 419
rect 60 418 61 419
rect 59 418 60 419
rect 58 418 59 419
rect 57 418 58 419
rect 56 418 57 419
rect 32 418 33 419
rect 31 418 32 419
rect 30 418 31 419
rect 29 418 30 419
rect 28 418 29 419
rect 27 418 28 419
rect 26 418 27 419
rect 25 418 26 419
rect 24 418 25 419
rect 23 418 24 419
rect 22 418 23 419
rect 21 418 22 419
rect 20 418 21 419
rect 19 418 20 419
rect 18 418 19 419
rect 17 418 18 419
rect 144 419 145 420
rect 143 419 144 420
rect 142 419 143 420
rect 141 419 142 420
rect 140 419 141 420
rect 139 419 140 420
rect 131 419 132 420
rect 130 419 131 420
rect 129 419 130 420
rect 128 419 129 420
rect 127 419 128 420
rect 126 419 127 420
rect 82 419 83 420
rect 81 419 82 420
rect 80 419 81 420
rect 79 419 80 420
rect 78 419 79 420
rect 77 419 78 420
rect 76 419 77 420
rect 75 419 76 420
rect 74 419 75 420
rect 73 419 74 420
rect 72 419 73 420
rect 71 419 72 420
rect 70 419 71 420
rect 69 419 70 420
rect 68 419 69 420
rect 67 419 68 420
rect 66 419 67 420
rect 65 419 66 420
rect 64 419 65 420
rect 63 419 64 420
rect 62 419 63 420
rect 61 419 62 420
rect 60 419 61 420
rect 59 419 60 420
rect 58 419 59 420
rect 57 419 58 420
rect 56 419 57 420
rect 31 419 32 420
rect 30 419 31 420
rect 29 419 30 420
rect 28 419 29 420
rect 27 419 28 420
rect 26 419 27 420
rect 25 419 26 420
rect 24 419 25 420
rect 23 419 24 420
rect 22 419 23 420
rect 21 419 22 420
rect 20 419 21 420
rect 19 419 20 420
rect 18 419 19 420
rect 17 419 18 420
rect 143 420 144 421
rect 142 420 143 421
rect 141 420 142 421
rect 140 420 141 421
rect 139 420 140 421
rect 138 420 139 421
rect 137 420 138 421
rect 136 420 137 421
rect 135 420 136 421
rect 134 420 135 421
rect 133 420 134 421
rect 132 420 133 421
rect 131 420 132 421
rect 130 420 131 421
rect 129 420 130 421
rect 128 420 129 421
rect 127 420 128 421
rect 82 420 83 421
rect 81 420 82 421
rect 80 420 81 421
rect 79 420 80 421
rect 78 420 79 421
rect 77 420 78 421
rect 76 420 77 421
rect 75 420 76 421
rect 74 420 75 421
rect 73 420 74 421
rect 72 420 73 421
rect 71 420 72 421
rect 70 420 71 421
rect 69 420 70 421
rect 68 420 69 421
rect 67 420 68 421
rect 66 420 67 421
rect 65 420 66 421
rect 64 420 65 421
rect 63 420 64 421
rect 62 420 63 421
rect 61 420 62 421
rect 60 420 61 421
rect 59 420 60 421
rect 58 420 59 421
rect 57 420 58 421
rect 56 420 57 421
rect 55 420 56 421
rect 31 420 32 421
rect 30 420 31 421
rect 29 420 30 421
rect 28 420 29 421
rect 27 420 28 421
rect 26 420 27 421
rect 25 420 26 421
rect 24 420 25 421
rect 23 420 24 421
rect 22 420 23 421
rect 21 420 22 421
rect 20 420 21 421
rect 19 420 20 421
rect 18 420 19 421
rect 17 420 18 421
rect 143 421 144 422
rect 142 421 143 422
rect 141 421 142 422
rect 140 421 141 422
rect 139 421 140 422
rect 138 421 139 422
rect 137 421 138 422
rect 136 421 137 422
rect 135 421 136 422
rect 134 421 135 422
rect 133 421 134 422
rect 132 421 133 422
rect 131 421 132 422
rect 130 421 131 422
rect 129 421 130 422
rect 128 421 129 422
rect 127 421 128 422
rect 82 421 83 422
rect 81 421 82 422
rect 80 421 81 422
rect 79 421 80 422
rect 78 421 79 422
rect 77 421 78 422
rect 76 421 77 422
rect 75 421 76 422
rect 74 421 75 422
rect 73 421 74 422
rect 72 421 73 422
rect 71 421 72 422
rect 70 421 71 422
rect 69 421 70 422
rect 68 421 69 422
rect 67 421 68 422
rect 66 421 67 422
rect 65 421 66 422
rect 64 421 65 422
rect 63 421 64 422
rect 62 421 63 422
rect 61 421 62 422
rect 60 421 61 422
rect 59 421 60 422
rect 58 421 59 422
rect 57 421 58 422
rect 56 421 57 422
rect 55 421 56 422
rect 54 421 55 422
rect 31 421 32 422
rect 30 421 31 422
rect 29 421 30 422
rect 28 421 29 422
rect 27 421 28 422
rect 26 421 27 422
rect 25 421 26 422
rect 24 421 25 422
rect 23 421 24 422
rect 22 421 23 422
rect 21 421 22 422
rect 20 421 21 422
rect 19 421 20 422
rect 18 421 19 422
rect 17 421 18 422
rect 16 421 17 422
rect 142 422 143 423
rect 141 422 142 423
rect 140 422 141 423
rect 139 422 140 423
rect 138 422 139 423
rect 137 422 138 423
rect 136 422 137 423
rect 135 422 136 423
rect 134 422 135 423
rect 133 422 134 423
rect 132 422 133 423
rect 131 422 132 423
rect 130 422 131 423
rect 129 422 130 423
rect 128 422 129 423
rect 82 422 83 423
rect 81 422 82 423
rect 80 422 81 423
rect 79 422 80 423
rect 78 422 79 423
rect 77 422 78 423
rect 76 422 77 423
rect 75 422 76 423
rect 74 422 75 423
rect 73 422 74 423
rect 72 422 73 423
rect 71 422 72 423
rect 70 422 71 423
rect 69 422 70 423
rect 68 422 69 423
rect 67 422 68 423
rect 66 422 67 423
rect 65 422 66 423
rect 64 422 65 423
rect 63 422 64 423
rect 62 422 63 423
rect 61 422 62 423
rect 60 422 61 423
rect 59 422 60 423
rect 58 422 59 423
rect 57 422 58 423
rect 56 422 57 423
rect 55 422 56 423
rect 54 422 55 423
rect 53 422 54 423
rect 31 422 32 423
rect 30 422 31 423
rect 29 422 30 423
rect 28 422 29 423
rect 27 422 28 423
rect 26 422 27 423
rect 25 422 26 423
rect 24 422 25 423
rect 23 422 24 423
rect 22 422 23 423
rect 21 422 22 423
rect 20 422 21 423
rect 19 422 20 423
rect 18 422 19 423
rect 17 422 18 423
rect 16 422 17 423
rect 141 423 142 424
rect 140 423 141 424
rect 139 423 140 424
rect 138 423 139 424
rect 137 423 138 424
rect 136 423 137 424
rect 135 423 136 424
rect 134 423 135 424
rect 133 423 134 424
rect 132 423 133 424
rect 131 423 132 424
rect 130 423 131 424
rect 129 423 130 424
rect 82 423 83 424
rect 81 423 82 424
rect 80 423 81 424
rect 79 423 80 424
rect 78 423 79 424
rect 77 423 78 424
rect 76 423 77 424
rect 75 423 76 424
rect 74 423 75 424
rect 73 423 74 424
rect 72 423 73 424
rect 71 423 72 424
rect 70 423 71 424
rect 69 423 70 424
rect 68 423 69 424
rect 67 423 68 424
rect 66 423 67 424
rect 65 423 66 424
rect 64 423 65 424
rect 63 423 64 424
rect 62 423 63 424
rect 61 423 62 424
rect 60 423 61 424
rect 59 423 60 424
rect 58 423 59 424
rect 57 423 58 424
rect 56 423 57 424
rect 55 423 56 424
rect 54 423 55 424
rect 53 423 54 424
rect 52 423 53 424
rect 30 423 31 424
rect 29 423 30 424
rect 28 423 29 424
rect 27 423 28 424
rect 26 423 27 424
rect 25 423 26 424
rect 24 423 25 424
rect 23 423 24 424
rect 22 423 23 424
rect 21 423 22 424
rect 20 423 21 424
rect 19 423 20 424
rect 18 423 19 424
rect 17 423 18 424
rect 16 423 17 424
rect 140 424 141 425
rect 139 424 140 425
rect 138 424 139 425
rect 137 424 138 425
rect 136 424 137 425
rect 135 424 136 425
rect 134 424 135 425
rect 133 424 134 425
rect 132 424 133 425
rect 131 424 132 425
rect 130 424 131 425
rect 82 424 83 425
rect 81 424 82 425
rect 80 424 81 425
rect 79 424 80 425
rect 78 424 79 425
rect 77 424 78 425
rect 76 424 77 425
rect 75 424 76 425
rect 74 424 75 425
rect 73 424 74 425
rect 72 424 73 425
rect 71 424 72 425
rect 70 424 71 425
rect 69 424 70 425
rect 68 424 69 425
rect 67 424 68 425
rect 66 424 67 425
rect 65 424 66 425
rect 64 424 65 425
rect 63 424 64 425
rect 62 424 63 425
rect 61 424 62 425
rect 60 424 61 425
rect 59 424 60 425
rect 58 424 59 425
rect 57 424 58 425
rect 56 424 57 425
rect 55 424 56 425
rect 54 424 55 425
rect 53 424 54 425
rect 52 424 53 425
rect 51 424 52 425
rect 30 424 31 425
rect 29 424 30 425
rect 28 424 29 425
rect 27 424 28 425
rect 26 424 27 425
rect 25 424 26 425
rect 24 424 25 425
rect 23 424 24 425
rect 22 424 23 425
rect 21 424 22 425
rect 20 424 21 425
rect 19 424 20 425
rect 18 424 19 425
rect 17 424 18 425
rect 16 424 17 425
rect 137 425 138 426
rect 136 425 137 426
rect 135 425 136 426
rect 134 425 135 426
rect 133 425 134 426
rect 132 425 133 426
rect 82 425 83 426
rect 81 425 82 426
rect 80 425 81 426
rect 79 425 80 426
rect 78 425 79 426
rect 77 425 78 426
rect 76 425 77 426
rect 75 425 76 426
rect 74 425 75 426
rect 73 425 74 426
rect 72 425 73 426
rect 71 425 72 426
rect 70 425 71 426
rect 69 425 70 426
rect 68 425 69 426
rect 67 425 68 426
rect 66 425 67 426
rect 65 425 66 426
rect 64 425 65 426
rect 63 425 64 426
rect 62 425 63 426
rect 61 425 62 426
rect 60 425 61 426
rect 59 425 60 426
rect 58 425 59 426
rect 57 425 58 426
rect 56 425 57 426
rect 55 425 56 426
rect 54 425 55 426
rect 53 425 54 426
rect 52 425 53 426
rect 51 425 52 426
rect 30 425 31 426
rect 29 425 30 426
rect 28 425 29 426
rect 27 425 28 426
rect 26 425 27 426
rect 25 425 26 426
rect 24 425 25 426
rect 23 425 24 426
rect 22 425 23 426
rect 21 425 22 426
rect 20 425 21 426
rect 19 425 20 426
rect 18 425 19 426
rect 17 425 18 426
rect 16 425 17 426
rect 82 426 83 427
rect 81 426 82 427
rect 80 426 81 427
rect 79 426 80 427
rect 78 426 79 427
rect 77 426 78 427
rect 76 426 77 427
rect 75 426 76 427
rect 74 426 75 427
rect 73 426 74 427
rect 72 426 73 427
rect 71 426 72 427
rect 70 426 71 427
rect 69 426 70 427
rect 68 426 69 427
rect 67 426 68 427
rect 66 426 67 427
rect 65 426 66 427
rect 64 426 65 427
rect 63 426 64 427
rect 62 426 63 427
rect 61 426 62 427
rect 60 426 61 427
rect 59 426 60 427
rect 58 426 59 427
rect 57 426 58 427
rect 56 426 57 427
rect 55 426 56 427
rect 54 426 55 427
rect 53 426 54 427
rect 52 426 53 427
rect 51 426 52 427
rect 50 426 51 427
rect 30 426 31 427
rect 29 426 30 427
rect 28 426 29 427
rect 27 426 28 427
rect 26 426 27 427
rect 25 426 26 427
rect 24 426 25 427
rect 23 426 24 427
rect 22 426 23 427
rect 21 426 22 427
rect 20 426 21 427
rect 19 426 20 427
rect 18 426 19 427
rect 17 426 18 427
rect 16 426 17 427
rect 82 427 83 428
rect 81 427 82 428
rect 80 427 81 428
rect 79 427 80 428
rect 78 427 79 428
rect 77 427 78 428
rect 76 427 77 428
rect 75 427 76 428
rect 74 427 75 428
rect 73 427 74 428
rect 72 427 73 428
rect 71 427 72 428
rect 70 427 71 428
rect 69 427 70 428
rect 68 427 69 428
rect 67 427 68 428
rect 66 427 67 428
rect 65 427 66 428
rect 64 427 65 428
rect 63 427 64 428
rect 62 427 63 428
rect 61 427 62 428
rect 60 427 61 428
rect 59 427 60 428
rect 58 427 59 428
rect 57 427 58 428
rect 56 427 57 428
rect 55 427 56 428
rect 54 427 55 428
rect 53 427 54 428
rect 52 427 53 428
rect 51 427 52 428
rect 50 427 51 428
rect 49 427 50 428
rect 30 427 31 428
rect 29 427 30 428
rect 28 427 29 428
rect 27 427 28 428
rect 26 427 27 428
rect 25 427 26 428
rect 24 427 25 428
rect 23 427 24 428
rect 22 427 23 428
rect 21 427 22 428
rect 20 427 21 428
rect 19 427 20 428
rect 18 427 19 428
rect 17 427 18 428
rect 16 427 17 428
rect 15 427 16 428
rect 82 428 83 429
rect 81 428 82 429
rect 80 428 81 429
rect 79 428 80 429
rect 78 428 79 429
rect 77 428 78 429
rect 76 428 77 429
rect 75 428 76 429
rect 74 428 75 429
rect 73 428 74 429
rect 72 428 73 429
rect 71 428 72 429
rect 70 428 71 429
rect 69 428 70 429
rect 68 428 69 429
rect 67 428 68 429
rect 66 428 67 429
rect 65 428 66 429
rect 64 428 65 429
rect 63 428 64 429
rect 62 428 63 429
rect 61 428 62 429
rect 60 428 61 429
rect 59 428 60 429
rect 58 428 59 429
rect 57 428 58 429
rect 56 428 57 429
rect 55 428 56 429
rect 54 428 55 429
rect 53 428 54 429
rect 52 428 53 429
rect 51 428 52 429
rect 50 428 51 429
rect 49 428 50 429
rect 48 428 49 429
rect 30 428 31 429
rect 29 428 30 429
rect 28 428 29 429
rect 27 428 28 429
rect 26 428 27 429
rect 25 428 26 429
rect 24 428 25 429
rect 23 428 24 429
rect 22 428 23 429
rect 21 428 22 429
rect 20 428 21 429
rect 19 428 20 429
rect 18 428 19 429
rect 17 428 18 429
rect 16 428 17 429
rect 15 428 16 429
rect 82 429 83 430
rect 81 429 82 430
rect 80 429 81 430
rect 79 429 80 430
rect 78 429 79 430
rect 77 429 78 430
rect 76 429 77 430
rect 75 429 76 430
rect 74 429 75 430
rect 73 429 74 430
rect 72 429 73 430
rect 71 429 72 430
rect 70 429 71 430
rect 69 429 70 430
rect 68 429 69 430
rect 67 429 68 430
rect 66 429 67 430
rect 65 429 66 430
rect 64 429 65 430
rect 63 429 64 430
rect 62 429 63 430
rect 61 429 62 430
rect 60 429 61 430
rect 59 429 60 430
rect 58 429 59 430
rect 57 429 58 430
rect 56 429 57 430
rect 55 429 56 430
rect 54 429 55 430
rect 53 429 54 430
rect 52 429 53 430
rect 51 429 52 430
rect 50 429 51 430
rect 49 429 50 430
rect 48 429 49 430
rect 47 429 48 430
rect 30 429 31 430
rect 29 429 30 430
rect 28 429 29 430
rect 27 429 28 430
rect 26 429 27 430
rect 25 429 26 430
rect 24 429 25 430
rect 23 429 24 430
rect 22 429 23 430
rect 21 429 22 430
rect 20 429 21 430
rect 19 429 20 430
rect 18 429 19 430
rect 17 429 18 430
rect 16 429 17 430
rect 15 429 16 430
rect 144 430 145 431
rect 143 430 144 431
rect 142 430 143 431
rect 141 430 142 431
rect 140 430 141 431
rect 139 430 140 431
rect 138 430 139 431
rect 137 430 138 431
rect 136 430 137 431
rect 135 430 136 431
rect 134 430 135 431
rect 133 430 134 431
rect 132 430 133 431
rect 131 430 132 431
rect 130 430 131 431
rect 129 430 130 431
rect 128 430 129 431
rect 127 430 128 431
rect 126 430 127 431
rect 125 430 126 431
rect 124 430 125 431
rect 123 430 124 431
rect 122 430 123 431
rect 121 430 122 431
rect 120 430 121 431
rect 119 430 120 431
rect 118 430 119 431
rect 117 430 118 431
rect 82 430 83 431
rect 81 430 82 431
rect 80 430 81 431
rect 79 430 80 431
rect 78 430 79 431
rect 77 430 78 431
rect 76 430 77 431
rect 75 430 76 431
rect 74 430 75 431
rect 73 430 74 431
rect 72 430 73 431
rect 71 430 72 431
rect 70 430 71 431
rect 69 430 70 431
rect 68 430 69 431
rect 67 430 68 431
rect 65 430 66 431
rect 64 430 65 431
rect 63 430 64 431
rect 62 430 63 431
rect 61 430 62 431
rect 60 430 61 431
rect 59 430 60 431
rect 58 430 59 431
rect 57 430 58 431
rect 56 430 57 431
rect 55 430 56 431
rect 54 430 55 431
rect 53 430 54 431
rect 52 430 53 431
rect 51 430 52 431
rect 50 430 51 431
rect 49 430 50 431
rect 48 430 49 431
rect 47 430 48 431
rect 30 430 31 431
rect 29 430 30 431
rect 28 430 29 431
rect 27 430 28 431
rect 26 430 27 431
rect 25 430 26 431
rect 24 430 25 431
rect 23 430 24 431
rect 22 430 23 431
rect 21 430 22 431
rect 20 430 21 431
rect 19 430 20 431
rect 18 430 19 431
rect 17 430 18 431
rect 16 430 17 431
rect 15 430 16 431
rect 144 431 145 432
rect 143 431 144 432
rect 142 431 143 432
rect 141 431 142 432
rect 140 431 141 432
rect 139 431 140 432
rect 138 431 139 432
rect 137 431 138 432
rect 136 431 137 432
rect 135 431 136 432
rect 134 431 135 432
rect 133 431 134 432
rect 132 431 133 432
rect 131 431 132 432
rect 130 431 131 432
rect 129 431 130 432
rect 128 431 129 432
rect 127 431 128 432
rect 126 431 127 432
rect 125 431 126 432
rect 124 431 125 432
rect 123 431 124 432
rect 122 431 123 432
rect 121 431 122 432
rect 120 431 121 432
rect 119 431 120 432
rect 118 431 119 432
rect 117 431 118 432
rect 82 431 83 432
rect 81 431 82 432
rect 80 431 81 432
rect 79 431 80 432
rect 78 431 79 432
rect 77 431 78 432
rect 76 431 77 432
rect 75 431 76 432
rect 74 431 75 432
rect 73 431 74 432
rect 72 431 73 432
rect 71 431 72 432
rect 70 431 71 432
rect 69 431 70 432
rect 68 431 69 432
rect 67 431 68 432
rect 64 431 65 432
rect 63 431 64 432
rect 62 431 63 432
rect 61 431 62 432
rect 60 431 61 432
rect 59 431 60 432
rect 58 431 59 432
rect 57 431 58 432
rect 56 431 57 432
rect 55 431 56 432
rect 54 431 55 432
rect 53 431 54 432
rect 52 431 53 432
rect 51 431 52 432
rect 50 431 51 432
rect 49 431 50 432
rect 48 431 49 432
rect 47 431 48 432
rect 46 431 47 432
rect 30 431 31 432
rect 29 431 30 432
rect 28 431 29 432
rect 27 431 28 432
rect 26 431 27 432
rect 25 431 26 432
rect 24 431 25 432
rect 23 431 24 432
rect 22 431 23 432
rect 21 431 22 432
rect 20 431 21 432
rect 19 431 20 432
rect 18 431 19 432
rect 17 431 18 432
rect 16 431 17 432
rect 15 431 16 432
rect 144 432 145 433
rect 143 432 144 433
rect 142 432 143 433
rect 141 432 142 433
rect 140 432 141 433
rect 139 432 140 433
rect 138 432 139 433
rect 137 432 138 433
rect 136 432 137 433
rect 135 432 136 433
rect 134 432 135 433
rect 133 432 134 433
rect 132 432 133 433
rect 131 432 132 433
rect 130 432 131 433
rect 129 432 130 433
rect 128 432 129 433
rect 127 432 128 433
rect 126 432 127 433
rect 125 432 126 433
rect 124 432 125 433
rect 123 432 124 433
rect 122 432 123 433
rect 121 432 122 433
rect 120 432 121 433
rect 119 432 120 433
rect 118 432 119 433
rect 117 432 118 433
rect 82 432 83 433
rect 81 432 82 433
rect 80 432 81 433
rect 79 432 80 433
rect 78 432 79 433
rect 77 432 78 433
rect 76 432 77 433
rect 75 432 76 433
rect 74 432 75 433
rect 73 432 74 433
rect 72 432 73 433
rect 71 432 72 433
rect 70 432 71 433
rect 69 432 70 433
rect 68 432 69 433
rect 67 432 68 433
rect 63 432 64 433
rect 62 432 63 433
rect 61 432 62 433
rect 60 432 61 433
rect 59 432 60 433
rect 58 432 59 433
rect 57 432 58 433
rect 56 432 57 433
rect 55 432 56 433
rect 54 432 55 433
rect 53 432 54 433
rect 52 432 53 433
rect 51 432 52 433
rect 50 432 51 433
rect 49 432 50 433
rect 48 432 49 433
rect 47 432 48 433
rect 46 432 47 433
rect 45 432 46 433
rect 31 432 32 433
rect 30 432 31 433
rect 29 432 30 433
rect 28 432 29 433
rect 27 432 28 433
rect 26 432 27 433
rect 25 432 26 433
rect 24 432 25 433
rect 23 432 24 433
rect 22 432 23 433
rect 21 432 22 433
rect 20 432 21 433
rect 19 432 20 433
rect 18 432 19 433
rect 17 432 18 433
rect 16 432 17 433
rect 15 432 16 433
rect 144 433 145 434
rect 143 433 144 434
rect 142 433 143 434
rect 141 433 142 434
rect 140 433 141 434
rect 139 433 140 434
rect 138 433 139 434
rect 137 433 138 434
rect 136 433 137 434
rect 135 433 136 434
rect 134 433 135 434
rect 133 433 134 434
rect 132 433 133 434
rect 131 433 132 434
rect 130 433 131 434
rect 129 433 130 434
rect 128 433 129 434
rect 127 433 128 434
rect 126 433 127 434
rect 125 433 126 434
rect 124 433 125 434
rect 123 433 124 434
rect 122 433 123 434
rect 121 433 122 434
rect 120 433 121 434
rect 119 433 120 434
rect 118 433 119 434
rect 117 433 118 434
rect 82 433 83 434
rect 81 433 82 434
rect 80 433 81 434
rect 79 433 80 434
rect 78 433 79 434
rect 77 433 78 434
rect 76 433 77 434
rect 75 433 76 434
rect 74 433 75 434
rect 73 433 74 434
rect 72 433 73 434
rect 71 433 72 434
rect 70 433 71 434
rect 69 433 70 434
rect 68 433 69 434
rect 67 433 68 434
rect 62 433 63 434
rect 61 433 62 434
rect 60 433 61 434
rect 59 433 60 434
rect 58 433 59 434
rect 57 433 58 434
rect 56 433 57 434
rect 55 433 56 434
rect 54 433 55 434
rect 53 433 54 434
rect 52 433 53 434
rect 51 433 52 434
rect 50 433 51 434
rect 49 433 50 434
rect 48 433 49 434
rect 47 433 48 434
rect 46 433 47 434
rect 45 433 46 434
rect 44 433 45 434
rect 31 433 32 434
rect 30 433 31 434
rect 29 433 30 434
rect 28 433 29 434
rect 27 433 28 434
rect 26 433 27 434
rect 25 433 26 434
rect 24 433 25 434
rect 23 433 24 434
rect 22 433 23 434
rect 21 433 22 434
rect 20 433 21 434
rect 19 433 20 434
rect 18 433 19 434
rect 17 433 18 434
rect 16 433 17 434
rect 15 433 16 434
rect 144 434 145 435
rect 143 434 144 435
rect 142 434 143 435
rect 141 434 142 435
rect 140 434 141 435
rect 139 434 140 435
rect 138 434 139 435
rect 137 434 138 435
rect 136 434 137 435
rect 135 434 136 435
rect 134 434 135 435
rect 133 434 134 435
rect 132 434 133 435
rect 131 434 132 435
rect 130 434 131 435
rect 129 434 130 435
rect 128 434 129 435
rect 127 434 128 435
rect 126 434 127 435
rect 125 434 126 435
rect 124 434 125 435
rect 123 434 124 435
rect 122 434 123 435
rect 121 434 122 435
rect 120 434 121 435
rect 119 434 120 435
rect 118 434 119 435
rect 117 434 118 435
rect 82 434 83 435
rect 81 434 82 435
rect 80 434 81 435
rect 79 434 80 435
rect 78 434 79 435
rect 77 434 78 435
rect 76 434 77 435
rect 75 434 76 435
rect 74 434 75 435
rect 73 434 74 435
rect 72 434 73 435
rect 71 434 72 435
rect 70 434 71 435
rect 69 434 70 435
rect 68 434 69 435
rect 67 434 68 435
rect 61 434 62 435
rect 60 434 61 435
rect 59 434 60 435
rect 58 434 59 435
rect 57 434 58 435
rect 56 434 57 435
rect 55 434 56 435
rect 54 434 55 435
rect 53 434 54 435
rect 52 434 53 435
rect 51 434 52 435
rect 50 434 51 435
rect 49 434 50 435
rect 48 434 49 435
rect 47 434 48 435
rect 46 434 47 435
rect 45 434 46 435
rect 44 434 45 435
rect 43 434 44 435
rect 42 434 43 435
rect 32 434 33 435
rect 31 434 32 435
rect 30 434 31 435
rect 29 434 30 435
rect 28 434 29 435
rect 27 434 28 435
rect 26 434 27 435
rect 25 434 26 435
rect 24 434 25 435
rect 23 434 24 435
rect 22 434 23 435
rect 21 434 22 435
rect 20 434 21 435
rect 19 434 20 435
rect 18 434 19 435
rect 17 434 18 435
rect 16 434 17 435
rect 15 434 16 435
rect 144 435 145 436
rect 143 435 144 436
rect 142 435 143 436
rect 141 435 142 436
rect 140 435 141 436
rect 139 435 140 436
rect 138 435 139 436
rect 137 435 138 436
rect 136 435 137 436
rect 135 435 136 436
rect 134 435 135 436
rect 133 435 134 436
rect 132 435 133 436
rect 131 435 132 436
rect 130 435 131 436
rect 129 435 130 436
rect 128 435 129 436
rect 127 435 128 436
rect 126 435 127 436
rect 125 435 126 436
rect 124 435 125 436
rect 123 435 124 436
rect 122 435 123 436
rect 121 435 122 436
rect 120 435 121 436
rect 119 435 120 436
rect 118 435 119 436
rect 117 435 118 436
rect 82 435 83 436
rect 81 435 82 436
rect 80 435 81 436
rect 79 435 80 436
rect 78 435 79 436
rect 77 435 78 436
rect 76 435 77 436
rect 75 435 76 436
rect 74 435 75 436
rect 73 435 74 436
rect 72 435 73 436
rect 71 435 72 436
rect 70 435 71 436
rect 69 435 70 436
rect 68 435 69 436
rect 67 435 68 436
rect 60 435 61 436
rect 59 435 60 436
rect 58 435 59 436
rect 57 435 58 436
rect 56 435 57 436
rect 55 435 56 436
rect 54 435 55 436
rect 53 435 54 436
rect 52 435 53 436
rect 51 435 52 436
rect 50 435 51 436
rect 49 435 50 436
rect 48 435 49 436
rect 47 435 48 436
rect 46 435 47 436
rect 45 435 46 436
rect 44 435 45 436
rect 43 435 44 436
rect 42 435 43 436
rect 41 435 42 436
rect 40 435 41 436
rect 34 435 35 436
rect 33 435 34 436
rect 32 435 33 436
rect 31 435 32 436
rect 30 435 31 436
rect 29 435 30 436
rect 28 435 29 436
rect 27 435 28 436
rect 26 435 27 436
rect 25 435 26 436
rect 24 435 25 436
rect 23 435 24 436
rect 22 435 23 436
rect 21 435 22 436
rect 20 435 21 436
rect 19 435 20 436
rect 18 435 19 436
rect 17 435 18 436
rect 16 435 17 436
rect 15 435 16 436
rect 136 436 137 437
rect 135 436 136 437
rect 134 436 135 437
rect 82 436 83 437
rect 81 436 82 437
rect 80 436 81 437
rect 79 436 80 437
rect 78 436 79 437
rect 77 436 78 437
rect 76 436 77 437
rect 75 436 76 437
rect 74 436 75 437
rect 73 436 74 437
rect 72 436 73 437
rect 71 436 72 437
rect 70 436 71 437
rect 69 436 70 437
rect 68 436 69 437
rect 67 436 68 437
rect 60 436 61 437
rect 59 436 60 437
rect 58 436 59 437
rect 57 436 58 437
rect 56 436 57 437
rect 55 436 56 437
rect 54 436 55 437
rect 53 436 54 437
rect 52 436 53 437
rect 51 436 52 437
rect 50 436 51 437
rect 49 436 50 437
rect 48 436 49 437
rect 47 436 48 437
rect 46 436 47 437
rect 45 436 46 437
rect 44 436 45 437
rect 43 436 44 437
rect 42 436 43 437
rect 41 436 42 437
rect 40 436 41 437
rect 39 436 40 437
rect 38 436 39 437
rect 37 436 38 437
rect 36 436 37 437
rect 35 436 36 437
rect 34 436 35 437
rect 33 436 34 437
rect 32 436 33 437
rect 31 436 32 437
rect 30 436 31 437
rect 29 436 30 437
rect 28 436 29 437
rect 27 436 28 437
rect 26 436 27 437
rect 25 436 26 437
rect 24 436 25 437
rect 23 436 24 437
rect 22 436 23 437
rect 21 436 22 437
rect 20 436 21 437
rect 19 436 20 437
rect 18 436 19 437
rect 17 436 18 437
rect 16 436 17 437
rect 15 436 16 437
rect 137 437 138 438
rect 136 437 137 438
rect 135 437 136 438
rect 134 437 135 438
rect 133 437 134 438
rect 132 437 133 438
rect 82 437 83 438
rect 81 437 82 438
rect 80 437 81 438
rect 79 437 80 438
rect 78 437 79 438
rect 77 437 78 438
rect 76 437 77 438
rect 75 437 76 438
rect 74 437 75 438
rect 73 437 74 438
rect 72 437 73 438
rect 71 437 72 438
rect 70 437 71 438
rect 69 437 70 438
rect 68 437 69 438
rect 67 437 68 438
rect 59 437 60 438
rect 58 437 59 438
rect 57 437 58 438
rect 56 437 57 438
rect 55 437 56 438
rect 54 437 55 438
rect 53 437 54 438
rect 52 437 53 438
rect 51 437 52 438
rect 50 437 51 438
rect 49 437 50 438
rect 48 437 49 438
rect 47 437 48 438
rect 46 437 47 438
rect 45 437 46 438
rect 44 437 45 438
rect 43 437 44 438
rect 42 437 43 438
rect 41 437 42 438
rect 40 437 41 438
rect 39 437 40 438
rect 38 437 39 438
rect 37 437 38 438
rect 36 437 37 438
rect 35 437 36 438
rect 34 437 35 438
rect 33 437 34 438
rect 32 437 33 438
rect 31 437 32 438
rect 30 437 31 438
rect 29 437 30 438
rect 28 437 29 438
rect 27 437 28 438
rect 26 437 27 438
rect 25 437 26 438
rect 24 437 25 438
rect 23 437 24 438
rect 22 437 23 438
rect 21 437 22 438
rect 20 437 21 438
rect 19 437 20 438
rect 18 437 19 438
rect 17 437 18 438
rect 16 437 17 438
rect 15 437 16 438
rect 139 438 140 439
rect 138 438 139 439
rect 137 438 138 439
rect 136 438 137 439
rect 135 438 136 439
rect 134 438 135 439
rect 133 438 134 439
rect 132 438 133 439
rect 131 438 132 439
rect 82 438 83 439
rect 81 438 82 439
rect 80 438 81 439
rect 79 438 80 439
rect 78 438 79 439
rect 77 438 78 439
rect 76 438 77 439
rect 75 438 76 439
rect 74 438 75 439
rect 73 438 74 439
rect 72 438 73 439
rect 71 438 72 439
rect 70 438 71 439
rect 69 438 70 439
rect 68 438 69 439
rect 67 438 68 439
rect 58 438 59 439
rect 57 438 58 439
rect 56 438 57 439
rect 55 438 56 439
rect 54 438 55 439
rect 53 438 54 439
rect 52 438 53 439
rect 51 438 52 439
rect 50 438 51 439
rect 49 438 50 439
rect 48 438 49 439
rect 47 438 48 439
rect 46 438 47 439
rect 45 438 46 439
rect 44 438 45 439
rect 43 438 44 439
rect 42 438 43 439
rect 41 438 42 439
rect 40 438 41 439
rect 39 438 40 439
rect 38 438 39 439
rect 37 438 38 439
rect 36 438 37 439
rect 35 438 36 439
rect 34 438 35 439
rect 33 438 34 439
rect 32 438 33 439
rect 31 438 32 439
rect 30 438 31 439
rect 29 438 30 439
rect 28 438 29 439
rect 27 438 28 439
rect 26 438 27 439
rect 25 438 26 439
rect 24 438 25 439
rect 23 438 24 439
rect 22 438 23 439
rect 21 438 22 439
rect 20 438 21 439
rect 19 438 20 439
rect 18 438 19 439
rect 17 438 18 439
rect 16 438 17 439
rect 15 438 16 439
rect 140 439 141 440
rect 139 439 140 440
rect 138 439 139 440
rect 137 439 138 440
rect 136 439 137 440
rect 135 439 136 440
rect 134 439 135 440
rect 133 439 134 440
rect 132 439 133 440
rect 131 439 132 440
rect 130 439 131 440
rect 129 439 130 440
rect 82 439 83 440
rect 81 439 82 440
rect 80 439 81 440
rect 79 439 80 440
rect 78 439 79 440
rect 77 439 78 440
rect 76 439 77 440
rect 75 439 76 440
rect 74 439 75 440
rect 73 439 74 440
rect 72 439 73 440
rect 71 439 72 440
rect 70 439 71 440
rect 69 439 70 440
rect 68 439 69 440
rect 67 439 68 440
rect 57 439 58 440
rect 56 439 57 440
rect 55 439 56 440
rect 54 439 55 440
rect 53 439 54 440
rect 52 439 53 440
rect 51 439 52 440
rect 50 439 51 440
rect 49 439 50 440
rect 48 439 49 440
rect 47 439 48 440
rect 46 439 47 440
rect 45 439 46 440
rect 44 439 45 440
rect 43 439 44 440
rect 42 439 43 440
rect 41 439 42 440
rect 40 439 41 440
rect 39 439 40 440
rect 38 439 39 440
rect 37 439 38 440
rect 36 439 37 440
rect 35 439 36 440
rect 34 439 35 440
rect 33 439 34 440
rect 32 439 33 440
rect 31 439 32 440
rect 30 439 31 440
rect 29 439 30 440
rect 28 439 29 440
rect 27 439 28 440
rect 26 439 27 440
rect 25 439 26 440
rect 24 439 25 440
rect 23 439 24 440
rect 22 439 23 440
rect 21 439 22 440
rect 20 439 21 440
rect 19 439 20 440
rect 18 439 19 440
rect 17 439 18 440
rect 16 439 17 440
rect 142 440 143 441
rect 141 440 142 441
rect 140 440 141 441
rect 139 440 140 441
rect 138 440 139 441
rect 137 440 138 441
rect 136 440 137 441
rect 135 440 136 441
rect 134 440 135 441
rect 133 440 134 441
rect 132 440 133 441
rect 131 440 132 441
rect 130 440 131 441
rect 129 440 130 441
rect 128 440 129 441
rect 82 440 83 441
rect 81 440 82 441
rect 80 440 81 441
rect 79 440 80 441
rect 78 440 79 441
rect 77 440 78 441
rect 76 440 77 441
rect 75 440 76 441
rect 74 440 75 441
rect 73 440 74 441
rect 72 440 73 441
rect 71 440 72 441
rect 70 440 71 441
rect 69 440 70 441
rect 68 440 69 441
rect 67 440 68 441
rect 57 440 58 441
rect 56 440 57 441
rect 55 440 56 441
rect 54 440 55 441
rect 53 440 54 441
rect 52 440 53 441
rect 51 440 52 441
rect 50 440 51 441
rect 49 440 50 441
rect 48 440 49 441
rect 47 440 48 441
rect 46 440 47 441
rect 45 440 46 441
rect 44 440 45 441
rect 43 440 44 441
rect 42 440 43 441
rect 41 440 42 441
rect 40 440 41 441
rect 39 440 40 441
rect 38 440 39 441
rect 37 440 38 441
rect 36 440 37 441
rect 35 440 36 441
rect 34 440 35 441
rect 33 440 34 441
rect 32 440 33 441
rect 31 440 32 441
rect 30 440 31 441
rect 29 440 30 441
rect 28 440 29 441
rect 27 440 28 441
rect 26 440 27 441
rect 25 440 26 441
rect 24 440 25 441
rect 23 440 24 441
rect 22 440 23 441
rect 21 440 22 441
rect 20 440 21 441
rect 19 440 20 441
rect 18 440 19 441
rect 17 440 18 441
rect 16 440 17 441
rect 143 441 144 442
rect 142 441 143 442
rect 141 441 142 442
rect 140 441 141 442
rect 139 441 140 442
rect 138 441 139 442
rect 137 441 138 442
rect 136 441 137 442
rect 135 441 136 442
rect 134 441 135 442
rect 133 441 134 442
rect 132 441 133 442
rect 131 441 132 442
rect 130 441 131 442
rect 129 441 130 442
rect 128 441 129 442
rect 127 441 128 442
rect 126 441 127 442
rect 82 441 83 442
rect 81 441 82 442
rect 80 441 81 442
rect 79 441 80 442
rect 78 441 79 442
rect 77 441 78 442
rect 76 441 77 442
rect 75 441 76 442
rect 74 441 75 442
rect 73 441 74 442
rect 72 441 73 442
rect 71 441 72 442
rect 70 441 71 442
rect 69 441 70 442
rect 68 441 69 442
rect 67 441 68 442
rect 56 441 57 442
rect 55 441 56 442
rect 54 441 55 442
rect 53 441 54 442
rect 52 441 53 442
rect 51 441 52 442
rect 50 441 51 442
rect 49 441 50 442
rect 48 441 49 442
rect 47 441 48 442
rect 46 441 47 442
rect 45 441 46 442
rect 44 441 45 442
rect 43 441 44 442
rect 42 441 43 442
rect 41 441 42 442
rect 40 441 41 442
rect 39 441 40 442
rect 38 441 39 442
rect 37 441 38 442
rect 36 441 37 442
rect 35 441 36 442
rect 34 441 35 442
rect 33 441 34 442
rect 32 441 33 442
rect 31 441 32 442
rect 30 441 31 442
rect 29 441 30 442
rect 28 441 29 442
rect 27 441 28 442
rect 26 441 27 442
rect 25 441 26 442
rect 24 441 25 442
rect 23 441 24 442
rect 22 441 23 442
rect 21 441 22 442
rect 20 441 21 442
rect 19 441 20 442
rect 18 441 19 442
rect 17 441 18 442
rect 16 441 17 442
rect 144 442 145 443
rect 143 442 144 443
rect 142 442 143 443
rect 141 442 142 443
rect 140 442 141 443
rect 139 442 140 443
rect 138 442 139 443
rect 137 442 138 443
rect 136 442 137 443
rect 133 442 134 443
rect 132 442 133 443
rect 131 442 132 443
rect 130 442 131 443
rect 129 442 130 443
rect 128 442 129 443
rect 127 442 128 443
rect 126 442 127 443
rect 82 442 83 443
rect 81 442 82 443
rect 80 442 81 443
rect 79 442 80 443
rect 78 442 79 443
rect 77 442 78 443
rect 76 442 77 443
rect 75 442 76 443
rect 74 442 75 443
rect 73 442 74 443
rect 72 442 73 443
rect 71 442 72 443
rect 70 442 71 443
rect 69 442 70 443
rect 68 442 69 443
rect 67 442 68 443
rect 56 442 57 443
rect 55 442 56 443
rect 54 442 55 443
rect 53 442 54 443
rect 52 442 53 443
rect 51 442 52 443
rect 50 442 51 443
rect 49 442 50 443
rect 48 442 49 443
rect 47 442 48 443
rect 46 442 47 443
rect 45 442 46 443
rect 44 442 45 443
rect 43 442 44 443
rect 42 442 43 443
rect 41 442 42 443
rect 40 442 41 443
rect 39 442 40 443
rect 38 442 39 443
rect 37 442 38 443
rect 36 442 37 443
rect 35 442 36 443
rect 34 442 35 443
rect 33 442 34 443
rect 32 442 33 443
rect 31 442 32 443
rect 30 442 31 443
rect 29 442 30 443
rect 28 442 29 443
rect 27 442 28 443
rect 26 442 27 443
rect 25 442 26 443
rect 24 442 25 443
rect 23 442 24 443
rect 22 442 23 443
rect 21 442 22 443
rect 20 442 21 443
rect 19 442 20 443
rect 18 442 19 443
rect 17 442 18 443
rect 16 442 17 443
rect 144 443 145 444
rect 143 443 144 444
rect 142 443 143 444
rect 141 443 142 444
rect 140 443 141 444
rect 139 443 140 444
rect 138 443 139 444
rect 131 443 132 444
rect 130 443 131 444
rect 129 443 130 444
rect 128 443 129 444
rect 127 443 128 444
rect 126 443 127 444
rect 82 443 83 444
rect 81 443 82 444
rect 80 443 81 444
rect 79 443 80 444
rect 78 443 79 444
rect 77 443 78 444
rect 76 443 77 444
rect 75 443 76 444
rect 74 443 75 444
rect 73 443 74 444
rect 72 443 73 444
rect 71 443 72 444
rect 70 443 71 444
rect 69 443 70 444
rect 68 443 69 444
rect 67 443 68 444
rect 55 443 56 444
rect 54 443 55 444
rect 53 443 54 444
rect 52 443 53 444
rect 51 443 52 444
rect 50 443 51 444
rect 49 443 50 444
rect 48 443 49 444
rect 47 443 48 444
rect 46 443 47 444
rect 45 443 46 444
rect 44 443 45 444
rect 43 443 44 444
rect 42 443 43 444
rect 41 443 42 444
rect 40 443 41 444
rect 39 443 40 444
rect 38 443 39 444
rect 37 443 38 444
rect 36 443 37 444
rect 35 443 36 444
rect 34 443 35 444
rect 33 443 34 444
rect 32 443 33 444
rect 31 443 32 444
rect 30 443 31 444
rect 29 443 30 444
rect 28 443 29 444
rect 27 443 28 444
rect 26 443 27 444
rect 25 443 26 444
rect 24 443 25 444
rect 23 443 24 444
rect 22 443 23 444
rect 21 443 22 444
rect 20 443 21 444
rect 19 443 20 444
rect 18 443 19 444
rect 17 443 18 444
rect 144 444 145 445
rect 143 444 144 445
rect 142 444 143 445
rect 141 444 142 445
rect 140 444 141 445
rect 139 444 140 445
rect 130 444 131 445
rect 129 444 130 445
rect 128 444 129 445
rect 127 444 128 445
rect 126 444 127 445
rect 82 444 83 445
rect 81 444 82 445
rect 80 444 81 445
rect 79 444 80 445
rect 78 444 79 445
rect 77 444 78 445
rect 76 444 77 445
rect 75 444 76 445
rect 74 444 75 445
rect 73 444 74 445
rect 72 444 73 445
rect 71 444 72 445
rect 70 444 71 445
rect 69 444 70 445
rect 68 444 69 445
rect 67 444 68 445
rect 54 444 55 445
rect 53 444 54 445
rect 52 444 53 445
rect 51 444 52 445
rect 50 444 51 445
rect 49 444 50 445
rect 48 444 49 445
rect 47 444 48 445
rect 46 444 47 445
rect 45 444 46 445
rect 44 444 45 445
rect 43 444 44 445
rect 42 444 43 445
rect 41 444 42 445
rect 40 444 41 445
rect 39 444 40 445
rect 38 444 39 445
rect 37 444 38 445
rect 36 444 37 445
rect 35 444 36 445
rect 34 444 35 445
rect 33 444 34 445
rect 32 444 33 445
rect 31 444 32 445
rect 30 444 31 445
rect 29 444 30 445
rect 28 444 29 445
rect 27 444 28 445
rect 26 444 27 445
rect 25 444 26 445
rect 24 444 25 445
rect 23 444 24 445
rect 22 444 23 445
rect 21 444 22 445
rect 20 444 21 445
rect 19 444 20 445
rect 18 444 19 445
rect 17 444 18 445
rect 144 445 145 446
rect 143 445 144 446
rect 142 445 143 446
rect 141 445 142 446
rect 140 445 141 446
rect 129 445 130 446
rect 128 445 129 446
rect 127 445 128 446
rect 126 445 127 446
rect 82 445 83 446
rect 81 445 82 446
rect 80 445 81 446
rect 79 445 80 446
rect 78 445 79 446
rect 77 445 78 446
rect 76 445 77 446
rect 75 445 76 446
rect 74 445 75 446
rect 73 445 74 446
rect 72 445 73 446
rect 71 445 72 446
rect 70 445 71 446
rect 69 445 70 446
rect 68 445 69 446
rect 67 445 68 446
rect 53 445 54 446
rect 52 445 53 446
rect 51 445 52 446
rect 50 445 51 446
rect 49 445 50 446
rect 48 445 49 446
rect 47 445 48 446
rect 46 445 47 446
rect 45 445 46 446
rect 44 445 45 446
rect 43 445 44 446
rect 42 445 43 446
rect 41 445 42 446
rect 40 445 41 446
rect 39 445 40 446
rect 38 445 39 446
rect 37 445 38 446
rect 36 445 37 446
rect 35 445 36 446
rect 34 445 35 446
rect 33 445 34 446
rect 32 445 33 446
rect 31 445 32 446
rect 30 445 31 446
rect 29 445 30 446
rect 28 445 29 446
rect 27 445 28 446
rect 26 445 27 446
rect 25 445 26 446
rect 24 445 25 446
rect 23 445 24 446
rect 22 445 23 446
rect 21 445 22 446
rect 20 445 21 446
rect 19 445 20 446
rect 18 445 19 446
rect 144 446 145 447
rect 143 446 144 447
rect 142 446 143 447
rect 127 446 128 447
rect 126 446 127 447
rect 82 446 83 447
rect 81 446 82 447
rect 80 446 81 447
rect 79 446 80 447
rect 78 446 79 447
rect 77 446 78 447
rect 76 446 77 447
rect 75 446 76 447
rect 74 446 75 447
rect 73 446 74 447
rect 72 446 73 447
rect 71 446 72 447
rect 70 446 71 447
rect 69 446 70 447
rect 68 446 69 447
rect 67 446 68 447
rect 53 446 54 447
rect 52 446 53 447
rect 51 446 52 447
rect 50 446 51 447
rect 49 446 50 447
rect 48 446 49 447
rect 47 446 48 447
rect 46 446 47 447
rect 45 446 46 447
rect 44 446 45 447
rect 43 446 44 447
rect 42 446 43 447
rect 41 446 42 447
rect 40 446 41 447
rect 39 446 40 447
rect 38 446 39 447
rect 37 446 38 447
rect 36 446 37 447
rect 35 446 36 447
rect 34 446 35 447
rect 33 446 34 447
rect 32 446 33 447
rect 31 446 32 447
rect 30 446 31 447
rect 29 446 30 447
rect 28 446 29 447
rect 27 446 28 447
rect 26 446 27 447
rect 25 446 26 447
rect 24 446 25 447
rect 23 446 24 447
rect 22 446 23 447
rect 21 446 22 447
rect 20 446 21 447
rect 19 446 20 447
rect 18 446 19 447
rect 144 447 145 448
rect 143 447 144 448
rect 126 447 127 448
rect 82 447 83 448
rect 81 447 82 448
rect 80 447 81 448
rect 79 447 80 448
rect 78 447 79 448
rect 77 447 78 448
rect 76 447 77 448
rect 75 447 76 448
rect 74 447 75 448
rect 73 447 74 448
rect 72 447 73 448
rect 71 447 72 448
rect 70 447 71 448
rect 69 447 70 448
rect 68 447 69 448
rect 67 447 68 448
rect 52 447 53 448
rect 51 447 52 448
rect 50 447 51 448
rect 49 447 50 448
rect 48 447 49 448
rect 47 447 48 448
rect 46 447 47 448
rect 45 447 46 448
rect 44 447 45 448
rect 43 447 44 448
rect 42 447 43 448
rect 41 447 42 448
rect 40 447 41 448
rect 39 447 40 448
rect 38 447 39 448
rect 37 447 38 448
rect 36 447 37 448
rect 35 447 36 448
rect 34 447 35 448
rect 33 447 34 448
rect 32 447 33 448
rect 31 447 32 448
rect 30 447 31 448
rect 29 447 30 448
rect 28 447 29 448
rect 27 447 28 448
rect 26 447 27 448
rect 25 447 26 448
rect 24 447 25 448
rect 23 447 24 448
rect 22 447 23 448
rect 21 447 22 448
rect 20 447 21 448
rect 19 447 20 448
rect 82 448 83 449
rect 81 448 82 449
rect 80 448 81 449
rect 79 448 80 449
rect 78 448 79 449
rect 77 448 78 449
rect 76 448 77 449
rect 75 448 76 449
rect 74 448 75 449
rect 73 448 74 449
rect 72 448 73 449
rect 71 448 72 449
rect 70 448 71 449
rect 69 448 70 449
rect 68 448 69 449
rect 67 448 68 449
rect 51 448 52 449
rect 50 448 51 449
rect 49 448 50 449
rect 48 448 49 449
rect 47 448 48 449
rect 46 448 47 449
rect 45 448 46 449
rect 44 448 45 449
rect 43 448 44 449
rect 42 448 43 449
rect 41 448 42 449
rect 40 448 41 449
rect 39 448 40 449
rect 38 448 39 449
rect 37 448 38 449
rect 36 448 37 449
rect 35 448 36 449
rect 34 448 35 449
rect 33 448 34 449
rect 32 448 33 449
rect 31 448 32 449
rect 30 448 31 449
rect 29 448 30 449
rect 28 448 29 449
rect 27 448 28 449
rect 26 448 27 449
rect 25 448 26 449
rect 24 448 25 449
rect 23 448 24 449
rect 22 448 23 449
rect 21 448 22 449
rect 20 448 21 449
rect 19 448 20 449
rect 82 449 83 450
rect 81 449 82 450
rect 80 449 81 450
rect 79 449 80 450
rect 78 449 79 450
rect 77 449 78 450
rect 76 449 77 450
rect 75 449 76 450
rect 74 449 75 450
rect 73 449 74 450
rect 72 449 73 450
rect 71 449 72 450
rect 70 449 71 450
rect 69 449 70 450
rect 68 449 69 450
rect 67 449 68 450
rect 50 449 51 450
rect 49 449 50 450
rect 48 449 49 450
rect 47 449 48 450
rect 46 449 47 450
rect 45 449 46 450
rect 44 449 45 450
rect 43 449 44 450
rect 42 449 43 450
rect 41 449 42 450
rect 40 449 41 450
rect 39 449 40 450
rect 38 449 39 450
rect 37 449 38 450
rect 36 449 37 450
rect 35 449 36 450
rect 34 449 35 450
rect 33 449 34 450
rect 32 449 33 450
rect 31 449 32 450
rect 30 449 31 450
rect 29 449 30 450
rect 28 449 29 450
rect 27 449 28 450
rect 26 449 27 450
rect 25 449 26 450
rect 24 449 25 450
rect 23 449 24 450
rect 22 449 23 450
rect 21 449 22 450
rect 20 449 21 450
rect 82 450 83 451
rect 81 450 82 451
rect 80 450 81 451
rect 79 450 80 451
rect 78 450 79 451
rect 77 450 78 451
rect 76 450 77 451
rect 75 450 76 451
rect 74 450 75 451
rect 73 450 74 451
rect 72 450 73 451
rect 71 450 72 451
rect 70 450 71 451
rect 69 450 70 451
rect 68 450 69 451
rect 67 450 68 451
rect 49 450 50 451
rect 48 450 49 451
rect 47 450 48 451
rect 46 450 47 451
rect 45 450 46 451
rect 44 450 45 451
rect 43 450 44 451
rect 42 450 43 451
rect 41 450 42 451
rect 40 450 41 451
rect 39 450 40 451
rect 38 450 39 451
rect 37 450 38 451
rect 36 450 37 451
rect 35 450 36 451
rect 34 450 35 451
rect 33 450 34 451
rect 32 450 33 451
rect 31 450 32 451
rect 30 450 31 451
rect 29 450 30 451
rect 28 450 29 451
rect 27 450 28 451
rect 26 450 27 451
rect 25 450 26 451
rect 24 450 25 451
rect 23 450 24 451
rect 22 450 23 451
rect 21 450 22 451
rect 82 451 83 452
rect 81 451 82 452
rect 80 451 81 452
rect 79 451 80 452
rect 78 451 79 452
rect 77 451 78 452
rect 76 451 77 452
rect 75 451 76 452
rect 74 451 75 452
rect 73 451 74 452
rect 72 451 73 452
rect 71 451 72 452
rect 70 451 71 452
rect 69 451 70 452
rect 68 451 69 452
rect 67 451 68 452
rect 48 451 49 452
rect 47 451 48 452
rect 46 451 47 452
rect 45 451 46 452
rect 44 451 45 452
rect 43 451 44 452
rect 42 451 43 452
rect 41 451 42 452
rect 40 451 41 452
rect 39 451 40 452
rect 38 451 39 452
rect 37 451 38 452
rect 36 451 37 452
rect 35 451 36 452
rect 34 451 35 452
rect 33 451 34 452
rect 32 451 33 452
rect 31 451 32 452
rect 30 451 31 452
rect 29 451 30 452
rect 28 451 29 452
rect 27 451 28 452
rect 26 451 27 452
rect 25 451 26 452
rect 24 451 25 452
rect 23 451 24 452
rect 22 451 23 452
rect 82 452 83 453
rect 81 452 82 453
rect 80 452 81 453
rect 79 452 80 453
rect 78 452 79 453
rect 77 452 78 453
rect 76 452 77 453
rect 75 452 76 453
rect 74 452 75 453
rect 73 452 74 453
rect 72 452 73 453
rect 71 452 72 453
rect 70 452 71 453
rect 69 452 70 453
rect 68 452 69 453
rect 67 452 68 453
rect 46 452 47 453
rect 45 452 46 453
rect 44 452 45 453
rect 43 452 44 453
rect 42 452 43 453
rect 41 452 42 453
rect 40 452 41 453
rect 39 452 40 453
rect 38 452 39 453
rect 37 452 38 453
rect 36 452 37 453
rect 35 452 36 453
rect 34 452 35 453
rect 33 452 34 453
rect 32 452 33 453
rect 31 452 32 453
rect 30 452 31 453
rect 29 452 30 453
rect 28 452 29 453
rect 27 452 28 453
rect 26 452 27 453
rect 25 452 26 453
rect 24 452 25 453
rect 23 452 24 453
rect 82 453 83 454
rect 81 453 82 454
rect 80 453 81 454
rect 79 453 80 454
rect 78 453 79 454
rect 77 453 78 454
rect 76 453 77 454
rect 75 453 76 454
rect 74 453 75 454
rect 73 453 74 454
rect 72 453 73 454
rect 71 453 72 454
rect 70 453 71 454
rect 69 453 70 454
rect 68 453 69 454
rect 67 453 68 454
rect 44 453 45 454
rect 43 453 44 454
rect 42 453 43 454
rect 41 453 42 454
rect 40 453 41 454
rect 39 453 40 454
rect 38 453 39 454
rect 37 453 38 454
rect 36 453 37 454
rect 35 453 36 454
rect 34 453 35 454
rect 33 453 34 454
rect 32 453 33 454
rect 31 453 32 454
rect 30 453 31 454
rect 29 453 30 454
rect 28 453 29 454
rect 27 453 28 454
rect 26 453 27 454
rect 25 453 26 454
rect 82 454 83 455
rect 81 454 82 455
rect 80 454 81 455
rect 79 454 80 455
rect 78 454 79 455
rect 77 454 78 455
rect 76 454 77 455
rect 75 454 76 455
rect 74 454 75 455
rect 73 454 74 455
rect 72 454 73 455
rect 71 454 72 455
rect 70 454 71 455
rect 69 454 70 455
rect 68 454 69 455
rect 67 454 68 455
rect 42 454 43 455
rect 41 454 42 455
rect 40 454 41 455
rect 39 454 40 455
rect 38 454 39 455
rect 37 454 38 455
rect 36 454 37 455
rect 35 454 36 455
rect 34 454 35 455
rect 33 454 34 455
rect 32 454 33 455
rect 31 454 32 455
rect 30 454 31 455
rect 29 454 30 455
rect 28 454 29 455
rect 27 454 28 455
rect 82 455 83 456
rect 81 455 82 456
rect 80 455 81 456
rect 79 455 80 456
rect 78 455 79 456
rect 77 455 78 456
rect 76 455 77 456
rect 75 455 76 456
rect 74 455 75 456
rect 73 455 74 456
rect 72 455 73 456
rect 71 455 72 456
rect 70 455 71 456
rect 69 455 70 456
rect 68 455 69 456
rect 67 455 68 456
rect 37 455 38 456
rect 36 455 37 456
rect 35 455 36 456
rect 34 455 35 456
rect 33 455 34 456
rect 32 455 33 456
<< metal3 >>
rect 59 16 60 17
rect 58 16 59 17
rect 57 16 58 17
rect 56 16 57 17
rect 55 16 56 17
rect 54 16 55 17
rect 53 16 54 17
rect 52 16 53 17
rect 51 16 52 17
rect 50 16 51 17
rect 49 16 50 17
rect 48 16 49 17
rect 47 16 48 17
rect 46 16 47 17
rect 63 17 64 18
rect 62 17 63 18
rect 61 17 62 18
rect 60 17 61 18
rect 59 17 60 18
rect 58 17 59 18
rect 57 17 58 18
rect 56 17 57 18
rect 55 17 56 18
rect 54 17 55 18
rect 53 17 54 18
rect 52 17 53 18
rect 51 17 52 18
rect 50 17 51 18
rect 49 17 50 18
rect 48 17 49 18
rect 47 17 48 18
rect 46 17 47 18
rect 45 17 46 18
rect 44 17 45 18
rect 43 17 44 18
rect 42 17 43 18
rect 41 17 42 18
rect 66 18 67 19
rect 65 18 66 19
rect 64 18 65 19
rect 63 18 64 19
rect 62 18 63 19
rect 61 18 62 19
rect 60 18 61 19
rect 59 18 60 19
rect 58 18 59 19
rect 57 18 58 19
rect 56 18 57 19
rect 55 18 56 19
rect 54 18 55 19
rect 53 18 54 19
rect 52 18 53 19
rect 51 18 52 19
rect 50 18 51 19
rect 49 18 50 19
rect 48 18 49 19
rect 47 18 48 19
rect 46 18 47 19
rect 45 18 46 19
rect 44 18 45 19
rect 43 18 44 19
rect 42 18 43 19
rect 41 18 42 19
rect 40 18 41 19
rect 39 18 40 19
rect 38 18 39 19
rect 68 19 69 20
rect 67 19 68 20
rect 66 19 67 20
rect 65 19 66 20
rect 64 19 65 20
rect 63 19 64 20
rect 62 19 63 20
rect 61 19 62 20
rect 60 19 61 20
rect 59 19 60 20
rect 58 19 59 20
rect 57 19 58 20
rect 56 19 57 20
rect 55 19 56 20
rect 54 19 55 20
rect 53 19 54 20
rect 52 19 53 20
rect 51 19 52 20
rect 50 19 51 20
rect 49 19 50 20
rect 48 19 49 20
rect 47 19 48 20
rect 46 19 47 20
rect 45 19 46 20
rect 44 19 45 20
rect 43 19 44 20
rect 42 19 43 20
rect 41 19 42 20
rect 40 19 41 20
rect 39 19 40 20
rect 38 19 39 20
rect 37 19 38 20
rect 36 19 37 20
rect 70 20 71 21
rect 69 20 70 21
rect 68 20 69 21
rect 67 20 68 21
rect 66 20 67 21
rect 65 20 66 21
rect 64 20 65 21
rect 63 20 64 21
rect 62 20 63 21
rect 61 20 62 21
rect 60 20 61 21
rect 59 20 60 21
rect 58 20 59 21
rect 57 20 58 21
rect 56 20 57 21
rect 55 20 56 21
rect 54 20 55 21
rect 53 20 54 21
rect 52 20 53 21
rect 51 20 52 21
rect 50 20 51 21
rect 49 20 50 21
rect 48 20 49 21
rect 47 20 48 21
rect 46 20 47 21
rect 45 20 46 21
rect 44 20 45 21
rect 43 20 44 21
rect 42 20 43 21
rect 41 20 42 21
rect 40 20 41 21
rect 39 20 40 21
rect 38 20 39 21
rect 37 20 38 21
rect 36 20 37 21
rect 35 20 36 21
rect 34 20 35 21
rect 72 21 73 22
rect 71 21 72 22
rect 70 21 71 22
rect 69 21 70 22
rect 68 21 69 22
rect 67 21 68 22
rect 66 21 67 22
rect 65 21 66 22
rect 64 21 65 22
rect 63 21 64 22
rect 62 21 63 22
rect 61 21 62 22
rect 60 21 61 22
rect 59 21 60 22
rect 58 21 59 22
rect 57 21 58 22
rect 56 21 57 22
rect 55 21 56 22
rect 54 21 55 22
rect 53 21 54 22
rect 52 21 53 22
rect 51 21 52 22
rect 50 21 51 22
rect 49 21 50 22
rect 48 21 49 22
rect 47 21 48 22
rect 46 21 47 22
rect 45 21 46 22
rect 44 21 45 22
rect 43 21 44 22
rect 42 21 43 22
rect 41 21 42 22
rect 40 21 41 22
rect 39 21 40 22
rect 38 21 39 22
rect 37 21 38 22
rect 36 21 37 22
rect 35 21 36 22
rect 34 21 35 22
rect 33 21 34 22
rect 73 22 74 23
rect 72 22 73 23
rect 71 22 72 23
rect 70 22 71 23
rect 69 22 70 23
rect 68 22 69 23
rect 67 22 68 23
rect 66 22 67 23
rect 65 22 66 23
rect 64 22 65 23
rect 63 22 64 23
rect 62 22 63 23
rect 61 22 62 23
rect 60 22 61 23
rect 59 22 60 23
rect 58 22 59 23
rect 57 22 58 23
rect 56 22 57 23
rect 55 22 56 23
rect 54 22 55 23
rect 53 22 54 23
rect 52 22 53 23
rect 51 22 52 23
rect 50 22 51 23
rect 49 22 50 23
rect 48 22 49 23
rect 47 22 48 23
rect 46 22 47 23
rect 45 22 46 23
rect 44 22 45 23
rect 43 22 44 23
rect 42 22 43 23
rect 41 22 42 23
rect 40 22 41 23
rect 39 22 40 23
rect 38 22 39 23
rect 37 22 38 23
rect 36 22 37 23
rect 35 22 36 23
rect 34 22 35 23
rect 33 22 34 23
rect 32 22 33 23
rect 31 22 32 23
rect 74 23 75 24
rect 73 23 74 24
rect 72 23 73 24
rect 71 23 72 24
rect 70 23 71 24
rect 69 23 70 24
rect 68 23 69 24
rect 67 23 68 24
rect 66 23 67 24
rect 65 23 66 24
rect 64 23 65 24
rect 63 23 64 24
rect 62 23 63 24
rect 61 23 62 24
rect 60 23 61 24
rect 59 23 60 24
rect 58 23 59 24
rect 57 23 58 24
rect 56 23 57 24
rect 55 23 56 24
rect 54 23 55 24
rect 53 23 54 24
rect 52 23 53 24
rect 51 23 52 24
rect 50 23 51 24
rect 49 23 50 24
rect 48 23 49 24
rect 47 23 48 24
rect 46 23 47 24
rect 45 23 46 24
rect 44 23 45 24
rect 43 23 44 24
rect 42 23 43 24
rect 41 23 42 24
rect 40 23 41 24
rect 39 23 40 24
rect 38 23 39 24
rect 37 23 38 24
rect 36 23 37 24
rect 35 23 36 24
rect 34 23 35 24
rect 33 23 34 24
rect 32 23 33 24
rect 31 23 32 24
rect 30 23 31 24
rect 75 24 76 25
rect 74 24 75 25
rect 73 24 74 25
rect 72 24 73 25
rect 71 24 72 25
rect 70 24 71 25
rect 69 24 70 25
rect 68 24 69 25
rect 67 24 68 25
rect 66 24 67 25
rect 65 24 66 25
rect 64 24 65 25
rect 63 24 64 25
rect 62 24 63 25
rect 61 24 62 25
rect 60 24 61 25
rect 59 24 60 25
rect 58 24 59 25
rect 57 24 58 25
rect 56 24 57 25
rect 55 24 56 25
rect 54 24 55 25
rect 53 24 54 25
rect 52 24 53 25
rect 51 24 52 25
rect 50 24 51 25
rect 49 24 50 25
rect 48 24 49 25
rect 47 24 48 25
rect 46 24 47 25
rect 45 24 46 25
rect 44 24 45 25
rect 43 24 44 25
rect 42 24 43 25
rect 41 24 42 25
rect 40 24 41 25
rect 39 24 40 25
rect 38 24 39 25
rect 37 24 38 25
rect 36 24 37 25
rect 35 24 36 25
rect 34 24 35 25
rect 33 24 34 25
rect 32 24 33 25
rect 31 24 32 25
rect 30 24 31 25
rect 29 24 30 25
rect 76 25 77 26
rect 75 25 76 26
rect 74 25 75 26
rect 73 25 74 26
rect 72 25 73 26
rect 71 25 72 26
rect 70 25 71 26
rect 69 25 70 26
rect 68 25 69 26
rect 67 25 68 26
rect 66 25 67 26
rect 65 25 66 26
rect 64 25 65 26
rect 63 25 64 26
rect 62 25 63 26
rect 61 25 62 26
rect 60 25 61 26
rect 59 25 60 26
rect 58 25 59 26
rect 57 25 58 26
rect 56 25 57 26
rect 55 25 56 26
rect 54 25 55 26
rect 53 25 54 26
rect 52 25 53 26
rect 51 25 52 26
rect 50 25 51 26
rect 49 25 50 26
rect 48 25 49 26
rect 47 25 48 26
rect 46 25 47 26
rect 45 25 46 26
rect 44 25 45 26
rect 43 25 44 26
rect 42 25 43 26
rect 41 25 42 26
rect 40 25 41 26
rect 39 25 40 26
rect 38 25 39 26
rect 37 25 38 26
rect 36 25 37 26
rect 35 25 36 26
rect 34 25 35 26
rect 33 25 34 26
rect 32 25 33 26
rect 31 25 32 26
rect 30 25 31 26
rect 29 25 30 26
rect 28 25 29 26
rect 27 25 28 26
rect 77 26 78 27
rect 76 26 77 27
rect 75 26 76 27
rect 74 26 75 27
rect 73 26 74 27
rect 72 26 73 27
rect 71 26 72 27
rect 70 26 71 27
rect 69 26 70 27
rect 68 26 69 27
rect 67 26 68 27
rect 66 26 67 27
rect 65 26 66 27
rect 64 26 65 27
rect 63 26 64 27
rect 62 26 63 27
rect 61 26 62 27
rect 60 26 61 27
rect 59 26 60 27
rect 58 26 59 27
rect 57 26 58 27
rect 56 26 57 27
rect 55 26 56 27
rect 54 26 55 27
rect 53 26 54 27
rect 52 26 53 27
rect 51 26 52 27
rect 50 26 51 27
rect 49 26 50 27
rect 48 26 49 27
rect 47 26 48 27
rect 46 26 47 27
rect 45 26 46 27
rect 44 26 45 27
rect 43 26 44 27
rect 42 26 43 27
rect 41 26 42 27
rect 40 26 41 27
rect 39 26 40 27
rect 38 26 39 27
rect 37 26 38 27
rect 36 26 37 27
rect 35 26 36 27
rect 34 26 35 27
rect 33 26 34 27
rect 32 26 33 27
rect 31 26 32 27
rect 30 26 31 27
rect 29 26 30 27
rect 28 26 29 27
rect 27 26 28 27
rect 26 26 27 27
rect 78 27 79 28
rect 77 27 78 28
rect 76 27 77 28
rect 75 27 76 28
rect 74 27 75 28
rect 73 27 74 28
rect 72 27 73 28
rect 71 27 72 28
rect 70 27 71 28
rect 69 27 70 28
rect 68 27 69 28
rect 67 27 68 28
rect 66 27 67 28
rect 65 27 66 28
rect 64 27 65 28
rect 63 27 64 28
rect 62 27 63 28
rect 61 27 62 28
rect 60 27 61 28
rect 59 27 60 28
rect 58 27 59 28
rect 57 27 58 28
rect 56 27 57 28
rect 55 27 56 28
rect 54 27 55 28
rect 53 27 54 28
rect 52 27 53 28
rect 51 27 52 28
rect 50 27 51 28
rect 49 27 50 28
rect 48 27 49 28
rect 47 27 48 28
rect 46 27 47 28
rect 45 27 46 28
rect 44 27 45 28
rect 43 27 44 28
rect 42 27 43 28
rect 41 27 42 28
rect 40 27 41 28
rect 39 27 40 28
rect 38 27 39 28
rect 37 27 38 28
rect 36 27 37 28
rect 35 27 36 28
rect 34 27 35 28
rect 33 27 34 28
rect 32 27 33 28
rect 31 27 32 28
rect 30 27 31 28
rect 29 27 30 28
rect 28 27 29 28
rect 27 27 28 28
rect 26 27 27 28
rect 79 28 80 29
rect 78 28 79 29
rect 77 28 78 29
rect 76 28 77 29
rect 75 28 76 29
rect 74 28 75 29
rect 73 28 74 29
rect 72 28 73 29
rect 71 28 72 29
rect 70 28 71 29
rect 69 28 70 29
rect 68 28 69 29
rect 67 28 68 29
rect 66 28 67 29
rect 65 28 66 29
rect 64 28 65 29
rect 63 28 64 29
rect 62 28 63 29
rect 61 28 62 29
rect 60 28 61 29
rect 59 28 60 29
rect 58 28 59 29
rect 57 28 58 29
rect 56 28 57 29
rect 55 28 56 29
rect 54 28 55 29
rect 53 28 54 29
rect 52 28 53 29
rect 51 28 52 29
rect 50 28 51 29
rect 49 28 50 29
rect 48 28 49 29
rect 47 28 48 29
rect 46 28 47 29
rect 45 28 46 29
rect 44 28 45 29
rect 43 28 44 29
rect 42 28 43 29
rect 41 28 42 29
rect 40 28 41 29
rect 39 28 40 29
rect 38 28 39 29
rect 37 28 38 29
rect 36 28 37 29
rect 35 28 36 29
rect 34 28 35 29
rect 33 28 34 29
rect 32 28 33 29
rect 31 28 32 29
rect 30 28 31 29
rect 29 28 30 29
rect 28 28 29 29
rect 27 28 28 29
rect 26 28 27 29
rect 25 28 26 29
rect 80 29 81 30
rect 79 29 80 30
rect 78 29 79 30
rect 77 29 78 30
rect 76 29 77 30
rect 75 29 76 30
rect 74 29 75 30
rect 73 29 74 30
rect 72 29 73 30
rect 71 29 72 30
rect 70 29 71 30
rect 69 29 70 30
rect 68 29 69 30
rect 67 29 68 30
rect 66 29 67 30
rect 65 29 66 30
rect 64 29 65 30
rect 63 29 64 30
rect 62 29 63 30
rect 61 29 62 30
rect 60 29 61 30
rect 59 29 60 30
rect 58 29 59 30
rect 57 29 58 30
rect 56 29 57 30
rect 55 29 56 30
rect 54 29 55 30
rect 53 29 54 30
rect 52 29 53 30
rect 51 29 52 30
rect 50 29 51 30
rect 49 29 50 30
rect 48 29 49 30
rect 47 29 48 30
rect 46 29 47 30
rect 45 29 46 30
rect 44 29 45 30
rect 43 29 44 30
rect 42 29 43 30
rect 41 29 42 30
rect 40 29 41 30
rect 39 29 40 30
rect 38 29 39 30
rect 37 29 38 30
rect 36 29 37 30
rect 35 29 36 30
rect 34 29 35 30
rect 33 29 34 30
rect 32 29 33 30
rect 31 29 32 30
rect 30 29 31 30
rect 29 29 30 30
rect 28 29 29 30
rect 27 29 28 30
rect 26 29 27 30
rect 25 29 26 30
rect 24 29 25 30
rect 80 30 81 31
rect 79 30 80 31
rect 78 30 79 31
rect 77 30 78 31
rect 76 30 77 31
rect 75 30 76 31
rect 74 30 75 31
rect 73 30 74 31
rect 72 30 73 31
rect 71 30 72 31
rect 70 30 71 31
rect 69 30 70 31
rect 68 30 69 31
rect 67 30 68 31
rect 66 30 67 31
rect 65 30 66 31
rect 64 30 65 31
rect 63 30 64 31
rect 62 30 63 31
rect 61 30 62 31
rect 60 30 61 31
rect 59 30 60 31
rect 58 30 59 31
rect 57 30 58 31
rect 56 30 57 31
rect 55 30 56 31
rect 54 30 55 31
rect 53 30 54 31
rect 52 30 53 31
rect 51 30 52 31
rect 50 30 51 31
rect 49 30 50 31
rect 48 30 49 31
rect 47 30 48 31
rect 46 30 47 31
rect 45 30 46 31
rect 44 30 45 31
rect 43 30 44 31
rect 42 30 43 31
rect 41 30 42 31
rect 40 30 41 31
rect 39 30 40 31
rect 38 30 39 31
rect 37 30 38 31
rect 36 30 37 31
rect 35 30 36 31
rect 34 30 35 31
rect 33 30 34 31
rect 32 30 33 31
rect 31 30 32 31
rect 30 30 31 31
rect 29 30 30 31
rect 28 30 29 31
rect 27 30 28 31
rect 26 30 27 31
rect 25 30 26 31
rect 24 30 25 31
rect 23 30 24 31
rect 81 31 82 32
rect 80 31 81 32
rect 79 31 80 32
rect 78 31 79 32
rect 77 31 78 32
rect 76 31 77 32
rect 75 31 76 32
rect 74 31 75 32
rect 73 31 74 32
rect 72 31 73 32
rect 71 31 72 32
rect 70 31 71 32
rect 69 31 70 32
rect 68 31 69 32
rect 67 31 68 32
rect 66 31 67 32
rect 65 31 66 32
rect 64 31 65 32
rect 63 31 64 32
rect 62 31 63 32
rect 61 31 62 32
rect 60 31 61 32
rect 59 31 60 32
rect 58 31 59 32
rect 57 31 58 32
rect 56 31 57 32
rect 55 31 56 32
rect 54 31 55 32
rect 53 31 54 32
rect 52 31 53 32
rect 51 31 52 32
rect 50 31 51 32
rect 49 31 50 32
rect 48 31 49 32
rect 47 31 48 32
rect 46 31 47 32
rect 45 31 46 32
rect 44 31 45 32
rect 43 31 44 32
rect 42 31 43 32
rect 41 31 42 32
rect 40 31 41 32
rect 39 31 40 32
rect 38 31 39 32
rect 37 31 38 32
rect 36 31 37 32
rect 35 31 36 32
rect 34 31 35 32
rect 33 31 34 32
rect 32 31 33 32
rect 31 31 32 32
rect 30 31 31 32
rect 29 31 30 32
rect 28 31 29 32
rect 27 31 28 32
rect 26 31 27 32
rect 25 31 26 32
rect 24 31 25 32
rect 23 31 24 32
rect 81 32 82 33
rect 80 32 81 33
rect 79 32 80 33
rect 78 32 79 33
rect 77 32 78 33
rect 76 32 77 33
rect 75 32 76 33
rect 74 32 75 33
rect 73 32 74 33
rect 72 32 73 33
rect 71 32 72 33
rect 70 32 71 33
rect 69 32 70 33
rect 68 32 69 33
rect 67 32 68 33
rect 66 32 67 33
rect 65 32 66 33
rect 64 32 65 33
rect 63 32 64 33
rect 62 32 63 33
rect 61 32 62 33
rect 60 32 61 33
rect 59 32 60 33
rect 58 32 59 33
rect 57 32 58 33
rect 56 32 57 33
rect 55 32 56 33
rect 54 32 55 33
rect 53 32 54 33
rect 52 32 53 33
rect 51 32 52 33
rect 50 32 51 33
rect 49 32 50 33
rect 48 32 49 33
rect 47 32 48 33
rect 46 32 47 33
rect 45 32 46 33
rect 44 32 45 33
rect 43 32 44 33
rect 42 32 43 33
rect 41 32 42 33
rect 40 32 41 33
rect 39 32 40 33
rect 38 32 39 33
rect 37 32 38 33
rect 36 32 37 33
rect 35 32 36 33
rect 34 32 35 33
rect 33 32 34 33
rect 32 32 33 33
rect 31 32 32 33
rect 30 32 31 33
rect 29 32 30 33
rect 28 32 29 33
rect 27 32 28 33
rect 26 32 27 33
rect 25 32 26 33
rect 24 32 25 33
rect 23 32 24 33
rect 22 32 23 33
rect 82 33 83 34
rect 81 33 82 34
rect 80 33 81 34
rect 79 33 80 34
rect 78 33 79 34
rect 77 33 78 34
rect 76 33 77 34
rect 75 33 76 34
rect 74 33 75 34
rect 73 33 74 34
rect 72 33 73 34
rect 71 33 72 34
rect 70 33 71 34
rect 69 33 70 34
rect 68 33 69 34
rect 67 33 68 34
rect 66 33 67 34
rect 65 33 66 34
rect 64 33 65 34
rect 63 33 64 34
rect 62 33 63 34
rect 61 33 62 34
rect 60 33 61 34
rect 59 33 60 34
rect 58 33 59 34
rect 57 33 58 34
rect 56 33 57 34
rect 55 33 56 34
rect 54 33 55 34
rect 53 33 54 34
rect 52 33 53 34
rect 51 33 52 34
rect 50 33 51 34
rect 49 33 50 34
rect 48 33 49 34
rect 47 33 48 34
rect 46 33 47 34
rect 45 33 46 34
rect 44 33 45 34
rect 43 33 44 34
rect 42 33 43 34
rect 41 33 42 34
rect 40 33 41 34
rect 39 33 40 34
rect 38 33 39 34
rect 37 33 38 34
rect 36 33 37 34
rect 35 33 36 34
rect 34 33 35 34
rect 33 33 34 34
rect 32 33 33 34
rect 31 33 32 34
rect 30 33 31 34
rect 29 33 30 34
rect 28 33 29 34
rect 27 33 28 34
rect 26 33 27 34
rect 25 33 26 34
rect 24 33 25 34
rect 23 33 24 34
rect 22 33 23 34
rect 82 34 83 35
rect 81 34 82 35
rect 80 34 81 35
rect 79 34 80 35
rect 78 34 79 35
rect 77 34 78 35
rect 76 34 77 35
rect 75 34 76 35
rect 74 34 75 35
rect 73 34 74 35
rect 72 34 73 35
rect 71 34 72 35
rect 70 34 71 35
rect 69 34 70 35
rect 68 34 69 35
rect 67 34 68 35
rect 66 34 67 35
rect 65 34 66 35
rect 64 34 65 35
rect 63 34 64 35
rect 62 34 63 35
rect 61 34 62 35
rect 60 34 61 35
rect 59 34 60 35
rect 58 34 59 35
rect 57 34 58 35
rect 56 34 57 35
rect 55 34 56 35
rect 54 34 55 35
rect 53 34 54 35
rect 52 34 53 35
rect 51 34 52 35
rect 50 34 51 35
rect 49 34 50 35
rect 48 34 49 35
rect 47 34 48 35
rect 46 34 47 35
rect 45 34 46 35
rect 44 34 45 35
rect 43 34 44 35
rect 42 34 43 35
rect 41 34 42 35
rect 40 34 41 35
rect 39 34 40 35
rect 38 34 39 35
rect 37 34 38 35
rect 36 34 37 35
rect 35 34 36 35
rect 34 34 35 35
rect 33 34 34 35
rect 32 34 33 35
rect 31 34 32 35
rect 30 34 31 35
rect 29 34 30 35
rect 28 34 29 35
rect 27 34 28 35
rect 26 34 27 35
rect 25 34 26 35
rect 24 34 25 35
rect 23 34 24 35
rect 22 34 23 35
rect 21 34 22 35
rect 146 35 147 36
rect 145 35 146 36
rect 144 35 145 36
rect 143 35 144 36
rect 142 35 143 36
rect 141 35 142 36
rect 83 35 84 36
rect 82 35 83 36
rect 81 35 82 36
rect 80 35 81 36
rect 79 35 80 36
rect 78 35 79 36
rect 77 35 78 36
rect 76 35 77 36
rect 75 35 76 36
rect 74 35 75 36
rect 73 35 74 36
rect 72 35 73 36
rect 71 35 72 36
rect 70 35 71 36
rect 69 35 70 36
rect 68 35 69 36
rect 67 35 68 36
rect 66 35 67 36
rect 65 35 66 36
rect 64 35 65 36
rect 63 35 64 36
rect 62 35 63 36
rect 61 35 62 36
rect 60 35 61 36
rect 59 35 60 36
rect 58 35 59 36
rect 57 35 58 36
rect 56 35 57 36
rect 55 35 56 36
rect 54 35 55 36
rect 53 35 54 36
rect 52 35 53 36
rect 51 35 52 36
rect 50 35 51 36
rect 49 35 50 36
rect 48 35 49 36
rect 47 35 48 36
rect 46 35 47 36
rect 45 35 46 36
rect 44 35 45 36
rect 43 35 44 36
rect 42 35 43 36
rect 41 35 42 36
rect 40 35 41 36
rect 39 35 40 36
rect 38 35 39 36
rect 37 35 38 36
rect 36 35 37 36
rect 35 35 36 36
rect 34 35 35 36
rect 33 35 34 36
rect 32 35 33 36
rect 31 35 32 36
rect 30 35 31 36
rect 29 35 30 36
rect 28 35 29 36
rect 27 35 28 36
rect 26 35 27 36
rect 25 35 26 36
rect 24 35 25 36
rect 23 35 24 36
rect 22 35 23 36
rect 21 35 22 36
rect 146 36 147 37
rect 145 36 146 37
rect 144 36 145 37
rect 143 36 144 37
rect 142 36 143 37
rect 141 36 142 37
rect 140 36 141 37
rect 139 36 140 37
rect 126 36 127 37
rect 125 36 126 37
rect 124 36 125 37
rect 123 36 124 37
rect 83 36 84 37
rect 82 36 83 37
rect 81 36 82 37
rect 80 36 81 37
rect 79 36 80 37
rect 78 36 79 37
rect 77 36 78 37
rect 76 36 77 37
rect 75 36 76 37
rect 74 36 75 37
rect 73 36 74 37
rect 72 36 73 37
rect 71 36 72 37
rect 70 36 71 37
rect 69 36 70 37
rect 68 36 69 37
rect 67 36 68 37
rect 66 36 67 37
rect 65 36 66 37
rect 64 36 65 37
rect 63 36 64 37
rect 62 36 63 37
rect 61 36 62 37
rect 60 36 61 37
rect 59 36 60 37
rect 58 36 59 37
rect 57 36 58 37
rect 56 36 57 37
rect 55 36 56 37
rect 54 36 55 37
rect 53 36 54 37
rect 52 36 53 37
rect 51 36 52 37
rect 50 36 51 37
rect 49 36 50 37
rect 48 36 49 37
rect 47 36 48 37
rect 46 36 47 37
rect 45 36 46 37
rect 44 36 45 37
rect 43 36 44 37
rect 42 36 43 37
rect 41 36 42 37
rect 40 36 41 37
rect 39 36 40 37
rect 38 36 39 37
rect 37 36 38 37
rect 36 36 37 37
rect 35 36 36 37
rect 34 36 35 37
rect 33 36 34 37
rect 32 36 33 37
rect 31 36 32 37
rect 30 36 31 37
rect 29 36 30 37
rect 28 36 29 37
rect 27 36 28 37
rect 26 36 27 37
rect 25 36 26 37
rect 24 36 25 37
rect 23 36 24 37
rect 22 36 23 37
rect 21 36 22 37
rect 20 36 21 37
rect 146 37 147 38
rect 145 37 146 38
rect 144 37 145 38
rect 143 37 144 38
rect 142 37 143 38
rect 141 37 142 38
rect 140 37 141 38
rect 139 37 140 38
rect 138 37 139 38
rect 126 37 127 38
rect 125 37 126 38
rect 124 37 125 38
rect 123 37 124 38
rect 122 37 123 38
rect 83 37 84 38
rect 82 37 83 38
rect 81 37 82 38
rect 80 37 81 38
rect 79 37 80 38
rect 78 37 79 38
rect 77 37 78 38
rect 76 37 77 38
rect 75 37 76 38
rect 74 37 75 38
rect 73 37 74 38
rect 72 37 73 38
rect 71 37 72 38
rect 70 37 71 38
rect 69 37 70 38
rect 68 37 69 38
rect 67 37 68 38
rect 66 37 67 38
rect 65 37 66 38
rect 64 37 65 38
rect 63 37 64 38
rect 62 37 63 38
rect 61 37 62 38
rect 60 37 61 38
rect 59 37 60 38
rect 58 37 59 38
rect 57 37 58 38
rect 56 37 57 38
rect 55 37 56 38
rect 47 37 48 38
rect 46 37 47 38
rect 45 37 46 38
rect 44 37 45 38
rect 43 37 44 38
rect 42 37 43 38
rect 41 37 42 38
rect 40 37 41 38
rect 39 37 40 38
rect 38 37 39 38
rect 37 37 38 38
rect 36 37 37 38
rect 35 37 36 38
rect 34 37 35 38
rect 33 37 34 38
rect 32 37 33 38
rect 31 37 32 38
rect 30 37 31 38
rect 29 37 30 38
rect 28 37 29 38
rect 27 37 28 38
rect 26 37 27 38
rect 25 37 26 38
rect 24 37 25 38
rect 23 37 24 38
rect 22 37 23 38
rect 21 37 22 38
rect 20 37 21 38
rect 146 38 147 39
rect 145 38 146 39
rect 144 38 145 39
rect 143 38 144 39
rect 142 38 143 39
rect 141 38 142 39
rect 140 38 141 39
rect 139 38 140 39
rect 138 38 139 39
rect 137 38 138 39
rect 125 38 126 39
rect 124 38 125 39
rect 123 38 124 39
rect 122 38 123 39
rect 83 38 84 39
rect 82 38 83 39
rect 81 38 82 39
rect 80 38 81 39
rect 79 38 80 39
rect 78 38 79 39
rect 77 38 78 39
rect 76 38 77 39
rect 75 38 76 39
rect 74 38 75 39
rect 73 38 74 39
rect 72 38 73 39
rect 71 38 72 39
rect 70 38 71 39
rect 69 38 70 39
rect 68 38 69 39
rect 67 38 68 39
rect 66 38 67 39
rect 65 38 66 39
rect 64 38 65 39
rect 63 38 64 39
rect 62 38 63 39
rect 61 38 62 39
rect 60 38 61 39
rect 59 38 60 39
rect 43 38 44 39
rect 42 38 43 39
rect 41 38 42 39
rect 40 38 41 39
rect 39 38 40 39
rect 38 38 39 39
rect 37 38 38 39
rect 36 38 37 39
rect 35 38 36 39
rect 34 38 35 39
rect 33 38 34 39
rect 32 38 33 39
rect 31 38 32 39
rect 30 38 31 39
rect 29 38 30 39
rect 28 38 29 39
rect 27 38 28 39
rect 26 38 27 39
rect 25 38 26 39
rect 24 38 25 39
rect 23 38 24 39
rect 22 38 23 39
rect 21 38 22 39
rect 20 38 21 39
rect 19 38 20 39
rect 146 39 147 40
rect 145 39 146 40
rect 144 39 145 40
rect 143 39 144 40
rect 142 39 143 40
rect 141 39 142 40
rect 140 39 141 40
rect 139 39 140 40
rect 138 39 139 40
rect 137 39 138 40
rect 136 39 137 40
rect 125 39 126 40
rect 124 39 125 40
rect 123 39 124 40
rect 122 39 123 40
rect 84 39 85 40
rect 83 39 84 40
rect 82 39 83 40
rect 81 39 82 40
rect 80 39 81 40
rect 79 39 80 40
rect 78 39 79 40
rect 77 39 78 40
rect 76 39 77 40
rect 75 39 76 40
rect 74 39 75 40
rect 73 39 74 40
rect 72 39 73 40
rect 71 39 72 40
rect 70 39 71 40
rect 69 39 70 40
rect 68 39 69 40
rect 67 39 68 40
rect 66 39 67 40
rect 65 39 66 40
rect 64 39 65 40
rect 63 39 64 40
rect 62 39 63 40
rect 61 39 62 40
rect 41 39 42 40
rect 40 39 41 40
rect 39 39 40 40
rect 38 39 39 40
rect 37 39 38 40
rect 36 39 37 40
rect 35 39 36 40
rect 34 39 35 40
rect 33 39 34 40
rect 32 39 33 40
rect 31 39 32 40
rect 30 39 31 40
rect 29 39 30 40
rect 28 39 29 40
rect 27 39 28 40
rect 26 39 27 40
rect 25 39 26 40
rect 24 39 25 40
rect 23 39 24 40
rect 22 39 23 40
rect 21 39 22 40
rect 20 39 21 40
rect 19 39 20 40
rect 146 40 147 41
rect 145 40 146 41
rect 144 40 145 41
rect 143 40 144 41
rect 142 40 143 41
rect 141 40 142 41
rect 140 40 141 41
rect 139 40 140 41
rect 138 40 139 41
rect 137 40 138 41
rect 136 40 137 41
rect 125 40 126 41
rect 124 40 125 41
rect 123 40 124 41
rect 122 40 123 41
rect 121 40 122 41
rect 84 40 85 41
rect 83 40 84 41
rect 82 40 83 41
rect 81 40 82 41
rect 80 40 81 41
rect 79 40 80 41
rect 78 40 79 41
rect 77 40 78 41
rect 76 40 77 41
rect 75 40 76 41
rect 74 40 75 41
rect 73 40 74 41
rect 72 40 73 41
rect 71 40 72 41
rect 70 40 71 41
rect 69 40 70 41
rect 68 40 69 41
rect 67 40 68 41
rect 66 40 67 41
rect 65 40 66 41
rect 64 40 65 41
rect 63 40 64 41
rect 62 40 63 41
rect 40 40 41 41
rect 39 40 40 41
rect 38 40 39 41
rect 37 40 38 41
rect 36 40 37 41
rect 35 40 36 41
rect 34 40 35 41
rect 33 40 34 41
rect 32 40 33 41
rect 31 40 32 41
rect 30 40 31 41
rect 29 40 30 41
rect 28 40 29 41
rect 27 40 28 41
rect 26 40 27 41
rect 25 40 26 41
rect 24 40 25 41
rect 23 40 24 41
rect 22 40 23 41
rect 21 40 22 41
rect 20 40 21 41
rect 19 40 20 41
rect 146 41 147 42
rect 145 41 146 42
rect 144 41 145 42
rect 143 41 144 42
rect 142 41 143 42
rect 140 41 141 42
rect 139 41 140 42
rect 138 41 139 42
rect 137 41 138 42
rect 136 41 137 42
rect 135 41 136 42
rect 124 41 125 42
rect 123 41 124 42
rect 122 41 123 42
rect 121 41 122 42
rect 84 41 85 42
rect 83 41 84 42
rect 82 41 83 42
rect 81 41 82 42
rect 80 41 81 42
rect 79 41 80 42
rect 78 41 79 42
rect 77 41 78 42
rect 76 41 77 42
rect 75 41 76 42
rect 74 41 75 42
rect 73 41 74 42
rect 72 41 73 42
rect 71 41 72 42
rect 70 41 71 42
rect 69 41 70 42
rect 68 41 69 42
rect 67 41 68 42
rect 66 41 67 42
rect 65 41 66 42
rect 64 41 65 42
rect 38 41 39 42
rect 37 41 38 42
rect 36 41 37 42
rect 35 41 36 42
rect 34 41 35 42
rect 33 41 34 42
rect 32 41 33 42
rect 31 41 32 42
rect 30 41 31 42
rect 29 41 30 42
rect 28 41 29 42
rect 27 41 28 42
rect 26 41 27 42
rect 25 41 26 42
rect 24 41 25 42
rect 23 41 24 42
rect 22 41 23 42
rect 21 41 22 42
rect 20 41 21 42
rect 19 41 20 42
rect 18 41 19 42
rect 146 42 147 43
rect 145 42 146 43
rect 144 42 145 43
rect 143 42 144 43
rect 142 42 143 43
rect 139 42 140 43
rect 138 42 139 43
rect 137 42 138 43
rect 136 42 137 43
rect 135 42 136 43
rect 134 42 135 43
rect 124 42 125 43
rect 123 42 124 43
rect 122 42 123 43
rect 121 42 122 43
rect 84 42 85 43
rect 83 42 84 43
rect 82 42 83 43
rect 81 42 82 43
rect 80 42 81 43
rect 79 42 80 43
rect 78 42 79 43
rect 77 42 78 43
rect 76 42 77 43
rect 75 42 76 43
rect 74 42 75 43
rect 73 42 74 43
rect 72 42 73 43
rect 71 42 72 43
rect 70 42 71 43
rect 69 42 70 43
rect 68 42 69 43
rect 67 42 68 43
rect 66 42 67 43
rect 65 42 66 43
rect 37 42 38 43
rect 36 42 37 43
rect 35 42 36 43
rect 34 42 35 43
rect 33 42 34 43
rect 32 42 33 43
rect 31 42 32 43
rect 30 42 31 43
rect 29 42 30 43
rect 28 42 29 43
rect 27 42 28 43
rect 26 42 27 43
rect 25 42 26 43
rect 24 42 25 43
rect 23 42 24 43
rect 22 42 23 43
rect 21 42 22 43
rect 20 42 21 43
rect 19 42 20 43
rect 18 42 19 43
rect 146 43 147 44
rect 145 43 146 44
rect 144 43 145 44
rect 143 43 144 44
rect 142 43 143 44
rect 138 43 139 44
rect 137 43 138 44
rect 136 43 137 44
rect 135 43 136 44
rect 134 43 135 44
rect 133 43 134 44
rect 125 43 126 44
rect 124 43 125 44
rect 123 43 124 44
rect 122 43 123 44
rect 121 43 122 44
rect 84 43 85 44
rect 83 43 84 44
rect 82 43 83 44
rect 81 43 82 44
rect 80 43 81 44
rect 79 43 80 44
rect 78 43 79 44
rect 77 43 78 44
rect 76 43 77 44
rect 75 43 76 44
rect 74 43 75 44
rect 73 43 74 44
rect 72 43 73 44
rect 71 43 72 44
rect 70 43 71 44
rect 69 43 70 44
rect 68 43 69 44
rect 67 43 68 44
rect 66 43 67 44
rect 36 43 37 44
rect 35 43 36 44
rect 34 43 35 44
rect 33 43 34 44
rect 32 43 33 44
rect 31 43 32 44
rect 30 43 31 44
rect 29 43 30 44
rect 28 43 29 44
rect 27 43 28 44
rect 26 43 27 44
rect 25 43 26 44
rect 24 43 25 44
rect 23 43 24 44
rect 22 43 23 44
rect 21 43 22 44
rect 20 43 21 44
rect 19 43 20 44
rect 18 43 19 44
rect 146 44 147 45
rect 145 44 146 45
rect 144 44 145 45
rect 143 44 144 45
rect 142 44 143 45
rect 137 44 138 45
rect 136 44 137 45
rect 135 44 136 45
rect 134 44 135 45
rect 133 44 134 45
rect 132 44 133 45
rect 125 44 126 45
rect 124 44 125 45
rect 123 44 124 45
rect 122 44 123 45
rect 121 44 122 45
rect 85 44 86 45
rect 84 44 85 45
rect 83 44 84 45
rect 82 44 83 45
rect 81 44 82 45
rect 80 44 81 45
rect 79 44 80 45
rect 78 44 79 45
rect 77 44 78 45
rect 76 44 77 45
rect 75 44 76 45
rect 74 44 75 45
rect 73 44 74 45
rect 72 44 73 45
rect 71 44 72 45
rect 70 44 71 45
rect 69 44 70 45
rect 68 44 69 45
rect 67 44 68 45
rect 66 44 67 45
rect 36 44 37 45
rect 35 44 36 45
rect 34 44 35 45
rect 33 44 34 45
rect 32 44 33 45
rect 31 44 32 45
rect 30 44 31 45
rect 29 44 30 45
rect 28 44 29 45
rect 27 44 28 45
rect 26 44 27 45
rect 25 44 26 45
rect 24 44 25 45
rect 23 44 24 45
rect 22 44 23 45
rect 21 44 22 45
rect 20 44 21 45
rect 19 44 20 45
rect 18 44 19 45
rect 146 45 147 46
rect 145 45 146 46
rect 144 45 145 46
rect 143 45 144 46
rect 142 45 143 46
rect 137 45 138 46
rect 136 45 137 46
rect 135 45 136 46
rect 134 45 135 46
rect 133 45 134 46
rect 132 45 133 46
rect 131 45 132 46
rect 126 45 127 46
rect 125 45 126 46
rect 124 45 125 46
rect 123 45 124 46
rect 122 45 123 46
rect 121 45 122 46
rect 85 45 86 46
rect 84 45 85 46
rect 83 45 84 46
rect 82 45 83 46
rect 81 45 82 46
rect 80 45 81 46
rect 79 45 80 46
rect 78 45 79 46
rect 77 45 78 46
rect 76 45 77 46
rect 75 45 76 46
rect 74 45 75 46
rect 73 45 74 46
rect 72 45 73 46
rect 71 45 72 46
rect 70 45 71 46
rect 69 45 70 46
rect 68 45 69 46
rect 67 45 68 46
rect 35 45 36 46
rect 34 45 35 46
rect 33 45 34 46
rect 32 45 33 46
rect 31 45 32 46
rect 30 45 31 46
rect 29 45 30 46
rect 28 45 29 46
rect 27 45 28 46
rect 26 45 27 46
rect 25 45 26 46
rect 24 45 25 46
rect 23 45 24 46
rect 22 45 23 46
rect 21 45 22 46
rect 20 45 21 46
rect 19 45 20 46
rect 18 45 19 46
rect 146 46 147 47
rect 145 46 146 47
rect 144 46 145 47
rect 143 46 144 47
rect 142 46 143 47
rect 136 46 137 47
rect 135 46 136 47
rect 134 46 135 47
rect 133 46 134 47
rect 132 46 133 47
rect 131 46 132 47
rect 130 46 131 47
rect 129 46 130 47
rect 128 46 129 47
rect 127 46 128 47
rect 126 46 127 47
rect 125 46 126 47
rect 124 46 125 47
rect 123 46 124 47
rect 122 46 123 47
rect 121 46 122 47
rect 85 46 86 47
rect 84 46 85 47
rect 83 46 84 47
rect 82 46 83 47
rect 81 46 82 47
rect 80 46 81 47
rect 79 46 80 47
rect 78 46 79 47
rect 77 46 78 47
rect 76 46 77 47
rect 75 46 76 47
rect 74 46 75 47
rect 73 46 74 47
rect 72 46 73 47
rect 71 46 72 47
rect 70 46 71 47
rect 69 46 70 47
rect 68 46 69 47
rect 67 46 68 47
rect 35 46 36 47
rect 34 46 35 47
rect 33 46 34 47
rect 32 46 33 47
rect 31 46 32 47
rect 30 46 31 47
rect 29 46 30 47
rect 28 46 29 47
rect 27 46 28 47
rect 26 46 27 47
rect 25 46 26 47
rect 24 46 25 47
rect 23 46 24 47
rect 22 46 23 47
rect 21 46 22 47
rect 20 46 21 47
rect 19 46 20 47
rect 18 46 19 47
rect 17 46 18 47
rect 146 47 147 48
rect 145 47 146 48
rect 144 47 145 48
rect 143 47 144 48
rect 142 47 143 48
rect 135 47 136 48
rect 134 47 135 48
rect 133 47 134 48
rect 132 47 133 48
rect 131 47 132 48
rect 130 47 131 48
rect 129 47 130 48
rect 128 47 129 48
rect 127 47 128 48
rect 126 47 127 48
rect 125 47 126 48
rect 124 47 125 48
rect 123 47 124 48
rect 122 47 123 48
rect 85 47 86 48
rect 84 47 85 48
rect 83 47 84 48
rect 82 47 83 48
rect 81 47 82 48
rect 80 47 81 48
rect 79 47 80 48
rect 78 47 79 48
rect 77 47 78 48
rect 76 47 77 48
rect 75 47 76 48
rect 74 47 75 48
rect 73 47 74 48
rect 72 47 73 48
rect 71 47 72 48
rect 70 47 71 48
rect 69 47 70 48
rect 68 47 69 48
rect 34 47 35 48
rect 33 47 34 48
rect 32 47 33 48
rect 31 47 32 48
rect 30 47 31 48
rect 29 47 30 48
rect 28 47 29 48
rect 27 47 28 48
rect 26 47 27 48
rect 25 47 26 48
rect 24 47 25 48
rect 23 47 24 48
rect 22 47 23 48
rect 21 47 22 48
rect 20 47 21 48
rect 19 47 20 48
rect 18 47 19 48
rect 17 47 18 48
rect 146 48 147 49
rect 145 48 146 49
rect 144 48 145 49
rect 143 48 144 49
rect 142 48 143 49
rect 134 48 135 49
rect 133 48 134 49
rect 132 48 133 49
rect 131 48 132 49
rect 130 48 131 49
rect 129 48 130 49
rect 128 48 129 49
rect 127 48 128 49
rect 126 48 127 49
rect 125 48 126 49
rect 124 48 125 49
rect 123 48 124 49
rect 122 48 123 49
rect 85 48 86 49
rect 84 48 85 49
rect 83 48 84 49
rect 82 48 83 49
rect 81 48 82 49
rect 80 48 81 49
rect 79 48 80 49
rect 78 48 79 49
rect 77 48 78 49
rect 76 48 77 49
rect 75 48 76 49
rect 74 48 75 49
rect 73 48 74 49
rect 72 48 73 49
rect 71 48 72 49
rect 70 48 71 49
rect 69 48 70 49
rect 68 48 69 49
rect 34 48 35 49
rect 33 48 34 49
rect 32 48 33 49
rect 31 48 32 49
rect 30 48 31 49
rect 29 48 30 49
rect 28 48 29 49
rect 27 48 28 49
rect 26 48 27 49
rect 25 48 26 49
rect 24 48 25 49
rect 23 48 24 49
rect 22 48 23 49
rect 21 48 22 49
rect 20 48 21 49
rect 19 48 20 49
rect 18 48 19 49
rect 17 48 18 49
rect 146 49 147 50
rect 145 49 146 50
rect 144 49 145 50
rect 143 49 144 50
rect 142 49 143 50
rect 133 49 134 50
rect 132 49 133 50
rect 131 49 132 50
rect 130 49 131 50
rect 129 49 130 50
rect 128 49 129 50
rect 127 49 128 50
rect 126 49 127 50
rect 125 49 126 50
rect 124 49 125 50
rect 123 49 124 50
rect 85 49 86 50
rect 84 49 85 50
rect 83 49 84 50
rect 82 49 83 50
rect 81 49 82 50
rect 80 49 81 50
rect 79 49 80 50
rect 78 49 79 50
rect 77 49 78 50
rect 76 49 77 50
rect 75 49 76 50
rect 74 49 75 50
rect 73 49 74 50
rect 72 49 73 50
rect 71 49 72 50
rect 70 49 71 50
rect 69 49 70 50
rect 68 49 69 50
rect 34 49 35 50
rect 33 49 34 50
rect 32 49 33 50
rect 31 49 32 50
rect 30 49 31 50
rect 29 49 30 50
rect 28 49 29 50
rect 27 49 28 50
rect 26 49 27 50
rect 25 49 26 50
rect 24 49 25 50
rect 23 49 24 50
rect 22 49 23 50
rect 21 49 22 50
rect 20 49 21 50
rect 19 49 20 50
rect 18 49 19 50
rect 17 49 18 50
rect 146 50 147 51
rect 145 50 146 51
rect 144 50 145 51
rect 143 50 144 51
rect 142 50 143 51
rect 132 50 133 51
rect 131 50 132 51
rect 130 50 131 51
rect 129 50 130 51
rect 128 50 129 51
rect 127 50 128 51
rect 126 50 127 51
rect 125 50 126 51
rect 124 50 125 51
rect 85 50 86 51
rect 84 50 85 51
rect 83 50 84 51
rect 82 50 83 51
rect 81 50 82 51
rect 80 50 81 51
rect 79 50 80 51
rect 78 50 79 51
rect 77 50 78 51
rect 76 50 77 51
rect 75 50 76 51
rect 74 50 75 51
rect 73 50 74 51
rect 72 50 73 51
rect 71 50 72 51
rect 70 50 71 51
rect 69 50 70 51
rect 33 50 34 51
rect 32 50 33 51
rect 31 50 32 51
rect 30 50 31 51
rect 29 50 30 51
rect 28 50 29 51
rect 27 50 28 51
rect 26 50 27 51
rect 25 50 26 51
rect 24 50 25 51
rect 23 50 24 51
rect 22 50 23 51
rect 21 50 22 51
rect 20 50 21 51
rect 19 50 20 51
rect 18 50 19 51
rect 17 50 18 51
rect 146 51 147 52
rect 145 51 146 52
rect 144 51 145 52
rect 143 51 144 52
rect 142 51 143 52
rect 129 51 130 52
rect 128 51 129 52
rect 127 51 128 52
rect 85 51 86 52
rect 84 51 85 52
rect 83 51 84 52
rect 82 51 83 52
rect 81 51 82 52
rect 80 51 81 52
rect 79 51 80 52
rect 78 51 79 52
rect 77 51 78 52
rect 76 51 77 52
rect 75 51 76 52
rect 74 51 75 52
rect 73 51 74 52
rect 72 51 73 52
rect 71 51 72 52
rect 70 51 71 52
rect 69 51 70 52
rect 33 51 34 52
rect 32 51 33 52
rect 31 51 32 52
rect 30 51 31 52
rect 29 51 30 52
rect 28 51 29 52
rect 27 51 28 52
rect 26 51 27 52
rect 25 51 26 52
rect 24 51 25 52
rect 23 51 24 52
rect 22 51 23 52
rect 21 51 22 52
rect 20 51 21 52
rect 19 51 20 52
rect 18 51 19 52
rect 17 51 18 52
rect 85 52 86 53
rect 84 52 85 53
rect 83 52 84 53
rect 82 52 83 53
rect 81 52 82 53
rect 80 52 81 53
rect 79 52 80 53
rect 78 52 79 53
rect 77 52 78 53
rect 76 52 77 53
rect 75 52 76 53
rect 74 52 75 53
rect 73 52 74 53
rect 72 52 73 53
rect 71 52 72 53
rect 70 52 71 53
rect 69 52 70 53
rect 33 52 34 53
rect 32 52 33 53
rect 31 52 32 53
rect 30 52 31 53
rect 29 52 30 53
rect 28 52 29 53
rect 27 52 28 53
rect 26 52 27 53
rect 25 52 26 53
rect 24 52 25 53
rect 23 52 24 53
rect 22 52 23 53
rect 21 52 22 53
rect 20 52 21 53
rect 19 52 20 53
rect 18 52 19 53
rect 17 52 18 53
rect 85 53 86 54
rect 84 53 85 54
rect 83 53 84 54
rect 82 53 83 54
rect 81 53 82 54
rect 80 53 81 54
rect 79 53 80 54
rect 78 53 79 54
rect 77 53 78 54
rect 76 53 77 54
rect 75 53 76 54
rect 74 53 75 54
rect 73 53 74 54
rect 72 53 73 54
rect 71 53 72 54
rect 70 53 71 54
rect 69 53 70 54
rect 33 53 34 54
rect 32 53 33 54
rect 31 53 32 54
rect 30 53 31 54
rect 29 53 30 54
rect 28 53 29 54
rect 27 53 28 54
rect 26 53 27 54
rect 25 53 26 54
rect 24 53 25 54
rect 23 53 24 54
rect 22 53 23 54
rect 21 53 22 54
rect 20 53 21 54
rect 19 53 20 54
rect 18 53 19 54
rect 17 53 18 54
rect 85 54 86 55
rect 84 54 85 55
rect 83 54 84 55
rect 82 54 83 55
rect 81 54 82 55
rect 80 54 81 55
rect 79 54 80 55
rect 78 54 79 55
rect 77 54 78 55
rect 76 54 77 55
rect 75 54 76 55
rect 74 54 75 55
rect 73 54 74 55
rect 72 54 73 55
rect 71 54 72 55
rect 70 54 71 55
rect 69 54 70 55
rect 33 54 34 55
rect 32 54 33 55
rect 31 54 32 55
rect 30 54 31 55
rect 29 54 30 55
rect 28 54 29 55
rect 27 54 28 55
rect 26 54 27 55
rect 25 54 26 55
rect 24 54 25 55
rect 23 54 24 55
rect 22 54 23 55
rect 21 54 22 55
rect 20 54 21 55
rect 19 54 20 55
rect 18 54 19 55
rect 17 54 18 55
rect 85 55 86 56
rect 84 55 85 56
rect 83 55 84 56
rect 82 55 83 56
rect 81 55 82 56
rect 80 55 81 56
rect 79 55 80 56
rect 78 55 79 56
rect 77 55 78 56
rect 76 55 77 56
rect 75 55 76 56
rect 74 55 75 56
rect 73 55 74 56
rect 72 55 73 56
rect 71 55 72 56
rect 70 55 71 56
rect 69 55 70 56
rect 33 55 34 56
rect 32 55 33 56
rect 31 55 32 56
rect 30 55 31 56
rect 29 55 30 56
rect 28 55 29 56
rect 27 55 28 56
rect 26 55 27 56
rect 25 55 26 56
rect 24 55 25 56
rect 23 55 24 56
rect 22 55 23 56
rect 21 55 22 56
rect 20 55 21 56
rect 19 55 20 56
rect 18 55 19 56
rect 17 55 18 56
rect 139 56 140 57
rect 138 56 139 57
rect 137 56 138 57
rect 136 56 137 57
rect 135 56 136 57
rect 134 56 135 57
rect 133 56 134 57
rect 132 56 133 57
rect 131 56 132 57
rect 130 56 131 57
rect 129 56 130 57
rect 128 56 129 57
rect 85 56 86 57
rect 84 56 85 57
rect 83 56 84 57
rect 82 56 83 57
rect 81 56 82 57
rect 80 56 81 57
rect 79 56 80 57
rect 78 56 79 57
rect 77 56 78 57
rect 76 56 77 57
rect 75 56 76 57
rect 74 56 75 57
rect 73 56 74 57
rect 72 56 73 57
rect 71 56 72 57
rect 70 56 71 57
rect 69 56 70 57
rect 33 56 34 57
rect 32 56 33 57
rect 31 56 32 57
rect 30 56 31 57
rect 29 56 30 57
rect 28 56 29 57
rect 27 56 28 57
rect 26 56 27 57
rect 25 56 26 57
rect 24 56 25 57
rect 23 56 24 57
rect 22 56 23 57
rect 21 56 22 57
rect 20 56 21 57
rect 19 56 20 57
rect 18 56 19 57
rect 17 56 18 57
rect 142 57 143 58
rect 141 57 142 58
rect 140 57 141 58
rect 139 57 140 58
rect 138 57 139 58
rect 137 57 138 58
rect 136 57 137 58
rect 135 57 136 58
rect 134 57 135 58
rect 133 57 134 58
rect 132 57 133 58
rect 131 57 132 58
rect 130 57 131 58
rect 129 57 130 58
rect 128 57 129 58
rect 127 57 128 58
rect 126 57 127 58
rect 85 57 86 58
rect 84 57 85 58
rect 83 57 84 58
rect 82 57 83 58
rect 81 57 82 58
rect 80 57 81 58
rect 79 57 80 58
rect 78 57 79 58
rect 77 57 78 58
rect 76 57 77 58
rect 75 57 76 58
rect 74 57 75 58
rect 73 57 74 58
rect 72 57 73 58
rect 71 57 72 58
rect 70 57 71 58
rect 69 57 70 58
rect 33 57 34 58
rect 32 57 33 58
rect 31 57 32 58
rect 30 57 31 58
rect 29 57 30 58
rect 28 57 29 58
rect 27 57 28 58
rect 26 57 27 58
rect 25 57 26 58
rect 24 57 25 58
rect 23 57 24 58
rect 22 57 23 58
rect 21 57 22 58
rect 20 57 21 58
rect 19 57 20 58
rect 18 57 19 58
rect 17 57 18 58
rect 143 58 144 59
rect 142 58 143 59
rect 141 58 142 59
rect 140 58 141 59
rect 139 58 140 59
rect 138 58 139 59
rect 137 58 138 59
rect 136 58 137 59
rect 135 58 136 59
rect 134 58 135 59
rect 133 58 134 59
rect 132 58 133 59
rect 131 58 132 59
rect 130 58 131 59
rect 129 58 130 59
rect 128 58 129 59
rect 127 58 128 59
rect 126 58 127 59
rect 125 58 126 59
rect 124 58 125 59
rect 84 58 85 59
rect 83 58 84 59
rect 82 58 83 59
rect 81 58 82 59
rect 80 58 81 59
rect 79 58 80 59
rect 78 58 79 59
rect 77 58 78 59
rect 76 58 77 59
rect 75 58 76 59
rect 74 58 75 59
rect 73 58 74 59
rect 72 58 73 59
rect 71 58 72 59
rect 70 58 71 59
rect 69 58 70 59
rect 33 58 34 59
rect 32 58 33 59
rect 31 58 32 59
rect 30 58 31 59
rect 29 58 30 59
rect 28 58 29 59
rect 27 58 28 59
rect 26 58 27 59
rect 25 58 26 59
rect 24 58 25 59
rect 23 58 24 59
rect 22 58 23 59
rect 21 58 22 59
rect 20 58 21 59
rect 19 58 20 59
rect 18 58 19 59
rect 17 58 18 59
rect 144 59 145 60
rect 143 59 144 60
rect 142 59 143 60
rect 141 59 142 60
rect 140 59 141 60
rect 139 59 140 60
rect 138 59 139 60
rect 137 59 138 60
rect 136 59 137 60
rect 135 59 136 60
rect 134 59 135 60
rect 133 59 134 60
rect 132 59 133 60
rect 131 59 132 60
rect 130 59 131 60
rect 129 59 130 60
rect 128 59 129 60
rect 127 59 128 60
rect 126 59 127 60
rect 125 59 126 60
rect 124 59 125 60
rect 123 59 124 60
rect 84 59 85 60
rect 83 59 84 60
rect 82 59 83 60
rect 81 59 82 60
rect 80 59 81 60
rect 79 59 80 60
rect 78 59 79 60
rect 77 59 78 60
rect 76 59 77 60
rect 75 59 76 60
rect 74 59 75 60
rect 73 59 74 60
rect 72 59 73 60
rect 71 59 72 60
rect 70 59 71 60
rect 69 59 70 60
rect 33 59 34 60
rect 32 59 33 60
rect 31 59 32 60
rect 30 59 31 60
rect 29 59 30 60
rect 28 59 29 60
rect 27 59 28 60
rect 26 59 27 60
rect 25 59 26 60
rect 24 59 25 60
rect 23 59 24 60
rect 22 59 23 60
rect 21 59 22 60
rect 20 59 21 60
rect 19 59 20 60
rect 18 59 19 60
rect 17 59 18 60
rect 145 60 146 61
rect 144 60 145 61
rect 143 60 144 61
rect 142 60 143 61
rect 141 60 142 61
rect 140 60 141 61
rect 139 60 140 61
rect 138 60 139 61
rect 137 60 138 61
rect 136 60 137 61
rect 135 60 136 61
rect 134 60 135 61
rect 133 60 134 61
rect 132 60 133 61
rect 131 60 132 61
rect 130 60 131 61
rect 129 60 130 61
rect 128 60 129 61
rect 127 60 128 61
rect 126 60 127 61
rect 125 60 126 61
rect 124 60 125 61
rect 123 60 124 61
rect 122 60 123 61
rect 84 60 85 61
rect 83 60 84 61
rect 82 60 83 61
rect 81 60 82 61
rect 80 60 81 61
rect 79 60 80 61
rect 78 60 79 61
rect 77 60 78 61
rect 76 60 77 61
rect 75 60 76 61
rect 74 60 75 61
rect 73 60 74 61
rect 72 60 73 61
rect 71 60 72 61
rect 70 60 71 61
rect 69 60 70 61
rect 68 60 69 61
rect 33 60 34 61
rect 32 60 33 61
rect 31 60 32 61
rect 30 60 31 61
rect 29 60 30 61
rect 28 60 29 61
rect 27 60 28 61
rect 26 60 27 61
rect 25 60 26 61
rect 24 60 25 61
rect 23 60 24 61
rect 22 60 23 61
rect 21 60 22 61
rect 20 60 21 61
rect 19 60 20 61
rect 18 60 19 61
rect 145 61 146 62
rect 144 61 145 62
rect 143 61 144 62
rect 142 61 143 62
rect 141 61 142 62
rect 140 61 141 62
rect 139 61 140 62
rect 138 61 139 62
rect 137 61 138 62
rect 130 61 131 62
rect 129 61 130 62
rect 128 61 129 62
rect 127 61 128 62
rect 126 61 127 62
rect 125 61 126 62
rect 124 61 125 62
rect 123 61 124 62
rect 122 61 123 62
rect 84 61 85 62
rect 83 61 84 62
rect 82 61 83 62
rect 81 61 82 62
rect 80 61 81 62
rect 79 61 80 62
rect 78 61 79 62
rect 77 61 78 62
rect 76 61 77 62
rect 75 61 76 62
rect 74 61 75 62
rect 73 61 74 62
rect 72 61 73 62
rect 71 61 72 62
rect 70 61 71 62
rect 69 61 70 62
rect 68 61 69 62
rect 34 61 35 62
rect 33 61 34 62
rect 32 61 33 62
rect 31 61 32 62
rect 30 61 31 62
rect 29 61 30 62
rect 28 61 29 62
rect 27 61 28 62
rect 26 61 27 62
rect 25 61 26 62
rect 24 61 25 62
rect 23 61 24 62
rect 22 61 23 62
rect 21 61 22 62
rect 20 61 21 62
rect 19 61 20 62
rect 18 61 19 62
rect 146 62 147 63
rect 145 62 146 63
rect 144 62 145 63
rect 143 62 144 63
rect 142 62 143 63
rect 141 62 142 63
rect 126 62 127 63
rect 125 62 126 63
rect 124 62 125 63
rect 123 62 124 63
rect 122 62 123 63
rect 121 62 122 63
rect 84 62 85 63
rect 83 62 84 63
rect 82 62 83 63
rect 81 62 82 63
rect 80 62 81 63
rect 79 62 80 63
rect 78 62 79 63
rect 77 62 78 63
rect 76 62 77 63
rect 75 62 76 63
rect 74 62 75 63
rect 73 62 74 63
rect 72 62 73 63
rect 71 62 72 63
rect 70 62 71 63
rect 69 62 70 63
rect 68 62 69 63
rect 34 62 35 63
rect 33 62 34 63
rect 32 62 33 63
rect 31 62 32 63
rect 30 62 31 63
rect 29 62 30 63
rect 28 62 29 63
rect 27 62 28 63
rect 26 62 27 63
rect 25 62 26 63
rect 24 62 25 63
rect 23 62 24 63
rect 22 62 23 63
rect 21 62 22 63
rect 20 62 21 63
rect 19 62 20 63
rect 18 62 19 63
rect 146 63 147 64
rect 145 63 146 64
rect 144 63 145 64
rect 143 63 144 64
rect 142 63 143 64
rect 125 63 126 64
rect 124 63 125 64
rect 123 63 124 64
rect 122 63 123 64
rect 121 63 122 64
rect 84 63 85 64
rect 83 63 84 64
rect 82 63 83 64
rect 81 63 82 64
rect 80 63 81 64
rect 79 63 80 64
rect 78 63 79 64
rect 77 63 78 64
rect 76 63 77 64
rect 75 63 76 64
rect 74 63 75 64
rect 73 63 74 64
rect 72 63 73 64
rect 71 63 72 64
rect 70 63 71 64
rect 69 63 70 64
rect 68 63 69 64
rect 34 63 35 64
rect 33 63 34 64
rect 32 63 33 64
rect 31 63 32 64
rect 30 63 31 64
rect 29 63 30 64
rect 28 63 29 64
rect 27 63 28 64
rect 26 63 27 64
rect 25 63 26 64
rect 24 63 25 64
rect 23 63 24 64
rect 22 63 23 64
rect 21 63 22 64
rect 20 63 21 64
rect 19 63 20 64
rect 18 63 19 64
rect 146 64 147 65
rect 145 64 146 65
rect 144 64 145 65
rect 143 64 144 65
rect 124 64 125 65
rect 123 64 124 65
rect 122 64 123 65
rect 121 64 122 65
rect 83 64 84 65
rect 82 64 83 65
rect 81 64 82 65
rect 80 64 81 65
rect 79 64 80 65
rect 78 64 79 65
rect 77 64 78 65
rect 76 64 77 65
rect 75 64 76 65
rect 74 64 75 65
rect 73 64 74 65
rect 72 64 73 65
rect 71 64 72 65
rect 70 64 71 65
rect 69 64 70 65
rect 68 64 69 65
rect 67 64 68 65
rect 35 64 36 65
rect 34 64 35 65
rect 33 64 34 65
rect 32 64 33 65
rect 31 64 32 65
rect 30 64 31 65
rect 29 64 30 65
rect 28 64 29 65
rect 27 64 28 65
rect 26 64 27 65
rect 25 64 26 65
rect 24 64 25 65
rect 23 64 24 65
rect 22 64 23 65
rect 21 64 22 65
rect 20 64 21 65
rect 19 64 20 65
rect 18 64 19 65
rect 146 65 147 66
rect 145 65 146 66
rect 144 65 145 66
rect 143 65 144 66
rect 124 65 125 66
rect 123 65 124 66
rect 122 65 123 66
rect 121 65 122 66
rect 83 65 84 66
rect 82 65 83 66
rect 81 65 82 66
rect 80 65 81 66
rect 79 65 80 66
rect 78 65 79 66
rect 77 65 78 66
rect 76 65 77 66
rect 75 65 76 66
rect 74 65 75 66
rect 73 65 74 66
rect 72 65 73 66
rect 71 65 72 66
rect 70 65 71 66
rect 69 65 70 66
rect 68 65 69 66
rect 67 65 68 66
rect 35 65 36 66
rect 34 65 35 66
rect 33 65 34 66
rect 32 65 33 66
rect 31 65 32 66
rect 30 65 31 66
rect 29 65 30 66
rect 28 65 29 66
rect 27 65 28 66
rect 26 65 27 66
rect 25 65 26 66
rect 24 65 25 66
rect 23 65 24 66
rect 22 65 23 66
rect 21 65 22 66
rect 20 65 21 66
rect 19 65 20 66
rect 18 65 19 66
rect 146 66 147 67
rect 145 66 146 67
rect 144 66 145 67
rect 143 66 144 67
rect 142 66 143 67
rect 125 66 126 67
rect 124 66 125 67
rect 123 66 124 67
rect 122 66 123 67
rect 121 66 122 67
rect 83 66 84 67
rect 82 66 83 67
rect 81 66 82 67
rect 80 66 81 67
rect 79 66 80 67
rect 78 66 79 67
rect 77 66 78 67
rect 76 66 77 67
rect 75 66 76 67
rect 74 66 75 67
rect 73 66 74 67
rect 72 66 73 67
rect 71 66 72 67
rect 70 66 71 67
rect 69 66 70 67
rect 68 66 69 67
rect 67 66 68 67
rect 35 66 36 67
rect 34 66 35 67
rect 33 66 34 67
rect 32 66 33 67
rect 31 66 32 67
rect 30 66 31 67
rect 29 66 30 67
rect 28 66 29 67
rect 27 66 28 67
rect 26 66 27 67
rect 25 66 26 67
rect 24 66 25 67
rect 23 66 24 67
rect 22 66 23 67
rect 21 66 22 67
rect 20 66 21 67
rect 19 66 20 67
rect 18 66 19 67
rect 146 67 147 68
rect 145 67 146 68
rect 144 67 145 68
rect 143 67 144 68
rect 142 67 143 68
rect 141 67 142 68
rect 126 67 127 68
rect 125 67 126 68
rect 124 67 125 68
rect 123 67 124 68
rect 122 67 123 68
rect 121 67 122 68
rect 83 67 84 68
rect 82 67 83 68
rect 81 67 82 68
rect 80 67 81 68
rect 79 67 80 68
rect 78 67 79 68
rect 77 67 78 68
rect 76 67 77 68
rect 75 67 76 68
rect 74 67 75 68
rect 73 67 74 68
rect 72 67 73 68
rect 71 67 72 68
rect 70 67 71 68
rect 69 67 70 68
rect 68 67 69 68
rect 67 67 68 68
rect 66 67 67 68
rect 36 67 37 68
rect 35 67 36 68
rect 34 67 35 68
rect 33 67 34 68
rect 32 67 33 68
rect 31 67 32 68
rect 30 67 31 68
rect 29 67 30 68
rect 28 67 29 68
rect 27 67 28 68
rect 26 67 27 68
rect 25 67 26 68
rect 24 67 25 68
rect 23 67 24 68
rect 22 67 23 68
rect 21 67 22 68
rect 20 67 21 68
rect 19 67 20 68
rect 145 68 146 69
rect 144 68 145 69
rect 143 68 144 69
rect 142 68 143 69
rect 141 68 142 69
rect 140 68 141 69
rect 139 68 140 69
rect 138 68 139 69
rect 129 68 130 69
rect 128 68 129 69
rect 127 68 128 69
rect 126 68 127 69
rect 125 68 126 69
rect 124 68 125 69
rect 123 68 124 69
rect 122 68 123 69
rect 121 68 122 69
rect 82 68 83 69
rect 81 68 82 69
rect 80 68 81 69
rect 79 68 80 69
rect 78 68 79 69
rect 77 68 78 69
rect 76 68 77 69
rect 75 68 76 69
rect 74 68 75 69
rect 73 68 74 69
rect 72 68 73 69
rect 71 68 72 69
rect 70 68 71 69
rect 69 68 70 69
rect 68 68 69 69
rect 67 68 68 69
rect 66 68 67 69
rect 36 68 37 69
rect 35 68 36 69
rect 34 68 35 69
rect 33 68 34 69
rect 32 68 33 69
rect 31 68 32 69
rect 30 68 31 69
rect 29 68 30 69
rect 28 68 29 69
rect 27 68 28 69
rect 26 68 27 69
rect 25 68 26 69
rect 24 68 25 69
rect 23 68 24 69
rect 22 68 23 69
rect 21 68 22 69
rect 20 68 21 69
rect 19 68 20 69
rect 145 69 146 70
rect 144 69 145 70
rect 143 69 144 70
rect 142 69 143 70
rect 141 69 142 70
rect 140 69 141 70
rect 139 69 140 70
rect 138 69 139 70
rect 137 69 138 70
rect 136 69 137 70
rect 135 69 136 70
rect 134 69 135 70
rect 133 69 134 70
rect 132 69 133 70
rect 131 69 132 70
rect 130 69 131 70
rect 129 69 130 70
rect 128 69 129 70
rect 127 69 128 70
rect 126 69 127 70
rect 125 69 126 70
rect 124 69 125 70
rect 123 69 124 70
rect 122 69 123 70
rect 82 69 83 70
rect 81 69 82 70
rect 80 69 81 70
rect 79 69 80 70
rect 78 69 79 70
rect 77 69 78 70
rect 76 69 77 70
rect 75 69 76 70
rect 74 69 75 70
rect 73 69 74 70
rect 72 69 73 70
rect 71 69 72 70
rect 70 69 71 70
rect 69 69 70 70
rect 68 69 69 70
rect 67 69 68 70
rect 66 69 67 70
rect 65 69 66 70
rect 37 69 38 70
rect 36 69 37 70
rect 35 69 36 70
rect 34 69 35 70
rect 33 69 34 70
rect 32 69 33 70
rect 31 69 32 70
rect 30 69 31 70
rect 29 69 30 70
rect 28 69 29 70
rect 27 69 28 70
rect 26 69 27 70
rect 25 69 26 70
rect 24 69 25 70
rect 23 69 24 70
rect 22 69 23 70
rect 21 69 22 70
rect 20 69 21 70
rect 19 69 20 70
rect 144 70 145 71
rect 143 70 144 71
rect 142 70 143 71
rect 141 70 142 71
rect 140 70 141 71
rect 139 70 140 71
rect 138 70 139 71
rect 137 70 138 71
rect 136 70 137 71
rect 135 70 136 71
rect 134 70 135 71
rect 133 70 134 71
rect 132 70 133 71
rect 131 70 132 71
rect 130 70 131 71
rect 129 70 130 71
rect 128 70 129 71
rect 127 70 128 71
rect 126 70 127 71
rect 125 70 126 71
rect 124 70 125 71
rect 123 70 124 71
rect 122 70 123 71
rect 143 71 144 72
rect 142 71 143 72
rect 141 71 142 72
rect 140 71 141 72
rect 139 71 140 72
rect 138 71 139 72
rect 137 71 138 72
rect 136 71 137 72
rect 135 71 136 72
rect 134 71 135 72
rect 133 71 134 72
rect 132 71 133 72
rect 131 71 132 72
rect 130 71 131 72
rect 129 71 130 72
rect 128 71 129 72
rect 127 71 128 72
rect 126 71 127 72
rect 125 71 126 72
rect 124 71 125 72
rect 123 71 124 72
rect 142 72 143 73
rect 141 72 142 73
rect 140 72 141 73
rect 139 72 140 73
rect 138 72 139 73
rect 137 72 138 73
rect 136 72 137 73
rect 135 72 136 73
rect 134 72 135 73
rect 133 72 134 73
rect 132 72 133 73
rect 131 72 132 73
rect 130 72 131 73
rect 129 72 130 73
rect 128 72 129 73
rect 127 72 128 73
rect 126 72 127 73
rect 125 72 126 73
rect 140 73 141 74
rect 139 73 140 74
rect 138 73 139 74
rect 137 73 138 74
rect 136 73 137 74
rect 135 73 136 74
rect 134 73 135 74
rect 133 73 134 74
rect 132 73 133 74
rect 131 73 132 74
rect 130 73 131 74
rect 129 73 130 74
rect 128 73 129 74
rect 127 73 128 74
rect 146 78 147 79
rect 145 78 146 79
rect 144 78 145 79
rect 143 78 144 79
rect 142 78 143 79
rect 141 78 142 79
rect 146 79 147 80
rect 145 79 146 80
rect 144 79 145 80
rect 143 79 144 80
rect 142 79 143 80
rect 141 79 142 80
rect 140 79 141 80
rect 139 79 140 80
rect 126 79 127 80
rect 125 79 126 80
rect 124 79 125 80
rect 123 79 124 80
rect 146 80 147 81
rect 145 80 146 81
rect 144 80 145 81
rect 143 80 144 81
rect 142 80 143 81
rect 141 80 142 81
rect 140 80 141 81
rect 139 80 140 81
rect 138 80 139 81
rect 126 80 127 81
rect 125 80 126 81
rect 124 80 125 81
rect 123 80 124 81
rect 122 80 123 81
rect 84 80 85 81
rect 83 80 84 81
rect 82 80 83 81
rect 81 80 82 81
rect 80 80 81 81
rect 79 80 80 81
rect 78 80 79 81
rect 77 80 78 81
rect 76 80 77 81
rect 75 80 76 81
rect 74 80 75 81
rect 73 80 74 81
rect 72 80 73 81
rect 71 80 72 81
rect 70 80 71 81
rect 69 80 70 81
rect 68 80 69 81
rect 67 80 68 81
rect 66 80 67 81
rect 65 80 66 81
rect 64 80 65 81
rect 63 80 64 81
rect 62 80 63 81
rect 61 80 62 81
rect 60 80 61 81
rect 59 80 60 81
rect 58 80 59 81
rect 57 80 58 81
rect 56 80 57 81
rect 55 80 56 81
rect 54 80 55 81
rect 53 80 54 81
rect 52 80 53 81
rect 51 80 52 81
rect 50 80 51 81
rect 49 80 50 81
rect 48 80 49 81
rect 47 80 48 81
rect 46 80 47 81
rect 45 80 46 81
rect 44 80 45 81
rect 43 80 44 81
rect 42 80 43 81
rect 41 80 42 81
rect 40 80 41 81
rect 39 80 40 81
rect 38 80 39 81
rect 37 80 38 81
rect 36 80 37 81
rect 35 80 36 81
rect 34 80 35 81
rect 33 80 34 81
rect 32 80 33 81
rect 31 80 32 81
rect 30 80 31 81
rect 29 80 30 81
rect 28 80 29 81
rect 27 80 28 81
rect 26 80 27 81
rect 25 80 26 81
rect 24 80 25 81
rect 23 80 24 81
rect 22 80 23 81
rect 21 80 22 81
rect 20 80 21 81
rect 19 80 20 81
rect 18 80 19 81
rect 146 81 147 82
rect 145 81 146 82
rect 144 81 145 82
rect 143 81 144 82
rect 142 81 143 82
rect 141 81 142 82
rect 140 81 141 82
rect 139 81 140 82
rect 138 81 139 82
rect 137 81 138 82
rect 125 81 126 82
rect 124 81 125 82
rect 123 81 124 82
rect 122 81 123 82
rect 84 81 85 82
rect 83 81 84 82
rect 82 81 83 82
rect 81 81 82 82
rect 80 81 81 82
rect 79 81 80 82
rect 78 81 79 82
rect 77 81 78 82
rect 76 81 77 82
rect 75 81 76 82
rect 74 81 75 82
rect 73 81 74 82
rect 72 81 73 82
rect 71 81 72 82
rect 70 81 71 82
rect 69 81 70 82
rect 68 81 69 82
rect 67 81 68 82
rect 66 81 67 82
rect 65 81 66 82
rect 64 81 65 82
rect 63 81 64 82
rect 62 81 63 82
rect 61 81 62 82
rect 60 81 61 82
rect 59 81 60 82
rect 58 81 59 82
rect 57 81 58 82
rect 56 81 57 82
rect 55 81 56 82
rect 54 81 55 82
rect 53 81 54 82
rect 52 81 53 82
rect 51 81 52 82
rect 50 81 51 82
rect 49 81 50 82
rect 48 81 49 82
rect 47 81 48 82
rect 46 81 47 82
rect 45 81 46 82
rect 44 81 45 82
rect 43 81 44 82
rect 42 81 43 82
rect 41 81 42 82
rect 40 81 41 82
rect 39 81 40 82
rect 38 81 39 82
rect 37 81 38 82
rect 36 81 37 82
rect 35 81 36 82
rect 34 81 35 82
rect 33 81 34 82
rect 32 81 33 82
rect 31 81 32 82
rect 30 81 31 82
rect 29 81 30 82
rect 28 81 29 82
rect 27 81 28 82
rect 26 81 27 82
rect 25 81 26 82
rect 24 81 25 82
rect 23 81 24 82
rect 22 81 23 82
rect 21 81 22 82
rect 20 81 21 82
rect 19 81 20 82
rect 18 81 19 82
rect 146 82 147 83
rect 145 82 146 83
rect 144 82 145 83
rect 143 82 144 83
rect 142 82 143 83
rect 141 82 142 83
rect 140 82 141 83
rect 139 82 140 83
rect 138 82 139 83
rect 137 82 138 83
rect 136 82 137 83
rect 125 82 126 83
rect 124 82 125 83
rect 123 82 124 83
rect 122 82 123 83
rect 84 82 85 83
rect 83 82 84 83
rect 82 82 83 83
rect 81 82 82 83
rect 80 82 81 83
rect 79 82 80 83
rect 78 82 79 83
rect 77 82 78 83
rect 76 82 77 83
rect 75 82 76 83
rect 74 82 75 83
rect 73 82 74 83
rect 72 82 73 83
rect 71 82 72 83
rect 70 82 71 83
rect 69 82 70 83
rect 68 82 69 83
rect 67 82 68 83
rect 66 82 67 83
rect 65 82 66 83
rect 64 82 65 83
rect 63 82 64 83
rect 62 82 63 83
rect 61 82 62 83
rect 60 82 61 83
rect 59 82 60 83
rect 58 82 59 83
rect 57 82 58 83
rect 56 82 57 83
rect 55 82 56 83
rect 54 82 55 83
rect 53 82 54 83
rect 52 82 53 83
rect 51 82 52 83
rect 50 82 51 83
rect 49 82 50 83
rect 48 82 49 83
rect 47 82 48 83
rect 46 82 47 83
rect 45 82 46 83
rect 44 82 45 83
rect 43 82 44 83
rect 42 82 43 83
rect 41 82 42 83
rect 40 82 41 83
rect 39 82 40 83
rect 38 82 39 83
rect 37 82 38 83
rect 36 82 37 83
rect 35 82 36 83
rect 34 82 35 83
rect 33 82 34 83
rect 32 82 33 83
rect 31 82 32 83
rect 30 82 31 83
rect 29 82 30 83
rect 28 82 29 83
rect 27 82 28 83
rect 26 82 27 83
rect 25 82 26 83
rect 24 82 25 83
rect 23 82 24 83
rect 22 82 23 83
rect 21 82 22 83
rect 20 82 21 83
rect 19 82 20 83
rect 18 82 19 83
rect 146 83 147 84
rect 145 83 146 84
rect 144 83 145 84
rect 143 83 144 84
rect 142 83 143 84
rect 141 83 142 84
rect 140 83 141 84
rect 139 83 140 84
rect 138 83 139 84
rect 137 83 138 84
rect 136 83 137 84
rect 125 83 126 84
rect 124 83 125 84
rect 123 83 124 84
rect 122 83 123 84
rect 121 83 122 84
rect 84 83 85 84
rect 83 83 84 84
rect 82 83 83 84
rect 81 83 82 84
rect 80 83 81 84
rect 79 83 80 84
rect 78 83 79 84
rect 77 83 78 84
rect 76 83 77 84
rect 75 83 76 84
rect 74 83 75 84
rect 73 83 74 84
rect 72 83 73 84
rect 71 83 72 84
rect 70 83 71 84
rect 69 83 70 84
rect 68 83 69 84
rect 67 83 68 84
rect 66 83 67 84
rect 65 83 66 84
rect 64 83 65 84
rect 63 83 64 84
rect 62 83 63 84
rect 61 83 62 84
rect 60 83 61 84
rect 59 83 60 84
rect 58 83 59 84
rect 57 83 58 84
rect 56 83 57 84
rect 55 83 56 84
rect 54 83 55 84
rect 53 83 54 84
rect 52 83 53 84
rect 51 83 52 84
rect 50 83 51 84
rect 49 83 50 84
rect 48 83 49 84
rect 47 83 48 84
rect 46 83 47 84
rect 45 83 46 84
rect 44 83 45 84
rect 43 83 44 84
rect 42 83 43 84
rect 41 83 42 84
rect 40 83 41 84
rect 39 83 40 84
rect 38 83 39 84
rect 37 83 38 84
rect 36 83 37 84
rect 35 83 36 84
rect 34 83 35 84
rect 33 83 34 84
rect 32 83 33 84
rect 31 83 32 84
rect 30 83 31 84
rect 29 83 30 84
rect 28 83 29 84
rect 27 83 28 84
rect 26 83 27 84
rect 25 83 26 84
rect 24 83 25 84
rect 23 83 24 84
rect 22 83 23 84
rect 21 83 22 84
rect 20 83 21 84
rect 19 83 20 84
rect 18 83 19 84
rect 146 84 147 85
rect 145 84 146 85
rect 144 84 145 85
rect 143 84 144 85
rect 142 84 143 85
rect 140 84 141 85
rect 139 84 140 85
rect 138 84 139 85
rect 137 84 138 85
rect 136 84 137 85
rect 135 84 136 85
rect 124 84 125 85
rect 123 84 124 85
rect 122 84 123 85
rect 121 84 122 85
rect 84 84 85 85
rect 83 84 84 85
rect 82 84 83 85
rect 81 84 82 85
rect 80 84 81 85
rect 79 84 80 85
rect 78 84 79 85
rect 77 84 78 85
rect 76 84 77 85
rect 75 84 76 85
rect 74 84 75 85
rect 73 84 74 85
rect 72 84 73 85
rect 71 84 72 85
rect 70 84 71 85
rect 69 84 70 85
rect 68 84 69 85
rect 67 84 68 85
rect 66 84 67 85
rect 65 84 66 85
rect 64 84 65 85
rect 63 84 64 85
rect 62 84 63 85
rect 61 84 62 85
rect 60 84 61 85
rect 59 84 60 85
rect 58 84 59 85
rect 57 84 58 85
rect 56 84 57 85
rect 55 84 56 85
rect 54 84 55 85
rect 53 84 54 85
rect 52 84 53 85
rect 51 84 52 85
rect 50 84 51 85
rect 49 84 50 85
rect 48 84 49 85
rect 47 84 48 85
rect 46 84 47 85
rect 45 84 46 85
rect 44 84 45 85
rect 43 84 44 85
rect 42 84 43 85
rect 41 84 42 85
rect 40 84 41 85
rect 39 84 40 85
rect 38 84 39 85
rect 37 84 38 85
rect 36 84 37 85
rect 35 84 36 85
rect 34 84 35 85
rect 33 84 34 85
rect 32 84 33 85
rect 31 84 32 85
rect 30 84 31 85
rect 29 84 30 85
rect 28 84 29 85
rect 27 84 28 85
rect 26 84 27 85
rect 25 84 26 85
rect 24 84 25 85
rect 23 84 24 85
rect 22 84 23 85
rect 21 84 22 85
rect 20 84 21 85
rect 19 84 20 85
rect 18 84 19 85
rect 146 85 147 86
rect 145 85 146 86
rect 144 85 145 86
rect 143 85 144 86
rect 142 85 143 86
rect 139 85 140 86
rect 138 85 139 86
rect 137 85 138 86
rect 136 85 137 86
rect 135 85 136 86
rect 134 85 135 86
rect 124 85 125 86
rect 123 85 124 86
rect 122 85 123 86
rect 121 85 122 86
rect 84 85 85 86
rect 83 85 84 86
rect 82 85 83 86
rect 81 85 82 86
rect 80 85 81 86
rect 79 85 80 86
rect 78 85 79 86
rect 77 85 78 86
rect 76 85 77 86
rect 75 85 76 86
rect 74 85 75 86
rect 73 85 74 86
rect 72 85 73 86
rect 71 85 72 86
rect 70 85 71 86
rect 69 85 70 86
rect 68 85 69 86
rect 67 85 68 86
rect 66 85 67 86
rect 65 85 66 86
rect 64 85 65 86
rect 63 85 64 86
rect 62 85 63 86
rect 61 85 62 86
rect 60 85 61 86
rect 59 85 60 86
rect 58 85 59 86
rect 57 85 58 86
rect 56 85 57 86
rect 55 85 56 86
rect 54 85 55 86
rect 53 85 54 86
rect 52 85 53 86
rect 51 85 52 86
rect 50 85 51 86
rect 49 85 50 86
rect 48 85 49 86
rect 47 85 48 86
rect 46 85 47 86
rect 45 85 46 86
rect 44 85 45 86
rect 43 85 44 86
rect 42 85 43 86
rect 41 85 42 86
rect 40 85 41 86
rect 39 85 40 86
rect 38 85 39 86
rect 37 85 38 86
rect 36 85 37 86
rect 35 85 36 86
rect 34 85 35 86
rect 33 85 34 86
rect 32 85 33 86
rect 31 85 32 86
rect 30 85 31 86
rect 29 85 30 86
rect 28 85 29 86
rect 27 85 28 86
rect 26 85 27 86
rect 25 85 26 86
rect 24 85 25 86
rect 23 85 24 86
rect 22 85 23 86
rect 21 85 22 86
rect 20 85 21 86
rect 19 85 20 86
rect 18 85 19 86
rect 146 86 147 87
rect 145 86 146 87
rect 144 86 145 87
rect 143 86 144 87
rect 142 86 143 87
rect 138 86 139 87
rect 137 86 138 87
rect 136 86 137 87
rect 135 86 136 87
rect 134 86 135 87
rect 133 86 134 87
rect 125 86 126 87
rect 124 86 125 87
rect 123 86 124 87
rect 122 86 123 87
rect 121 86 122 87
rect 84 86 85 87
rect 83 86 84 87
rect 82 86 83 87
rect 81 86 82 87
rect 80 86 81 87
rect 79 86 80 87
rect 78 86 79 87
rect 77 86 78 87
rect 76 86 77 87
rect 75 86 76 87
rect 74 86 75 87
rect 73 86 74 87
rect 72 86 73 87
rect 71 86 72 87
rect 70 86 71 87
rect 69 86 70 87
rect 68 86 69 87
rect 67 86 68 87
rect 66 86 67 87
rect 65 86 66 87
rect 64 86 65 87
rect 63 86 64 87
rect 62 86 63 87
rect 61 86 62 87
rect 60 86 61 87
rect 59 86 60 87
rect 58 86 59 87
rect 57 86 58 87
rect 56 86 57 87
rect 55 86 56 87
rect 54 86 55 87
rect 53 86 54 87
rect 52 86 53 87
rect 51 86 52 87
rect 50 86 51 87
rect 49 86 50 87
rect 48 86 49 87
rect 47 86 48 87
rect 46 86 47 87
rect 45 86 46 87
rect 44 86 45 87
rect 43 86 44 87
rect 42 86 43 87
rect 41 86 42 87
rect 40 86 41 87
rect 39 86 40 87
rect 38 86 39 87
rect 37 86 38 87
rect 36 86 37 87
rect 35 86 36 87
rect 34 86 35 87
rect 33 86 34 87
rect 32 86 33 87
rect 31 86 32 87
rect 30 86 31 87
rect 29 86 30 87
rect 28 86 29 87
rect 27 86 28 87
rect 26 86 27 87
rect 25 86 26 87
rect 24 86 25 87
rect 23 86 24 87
rect 22 86 23 87
rect 21 86 22 87
rect 20 86 21 87
rect 19 86 20 87
rect 18 86 19 87
rect 146 87 147 88
rect 145 87 146 88
rect 144 87 145 88
rect 143 87 144 88
rect 142 87 143 88
rect 137 87 138 88
rect 136 87 137 88
rect 135 87 136 88
rect 134 87 135 88
rect 133 87 134 88
rect 132 87 133 88
rect 125 87 126 88
rect 124 87 125 88
rect 123 87 124 88
rect 122 87 123 88
rect 121 87 122 88
rect 84 87 85 88
rect 83 87 84 88
rect 82 87 83 88
rect 81 87 82 88
rect 80 87 81 88
rect 79 87 80 88
rect 78 87 79 88
rect 77 87 78 88
rect 76 87 77 88
rect 75 87 76 88
rect 74 87 75 88
rect 73 87 74 88
rect 72 87 73 88
rect 71 87 72 88
rect 70 87 71 88
rect 69 87 70 88
rect 68 87 69 88
rect 67 87 68 88
rect 66 87 67 88
rect 65 87 66 88
rect 64 87 65 88
rect 63 87 64 88
rect 62 87 63 88
rect 61 87 62 88
rect 60 87 61 88
rect 59 87 60 88
rect 58 87 59 88
rect 57 87 58 88
rect 56 87 57 88
rect 55 87 56 88
rect 54 87 55 88
rect 53 87 54 88
rect 52 87 53 88
rect 51 87 52 88
rect 50 87 51 88
rect 49 87 50 88
rect 48 87 49 88
rect 47 87 48 88
rect 46 87 47 88
rect 45 87 46 88
rect 44 87 45 88
rect 43 87 44 88
rect 42 87 43 88
rect 41 87 42 88
rect 40 87 41 88
rect 39 87 40 88
rect 38 87 39 88
rect 37 87 38 88
rect 36 87 37 88
rect 35 87 36 88
rect 34 87 35 88
rect 33 87 34 88
rect 32 87 33 88
rect 31 87 32 88
rect 30 87 31 88
rect 29 87 30 88
rect 28 87 29 88
rect 27 87 28 88
rect 26 87 27 88
rect 25 87 26 88
rect 24 87 25 88
rect 23 87 24 88
rect 22 87 23 88
rect 21 87 22 88
rect 20 87 21 88
rect 19 87 20 88
rect 18 87 19 88
rect 146 88 147 89
rect 145 88 146 89
rect 144 88 145 89
rect 143 88 144 89
rect 142 88 143 89
rect 137 88 138 89
rect 136 88 137 89
rect 135 88 136 89
rect 134 88 135 89
rect 133 88 134 89
rect 132 88 133 89
rect 131 88 132 89
rect 126 88 127 89
rect 125 88 126 89
rect 124 88 125 89
rect 123 88 124 89
rect 122 88 123 89
rect 121 88 122 89
rect 84 88 85 89
rect 83 88 84 89
rect 82 88 83 89
rect 81 88 82 89
rect 80 88 81 89
rect 79 88 80 89
rect 78 88 79 89
rect 77 88 78 89
rect 76 88 77 89
rect 75 88 76 89
rect 74 88 75 89
rect 73 88 74 89
rect 72 88 73 89
rect 71 88 72 89
rect 70 88 71 89
rect 69 88 70 89
rect 68 88 69 89
rect 67 88 68 89
rect 66 88 67 89
rect 65 88 66 89
rect 64 88 65 89
rect 63 88 64 89
rect 62 88 63 89
rect 61 88 62 89
rect 60 88 61 89
rect 59 88 60 89
rect 58 88 59 89
rect 57 88 58 89
rect 56 88 57 89
rect 55 88 56 89
rect 54 88 55 89
rect 53 88 54 89
rect 52 88 53 89
rect 51 88 52 89
rect 50 88 51 89
rect 49 88 50 89
rect 48 88 49 89
rect 47 88 48 89
rect 46 88 47 89
rect 45 88 46 89
rect 44 88 45 89
rect 43 88 44 89
rect 42 88 43 89
rect 41 88 42 89
rect 40 88 41 89
rect 39 88 40 89
rect 38 88 39 89
rect 37 88 38 89
rect 36 88 37 89
rect 35 88 36 89
rect 34 88 35 89
rect 33 88 34 89
rect 32 88 33 89
rect 31 88 32 89
rect 30 88 31 89
rect 29 88 30 89
rect 28 88 29 89
rect 27 88 28 89
rect 26 88 27 89
rect 25 88 26 89
rect 24 88 25 89
rect 23 88 24 89
rect 22 88 23 89
rect 21 88 22 89
rect 20 88 21 89
rect 19 88 20 89
rect 18 88 19 89
rect 146 89 147 90
rect 145 89 146 90
rect 144 89 145 90
rect 143 89 144 90
rect 142 89 143 90
rect 136 89 137 90
rect 135 89 136 90
rect 134 89 135 90
rect 133 89 134 90
rect 132 89 133 90
rect 131 89 132 90
rect 130 89 131 90
rect 129 89 130 90
rect 128 89 129 90
rect 127 89 128 90
rect 126 89 127 90
rect 125 89 126 90
rect 124 89 125 90
rect 123 89 124 90
rect 122 89 123 90
rect 121 89 122 90
rect 84 89 85 90
rect 83 89 84 90
rect 82 89 83 90
rect 81 89 82 90
rect 80 89 81 90
rect 79 89 80 90
rect 78 89 79 90
rect 77 89 78 90
rect 76 89 77 90
rect 75 89 76 90
rect 74 89 75 90
rect 73 89 74 90
rect 72 89 73 90
rect 71 89 72 90
rect 70 89 71 90
rect 69 89 70 90
rect 68 89 69 90
rect 67 89 68 90
rect 66 89 67 90
rect 65 89 66 90
rect 64 89 65 90
rect 63 89 64 90
rect 62 89 63 90
rect 61 89 62 90
rect 60 89 61 90
rect 59 89 60 90
rect 58 89 59 90
rect 57 89 58 90
rect 56 89 57 90
rect 55 89 56 90
rect 54 89 55 90
rect 53 89 54 90
rect 52 89 53 90
rect 51 89 52 90
rect 50 89 51 90
rect 49 89 50 90
rect 48 89 49 90
rect 47 89 48 90
rect 46 89 47 90
rect 45 89 46 90
rect 44 89 45 90
rect 43 89 44 90
rect 42 89 43 90
rect 41 89 42 90
rect 40 89 41 90
rect 39 89 40 90
rect 38 89 39 90
rect 37 89 38 90
rect 36 89 37 90
rect 35 89 36 90
rect 34 89 35 90
rect 33 89 34 90
rect 32 89 33 90
rect 31 89 32 90
rect 30 89 31 90
rect 29 89 30 90
rect 28 89 29 90
rect 27 89 28 90
rect 26 89 27 90
rect 25 89 26 90
rect 24 89 25 90
rect 23 89 24 90
rect 22 89 23 90
rect 21 89 22 90
rect 20 89 21 90
rect 19 89 20 90
rect 18 89 19 90
rect 146 90 147 91
rect 145 90 146 91
rect 144 90 145 91
rect 143 90 144 91
rect 142 90 143 91
rect 135 90 136 91
rect 134 90 135 91
rect 133 90 134 91
rect 132 90 133 91
rect 131 90 132 91
rect 130 90 131 91
rect 129 90 130 91
rect 128 90 129 91
rect 127 90 128 91
rect 126 90 127 91
rect 125 90 126 91
rect 124 90 125 91
rect 123 90 124 91
rect 122 90 123 91
rect 84 90 85 91
rect 83 90 84 91
rect 82 90 83 91
rect 81 90 82 91
rect 80 90 81 91
rect 79 90 80 91
rect 78 90 79 91
rect 77 90 78 91
rect 76 90 77 91
rect 75 90 76 91
rect 74 90 75 91
rect 73 90 74 91
rect 72 90 73 91
rect 71 90 72 91
rect 70 90 71 91
rect 69 90 70 91
rect 68 90 69 91
rect 67 90 68 91
rect 66 90 67 91
rect 65 90 66 91
rect 64 90 65 91
rect 63 90 64 91
rect 62 90 63 91
rect 61 90 62 91
rect 60 90 61 91
rect 59 90 60 91
rect 58 90 59 91
rect 57 90 58 91
rect 56 90 57 91
rect 55 90 56 91
rect 54 90 55 91
rect 53 90 54 91
rect 52 90 53 91
rect 51 90 52 91
rect 50 90 51 91
rect 49 90 50 91
rect 48 90 49 91
rect 47 90 48 91
rect 46 90 47 91
rect 45 90 46 91
rect 44 90 45 91
rect 43 90 44 91
rect 42 90 43 91
rect 41 90 42 91
rect 40 90 41 91
rect 39 90 40 91
rect 38 90 39 91
rect 37 90 38 91
rect 36 90 37 91
rect 35 90 36 91
rect 34 90 35 91
rect 33 90 34 91
rect 32 90 33 91
rect 31 90 32 91
rect 30 90 31 91
rect 29 90 30 91
rect 28 90 29 91
rect 27 90 28 91
rect 26 90 27 91
rect 25 90 26 91
rect 24 90 25 91
rect 23 90 24 91
rect 22 90 23 91
rect 21 90 22 91
rect 20 90 21 91
rect 19 90 20 91
rect 18 90 19 91
rect 146 91 147 92
rect 145 91 146 92
rect 144 91 145 92
rect 143 91 144 92
rect 142 91 143 92
rect 134 91 135 92
rect 133 91 134 92
rect 132 91 133 92
rect 131 91 132 92
rect 130 91 131 92
rect 129 91 130 92
rect 128 91 129 92
rect 127 91 128 92
rect 126 91 127 92
rect 125 91 126 92
rect 124 91 125 92
rect 123 91 124 92
rect 122 91 123 92
rect 84 91 85 92
rect 83 91 84 92
rect 82 91 83 92
rect 81 91 82 92
rect 80 91 81 92
rect 79 91 80 92
rect 78 91 79 92
rect 77 91 78 92
rect 76 91 77 92
rect 75 91 76 92
rect 74 91 75 92
rect 73 91 74 92
rect 72 91 73 92
rect 71 91 72 92
rect 70 91 71 92
rect 69 91 70 92
rect 68 91 69 92
rect 67 91 68 92
rect 66 91 67 92
rect 65 91 66 92
rect 64 91 65 92
rect 63 91 64 92
rect 62 91 63 92
rect 61 91 62 92
rect 60 91 61 92
rect 59 91 60 92
rect 58 91 59 92
rect 57 91 58 92
rect 56 91 57 92
rect 55 91 56 92
rect 54 91 55 92
rect 53 91 54 92
rect 52 91 53 92
rect 51 91 52 92
rect 50 91 51 92
rect 49 91 50 92
rect 48 91 49 92
rect 47 91 48 92
rect 46 91 47 92
rect 45 91 46 92
rect 44 91 45 92
rect 43 91 44 92
rect 42 91 43 92
rect 41 91 42 92
rect 40 91 41 92
rect 39 91 40 92
rect 38 91 39 92
rect 37 91 38 92
rect 36 91 37 92
rect 35 91 36 92
rect 34 91 35 92
rect 33 91 34 92
rect 32 91 33 92
rect 31 91 32 92
rect 30 91 31 92
rect 29 91 30 92
rect 28 91 29 92
rect 27 91 28 92
rect 26 91 27 92
rect 25 91 26 92
rect 24 91 25 92
rect 23 91 24 92
rect 22 91 23 92
rect 21 91 22 92
rect 20 91 21 92
rect 19 91 20 92
rect 18 91 19 92
rect 146 92 147 93
rect 145 92 146 93
rect 144 92 145 93
rect 143 92 144 93
rect 142 92 143 93
rect 133 92 134 93
rect 132 92 133 93
rect 131 92 132 93
rect 130 92 131 93
rect 129 92 130 93
rect 128 92 129 93
rect 127 92 128 93
rect 126 92 127 93
rect 125 92 126 93
rect 124 92 125 93
rect 123 92 124 93
rect 84 92 85 93
rect 83 92 84 93
rect 82 92 83 93
rect 81 92 82 93
rect 80 92 81 93
rect 79 92 80 93
rect 78 92 79 93
rect 77 92 78 93
rect 76 92 77 93
rect 75 92 76 93
rect 74 92 75 93
rect 73 92 74 93
rect 72 92 73 93
rect 71 92 72 93
rect 70 92 71 93
rect 69 92 70 93
rect 68 92 69 93
rect 67 92 68 93
rect 66 92 67 93
rect 65 92 66 93
rect 64 92 65 93
rect 63 92 64 93
rect 62 92 63 93
rect 61 92 62 93
rect 60 92 61 93
rect 59 92 60 93
rect 58 92 59 93
rect 57 92 58 93
rect 56 92 57 93
rect 55 92 56 93
rect 54 92 55 93
rect 53 92 54 93
rect 52 92 53 93
rect 51 92 52 93
rect 50 92 51 93
rect 49 92 50 93
rect 48 92 49 93
rect 47 92 48 93
rect 46 92 47 93
rect 45 92 46 93
rect 44 92 45 93
rect 43 92 44 93
rect 42 92 43 93
rect 41 92 42 93
rect 40 92 41 93
rect 39 92 40 93
rect 38 92 39 93
rect 37 92 38 93
rect 36 92 37 93
rect 35 92 36 93
rect 34 92 35 93
rect 33 92 34 93
rect 32 92 33 93
rect 31 92 32 93
rect 30 92 31 93
rect 29 92 30 93
rect 28 92 29 93
rect 27 92 28 93
rect 26 92 27 93
rect 25 92 26 93
rect 24 92 25 93
rect 23 92 24 93
rect 22 92 23 93
rect 21 92 22 93
rect 20 92 21 93
rect 19 92 20 93
rect 18 92 19 93
rect 146 93 147 94
rect 145 93 146 94
rect 144 93 145 94
rect 143 93 144 94
rect 142 93 143 94
rect 132 93 133 94
rect 131 93 132 94
rect 130 93 131 94
rect 129 93 130 94
rect 128 93 129 94
rect 127 93 128 94
rect 126 93 127 94
rect 125 93 126 94
rect 124 93 125 94
rect 84 93 85 94
rect 83 93 84 94
rect 82 93 83 94
rect 81 93 82 94
rect 80 93 81 94
rect 79 93 80 94
rect 78 93 79 94
rect 77 93 78 94
rect 76 93 77 94
rect 75 93 76 94
rect 74 93 75 94
rect 73 93 74 94
rect 72 93 73 94
rect 71 93 72 94
rect 70 93 71 94
rect 69 93 70 94
rect 68 93 69 94
rect 67 93 68 94
rect 66 93 67 94
rect 65 93 66 94
rect 64 93 65 94
rect 63 93 64 94
rect 62 93 63 94
rect 61 93 62 94
rect 60 93 61 94
rect 59 93 60 94
rect 58 93 59 94
rect 57 93 58 94
rect 56 93 57 94
rect 55 93 56 94
rect 54 93 55 94
rect 53 93 54 94
rect 52 93 53 94
rect 51 93 52 94
rect 50 93 51 94
rect 49 93 50 94
rect 48 93 49 94
rect 47 93 48 94
rect 46 93 47 94
rect 45 93 46 94
rect 44 93 45 94
rect 43 93 44 94
rect 42 93 43 94
rect 41 93 42 94
rect 40 93 41 94
rect 39 93 40 94
rect 38 93 39 94
rect 37 93 38 94
rect 36 93 37 94
rect 35 93 36 94
rect 34 93 35 94
rect 33 93 34 94
rect 32 93 33 94
rect 31 93 32 94
rect 30 93 31 94
rect 29 93 30 94
rect 28 93 29 94
rect 27 93 28 94
rect 26 93 27 94
rect 25 93 26 94
rect 24 93 25 94
rect 23 93 24 94
rect 22 93 23 94
rect 21 93 22 94
rect 20 93 21 94
rect 19 93 20 94
rect 18 93 19 94
rect 146 94 147 95
rect 145 94 146 95
rect 144 94 145 95
rect 143 94 144 95
rect 142 94 143 95
rect 129 94 130 95
rect 128 94 129 95
rect 127 94 128 95
rect 84 94 85 95
rect 83 94 84 95
rect 82 94 83 95
rect 81 94 82 95
rect 80 94 81 95
rect 79 94 80 95
rect 78 94 79 95
rect 77 94 78 95
rect 76 94 77 95
rect 75 94 76 95
rect 74 94 75 95
rect 73 94 74 95
rect 72 94 73 95
rect 71 94 72 95
rect 70 94 71 95
rect 69 94 70 95
rect 68 94 69 95
rect 67 94 68 95
rect 66 94 67 95
rect 65 94 66 95
rect 64 94 65 95
rect 63 94 64 95
rect 62 94 63 95
rect 61 94 62 95
rect 60 94 61 95
rect 59 94 60 95
rect 58 94 59 95
rect 57 94 58 95
rect 56 94 57 95
rect 55 94 56 95
rect 54 94 55 95
rect 53 94 54 95
rect 52 94 53 95
rect 51 94 52 95
rect 50 94 51 95
rect 49 94 50 95
rect 48 94 49 95
rect 47 94 48 95
rect 46 94 47 95
rect 45 94 46 95
rect 44 94 45 95
rect 43 94 44 95
rect 42 94 43 95
rect 41 94 42 95
rect 40 94 41 95
rect 39 94 40 95
rect 38 94 39 95
rect 37 94 38 95
rect 36 94 37 95
rect 35 94 36 95
rect 34 94 35 95
rect 33 94 34 95
rect 32 94 33 95
rect 31 94 32 95
rect 30 94 31 95
rect 29 94 30 95
rect 28 94 29 95
rect 27 94 28 95
rect 26 94 27 95
rect 25 94 26 95
rect 24 94 25 95
rect 23 94 24 95
rect 22 94 23 95
rect 21 94 22 95
rect 20 94 21 95
rect 19 94 20 95
rect 18 94 19 95
rect 84 95 85 96
rect 83 95 84 96
rect 82 95 83 96
rect 81 95 82 96
rect 80 95 81 96
rect 79 95 80 96
rect 78 95 79 96
rect 77 95 78 96
rect 76 95 77 96
rect 75 95 76 96
rect 74 95 75 96
rect 73 95 74 96
rect 72 95 73 96
rect 71 95 72 96
rect 70 95 71 96
rect 69 95 70 96
rect 68 95 69 96
rect 67 95 68 96
rect 66 95 67 96
rect 65 95 66 96
rect 64 95 65 96
rect 63 95 64 96
rect 62 95 63 96
rect 61 95 62 96
rect 60 95 61 96
rect 59 95 60 96
rect 58 95 59 96
rect 57 95 58 96
rect 56 95 57 96
rect 55 95 56 96
rect 54 95 55 96
rect 53 95 54 96
rect 52 95 53 96
rect 51 95 52 96
rect 50 95 51 96
rect 49 95 50 96
rect 48 95 49 96
rect 47 95 48 96
rect 46 95 47 96
rect 45 95 46 96
rect 44 95 45 96
rect 43 95 44 96
rect 42 95 43 96
rect 41 95 42 96
rect 40 95 41 96
rect 39 95 40 96
rect 38 95 39 96
rect 37 95 38 96
rect 36 95 37 96
rect 35 95 36 96
rect 34 95 35 96
rect 33 95 34 96
rect 32 95 33 96
rect 31 95 32 96
rect 30 95 31 96
rect 29 95 30 96
rect 28 95 29 96
rect 27 95 28 96
rect 26 95 27 96
rect 25 95 26 96
rect 24 95 25 96
rect 23 95 24 96
rect 22 95 23 96
rect 21 95 22 96
rect 20 95 21 96
rect 19 95 20 96
rect 18 95 19 96
rect 84 96 85 97
rect 83 96 84 97
rect 82 96 83 97
rect 81 96 82 97
rect 80 96 81 97
rect 79 96 80 97
rect 78 96 79 97
rect 77 96 78 97
rect 76 96 77 97
rect 75 96 76 97
rect 74 96 75 97
rect 73 96 74 97
rect 72 96 73 97
rect 71 96 72 97
rect 70 96 71 97
rect 69 96 70 97
rect 68 96 69 97
rect 67 96 68 97
rect 66 96 67 97
rect 65 96 66 97
rect 64 96 65 97
rect 63 96 64 97
rect 62 96 63 97
rect 61 96 62 97
rect 60 96 61 97
rect 59 96 60 97
rect 58 96 59 97
rect 57 96 58 97
rect 56 96 57 97
rect 55 96 56 97
rect 54 96 55 97
rect 53 96 54 97
rect 52 96 53 97
rect 51 96 52 97
rect 50 96 51 97
rect 49 96 50 97
rect 48 96 49 97
rect 47 96 48 97
rect 46 96 47 97
rect 45 96 46 97
rect 44 96 45 97
rect 43 96 44 97
rect 42 96 43 97
rect 41 96 42 97
rect 40 96 41 97
rect 39 96 40 97
rect 38 96 39 97
rect 37 96 38 97
rect 36 96 37 97
rect 35 96 36 97
rect 34 96 35 97
rect 33 96 34 97
rect 32 96 33 97
rect 31 96 32 97
rect 30 96 31 97
rect 29 96 30 97
rect 28 96 29 97
rect 27 96 28 97
rect 26 96 27 97
rect 25 96 26 97
rect 24 96 25 97
rect 23 96 24 97
rect 22 96 23 97
rect 21 96 22 97
rect 20 96 21 97
rect 19 96 20 97
rect 18 96 19 97
rect 84 97 85 98
rect 83 97 84 98
rect 82 97 83 98
rect 81 97 82 98
rect 80 97 81 98
rect 79 97 80 98
rect 78 97 79 98
rect 77 97 78 98
rect 76 97 77 98
rect 75 97 76 98
rect 74 97 75 98
rect 73 97 74 98
rect 72 97 73 98
rect 71 97 72 98
rect 70 97 71 98
rect 69 97 70 98
rect 68 97 69 98
rect 67 97 68 98
rect 66 97 67 98
rect 65 97 66 98
rect 64 97 65 98
rect 63 97 64 98
rect 62 97 63 98
rect 61 97 62 98
rect 60 97 61 98
rect 59 97 60 98
rect 58 97 59 98
rect 57 97 58 98
rect 56 97 57 98
rect 55 97 56 98
rect 54 97 55 98
rect 53 97 54 98
rect 52 97 53 98
rect 51 97 52 98
rect 50 97 51 98
rect 49 97 50 98
rect 48 97 49 98
rect 47 97 48 98
rect 46 97 47 98
rect 45 97 46 98
rect 44 97 45 98
rect 43 97 44 98
rect 42 97 43 98
rect 41 97 42 98
rect 40 97 41 98
rect 39 97 40 98
rect 38 97 39 98
rect 37 97 38 98
rect 36 97 37 98
rect 35 97 36 98
rect 34 97 35 98
rect 33 97 34 98
rect 32 97 33 98
rect 31 97 32 98
rect 30 97 31 98
rect 29 97 30 98
rect 28 97 29 98
rect 27 97 28 98
rect 26 97 27 98
rect 25 97 26 98
rect 24 97 25 98
rect 23 97 24 98
rect 22 97 23 98
rect 21 97 22 98
rect 20 97 21 98
rect 19 97 20 98
rect 18 97 19 98
rect 141 98 142 99
rect 140 98 141 99
rect 139 98 140 99
rect 138 98 139 99
rect 137 98 138 99
rect 84 98 85 99
rect 83 98 84 99
rect 82 98 83 99
rect 81 98 82 99
rect 80 98 81 99
rect 79 98 80 99
rect 78 98 79 99
rect 77 98 78 99
rect 76 98 77 99
rect 75 98 76 99
rect 74 98 75 99
rect 73 98 74 99
rect 72 98 73 99
rect 71 98 72 99
rect 70 98 71 99
rect 69 98 70 99
rect 68 98 69 99
rect 67 98 68 99
rect 66 98 67 99
rect 65 98 66 99
rect 64 98 65 99
rect 63 98 64 99
rect 62 98 63 99
rect 61 98 62 99
rect 60 98 61 99
rect 59 98 60 99
rect 58 98 59 99
rect 57 98 58 99
rect 56 98 57 99
rect 55 98 56 99
rect 54 98 55 99
rect 53 98 54 99
rect 52 98 53 99
rect 51 98 52 99
rect 50 98 51 99
rect 49 98 50 99
rect 48 98 49 99
rect 47 98 48 99
rect 46 98 47 99
rect 45 98 46 99
rect 44 98 45 99
rect 43 98 44 99
rect 42 98 43 99
rect 41 98 42 99
rect 40 98 41 99
rect 39 98 40 99
rect 38 98 39 99
rect 37 98 38 99
rect 36 98 37 99
rect 35 98 36 99
rect 34 98 35 99
rect 33 98 34 99
rect 32 98 33 99
rect 31 98 32 99
rect 30 98 31 99
rect 29 98 30 99
rect 28 98 29 99
rect 27 98 28 99
rect 26 98 27 99
rect 25 98 26 99
rect 24 98 25 99
rect 23 98 24 99
rect 22 98 23 99
rect 21 98 22 99
rect 20 98 21 99
rect 19 98 20 99
rect 18 98 19 99
rect 141 99 142 100
rect 140 99 141 100
rect 139 99 140 100
rect 138 99 139 100
rect 137 99 138 100
rect 136 99 137 100
rect 84 99 85 100
rect 83 99 84 100
rect 82 99 83 100
rect 81 99 82 100
rect 80 99 81 100
rect 79 99 80 100
rect 78 99 79 100
rect 77 99 78 100
rect 76 99 77 100
rect 75 99 76 100
rect 74 99 75 100
rect 73 99 74 100
rect 72 99 73 100
rect 71 99 72 100
rect 70 99 71 100
rect 69 99 70 100
rect 68 99 69 100
rect 67 99 68 100
rect 66 99 67 100
rect 65 99 66 100
rect 64 99 65 100
rect 63 99 64 100
rect 62 99 63 100
rect 61 99 62 100
rect 60 99 61 100
rect 59 99 60 100
rect 58 99 59 100
rect 57 99 58 100
rect 56 99 57 100
rect 55 99 56 100
rect 54 99 55 100
rect 53 99 54 100
rect 52 99 53 100
rect 51 99 52 100
rect 50 99 51 100
rect 49 99 50 100
rect 48 99 49 100
rect 47 99 48 100
rect 46 99 47 100
rect 45 99 46 100
rect 44 99 45 100
rect 43 99 44 100
rect 42 99 43 100
rect 41 99 42 100
rect 40 99 41 100
rect 39 99 40 100
rect 38 99 39 100
rect 37 99 38 100
rect 36 99 37 100
rect 35 99 36 100
rect 34 99 35 100
rect 33 99 34 100
rect 32 99 33 100
rect 31 99 32 100
rect 30 99 31 100
rect 29 99 30 100
rect 28 99 29 100
rect 27 99 28 100
rect 26 99 27 100
rect 25 99 26 100
rect 24 99 25 100
rect 23 99 24 100
rect 22 99 23 100
rect 21 99 22 100
rect 20 99 21 100
rect 19 99 20 100
rect 18 99 19 100
rect 141 100 142 101
rect 140 100 141 101
rect 139 100 140 101
rect 138 100 139 101
rect 137 100 138 101
rect 136 100 137 101
rect 135 100 136 101
rect 62 100 63 101
rect 61 100 62 101
rect 60 100 61 101
rect 59 100 60 101
rect 58 100 59 101
rect 57 100 58 101
rect 56 100 57 101
rect 55 100 56 101
rect 54 100 55 101
rect 53 100 54 101
rect 52 100 53 101
rect 51 100 52 101
rect 50 100 51 101
rect 49 100 50 101
rect 31 100 32 101
rect 30 100 31 101
rect 29 100 30 101
rect 28 100 29 101
rect 27 100 28 101
rect 26 100 27 101
rect 25 100 26 101
rect 24 100 25 101
rect 23 100 24 101
rect 22 100 23 101
rect 21 100 22 101
rect 20 100 21 101
rect 19 100 20 101
rect 18 100 19 101
rect 141 101 142 102
rect 140 101 141 102
rect 139 101 140 102
rect 138 101 139 102
rect 137 101 138 102
rect 136 101 137 102
rect 135 101 136 102
rect 134 101 135 102
rect 62 101 63 102
rect 61 101 62 102
rect 60 101 61 102
rect 59 101 60 102
rect 58 101 59 102
rect 57 101 58 102
rect 56 101 57 102
rect 55 101 56 102
rect 54 101 55 102
rect 53 101 54 102
rect 52 101 53 102
rect 51 101 52 102
rect 50 101 51 102
rect 49 101 50 102
rect 31 101 32 102
rect 30 101 31 102
rect 29 101 30 102
rect 28 101 29 102
rect 27 101 28 102
rect 26 101 27 102
rect 25 101 26 102
rect 24 101 25 102
rect 23 101 24 102
rect 22 101 23 102
rect 21 101 22 102
rect 20 101 21 102
rect 19 101 20 102
rect 18 101 19 102
rect 141 102 142 103
rect 140 102 141 103
rect 139 102 140 103
rect 138 102 139 103
rect 137 102 138 103
rect 136 102 137 103
rect 135 102 136 103
rect 134 102 135 103
rect 133 102 134 103
rect 132 102 133 103
rect 62 102 63 103
rect 61 102 62 103
rect 60 102 61 103
rect 59 102 60 103
rect 58 102 59 103
rect 57 102 58 103
rect 56 102 57 103
rect 55 102 56 103
rect 54 102 55 103
rect 53 102 54 103
rect 52 102 53 103
rect 51 102 52 103
rect 50 102 51 103
rect 49 102 50 103
rect 31 102 32 103
rect 30 102 31 103
rect 29 102 30 103
rect 28 102 29 103
rect 27 102 28 103
rect 26 102 27 103
rect 25 102 26 103
rect 24 102 25 103
rect 23 102 24 103
rect 22 102 23 103
rect 21 102 22 103
rect 20 102 21 103
rect 19 102 20 103
rect 18 102 19 103
rect 141 103 142 104
rect 140 103 141 104
rect 139 103 140 104
rect 138 103 139 104
rect 137 103 138 104
rect 136 103 137 104
rect 135 103 136 104
rect 134 103 135 104
rect 133 103 134 104
rect 132 103 133 104
rect 131 103 132 104
rect 62 103 63 104
rect 61 103 62 104
rect 60 103 61 104
rect 59 103 60 104
rect 58 103 59 104
rect 57 103 58 104
rect 56 103 57 104
rect 55 103 56 104
rect 54 103 55 104
rect 53 103 54 104
rect 52 103 53 104
rect 51 103 52 104
rect 50 103 51 104
rect 49 103 50 104
rect 31 103 32 104
rect 30 103 31 104
rect 29 103 30 104
rect 28 103 29 104
rect 27 103 28 104
rect 26 103 27 104
rect 25 103 26 104
rect 24 103 25 104
rect 23 103 24 104
rect 22 103 23 104
rect 21 103 22 104
rect 20 103 21 104
rect 19 103 20 104
rect 18 103 19 104
rect 141 104 142 105
rect 140 104 141 105
rect 139 104 140 105
rect 138 104 139 105
rect 135 104 136 105
rect 134 104 135 105
rect 133 104 134 105
rect 132 104 133 105
rect 131 104 132 105
rect 130 104 131 105
rect 129 104 130 105
rect 62 104 63 105
rect 61 104 62 105
rect 60 104 61 105
rect 59 104 60 105
rect 58 104 59 105
rect 57 104 58 105
rect 56 104 57 105
rect 55 104 56 105
rect 54 104 55 105
rect 53 104 54 105
rect 52 104 53 105
rect 51 104 52 105
rect 50 104 51 105
rect 49 104 50 105
rect 31 104 32 105
rect 30 104 31 105
rect 29 104 30 105
rect 28 104 29 105
rect 27 104 28 105
rect 26 104 27 105
rect 25 104 26 105
rect 24 104 25 105
rect 23 104 24 105
rect 22 104 23 105
rect 21 104 22 105
rect 20 104 21 105
rect 19 104 20 105
rect 18 104 19 105
rect 141 105 142 106
rect 140 105 141 106
rect 139 105 140 106
rect 138 105 139 106
rect 134 105 135 106
rect 133 105 134 106
rect 132 105 133 106
rect 131 105 132 106
rect 130 105 131 106
rect 129 105 130 106
rect 128 105 129 106
rect 62 105 63 106
rect 61 105 62 106
rect 60 105 61 106
rect 59 105 60 106
rect 58 105 59 106
rect 57 105 58 106
rect 56 105 57 106
rect 55 105 56 106
rect 54 105 55 106
rect 53 105 54 106
rect 52 105 53 106
rect 51 105 52 106
rect 50 105 51 106
rect 49 105 50 106
rect 31 105 32 106
rect 30 105 31 106
rect 29 105 30 106
rect 28 105 29 106
rect 27 105 28 106
rect 26 105 27 106
rect 25 105 26 106
rect 24 105 25 106
rect 23 105 24 106
rect 22 105 23 106
rect 21 105 22 106
rect 20 105 21 106
rect 19 105 20 106
rect 18 105 19 106
rect 141 106 142 107
rect 140 106 141 107
rect 139 106 140 107
rect 138 106 139 107
rect 132 106 133 107
rect 131 106 132 107
rect 130 106 131 107
rect 129 106 130 107
rect 128 106 129 107
rect 127 106 128 107
rect 126 106 127 107
rect 62 106 63 107
rect 61 106 62 107
rect 60 106 61 107
rect 59 106 60 107
rect 58 106 59 107
rect 57 106 58 107
rect 56 106 57 107
rect 55 106 56 107
rect 54 106 55 107
rect 53 106 54 107
rect 52 106 53 107
rect 51 106 52 107
rect 50 106 51 107
rect 49 106 50 107
rect 31 106 32 107
rect 30 106 31 107
rect 29 106 30 107
rect 28 106 29 107
rect 27 106 28 107
rect 26 106 27 107
rect 25 106 26 107
rect 24 106 25 107
rect 23 106 24 107
rect 22 106 23 107
rect 21 106 22 107
rect 20 106 21 107
rect 19 106 20 107
rect 18 106 19 107
rect 141 107 142 108
rect 140 107 141 108
rect 139 107 140 108
rect 138 107 139 108
rect 131 107 132 108
rect 130 107 131 108
rect 129 107 130 108
rect 128 107 129 108
rect 127 107 128 108
rect 126 107 127 108
rect 125 107 126 108
rect 62 107 63 108
rect 61 107 62 108
rect 60 107 61 108
rect 59 107 60 108
rect 58 107 59 108
rect 57 107 58 108
rect 56 107 57 108
rect 55 107 56 108
rect 54 107 55 108
rect 53 107 54 108
rect 52 107 53 108
rect 51 107 52 108
rect 50 107 51 108
rect 49 107 50 108
rect 31 107 32 108
rect 30 107 31 108
rect 29 107 30 108
rect 28 107 29 108
rect 27 107 28 108
rect 26 107 27 108
rect 25 107 26 108
rect 24 107 25 108
rect 23 107 24 108
rect 22 107 23 108
rect 21 107 22 108
rect 20 107 21 108
rect 19 107 20 108
rect 18 107 19 108
rect 141 108 142 109
rect 140 108 141 109
rect 139 108 140 109
rect 138 108 139 109
rect 129 108 130 109
rect 128 108 129 109
rect 127 108 128 109
rect 126 108 127 109
rect 125 108 126 109
rect 124 108 125 109
rect 123 108 124 109
rect 62 108 63 109
rect 61 108 62 109
rect 60 108 61 109
rect 59 108 60 109
rect 58 108 59 109
rect 57 108 58 109
rect 56 108 57 109
rect 55 108 56 109
rect 54 108 55 109
rect 53 108 54 109
rect 52 108 53 109
rect 51 108 52 109
rect 50 108 51 109
rect 49 108 50 109
rect 32 108 33 109
rect 31 108 32 109
rect 30 108 31 109
rect 29 108 30 109
rect 28 108 29 109
rect 27 108 28 109
rect 26 108 27 109
rect 25 108 26 109
rect 24 108 25 109
rect 23 108 24 109
rect 22 108 23 109
rect 21 108 22 109
rect 20 108 21 109
rect 19 108 20 109
rect 18 108 19 109
rect 141 109 142 110
rect 140 109 141 110
rect 139 109 140 110
rect 138 109 139 110
rect 137 109 138 110
rect 128 109 129 110
rect 127 109 128 110
rect 126 109 127 110
rect 125 109 126 110
rect 124 109 125 110
rect 123 109 124 110
rect 122 109 123 110
rect 121 109 122 110
rect 62 109 63 110
rect 61 109 62 110
rect 60 109 61 110
rect 59 109 60 110
rect 58 109 59 110
rect 57 109 58 110
rect 56 109 57 110
rect 55 109 56 110
rect 54 109 55 110
rect 53 109 54 110
rect 52 109 53 110
rect 51 109 52 110
rect 50 109 51 110
rect 49 109 50 110
rect 48 109 49 110
rect 32 109 33 110
rect 31 109 32 110
rect 30 109 31 110
rect 29 109 30 110
rect 28 109 29 110
rect 27 109 28 110
rect 26 109 27 110
rect 25 109 26 110
rect 24 109 25 110
rect 23 109 24 110
rect 22 109 23 110
rect 21 109 22 110
rect 20 109 21 110
rect 19 109 20 110
rect 18 109 19 110
rect 146 110 147 111
rect 145 110 146 111
rect 144 110 145 111
rect 143 110 144 111
rect 142 110 143 111
rect 141 110 142 111
rect 140 110 141 111
rect 139 110 140 111
rect 138 110 139 111
rect 137 110 138 111
rect 136 110 137 111
rect 135 110 136 111
rect 134 110 135 111
rect 133 110 134 111
rect 132 110 133 111
rect 131 110 132 111
rect 130 110 131 111
rect 129 110 130 111
rect 128 110 129 111
rect 127 110 128 111
rect 126 110 127 111
rect 125 110 126 111
rect 124 110 125 111
rect 123 110 124 111
rect 122 110 123 111
rect 121 110 122 111
rect 62 110 63 111
rect 61 110 62 111
rect 60 110 61 111
rect 59 110 60 111
rect 58 110 59 111
rect 57 110 58 111
rect 56 110 57 111
rect 55 110 56 111
rect 54 110 55 111
rect 53 110 54 111
rect 52 110 53 111
rect 51 110 52 111
rect 50 110 51 111
rect 49 110 50 111
rect 48 110 49 111
rect 33 110 34 111
rect 32 110 33 111
rect 31 110 32 111
rect 30 110 31 111
rect 29 110 30 111
rect 28 110 29 111
rect 27 110 28 111
rect 26 110 27 111
rect 25 110 26 111
rect 24 110 25 111
rect 23 110 24 111
rect 22 110 23 111
rect 21 110 22 111
rect 20 110 21 111
rect 19 110 20 111
rect 18 110 19 111
rect 146 111 147 112
rect 145 111 146 112
rect 144 111 145 112
rect 143 111 144 112
rect 142 111 143 112
rect 141 111 142 112
rect 140 111 141 112
rect 139 111 140 112
rect 138 111 139 112
rect 137 111 138 112
rect 136 111 137 112
rect 135 111 136 112
rect 134 111 135 112
rect 133 111 134 112
rect 132 111 133 112
rect 131 111 132 112
rect 130 111 131 112
rect 129 111 130 112
rect 128 111 129 112
rect 127 111 128 112
rect 126 111 127 112
rect 125 111 126 112
rect 124 111 125 112
rect 123 111 124 112
rect 122 111 123 112
rect 121 111 122 112
rect 62 111 63 112
rect 61 111 62 112
rect 60 111 61 112
rect 59 111 60 112
rect 58 111 59 112
rect 57 111 58 112
rect 56 111 57 112
rect 55 111 56 112
rect 54 111 55 112
rect 53 111 54 112
rect 52 111 53 112
rect 51 111 52 112
rect 50 111 51 112
rect 49 111 50 112
rect 48 111 49 112
rect 47 111 48 112
rect 33 111 34 112
rect 32 111 33 112
rect 31 111 32 112
rect 30 111 31 112
rect 29 111 30 112
rect 28 111 29 112
rect 27 111 28 112
rect 26 111 27 112
rect 25 111 26 112
rect 24 111 25 112
rect 23 111 24 112
rect 22 111 23 112
rect 21 111 22 112
rect 20 111 21 112
rect 19 111 20 112
rect 18 111 19 112
rect 146 112 147 113
rect 145 112 146 113
rect 144 112 145 113
rect 143 112 144 113
rect 142 112 143 113
rect 141 112 142 113
rect 140 112 141 113
rect 139 112 140 113
rect 138 112 139 113
rect 137 112 138 113
rect 136 112 137 113
rect 135 112 136 113
rect 134 112 135 113
rect 133 112 134 113
rect 132 112 133 113
rect 131 112 132 113
rect 130 112 131 113
rect 129 112 130 113
rect 128 112 129 113
rect 127 112 128 113
rect 126 112 127 113
rect 125 112 126 113
rect 124 112 125 113
rect 123 112 124 113
rect 122 112 123 113
rect 121 112 122 113
rect 62 112 63 113
rect 61 112 62 113
rect 60 112 61 113
rect 59 112 60 113
rect 58 112 59 113
rect 57 112 58 113
rect 56 112 57 113
rect 55 112 56 113
rect 54 112 55 113
rect 53 112 54 113
rect 52 112 53 113
rect 51 112 52 113
rect 50 112 51 113
rect 49 112 50 113
rect 48 112 49 113
rect 47 112 48 113
rect 46 112 47 113
rect 35 112 36 113
rect 34 112 35 113
rect 33 112 34 113
rect 32 112 33 113
rect 31 112 32 113
rect 30 112 31 113
rect 29 112 30 113
rect 28 112 29 113
rect 27 112 28 113
rect 26 112 27 113
rect 25 112 26 113
rect 24 112 25 113
rect 23 112 24 113
rect 22 112 23 113
rect 21 112 22 113
rect 20 112 21 113
rect 19 112 20 113
rect 18 112 19 113
rect 146 113 147 114
rect 145 113 146 114
rect 144 113 145 114
rect 143 113 144 114
rect 142 113 143 114
rect 141 113 142 114
rect 140 113 141 114
rect 139 113 140 114
rect 138 113 139 114
rect 137 113 138 114
rect 136 113 137 114
rect 135 113 136 114
rect 134 113 135 114
rect 133 113 134 114
rect 132 113 133 114
rect 131 113 132 114
rect 130 113 131 114
rect 129 113 130 114
rect 128 113 129 114
rect 127 113 128 114
rect 126 113 127 114
rect 125 113 126 114
rect 124 113 125 114
rect 123 113 124 114
rect 122 113 123 114
rect 121 113 122 114
rect 61 113 62 114
rect 60 113 61 114
rect 59 113 60 114
rect 58 113 59 114
rect 57 113 58 114
rect 56 113 57 114
rect 55 113 56 114
rect 54 113 55 114
rect 53 113 54 114
rect 52 113 53 114
rect 51 113 52 114
rect 50 113 51 114
rect 49 113 50 114
rect 48 113 49 114
rect 47 113 48 114
rect 46 113 47 114
rect 45 113 46 114
rect 44 113 45 114
rect 43 113 44 114
rect 37 113 38 114
rect 36 113 37 114
rect 35 113 36 114
rect 34 113 35 114
rect 33 113 34 114
rect 32 113 33 114
rect 31 113 32 114
rect 30 113 31 114
rect 29 113 30 114
rect 28 113 29 114
rect 27 113 28 114
rect 26 113 27 114
rect 25 113 26 114
rect 24 113 25 114
rect 23 113 24 114
rect 22 113 23 114
rect 21 113 22 114
rect 20 113 21 114
rect 19 113 20 114
rect 18 113 19 114
rect 146 114 147 115
rect 145 114 146 115
rect 144 114 145 115
rect 143 114 144 115
rect 142 114 143 115
rect 141 114 142 115
rect 140 114 141 115
rect 139 114 140 115
rect 138 114 139 115
rect 137 114 138 115
rect 136 114 137 115
rect 135 114 136 115
rect 134 114 135 115
rect 133 114 134 115
rect 132 114 133 115
rect 131 114 132 115
rect 130 114 131 115
rect 129 114 130 115
rect 128 114 129 115
rect 127 114 128 115
rect 126 114 127 115
rect 125 114 126 115
rect 124 114 125 115
rect 123 114 124 115
rect 122 114 123 115
rect 121 114 122 115
rect 61 114 62 115
rect 60 114 61 115
rect 59 114 60 115
rect 58 114 59 115
rect 57 114 58 115
rect 56 114 57 115
rect 55 114 56 115
rect 54 114 55 115
rect 53 114 54 115
rect 52 114 53 115
rect 51 114 52 115
rect 50 114 51 115
rect 49 114 50 115
rect 48 114 49 115
rect 47 114 48 115
rect 46 114 47 115
rect 45 114 46 115
rect 44 114 45 115
rect 43 114 44 115
rect 42 114 43 115
rect 41 114 42 115
rect 40 114 41 115
rect 39 114 40 115
rect 38 114 39 115
rect 37 114 38 115
rect 36 114 37 115
rect 35 114 36 115
rect 34 114 35 115
rect 33 114 34 115
rect 32 114 33 115
rect 31 114 32 115
rect 30 114 31 115
rect 29 114 30 115
rect 28 114 29 115
rect 27 114 28 115
rect 26 114 27 115
rect 25 114 26 115
rect 24 114 25 115
rect 23 114 24 115
rect 22 114 23 115
rect 21 114 22 115
rect 20 114 21 115
rect 19 114 20 115
rect 18 114 19 115
rect 141 115 142 116
rect 140 115 141 116
rect 139 115 140 116
rect 138 115 139 116
rect 61 115 62 116
rect 60 115 61 116
rect 59 115 60 116
rect 58 115 59 116
rect 57 115 58 116
rect 56 115 57 116
rect 55 115 56 116
rect 54 115 55 116
rect 53 115 54 116
rect 52 115 53 116
rect 51 115 52 116
rect 50 115 51 116
rect 49 115 50 116
rect 48 115 49 116
rect 47 115 48 116
rect 46 115 47 116
rect 45 115 46 116
rect 44 115 45 116
rect 43 115 44 116
rect 42 115 43 116
rect 41 115 42 116
rect 40 115 41 116
rect 39 115 40 116
rect 38 115 39 116
rect 37 115 38 116
rect 36 115 37 116
rect 35 115 36 116
rect 34 115 35 116
rect 33 115 34 116
rect 32 115 33 116
rect 31 115 32 116
rect 30 115 31 116
rect 29 115 30 116
rect 28 115 29 116
rect 27 115 28 116
rect 26 115 27 116
rect 25 115 26 116
rect 24 115 25 116
rect 23 115 24 116
rect 22 115 23 116
rect 21 115 22 116
rect 20 115 21 116
rect 19 115 20 116
rect 141 116 142 117
rect 140 116 141 117
rect 139 116 140 117
rect 138 116 139 117
rect 61 116 62 117
rect 60 116 61 117
rect 59 116 60 117
rect 58 116 59 117
rect 57 116 58 117
rect 56 116 57 117
rect 55 116 56 117
rect 54 116 55 117
rect 53 116 54 117
rect 52 116 53 117
rect 51 116 52 117
rect 50 116 51 117
rect 49 116 50 117
rect 48 116 49 117
rect 47 116 48 117
rect 46 116 47 117
rect 45 116 46 117
rect 44 116 45 117
rect 43 116 44 117
rect 42 116 43 117
rect 41 116 42 117
rect 40 116 41 117
rect 39 116 40 117
rect 38 116 39 117
rect 37 116 38 117
rect 36 116 37 117
rect 35 116 36 117
rect 34 116 35 117
rect 33 116 34 117
rect 32 116 33 117
rect 31 116 32 117
rect 30 116 31 117
rect 29 116 30 117
rect 28 116 29 117
rect 27 116 28 117
rect 26 116 27 117
rect 25 116 26 117
rect 24 116 25 117
rect 23 116 24 117
rect 22 116 23 117
rect 21 116 22 117
rect 20 116 21 117
rect 19 116 20 117
rect 141 117 142 118
rect 140 117 141 118
rect 139 117 140 118
rect 138 117 139 118
rect 61 117 62 118
rect 60 117 61 118
rect 59 117 60 118
rect 58 117 59 118
rect 57 117 58 118
rect 56 117 57 118
rect 55 117 56 118
rect 54 117 55 118
rect 53 117 54 118
rect 52 117 53 118
rect 51 117 52 118
rect 50 117 51 118
rect 49 117 50 118
rect 48 117 49 118
rect 47 117 48 118
rect 46 117 47 118
rect 45 117 46 118
rect 44 117 45 118
rect 43 117 44 118
rect 42 117 43 118
rect 41 117 42 118
rect 40 117 41 118
rect 39 117 40 118
rect 38 117 39 118
rect 37 117 38 118
rect 36 117 37 118
rect 35 117 36 118
rect 34 117 35 118
rect 33 117 34 118
rect 32 117 33 118
rect 31 117 32 118
rect 30 117 31 118
rect 29 117 30 118
rect 28 117 29 118
rect 27 117 28 118
rect 26 117 27 118
rect 25 117 26 118
rect 24 117 25 118
rect 23 117 24 118
rect 22 117 23 118
rect 21 117 22 118
rect 20 117 21 118
rect 19 117 20 118
rect 60 118 61 119
rect 59 118 60 119
rect 58 118 59 119
rect 57 118 58 119
rect 56 118 57 119
rect 55 118 56 119
rect 54 118 55 119
rect 53 118 54 119
rect 52 118 53 119
rect 51 118 52 119
rect 50 118 51 119
rect 49 118 50 119
rect 48 118 49 119
rect 47 118 48 119
rect 46 118 47 119
rect 45 118 46 119
rect 44 118 45 119
rect 43 118 44 119
rect 42 118 43 119
rect 41 118 42 119
rect 40 118 41 119
rect 39 118 40 119
rect 38 118 39 119
rect 37 118 38 119
rect 36 118 37 119
rect 35 118 36 119
rect 34 118 35 119
rect 33 118 34 119
rect 32 118 33 119
rect 31 118 32 119
rect 30 118 31 119
rect 29 118 30 119
rect 28 118 29 119
rect 27 118 28 119
rect 26 118 27 119
rect 25 118 26 119
rect 24 118 25 119
rect 23 118 24 119
rect 22 118 23 119
rect 21 118 22 119
rect 20 118 21 119
rect 19 118 20 119
rect 60 119 61 120
rect 59 119 60 120
rect 58 119 59 120
rect 57 119 58 120
rect 56 119 57 120
rect 55 119 56 120
rect 54 119 55 120
rect 53 119 54 120
rect 52 119 53 120
rect 51 119 52 120
rect 50 119 51 120
rect 49 119 50 120
rect 48 119 49 120
rect 47 119 48 120
rect 46 119 47 120
rect 45 119 46 120
rect 44 119 45 120
rect 43 119 44 120
rect 42 119 43 120
rect 41 119 42 120
rect 40 119 41 120
rect 39 119 40 120
rect 38 119 39 120
rect 37 119 38 120
rect 36 119 37 120
rect 35 119 36 120
rect 34 119 35 120
rect 33 119 34 120
rect 32 119 33 120
rect 31 119 32 120
rect 30 119 31 120
rect 29 119 30 120
rect 28 119 29 120
rect 27 119 28 120
rect 26 119 27 120
rect 25 119 26 120
rect 24 119 25 120
rect 23 119 24 120
rect 22 119 23 120
rect 21 119 22 120
rect 20 119 21 120
rect 19 119 20 120
rect 151 120 152 121
rect 150 120 151 121
rect 149 120 150 121
rect 148 120 149 121
rect 60 120 61 121
rect 59 120 60 121
rect 58 120 59 121
rect 57 120 58 121
rect 56 120 57 121
rect 55 120 56 121
rect 54 120 55 121
rect 53 120 54 121
rect 52 120 53 121
rect 51 120 52 121
rect 50 120 51 121
rect 49 120 50 121
rect 48 120 49 121
rect 47 120 48 121
rect 46 120 47 121
rect 45 120 46 121
rect 44 120 45 121
rect 43 120 44 121
rect 42 120 43 121
rect 41 120 42 121
rect 40 120 41 121
rect 39 120 40 121
rect 38 120 39 121
rect 37 120 38 121
rect 36 120 37 121
rect 35 120 36 121
rect 34 120 35 121
rect 33 120 34 121
rect 32 120 33 121
rect 31 120 32 121
rect 30 120 31 121
rect 29 120 30 121
rect 28 120 29 121
rect 27 120 28 121
rect 26 120 27 121
rect 25 120 26 121
rect 24 120 25 121
rect 23 120 24 121
rect 22 120 23 121
rect 21 120 22 121
rect 20 120 21 121
rect 19 120 20 121
rect 151 121 152 122
rect 150 121 151 122
rect 149 121 150 122
rect 148 121 149 122
rect 147 121 148 122
rect 146 121 147 122
rect 145 121 146 122
rect 144 121 145 122
rect 143 121 144 122
rect 59 121 60 122
rect 58 121 59 122
rect 57 121 58 122
rect 56 121 57 122
rect 55 121 56 122
rect 54 121 55 122
rect 53 121 54 122
rect 52 121 53 122
rect 51 121 52 122
rect 50 121 51 122
rect 49 121 50 122
rect 48 121 49 122
rect 47 121 48 122
rect 46 121 47 122
rect 45 121 46 122
rect 44 121 45 122
rect 43 121 44 122
rect 42 121 43 122
rect 41 121 42 122
rect 40 121 41 122
rect 39 121 40 122
rect 38 121 39 122
rect 37 121 38 122
rect 36 121 37 122
rect 35 121 36 122
rect 34 121 35 122
rect 33 121 34 122
rect 32 121 33 122
rect 31 121 32 122
rect 30 121 31 122
rect 29 121 30 122
rect 28 121 29 122
rect 27 121 28 122
rect 26 121 27 122
rect 25 121 26 122
rect 24 121 25 122
rect 23 121 24 122
rect 22 121 23 122
rect 21 121 22 122
rect 20 121 21 122
rect 151 122 152 123
rect 150 122 151 123
rect 149 122 150 123
rect 148 122 149 123
rect 147 122 148 123
rect 146 122 147 123
rect 145 122 146 123
rect 144 122 145 123
rect 143 122 144 123
rect 59 122 60 123
rect 58 122 59 123
rect 57 122 58 123
rect 56 122 57 123
rect 55 122 56 123
rect 54 122 55 123
rect 53 122 54 123
rect 52 122 53 123
rect 51 122 52 123
rect 50 122 51 123
rect 49 122 50 123
rect 48 122 49 123
rect 47 122 48 123
rect 46 122 47 123
rect 45 122 46 123
rect 44 122 45 123
rect 43 122 44 123
rect 42 122 43 123
rect 41 122 42 123
rect 40 122 41 123
rect 39 122 40 123
rect 38 122 39 123
rect 37 122 38 123
rect 36 122 37 123
rect 35 122 36 123
rect 34 122 35 123
rect 33 122 34 123
rect 32 122 33 123
rect 31 122 32 123
rect 30 122 31 123
rect 29 122 30 123
rect 28 122 29 123
rect 27 122 28 123
rect 26 122 27 123
rect 25 122 26 123
rect 24 122 25 123
rect 23 122 24 123
rect 22 122 23 123
rect 21 122 22 123
rect 20 122 21 123
rect 151 123 152 124
rect 150 123 151 124
rect 149 123 150 124
rect 148 123 149 124
rect 147 123 148 124
rect 146 123 147 124
rect 145 123 146 124
rect 144 123 145 124
rect 143 123 144 124
rect 58 123 59 124
rect 57 123 58 124
rect 56 123 57 124
rect 55 123 56 124
rect 54 123 55 124
rect 53 123 54 124
rect 52 123 53 124
rect 51 123 52 124
rect 50 123 51 124
rect 49 123 50 124
rect 48 123 49 124
rect 47 123 48 124
rect 46 123 47 124
rect 45 123 46 124
rect 44 123 45 124
rect 43 123 44 124
rect 42 123 43 124
rect 41 123 42 124
rect 40 123 41 124
rect 39 123 40 124
rect 38 123 39 124
rect 37 123 38 124
rect 36 123 37 124
rect 35 123 36 124
rect 34 123 35 124
rect 33 123 34 124
rect 32 123 33 124
rect 31 123 32 124
rect 30 123 31 124
rect 29 123 30 124
rect 28 123 29 124
rect 27 123 28 124
rect 26 123 27 124
rect 25 123 26 124
rect 24 123 25 124
rect 23 123 24 124
rect 22 123 23 124
rect 21 123 22 124
rect 20 123 21 124
rect 149 124 150 125
rect 148 124 149 125
rect 147 124 148 125
rect 146 124 147 125
rect 145 124 146 125
rect 144 124 145 125
rect 143 124 144 125
rect 58 124 59 125
rect 57 124 58 125
rect 56 124 57 125
rect 55 124 56 125
rect 54 124 55 125
rect 53 124 54 125
rect 52 124 53 125
rect 51 124 52 125
rect 50 124 51 125
rect 49 124 50 125
rect 48 124 49 125
rect 47 124 48 125
rect 46 124 47 125
rect 45 124 46 125
rect 44 124 45 125
rect 43 124 44 125
rect 42 124 43 125
rect 41 124 42 125
rect 40 124 41 125
rect 39 124 40 125
rect 38 124 39 125
rect 37 124 38 125
rect 36 124 37 125
rect 35 124 36 125
rect 34 124 35 125
rect 33 124 34 125
rect 32 124 33 125
rect 31 124 32 125
rect 30 124 31 125
rect 29 124 30 125
rect 28 124 29 125
rect 27 124 28 125
rect 26 124 27 125
rect 25 124 26 125
rect 24 124 25 125
rect 23 124 24 125
rect 22 124 23 125
rect 21 124 22 125
rect 146 125 147 126
rect 145 125 146 126
rect 144 125 145 126
rect 143 125 144 126
rect 57 125 58 126
rect 56 125 57 126
rect 55 125 56 126
rect 54 125 55 126
rect 53 125 54 126
rect 52 125 53 126
rect 51 125 52 126
rect 50 125 51 126
rect 49 125 50 126
rect 48 125 49 126
rect 47 125 48 126
rect 46 125 47 126
rect 45 125 46 126
rect 44 125 45 126
rect 43 125 44 126
rect 42 125 43 126
rect 41 125 42 126
rect 40 125 41 126
rect 39 125 40 126
rect 38 125 39 126
rect 37 125 38 126
rect 36 125 37 126
rect 35 125 36 126
rect 34 125 35 126
rect 33 125 34 126
rect 32 125 33 126
rect 31 125 32 126
rect 30 125 31 126
rect 29 125 30 126
rect 28 125 29 126
rect 27 125 28 126
rect 26 125 27 126
rect 25 125 26 126
rect 24 125 25 126
rect 23 125 24 126
rect 22 125 23 126
rect 21 125 22 126
rect 143 126 144 127
rect 56 126 57 127
rect 55 126 56 127
rect 54 126 55 127
rect 53 126 54 127
rect 52 126 53 127
rect 51 126 52 127
rect 50 126 51 127
rect 49 126 50 127
rect 48 126 49 127
rect 47 126 48 127
rect 46 126 47 127
rect 45 126 46 127
rect 44 126 45 127
rect 43 126 44 127
rect 42 126 43 127
rect 41 126 42 127
rect 40 126 41 127
rect 39 126 40 127
rect 38 126 39 127
rect 37 126 38 127
rect 36 126 37 127
rect 35 126 36 127
rect 34 126 35 127
rect 33 126 34 127
rect 32 126 33 127
rect 31 126 32 127
rect 30 126 31 127
rect 29 126 30 127
rect 28 126 29 127
rect 27 126 28 127
rect 26 126 27 127
rect 25 126 26 127
rect 24 126 25 127
rect 23 126 24 127
rect 22 126 23 127
rect 55 127 56 128
rect 54 127 55 128
rect 53 127 54 128
rect 52 127 53 128
rect 51 127 52 128
rect 50 127 51 128
rect 49 127 50 128
rect 48 127 49 128
rect 47 127 48 128
rect 46 127 47 128
rect 45 127 46 128
rect 44 127 45 128
rect 43 127 44 128
rect 42 127 43 128
rect 41 127 42 128
rect 40 127 41 128
rect 39 127 40 128
rect 38 127 39 128
rect 37 127 38 128
rect 36 127 37 128
rect 35 127 36 128
rect 34 127 35 128
rect 33 127 34 128
rect 32 127 33 128
rect 31 127 32 128
rect 30 127 31 128
rect 29 127 30 128
rect 28 127 29 128
rect 27 127 28 128
rect 26 127 27 128
rect 25 127 26 128
rect 24 127 25 128
rect 23 127 24 128
rect 55 128 56 129
rect 54 128 55 129
rect 53 128 54 129
rect 52 128 53 129
rect 51 128 52 129
rect 50 128 51 129
rect 49 128 50 129
rect 48 128 49 129
rect 47 128 48 129
rect 46 128 47 129
rect 45 128 46 129
rect 44 128 45 129
rect 43 128 44 129
rect 42 128 43 129
rect 41 128 42 129
rect 40 128 41 129
rect 39 128 40 129
rect 38 128 39 129
rect 37 128 38 129
rect 36 128 37 129
rect 35 128 36 129
rect 34 128 35 129
rect 33 128 34 129
rect 32 128 33 129
rect 31 128 32 129
rect 30 128 31 129
rect 29 128 30 129
rect 28 128 29 129
rect 27 128 28 129
rect 26 128 27 129
rect 25 128 26 129
rect 24 128 25 129
rect 23 128 24 129
rect 54 129 55 130
rect 53 129 54 130
rect 52 129 53 130
rect 51 129 52 130
rect 50 129 51 130
rect 49 129 50 130
rect 48 129 49 130
rect 47 129 48 130
rect 46 129 47 130
rect 45 129 46 130
rect 44 129 45 130
rect 43 129 44 130
rect 42 129 43 130
rect 41 129 42 130
rect 40 129 41 130
rect 39 129 40 130
rect 38 129 39 130
rect 37 129 38 130
rect 36 129 37 130
rect 35 129 36 130
rect 34 129 35 130
rect 33 129 34 130
rect 32 129 33 130
rect 31 129 32 130
rect 30 129 31 130
rect 29 129 30 130
rect 28 129 29 130
rect 27 129 28 130
rect 26 129 27 130
rect 25 129 26 130
rect 24 129 25 130
rect 52 130 53 131
rect 51 130 52 131
rect 50 130 51 131
rect 49 130 50 131
rect 48 130 49 131
rect 47 130 48 131
rect 46 130 47 131
rect 45 130 46 131
rect 44 130 45 131
rect 43 130 44 131
rect 42 130 43 131
rect 41 130 42 131
rect 40 130 41 131
rect 39 130 40 131
rect 38 130 39 131
rect 37 130 38 131
rect 36 130 37 131
rect 35 130 36 131
rect 34 130 35 131
rect 33 130 34 131
rect 32 130 33 131
rect 31 130 32 131
rect 30 130 31 131
rect 29 130 30 131
rect 28 130 29 131
rect 27 130 28 131
rect 26 130 27 131
rect 25 130 26 131
rect 51 131 52 132
rect 50 131 51 132
rect 49 131 50 132
rect 48 131 49 132
rect 47 131 48 132
rect 46 131 47 132
rect 45 131 46 132
rect 44 131 45 132
rect 43 131 44 132
rect 42 131 43 132
rect 41 131 42 132
rect 40 131 41 132
rect 39 131 40 132
rect 38 131 39 132
rect 37 131 38 132
rect 36 131 37 132
rect 35 131 36 132
rect 34 131 35 132
rect 33 131 34 132
rect 32 131 33 132
rect 31 131 32 132
rect 30 131 31 132
rect 29 131 30 132
rect 28 131 29 132
rect 27 131 28 132
rect 49 132 50 133
rect 48 132 49 133
rect 47 132 48 133
rect 46 132 47 133
rect 45 132 46 133
rect 44 132 45 133
rect 43 132 44 133
rect 42 132 43 133
rect 41 132 42 133
rect 40 132 41 133
rect 39 132 40 133
rect 38 132 39 133
rect 37 132 38 133
rect 36 132 37 133
rect 35 132 36 133
rect 34 132 35 133
rect 33 132 34 133
rect 32 132 33 133
rect 31 132 32 133
rect 30 132 31 133
rect 29 132 30 133
rect 28 132 29 133
rect 47 133 48 134
rect 46 133 47 134
rect 45 133 46 134
rect 44 133 45 134
rect 43 133 44 134
rect 42 133 43 134
rect 41 133 42 134
rect 40 133 41 134
rect 39 133 40 134
rect 38 133 39 134
rect 37 133 38 134
rect 36 133 37 134
rect 35 133 36 134
rect 34 133 35 134
rect 33 133 34 134
rect 32 133 33 134
rect 31 133 32 134
rect 30 133 31 134
rect 44 134 45 135
rect 43 134 44 135
rect 42 134 43 135
rect 41 134 42 135
rect 40 134 41 135
rect 39 134 40 135
rect 38 134 39 135
rect 37 134 38 135
rect 36 134 37 135
rect 35 134 36 135
rect 34 134 35 135
rect 146 140 147 141
rect 145 140 146 141
rect 144 140 145 141
rect 143 140 144 141
rect 142 140 143 141
rect 141 140 142 141
rect 146 141 147 142
rect 145 141 146 142
rect 144 141 145 142
rect 143 141 144 142
rect 142 141 143 142
rect 146 142 147 143
rect 145 142 146 143
rect 144 142 145 143
rect 143 142 144 143
rect 142 142 143 143
rect 54 142 55 143
rect 53 142 54 143
rect 52 142 53 143
rect 51 142 52 143
rect 50 142 51 143
rect 49 142 50 143
rect 48 142 49 143
rect 47 142 48 143
rect 46 142 47 143
rect 45 142 46 143
rect 44 142 45 143
rect 43 142 44 143
rect 42 142 43 143
rect 41 142 42 143
rect 40 142 41 143
rect 39 142 40 143
rect 38 142 39 143
rect 37 142 38 143
rect 36 142 37 143
rect 35 142 36 143
rect 34 142 35 143
rect 33 142 34 143
rect 32 142 33 143
rect 31 142 32 143
rect 30 142 31 143
rect 29 142 30 143
rect 28 142 29 143
rect 27 142 28 143
rect 26 142 27 143
rect 25 142 26 143
rect 24 142 25 143
rect 23 142 24 143
rect 22 142 23 143
rect 21 142 22 143
rect 20 142 21 143
rect 19 142 20 143
rect 18 142 19 143
rect 146 143 147 144
rect 145 143 146 144
rect 144 143 145 144
rect 143 143 144 144
rect 142 143 143 144
rect 65 143 66 144
rect 64 143 65 144
rect 63 143 64 144
rect 62 143 63 144
rect 61 143 62 144
rect 60 143 61 144
rect 59 143 60 144
rect 58 143 59 144
rect 57 143 58 144
rect 56 143 57 144
rect 55 143 56 144
rect 54 143 55 144
rect 53 143 54 144
rect 52 143 53 144
rect 51 143 52 144
rect 50 143 51 144
rect 49 143 50 144
rect 48 143 49 144
rect 47 143 48 144
rect 46 143 47 144
rect 45 143 46 144
rect 44 143 45 144
rect 43 143 44 144
rect 42 143 43 144
rect 41 143 42 144
rect 40 143 41 144
rect 39 143 40 144
rect 38 143 39 144
rect 37 143 38 144
rect 36 143 37 144
rect 35 143 36 144
rect 34 143 35 144
rect 33 143 34 144
rect 32 143 33 144
rect 31 143 32 144
rect 30 143 31 144
rect 29 143 30 144
rect 28 143 29 144
rect 27 143 28 144
rect 26 143 27 144
rect 25 143 26 144
rect 24 143 25 144
rect 23 143 24 144
rect 22 143 23 144
rect 21 143 22 144
rect 20 143 21 144
rect 19 143 20 144
rect 18 143 19 144
rect 146 144 147 145
rect 145 144 146 145
rect 144 144 145 145
rect 143 144 144 145
rect 142 144 143 145
rect 68 144 69 145
rect 67 144 68 145
rect 66 144 67 145
rect 65 144 66 145
rect 64 144 65 145
rect 63 144 64 145
rect 62 144 63 145
rect 61 144 62 145
rect 60 144 61 145
rect 59 144 60 145
rect 58 144 59 145
rect 57 144 58 145
rect 56 144 57 145
rect 55 144 56 145
rect 54 144 55 145
rect 53 144 54 145
rect 52 144 53 145
rect 51 144 52 145
rect 50 144 51 145
rect 49 144 50 145
rect 48 144 49 145
rect 47 144 48 145
rect 46 144 47 145
rect 45 144 46 145
rect 44 144 45 145
rect 43 144 44 145
rect 42 144 43 145
rect 41 144 42 145
rect 40 144 41 145
rect 39 144 40 145
rect 38 144 39 145
rect 37 144 38 145
rect 36 144 37 145
rect 35 144 36 145
rect 34 144 35 145
rect 33 144 34 145
rect 32 144 33 145
rect 31 144 32 145
rect 30 144 31 145
rect 29 144 30 145
rect 28 144 29 145
rect 27 144 28 145
rect 26 144 27 145
rect 25 144 26 145
rect 24 144 25 145
rect 23 144 24 145
rect 22 144 23 145
rect 21 144 22 145
rect 20 144 21 145
rect 19 144 20 145
rect 18 144 19 145
rect 146 145 147 146
rect 145 145 146 146
rect 144 145 145 146
rect 143 145 144 146
rect 142 145 143 146
rect 141 145 142 146
rect 71 145 72 146
rect 70 145 71 146
rect 69 145 70 146
rect 68 145 69 146
rect 67 145 68 146
rect 66 145 67 146
rect 65 145 66 146
rect 64 145 65 146
rect 63 145 64 146
rect 62 145 63 146
rect 61 145 62 146
rect 60 145 61 146
rect 59 145 60 146
rect 58 145 59 146
rect 57 145 58 146
rect 56 145 57 146
rect 55 145 56 146
rect 54 145 55 146
rect 53 145 54 146
rect 52 145 53 146
rect 51 145 52 146
rect 50 145 51 146
rect 49 145 50 146
rect 48 145 49 146
rect 47 145 48 146
rect 46 145 47 146
rect 45 145 46 146
rect 44 145 45 146
rect 43 145 44 146
rect 42 145 43 146
rect 41 145 42 146
rect 40 145 41 146
rect 39 145 40 146
rect 38 145 39 146
rect 37 145 38 146
rect 36 145 37 146
rect 35 145 36 146
rect 34 145 35 146
rect 33 145 34 146
rect 32 145 33 146
rect 31 145 32 146
rect 30 145 31 146
rect 29 145 30 146
rect 28 145 29 146
rect 27 145 28 146
rect 26 145 27 146
rect 25 145 26 146
rect 24 145 25 146
rect 23 145 24 146
rect 22 145 23 146
rect 21 145 22 146
rect 20 145 21 146
rect 19 145 20 146
rect 18 145 19 146
rect 146 146 147 147
rect 145 146 146 147
rect 144 146 145 147
rect 143 146 144 147
rect 142 146 143 147
rect 141 146 142 147
rect 140 146 141 147
rect 73 146 74 147
rect 72 146 73 147
rect 71 146 72 147
rect 70 146 71 147
rect 69 146 70 147
rect 68 146 69 147
rect 67 146 68 147
rect 66 146 67 147
rect 65 146 66 147
rect 64 146 65 147
rect 63 146 64 147
rect 62 146 63 147
rect 61 146 62 147
rect 60 146 61 147
rect 59 146 60 147
rect 58 146 59 147
rect 57 146 58 147
rect 56 146 57 147
rect 55 146 56 147
rect 54 146 55 147
rect 53 146 54 147
rect 52 146 53 147
rect 51 146 52 147
rect 50 146 51 147
rect 49 146 50 147
rect 48 146 49 147
rect 47 146 48 147
rect 46 146 47 147
rect 45 146 46 147
rect 44 146 45 147
rect 43 146 44 147
rect 42 146 43 147
rect 41 146 42 147
rect 40 146 41 147
rect 39 146 40 147
rect 38 146 39 147
rect 37 146 38 147
rect 36 146 37 147
rect 35 146 36 147
rect 34 146 35 147
rect 33 146 34 147
rect 32 146 33 147
rect 31 146 32 147
rect 30 146 31 147
rect 29 146 30 147
rect 28 146 29 147
rect 27 146 28 147
rect 26 146 27 147
rect 25 146 26 147
rect 24 146 25 147
rect 23 146 24 147
rect 22 146 23 147
rect 21 146 22 147
rect 20 146 21 147
rect 19 146 20 147
rect 18 146 19 147
rect 145 147 146 148
rect 144 147 145 148
rect 143 147 144 148
rect 142 147 143 148
rect 141 147 142 148
rect 140 147 141 148
rect 139 147 140 148
rect 138 147 139 148
rect 137 147 138 148
rect 136 147 137 148
rect 135 147 136 148
rect 134 147 135 148
rect 133 147 134 148
rect 132 147 133 148
rect 131 147 132 148
rect 130 147 131 148
rect 129 147 130 148
rect 128 147 129 148
rect 127 147 128 148
rect 126 147 127 148
rect 125 147 126 148
rect 124 147 125 148
rect 123 147 124 148
rect 122 147 123 148
rect 121 147 122 148
rect 74 147 75 148
rect 73 147 74 148
rect 72 147 73 148
rect 71 147 72 148
rect 70 147 71 148
rect 69 147 70 148
rect 68 147 69 148
rect 67 147 68 148
rect 66 147 67 148
rect 65 147 66 148
rect 64 147 65 148
rect 63 147 64 148
rect 62 147 63 148
rect 61 147 62 148
rect 60 147 61 148
rect 59 147 60 148
rect 58 147 59 148
rect 57 147 58 148
rect 56 147 57 148
rect 55 147 56 148
rect 54 147 55 148
rect 53 147 54 148
rect 52 147 53 148
rect 51 147 52 148
rect 50 147 51 148
rect 49 147 50 148
rect 48 147 49 148
rect 47 147 48 148
rect 46 147 47 148
rect 45 147 46 148
rect 44 147 45 148
rect 43 147 44 148
rect 42 147 43 148
rect 41 147 42 148
rect 40 147 41 148
rect 39 147 40 148
rect 38 147 39 148
rect 37 147 38 148
rect 36 147 37 148
rect 35 147 36 148
rect 34 147 35 148
rect 33 147 34 148
rect 32 147 33 148
rect 31 147 32 148
rect 30 147 31 148
rect 29 147 30 148
rect 28 147 29 148
rect 27 147 28 148
rect 26 147 27 148
rect 25 147 26 148
rect 24 147 25 148
rect 23 147 24 148
rect 22 147 23 148
rect 21 147 22 148
rect 20 147 21 148
rect 19 147 20 148
rect 18 147 19 148
rect 145 148 146 149
rect 144 148 145 149
rect 143 148 144 149
rect 142 148 143 149
rect 141 148 142 149
rect 140 148 141 149
rect 139 148 140 149
rect 138 148 139 149
rect 137 148 138 149
rect 136 148 137 149
rect 135 148 136 149
rect 134 148 135 149
rect 133 148 134 149
rect 132 148 133 149
rect 131 148 132 149
rect 130 148 131 149
rect 129 148 130 149
rect 128 148 129 149
rect 127 148 128 149
rect 126 148 127 149
rect 125 148 126 149
rect 124 148 125 149
rect 123 148 124 149
rect 122 148 123 149
rect 121 148 122 149
rect 76 148 77 149
rect 75 148 76 149
rect 74 148 75 149
rect 73 148 74 149
rect 72 148 73 149
rect 71 148 72 149
rect 70 148 71 149
rect 69 148 70 149
rect 68 148 69 149
rect 67 148 68 149
rect 66 148 67 149
rect 65 148 66 149
rect 64 148 65 149
rect 63 148 64 149
rect 62 148 63 149
rect 61 148 62 149
rect 60 148 61 149
rect 59 148 60 149
rect 58 148 59 149
rect 57 148 58 149
rect 56 148 57 149
rect 55 148 56 149
rect 54 148 55 149
rect 53 148 54 149
rect 52 148 53 149
rect 51 148 52 149
rect 50 148 51 149
rect 49 148 50 149
rect 48 148 49 149
rect 47 148 48 149
rect 46 148 47 149
rect 45 148 46 149
rect 44 148 45 149
rect 43 148 44 149
rect 42 148 43 149
rect 41 148 42 149
rect 40 148 41 149
rect 39 148 40 149
rect 38 148 39 149
rect 37 148 38 149
rect 36 148 37 149
rect 35 148 36 149
rect 34 148 35 149
rect 33 148 34 149
rect 32 148 33 149
rect 31 148 32 149
rect 30 148 31 149
rect 29 148 30 149
rect 28 148 29 149
rect 27 148 28 149
rect 26 148 27 149
rect 25 148 26 149
rect 24 148 25 149
rect 23 148 24 149
rect 22 148 23 149
rect 21 148 22 149
rect 20 148 21 149
rect 19 148 20 149
rect 18 148 19 149
rect 144 149 145 150
rect 143 149 144 150
rect 142 149 143 150
rect 141 149 142 150
rect 140 149 141 150
rect 139 149 140 150
rect 138 149 139 150
rect 137 149 138 150
rect 136 149 137 150
rect 135 149 136 150
rect 134 149 135 150
rect 133 149 134 150
rect 132 149 133 150
rect 131 149 132 150
rect 130 149 131 150
rect 129 149 130 150
rect 128 149 129 150
rect 127 149 128 150
rect 126 149 127 150
rect 125 149 126 150
rect 124 149 125 150
rect 123 149 124 150
rect 122 149 123 150
rect 121 149 122 150
rect 77 149 78 150
rect 76 149 77 150
rect 75 149 76 150
rect 74 149 75 150
rect 73 149 74 150
rect 72 149 73 150
rect 71 149 72 150
rect 70 149 71 150
rect 69 149 70 150
rect 68 149 69 150
rect 67 149 68 150
rect 66 149 67 150
rect 65 149 66 150
rect 64 149 65 150
rect 63 149 64 150
rect 62 149 63 150
rect 61 149 62 150
rect 60 149 61 150
rect 59 149 60 150
rect 58 149 59 150
rect 57 149 58 150
rect 56 149 57 150
rect 55 149 56 150
rect 54 149 55 150
rect 53 149 54 150
rect 52 149 53 150
rect 51 149 52 150
rect 50 149 51 150
rect 49 149 50 150
rect 48 149 49 150
rect 47 149 48 150
rect 46 149 47 150
rect 45 149 46 150
rect 44 149 45 150
rect 43 149 44 150
rect 42 149 43 150
rect 41 149 42 150
rect 40 149 41 150
rect 39 149 40 150
rect 38 149 39 150
rect 37 149 38 150
rect 36 149 37 150
rect 35 149 36 150
rect 34 149 35 150
rect 33 149 34 150
rect 32 149 33 150
rect 31 149 32 150
rect 30 149 31 150
rect 29 149 30 150
rect 28 149 29 150
rect 27 149 28 150
rect 26 149 27 150
rect 25 149 26 150
rect 24 149 25 150
rect 23 149 24 150
rect 22 149 23 150
rect 21 149 22 150
rect 20 149 21 150
rect 19 149 20 150
rect 18 149 19 150
rect 143 150 144 151
rect 142 150 143 151
rect 141 150 142 151
rect 140 150 141 151
rect 139 150 140 151
rect 138 150 139 151
rect 137 150 138 151
rect 136 150 137 151
rect 135 150 136 151
rect 134 150 135 151
rect 133 150 134 151
rect 132 150 133 151
rect 131 150 132 151
rect 130 150 131 151
rect 129 150 130 151
rect 128 150 129 151
rect 127 150 128 151
rect 126 150 127 151
rect 125 150 126 151
rect 124 150 125 151
rect 123 150 124 151
rect 122 150 123 151
rect 121 150 122 151
rect 78 150 79 151
rect 77 150 78 151
rect 76 150 77 151
rect 75 150 76 151
rect 74 150 75 151
rect 73 150 74 151
rect 72 150 73 151
rect 71 150 72 151
rect 70 150 71 151
rect 69 150 70 151
rect 68 150 69 151
rect 67 150 68 151
rect 66 150 67 151
rect 65 150 66 151
rect 64 150 65 151
rect 63 150 64 151
rect 62 150 63 151
rect 61 150 62 151
rect 60 150 61 151
rect 59 150 60 151
rect 58 150 59 151
rect 57 150 58 151
rect 56 150 57 151
rect 55 150 56 151
rect 54 150 55 151
rect 53 150 54 151
rect 52 150 53 151
rect 51 150 52 151
rect 50 150 51 151
rect 49 150 50 151
rect 48 150 49 151
rect 47 150 48 151
rect 46 150 47 151
rect 45 150 46 151
rect 44 150 45 151
rect 43 150 44 151
rect 42 150 43 151
rect 41 150 42 151
rect 40 150 41 151
rect 39 150 40 151
rect 38 150 39 151
rect 37 150 38 151
rect 36 150 37 151
rect 35 150 36 151
rect 34 150 35 151
rect 33 150 34 151
rect 32 150 33 151
rect 31 150 32 151
rect 30 150 31 151
rect 29 150 30 151
rect 28 150 29 151
rect 27 150 28 151
rect 26 150 27 151
rect 25 150 26 151
rect 24 150 25 151
rect 23 150 24 151
rect 22 150 23 151
rect 21 150 22 151
rect 20 150 21 151
rect 19 150 20 151
rect 18 150 19 151
rect 142 151 143 152
rect 141 151 142 152
rect 140 151 141 152
rect 139 151 140 152
rect 138 151 139 152
rect 137 151 138 152
rect 136 151 137 152
rect 135 151 136 152
rect 134 151 135 152
rect 133 151 134 152
rect 132 151 133 152
rect 131 151 132 152
rect 130 151 131 152
rect 129 151 130 152
rect 128 151 129 152
rect 127 151 128 152
rect 126 151 127 152
rect 125 151 126 152
rect 124 151 125 152
rect 123 151 124 152
rect 122 151 123 152
rect 121 151 122 152
rect 79 151 80 152
rect 78 151 79 152
rect 77 151 78 152
rect 76 151 77 152
rect 75 151 76 152
rect 74 151 75 152
rect 73 151 74 152
rect 72 151 73 152
rect 71 151 72 152
rect 70 151 71 152
rect 69 151 70 152
rect 68 151 69 152
rect 67 151 68 152
rect 66 151 67 152
rect 65 151 66 152
rect 64 151 65 152
rect 63 151 64 152
rect 62 151 63 152
rect 61 151 62 152
rect 60 151 61 152
rect 59 151 60 152
rect 58 151 59 152
rect 57 151 58 152
rect 56 151 57 152
rect 55 151 56 152
rect 54 151 55 152
rect 53 151 54 152
rect 52 151 53 152
rect 51 151 52 152
rect 50 151 51 152
rect 49 151 50 152
rect 48 151 49 152
rect 47 151 48 152
rect 46 151 47 152
rect 45 151 46 152
rect 44 151 45 152
rect 43 151 44 152
rect 42 151 43 152
rect 41 151 42 152
rect 40 151 41 152
rect 39 151 40 152
rect 38 151 39 152
rect 37 151 38 152
rect 36 151 37 152
rect 35 151 36 152
rect 34 151 35 152
rect 33 151 34 152
rect 32 151 33 152
rect 31 151 32 152
rect 30 151 31 152
rect 29 151 30 152
rect 28 151 29 152
rect 27 151 28 152
rect 26 151 27 152
rect 25 151 26 152
rect 24 151 25 152
rect 23 151 24 152
rect 22 151 23 152
rect 21 151 22 152
rect 20 151 21 152
rect 19 151 20 152
rect 18 151 19 152
rect 139 152 140 153
rect 138 152 139 153
rect 137 152 138 153
rect 136 152 137 153
rect 135 152 136 153
rect 134 152 135 153
rect 133 152 134 153
rect 132 152 133 153
rect 131 152 132 153
rect 130 152 131 153
rect 129 152 130 153
rect 128 152 129 153
rect 127 152 128 153
rect 126 152 127 153
rect 125 152 126 153
rect 124 152 125 153
rect 123 152 124 153
rect 122 152 123 153
rect 121 152 122 153
rect 80 152 81 153
rect 79 152 80 153
rect 78 152 79 153
rect 77 152 78 153
rect 76 152 77 153
rect 75 152 76 153
rect 74 152 75 153
rect 73 152 74 153
rect 72 152 73 153
rect 71 152 72 153
rect 70 152 71 153
rect 69 152 70 153
rect 68 152 69 153
rect 67 152 68 153
rect 66 152 67 153
rect 65 152 66 153
rect 64 152 65 153
rect 63 152 64 153
rect 62 152 63 153
rect 61 152 62 153
rect 60 152 61 153
rect 59 152 60 153
rect 58 152 59 153
rect 57 152 58 153
rect 56 152 57 153
rect 55 152 56 153
rect 54 152 55 153
rect 53 152 54 153
rect 52 152 53 153
rect 51 152 52 153
rect 50 152 51 153
rect 49 152 50 153
rect 48 152 49 153
rect 47 152 48 153
rect 46 152 47 153
rect 45 152 46 153
rect 44 152 45 153
rect 43 152 44 153
rect 42 152 43 153
rect 41 152 42 153
rect 40 152 41 153
rect 39 152 40 153
rect 38 152 39 153
rect 37 152 38 153
rect 36 152 37 153
rect 35 152 36 153
rect 34 152 35 153
rect 33 152 34 153
rect 32 152 33 153
rect 31 152 32 153
rect 30 152 31 153
rect 29 152 30 153
rect 28 152 29 153
rect 27 152 28 153
rect 26 152 27 153
rect 25 152 26 153
rect 24 152 25 153
rect 23 152 24 153
rect 22 152 23 153
rect 21 152 22 153
rect 20 152 21 153
rect 19 152 20 153
rect 18 152 19 153
rect 80 153 81 154
rect 79 153 80 154
rect 78 153 79 154
rect 77 153 78 154
rect 76 153 77 154
rect 75 153 76 154
rect 74 153 75 154
rect 73 153 74 154
rect 72 153 73 154
rect 71 153 72 154
rect 70 153 71 154
rect 69 153 70 154
rect 68 153 69 154
rect 67 153 68 154
rect 66 153 67 154
rect 65 153 66 154
rect 64 153 65 154
rect 63 153 64 154
rect 62 153 63 154
rect 61 153 62 154
rect 60 153 61 154
rect 59 153 60 154
rect 58 153 59 154
rect 57 153 58 154
rect 56 153 57 154
rect 55 153 56 154
rect 54 153 55 154
rect 53 153 54 154
rect 52 153 53 154
rect 51 153 52 154
rect 50 153 51 154
rect 49 153 50 154
rect 48 153 49 154
rect 47 153 48 154
rect 46 153 47 154
rect 45 153 46 154
rect 44 153 45 154
rect 43 153 44 154
rect 42 153 43 154
rect 41 153 42 154
rect 40 153 41 154
rect 39 153 40 154
rect 38 153 39 154
rect 37 153 38 154
rect 36 153 37 154
rect 35 153 36 154
rect 34 153 35 154
rect 33 153 34 154
rect 32 153 33 154
rect 31 153 32 154
rect 30 153 31 154
rect 29 153 30 154
rect 28 153 29 154
rect 27 153 28 154
rect 26 153 27 154
rect 25 153 26 154
rect 24 153 25 154
rect 23 153 24 154
rect 22 153 23 154
rect 21 153 22 154
rect 20 153 21 154
rect 19 153 20 154
rect 18 153 19 154
rect 81 154 82 155
rect 80 154 81 155
rect 79 154 80 155
rect 78 154 79 155
rect 77 154 78 155
rect 76 154 77 155
rect 75 154 76 155
rect 74 154 75 155
rect 73 154 74 155
rect 72 154 73 155
rect 71 154 72 155
rect 70 154 71 155
rect 69 154 70 155
rect 68 154 69 155
rect 67 154 68 155
rect 66 154 67 155
rect 65 154 66 155
rect 64 154 65 155
rect 63 154 64 155
rect 62 154 63 155
rect 61 154 62 155
rect 60 154 61 155
rect 59 154 60 155
rect 58 154 59 155
rect 57 154 58 155
rect 56 154 57 155
rect 55 154 56 155
rect 54 154 55 155
rect 53 154 54 155
rect 52 154 53 155
rect 51 154 52 155
rect 50 154 51 155
rect 49 154 50 155
rect 48 154 49 155
rect 47 154 48 155
rect 46 154 47 155
rect 45 154 46 155
rect 44 154 45 155
rect 43 154 44 155
rect 42 154 43 155
rect 41 154 42 155
rect 40 154 41 155
rect 39 154 40 155
rect 38 154 39 155
rect 37 154 38 155
rect 36 154 37 155
rect 35 154 36 155
rect 34 154 35 155
rect 33 154 34 155
rect 32 154 33 155
rect 31 154 32 155
rect 30 154 31 155
rect 29 154 30 155
rect 28 154 29 155
rect 27 154 28 155
rect 26 154 27 155
rect 25 154 26 155
rect 24 154 25 155
rect 23 154 24 155
rect 22 154 23 155
rect 21 154 22 155
rect 20 154 21 155
rect 19 154 20 155
rect 18 154 19 155
rect 81 155 82 156
rect 80 155 81 156
rect 79 155 80 156
rect 78 155 79 156
rect 77 155 78 156
rect 76 155 77 156
rect 75 155 76 156
rect 74 155 75 156
rect 73 155 74 156
rect 72 155 73 156
rect 71 155 72 156
rect 70 155 71 156
rect 69 155 70 156
rect 68 155 69 156
rect 67 155 68 156
rect 66 155 67 156
rect 65 155 66 156
rect 64 155 65 156
rect 63 155 64 156
rect 62 155 63 156
rect 61 155 62 156
rect 60 155 61 156
rect 59 155 60 156
rect 58 155 59 156
rect 57 155 58 156
rect 56 155 57 156
rect 55 155 56 156
rect 54 155 55 156
rect 53 155 54 156
rect 52 155 53 156
rect 51 155 52 156
rect 50 155 51 156
rect 49 155 50 156
rect 48 155 49 156
rect 47 155 48 156
rect 46 155 47 156
rect 45 155 46 156
rect 44 155 45 156
rect 43 155 44 156
rect 42 155 43 156
rect 41 155 42 156
rect 40 155 41 156
rect 39 155 40 156
rect 38 155 39 156
rect 37 155 38 156
rect 36 155 37 156
rect 35 155 36 156
rect 34 155 35 156
rect 33 155 34 156
rect 32 155 33 156
rect 31 155 32 156
rect 30 155 31 156
rect 29 155 30 156
rect 28 155 29 156
rect 27 155 28 156
rect 26 155 27 156
rect 25 155 26 156
rect 24 155 25 156
rect 23 155 24 156
rect 22 155 23 156
rect 21 155 22 156
rect 20 155 21 156
rect 19 155 20 156
rect 18 155 19 156
rect 82 156 83 157
rect 81 156 82 157
rect 80 156 81 157
rect 79 156 80 157
rect 78 156 79 157
rect 77 156 78 157
rect 76 156 77 157
rect 75 156 76 157
rect 74 156 75 157
rect 73 156 74 157
rect 72 156 73 157
rect 71 156 72 157
rect 70 156 71 157
rect 69 156 70 157
rect 68 156 69 157
rect 67 156 68 157
rect 66 156 67 157
rect 65 156 66 157
rect 64 156 65 157
rect 63 156 64 157
rect 62 156 63 157
rect 61 156 62 157
rect 60 156 61 157
rect 59 156 60 157
rect 58 156 59 157
rect 57 156 58 157
rect 56 156 57 157
rect 55 156 56 157
rect 54 156 55 157
rect 53 156 54 157
rect 52 156 53 157
rect 51 156 52 157
rect 50 156 51 157
rect 49 156 50 157
rect 48 156 49 157
rect 47 156 48 157
rect 46 156 47 157
rect 45 156 46 157
rect 44 156 45 157
rect 43 156 44 157
rect 42 156 43 157
rect 41 156 42 157
rect 40 156 41 157
rect 39 156 40 157
rect 38 156 39 157
rect 37 156 38 157
rect 36 156 37 157
rect 35 156 36 157
rect 34 156 35 157
rect 33 156 34 157
rect 32 156 33 157
rect 31 156 32 157
rect 30 156 31 157
rect 29 156 30 157
rect 28 156 29 157
rect 27 156 28 157
rect 26 156 27 157
rect 25 156 26 157
rect 24 156 25 157
rect 23 156 24 157
rect 22 156 23 157
rect 21 156 22 157
rect 20 156 21 157
rect 19 156 20 157
rect 18 156 19 157
rect 143 157 144 158
rect 142 157 143 158
rect 141 157 142 158
rect 140 157 141 158
rect 139 157 140 158
rect 82 157 83 158
rect 81 157 82 158
rect 80 157 81 158
rect 79 157 80 158
rect 78 157 79 158
rect 77 157 78 158
rect 76 157 77 158
rect 75 157 76 158
rect 74 157 75 158
rect 73 157 74 158
rect 72 157 73 158
rect 71 157 72 158
rect 70 157 71 158
rect 69 157 70 158
rect 68 157 69 158
rect 67 157 68 158
rect 66 157 67 158
rect 65 157 66 158
rect 64 157 65 158
rect 63 157 64 158
rect 62 157 63 158
rect 61 157 62 158
rect 60 157 61 158
rect 59 157 60 158
rect 58 157 59 158
rect 57 157 58 158
rect 56 157 57 158
rect 55 157 56 158
rect 54 157 55 158
rect 53 157 54 158
rect 52 157 53 158
rect 51 157 52 158
rect 50 157 51 158
rect 49 157 50 158
rect 48 157 49 158
rect 47 157 48 158
rect 46 157 47 158
rect 45 157 46 158
rect 44 157 45 158
rect 43 157 44 158
rect 42 157 43 158
rect 41 157 42 158
rect 40 157 41 158
rect 39 157 40 158
rect 38 157 39 158
rect 37 157 38 158
rect 36 157 37 158
rect 35 157 36 158
rect 34 157 35 158
rect 33 157 34 158
rect 32 157 33 158
rect 31 157 32 158
rect 30 157 31 158
rect 29 157 30 158
rect 28 157 29 158
rect 27 157 28 158
rect 26 157 27 158
rect 25 157 26 158
rect 24 157 25 158
rect 23 157 24 158
rect 22 157 23 158
rect 21 157 22 158
rect 20 157 21 158
rect 19 157 20 158
rect 18 157 19 158
rect 144 158 145 159
rect 143 158 144 159
rect 142 158 143 159
rect 141 158 142 159
rect 140 158 141 159
rect 139 158 140 159
rect 138 158 139 159
rect 83 158 84 159
rect 82 158 83 159
rect 81 158 82 159
rect 80 158 81 159
rect 79 158 80 159
rect 78 158 79 159
rect 77 158 78 159
rect 76 158 77 159
rect 75 158 76 159
rect 74 158 75 159
rect 73 158 74 159
rect 72 158 73 159
rect 71 158 72 159
rect 70 158 71 159
rect 69 158 70 159
rect 68 158 69 159
rect 67 158 68 159
rect 66 158 67 159
rect 65 158 66 159
rect 64 158 65 159
rect 63 158 64 159
rect 62 158 63 159
rect 61 158 62 159
rect 60 158 61 159
rect 59 158 60 159
rect 58 158 59 159
rect 57 158 58 159
rect 56 158 57 159
rect 55 158 56 159
rect 54 158 55 159
rect 53 158 54 159
rect 52 158 53 159
rect 51 158 52 159
rect 50 158 51 159
rect 49 158 50 159
rect 48 158 49 159
rect 47 158 48 159
rect 46 158 47 159
rect 45 158 46 159
rect 44 158 45 159
rect 43 158 44 159
rect 42 158 43 159
rect 41 158 42 159
rect 40 158 41 159
rect 39 158 40 159
rect 38 158 39 159
rect 37 158 38 159
rect 36 158 37 159
rect 35 158 36 159
rect 34 158 35 159
rect 33 158 34 159
rect 32 158 33 159
rect 31 158 32 159
rect 30 158 31 159
rect 29 158 30 159
rect 28 158 29 159
rect 27 158 28 159
rect 26 158 27 159
rect 25 158 26 159
rect 24 158 25 159
rect 23 158 24 159
rect 22 158 23 159
rect 21 158 22 159
rect 20 158 21 159
rect 19 158 20 159
rect 18 158 19 159
rect 145 159 146 160
rect 144 159 145 160
rect 143 159 144 160
rect 142 159 143 160
rect 141 159 142 160
rect 140 159 141 160
rect 139 159 140 160
rect 138 159 139 160
rect 137 159 138 160
rect 133 159 134 160
rect 132 159 133 160
rect 131 159 132 160
rect 130 159 131 160
rect 129 159 130 160
rect 83 159 84 160
rect 82 159 83 160
rect 81 159 82 160
rect 80 159 81 160
rect 79 159 80 160
rect 78 159 79 160
rect 77 159 78 160
rect 76 159 77 160
rect 75 159 76 160
rect 74 159 75 160
rect 73 159 74 160
rect 72 159 73 160
rect 71 159 72 160
rect 70 159 71 160
rect 69 159 70 160
rect 68 159 69 160
rect 67 159 68 160
rect 66 159 67 160
rect 65 159 66 160
rect 64 159 65 160
rect 63 159 64 160
rect 62 159 63 160
rect 61 159 62 160
rect 60 159 61 160
rect 59 159 60 160
rect 58 159 59 160
rect 57 159 58 160
rect 56 159 57 160
rect 55 159 56 160
rect 54 159 55 160
rect 53 159 54 160
rect 52 159 53 160
rect 51 159 52 160
rect 50 159 51 160
rect 49 159 50 160
rect 48 159 49 160
rect 47 159 48 160
rect 46 159 47 160
rect 45 159 46 160
rect 44 159 45 160
rect 43 159 44 160
rect 42 159 43 160
rect 41 159 42 160
rect 40 159 41 160
rect 39 159 40 160
rect 38 159 39 160
rect 37 159 38 160
rect 36 159 37 160
rect 35 159 36 160
rect 34 159 35 160
rect 33 159 34 160
rect 32 159 33 160
rect 31 159 32 160
rect 30 159 31 160
rect 29 159 30 160
rect 28 159 29 160
rect 27 159 28 160
rect 26 159 27 160
rect 25 159 26 160
rect 24 159 25 160
rect 23 159 24 160
rect 22 159 23 160
rect 21 159 22 160
rect 20 159 21 160
rect 19 159 20 160
rect 18 159 19 160
rect 146 160 147 161
rect 145 160 146 161
rect 144 160 145 161
rect 143 160 144 161
rect 142 160 143 161
rect 141 160 142 161
rect 140 160 141 161
rect 139 160 140 161
rect 138 160 139 161
rect 137 160 138 161
rect 136 160 137 161
rect 132 160 133 161
rect 131 160 132 161
rect 130 160 131 161
rect 129 160 130 161
rect 84 160 85 161
rect 83 160 84 161
rect 82 160 83 161
rect 81 160 82 161
rect 80 160 81 161
rect 79 160 80 161
rect 78 160 79 161
rect 77 160 78 161
rect 76 160 77 161
rect 75 160 76 161
rect 74 160 75 161
rect 73 160 74 161
rect 72 160 73 161
rect 71 160 72 161
rect 70 160 71 161
rect 69 160 70 161
rect 68 160 69 161
rect 67 160 68 161
rect 66 160 67 161
rect 65 160 66 161
rect 64 160 65 161
rect 63 160 64 161
rect 62 160 63 161
rect 61 160 62 161
rect 60 160 61 161
rect 59 160 60 161
rect 58 160 59 161
rect 57 160 58 161
rect 56 160 57 161
rect 55 160 56 161
rect 54 160 55 161
rect 53 160 54 161
rect 52 160 53 161
rect 51 160 52 161
rect 50 160 51 161
rect 49 160 50 161
rect 48 160 49 161
rect 47 160 48 161
rect 46 160 47 161
rect 45 160 46 161
rect 44 160 45 161
rect 43 160 44 161
rect 42 160 43 161
rect 41 160 42 161
rect 40 160 41 161
rect 39 160 40 161
rect 38 160 39 161
rect 37 160 38 161
rect 36 160 37 161
rect 35 160 36 161
rect 34 160 35 161
rect 33 160 34 161
rect 32 160 33 161
rect 31 160 32 161
rect 30 160 31 161
rect 29 160 30 161
rect 28 160 29 161
rect 27 160 28 161
rect 26 160 27 161
rect 25 160 26 161
rect 24 160 25 161
rect 23 160 24 161
rect 22 160 23 161
rect 21 160 22 161
rect 20 160 21 161
rect 19 160 20 161
rect 18 160 19 161
rect 146 161 147 162
rect 145 161 146 162
rect 144 161 145 162
rect 143 161 144 162
rect 142 161 143 162
rect 141 161 142 162
rect 140 161 141 162
rect 139 161 140 162
rect 138 161 139 162
rect 137 161 138 162
rect 136 161 137 162
rect 132 161 133 162
rect 131 161 132 162
rect 130 161 131 162
rect 129 161 130 162
rect 84 161 85 162
rect 83 161 84 162
rect 82 161 83 162
rect 81 161 82 162
rect 80 161 81 162
rect 79 161 80 162
rect 78 161 79 162
rect 77 161 78 162
rect 76 161 77 162
rect 75 161 76 162
rect 74 161 75 162
rect 73 161 74 162
rect 72 161 73 162
rect 71 161 72 162
rect 70 161 71 162
rect 69 161 70 162
rect 68 161 69 162
rect 67 161 68 162
rect 66 161 67 162
rect 65 161 66 162
rect 64 161 65 162
rect 63 161 64 162
rect 62 161 63 162
rect 61 161 62 162
rect 60 161 61 162
rect 59 161 60 162
rect 58 161 59 162
rect 57 161 58 162
rect 56 161 57 162
rect 55 161 56 162
rect 54 161 55 162
rect 53 161 54 162
rect 52 161 53 162
rect 51 161 52 162
rect 50 161 51 162
rect 49 161 50 162
rect 48 161 49 162
rect 47 161 48 162
rect 46 161 47 162
rect 45 161 46 162
rect 44 161 45 162
rect 43 161 44 162
rect 42 161 43 162
rect 41 161 42 162
rect 40 161 41 162
rect 39 161 40 162
rect 38 161 39 162
rect 37 161 38 162
rect 36 161 37 162
rect 35 161 36 162
rect 34 161 35 162
rect 33 161 34 162
rect 32 161 33 162
rect 31 161 32 162
rect 30 161 31 162
rect 29 161 30 162
rect 28 161 29 162
rect 27 161 28 162
rect 26 161 27 162
rect 25 161 26 162
rect 24 161 25 162
rect 23 161 24 162
rect 22 161 23 162
rect 21 161 22 162
rect 20 161 21 162
rect 19 161 20 162
rect 18 161 19 162
rect 146 162 147 163
rect 145 162 146 163
rect 144 162 145 163
rect 143 162 144 163
rect 142 162 143 163
rect 139 162 140 163
rect 138 162 139 163
rect 137 162 138 163
rect 136 162 137 163
rect 131 162 132 163
rect 130 162 131 163
rect 129 162 130 163
rect 128 162 129 163
rect 84 162 85 163
rect 83 162 84 163
rect 82 162 83 163
rect 81 162 82 163
rect 80 162 81 163
rect 79 162 80 163
rect 78 162 79 163
rect 77 162 78 163
rect 76 162 77 163
rect 75 162 76 163
rect 74 162 75 163
rect 73 162 74 163
rect 72 162 73 163
rect 71 162 72 163
rect 70 162 71 163
rect 69 162 70 163
rect 68 162 69 163
rect 67 162 68 163
rect 66 162 67 163
rect 65 162 66 163
rect 64 162 65 163
rect 63 162 64 163
rect 62 162 63 163
rect 61 162 62 163
rect 60 162 61 163
rect 59 162 60 163
rect 58 162 59 163
rect 57 162 58 163
rect 56 162 57 163
rect 55 162 56 163
rect 54 162 55 163
rect 53 162 54 163
rect 52 162 53 163
rect 51 162 52 163
rect 50 162 51 163
rect 49 162 50 163
rect 48 162 49 163
rect 47 162 48 163
rect 46 162 47 163
rect 45 162 46 163
rect 44 162 45 163
rect 43 162 44 163
rect 42 162 43 163
rect 41 162 42 163
rect 40 162 41 163
rect 39 162 40 163
rect 38 162 39 163
rect 37 162 38 163
rect 36 162 37 163
rect 35 162 36 163
rect 34 162 35 163
rect 33 162 34 163
rect 32 162 33 163
rect 31 162 32 163
rect 30 162 31 163
rect 29 162 30 163
rect 28 162 29 163
rect 27 162 28 163
rect 26 162 27 163
rect 25 162 26 163
rect 24 162 25 163
rect 23 162 24 163
rect 22 162 23 163
rect 21 162 22 163
rect 20 162 21 163
rect 19 162 20 163
rect 18 162 19 163
rect 146 163 147 164
rect 145 163 146 164
rect 144 163 145 164
rect 143 163 144 164
rect 138 163 139 164
rect 137 163 138 164
rect 136 163 137 164
rect 135 163 136 164
rect 131 163 132 164
rect 130 163 131 164
rect 129 163 130 164
rect 128 163 129 164
rect 84 163 85 164
rect 83 163 84 164
rect 82 163 83 164
rect 81 163 82 164
rect 80 163 81 164
rect 79 163 80 164
rect 78 163 79 164
rect 77 163 78 164
rect 76 163 77 164
rect 75 163 76 164
rect 74 163 75 164
rect 73 163 74 164
rect 72 163 73 164
rect 71 163 72 164
rect 70 163 71 164
rect 69 163 70 164
rect 68 163 69 164
rect 67 163 68 164
rect 66 163 67 164
rect 65 163 66 164
rect 64 163 65 164
rect 63 163 64 164
rect 62 163 63 164
rect 146 164 147 165
rect 145 164 146 165
rect 144 164 145 165
rect 143 164 144 165
rect 137 164 138 165
rect 136 164 137 165
rect 135 164 136 165
rect 131 164 132 165
rect 130 164 131 165
rect 129 164 130 165
rect 128 164 129 165
rect 84 164 85 165
rect 83 164 84 165
rect 82 164 83 165
rect 81 164 82 165
rect 80 164 81 165
rect 79 164 80 165
rect 78 164 79 165
rect 77 164 78 165
rect 76 164 77 165
rect 75 164 76 165
rect 74 164 75 165
rect 73 164 74 165
rect 72 164 73 165
rect 71 164 72 165
rect 70 164 71 165
rect 69 164 70 165
rect 68 164 69 165
rect 67 164 68 165
rect 66 164 67 165
rect 65 164 66 165
rect 145 165 146 166
rect 144 165 145 166
rect 143 165 144 166
rect 137 165 138 166
rect 136 165 137 166
rect 135 165 136 166
rect 131 165 132 166
rect 130 165 131 166
rect 129 165 130 166
rect 128 165 129 166
rect 85 165 86 166
rect 84 165 85 166
rect 83 165 84 166
rect 82 165 83 166
rect 81 165 82 166
rect 80 165 81 166
rect 79 165 80 166
rect 78 165 79 166
rect 77 165 78 166
rect 76 165 77 166
rect 75 165 76 166
rect 74 165 75 166
rect 73 165 74 166
rect 72 165 73 166
rect 71 165 72 166
rect 70 165 71 166
rect 69 165 70 166
rect 68 165 69 166
rect 67 165 68 166
rect 66 165 67 166
rect 145 166 146 167
rect 144 166 145 167
rect 143 166 144 167
rect 137 166 138 167
rect 136 166 137 167
rect 135 166 136 167
rect 131 166 132 167
rect 130 166 131 167
rect 129 166 130 167
rect 128 166 129 167
rect 85 166 86 167
rect 84 166 85 167
rect 83 166 84 167
rect 82 166 83 167
rect 81 166 82 167
rect 80 166 81 167
rect 79 166 80 167
rect 78 166 79 167
rect 77 166 78 167
rect 76 166 77 167
rect 75 166 76 167
rect 74 166 75 167
rect 73 166 74 167
rect 72 166 73 167
rect 71 166 72 167
rect 70 166 71 167
rect 69 166 70 167
rect 68 166 69 167
rect 67 166 68 167
rect 144 167 145 168
rect 143 167 144 168
rect 142 167 143 168
rect 137 167 138 168
rect 136 167 137 168
rect 135 167 136 168
rect 131 167 132 168
rect 130 167 131 168
rect 129 167 130 168
rect 128 167 129 168
rect 85 167 86 168
rect 84 167 85 168
rect 83 167 84 168
rect 82 167 83 168
rect 81 167 82 168
rect 80 167 81 168
rect 79 167 80 168
rect 78 167 79 168
rect 77 167 78 168
rect 76 167 77 168
rect 75 167 76 168
rect 74 167 75 168
rect 73 167 74 168
rect 72 167 73 168
rect 71 167 72 168
rect 70 167 71 168
rect 69 167 70 168
rect 68 167 69 168
rect 144 168 145 169
rect 143 168 144 169
rect 142 168 143 169
rect 141 168 142 169
rect 140 168 141 169
rect 137 168 138 169
rect 136 168 137 169
rect 135 168 136 169
rect 134 168 135 169
rect 133 168 134 169
rect 132 168 133 169
rect 131 168 132 169
rect 130 168 131 169
rect 129 168 130 169
rect 128 168 129 169
rect 85 168 86 169
rect 84 168 85 169
rect 83 168 84 169
rect 82 168 83 169
rect 81 168 82 169
rect 80 168 81 169
rect 79 168 80 169
rect 78 168 79 169
rect 77 168 78 169
rect 76 168 77 169
rect 75 168 76 169
rect 74 168 75 169
rect 73 168 74 169
rect 72 168 73 169
rect 71 168 72 169
rect 70 168 71 169
rect 69 168 70 169
rect 68 168 69 169
rect 146 169 147 170
rect 145 169 146 170
rect 144 169 145 170
rect 143 169 144 170
rect 142 169 143 170
rect 141 169 142 170
rect 140 169 141 170
rect 139 169 140 170
rect 138 169 139 170
rect 137 169 138 170
rect 136 169 137 170
rect 135 169 136 170
rect 134 169 135 170
rect 133 169 134 170
rect 132 169 133 170
rect 131 169 132 170
rect 130 169 131 170
rect 129 169 130 170
rect 85 169 86 170
rect 84 169 85 170
rect 83 169 84 170
rect 82 169 83 170
rect 81 169 82 170
rect 80 169 81 170
rect 79 169 80 170
rect 78 169 79 170
rect 77 169 78 170
rect 76 169 77 170
rect 75 169 76 170
rect 74 169 75 170
rect 73 169 74 170
rect 72 169 73 170
rect 71 169 72 170
rect 70 169 71 170
rect 69 169 70 170
rect 146 170 147 171
rect 145 170 146 171
rect 144 170 145 171
rect 143 170 144 171
rect 142 170 143 171
rect 141 170 142 171
rect 140 170 141 171
rect 139 170 140 171
rect 138 170 139 171
rect 137 170 138 171
rect 136 170 137 171
rect 135 170 136 171
rect 134 170 135 171
rect 133 170 134 171
rect 132 170 133 171
rect 131 170 132 171
rect 130 170 131 171
rect 129 170 130 171
rect 85 170 86 171
rect 84 170 85 171
rect 83 170 84 171
rect 82 170 83 171
rect 81 170 82 171
rect 80 170 81 171
rect 79 170 80 171
rect 78 170 79 171
rect 77 170 78 171
rect 76 170 77 171
rect 75 170 76 171
rect 74 170 75 171
rect 73 170 74 171
rect 72 170 73 171
rect 71 170 72 171
rect 70 170 71 171
rect 69 170 70 171
rect 146 171 147 172
rect 145 171 146 172
rect 144 171 145 172
rect 143 171 144 172
rect 142 171 143 172
rect 141 171 142 172
rect 140 171 141 172
rect 139 171 140 172
rect 138 171 139 172
rect 137 171 138 172
rect 136 171 137 172
rect 135 171 136 172
rect 134 171 135 172
rect 133 171 134 172
rect 132 171 133 172
rect 131 171 132 172
rect 130 171 131 172
rect 85 171 86 172
rect 84 171 85 172
rect 83 171 84 172
rect 82 171 83 172
rect 81 171 82 172
rect 80 171 81 172
rect 79 171 80 172
rect 78 171 79 172
rect 77 171 78 172
rect 76 171 77 172
rect 75 171 76 172
rect 74 171 75 172
rect 73 171 74 172
rect 72 171 73 172
rect 71 171 72 172
rect 70 171 71 172
rect 69 171 70 172
rect 146 172 147 173
rect 145 172 146 173
rect 144 172 145 173
rect 143 172 144 173
rect 142 172 143 173
rect 141 172 142 173
rect 140 172 141 173
rect 139 172 140 173
rect 138 172 139 173
rect 137 172 138 173
rect 136 172 137 173
rect 135 172 136 173
rect 134 172 135 173
rect 133 172 134 173
rect 132 172 133 173
rect 131 172 132 173
rect 85 172 86 173
rect 84 172 85 173
rect 83 172 84 173
rect 82 172 83 173
rect 81 172 82 173
rect 80 172 81 173
rect 79 172 80 173
rect 78 172 79 173
rect 77 172 78 173
rect 76 172 77 173
rect 75 172 76 173
rect 74 172 75 173
rect 73 172 74 173
rect 72 172 73 173
rect 71 172 72 173
rect 70 172 71 173
rect 69 172 70 173
rect 146 173 147 174
rect 145 173 146 174
rect 144 173 145 174
rect 143 173 144 174
rect 142 173 143 174
rect 141 173 142 174
rect 140 173 141 174
rect 139 173 140 174
rect 138 173 139 174
rect 137 173 138 174
rect 136 173 137 174
rect 135 173 136 174
rect 134 173 135 174
rect 133 173 134 174
rect 85 173 86 174
rect 84 173 85 174
rect 83 173 84 174
rect 82 173 83 174
rect 81 173 82 174
rect 80 173 81 174
rect 79 173 80 174
rect 78 173 79 174
rect 77 173 78 174
rect 76 173 77 174
rect 75 173 76 174
rect 74 173 75 174
rect 73 173 74 174
rect 72 173 73 174
rect 71 173 72 174
rect 70 173 71 174
rect 69 173 70 174
rect 85 174 86 175
rect 84 174 85 175
rect 83 174 84 175
rect 82 174 83 175
rect 81 174 82 175
rect 80 174 81 175
rect 79 174 80 175
rect 78 174 79 175
rect 77 174 78 175
rect 76 174 77 175
rect 75 174 76 175
rect 74 174 75 175
rect 73 174 74 175
rect 72 174 73 175
rect 71 174 72 175
rect 70 174 71 175
rect 69 174 70 175
rect 85 175 86 176
rect 84 175 85 176
rect 83 175 84 176
rect 82 175 83 176
rect 81 175 82 176
rect 80 175 81 176
rect 79 175 80 176
rect 78 175 79 176
rect 77 175 78 176
rect 76 175 77 176
rect 75 175 76 176
rect 74 175 75 176
rect 73 175 74 176
rect 72 175 73 176
rect 71 175 72 176
rect 70 175 71 176
rect 69 175 70 176
rect 68 175 69 176
rect 85 176 86 177
rect 84 176 85 177
rect 83 176 84 177
rect 82 176 83 177
rect 81 176 82 177
rect 80 176 81 177
rect 79 176 80 177
rect 78 176 79 177
rect 77 176 78 177
rect 76 176 77 177
rect 75 176 76 177
rect 74 176 75 177
rect 73 176 74 177
rect 72 176 73 177
rect 71 176 72 177
rect 70 176 71 177
rect 69 176 70 177
rect 68 176 69 177
rect 85 177 86 178
rect 84 177 85 178
rect 83 177 84 178
rect 82 177 83 178
rect 81 177 82 178
rect 80 177 81 178
rect 79 177 80 178
rect 78 177 79 178
rect 77 177 78 178
rect 76 177 77 178
rect 75 177 76 178
rect 74 177 75 178
rect 73 177 74 178
rect 72 177 73 178
rect 71 177 72 178
rect 70 177 71 178
rect 69 177 70 178
rect 68 177 69 178
rect 67 177 68 178
rect 84 178 85 179
rect 83 178 84 179
rect 82 178 83 179
rect 81 178 82 179
rect 80 178 81 179
rect 79 178 80 179
rect 78 178 79 179
rect 77 178 78 179
rect 76 178 77 179
rect 75 178 76 179
rect 74 178 75 179
rect 73 178 74 179
rect 72 178 73 179
rect 71 178 72 179
rect 70 178 71 179
rect 69 178 70 179
rect 68 178 69 179
rect 67 178 68 179
rect 66 178 67 179
rect 146 179 147 180
rect 145 179 146 180
rect 144 179 145 180
rect 143 179 144 180
rect 142 179 143 180
rect 141 179 142 180
rect 140 179 141 180
rect 139 179 140 180
rect 138 179 139 180
rect 137 179 138 180
rect 136 179 137 180
rect 135 179 136 180
rect 134 179 135 180
rect 133 179 134 180
rect 132 179 133 180
rect 131 179 132 180
rect 130 179 131 180
rect 129 179 130 180
rect 128 179 129 180
rect 84 179 85 180
rect 83 179 84 180
rect 82 179 83 180
rect 81 179 82 180
rect 80 179 81 180
rect 79 179 80 180
rect 78 179 79 180
rect 77 179 78 180
rect 76 179 77 180
rect 75 179 76 180
rect 74 179 75 180
rect 73 179 74 180
rect 72 179 73 180
rect 71 179 72 180
rect 70 179 71 180
rect 69 179 70 180
rect 68 179 69 180
rect 67 179 68 180
rect 66 179 67 180
rect 65 179 66 180
rect 146 180 147 181
rect 145 180 146 181
rect 144 180 145 181
rect 143 180 144 181
rect 142 180 143 181
rect 141 180 142 181
rect 140 180 141 181
rect 139 180 140 181
rect 138 180 139 181
rect 137 180 138 181
rect 136 180 137 181
rect 135 180 136 181
rect 134 180 135 181
rect 133 180 134 181
rect 132 180 133 181
rect 131 180 132 181
rect 130 180 131 181
rect 129 180 130 181
rect 128 180 129 181
rect 84 180 85 181
rect 83 180 84 181
rect 82 180 83 181
rect 81 180 82 181
rect 80 180 81 181
rect 79 180 80 181
rect 78 180 79 181
rect 77 180 78 181
rect 76 180 77 181
rect 75 180 76 181
rect 74 180 75 181
rect 73 180 74 181
rect 72 180 73 181
rect 71 180 72 181
rect 70 180 71 181
rect 69 180 70 181
rect 68 180 69 181
rect 67 180 68 181
rect 66 180 67 181
rect 65 180 66 181
rect 64 180 65 181
rect 63 180 64 181
rect 62 180 63 181
rect 146 181 147 182
rect 145 181 146 182
rect 144 181 145 182
rect 143 181 144 182
rect 142 181 143 182
rect 141 181 142 182
rect 140 181 141 182
rect 139 181 140 182
rect 138 181 139 182
rect 137 181 138 182
rect 136 181 137 182
rect 135 181 136 182
rect 134 181 135 182
rect 133 181 134 182
rect 132 181 133 182
rect 131 181 132 182
rect 130 181 131 182
rect 129 181 130 182
rect 128 181 129 182
rect 84 181 85 182
rect 83 181 84 182
rect 82 181 83 182
rect 81 181 82 182
rect 80 181 81 182
rect 79 181 80 182
rect 78 181 79 182
rect 77 181 78 182
rect 76 181 77 182
rect 75 181 76 182
rect 74 181 75 182
rect 73 181 74 182
rect 72 181 73 182
rect 71 181 72 182
rect 70 181 71 182
rect 69 181 70 182
rect 68 181 69 182
rect 67 181 68 182
rect 66 181 67 182
rect 65 181 66 182
rect 64 181 65 182
rect 63 181 64 182
rect 62 181 63 182
rect 61 181 62 182
rect 60 181 61 182
rect 59 181 60 182
rect 58 181 59 182
rect 57 181 58 182
rect 56 181 57 182
rect 55 181 56 182
rect 54 181 55 182
rect 53 181 54 182
rect 52 181 53 182
rect 51 181 52 182
rect 50 181 51 182
rect 49 181 50 182
rect 48 181 49 182
rect 47 181 48 182
rect 46 181 47 182
rect 45 181 46 182
rect 44 181 45 182
rect 43 181 44 182
rect 42 181 43 182
rect 41 181 42 182
rect 40 181 41 182
rect 39 181 40 182
rect 38 181 39 182
rect 37 181 38 182
rect 36 181 37 182
rect 35 181 36 182
rect 34 181 35 182
rect 33 181 34 182
rect 32 181 33 182
rect 31 181 32 182
rect 30 181 31 182
rect 29 181 30 182
rect 28 181 29 182
rect 27 181 28 182
rect 26 181 27 182
rect 25 181 26 182
rect 24 181 25 182
rect 23 181 24 182
rect 22 181 23 182
rect 21 181 22 182
rect 20 181 21 182
rect 19 181 20 182
rect 18 181 19 182
rect 146 182 147 183
rect 145 182 146 183
rect 144 182 145 183
rect 143 182 144 183
rect 142 182 143 183
rect 141 182 142 183
rect 140 182 141 183
rect 139 182 140 183
rect 138 182 139 183
rect 137 182 138 183
rect 136 182 137 183
rect 135 182 136 183
rect 134 182 135 183
rect 133 182 134 183
rect 132 182 133 183
rect 131 182 132 183
rect 130 182 131 183
rect 129 182 130 183
rect 128 182 129 183
rect 84 182 85 183
rect 83 182 84 183
rect 82 182 83 183
rect 81 182 82 183
rect 80 182 81 183
rect 79 182 80 183
rect 78 182 79 183
rect 77 182 78 183
rect 76 182 77 183
rect 75 182 76 183
rect 74 182 75 183
rect 73 182 74 183
rect 72 182 73 183
rect 71 182 72 183
rect 70 182 71 183
rect 69 182 70 183
rect 68 182 69 183
rect 67 182 68 183
rect 66 182 67 183
rect 65 182 66 183
rect 64 182 65 183
rect 63 182 64 183
rect 62 182 63 183
rect 61 182 62 183
rect 60 182 61 183
rect 59 182 60 183
rect 58 182 59 183
rect 57 182 58 183
rect 56 182 57 183
rect 55 182 56 183
rect 54 182 55 183
rect 53 182 54 183
rect 52 182 53 183
rect 51 182 52 183
rect 50 182 51 183
rect 49 182 50 183
rect 48 182 49 183
rect 47 182 48 183
rect 46 182 47 183
rect 45 182 46 183
rect 44 182 45 183
rect 43 182 44 183
rect 42 182 43 183
rect 41 182 42 183
rect 40 182 41 183
rect 39 182 40 183
rect 38 182 39 183
rect 37 182 38 183
rect 36 182 37 183
rect 35 182 36 183
rect 34 182 35 183
rect 33 182 34 183
rect 32 182 33 183
rect 31 182 32 183
rect 30 182 31 183
rect 29 182 30 183
rect 28 182 29 183
rect 27 182 28 183
rect 26 182 27 183
rect 25 182 26 183
rect 24 182 25 183
rect 23 182 24 183
rect 22 182 23 183
rect 21 182 22 183
rect 20 182 21 183
rect 19 182 20 183
rect 18 182 19 183
rect 146 183 147 184
rect 145 183 146 184
rect 144 183 145 184
rect 143 183 144 184
rect 142 183 143 184
rect 141 183 142 184
rect 140 183 141 184
rect 139 183 140 184
rect 138 183 139 184
rect 137 183 138 184
rect 136 183 137 184
rect 135 183 136 184
rect 134 183 135 184
rect 133 183 134 184
rect 132 183 133 184
rect 131 183 132 184
rect 130 183 131 184
rect 129 183 130 184
rect 128 183 129 184
rect 83 183 84 184
rect 82 183 83 184
rect 81 183 82 184
rect 80 183 81 184
rect 79 183 80 184
rect 78 183 79 184
rect 77 183 78 184
rect 76 183 77 184
rect 75 183 76 184
rect 74 183 75 184
rect 73 183 74 184
rect 72 183 73 184
rect 71 183 72 184
rect 70 183 71 184
rect 69 183 70 184
rect 68 183 69 184
rect 67 183 68 184
rect 66 183 67 184
rect 65 183 66 184
rect 64 183 65 184
rect 63 183 64 184
rect 62 183 63 184
rect 61 183 62 184
rect 60 183 61 184
rect 59 183 60 184
rect 58 183 59 184
rect 57 183 58 184
rect 56 183 57 184
rect 55 183 56 184
rect 54 183 55 184
rect 53 183 54 184
rect 52 183 53 184
rect 51 183 52 184
rect 50 183 51 184
rect 49 183 50 184
rect 48 183 49 184
rect 47 183 48 184
rect 46 183 47 184
rect 45 183 46 184
rect 44 183 45 184
rect 43 183 44 184
rect 42 183 43 184
rect 41 183 42 184
rect 40 183 41 184
rect 39 183 40 184
rect 38 183 39 184
rect 37 183 38 184
rect 36 183 37 184
rect 35 183 36 184
rect 34 183 35 184
rect 33 183 34 184
rect 32 183 33 184
rect 31 183 32 184
rect 30 183 31 184
rect 29 183 30 184
rect 28 183 29 184
rect 27 183 28 184
rect 26 183 27 184
rect 25 183 26 184
rect 24 183 25 184
rect 23 183 24 184
rect 22 183 23 184
rect 21 183 22 184
rect 20 183 21 184
rect 19 183 20 184
rect 18 183 19 184
rect 133 184 134 185
rect 132 184 133 185
rect 131 184 132 185
rect 83 184 84 185
rect 82 184 83 185
rect 81 184 82 185
rect 80 184 81 185
rect 79 184 80 185
rect 78 184 79 185
rect 77 184 78 185
rect 76 184 77 185
rect 75 184 76 185
rect 74 184 75 185
rect 73 184 74 185
rect 72 184 73 185
rect 71 184 72 185
rect 70 184 71 185
rect 69 184 70 185
rect 68 184 69 185
rect 67 184 68 185
rect 66 184 67 185
rect 65 184 66 185
rect 64 184 65 185
rect 63 184 64 185
rect 62 184 63 185
rect 61 184 62 185
rect 60 184 61 185
rect 59 184 60 185
rect 58 184 59 185
rect 57 184 58 185
rect 56 184 57 185
rect 55 184 56 185
rect 54 184 55 185
rect 53 184 54 185
rect 52 184 53 185
rect 51 184 52 185
rect 50 184 51 185
rect 49 184 50 185
rect 48 184 49 185
rect 47 184 48 185
rect 46 184 47 185
rect 45 184 46 185
rect 44 184 45 185
rect 43 184 44 185
rect 42 184 43 185
rect 41 184 42 185
rect 40 184 41 185
rect 39 184 40 185
rect 38 184 39 185
rect 37 184 38 185
rect 36 184 37 185
rect 35 184 36 185
rect 34 184 35 185
rect 33 184 34 185
rect 32 184 33 185
rect 31 184 32 185
rect 30 184 31 185
rect 29 184 30 185
rect 28 184 29 185
rect 27 184 28 185
rect 26 184 27 185
rect 25 184 26 185
rect 24 184 25 185
rect 23 184 24 185
rect 22 184 23 185
rect 21 184 22 185
rect 20 184 21 185
rect 19 184 20 185
rect 18 184 19 185
rect 132 185 133 186
rect 131 185 132 186
rect 130 185 131 186
rect 83 185 84 186
rect 82 185 83 186
rect 81 185 82 186
rect 80 185 81 186
rect 79 185 80 186
rect 78 185 79 186
rect 77 185 78 186
rect 76 185 77 186
rect 75 185 76 186
rect 74 185 75 186
rect 73 185 74 186
rect 72 185 73 186
rect 71 185 72 186
rect 70 185 71 186
rect 69 185 70 186
rect 68 185 69 186
rect 67 185 68 186
rect 66 185 67 186
rect 65 185 66 186
rect 64 185 65 186
rect 63 185 64 186
rect 62 185 63 186
rect 61 185 62 186
rect 60 185 61 186
rect 59 185 60 186
rect 58 185 59 186
rect 57 185 58 186
rect 56 185 57 186
rect 55 185 56 186
rect 54 185 55 186
rect 53 185 54 186
rect 52 185 53 186
rect 51 185 52 186
rect 50 185 51 186
rect 49 185 50 186
rect 48 185 49 186
rect 47 185 48 186
rect 46 185 47 186
rect 45 185 46 186
rect 44 185 45 186
rect 43 185 44 186
rect 42 185 43 186
rect 41 185 42 186
rect 40 185 41 186
rect 39 185 40 186
rect 38 185 39 186
rect 37 185 38 186
rect 36 185 37 186
rect 35 185 36 186
rect 34 185 35 186
rect 33 185 34 186
rect 32 185 33 186
rect 31 185 32 186
rect 30 185 31 186
rect 29 185 30 186
rect 28 185 29 186
rect 27 185 28 186
rect 26 185 27 186
rect 25 185 26 186
rect 24 185 25 186
rect 23 185 24 186
rect 22 185 23 186
rect 21 185 22 186
rect 20 185 21 186
rect 19 185 20 186
rect 18 185 19 186
rect 132 186 133 187
rect 131 186 132 187
rect 130 186 131 187
rect 129 186 130 187
rect 82 186 83 187
rect 81 186 82 187
rect 80 186 81 187
rect 79 186 80 187
rect 78 186 79 187
rect 77 186 78 187
rect 76 186 77 187
rect 75 186 76 187
rect 74 186 75 187
rect 73 186 74 187
rect 72 186 73 187
rect 71 186 72 187
rect 70 186 71 187
rect 69 186 70 187
rect 68 186 69 187
rect 67 186 68 187
rect 66 186 67 187
rect 65 186 66 187
rect 64 186 65 187
rect 63 186 64 187
rect 62 186 63 187
rect 61 186 62 187
rect 60 186 61 187
rect 59 186 60 187
rect 58 186 59 187
rect 57 186 58 187
rect 56 186 57 187
rect 55 186 56 187
rect 54 186 55 187
rect 53 186 54 187
rect 52 186 53 187
rect 51 186 52 187
rect 50 186 51 187
rect 49 186 50 187
rect 48 186 49 187
rect 47 186 48 187
rect 46 186 47 187
rect 45 186 46 187
rect 44 186 45 187
rect 43 186 44 187
rect 42 186 43 187
rect 41 186 42 187
rect 40 186 41 187
rect 39 186 40 187
rect 38 186 39 187
rect 37 186 38 187
rect 36 186 37 187
rect 35 186 36 187
rect 34 186 35 187
rect 33 186 34 187
rect 32 186 33 187
rect 31 186 32 187
rect 30 186 31 187
rect 29 186 30 187
rect 28 186 29 187
rect 27 186 28 187
rect 26 186 27 187
rect 25 186 26 187
rect 24 186 25 187
rect 23 186 24 187
rect 22 186 23 187
rect 21 186 22 187
rect 20 186 21 187
rect 19 186 20 187
rect 18 186 19 187
rect 131 187 132 188
rect 130 187 131 188
rect 129 187 130 188
rect 82 187 83 188
rect 81 187 82 188
rect 80 187 81 188
rect 79 187 80 188
rect 78 187 79 188
rect 77 187 78 188
rect 76 187 77 188
rect 75 187 76 188
rect 74 187 75 188
rect 73 187 74 188
rect 72 187 73 188
rect 71 187 72 188
rect 70 187 71 188
rect 69 187 70 188
rect 68 187 69 188
rect 67 187 68 188
rect 66 187 67 188
rect 65 187 66 188
rect 64 187 65 188
rect 63 187 64 188
rect 62 187 63 188
rect 61 187 62 188
rect 60 187 61 188
rect 59 187 60 188
rect 58 187 59 188
rect 57 187 58 188
rect 56 187 57 188
rect 55 187 56 188
rect 54 187 55 188
rect 53 187 54 188
rect 52 187 53 188
rect 51 187 52 188
rect 50 187 51 188
rect 49 187 50 188
rect 48 187 49 188
rect 47 187 48 188
rect 46 187 47 188
rect 45 187 46 188
rect 44 187 45 188
rect 43 187 44 188
rect 42 187 43 188
rect 41 187 42 188
rect 40 187 41 188
rect 39 187 40 188
rect 38 187 39 188
rect 37 187 38 188
rect 36 187 37 188
rect 35 187 36 188
rect 34 187 35 188
rect 33 187 34 188
rect 32 187 33 188
rect 31 187 32 188
rect 30 187 31 188
rect 29 187 30 188
rect 28 187 29 188
rect 27 187 28 188
rect 26 187 27 188
rect 25 187 26 188
rect 24 187 25 188
rect 23 187 24 188
rect 22 187 23 188
rect 21 187 22 188
rect 20 187 21 188
rect 19 187 20 188
rect 18 187 19 188
rect 132 188 133 189
rect 131 188 132 189
rect 130 188 131 189
rect 129 188 130 189
rect 128 188 129 189
rect 81 188 82 189
rect 80 188 81 189
rect 79 188 80 189
rect 78 188 79 189
rect 77 188 78 189
rect 76 188 77 189
rect 75 188 76 189
rect 74 188 75 189
rect 73 188 74 189
rect 72 188 73 189
rect 71 188 72 189
rect 70 188 71 189
rect 69 188 70 189
rect 68 188 69 189
rect 67 188 68 189
rect 66 188 67 189
rect 65 188 66 189
rect 64 188 65 189
rect 63 188 64 189
rect 62 188 63 189
rect 61 188 62 189
rect 60 188 61 189
rect 59 188 60 189
rect 58 188 59 189
rect 57 188 58 189
rect 56 188 57 189
rect 55 188 56 189
rect 54 188 55 189
rect 53 188 54 189
rect 52 188 53 189
rect 51 188 52 189
rect 50 188 51 189
rect 49 188 50 189
rect 48 188 49 189
rect 47 188 48 189
rect 46 188 47 189
rect 45 188 46 189
rect 44 188 45 189
rect 43 188 44 189
rect 42 188 43 189
rect 41 188 42 189
rect 40 188 41 189
rect 39 188 40 189
rect 38 188 39 189
rect 37 188 38 189
rect 36 188 37 189
rect 35 188 36 189
rect 34 188 35 189
rect 33 188 34 189
rect 32 188 33 189
rect 31 188 32 189
rect 30 188 31 189
rect 29 188 30 189
rect 28 188 29 189
rect 27 188 28 189
rect 26 188 27 189
rect 25 188 26 189
rect 24 188 25 189
rect 23 188 24 189
rect 22 188 23 189
rect 21 188 22 189
rect 20 188 21 189
rect 19 188 20 189
rect 18 188 19 189
rect 132 189 133 190
rect 131 189 132 190
rect 130 189 131 190
rect 129 189 130 190
rect 128 189 129 190
rect 81 189 82 190
rect 80 189 81 190
rect 79 189 80 190
rect 78 189 79 190
rect 77 189 78 190
rect 76 189 77 190
rect 75 189 76 190
rect 74 189 75 190
rect 73 189 74 190
rect 72 189 73 190
rect 71 189 72 190
rect 70 189 71 190
rect 69 189 70 190
rect 68 189 69 190
rect 67 189 68 190
rect 66 189 67 190
rect 65 189 66 190
rect 64 189 65 190
rect 63 189 64 190
rect 62 189 63 190
rect 61 189 62 190
rect 60 189 61 190
rect 59 189 60 190
rect 58 189 59 190
rect 57 189 58 190
rect 56 189 57 190
rect 55 189 56 190
rect 54 189 55 190
rect 53 189 54 190
rect 52 189 53 190
rect 51 189 52 190
rect 50 189 51 190
rect 49 189 50 190
rect 48 189 49 190
rect 47 189 48 190
rect 46 189 47 190
rect 45 189 46 190
rect 44 189 45 190
rect 43 189 44 190
rect 42 189 43 190
rect 41 189 42 190
rect 40 189 41 190
rect 39 189 40 190
rect 38 189 39 190
rect 37 189 38 190
rect 36 189 37 190
rect 35 189 36 190
rect 34 189 35 190
rect 33 189 34 190
rect 32 189 33 190
rect 31 189 32 190
rect 30 189 31 190
rect 29 189 30 190
rect 28 189 29 190
rect 27 189 28 190
rect 26 189 27 190
rect 25 189 26 190
rect 24 189 25 190
rect 23 189 24 190
rect 22 189 23 190
rect 21 189 22 190
rect 20 189 21 190
rect 19 189 20 190
rect 18 189 19 190
rect 134 190 135 191
rect 133 190 134 191
rect 132 190 133 191
rect 131 190 132 191
rect 130 190 131 191
rect 129 190 130 191
rect 128 190 129 191
rect 80 190 81 191
rect 79 190 80 191
rect 78 190 79 191
rect 77 190 78 191
rect 76 190 77 191
rect 75 190 76 191
rect 74 190 75 191
rect 73 190 74 191
rect 72 190 73 191
rect 71 190 72 191
rect 70 190 71 191
rect 69 190 70 191
rect 68 190 69 191
rect 67 190 68 191
rect 66 190 67 191
rect 65 190 66 191
rect 64 190 65 191
rect 63 190 64 191
rect 62 190 63 191
rect 61 190 62 191
rect 60 190 61 191
rect 59 190 60 191
rect 58 190 59 191
rect 57 190 58 191
rect 56 190 57 191
rect 55 190 56 191
rect 54 190 55 191
rect 53 190 54 191
rect 52 190 53 191
rect 51 190 52 191
rect 50 190 51 191
rect 49 190 50 191
rect 48 190 49 191
rect 47 190 48 191
rect 46 190 47 191
rect 45 190 46 191
rect 44 190 45 191
rect 43 190 44 191
rect 42 190 43 191
rect 41 190 42 191
rect 40 190 41 191
rect 39 190 40 191
rect 38 190 39 191
rect 37 190 38 191
rect 36 190 37 191
rect 35 190 36 191
rect 34 190 35 191
rect 33 190 34 191
rect 32 190 33 191
rect 31 190 32 191
rect 30 190 31 191
rect 29 190 30 191
rect 28 190 29 191
rect 27 190 28 191
rect 26 190 27 191
rect 25 190 26 191
rect 24 190 25 191
rect 23 190 24 191
rect 22 190 23 191
rect 21 190 22 191
rect 20 190 21 191
rect 19 190 20 191
rect 18 190 19 191
rect 146 191 147 192
rect 145 191 146 192
rect 144 191 145 192
rect 143 191 144 192
rect 142 191 143 192
rect 141 191 142 192
rect 140 191 141 192
rect 139 191 140 192
rect 138 191 139 192
rect 137 191 138 192
rect 136 191 137 192
rect 135 191 136 192
rect 134 191 135 192
rect 133 191 134 192
rect 132 191 133 192
rect 131 191 132 192
rect 130 191 131 192
rect 129 191 130 192
rect 128 191 129 192
rect 80 191 81 192
rect 79 191 80 192
rect 78 191 79 192
rect 77 191 78 192
rect 76 191 77 192
rect 75 191 76 192
rect 74 191 75 192
rect 73 191 74 192
rect 72 191 73 192
rect 71 191 72 192
rect 70 191 71 192
rect 69 191 70 192
rect 68 191 69 192
rect 67 191 68 192
rect 66 191 67 192
rect 65 191 66 192
rect 64 191 65 192
rect 63 191 64 192
rect 62 191 63 192
rect 61 191 62 192
rect 60 191 61 192
rect 59 191 60 192
rect 58 191 59 192
rect 57 191 58 192
rect 56 191 57 192
rect 55 191 56 192
rect 54 191 55 192
rect 53 191 54 192
rect 52 191 53 192
rect 51 191 52 192
rect 50 191 51 192
rect 49 191 50 192
rect 48 191 49 192
rect 47 191 48 192
rect 46 191 47 192
rect 45 191 46 192
rect 44 191 45 192
rect 43 191 44 192
rect 42 191 43 192
rect 41 191 42 192
rect 40 191 41 192
rect 39 191 40 192
rect 38 191 39 192
rect 37 191 38 192
rect 36 191 37 192
rect 35 191 36 192
rect 34 191 35 192
rect 33 191 34 192
rect 32 191 33 192
rect 31 191 32 192
rect 30 191 31 192
rect 29 191 30 192
rect 28 191 29 192
rect 27 191 28 192
rect 26 191 27 192
rect 25 191 26 192
rect 24 191 25 192
rect 23 191 24 192
rect 22 191 23 192
rect 21 191 22 192
rect 20 191 21 192
rect 19 191 20 192
rect 18 191 19 192
rect 146 192 147 193
rect 145 192 146 193
rect 144 192 145 193
rect 143 192 144 193
rect 142 192 143 193
rect 141 192 142 193
rect 140 192 141 193
rect 139 192 140 193
rect 138 192 139 193
rect 137 192 138 193
rect 136 192 137 193
rect 135 192 136 193
rect 134 192 135 193
rect 133 192 134 193
rect 132 192 133 193
rect 131 192 132 193
rect 130 192 131 193
rect 129 192 130 193
rect 128 192 129 193
rect 79 192 80 193
rect 78 192 79 193
rect 77 192 78 193
rect 76 192 77 193
rect 75 192 76 193
rect 74 192 75 193
rect 73 192 74 193
rect 72 192 73 193
rect 71 192 72 193
rect 70 192 71 193
rect 69 192 70 193
rect 68 192 69 193
rect 67 192 68 193
rect 66 192 67 193
rect 65 192 66 193
rect 64 192 65 193
rect 63 192 64 193
rect 62 192 63 193
rect 61 192 62 193
rect 60 192 61 193
rect 59 192 60 193
rect 58 192 59 193
rect 57 192 58 193
rect 56 192 57 193
rect 55 192 56 193
rect 54 192 55 193
rect 53 192 54 193
rect 52 192 53 193
rect 51 192 52 193
rect 50 192 51 193
rect 49 192 50 193
rect 48 192 49 193
rect 47 192 48 193
rect 46 192 47 193
rect 45 192 46 193
rect 44 192 45 193
rect 43 192 44 193
rect 42 192 43 193
rect 41 192 42 193
rect 40 192 41 193
rect 39 192 40 193
rect 38 192 39 193
rect 37 192 38 193
rect 36 192 37 193
rect 35 192 36 193
rect 34 192 35 193
rect 33 192 34 193
rect 32 192 33 193
rect 31 192 32 193
rect 30 192 31 193
rect 29 192 30 193
rect 28 192 29 193
rect 27 192 28 193
rect 26 192 27 193
rect 25 192 26 193
rect 24 192 25 193
rect 23 192 24 193
rect 22 192 23 193
rect 21 192 22 193
rect 20 192 21 193
rect 19 192 20 193
rect 18 192 19 193
rect 146 193 147 194
rect 145 193 146 194
rect 144 193 145 194
rect 143 193 144 194
rect 142 193 143 194
rect 141 193 142 194
rect 140 193 141 194
rect 139 193 140 194
rect 138 193 139 194
rect 137 193 138 194
rect 136 193 137 194
rect 135 193 136 194
rect 134 193 135 194
rect 133 193 134 194
rect 132 193 133 194
rect 131 193 132 194
rect 130 193 131 194
rect 129 193 130 194
rect 78 193 79 194
rect 77 193 78 194
rect 76 193 77 194
rect 75 193 76 194
rect 74 193 75 194
rect 73 193 74 194
rect 72 193 73 194
rect 71 193 72 194
rect 70 193 71 194
rect 69 193 70 194
rect 68 193 69 194
rect 67 193 68 194
rect 66 193 67 194
rect 65 193 66 194
rect 64 193 65 194
rect 63 193 64 194
rect 62 193 63 194
rect 61 193 62 194
rect 60 193 61 194
rect 59 193 60 194
rect 58 193 59 194
rect 57 193 58 194
rect 56 193 57 194
rect 55 193 56 194
rect 54 193 55 194
rect 53 193 54 194
rect 52 193 53 194
rect 51 193 52 194
rect 50 193 51 194
rect 49 193 50 194
rect 48 193 49 194
rect 47 193 48 194
rect 46 193 47 194
rect 45 193 46 194
rect 44 193 45 194
rect 43 193 44 194
rect 42 193 43 194
rect 41 193 42 194
rect 40 193 41 194
rect 39 193 40 194
rect 38 193 39 194
rect 37 193 38 194
rect 36 193 37 194
rect 35 193 36 194
rect 34 193 35 194
rect 33 193 34 194
rect 32 193 33 194
rect 31 193 32 194
rect 30 193 31 194
rect 29 193 30 194
rect 28 193 29 194
rect 27 193 28 194
rect 26 193 27 194
rect 25 193 26 194
rect 24 193 25 194
rect 23 193 24 194
rect 22 193 23 194
rect 21 193 22 194
rect 20 193 21 194
rect 19 193 20 194
rect 18 193 19 194
rect 146 194 147 195
rect 145 194 146 195
rect 144 194 145 195
rect 143 194 144 195
rect 142 194 143 195
rect 141 194 142 195
rect 140 194 141 195
rect 139 194 140 195
rect 138 194 139 195
rect 137 194 138 195
rect 136 194 137 195
rect 135 194 136 195
rect 134 194 135 195
rect 133 194 134 195
rect 132 194 133 195
rect 131 194 132 195
rect 130 194 131 195
rect 77 194 78 195
rect 76 194 77 195
rect 75 194 76 195
rect 74 194 75 195
rect 73 194 74 195
rect 72 194 73 195
rect 71 194 72 195
rect 70 194 71 195
rect 69 194 70 195
rect 68 194 69 195
rect 67 194 68 195
rect 66 194 67 195
rect 65 194 66 195
rect 64 194 65 195
rect 63 194 64 195
rect 62 194 63 195
rect 61 194 62 195
rect 60 194 61 195
rect 59 194 60 195
rect 58 194 59 195
rect 57 194 58 195
rect 56 194 57 195
rect 55 194 56 195
rect 54 194 55 195
rect 53 194 54 195
rect 52 194 53 195
rect 51 194 52 195
rect 50 194 51 195
rect 49 194 50 195
rect 48 194 49 195
rect 47 194 48 195
rect 46 194 47 195
rect 45 194 46 195
rect 44 194 45 195
rect 43 194 44 195
rect 42 194 43 195
rect 41 194 42 195
rect 40 194 41 195
rect 39 194 40 195
rect 38 194 39 195
rect 37 194 38 195
rect 36 194 37 195
rect 35 194 36 195
rect 34 194 35 195
rect 33 194 34 195
rect 32 194 33 195
rect 31 194 32 195
rect 30 194 31 195
rect 29 194 30 195
rect 28 194 29 195
rect 27 194 28 195
rect 26 194 27 195
rect 25 194 26 195
rect 24 194 25 195
rect 23 194 24 195
rect 22 194 23 195
rect 21 194 22 195
rect 20 194 21 195
rect 19 194 20 195
rect 18 194 19 195
rect 146 195 147 196
rect 145 195 146 196
rect 144 195 145 196
rect 143 195 144 196
rect 142 195 143 196
rect 141 195 142 196
rect 140 195 141 196
rect 139 195 140 196
rect 138 195 139 196
rect 137 195 138 196
rect 136 195 137 196
rect 135 195 136 196
rect 134 195 135 196
rect 133 195 134 196
rect 132 195 133 196
rect 131 195 132 196
rect 76 195 77 196
rect 75 195 76 196
rect 74 195 75 196
rect 73 195 74 196
rect 72 195 73 196
rect 71 195 72 196
rect 70 195 71 196
rect 69 195 70 196
rect 68 195 69 196
rect 67 195 68 196
rect 66 195 67 196
rect 65 195 66 196
rect 64 195 65 196
rect 63 195 64 196
rect 62 195 63 196
rect 61 195 62 196
rect 60 195 61 196
rect 59 195 60 196
rect 58 195 59 196
rect 57 195 58 196
rect 56 195 57 196
rect 55 195 56 196
rect 54 195 55 196
rect 53 195 54 196
rect 52 195 53 196
rect 51 195 52 196
rect 50 195 51 196
rect 49 195 50 196
rect 48 195 49 196
rect 47 195 48 196
rect 46 195 47 196
rect 45 195 46 196
rect 44 195 45 196
rect 43 195 44 196
rect 42 195 43 196
rect 41 195 42 196
rect 40 195 41 196
rect 39 195 40 196
rect 38 195 39 196
rect 37 195 38 196
rect 36 195 37 196
rect 35 195 36 196
rect 34 195 35 196
rect 33 195 34 196
rect 32 195 33 196
rect 31 195 32 196
rect 30 195 31 196
rect 29 195 30 196
rect 28 195 29 196
rect 27 195 28 196
rect 26 195 27 196
rect 25 195 26 196
rect 24 195 25 196
rect 23 195 24 196
rect 22 195 23 196
rect 21 195 22 196
rect 20 195 21 196
rect 19 195 20 196
rect 18 195 19 196
rect 74 196 75 197
rect 73 196 74 197
rect 72 196 73 197
rect 71 196 72 197
rect 70 196 71 197
rect 69 196 70 197
rect 68 196 69 197
rect 67 196 68 197
rect 66 196 67 197
rect 65 196 66 197
rect 64 196 65 197
rect 63 196 64 197
rect 62 196 63 197
rect 61 196 62 197
rect 60 196 61 197
rect 59 196 60 197
rect 58 196 59 197
rect 57 196 58 197
rect 56 196 57 197
rect 55 196 56 197
rect 54 196 55 197
rect 53 196 54 197
rect 52 196 53 197
rect 51 196 52 197
rect 50 196 51 197
rect 49 196 50 197
rect 48 196 49 197
rect 47 196 48 197
rect 46 196 47 197
rect 45 196 46 197
rect 44 196 45 197
rect 43 196 44 197
rect 42 196 43 197
rect 41 196 42 197
rect 40 196 41 197
rect 39 196 40 197
rect 38 196 39 197
rect 37 196 38 197
rect 36 196 37 197
rect 35 196 36 197
rect 34 196 35 197
rect 33 196 34 197
rect 32 196 33 197
rect 31 196 32 197
rect 30 196 31 197
rect 29 196 30 197
rect 28 196 29 197
rect 27 196 28 197
rect 26 196 27 197
rect 25 196 26 197
rect 24 196 25 197
rect 23 196 24 197
rect 22 196 23 197
rect 21 196 22 197
rect 20 196 21 197
rect 19 196 20 197
rect 18 196 19 197
rect 73 197 74 198
rect 72 197 73 198
rect 71 197 72 198
rect 70 197 71 198
rect 69 197 70 198
rect 68 197 69 198
rect 67 197 68 198
rect 66 197 67 198
rect 65 197 66 198
rect 64 197 65 198
rect 63 197 64 198
rect 62 197 63 198
rect 61 197 62 198
rect 60 197 61 198
rect 59 197 60 198
rect 58 197 59 198
rect 57 197 58 198
rect 56 197 57 198
rect 55 197 56 198
rect 54 197 55 198
rect 53 197 54 198
rect 52 197 53 198
rect 51 197 52 198
rect 50 197 51 198
rect 49 197 50 198
rect 48 197 49 198
rect 47 197 48 198
rect 46 197 47 198
rect 45 197 46 198
rect 44 197 45 198
rect 43 197 44 198
rect 42 197 43 198
rect 41 197 42 198
rect 40 197 41 198
rect 39 197 40 198
rect 38 197 39 198
rect 37 197 38 198
rect 36 197 37 198
rect 35 197 36 198
rect 34 197 35 198
rect 33 197 34 198
rect 32 197 33 198
rect 31 197 32 198
rect 30 197 31 198
rect 29 197 30 198
rect 28 197 29 198
rect 27 197 28 198
rect 26 197 27 198
rect 25 197 26 198
rect 24 197 25 198
rect 23 197 24 198
rect 22 197 23 198
rect 21 197 22 198
rect 20 197 21 198
rect 19 197 20 198
rect 18 197 19 198
rect 71 198 72 199
rect 70 198 71 199
rect 69 198 70 199
rect 68 198 69 199
rect 67 198 68 199
rect 66 198 67 199
rect 65 198 66 199
rect 64 198 65 199
rect 63 198 64 199
rect 62 198 63 199
rect 61 198 62 199
rect 60 198 61 199
rect 59 198 60 199
rect 58 198 59 199
rect 57 198 58 199
rect 56 198 57 199
rect 55 198 56 199
rect 54 198 55 199
rect 53 198 54 199
rect 52 198 53 199
rect 51 198 52 199
rect 50 198 51 199
rect 49 198 50 199
rect 48 198 49 199
rect 47 198 48 199
rect 46 198 47 199
rect 45 198 46 199
rect 44 198 45 199
rect 43 198 44 199
rect 42 198 43 199
rect 41 198 42 199
rect 40 198 41 199
rect 39 198 40 199
rect 38 198 39 199
rect 37 198 38 199
rect 36 198 37 199
rect 35 198 36 199
rect 34 198 35 199
rect 33 198 34 199
rect 32 198 33 199
rect 31 198 32 199
rect 30 198 31 199
rect 29 198 30 199
rect 28 198 29 199
rect 27 198 28 199
rect 26 198 27 199
rect 25 198 26 199
rect 24 198 25 199
rect 23 198 24 199
rect 22 198 23 199
rect 21 198 22 199
rect 20 198 21 199
rect 19 198 20 199
rect 18 198 19 199
rect 68 199 69 200
rect 67 199 68 200
rect 66 199 67 200
rect 65 199 66 200
rect 64 199 65 200
rect 63 199 64 200
rect 62 199 63 200
rect 61 199 62 200
rect 60 199 61 200
rect 59 199 60 200
rect 58 199 59 200
rect 57 199 58 200
rect 56 199 57 200
rect 55 199 56 200
rect 54 199 55 200
rect 53 199 54 200
rect 52 199 53 200
rect 51 199 52 200
rect 50 199 51 200
rect 49 199 50 200
rect 48 199 49 200
rect 47 199 48 200
rect 46 199 47 200
rect 45 199 46 200
rect 44 199 45 200
rect 43 199 44 200
rect 42 199 43 200
rect 41 199 42 200
rect 40 199 41 200
rect 39 199 40 200
rect 38 199 39 200
rect 37 199 38 200
rect 36 199 37 200
rect 35 199 36 200
rect 34 199 35 200
rect 33 199 34 200
rect 32 199 33 200
rect 31 199 32 200
rect 30 199 31 200
rect 29 199 30 200
rect 28 199 29 200
rect 27 199 28 200
rect 26 199 27 200
rect 25 199 26 200
rect 24 199 25 200
rect 23 199 24 200
rect 22 199 23 200
rect 21 199 22 200
rect 20 199 21 200
rect 19 199 20 200
rect 18 199 19 200
rect 144 200 145 201
rect 143 200 144 201
rect 65 200 66 201
rect 64 200 65 201
rect 63 200 64 201
rect 62 200 63 201
rect 61 200 62 201
rect 60 200 61 201
rect 59 200 60 201
rect 58 200 59 201
rect 57 200 58 201
rect 56 200 57 201
rect 55 200 56 201
rect 54 200 55 201
rect 53 200 54 201
rect 52 200 53 201
rect 51 200 52 201
rect 50 200 51 201
rect 49 200 50 201
rect 48 200 49 201
rect 47 200 48 201
rect 46 200 47 201
rect 45 200 46 201
rect 44 200 45 201
rect 43 200 44 201
rect 42 200 43 201
rect 41 200 42 201
rect 40 200 41 201
rect 39 200 40 201
rect 38 200 39 201
rect 37 200 38 201
rect 36 200 37 201
rect 35 200 36 201
rect 34 200 35 201
rect 33 200 34 201
rect 32 200 33 201
rect 31 200 32 201
rect 30 200 31 201
rect 29 200 30 201
rect 28 200 29 201
rect 27 200 28 201
rect 26 200 27 201
rect 25 200 26 201
rect 24 200 25 201
rect 23 200 24 201
rect 22 200 23 201
rect 21 200 22 201
rect 20 200 21 201
rect 19 200 20 201
rect 18 200 19 201
rect 145 201 146 202
rect 144 201 145 202
rect 143 201 144 202
rect 142 201 143 202
rect 57 201 58 202
rect 56 201 57 202
rect 55 201 56 202
rect 54 201 55 202
rect 53 201 54 202
rect 52 201 53 202
rect 51 201 52 202
rect 50 201 51 202
rect 49 201 50 202
rect 48 201 49 202
rect 47 201 48 202
rect 46 201 47 202
rect 45 201 46 202
rect 44 201 45 202
rect 43 201 44 202
rect 42 201 43 202
rect 41 201 42 202
rect 40 201 41 202
rect 39 201 40 202
rect 38 201 39 202
rect 37 201 38 202
rect 36 201 37 202
rect 35 201 36 202
rect 34 201 35 202
rect 33 201 34 202
rect 32 201 33 202
rect 31 201 32 202
rect 30 201 31 202
rect 29 201 30 202
rect 28 201 29 202
rect 27 201 28 202
rect 26 201 27 202
rect 25 201 26 202
rect 24 201 25 202
rect 23 201 24 202
rect 22 201 23 202
rect 21 201 22 202
rect 20 201 21 202
rect 19 201 20 202
rect 18 201 19 202
rect 146 202 147 203
rect 145 202 146 203
rect 144 202 145 203
rect 143 202 144 203
rect 142 202 143 203
rect 141 202 142 203
rect 146 203 147 204
rect 145 203 146 204
rect 144 203 145 204
rect 143 203 144 204
rect 142 203 143 204
rect 141 203 142 204
rect 146 204 147 205
rect 145 204 146 205
rect 144 204 145 205
rect 143 204 144 205
rect 142 204 143 205
rect 141 204 142 205
rect 145 205 146 206
rect 144 205 145 206
rect 143 205 144 206
rect 142 205 143 206
rect 144 206 145 207
rect 143 206 144 207
rect 142 222 143 223
rect 141 222 142 223
rect 140 222 141 223
rect 139 222 140 223
rect 138 222 139 223
rect 137 222 138 223
rect 136 222 137 223
rect 135 222 136 223
rect 134 222 135 223
rect 133 222 134 223
rect 132 222 133 223
rect 145 223 146 224
rect 144 223 145 224
rect 143 223 144 224
rect 142 223 143 224
rect 141 223 142 224
rect 140 223 141 224
rect 139 223 140 224
rect 138 223 139 224
rect 137 223 138 224
rect 136 223 137 224
rect 135 223 136 224
rect 134 223 135 224
rect 133 223 134 224
rect 132 223 133 224
rect 131 223 132 224
rect 130 223 131 224
rect 129 223 130 224
rect 128 223 129 224
rect 147 224 148 225
rect 146 224 147 225
rect 145 224 146 225
rect 144 224 145 225
rect 143 224 144 225
rect 142 224 143 225
rect 141 224 142 225
rect 140 224 141 225
rect 139 224 140 225
rect 138 224 139 225
rect 137 224 138 225
rect 136 224 137 225
rect 135 224 136 225
rect 134 224 135 225
rect 133 224 134 225
rect 132 224 133 225
rect 131 224 132 225
rect 130 224 131 225
rect 129 224 130 225
rect 128 224 129 225
rect 127 224 128 225
rect 126 224 127 225
rect 149 225 150 226
rect 148 225 149 226
rect 147 225 148 226
rect 146 225 147 226
rect 145 225 146 226
rect 144 225 145 226
rect 143 225 144 226
rect 142 225 143 226
rect 141 225 142 226
rect 140 225 141 226
rect 139 225 140 226
rect 138 225 139 226
rect 137 225 138 226
rect 136 225 137 226
rect 135 225 136 226
rect 134 225 135 226
rect 133 225 134 226
rect 132 225 133 226
rect 131 225 132 226
rect 130 225 131 226
rect 129 225 130 226
rect 128 225 129 226
rect 127 225 128 226
rect 126 225 127 226
rect 125 225 126 226
rect 124 225 125 226
rect 151 226 152 227
rect 150 226 151 227
rect 149 226 150 227
rect 148 226 149 227
rect 147 226 148 227
rect 146 226 147 227
rect 145 226 146 227
rect 144 226 145 227
rect 143 226 144 227
rect 142 226 143 227
rect 141 226 142 227
rect 140 226 141 227
rect 139 226 140 227
rect 138 226 139 227
rect 137 226 138 227
rect 136 226 137 227
rect 135 226 136 227
rect 134 226 135 227
rect 133 226 134 227
rect 132 226 133 227
rect 131 226 132 227
rect 130 226 131 227
rect 129 226 130 227
rect 128 226 129 227
rect 127 226 128 227
rect 126 226 127 227
rect 125 226 126 227
rect 124 226 125 227
rect 123 226 124 227
rect 152 227 153 228
rect 151 227 152 228
rect 150 227 151 228
rect 149 227 150 228
rect 148 227 149 228
rect 147 227 148 228
rect 146 227 147 228
rect 145 227 146 228
rect 144 227 145 228
rect 143 227 144 228
rect 130 227 131 228
rect 129 227 130 228
rect 128 227 129 228
rect 127 227 128 228
rect 126 227 127 228
rect 125 227 126 228
rect 124 227 125 228
rect 123 227 124 228
rect 122 227 123 228
rect 121 227 122 228
rect 152 228 153 229
rect 151 228 152 229
rect 150 228 151 229
rect 149 228 150 229
rect 148 228 149 229
rect 147 228 148 229
rect 146 228 147 229
rect 127 228 128 229
rect 126 228 127 229
rect 125 228 126 229
rect 124 228 125 229
rect 123 228 124 229
rect 122 228 123 229
rect 121 228 122 229
rect 152 229 153 230
rect 151 229 152 230
rect 150 229 151 230
rect 149 229 150 230
rect 125 229 126 230
rect 124 229 125 230
rect 123 229 124 230
rect 122 229 123 230
rect 121 229 122 230
rect 152 230 153 231
rect 151 230 152 231
rect 150 230 151 231
rect 123 230 124 231
rect 122 230 123 231
rect 121 230 122 231
rect 152 231 153 232
rect 121 231 122 232
rect 140 234 141 235
rect 139 234 140 235
rect 138 234 139 235
rect 137 234 138 235
rect 136 234 137 235
rect 135 234 136 235
rect 142 235 143 236
rect 141 235 142 236
rect 140 235 141 236
rect 139 235 140 236
rect 138 235 139 236
rect 137 235 138 236
rect 136 235 137 236
rect 135 235 136 236
rect 134 235 135 236
rect 133 235 134 236
rect 132 235 133 236
rect 143 236 144 237
rect 142 236 143 237
rect 141 236 142 237
rect 140 236 141 237
rect 139 236 140 237
rect 138 236 139 237
rect 137 236 138 237
rect 136 236 137 237
rect 135 236 136 237
rect 134 236 135 237
rect 133 236 134 237
rect 132 236 133 237
rect 131 236 132 237
rect 144 237 145 238
rect 143 237 144 238
rect 142 237 143 238
rect 141 237 142 238
rect 140 237 141 238
rect 139 237 140 238
rect 138 237 139 238
rect 137 237 138 238
rect 136 237 137 238
rect 135 237 136 238
rect 134 237 135 238
rect 133 237 134 238
rect 132 237 133 238
rect 131 237 132 238
rect 130 237 131 238
rect 145 238 146 239
rect 144 238 145 239
rect 143 238 144 239
rect 142 238 143 239
rect 141 238 142 239
rect 140 238 141 239
rect 139 238 140 239
rect 138 238 139 239
rect 137 238 138 239
rect 136 238 137 239
rect 135 238 136 239
rect 134 238 135 239
rect 133 238 134 239
rect 132 238 133 239
rect 131 238 132 239
rect 130 238 131 239
rect 145 239 146 240
rect 144 239 145 240
rect 143 239 144 240
rect 142 239 143 240
rect 141 239 142 240
rect 140 239 141 240
rect 139 239 140 240
rect 138 239 139 240
rect 137 239 138 240
rect 136 239 137 240
rect 135 239 136 240
rect 134 239 135 240
rect 133 239 134 240
rect 132 239 133 240
rect 131 239 132 240
rect 130 239 131 240
rect 129 239 130 240
rect 63 239 64 240
rect 62 239 63 240
rect 61 239 62 240
rect 60 239 61 240
rect 59 239 60 240
rect 58 239 59 240
rect 57 239 58 240
rect 56 239 57 240
rect 55 239 56 240
rect 54 239 55 240
rect 53 239 54 240
rect 52 239 53 240
rect 51 239 52 240
rect 50 239 51 240
rect 49 239 50 240
rect 48 239 49 240
rect 47 239 48 240
rect 46 239 47 240
rect 146 240 147 241
rect 145 240 146 241
rect 144 240 145 241
rect 143 240 144 241
rect 142 240 143 241
rect 141 240 142 241
rect 134 240 135 241
rect 133 240 134 241
rect 132 240 133 241
rect 131 240 132 241
rect 130 240 131 241
rect 129 240 130 241
rect 67 240 68 241
rect 66 240 67 241
rect 65 240 66 241
rect 64 240 65 241
rect 63 240 64 241
rect 62 240 63 241
rect 61 240 62 241
rect 60 240 61 241
rect 59 240 60 241
rect 58 240 59 241
rect 57 240 58 241
rect 56 240 57 241
rect 55 240 56 241
rect 54 240 55 241
rect 53 240 54 241
rect 52 240 53 241
rect 51 240 52 241
rect 50 240 51 241
rect 49 240 50 241
rect 48 240 49 241
rect 47 240 48 241
rect 46 240 47 241
rect 45 240 46 241
rect 44 240 45 241
rect 43 240 44 241
rect 42 240 43 241
rect 41 240 42 241
rect 146 241 147 242
rect 145 241 146 242
rect 144 241 145 242
rect 143 241 144 242
rect 142 241 143 242
rect 132 241 133 242
rect 131 241 132 242
rect 130 241 131 242
rect 129 241 130 242
rect 128 241 129 242
rect 70 241 71 242
rect 69 241 70 242
rect 68 241 69 242
rect 67 241 68 242
rect 66 241 67 242
rect 65 241 66 242
rect 64 241 65 242
rect 63 241 64 242
rect 62 241 63 242
rect 61 241 62 242
rect 60 241 61 242
rect 59 241 60 242
rect 58 241 59 242
rect 57 241 58 242
rect 56 241 57 242
rect 55 241 56 242
rect 54 241 55 242
rect 53 241 54 242
rect 52 241 53 242
rect 51 241 52 242
rect 50 241 51 242
rect 49 241 50 242
rect 48 241 49 242
rect 47 241 48 242
rect 46 241 47 242
rect 45 241 46 242
rect 44 241 45 242
rect 43 241 44 242
rect 42 241 43 242
rect 41 241 42 242
rect 40 241 41 242
rect 39 241 40 242
rect 38 241 39 242
rect 146 242 147 243
rect 145 242 146 243
rect 144 242 145 243
rect 143 242 144 243
rect 142 242 143 243
rect 132 242 133 243
rect 131 242 132 243
rect 130 242 131 243
rect 129 242 130 243
rect 128 242 129 243
rect 72 242 73 243
rect 71 242 72 243
rect 70 242 71 243
rect 69 242 70 243
rect 68 242 69 243
rect 67 242 68 243
rect 66 242 67 243
rect 65 242 66 243
rect 64 242 65 243
rect 63 242 64 243
rect 62 242 63 243
rect 61 242 62 243
rect 60 242 61 243
rect 59 242 60 243
rect 58 242 59 243
rect 57 242 58 243
rect 56 242 57 243
rect 55 242 56 243
rect 54 242 55 243
rect 53 242 54 243
rect 52 242 53 243
rect 51 242 52 243
rect 50 242 51 243
rect 49 242 50 243
rect 48 242 49 243
rect 47 242 48 243
rect 46 242 47 243
rect 45 242 46 243
rect 44 242 45 243
rect 43 242 44 243
rect 42 242 43 243
rect 41 242 42 243
rect 40 242 41 243
rect 39 242 40 243
rect 38 242 39 243
rect 37 242 38 243
rect 36 242 37 243
rect 35 242 36 243
rect 146 243 147 244
rect 145 243 146 244
rect 144 243 145 244
rect 143 243 144 244
rect 132 243 133 244
rect 131 243 132 244
rect 130 243 131 244
rect 129 243 130 244
rect 128 243 129 244
rect 74 243 75 244
rect 73 243 74 244
rect 72 243 73 244
rect 71 243 72 244
rect 70 243 71 244
rect 69 243 70 244
rect 68 243 69 244
rect 67 243 68 244
rect 66 243 67 244
rect 65 243 66 244
rect 64 243 65 244
rect 63 243 64 244
rect 62 243 63 244
rect 61 243 62 244
rect 60 243 61 244
rect 59 243 60 244
rect 58 243 59 244
rect 57 243 58 244
rect 56 243 57 244
rect 55 243 56 244
rect 54 243 55 244
rect 53 243 54 244
rect 52 243 53 244
rect 51 243 52 244
rect 50 243 51 244
rect 49 243 50 244
rect 48 243 49 244
rect 47 243 48 244
rect 46 243 47 244
rect 45 243 46 244
rect 44 243 45 244
rect 43 243 44 244
rect 42 243 43 244
rect 41 243 42 244
rect 40 243 41 244
rect 39 243 40 244
rect 38 243 39 244
rect 37 243 38 244
rect 36 243 37 244
rect 35 243 36 244
rect 34 243 35 244
rect 33 243 34 244
rect 146 244 147 245
rect 145 244 146 245
rect 144 244 145 245
rect 143 244 144 245
rect 131 244 132 245
rect 130 244 131 245
rect 129 244 130 245
rect 128 244 129 245
rect 76 244 77 245
rect 75 244 76 245
rect 74 244 75 245
rect 73 244 74 245
rect 72 244 73 245
rect 71 244 72 245
rect 70 244 71 245
rect 69 244 70 245
rect 68 244 69 245
rect 67 244 68 245
rect 66 244 67 245
rect 65 244 66 245
rect 64 244 65 245
rect 63 244 64 245
rect 62 244 63 245
rect 61 244 62 245
rect 60 244 61 245
rect 59 244 60 245
rect 58 244 59 245
rect 57 244 58 245
rect 56 244 57 245
rect 55 244 56 245
rect 54 244 55 245
rect 53 244 54 245
rect 52 244 53 245
rect 51 244 52 245
rect 50 244 51 245
rect 49 244 50 245
rect 48 244 49 245
rect 47 244 48 245
rect 46 244 47 245
rect 45 244 46 245
rect 44 244 45 245
rect 43 244 44 245
rect 42 244 43 245
rect 41 244 42 245
rect 40 244 41 245
rect 39 244 40 245
rect 38 244 39 245
rect 37 244 38 245
rect 36 244 37 245
rect 35 244 36 245
rect 34 244 35 245
rect 33 244 34 245
rect 32 244 33 245
rect 146 245 147 246
rect 145 245 146 246
rect 144 245 145 246
rect 143 245 144 246
rect 131 245 132 246
rect 130 245 131 246
rect 129 245 130 246
rect 128 245 129 246
rect 77 245 78 246
rect 76 245 77 246
rect 75 245 76 246
rect 74 245 75 246
rect 73 245 74 246
rect 72 245 73 246
rect 71 245 72 246
rect 70 245 71 246
rect 69 245 70 246
rect 68 245 69 246
rect 67 245 68 246
rect 66 245 67 246
rect 65 245 66 246
rect 64 245 65 246
rect 63 245 64 246
rect 62 245 63 246
rect 61 245 62 246
rect 60 245 61 246
rect 59 245 60 246
rect 58 245 59 246
rect 57 245 58 246
rect 56 245 57 246
rect 55 245 56 246
rect 54 245 55 246
rect 53 245 54 246
rect 52 245 53 246
rect 51 245 52 246
rect 50 245 51 246
rect 49 245 50 246
rect 48 245 49 246
rect 47 245 48 246
rect 46 245 47 246
rect 45 245 46 246
rect 44 245 45 246
rect 43 245 44 246
rect 42 245 43 246
rect 41 245 42 246
rect 40 245 41 246
rect 39 245 40 246
rect 38 245 39 246
rect 37 245 38 246
rect 36 245 37 246
rect 35 245 36 246
rect 34 245 35 246
rect 33 245 34 246
rect 32 245 33 246
rect 31 245 32 246
rect 30 245 31 246
rect 146 246 147 247
rect 145 246 146 247
rect 144 246 145 247
rect 143 246 144 247
rect 142 246 143 247
rect 132 246 133 247
rect 131 246 132 247
rect 130 246 131 247
rect 129 246 130 247
rect 128 246 129 247
rect 78 246 79 247
rect 77 246 78 247
rect 76 246 77 247
rect 75 246 76 247
rect 74 246 75 247
rect 73 246 74 247
rect 72 246 73 247
rect 71 246 72 247
rect 70 246 71 247
rect 69 246 70 247
rect 68 246 69 247
rect 67 246 68 247
rect 66 246 67 247
rect 65 246 66 247
rect 64 246 65 247
rect 63 246 64 247
rect 62 246 63 247
rect 61 246 62 247
rect 60 246 61 247
rect 59 246 60 247
rect 58 246 59 247
rect 57 246 58 247
rect 56 246 57 247
rect 55 246 56 247
rect 54 246 55 247
rect 53 246 54 247
rect 52 246 53 247
rect 51 246 52 247
rect 50 246 51 247
rect 49 246 50 247
rect 48 246 49 247
rect 47 246 48 247
rect 46 246 47 247
rect 45 246 46 247
rect 44 246 45 247
rect 43 246 44 247
rect 42 246 43 247
rect 41 246 42 247
rect 40 246 41 247
rect 39 246 40 247
rect 38 246 39 247
rect 37 246 38 247
rect 36 246 37 247
rect 35 246 36 247
rect 34 246 35 247
rect 33 246 34 247
rect 32 246 33 247
rect 31 246 32 247
rect 30 246 31 247
rect 29 246 30 247
rect 146 247 147 248
rect 145 247 146 248
rect 144 247 145 248
rect 143 247 144 248
rect 142 247 143 248
rect 132 247 133 248
rect 131 247 132 248
rect 130 247 131 248
rect 129 247 130 248
rect 128 247 129 248
rect 79 247 80 248
rect 78 247 79 248
rect 77 247 78 248
rect 76 247 77 248
rect 75 247 76 248
rect 74 247 75 248
rect 73 247 74 248
rect 72 247 73 248
rect 71 247 72 248
rect 70 247 71 248
rect 69 247 70 248
rect 68 247 69 248
rect 67 247 68 248
rect 66 247 67 248
rect 65 247 66 248
rect 64 247 65 248
rect 63 247 64 248
rect 62 247 63 248
rect 61 247 62 248
rect 60 247 61 248
rect 59 247 60 248
rect 58 247 59 248
rect 57 247 58 248
rect 56 247 57 248
rect 55 247 56 248
rect 54 247 55 248
rect 53 247 54 248
rect 52 247 53 248
rect 51 247 52 248
rect 50 247 51 248
rect 49 247 50 248
rect 48 247 49 248
rect 47 247 48 248
rect 46 247 47 248
rect 45 247 46 248
rect 44 247 45 248
rect 43 247 44 248
rect 42 247 43 248
rect 41 247 42 248
rect 40 247 41 248
rect 39 247 40 248
rect 38 247 39 248
rect 37 247 38 248
rect 36 247 37 248
rect 35 247 36 248
rect 34 247 35 248
rect 33 247 34 248
rect 32 247 33 248
rect 31 247 32 248
rect 30 247 31 248
rect 29 247 30 248
rect 28 247 29 248
rect 27 247 28 248
rect 145 248 146 249
rect 144 248 145 249
rect 143 248 144 249
rect 142 248 143 249
rect 132 248 133 249
rect 131 248 132 249
rect 130 248 131 249
rect 129 248 130 249
rect 80 248 81 249
rect 79 248 80 249
rect 78 248 79 249
rect 77 248 78 249
rect 76 248 77 249
rect 75 248 76 249
rect 74 248 75 249
rect 73 248 74 249
rect 72 248 73 249
rect 71 248 72 249
rect 70 248 71 249
rect 69 248 70 249
rect 68 248 69 249
rect 67 248 68 249
rect 66 248 67 249
rect 65 248 66 249
rect 64 248 65 249
rect 63 248 64 249
rect 62 248 63 249
rect 61 248 62 249
rect 60 248 61 249
rect 59 248 60 249
rect 58 248 59 249
rect 57 248 58 249
rect 56 248 57 249
rect 55 248 56 249
rect 54 248 55 249
rect 53 248 54 249
rect 52 248 53 249
rect 51 248 52 249
rect 50 248 51 249
rect 49 248 50 249
rect 48 248 49 249
rect 47 248 48 249
rect 46 248 47 249
rect 45 248 46 249
rect 44 248 45 249
rect 43 248 44 249
rect 42 248 43 249
rect 41 248 42 249
rect 40 248 41 249
rect 39 248 40 249
rect 38 248 39 249
rect 37 248 38 249
rect 36 248 37 249
rect 35 248 36 249
rect 34 248 35 249
rect 33 248 34 249
rect 32 248 33 249
rect 31 248 32 249
rect 30 248 31 249
rect 29 248 30 249
rect 28 248 29 249
rect 27 248 28 249
rect 26 248 27 249
rect 81 249 82 250
rect 80 249 81 250
rect 79 249 80 250
rect 78 249 79 250
rect 77 249 78 250
rect 76 249 77 250
rect 75 249 76 250
rect 74 249 75 250
rect 73 249 74 250
rect 72 249 73 250
rect 71 249 72 250
rect 70 249 71 250
rect 69 249 70 250
rect 68 249 69 250
rect 67 249 68 250
rect 66 249 67 250
rect 65 249 66 250
rect 64 249 65 250
rect 63 249 64 250
rect 62 249 63 250
rect 61 249 62 250
rect 60 249 61 250
rect 59 249 60 250
rect 58 249 59 250
rect 57 249 58 250
rect 56 249 57 250
rect 55 249 56 250
rect 54 249 55 250
rect 53 249 54 250
rect 52 249 53 250
rect 51 249 52 250
rect 50 249 51 250
rect 49 249 50 250
rect 48 249 49 250
rect 47 249 48 250
rect 46 249 47 250
rect 45 249 46 250
rect 44 249 45 250
rect 43 249 44 250
rect 42 249 43 250
rect 41 249 42 250
rect 40 249 41 250
rect 39 249 40 250
rect 38 249 39 250
rect 37 249 38 250
rect 36 249 37 250
rect 35 249 36 250
rect 34 249 35 250
rect 33 249 34 250
rect 32 249 33 250
rect 31 249 32 250
rect 30 249 31 250
rect 29 249 30 250
rect 28 249 29 250
rect 27 249 28 250
rect 26 249 27 250
rect 25 249 26 250
rect 81 250 82 251
rect 80 250 81 251
rect 79 250 80 251
rect 78 250 79 251
rect 77 250 78 251
rect 76 250 77 251
rect 75 250 76 251
rect 74 250 75 251
rect 73 250 74 251
rect 72 250 73 251
rect 71 250 72 251
rect 70 250 71 251
rect 69 250 70 251
rect 68 250 69 251
rect 67 250 68 251
rect 66 250 67 251
rect 65 250 66 251
rect 64 250 65 251
rect 63 250 64 251
rect 62 250 63 251
rect 61 250 62 251
rect 60 250 61 251
rect 59 250 60 251
rect 58 250 59 251
rect 57 250 58 251
rect 56 250 57 251
rect 55 250 56 251
rect 54 250 55 251
rect 53 250 54 251
rect 52 250 53 251
rect 51 250 52 251
rect 50 250 51 251
rect 49 250 50 251
rect 48 250 49 251
rect 47 250 48 251
rect 46 250 47 251
rect 45 250 46 251
rect 44 250 45 251
rect 43 250 44 251
rect 42 250 43 251
rect 41 250 42 251
rect 40 250 41 251
rect 39 250 40 251
rect 38 250 39 251
rect 37 250 38 251
rect 36 250 37 251
rect 35 250 36 251
rect 34 250 35 251
rect 33 250 34 251
rect 32 250 33 251
rect 31 250 32 251
rect 30 250 31 251
rect 29 250 30 251
rect 28 250 29 251
rect 27 250 28 251
rect 26 250 27 251
rect 25 250 26 251
rect 24 250 25 251
rect 152 251 153 252
rect 121 251 122 252
rect 82 251 83 252
rect 81 251 82 252
rect 80 251 81 252
rect 79 251 80 252
rect 78 251 79 252
rect 77 251 78 252
rect 76 251 77 252
rect 75 251 76 252
rect 74 251 75 252
rect 73 251 74 252
rect 72 251 73 252
rect 71 251 72 252
rect 70 251 71 252
rect 69 251 70 252
rect 68 251 69 252
rect 67 251 68 252
rect 66 251 67 252
rect 65 251 66 252
rect 64 251 65 252
rect 63 251 64 252
rect 62 251 63 252
rect 61 251 62 252
rect 60 251 61 252
rect 59 251 60 252
rect 58 251 59 252
rect 57 251 58 252
rect 56 251 57 252
rect 55 251 56 252
rect 54 251 55 252
rect 53 251 54 252
rect 52 251 53 252
rect 51 251 52 252
rect 50 251 51 252
rect 49 251 50 252
rect 48 251 49 252
rect 47 251 48 252
rect 46 251 47 252
rect 45 251 46 252
rect 44 251 45 252
rect 43 251 44 252
rect 42 251 43 252
rect 41 251 42 252
rect 40 251 41 252
rect 39 251 40 252
rect 38 251 39 252
rect 37 251 38 252
rect 36 251 37 252
rect 35 251 36 252
rect 34 251 35 252
rect 33 251 34 252
rect 32 251 33 252
rect 31 251 32 252
rect 30 251 31 252
rect 29 251 30 252
rect 28 251 29 252
rect 27 251 28 252
rect 26 251 27 252
rect 25 251 26 252
rect 24 251 25 252
rect 23 251 24 252
rect 152 252 153 253
rect 151 252 152 253
rect 122 252 123 253
rect 121 252 122 253
rect 82 252 83 253
rect 81 252 82 253
rect 80 252 81 253
rect 79 252 80 253
rect 78 252 79 253
rect 77 252 78 253
rect 76 252 77 253
rect 75 252 76 253
rect 74 252 75 253
rect 73 252 74 253
rect 72 252 73 253
rect 71 252 72 253
rect 70 252 71 253
rect 69 252 70 253
rect 68 252 69 253
rect 67 252 68 253
rect 66 252 67 253
rect 65 252 66 253
rect 64 252 65 253
rect 63 252 64 253
rect 62 252 63 253
rect 61 252 62 253
rect 60 252 61 253
rect 59 252 60 253
rect 58 252 59 253
rect 57 252 58 253
rect 56 252 57 253
rect 55 252 56 253
rect 54 252 55 253
rect 53 252 54 253
rect 52 252 53 253
rect 51 252 52 253
rect 50 252 51 253
rect 49 252 50 253
rect 48 252 49 253
rect 47 252 48 253
rect 46 252 47 253
rect 45 252 46 253
rect 44 252 45 253
rect 43 252 44 253
rect 42 252 43 253
rect 41 252 42 253
rect 40 252 41 253
rect 39 252 40 253
rect 38 252 39 253
rect 37 252 38 253
rect 36 252 37 253
rect 35 252 36 253
rect 34 252 35 253
rect 33 252 34 253
rect 32 252 33 253
rect 31 252 32 253
rect 30 252 31 253
rect 29 252 30 253
rect 28 252 29 253
rect 27 252 28 253
rect 26 252 27 253
rect 25 252 26 253
rect 24 252 25 253
rect 23 252 24 253
rect 152 253 153 254
rect 151 253 152 254
rect 150 253 151 254
rect 149 253 150 254
rect 124 253 125 254
rect 123 253 124 254
rect 122 253 123 254
rect 121 253 122 254
rect 83 253 84 254
rect 82 253 83 254
rect 81 253 82 254
rect 80 253 81 254
rect 79 253 80 254
rect 78 253 79 254
rect 77 253 78 254
rect 76 253 77 254
rect 75 253 76 254
rect 74 253 75 254
rect 73 253 74 254
rect 72 253 73 254
rect 71 253 72 254
rect 70 253 71 254
rect 69 253 70 254
rect 68 253 69 254
rect 67 253 68 254
rect 66 253 67 254
rect 65 253 66 254
rect 64 253 65 254
rect 63 253 64 254
rect 62 253 63 254
rect 61 253 62 254
rect 60 253 61 254
rect 59 253 60 254
rect 58 253 59 254
rect 57 253 58 254
rect 56 253 57 254
rect 55 253 56 254
rect 54 253 55 254
rect 53 253 54 254
rect 52 253 53 254
rect 51 253 52 254
rect 50 253 51 254
rect 49 253 50 254
rect 48 253 49 254
rect 47 253 48 254
rect 46 253 47 254
rect 45 253 46 254
rect 44 253 45 254
rect 43 253 44 254
rect 42 253 43 254
rect 41 253 42 254
rect 40 253 41 254
rect 39 253 40 254
rect 38 253 39 254
rect 37 253 38 254
rect 36 253 37 254
rect 35 253 36 254
rect 34 253 35 254
rect 33 253 34 254
rect 32 253 33 254
rect 31 253 32 254
rect 30 253 31 254
rect 29 253 30 254
rect 28 253 29 254
rect 27 253 28 254
rect 26 253 27 254
rect 25 253 26 254
rect 24 253 25 254
rect 23 253 24 254
rect 22 253 23 254
rect 152 254 153 255
rect 151 254 152 255
rect 150 254 151 255
rect 149 254 150 255
rect 148 254 149 255
rect 147 254 148 255
rect 126 254 127 255
rect 125 254 126 255
rect 124 254 125 255
rect 123 254 124 255
rect 122 254 123 255
rect 121 254 122 255
rect 83 254 84 255
rect 82 254 83 255
rect 81 254 82 255
rect 80 254 81 255
rect 79 254 80 255
rect 78 254 79 255
rect 77 254 78 255
rect 76 254 77 255
rect 75 254 76 255
rect 74 254 75 255
rect 73 254 74 255
rect 72 254 73 255
rect 71 254 72 255
rect 70 254 71 255
rect 69 254 70 255
rect 68 254 69 255
rect 67 254 68 255
rect 66 254 67 255
rect 65 254 66 255
rect 64 254 65 255
rect 63 254 64 255
rect 62 254 63 255
rect 61 254 62 255
rect 60 254 61 255
rect 59 254 60 255
rect 58 254 59 255
rect 57 254 58 255
rect 56 254 57 255
rect 55 254 56 255
rect 54 254 55 255
rect 53 254 54 255
rect 52 254 53 255
rect 51 254 52 255
rect 50 254 51 255
rect 49 254 50 255
rect 48 254 49 255
rect 47 254 48 255
rect 46 254 47 255
rect 45 254 46 255
rect 44 254 45 255
rect 43 254 44 255
rect 42 254 43 255
rect 41 254 42 255
rect 40 254 41 255
rect 39 254 40 255
rect 38 254 39 255
rect 37 254 38 255
rect 36 254 37 255
rect 35 254 36 255
rect 34 254 35 255
rect 33 254 34 255
rect 32 254 33 255
rect 31 254 32 255
rect 30 254 31 255
rect 29 254 30 255
rect 28 254 29 255
rect 27 254 28 255
rect 26 254 27 255
rect 25 254 26 255
rect 24 254 25 255
rect 23 254 24 255
rect 22 254 23 255
rect 21 254 22 255
rect 152 255 153 256
rect 151 255 152 256
rect 150 255 151 256
rect 149 255 150 256
rect 148 255 149 256
rect 147 255 148 256
rect 146 255 147 256
rect 145 255 146 256
rect 128 255 129 256
rect 127 255 128 256
rect 126 255 127 256
rect 125 255 126 256
rect 124 255 125 256
rect 123 255 124 256
rect 122 255 123 256
rect 121 255 122 256
rect 84 255 85 256
rect 83 255 84 256
rect 82 255 83 256
rect 81 255 82 256
rect 80 255 81 256
rect 79 255 80 256
rect 78 255 79 256
rect 77 255 78 256
rect 76 255 77 256
rect 75 255 76 256
rect 74 255 75 256
rect 73 255 74 256
rect 72 255 73 256
rect 71 255 72 256
rect 70 255 71 256
rect 69 255 70 256
rect 68 255 69 256
rect 67 255 68 256
rect 66 255 67 256
rect 65 255 66 256
rect 64 255 65 256
rect 63 255 64 256
rect 62 255 63 256
rect 61 255 62 256
rect 60 255 61 256
rect 59 255 60 256
rect 58 255 59 256
rect 57 255 58 256
rect 56 255 57 256
rect 55 255 56 256
rect 54 255 55 256
rect 53 255 54 256
rect 52 255 53 256
rect 51 255 52 256
rect 50 255 51 256
rect 49 255 50 256
rect 48 255 49 256
rect 47 255 48 256
rect 46 255 47 256
rect 45 255 46 256
rect 44 255 45 256
rect 43 255 44 256
rect 42 255 43 256
rect 41 255 42 256
rect 40 255 41 256
rect 39 255 40 256
rect 38 255 39 256
rect 37 255 38 256
rect 36 255 37 256
rect 35 255 36 256
rect 34 255 35 256
rect 33 255 34 256
rect 32 255 33 256
rect 31 255 32 256
rect 30 255 31 256
rect 29 255 30 256
rect 28 255 29 256
rect 27 255 28 256
rect 26 255 27 256
rect 25 255 26 256
rect 24 255 25 256
rect 23 255 24 256
rect 22 255 23 256
rect 21 255 22 256
rect 151 256 152 257
rect 150 256 151 257
rect 149 256 150 257
rect 148 256 149 257
rect 147 256 148 257
rect 146 256 147 257
rect 145 256 146 257
rect 144 256 145 257
rect 143 256 144 257
rect 142 256 143 257
rect 141 256 142 257
rect 140 256 141 257
rect 133 256 134 257
rect 132 256 133 257
rect 131 256 132 257
rect 130 256 131 257
rect 129 256 130 257
rect 128 256 129 257
rect 127 256 128 257
rect 126 256 127 257
rect 125 256 126 257
rect 124 256 125 257
rect 123 256 124 257
rect 122 256 123 257
rect 84 256 85 257
rect 83 256 84 257
rect 82 256 83 257
rect 81 256 82 257
rect 80 256 81 257
rect 79 256 80 257
rect 78 256 79 257
rect 77 256 78 257
rect 76 256 77 257
rect 75 256 76 257
rect 74 256 75 257
rect 73 256 74 257
rect 72 256 73 257
rect 71 256 72 257
rect 70 256 71 257
rect 69 256 70 257
rect 68 256 69 257
rect 67 256 68 257
rect 66 256 67 257
rect 65 256 66 257
rect 64 256 65 257
rect 63 256 64 257
rect 62 256 63 257
rect 61 256 62 257
rect 60 256 61 257
rect 59 256 60 257
rect 58 256 59 257
rect 57 256 58 257
rect 56 256 57 257
rect 55 256 56 257
rect 54 256 55 257
rect 53 256 54 257
rect 52 256 53 257
rect 51 256 52 257
rect 50 256 51 257
rect 49 256 50 257
rect 48 256 49 257
rect 47 256 48 257
rect 46 256 47 257
rect 45 256 46 257
rect 44 256 45 257
rect 43 256 44 257
rect 42 256 43 257
rect 41 256 42 257
rect 40 256 41 257
rect 39 256 40 257
rect 38 256 39 257
rect 37 256 38 257
rect 36 256 37 257
rect 35 256 36 257
rect 34 256 35 257
rect 33 256 34 257
rect 32 256 33 257
rect 31 256 32 257
rect 30 256 31 257
rect 29 256 30 257
rect 28 256 29 257
rect 27 256 28 257
rect 26 256 27 257
rect 25 256 26 257
rect 24 256 25 257
rect 23 256 24 257
rect 22 256 23 257
rect 21 256 22 257
rect 20 256 21 257
rect 150 257 151 258
rect 149 257 150 258
rect 148 257 149 258
rect 147 257 148 258
rect 146 257 147 258
rect 145 257 146 258
rect 144 257 145 258
rect 143 257 144 258
rect 142 257 143 258
rect 141 257 142 258
rect 140 257 141 258
rect 139 257 140 258
rect 138 257 139 258
rect 137 257 138 258
rect 136 257 137 258
rect 135 257 136 258
rect 134 257 135 258
rect 133 257 134 258
rect 132 257 133 258
rect 131 257 132 258
rect 130 257 131 258
rect 129 257 130 258
rect 128 257 129 258
rect 127 257 128 258
rect 126 257 127 258
rect 125 257 126 258
rect 124 257 125 258
rect 123 257 124 258
rect 84 257 85 258
rect 83 257 84 258
rect 82 257 83 258
rect 81 257 82 258
rect 80 257 81 258
rect 79 257 80 258
rect 78 257 79 258
rect 77 257 78 258
rect 76 257 77 258
rect 75 257 76 258
rect 74 257 75 258
rect 73 257 74 258
rect 72 257 73 258
rect 71 257 72 258
rect 70 257 71 258
rect 69 257 70 258
rect 68 257 69 258
rect 67 257 68 258
rect 66 257 67 258
rect 65 257 66 258
rect 64 257 65 258
rect 63 257 64 258
rect 62 257 63 258
rect 61 257 62 258
rect 60 257 61 258
rect 59 257 60 258
rect 58 257 59 258
rect 57 257 58 258
rect 56 257 57 258
rect 55 257 56 258
rect 54 257 55 258
rect 53 257 54 258
rect 52 257 53 258
rect 51 257 52 258
rect 50 257 51 258
rect 49 257 50 258
rect 48 257 49 258
rect 47 257 48 258
rect 46 257 47 258
rect 45 257 46 258
rect 44 257 45 258
rect 43 257 44 258
rect 42 257 43 258
rect 41 257 42 258
rect 40 257 41 258
rect 39 257 40 258
rect 38 257 39 258
rect 37 257 38 258
rect 36 257 37 258
rect 35 257 36 258
rect 34 257 35 258
rect 33 257 34 258
rect 32 257 33 258
rect 31 257 32 258
rect 30 257 31 258
rect 29 257 30 258
rect 28 257 29 258
rect 27 257 28 258
rect 26 257 27 258
rect 25 257 26 258
rect 24 257 25 258
rect 23 257 24 258
rect 22 257 23 258
rect 21 257 22 258
rect 20 257 21 258
rect 148 258 149 259
rect 147 258 148 259
rect 146 258 147 259
rect 145 258 146 259
rect 144 258 145 259
rect 143 258 144 259
rect 142 258 143 259
rect 141 258 142 259
rect 140 258 141 259
rect 139 258 140 259
rect 138 258 139 259
rect 137 258 138 259
rect 136 258 137 259
rect 135 258 136 259
rect 134 258 135 259
rect 133 258 134 259
rect 132 258 133 259
rect 131 258 132 259
rect 130 258 131 259
rect 129 258 130 259
rect 128 258 129 259
rect 127 258 128 259
rect 126 258 127 259
rect 125 258 126 259
rect 84 258 85 259
rect 83 258 84 259
rect 82 258 83 259
rect 81 258 82 259
rect 80 258 81 259
rect 79 258 80 259
rect 78 258 79 259
rect 77 258 78 259
rect 76 258 77 259
rect 75 258 76 259
rect 74 258 75 259
rect 73 258 74 259
rect 72 258 73 259
rect 71 258 72 259
rect 70 258 71 259
rect 69 258 70 259
rect 68 258 69 259
rect 67 258 68 259
rect 66 258 67 259
rect 65 258 66 259
rect 64 258 65 259
rect 61 258 62 259
rect 60 258 61 259
rect 59 258 60 259
rect 58 258 59 259
rect 57 258 58 259
rect 56 258 57 259
rect 55 258 56 259
rect 54 258 55 259
rect 53 258 54 259
rect 52 258 53 259
rect 51 258 52 259
rect 50 258 51 259
rect 49 258 50 259
rect 48 258 49 259
rect 47 258 48 259
rect 42 258 43 259
rect 41 258 42 259
rect 40 258 41 259
rect 39 258 40 259
rect 38 258 39 259
rect 37 258 38 259
rect 36 258 37 259
rect 35 258 36 259
rect 34 258 35 259
rect 33 258 34 259
rect 32 258 33 259
rect 31 258 32 259
rect 30 258 31 259
rect 29 258 30 259
rect 28 258 29 259
rect 27 258 28 259
rect 26 258 27 259
rect 25 258 26 259
rect 24 258 25 259
rect 23 258 24 259
rect 22 258 23 259
rect 21 258 22 259
rect 20 258 21 259
rect 19 258 20 259
rect 146 259 147 260
rect 145 259 146 260
rect 144 259 145 260
rect 143 259 144 260
rect 142 259 143 260
rect 141 259 142 260
rect 140 259 141 260
rect 139 259 140 260
rect 138 259 139 260
rect 137 259 138 260
rect 136 259 137 260
rect 135 259 136 260
rect 134 259 135 260
rect 133 259 134 260
rect 132 259 133 260
rect 131 259 132 260
rect 130 259 131 260
rect 129 259 130 260
rect 128 259 129 260
rect 127 259 128 260
rect 85 259 86 260
rect 84 259 85 260
rect 83 259 84 260
rect 82 259 83 260
rect 81 259 82 260
rect 80 259 81 260
rect 79 259 80 260
rect 78 259 79 260
rect 77 259 78 260
rect 76 259 77 260
rect 75 259 76 260
rect 74 259 75 260
rect 73 259 74 260
rect 72 259 73 260
rect 71 259 72 260
rect 70 259 71 260
rect 69 259 70 260
rect 68 259 69 260
rect 57 259 58 260
rect 56 259 57 260
rect 55 259 56 260
rect 54 259 55 260
rect 53 259 54 260
rect 52 259 53 260
rect 51 259 52 260
rect 50 259 51 260
rect 49 259 50 260
rect 48 259 49 260
rect 47 259 48 260
rect 46 259 47 260
rect 39 259 40 260
rect 38 259 39 260
rect 37 259 38 260
rect 36 259 37 260
rect 35 259 36 260
rect 34 259 35 260
rect 33 259 34 260
rect 32 259 33 260
rect 31 259 32 260
rect 30 259 31 260
rect 29 259 30 260
rect 28 259 29 260
rect 27 259 28 260
rect 26 259 27 260
rect 25 259 26 260
rect 24 259 25 260
rect 23 259 24 260
rect 22 259 23 260
rect 21 259 22 260
rect 20 259 21 260
rect 19 259 20 260
rect 144 260 145 261
rect 143 260 144 261
rect 142 260 143 261
rect 141 260 142 261
rect 140 260 141 261
rect 139 260 140 261
rect 138 260 139 261
rect 137 260 138 261
rect 136 260 137 261
rect 135 260 136 261
rect 134 260 135 261
rect 133 260 134 261
rect 132 260 133 261
rect 131 260 132 261
rect 130 260 131 261
rect 85 260 86 261
rect 84 260 85 261
rect 83 260 84 261
rect 82 260 83 261
rect 81 260 82 261
rect 80 260 81 261
rect 79 260 80 261
rect 78 260 79 261
rect 77 260 78 261
rect 76 260 77 261
rect 75 260 76 261
rect 74 260 75 261
rect 73 260 74 261
rect 72 260 73 261
rect 71 260 72 261
rect 70 260 71 261
rect 69 260 70 261
rect 56 260 57 261
rect 55 260 56 261
rect 54 260 55 261
rect 53 260 54 261
rect 52 260 53 261
rect 51 260 52 261
rect 50 260 51 261
rect 49 260 50 261
rect 48 260 49 261
rect 47 260 48 261
rect 46 260 47 261
rect 45 260 46 261
rect 38 260 39 261
rect 37 260 38 261
rect 36 260 37 261
rect 35 260 36 261
rect 34 260 35 261
rect 33 260 34 261
rect 32 260 33 261
rect 31 260 32 261
rect 30 260 31 261
rect 29 260 30 261
rect 28 260 29 261
rect 27 260 28 261
rect 26 260 27 261
rect 25 260 26 261
rect 24 260 25 261
rect 23 260 24 261
rect 22 260 23 261
rect 21 260 22 261
rect 20 260 21 261
rect 19 260 20 261
rect 85 261 86 262
rect 84 261 85 262
rect 83 261 84 262
rect 82 261 83 262
rect 81 261 82 262
rect 80 261 81 262
rect 79 261 80 262
rect 78 261 79 262
rect 77 261 78 262
rect 76 261 77 262
rect 75 261 76 262
rect 74 261 75 262
rect 73 261 74 262
rect 72 261 73 262
rect 71 261 72 262
rect 70 261 71 262
rect 55 261 56 262
rect 54 261 55 262
rect 53 261 54 262
rect 52 261 53 262
rect 51 261 52 262
rect 50 261 51 262
rect 49 261 50 262
rect 48 261 49 262
rect 47 261 48 262
rect 46 261 47 262
rect 45 261 46 262
rect 44 261 45 262
rect 36 261 37 262
rect 35 261 36 262
rect 34 261 35 262
rect 33 261 34 262
rect 32 261 33 262
rect 31 261 32 262
rect 30 261 31 262
rect 29 261 30 262
rect 28 261 29 262
rect 27 261 28 262
rect 26 261 27 262
rect 25 261 26 262
rect 24 261 25 262
rect 23 261 24 262
rect 22 261 23 262
rect 21 261 22 262
rect 20 261 21 262
rect 19 261 20 262
rect 18 261 19 262
rect 85 262 86 263
rect 84 262 85 263
rect 83 262 84 263
rect 82 262 83 263
rect 81 262 82 263
rect 80 262 81 263
rect 79 262 80 263
rect 78 262 79 263
rect 77 262 78 263
rect 76 262 77 263
rect 75 262 76 263
rect 74 262 75 263
rect 73 262 74 263
rect 72 262 73 263
rect 71 262 72 263
rect 54 262 55 263
rect 53 262 54 263
rect 52 262 53 263
rect 51 262 52 263
rect 50 262 51 263
rect 49 262 50 263
rect 48 262 49 263
rect 47 262 48 263
rect 46 262 47 263
rect 45 262 46 263
rect 44 262 45 263
rect 43 262 44 263
rect 35 262 36 263
rect 34 262 35 263
rect 33 262 34 263
rect 32 262 33 263
rect 31 262 32 263
rect 30 262 31 263
rect 29 262 30 263
rect 28 262 29 263
rect 27 262 28 263
rect 26 262 27 263
rect 25 262 26 263
rect 24 262 25 263
rect 23 262 24 263
rect 22 262 23 263
rect 21 262 22 263
rect 20 262 21 263
rect 19 262 20 263
rect 18 262 19 263
rect 85 263 86 264
rect 84 263 85 264
rect 83 263 84 264
rect 82 263 83 264
rect 81 263 82 264
rect 80 263 81 264
rect 79 263 80 264
rect 78 263 79 264
rect 77 263 78 264
rect 76 263 77 264
rect 75 263 76 264
rect 74 263 75 264
rect 73 263 74 264
rect 72 263 73 264
rect 71 263 72 264
rect 54 263 55 264
rect 53 263 54 264
rect 52 263 53 264
rect 51 263 52 264
rect 50 263 51 264
rect 49 263 50 264
rect 48 263 49 264
rect 47 263 48 264
rect 46 263 47 264
rect 45 263 46 264
rect 44 263 45 264
rect 43 263 44 264
rect 34 263 35 264
rect 33 263 34 264
rect 32 263 33 264
rect 31 263 32 264
rect 30 263 31 264
rect 29 263 30 264
rect 28 263 29 264
rect 27 263 28 264
rect 26 263 27 264
rect 25 263 26 264
rect 24 263 25 264
rect 23 263 24 264
rect 22 263 23 264
rect 21 263 22 264
rect 20 263 21 264
rect 19 263 20 264
rect 18 263 19 264
rect 85 264 86 265
rect 84 264 85 265
rect 83 264 84 265
rect 82 264 83 265
rect 81 264 82 265
rect 80 264 81 265
rect 79 264 80 265
rect 78 264 79 265
rect 77 264 78 265
rect 76 264 77 265
rect 75 264 76 265
rect 74 264 75 265
rect 73 264 74 265
rect 72 264 73 265
rect 71 264 72 265
rect 54 264 55 265
rect 53 264 54 265
rect 52 264 53 265
rect 51 264 52 265
rect 50 264 51 265
rect 49 264 50 265
rect 48 264 49 265
rect 47 264 48 265
rect 46 264 47 265
rect 45 264 46 265
rect 44 264 45 265
rect 43 264 44 265
rect 42 264 43 265
rect 33 264 34 265
rect 32 264 33 265
rect 31 264 32 265
rect 30 264 31 265
rect 29 264 30 265
rect 28 264 29 265
rect 27 264 28 265
rect 26 264 27 265
rect 25 264 26 265
rect 24 264 25 265
rect 23 264 24 265
rect 22 264 23 265
rect 21 264 22 265
rect 20 264 21 265
rect 19 264 20 265
rect 18 264 19 265
rect 85 265 86 266
rect 84 265 85 266
rect 83 265 84 266
rect 82 265 83 266
rect 81 265 82 266
rect 80 265 81 266
rect 79 265 80 266
rect 78 265 79 266
rect 77 265 78 266
rect 76 265 77 266
rect 75 265 76 266
rect 74 265 75 266
rect 73 265 74 266
rect 72 265 73 266
rect 71 265 72 266
rect 54 265 55 266
rect 53 265 54 266
rect 52 265 53 266
rect 51 265 52 266
rect 50 265 51 266
rect 49 265 50 266
rect 48 265 49 266
rect 47 265 48 266
rect 46 265 47 266
rect 45 265 46 266
rect 44 265 45 266
rect 43 265 44 266
rect 42 265 43 266
rect 33 265 34 266
rect 32 265 33 266
rect 31 265 32 266
rect 30 265 31 266
rect 29 265 30 266
rect 28 265 29 266
rect 27 265 28 266
rect 26 265 27 266
rect 25 265 26 266
rect 24 265 25 266
rect 23 265 24 266
rect 22 265 23 266
rect 21 265 22 266
rect 20 265 21 266
rect 19 265 20 266
rect 18 265 19 266
rect 138 266 139 267
rect 137 266 138 267
rect 136 266 137 267
rect 135 266 136 267
rect 134 266 135 267
rect 133 266 134 267
rect 132 266 133 267
rect 131 266 132 267
rect 130 266 131 267
rect 85 266 86 267
rect 84 266 85 267
rect 83 266 84 267
rect 82 266 83 267
rect 81 266 82 267
rect 80 266 81 267
rect 79 266 80 267
rect 78 266 79 267
rect 77 266 78 267
rect 76 266 77 267
rect 75 266 76 267
rect 74 266 75 267
rect 73 266 74 267
rect 72 266 73 267
rect 71 266 72 267
rect 54 266 55 267
rect 53 266 54 267
rect 52 266 53 267
rect 51 266 52 267
rect 50 266 51 267
rect 49 266 50 267
rect 48 266 49 267
rect 47 266 48 267
rect 46 266 47 267
rect 45 266 46 267
rect 44 266 45 267
rect 43 266 44 267
rect 42 266 43 267
rect 32 266 33 267
rect 31 266 32 267
rect 30 266 31 267
rect 29 266 30 267
rect 28 266 29 267
rect 27 266 28 267
rect 26 266 27 267
rect 25 266 26 267
rect 24 266 25 267
rect 23 266 24 267
rect 22 266 23 267
rect 21 266 22 267
rect 20 266 21 267
rect 19 266 20 267
rect 18 266 19 267
rect 17 266 18 267
rect 140 267 141 268
rect 139 267 140 268
rect 138 267 139 268
rect 137 267 138 268
rect 136 267 137 268
rect 135 267 136 268
rect 134 267 135 268
rect 133 267 134 268
rect 132 267 133 268
rect 131 267 132 268
rect 130 267 131 268
rect 129 267 130 268
rect 128 267 129 268
rect 85 267 86 268
rect 84 267 85 268
rect 83 267 84 268
rect 82 267 83 268
rect 81 267 82 268
rect 80 267 81 268
rect 79 267 80 268
rect 78 267 79 268
rect 77 267 78 268
rect 76 267 77 268
rect 75 267 76 268
rect 74 267 75 268
rect 73 267 74 268
rect 72 267 73 268
rect 71 267 72 268
rect 70 267 71 268
rect 55 267 56 268
rect 54 267 55 268
rect 53 267 54 268
rect 52 267 53 268
rect 51 267 52 268
rect 50 267 51 268
rect 49 267 50 268
rect 48 267 49 268
rect 47 267 48 268
rect 46 267 47 268
rect 45 267 46 268
rect 44 267 45 268
rect 43 267 44 268
rect 42 267 43 268
rect 41 267 42 268
rect 32 267 33 268
rect 31 267 32 268
rect 30 267 31 268
rect 29 267 30 268
rect 28 267 29 268
rect 27 267 28 268
rect 26 267 27 268
rect 25 267 26 268
rect 24 267 25 268
rect 23 267 24 268
rect 22 267 23 268
rect 21 267 22 268
rect 20 267 21 268
rect 19 267 20 268
rect 18 267 19 268
rect 17 267 18 268
rect 142 268 143 269
rect 141 268 142 269
rect 140 268 141 269
rect 139 268 140 269
rect 138 268 139 269
rect 137 268 138 269
rect 136 268 137 269
rect 135 268 136 269
rect 134 268 135 269
rect 133 268 134 269
rect 132 268 133 269
rect 131 268 132 269
rect 130 268 131 269
rect 129 268 130 269
rect 128 268 129 269
rect 127 268 128 269
rect 126 268 127 269
rect 85 268 86 269
rect 84 268 85 269
rect 83 268 84 269
rect 82 268 83 269
rect 81 268 82 269
rect 80 268 81 269
rect 79 268 80 269
rect 78 268 79 269
rect 77 268 78 269
rect 76 268 77 269
rect 75 268 76 269
rect 74 268 75 269
rect 73 268 74 269
rect 72 268 73 269
rect 71 268 72 269
rect 70 268 71 269
rect 69 268 70 269
rect 56 268 57 269
rect 55 268 56 269
rect 54 268 55 269
rect 53 268 54 269
rect 52 268 53 269
rect 51 268 52 269
rect 50 268 51 269
rect 49 268 50 269
rect 48 268 49 269
rect 47 268 48 269
rect 46 268 47 269
rect 45 268 46 269
rect 44 268 45 269
rect 43 268 44 269
rect 42 268 43 269
rect 41 268 42 269
rect 32 268 33 269
rect 31 268 32 269
rect 30 268 31 269
rect 29 268 30 269
rect 28 268 29 269
rect 27 268 28 269
rect 26 268 27 269
rect 25 268 26 269
rect 24 268 25 269
rect 23 268 24 269
rect 22 268 23 269
rect 21 268 22 269
rect 20 268 21 269
rect 19 268 20 269
rect 18 268 19 269
rect 17 268 18 269
rect 143 269 144 270
rect 142 269 143 270
rect 141 269 142 270
rect 140 269 141 270
rect 139 269 140 270
rect 138 269 139 270
rect 137 269 138 270
rect 136 269 137 270
rect 135 269 136 270
rect 134 269 135 270
rect 133 269 134 270
rect 132 269 133 270
rect 131 269 132 270
rect 130 269 131 270
rect 129 269 130 270
rect 128 269 129 270
rect 127 269 128 270
rect 126 269 127 270
rect 125 269 126 270
rect 84 269 85 270
rect 83 269 84 270
rect 82 269 83 270
rect 81 269 82 270
rect 80 269 81 270
rect 79 269 80 270
rect 78 269 79 270
rect 77 269 78 270
rect 76 269 77 270
rect 75 269 76 270
rect 74 269 75 270
rect 73 269 74 270
rect 72 269 73 270
rect 71 269 72 270
rect 70 269 71 270
rect 69 269 70 270
rect 68 269 69 270
rect 67 269 68 270
rect 58 269 59 270
rect 57 269 58 270
rect 56 269 57 270
rect 55 269 56 270
rect 54 269 55 270
rect 53 269 54 270
rect 52 269 53 270
rect 51 269 52 270
rect 50 269 51 270
rect 49 269 50 270
rect 48 269 49 270
rect 47 269 48 270
rect 46 269 47 270
rect 45 269 46 270
rect 44 269 45 270
rect 43 269 44 270
rect 42 269 43 270
rect 41 269 42 270
rect 31 269 32 270
rect 30 269 31 270
rect 29 269 30 270
rect 28 269 29 270
rect 27 269 28 270
rect 26 269 27 270
rect 25 269 26 270
rect 24 269 25 270
rect 23 269 24 270
rect 22 269 23 270
rect 21 269 22 270
rect 20 269 21 270
rect 19 269 20 270
rect 18 269 19 270
rect 17 269 18 270
rect 143 270 144 271
rect 142 270 143 271
rect 141 270 142 271
rect 140 270 141 271
rect 139 270 140 271
rect 138 270 139 271
rect 137 270 138 271
rect 136 270 137 271
rect 135 270 136 271
rect 134 270 135 271
rect 133 270 134 271
rect 132 270 133 271
rect 131 270 132 271
rect 130 270 131 271
rect 129 270 130 271
rect 128 270 129 271
rect 127 270 128 271
rect 126 270 127 271
rect 125 270 126 271
rect 124 270 125 271
rect 84 270 85 271
rect 83 270 84 271
rect 82 270 83 271
rect 81 270 82 271
rect 80 270 81 271
rect 79 270 80 271
rect 78 270 79 271
rect 77 270 78 271
rect 76 270 77 271
rect 75 270 76 271
rect 74 270 75 271
rect 73 270 74 271
rect 72 270 73 271
rect 71 270 72 271
rect 70 270 71 271
rect 69 270 70 271
rect 68 270 69 271
rect 67 270 68 271
rect 66 270 67 271
rect 65 270 66 271
rect 64 270 65 271
rect 63 270 64 271
rect 62 270 63 271
rect 61 270 62 271
rect 60 270 61 271
rect 59 270 60 271
rect 58 270 59 271
rect 57 270 58 271
rect 56 270 57 271
rect 55 270 56 271
rect 54 270 55 271
rect 53 270 54 271
rect 52 270 53 271
rect 51 270 52 271
rect 50 270 51 271
rect 49 270 50 271
rect 48 270 49 271
rect 47 270 48 271
rect 46 270 47 271
rect 45 270 46 271
rect 44 270 45 271
rect 43 270 44 271
rect 42 270 43 271
rect 41 270 42 271
rect 31 270 32 271
rect 30 270 31 271
rect 29 270 30 271
rect 28 270 29 271
rect 27 270 28 271
rect 26 270 27 271
rect 25 270 26 271
rect 24 270 25 271
rect 23 270 24 271
rect 22 270 23 271
rect 21 270 22 271
rect 20 270 21 271
rect 19 270 20 271
rect 18 270 19 271
rect 17 270 18 271
rect 144 271 145 272
rect 143 271 144 272
rect 142 271 143 272
rect 141 271 142 272
rect 140 271 141 272
rect 139 271 140 272
rect 138 271 139 272
rect 137 271 138 272
rect 136 271 137 272
rect 135 271 136 272
rect 134 271 135 272
rect 133 271 134 272
rect 132 271 133 272
rect 131 271 132 272
rect 130 271 131 272
rect 129 271 130 272
rect 128 271 129 272
rect 127 271 128 272
rect 126 271 127 272
rect 125 271 126 272
rect 124 271 125 272
rect 123 271 124 272
rect 84 271 85 272
rect 83 271 84 272
rect 82 271 83 272
rect 81 271 82 272
rect 80 271 81 272
rect 79 271 80 272
rect 78 271 79 272
rect 77 271 78 272
rect 76 271 77 272
rect 75 271 76 272
rect 74 271 75 272
rect 73 271 74 272
rect 72 271 73 272
rect 71 271 72 272
rect 70 271 71 272
rect 69 271 70 272
rect 68 271 69 272
rect 67 271 68 272
rect 66 271 67 272
rect 65 271 66 272
rect 64 271 65 272
rect 63 271 64 272
rect 62 271 63 272
rect 61 271 62 272
rect 60 271 61 272
rect 59 271 60 272
rect 58 271 59 272
rect 57 271 58 272
rect 56 271 57 272
rect 55 271 56 272
rect 54 271 55 272
rect 53 271 54 272
rect 52 271 53 272
rect 51 271 52 272
rect 50 271 51 272
rect 49 271 50 272
rect 48 271 49 272
rect 47 271 48 272
rect 46 271 47 272
rect 45 271 46 272
rect 44 271 45 272
rect 43 271 44 272
rect 42 271 43 272
rect 41 271 42 272
rect 31 271 32 272
rect 30 271 31 272
rect 29 271 30 272
rect 28 271 29 272
rect 27 271 28 272
rect 26 271 27 272
rect 25 271 26 272
rect 24 271 25 272
rect 23 271 24 272
rect 22 271 23 272
rect 21 271 22 272
rect 20 271 21 272
rect 19 271 20 272
rect 18 271 19 272
rect 17 271 18 272
rect 145 272 146 273
rect 144 272 145 273
rect 143 272 144 273
rect 142 272 143 273
rect 141 272 142 273
rect 140 272 141 273
rect 139 272 140 273
rect 138 272 139 273
rect 137 272 138 273
rect 130 272 131 273
rect 129 272 130 273
rect 128 272 129 273
rect 127 272 128 273
rect 126 272 127 273
rect 125 272 126 273
rect 124 272 125 273
rect 123 272 124 273
rect 84 272 85 273
rect 83 272 84 273
rect 82 272 83 273
rect 81 272 82 273
rect 80 272 81 273
rect 79 272 80 273
rect 78 272 79 273
rect 77 272 78 273
rect 76 272 77 273
rect 75 272 76 273
rect 74 272 75 273
rect 73 272 74 273
rect 72 272 73 273
rect 71 272 72 273
rect 70 272 71 273
rect 69 272 70 273
rect 68 272 69 273
rect 67 272 68 273
rect 66 272 67 273
rect 65 272 66 273
rect 64 272 65 273
rect 63 272 64 273
rect 62 272 63 273
rect 61 272 62 273
rect 60 272 61 273
rect 59 272 60 273
rect 58 272 59 273
rect 57 272 58 273
rect 56 272 57 273
rect 55 272 56 273
rect 54 272 55 273
rect 53 272 54 273
rect 52 272 53 273
rect 51 272 52 273
rect 50 272 51 273
rect 49 272 50 273
rect 48 272 49 273
rect 47 272 48 273
rect 46 272 47 273
rect 45 272 46 273
rect 44 272 45 273
rect 43 272 44 273
rect 42 272 43 273
rect 41 272 42 273
rect 31 272 32 273
rect 30 272 31 273
rect 29 272 30 273
rect 28 272 29 273
rect 27 272 28 273
rect 26 272 27 273
rect 25 272 26 273
rect 24 272 25 273
rect 23 272 24 273
rect 22 272 23 273
rect 21 272 22 273
rect 20 272 21 273
rect 19 272 20 273
rect 18 272 19 273
rect 17 272 18 273
rect 145 273 146 274
rect 144 273 145 274
rect 143 273 144 274
rect 142 273 143 274
rect 141 273 142 274
rect 140 273 141 274
rect 139 273 140 274
rect 128 273 129 274
rect 127 273 128 274
rect 126 273 127 274
rect 125 273 126 274
rect 124 273 125 274
rect 123 273 124 274
rect 122 273 123 274
rect 83 273 84 274
rect 82 273 83 274
rect 81 273 82 274
rect 80 273 81 274
rect 79 273 80 274
rect 78 273 79 274
rect 77 273 78 274
rect 76 273 77 274
rect 75 273 76 274
rect 74 273 75 274
rect 73 273 74 274
rect 72 273 73 274
rect 71 273 72 274
rect 70 273 71 274
rect 69 273 70 274
rect 68 273 69 274
rect 67 273 68 274
rect 66 273 67 274
rect 65 273 66 274
rect 64 273 65 274
rect 63 273 64 274
rect 62 273 63 274
rect 61 273 62 274
rect 60 273 61 274
rect 59 273 60 274
rect 58 273 59 274
rect 57 273 58 274
rect 56 273 57 274
rect 55 273 56 274
rect 54 273 55 274
rect 53 273 54 274
rect 52 273 53 274
rect 51 273 52 274
rect 50 273 51 274
rect 49 273 50 274
rect 48 273 49 274
rect 47 273 48 274
rect 46 273 47 274
rect 45 273 46 274
rect 44 273 45 274
rect 43 273 44 274
rect 42 273 43 274
rect 41 273 42 274
rect 31 273 32 274
rect 30 273 31 274
rect 29 273 30 274
rect 28 273 29 274
rect 27 273 28 274
rect 26 273 27 274
rect 25 273 26 274
rect 24 273 25 274
rect 23 273 24 274
rect 22 273 23 274
rect 21 273 22 274
rect 20 273 21 274
rect 19 273 20 274
rect 18 273 19 274
rect 17 273 18 274
rect 145 274 146 275
rect 144 274 145 275
rect 143 274 144 275
rect 142 274 143 275
rect 141 274 142 275
rect 140 274 141 275
rect 127 274 128 275
rect 126 274 127 275
rect 125 274 126 275
rect 124 274 125 275
rect 123 274 124 275
rect 122 274 123 275
rect 83 274 84 275
rect 82 274 83 275
rect 81 274 82 275
rect 80 274 81 275
rect 79 274 80 275
rect 78 274 79 275
rect 77 274 78 275
rect 76 274 77 275
rect 75 274 76 275
rect 74 274 75 275
rect 73 274 74 275
rect 72 274 73 275
rect 71 274 72 275
rect 70 274 71 275
rect 69 274 70 275
rect 68 274 69 275
rect 67 274 68 275
rect 66 274 67 275
rect 65 274 66 275
rect 64 274 65 275
rect 63 274 64 275
rect 62 274 63 275
rect 61 274 62 275
rect 60 274 61 275
rect 59 274 60 275
rect 58 274 59 275
rect 57 274 58 275
rect 56 274 57 275
rect 55 274 56 275
rect 54 274 55 275
rect 53 274 54 275
rect 52 274 53 275
rect 51 274 52 275
rect 50 274 51 275
rect 49 274 50 275
rect 48 274 49 275
rect 47 274 48 275
rect 46 274 47 275
rect 45 274 46 275
rect 44 274 45 275
rect 43 274 44 275
rect 42 274 43 275
rect 41 274 42 275
rect 31 274 32 275
rect 30 274 31 275
rect 29 274 30 275
rect 28 274 29 275
rect 27 274 28 275
rect 26 274 27 275
rect 25 274 26 275
rect 24 274 25 275
rect 23 274 24 275
rect 22 274 23 275
rect 21 274 22 275
rect 20 274 21 275
rect 19 274 20 275
rect 18 274 19 275
rect 17 274 18 275
rect 146 275 147 276
rect 145 275 146 276
rect 144 275 145 276
rect 143 275 144 276
rect 142 275 143 276
rect 141 275 142 276
rect 126 275 127 276
rect 125 275 126 276
rect 124 275 125 276
rect 123 275 124 276
rect 122 275 123 276
rect 83 275 84 276
rect 82 275 83 276
rect 81 275 82 276
rect 80 275 81 276
rect 79 275 80 276
rect 78 275 79 276
rect 77 275 78 276
rect 76 275 77 276
rect 75 275 76 276
rect 74 275 75 276
rect 73 275 74 276
rect 72 275 73 276
rect 71 275 72 276
rect 70 275 71 276
rect 69 275 70 276
rect 68 275 69 276
rect 67 275 68 276
rect 66 275 67 276
rect 65 275 66 276
rect 64 275 65 276
rect 63 275 64 276
rect 62 275 63 276
rect 61 275 62 276
rect 60 275 61 276
rect 59 275 60 276
rect 58 275 59 276
rect 57 275 58 276
rect 56 275 57 276
rect 55 275 56 276
rect 54 275 55 276
rect 53 275 54 276
rect 52 275 53 276
rect 51 275 52 276
rect 50 275 51 276
rect 49 275 50 276
rect 48 275 49 276
rect 47 275 48 276
rect 46 275 47 276
rect 45 275 46 276
rect 44 275 45 276
rect 43 275 44 276
rect 42 275 43 276
rect 41 275 42 276
rect 31 275 32 276
rect 30 275 31 276
rect 29 275 30 276
rect 28 275 29 276
rect 27 275 28 276
rect 26 275 27 276
rect 25 275 26 276
rect 24 275 25 276
rect 23 275 24 276
rect 22 275 23 276
rect 21 275 22 276
rect 20 275 21 276
rect 19 275 20 276
rect 18 275 19 276
rect 17 275 18 276
rect 146 276 147 277
rect 145 276 146 277
rect 144 276 145 277
rect 143 276 144 277
rect 142 276 143 277
rect 126 276 127 277
rect 125 276 126 277
rect 124 276 125 277
rect 123 276 124 277
rect 122 276 123 277
rect 121 276 122 277
rect 82 276 83 277
rect 81 276 82 277
rect 80 276 81 277
rect 79 276 80 277
rect 78 276 79 277
rect 77 276 78 277
rect 76 276 77 277
rect 75 276 76 277
rect 74 276 75 277
rect 73 276 74 277
rect 72 276 73 277
rect 71 276 72 277
rect 70 276 71 277
rect 69 276 70 277
rect 68 276 69 277
rect 67 276 68 277
rect 66 276 67 277
rect 65 276 66 277
rect 64 276 65 277
rect 63 276 64 277
rect 62 276 63 277
rect 61 276 62 277
rect 60 276 61 277
rect 59 276 60 277
rect 58 276 59 277
rect 57 276 58 277
rect 56 276 57 277
rect 55 276 56 277
rect 54 276 55 277
rect 53 276 54 277
rect 52 276 53 277
rect 51 276 52 277
rect 50 276 51 277
rect 49 276 50 277
rect 48 276 49 277
rect 47 276 48 277
rect 46 276 47 277
rect 45 276 46 277
rect 44 276 45 277
rect 43 276 44 277
rect 42 276 43 277
rect 31 276 32 277
rect 30 276 31 277
rect 29 276 30 277
rect 28 276 29 277
rect 27 276 28 277
rect 26 276 27 277
rect 25 276 26 277
rect 24 276 25 277
rect 23 276 24 277
rect 22 276 23 277
rect 21 276 22 277
rect 20 276 21 277
rect 19 276 20 277
rect 18 276 19 277
rect 17 276 18 277
rect 146 277 147 278
rect 145 277 146 278
rect 144 277 145 278
rect 143 277 144 278
rect 142 277 143 278
rect 125 277 126 278
rect 124 277 125 278
rect 123 277 124 278
rect 122 277 123 278
rect 121 277 122 278
rect 82 277 83 278
rect 81 277 82 278
rect 80 277 81 278
rect 79 277 80 278
rect 78 277 79 278
rect 77 277 78 278
rect 76 277 77 278
rect 75 277 76 278
rect 74 277 75 278
rect 73 277 74 278
rect 72 277 73 278
rect 71 277 72 278
rect 70 277 71 278
rect 69 277 70 278
rect 68 277 69 278
rect 67 277 68 278
rect 66 277 67 278
rect 65 277 66 278
rect 64 277 65 278
rect 63 277 64 278
rect 62 277 63 278
rect 61 277 62 278
rect 60 277 61 278
rect 59 277 60 278
rect 58 277 59 278
rect 57 277 58 278
rect 56 277 57 278
rect 55 277 56 278
rect 54 277 55 278
rect 53 277 54 278
rect 52 277 53 278
rect 51 277 52 278
rect 50 277 51 278
rect 49 277 50 278
rect 48 277 49 278
rect 47 277 48 278
rect 46 277 47 278
rect 45 277 46 278
rect 44 277 45 278
rect 43 277 44 278
rect 42 277 43 278
rect 31 277 32 278
rect 30 277 31 278
rect 29 277 30 278
rect 28 277 29 278
rect 27 277 28 278
rect 26 277 27 278
rect 25 277 26 278
rect 24 277 25 278
rect 23 277 24 278
rect 22 277 23 278
rect 21 277 22 278
rect 20 277 21 278
rect 19 277 20 278
rect 18 277 19 278
rect 17 277 18 278
rect 146 278 147 279
rect 145 278 146 279
rect 144 278 145 279
rect 143 278 144 279
rect 142 278 143 279
rect 136 278 137 279
rect 135 278 136 279
rect 134 278 135 279
rect 133 278 134 279
rect 132 278 133 279
rect 125 278 126 279
rect 124 278 125 279
rect 123 278 124 279
rect 122 278 123 279
rect 121 278 122 279
rect 81 278 82 279
rect 80 278 81 279
rect 79 278 80 279
rect 78 278 79 279
rect 77 278 78 279
rect 76 278 77 279
rect 75 278 76 279
rect 74 278 75 279
rect 73 278 74 279
rect 72 278 73 279
rect 71 278 72 279
rect 70 278 71 279
rect 69 278 70 279
rect 68 278 69 279
rect 67 278 68 279
rect 66 278 67 279
rect 65 278 66 279
rect 64 278 65 279
rect 63 278 64 279
rect 62 278 63 279
rect 61 278 62 279
rect 60 278 61 279
rect 59 278 60 279
rect 58 278 59 279
rect 57 278 58 279
rect 56 278 57 279
rect 55 278 56 279
rect 54 278 55 279
rect 53 278 54 279
rect 52 278 53 279
rect 51 278 52 279
rect 50 278 51 279
rect 49 278 50 279
rect 48 278 49 279
rect 47 278 48 279
rect 46 278 47 279
rect 45 278 46 279
rect 44 278 45 279
rect 43 278 44 279
rect 42 278 43 279
rect 31 278 32 279
rect 30 278 31 279
rect 29 278 30 279
rect 28 278 29 279
rect 27 278 28 279
rect 26 278 27 279
rect 25 278 26 279
rect 24 278 25 279
rect 23 278 24 279
rect 22 278 23 279
rect 21 278 22 279
rect 20 278 21 279
rect 19 278 20 279
rect 18 278 19 279
rect 17 278 18 279
rect 146 279 147 280
rect 145 279 146 280
rect 144 279 145 280
rect 143 279 144 280
rect 142 279 143 280
rect 136 279 137 280
rect 135 279 136 280
rect 134 279 135 280
rect 133 279 134 280
rect 132 279 133 280
rect 125 279 126 280
rect 124 279 125 280
rect 123 279 124 280
rect 122 279 123 280
rect 121 279 122 280
rect 80 279 81 280
rect 79 279 80 280
rect 78 279 79 280
rect 77 279 78 280
rect 76 279 77 280
rect 75 279 76 280
rect 74 279 75 280
rect 73 279 74 280
rect 72 279 73 280
rect 71 279 72 280
rect 70 279 71 280
rect 69 279 70 280
rect 68 279 69 280
rect 67 279 68 280
rect 66 279 67 280
rect 65 279 66 280
rect 64 279 65 280
rect 63 279 64 280
rect 62 279 63 280
rect 61 279 62 280
rect 60 279 61 280
rect 59 279 60 280
rect 58 279 59 280
rect 57 279 58 280
rect 56 279 57 280
rect 55 279 56 280
rect 54 279 55 280
rect 53 279 54 280
rect 52 279 53 280
rect 51 279 52 280
rect 50 279 51 280
rect 49 279 50 280
rect 48 279 49 280
rect 47 279 48 280
rect 46 279 47 280
rect 45 279 46 280
rect 44 279 45 280
rect 43 279 44 280
rect 31 279 32 280
rect 30 279 31 280
rect 29 279 30 280
rect 28 279 29 280
rect 27 279 28 280
rect 26 279 27 280
rect 25 279 26 280
rect 24 279 25 280
rect 23 279 24 280
rect 22 279 23 280
rect 21 279 22 280
rect 20 279 21 280
rect 19 279 20 280
rect 18 279 19 280
rect 146 280 147 281
rect 145 280 146 281
rect 144 280 145 281
rect 143 280 144 281
rect 142 280 143 281
rect 136 280 137 281
rect 135 280 136 281
rect 134 280 135 281
rect 133 280 134 281
rect 132 280 133 281
rect 125 280 126 281
rect 124 280 125 281
rect 123 280 124 281
rect 122 280 123 281
rect 121 280 122 281
rect 80 280 81 281
rect 79 280 80 281
rect 78 280 79 281
rect 77 280 78 281
rect 76 280 77 281
rect 75 280 76 281
rect 74 280 75 281
rect 73 280 74 281
rect 72 280 73 281
rect 71 280 72 281
rect 70 280 71 281
rect 69 280 70 281
rect 68 280 69 281
rect 67 280 68 281
rect 66 280 67 281
rect 65 280 66 281
rect 64 280 65 281
rect 63 280 64 281
rect 62 280 63 281
rect 61 280 62 281
rect 60 280 61 281
rect 59 280 60 281
rect 58 280 59 281
rect 57 280 58 281
rect 56 280 57 281
rect 55 280 56 281
rect 54 280 55 281
rect 53 280 54 281
rect 52 280 53 281
rect 51 280 52 281
rect 50 280 51 281
rect 49 280 50 281
rect 48 280 49 281
rect 47 280 48 281
rect 46 280 47 281
rect 45 280 46 281
rect 44 280 45 281
rect 43 280 44 281
rect 31 280 32 281
rect 30 280 31 281
rect 29 280 30 281
rect 28 280 29 281
rect 27 280 28 281
rect 26 280 27 281
rect 25 280 26 281
rect 24 280 25 281
rect 23 280 24 281
rect 22 280 23 281
rect 21 280 22 281
rect 20 280 21 281
rect 19 280 20 281
rect 18 280 19 281
rect 146 281 147 282
rect 145 281 146 282
rect 144 281 145 282
rect 143 281 144 282
rect 142 281 143 282
rect 136 281 137 282
rect 135 281 136 282
rect 134 281 135 282
rect 133 281 134 282
rect 132 281 133 282
rect 125 281 126 282
rect 124 281 125 282
rect 123 281 124 282
rect 122 281 123 282
rect 121 281 122 282
rect 79 281 80 282
rect 78 281 79 282
rect 77 281 78 282
rect 76 281 77 282
rect 75 281 76 282
rect 74 281 75 282
rect 73 281 74 282
rect 72 281 73 282
rect 71 281 72 282
rect 70 281 71 282
rect 69 281 70 282
rect 68 281 69 282
rect 67 281 68 282
rect 66 281 67 282
rect 65 281 66 282
rect 64 281 65 282
rect 63 281 64 282
rect 62 281 63 282
rect 61 281 62 282
rect 60 281 61 282
rect 59 281 60 282
rect 58 281 59 282
rect 57 281 58 282
rect 56 281 57 282
rect 55 281 56 282
rect 54 281 55 282
rect 53 281 54 282
rect 52 281 53 282
rect 51 281 52 282
rect 50 281 51 282
rect 49 281 50 282
rect 48 281 49 282
rect 47 281 48 282
rect 46 281 47 282
rect 45 281 46 282
rect 44 281 45 282
rect 32 281 33 282
rect 31 281 32 282
rect 30 281 31 282
rect 29 281 30 282
rect 28 281 29 282
rect 27 281 28 282
rect 26 281 27 282
rect 25 281 26 282
rect 24 281 25 282
rect 23 281 24 282
rect 22 281 23 282
rect 21 281 22 282
rect 20 281 21 282
rect 19 281 20 282
rect 18 281 19 282
rect 146 282 147 283
rect 145 282 146 283
rect 144 282 145 283
rect 143 282 144 283
rect 142 282 143 283
rect 136 282 137 283
rect 135 282 136 283
rect 134 282 135 283
rect 133 282 134 283
rect 132 282 133 283
rect 125 282 126 283
rect 124 282 125 283
rect 123 282 124 283
rect 122 282 123 283
rect 121 282 122 283
rect 78 282 79 283
rect 77 282 78 283
rect 76 282 77 283
rect 75 282 76 283
rect 74 282 75 283
rect 73 282 74 283
rect 72 282 73 283
rect 71 282 72 283
rect 70 282 71 283
rect 69 282 70 283
rect 68 282 69 283
rect 67 282 68 283
rect 66 282 67 283
rect 65 282 66 283
rect 64 282 65 283
rect 63 282 64 283
rect 62 282 63 283
rect 61 282 62 283
rect 60 282 61 283
rect 59 282 60 283
rect 58 282 59 283
rect 57 282 58 283
rect 56 282 57 283
rect 55 282 56 283
rect 54 282 55 283
rect 53 282 54 283
rect 52 282 53 283
rect 51 282 52 283
rect 50 282 51 283
rect 49 282 50 283
rect 48 282 49 283
rect 47 282 48 283
rect 46 282 47 283
rect 45 282 46 283
rect 32 282 33 283
rect 31 282 32 283
rect 30 282 31 283
rect 29 282 30 283
rect 28 282 29 283
rect 27 282 28 283
rect 26 282 27 283
rect 25 282 26 283
rect 24 282 25 283
rect 23 282 24 283
rect 22 282 23 283
rect 21 282 22 283
rect 20 282 21 283
rect 19 282 20 283
rect 18 282 19 283
rect 146 283 147 284
rect 145 283 146 284
rect 144 283 145 284
rect 143 283 144 284
rect 142 283 143 284
rect 141 283 142 284
rect 140 283 141 284
rect 139 283 140 284
rect 138 283 139 284
rect 137 283 138 284
rect 136 283 137 284
rect 135 283 136 284
rect 134 283 135 284
rect 133 283 134 284
rect 132 283 133 284
rect 125 283 126 284
rect 124 283 125 284
rect 123 283 124 284
rect 122 283 123 284
rect 121 283 122 284
rect 77 283 78 284
rect 76 283 77 284
rect 75 283 76 284
rect 74 283 75 284
rect 73 283 74 284
rect 72 283 73 284
rect 71 283 72 284
rect 70 283 71 284
rect 69 283 70 284
rect 68 283 69 284
rect 67 283 68 284
rect 66 283 67 284
rect 65 283 66 284
rect 64 283 65 284
rect 63 283 64 284
rect 62 283 63 284
rect 61 283 62 284
rect 60 283 61 284
rect 59 283 60 284
rect 58 283 59 284
rect 57 283 58 284
rect 56 283 57 284
rect 55 283 56 284
rect 54 283 55 284
rect 53 283 54 284
rect 52 283 53 284
rect 51 283 52 284
rect 50 283 51 284
rect 49 283 50 284
rect 48 283 49 284
rect 47 283 48 284
rect 46 283 47 284
rect 32 283 33 284
rect 31 283 32 284
rect 30 283 31 284
rect 29 283 30 284
rect 28 283 29 284
rect 27 283 28 284
rect 26 283 27 284
rect 25 283 26 284
rect 24 283 25 284
rect 23 283 24 284
rect 22 283 23 284
rect 21 283 22 284
rect 20 283 21 284
rect 19 283 20 284
rect 145 284 146 285
rect 144 284 145 285
rect 143 284 144 285
rect 142 284 143 285
rect 141 284 142 285
rect 140 284 141 285
rect 139 284 140 285
rect 138 284 139 285
rect 137 284 138 285
rect 136 284 137 285
rect 135 284 136 285
rect 134 284 135 285
rect 133 284 134 285
rect 132 284 133 285
rect 125 284 126 285
rect 124 284 125 285
rect 123 284 124 285
rect 122 284 123 285
rect 121 284 122 285
rect 75 284 76 285
rect 74 284 75 285
rect 73 284 74 285
rect 72 284 73 285
rect 71 284 72 285
rect 70 284 71 285
rect 69 284 70 285
rect 68 284 69 285
rect 67 284 68 285
rect 66 284 67 285
rect 65 284 66 285
rect 64 284 65 285
rect 63 284 64 285
rect 62 284 63 285
rect 61 284 62 285
rect 60 284 61 285
rect 59 284 60 285
rect 58 284 59 285
rect 57 284 58 285
rect 56 284 57 285
rect 55 284 56 285
rect 54 284 55 285
rect 53 284 54 285
rect 52 284 53 285
rect 51 284 52 285
rect 50 284 51 285
rect 49 284 50 285
rect 48 284 49 285
rect 47 284 48 285
rect 145 285 146 286
rect 144 285 145 286
rect 143 285 144 286
rect 142 285 143 286
rect 141 285 142 286
rect 140 285 141 286
rect 139 285 140 286
rect 138 285 139 286
rect 137 285 138 286
rect 136 285 137 286
rect 135 285 136 286
rect 134 285 135 286
rect 133 285 134 286
rect 132 285 133 286
rect 126 285 127 286
rect 125 285 126 286
rect 124 285 125 286
rect 123 285 124 286
rect 122 285 123 286
rect 74 285 75 286
rect 73 285 74 286
rect 72 285 73 286
rect 71 285 72 286
rect 70 285 71 286
rect 69 285 70 286
rect 68 285 69 286
rect 67 285 68 286
rect 66 285 67 286
rect 65 285 66 286
rect 64 285 65 286
rect 63 285 64 286
rect 62 285 63 286
rect 61 285 62 286
rect 60 285 61 286
rect 59 285 60 286
rect 58 285 59 286
rect 57 285 58 286
rect 56 285 57 286
rect 55 285 56 286
rect 54 285 55 286
rect 53 285 54 286
rect 52 285 53 286
rect 51 285 52 286
rect 50 285 51 286
rect 49 285 50 286
rect 48 285 49 286
rect 145 286 146 287
rect 144 286 145 287
rect 143 286 144 287
rect 142 286 143 287
rect 141 286 142 287
rect 140 286 141 287
rect 139 286 140 287
rect 138 286 139 287
rect 137 286 138 287
rect 136 286 137 287
rect 135 286 136 287
rect 134 286 135 287
rect 133 286 134 287
rect 132 286 133 287
rect 126 286 127 287
rect 125 286 126 287
rect 124 286 125 287
rect 123 286 124 287
rect 122 286 123 287
rect 72 286 73 287
rect 71 286 72 287
rect 70 286 71 287
rect 69 286 70 287
rect 68 286 69 287
rect 67 286 68 287
rect 66 286 67 287
rect 65 286 66 287
rect 64 286 65 287
rect 63 286 64 287
rect 62 286 63 287
rect 61 286 62 287
rect 60 286 61 287
rect 59 286 60 287
rect 58 286 59 287
rect 57 286 58 287
rect 56 286 57 287
rect 55 286 56 287
rect 54 286 55 287
rect 53 286 54 287
rect 52 286 53 287
rect 51 286 52 287
rect 50 286 51 287
rect 144 287 145 288
rect 143 287 144 288
rect 142 287 143 288
rect 141 287 142 288
rect 140 287 141 288
rect 139 287 140 288
rect 138 287 139 288
rect 137 287 138 288
rect 136 287 137 288
rect 135 287 136 288
rect 134 287 135 288
rect 133 287 134 288
rect 132 287 133 288
rect 70 287 71 288
rect 69 287 70 288
rect 68 287 69 288
rect 67 287 68 288
rect 66 287 67 288
rect 65 287 66 288
rect 64 287 65 288
rect 63 287 64 288
rect 62 287 63 288
rect 61 287 62 288
rect 60 287 61 288
rect 59 287 60 288
rect 58 287 59 288
rect 57 287 58 288
rect 56 287 57 288
rect 55 287 56 288
rect 54 287 55 288
rect 53 287 54 288
rect 52 287 53 288
rect 144 288 145 289
rect 143 288 144 289
rect 142 288 143 289
rect 141 288 142 289
rect 140 288 141 289
rect 139 288 140 289
rect 138 288 139 289
rect 137 288 138 289
rect 136 288 137 289
rect 135 288 136 289
rect 134 288 135 289
rect 133 288 134 289
rect 132 288 133 289
rect 66 288 67 289
rect 65 288 66 289
rect 64 288 65 289
rect 63 288 64 289
rect 62 288 63 289
rect 61 288 62 289
rect 60 288 61 289
rect 59 288 60 289
rect 58 288 59 289
rect 57 288 58 289
rect 56 288 57 289
rect 138 292 139 293
rect 137 292 138 293
rect 136 292 137 293
rect 141 293 142 294
rect 140 293 141 294
rect 139 293 140 294
rect 138 293 139 294
rect 137 293 138 294
rect 136 293 137 294
rect 135 293 136 294
rect 134 293 135 294
rect 133 293 134 294
rect 143 294 144 295
rect 142 294 143 295
rect 141 294 142 295
rect 140 294 141 295
rect 139 294 140 295
rect 138 294 139 295
rect 137 294 138 295
rect 136 294 137 295
rect 135 294 136 295
rect 134 294 135 295
rect 133 294 134 295
rect 132 294 133 295
rect 131 294 132 295
rect 144 295 145 296
rect 143 295 144 296
rect 142 295 143 296
rect 141 295 142 296
rect 140 295 141 296
rect 139 295 140 296
rect 138 295 139 296
rect 137 295 138 296
rect 136 295 137 296
rect 135 295 136 296
rect 134 295 135 296
rect 133 295 134 296
rect 132 295 133 296
rect 131 295 132 296
rect 130 295 131 296
rect 145 296 146 297
rect 144 296 145 297
rect 143 296 144 297
rect 142 296 143 297
rect 141 296 142 297
rect 140 296 141 297
rect 139 296 140 297
rect 138 296 139 297
rect 137 296 138 297
rect 136 296 137 297
rect 135 296 136 297
rect 134 296 135 297
rect 133 296 134 297
rect 132 296 133 297
rect 131 296 132 297
rect 130 296 131 297
rect 129 296 130 297
rect 145 297 146 298
rect 144 297 145 298
rect 143 297 144 298
rect 142 297 143 298
rect 141 297 142 298
rect 140 297 141 298
rect 139 297 140 298
rect 138 297 139 298
rect 137 297 138 298
rect 136 297 137 298
rect 135 297 136 298
rect 134 297 135 298
rect 133 297 134 298
rect 132 297 133 298
rect 131 297 132 298
rect 130 297 131 298
rect 129 297 130 298
rect 145 298 146 299
rect 144 298 145 299
rect 143 298 144 299
rect 142 298 143 299
rect 141 298 142 299
rect 140 298 141 299
rect 134 298 135 299
rect 133 298 134 299
rect 132 298 133 299
rect 131 298 132 299
rect 130 298 131 299
rect 129 298 130 299
rect 83 298 84 299
rect 82 298 83 299
rect 81 298 82 299
rect 80 298 81 299
rect 79 298 80 299
rect 78 298 79 299
rect 77 298 78 299
rect 76 298 77 299
rect 75 298 76 299
rect 74 298 75 299
rect 73 298 74 299
rect 72 298 73 299
rect 71 298 72 299
rect 70 298 71 299
rect 69 298 70 299
rect 68 298 69 299
rect 146 299 147 300
rect 145 299 146 300
rect 144 299 145 300
rect 143 299 144 300
rect 142 299 143 300
rect 132 299 133 300
rect 131 299 132 300
rect 130 299 131 300
rect 129 299 130 300
rect 128 299 129 300
rect 83 299 84 300
rect 82 299 83 300
rect 81 299 82 300
rect 80 299 81 300
rect 79 299 80 300
rect 78 299 79 300
rect 77 299 78 300
rect 76 299 77 300
rect 75 299 76 300
rect 74 299 75 300
rect 73 299 74 300
rect 72 299 73 300
rect 71 299 72 300
rect 70 299 71 300
rect 69 299 70 300
rect 146 300 147 301
rect 145 300 146 301
rect 144 300 145 301
rect 143 300 144 301
rect 142 300 143 301
rect 132 300 133 301
rect 131 300 132 301
rect 130 300 131 301
rect 129 300 130 301
rect 128 300 129 301
rect 83 300 84 301
rect 82 300 83 301
rect 81 300 82 301
rect 80 300 81 301
rect 79 300 80 301
rect 78 300 79 301
rect 77 300 78 301
rect 76 300 77 301
rect 75 300 76 301
rect 74 300 75 301
rect 73 300 74 301
rect 72 300 73 301
rect 71 300 72 301
rect 70 300 71 301
rect 69 300 70 301
rect 57 300 58 301
rect 56 300 57 301
rect 55 300 56 301
rect 54 300 55 301
rect 53 300 54 301
rect 52 300 53 301
rect 51 300 52 301
rect 50 300 51 301
rect 49 300 50 301
rect 48 300 49 301
rect 47 300 48 301
rect 46 300 47 301
rect 45 300 46 301
rect 44 300 45 301
rect 43 300 44 301
rect 42 300 43 301
rect 146 301 147 302
rect 145 301 146 302
rect 144 301 145 302
rect 143 301 144 302
rect 131 301 132 302
rect 130 301 131 302
rect 129 301 130 302
rect 128 301 129 302
rect 83 301 84 302
rect 82 301 83 302
rect 81 301 82 302
rect 80 301 81 302
rect 79 301 80 302
rect 78 301 79 302
rect 77 301 78 302
rect 76 301 77 302
rect 75 301 76 302
rect 74 301 75 302
rect 73 301 74 302
rect 72 301 73 302
rect 71 301 72 302
rect 70 301 71 302
rect 69 301 70 302
rect 57 301 58 302
rect 56 301 57 302
rect 55 301 56 302
rect 54 301 55 302
rect 53 301 54 302
rect 52 301 53 302
rect 51 301 52 302
rect 50 301 51 302
rect 49 301 50 302
rect 48 301 49 302
rect 47 301 48 302
rect 46 301 47 302
rect 45 301 46 302
rect 44 301 45 302
rect 43 301 44 302
rect 42 301 43 302
rect 41 301 42 302
rect 40 301 41 302
rect 39 301 40 302
rect 38 301 39 302
rect 37 301 38 302
rect 36 301 37 302
rect 35 301 36 302
rect 34 301 35 302
rect 33 301 34 302
rect 32 301 33 302
rect 31 301 32 302
rect 30 301 31 302
rect 29 301 30 302
rect 28 301 29 302
rect 27 301 28 302
rect 26 301 27 302
rect 146 302 147 303
rect 145 302 146 303
rect 144 302 145 303
rect 143 302 144 303
rect 131 302 132 303
rect 130 302 131 303
rect 129 302 130 303
rect 128 302 129 303
rect 84 302 85 303
rect 83 302 84 303
rect 82 302 83 303
rect 81 302 82 303
rect 80 302 81 303
rect 79 302 80 303
rect 78 302 79 303
rect 77 302 78 303
rect 76 302 77 303
rect 75 302 76 303
rect 74 302 75 303
rect 73 302 74 303
rect 72 302 73 303
rect 71 302 72 303
rect 70 302 71 303
rect 56 302 57 303
rect 55 302 56 303
rect 54 302 55 303
rect 53 302 54 303
rect 52 302 53 303
rect 51 302 52 303
rect 50 302 51 303
rect 49 302 50 303
rect 48 302 49 303
rect 47 302 48 303
rect 46 302 47 303
rect 45 302 46 303
rect 44 302 45 303
rect 43 302 44 303
rect 42 302 43 303
rect 41 302 42 303
rect 40 302 41 303
rect 39 302 40 303
rect 38 302 39 303
rect 37 302 38 303
rect 36 302 37 303
rect 35 302 36 303
rect 34 302 35 303
rect 33 302 34 303
rect 32 302 33 303
rect 31 302 32 303
rect 30 302 31 303
rect 29 302 30 303
rect 28 302 29 303
rect 27 302 28 303
rect 26 302 27 303
rect 25 302 26 303
rect 24 302 25 303
rect 23 302 24 303
rect 22 302 23 303
rect 21 302 22 303
rect 20 302 21 303
rect 19 302 20 303
rect 18 302 19 303
rect 146 303 147 304
rect 145 303 146 304
rect 144 303 145 304
rect 143 303 144 304
rect 131 303 132 304
rect 130 303 131 304
rect 129 303 130 304
rect 128 303 129 304
rect 84 303 85 304
rect 83 303 84 304
rect 82 303 83 304
rect 81 303 82 304
rect 80 303 81 304
rect 79 303 80 304
rect 78 303 79 304
rect 77 303 78 304
rect 76 303 77 304
rect 75 303 76 304
rect 74 303 75 304
rect 73 303 74 304
rect 72 303 73 304
rect 71 303 72 304
rect 70 303 71 304
rect 56 303 57 304
rect 55 303 56 304
rect 54 303 55 304
rect 53 303 54 304
rect 52 303 53 304
rect 51 303 52 304
rect 50 303 51 304
rect 49 303 50 304
rect 48 303 49 304
rect 47 303 48 304
rect 46 303 47 304
rect 45 303 46 304
rect 44 303 45 304
rect 43 303 44 304
rect 42 303 43 304
rect 41 303 42 304
rect 40 303 41 304
rect 39 303 40 304
rect 38 303 39 304
rect 37 303 38 304
rect 36 303 37 304
rect 35 303 36 304
rect 34 303 35 304
rect 33 303 34 304
rect 32 303 33 304
rect 31 303 32 304
rect 30 303 31 304
rect 29 303 30 304
rect 28 303 29 304
rect 27 303 28 304
rect 26 303 27 304
rect 25 303 26 304
rect 24 303 25 304
rect 23 303 24 304
rect 22 303 23 304
rect 21 303 22 304
rect 20 303 21 304
rect 19 303 20 304
rect 18 303 19 304
rect 146 304 147 305
rect 145 304 146 305
rect 144 304 145 305
rect 143 304 144 305
rect 142 304 143 305
rect 132 304 133 305
rect 131 304 132 305
rect 130 304 131 305
rect 129 304 130 305
rect 128 304 129 305
rect 84 304 85 305
rect 83 304 84 305
rect 82 304 83 305
rect 81 304 82 305
rect 80 304 81 305
rect 79 304 80 305
rect 78 304 79 305
rect 77 304 78 305
rect 76 304 77 305
rect 75 304 76 305
rect 74 304 75 305
rect 73 304 74 305
rect 72 304 73 305
rect 71 304 72 305
rect 70 304 71 305
rect 56 304 57 305
rect 55 304 56 305
rect 54 304 55 305
rect 53 304 54 305
rect 52 304 53 305
rect 51 304 52 305
rect 50 304 51 305
rect 49 304 50 305
rect 48 304 49 305
rect 47 304 48 305
rect 46 304 47 305
rect 45 304 46 305
rect 44 304 45 305
rect 43 304 44 305
rect 42 304 43 305
rect 41 304 42 305
rect 40 304 41 305
rect 39 304 40 305
rect 38 304 39 305
rect 37 304 38 305
rect 36 304 37 305
rect 35 304 36 305
rect 34 304 35 305
rect 33 304 34 305
rect 32 304 33 305
rect 31 304 32 305
rect 30 304 31 305
rect 29 304 30 305
rect 28 304 29 305
rect 27 304 28 305
rect 26 304 27 305
rect 25 304 26 305
rect 24 304 25 305
rect 23 304 24 305
rect 22 304 23 305
rect 21 304 22 305
rect 20 304 21 305
rect 19 304 20 305
rect 18 304 19 305
rect 146 305 147 306
rect 145 305 146 306
rect 144 305 145 306
rect 143 305 144 306
rect 142 305 143 306
rect 141 305 142 306
rect 133 305 134 306
rect 132 305 133 306
rect 131 305 132 306
rect 130 305 131 306
rect 129 305 130 306
rect 128 305 129 306
rect 84 305 85 306
rect 83 305 84 306
rect 82 305 83 306
rect 81 305 82 306
rect 80 305 81 306
rect 79 305 80 306
rect 78 305 79 306
rect 77 305 78 306
rect 76 305 77 306
rect 75 305 76 306
rect 74 305 75 306
rect 73 305 74 306
rect 72 305 73 306
rect 71 305 72 306
rect 70 305 71 306
rect 56 305 57 306
rect 55 305 56 306
rect 54 305 55 306
rect 53 305 54 306
rect 52 305 53 306
rect 51 305 52 306
rect 50 305 51 306
rect 49 305 50 306
rect 48 305 49 306
rect 47 305 48 306
rect 46 305 47 306
rect 45 305 46 306
rect 44 305 45 306
rect 43 305 44 306
rect 42 305 43 306
rect 41 305 42 306
rect 40 305 41 306
rect 39 305 40 306
rect 38 305 39 306
rect 37 305 38 306
rect 36 305 37 306
rect 35 305 36 306
rect 34 305 35 306
rect 33 305 34 306
rect 32 305 33 306
rect 31 305 32 306
rect 30 305 31 306
rect 29 305 30 306
rect 28 305 29 306
rect 27 305 28 306
rect 26 305 27 306
rect 25 305 26 306
rect 24 305 25 306
rect 23 305 24 306
rect 22 305 23 306
rect 21 305 22 306
rect 20 305 21 306
rect 19 305 20 306
rect 18 305 19 306
rect 145 306 146 307
rect 144 306 145 307
rect 143 306 144 307
rect 142 306 143 307
rect 141 306 142 307
rect 140 306 141 307
rect 139 306 140 307
rect 135 306 136 307
rect 134 306 135 307
rect 133 306 134 307
rect 132 306 133 307
rect 131 306 132 307
rect 130 306 131 307
rect 129 306 130 307
rect 84 306 85 307
rect 83 306 84 307
rect 82 306 83 307
rect 81 306 82 307
rect 80 306 81 307
rect 79 306 80 307
rect 78 306 79 307
rect 77 306 78 307
rect 76 306 77 307
rect 75 306 76 307
rect 74 306 75 307
rect 73 306 74 307
rect 72 306 73 307
rect 71 306 72 307
rect 56 306 57 307
rect 55 306 56 307
rect 54 306 55 307
rect 53 306 54 307
rect 52 306 53 307
rect 51 306 52 307
rect 50 306 51 307
rect 49 306 50 307
rect 48 306 49 307
rect 47 306 48 307
rect 46 306 47 307
rect 45 306 46 307
rect 44 306 45 307
rect 43 306 44 307
rect 42 306 43 307
rect 41 306 42 307
rect 40 306 41 307
rect 39 306 40 307
rect 38 306 39 307
rect 37 306 38 307
rect 36 306 37 307
rect 35 306 36 307
rect 34 306 35 307
rect 33 306 34 307
rect 32 306 33 307
rect 31 306 32 307
rect 30 306 31 307
rect 29 306 30 307
rect 28 306 29 307
rect 27 306 28 307
rect 26 306 27 307
rect 25 306 26 307
rect 24 306 25 307
rect 23 306 24 307
rect 22 306 23 307
rect 21 306 22 307
rect 20 306 21 307
rect 19 306 20 307
rect 18 306 19 307
rect 145 307 146 308
rect 144 307 145 308
rect 143 307 144 308
rect 142 307 143 308
rect 141 307 142 308
rect 140 307 141 308
rect 139 307 140 308
rect 138 307 139 308
rect 137 307 138 308
rect 136 307 137 308
rect 135 307 136 308
rect 134 307 135 308
rect 133 307 134 308
rect 132 307 133 308
rect 131 307 132 308
rect 130 307 131 308
rect 129 307 130 308
rect 84 307 85 308
rect 83 307 84 308
rect 82 307 83 308
rect 81 307 82 308
rect 80 307 81 308
rect 79 307 80 308
rect 78 307 79 308
rect 77 307 78 308
rect 76 307 77 308
rect 75 307 76 308
rect 74 307 75 308
rect 73 307 74 308
rect 72 307 73 308
rect 71 307 72 308
rect 56 307 57 308
rect 55 307 56 308
rect 54 307 55 308
rect 53 307 54 308
rect 52 307 53 308
rect 51 307 52 308
rect 50 307 51 308
rect 49 307 50 308
rect 48 307 49 308
rect 47 307 48 308
rect 46 307 47 308
rect 45 307 46 308
rect 44 307 45 308
rect 43 307 44 308
rect 42 307 43 308
rect 41 307 42 308
rect 40 307 41 308
rect 39 307 40 308
rect 38 307 39 308
rect 37 307 38 308
rect 36 307 37 308
rect 35 307 36 308
rect 34 307 35 308
rect 33 307 34 308
rect 32 307 33 308
rect 31 307 32 308
rect 30 307 31 308
rect 29 307 30 308
rect 28 307 29 308
rect 27 307 28 308
rect 26 307 27 308
rect 25 307 26 308
rect 24 307 25 308
rect 23 307 24 308
rect 22 307 23 308
rect 21 307 22 308
rect 20 307 21 308
rect 19 307 20 308
rect 18 307 19 308
rect 144 308 145 309
rect 143 308 144 309
rect 142 308 143 309
rect 141 308 142 309
rect 140 308 141 309
rect 139 308 140 309
rect 138 308 139 309
rect 137 308 138 309
rect 136 308 137 309
rect 135 308 136 309
rect 134 308 135 309
rect 133 308 134 309
rect 132 308 133 309
rect 131 308 132 309
rect 130 308 131 309
rect 84 308 85 309
rect 83 308 84 309
rect 82 308 83 309
rect 81 308 82 309
rect 80 308 81 309
rect 79 308 80 309
rect 78 308 79 309
rect 77 308 78 309
rect 76 308 77 309
rect 75 308 76 309
rect 74 308 75 309
rect 73 308 74 309
rect 72 308 73 309
rect 71 308 72 309
rect 56 308 57 309
rect 55 308 56 309
rect 54 308 55 309
rect 53 308 54 309
rect 52 308 53 309
rect 51 308 52 309
rect 50 308 51 309
rect 49 308 50 309
rect 48 308 49 309
rect 47 308 48 309
rect 46 308 47 309
rect 45 308 46 309
rect 44 308 45 309
rect 43 308 44 309
rect 42 308 43 309
rect 41 308 42 309
rect 40 308 41 309
rect 39 308 40 309
rect 38 308 39 309
rect 37 308 38 309
rect 36 308 37 309
rect 35 308 36 309
rect 34 308 35 309
rect 33 308 34 309
rect 32 308 33 309
rect 31 308 32 309
rect 30 308 31 309
rect 29 308 30 309
rect 28 308 29 309
rect 27 308 28 309
rect 26 308 27 309
rect 25 308 26 309
rect 24 308 25 309
rect 23 308 24 309
rect 22 308 23 309
rect 21 308 22 309
rect 20 308 21 309
rect 19 308 20 309
rect 18 308 19 309
rect 143 309 144 310
rect 142 309 143 310
rect 141 309 142 310
rect 140 309 141 310
rect 139 309 140 310
rect 138 309 139 310
rect 137 309 138 310
rect 136 309 137 310
rect 135 309 136 310
rect 134 309 135 310
rect 133 309 134 310
rect 132 309 133 310
rect 131 309 132 310
rect 130 309 131 310
rect 85 309 86 310
rect 84 309 85 310
rect 83 309 84 310
rect 82 309 83 310
rect 81 309 82 310
rect 80 309 81 310
rect 79 309 80 310
rect 78 309 79 310
rect 77 309 78 310
rect 76 309 77 310
rect 75 309 76 310
rect 74 309 75 310
rect 73 309 74 310
rect 72 309 73 310
rect 71 309 72 310
rect 56 309 57 310
rect 55 309 56 310
rect 54 309 55 310
rect 53 309 54 310
rect 52 309 53 310
rect 51 309 52 310
rect 50 309 51 310
rect 49 309 50 310
rect 48 309 49 310
rect 47 309 48 310
rect 46 309 47 310
rect 45 309 46 310
rect 44 309 45 310
rect 43 309 44 310
rect 42 309 43 310
rect 41 309 42 310
rect 40 309 41 310
rect 39 309 40 310
rect 38 309 39 310
rect 37 309 38 310
rect 36 309 37 310
rect 35 309 36 310
rect 34 309 35 310
rect 33 309 34 310
rect 32 309 33 310
rect 31 309 32 310
rect 30 309 31 310
rect 29 309 30 310
rect 28 309 29 310
rect 27 309 28 310
rect 26 309 27 310
rect 25 309 26 310
rect 24 309 25 310
rect 23 309 24 310
rect 22 309 23 310
rect 21 309 22 310
rect 20 309 21 310
rect 19 309 20 310
rect 18 309 19 310
rect 142 310 143 311
rect 141 310 142 311
rect 140 310 141 311
rect 139 310 140 311
rect 138 310 139 311
rect 137 310 138 311
rect 136 310 137 311
rect 135 310 136 311
rect 134 310 135 311
rect 133 310 134 311
rect 132 310 133 311
rect 85 310 86 311
rect 84 310 85 311
rect 83 310 84 311
rect 82 310 83 311
rect 81 310 82 311
rect 80 310 81 311
rect 79 310 80 311
rect 78 310 79 311
rect 77 310 78 311
rect 76 310 77 311
rect 75 310 76 311
rect 74 310 75 311
rect 73 310 74 311
rect 72 310 73 311
rect 71 310 72 311
rect 56 310 57 311
rect 55 310 56 311
rect 54 310 55 311
rect 53 310 54 311
rect 52 310 53 311
rect 51 310 52 311
rect 50 310 51 311
rect 49 310 50 311
rect 48 310 49 311
rect 47 310 48 311
rect 46 310 47 311
rect 45 310 46 311
rect 44 310 45 311
rect 43 310 44 311
rect 42 310 43 311
rect 41 310 42 311
rect 40 310 41 311
rect 39 310 40 311
rect 38 310 39 311
rect 37 310 38 311
rect 36 310 37 311
rect 35 310 36 311
rect 34 310 35 311
rect 33 310 34 311
rect 32 310 33 311
rect 31 310 32 311
rect 30 310 31 311
rect 29 310 30 311
rect 28 310 29 311
rect 27 310 28 311
rect 26 310 27 311
rect 25 310 26 311
rect 24 310 25 311
rect 23 310 24 311
rect 22 310 23 311
rect 21 310 22 311
rect 20 310 21 311
rect 19 310 20 311
rect 18 310 19 311
rect 140 311 141 312
rect 139 311 140 312
rect 138 311 139 312
rect 137 311 138 312
rect 136 311 137 312
rect 135 311 136 312
rect 134 311 135 312
rect 133 311 134 312
rect 85 311 86 312
rect 84 311 85 312
rect 83 311 84 312
rect 82 311 83 312
rect 81 311 82 312
rect 80 311 81 312
rect 79 311 80 312
rect 78 311 79 312
rect 77 311 78 312
rect 76 311 77 312
rect 75 311 76 312
rect 74 311 75 312
rect 73 311 74 312
rect 72 311 73 312
rect 71 311 72 312
rect 56 311 57 312
rect 55 311 56 312
rect 54 311 55 312
rect 53 311 54 312
rect 52 311 53 312
rect 51 311 52 312
rect 50 311 51 312
rect 49 311 50 312
rect 48 311 49 312
rect 47 311 48 312
rect 46 311 47 312
rect 45 311 46 312
rect 44 311 45 312
rect 43 311 44 312
rect 42 311 43 312
rect 41 311 42 312
rect 40 311 41 312
rect 39 311 40 312
rect 38 311 39 312
rect 37 311 38 312
rect 36 311 37 312
rect 35 311 36 312
rect 34 311 35 312
rect 33 311 34 312
rect 32 311 33 312
rect 31 311 32 312
rect 30 311 31 312
rect 29 311 30 312
rect 28 311 29 312
rect 27 311 28 312
rect 26 311 27 312
rect 25 311 26 312
rect 24 311 25 312
rect 23 311 24 312
rect 22 311 23 312
rect 21 311 22 312
rect 20 311 21 312
rect 19 311 20 312
rect 18 311 19 312
rect 85 312 86 313
rect 84 312 85 313
rect 83 312 84 313
rect 82 312 83 313
rect 81 312 82 313
rect 80 312 81 313
rect 79 312 80 313
rect 78 312 79 313
rect 77 312 78 313
rect 76 312 77 313
rect 75 312 76 313
rect 74 312 75 313
rect 73 312 74 313
rect 72 312 73 313
rect 71 312 72 313
rect 56 312 57 313
rect 55 312 56 313
rect 54 312 55 313
rect 53 312 54 313
rect 52 312 53 313
rect 51 312 52 313
rect 50 312 51 313
rect 49 312 50 313
rect 48 312 49 313
rect 47 312 48 313
rect 46 312 47 313
rect 45 312 46 313
rect 44 312 45 313
rect 43 312 44 313
rect 42 312 43 313
rect 41 312 42 313
rect 40 312 41 313
rect 39 312 40 313
rect 38 312 39 313
rect 37 312 38 313
rect 36 312 37 313
rect 35 312 36 313
rect 34 312 35 313
rect 33 312 34 313
rect 32 312 33 313
rect 31 312 32 313
rect 30 312 31 313
rect 29 312 30 313
rect 28 312 29 313
rect 27 312 28 313
rect 26 312 27 313
rect 25 312 26 313
rect 24 312 25 313
rect 23 312 24 313
rect 22 312 23 313
rect 21 312 22 313
rect 20 312 21 313
rect 19 312 20 313
rect 18 312 19 313
rect 85 313 86 314
rect 84 313 85 314
rect 83 313 84 314
rect 82 313 83 314
rect 81 313 82 314
rect 80 313 81 314
rect 79 313 80 314
rect 78 313 79 314
rect 77 313 78 314
rect 76 313 77 314
rect 75 313 76 314
rect 74 313 75 314
rect 73 313 74 314
rect 72 313 73 314
rect 71 313 72 314
rect 56 313 57 314
rect 55 313 56 314
rect 54 313 55 314
rect 53 313 54 314
rect 52 313 53 314
rect 51 313 52 314
rect 50 313 51 314
rect 49 313 50 314
rect 48 313 49 314
rect 47 313 48 314
rect 46 313 47 314
rect 45 313 46 314
rect 44 313 45 314
rect 43 313 44 314
rect 42 313 43 314
rect 41 313 42 314
rect 40 313 41 314
rect 39 313 40 314
rect 38 313 39 314
rect 37 313 38 314
rect 36 313 37 314
rect 35 313 36 314
rect 34 313 35 314
rect 33 313 34 314
rect 32 313 33 314
rect 31 313 32 314
rect 30 313 31 314
rect 29 313 30 314
rect 28 313 29 314
rect 27 313 28 314
rect 26 313 27 314
rect 25 313 26 314
rect 24 313 25 314
rect 23 313 24 314
rect 22 313 23 314
rect 21 313 22 314
rect 20 313 21 314
rect 19 313 20 314
rect 18 313 19 314
rect 85 314 86 315
rect 84 314 85 315
rect 83 314 84 315
rect 82 314 83 315
rect 81 314 82 315
rect 80 314 81 315
rect 79 314 80 315
rect 78 314 79 315
rect 77 314 78 315
rect 76 314 77 315
rect 75 314 76 315
rect 74 314 75 315
rect 73 314 74 315
rect 72 314 73 315
rect 71 314 72 315
rect 56 314 57 315
rect 55 314 56 315
rect 54 314 55 315
rect 53 314 54 315
rect 52 314 53 315
rect 51 314 52 315
rect 50 314 51 315
rect 49 314 50 315
rect 48 314 49 315
rect 47 314 48 315
rect 46 314 47 315
rect 45 314 46 315
rect 44 314 45 315
rect 43 314 44 315
rect 42 314 43 315
rect 41 314 42 315
rect 40 314 41 315
rect 39 314 40 315
rect 38 314 39 315
rect 37 314 38 315
rect 36 314 37 315
rect 35 314 36 315
rect 34 314 35 315
rect 33 314 34 315
rect 32 314 33 315
rect 31 314 32 315
rect 30 314 31 315
rect 29 314 30 315
rect 28 314 29 315
rect 27 314 28 315
rect 26 314 27 315
rect 25 314 26 315
rect 24 314 25 315
rect 23 314 24 315
rect 22 314 23 315
rect 21 314 22 315
rect 20 314 21 315
rect 19 314 20 315
rect 18 314 19 315
rect 140 315 141 316
rect 139 315 140 316
rect 138 315 139 316
rect 137 315 138 316
rect 136 315 137 316
rect 135 315 136 316
rect 134 315 135 316
rect 85 315 86 316
rect 84 315 85 316
rect 83 315 84 316
rect 82 315 83 316
rect 81 315 82 316
rect 80 315 81 316
rect 79 315 80 316
rect 78 315 79 316
rect 77 315 78 316
rect 76 315 77 316
rect 75 315 76 316
rect 74 315 75 316
rect 73 315 74 316
rect 72 315 73 316
rect 71 315 72 316
rect 56 315 57 316
rect 55 315 56 316
rect 54 315 55 316
rect 53 315 54 316
rect 52 315 53 316
rect 51 315 52 316
rect 50 315 51 316
rect 49 315 50 316
rect 48 315 49 316
rect 47 315 48 316
rect 46 315 47 316
rect 45 315 46 316
rect 44 315 45 316
rect 43 315 44 316
rect 42 315 43 316
rect 41 315 42 316
rect 40 315 41 316
rect 39 315 40 316
rect 38 315 39 316
rect 37 315 38 316
rect 36 315 37 316
rect 35 315 36 316
rect 34 315 35 316
rect 33 315 34 316
rect 32 315 33 316
rect 31 315 32 316
rect 30 315 31 316
rect 29 315 30 316
rect 28 315 29 316
rect 27 315 28 316
rect 26 315 27 316
rect 25 315 26 316
rect 24 315 25 316
rect 23 315 24 316
rect 22 315 23 316
rect 21 315 22 316
rect 20 315 21 316
rect 19 315 20 316
rect 18 315 19 316
rect 142 316 143 317
rect 141 316 142 317
rect 140 316 141 317
rect 139 316 140 317
rect 138 316 139 317
rect 137 316 138 317
rect 136 316 137 317
rect 135 316 136 317
rect 134 316 135 317
rect 133 316 134 317
rect 132 316 133 317
rect 85 316 86 317
rect 84 316 85 317
rect 83 316 84 317
rect 82 316 83 317
rect 81 316 82 317
rect 80 316 81 317
rect 79 316 80 317
rect 78 316 79 317
rect 77 316 78 317
rect 76 316 77 317
rect 75 316 76 317
rect 74 316 75 317
rect 73 316 74 317
rect 72 316 73 317
rect 71 316 72 317
rect 56 316 57 317
rect 55 316 56 317
rect 54 316 55 317
rect 53 316 54 317
rect 52 316 53 317
rect 51 316 52 317
rect 50 316 51 317
rect 49 316 50 317
rect 48 316 49 317
rect 47 316 48 317
rect 46 316 47 317
rect 45 316 46 317
rect 44 316 45 317
rect 43 316 44 317
rect 42 316 43 317
rect 41 316 42 317
rect 40 316 41 317
rect 39 316 40 317
rect 38 316 39 317
rect 37 316 38 317
rect 36 316 37 317
rect 35 316 36 317
rect 34 316 35 317
rect 33 316 34 317
rect 32 316 33 317
rect 31 316 32 317
rect 30 316 31 317
rect 29 316 30 317
rect 28 316 29 317
rect 27 316 28 317
rect 26 316 27 317
rect 25 316 26 317
rect 24 316 25 317
rect 23 316 24 317
rect 22 316 23 317
rect 21 316 22 317
rect 20 316 21 317
rect 19 316 20 317
rect 18 316 19 317
rect 143 317 144 318
rect 142 317 143 318
rect 141 317 142 318
rect 140 317 141 318
rect 139 317 140 318
rect 138 317 139 318
rect 137 317 138 318
rect 136 317 137 318
rect 135 317 136 318
rect 134 317 135 318
rect 133 317 134 318
rect 132 317 133 318
rect 131 317 132 318
rect 85 317 86 318
rect 84 317 85 318
rect 83 317 84 318
rect 82 317 83 318
rect 81 317 82 318
rect 80 317 81 318
rect 79 317 80 318
rect 78 317 79 318
rect 77 317 78 318
rect 76 317 77 318
rect 75 317 76 318
rect 74 317 75 318
rect 73 317 74 318
rect 72 317 73 318
rect 71 317 72 318
rect 70 317 71 318
rect 57 317 58 318
rect 56 317 57 318
rect 55 317 56 318
rect 54 317 55 318
rect 53 317 54 318
rect 52 317 53 318
rect 51 317 52 318
rect 50 317 51 318
rect 49 317 50 318
rect 48 317 49 318
rect 47 317 48 318
rect 46 317 47 318
rect 45 317 46 318
rect 44 317 45 318
rect 43 317 44 318
rect 33 317 34 318
rect 32 317 33 318
rect 31 317 32 318
rect 30 317 31 318
rect 29 317 30 318
rect 28 317 29 318
rect 27 317 28 318
rect 26 317 27 318
rect 25 317 26 318
rect 24 317 25 318
rect 23 317 24 318
rect 22 317 23 318
rect 21 317 22 318
rect 20 317 21 318
rect 19 317 20 318
rect 18 317 19 318
rect 144 318 145 319
rect 143 318 144 319
rect 142 318 143 319
rect 141 318 142 319
rect 140 318 141 319
rect 139 318 140 319
rect 138 318 139 319
rect 137 318 138 319
rect 136 318 137 319
rect 135 318 136 319
rect 134 318 135 319
rect 133 318 134 319
rect 132 318 133 319
rect 131 318 132 319
rect 130 318 131 319
rect 85 318 86 319
rect 84 318 85 319
rect 83 318 84 319
rect 82 318 83 319
rect 81 318 82 319
rect 80 318 81 319
rect 79 318 80 319
rect 78 318 79 319
rect 77 318 78 319
rect 76 318 77 319
rect 75 318 76 319
rect 74 318 75 319
rect 73 318 74 319
rect 72 318 73 319
rect 71 318 72 319
rect 70 318 71 319
rect 57 318 58 319
rect 56 318 57 319
rect 55 318 56 319
rect 54 318 55 319
rect 53 318 54 319
rect 52 318 53 319
rect 51 318 52 319
rect 50 318 51 319
rect 49 318 50 319
rect 48 318 49 319
rect 47 318 48 319
rect 46 318 47 319
rect 45 318 46 319
rect 44 318 45 319
rect 43 318 44 319
rect 33 318 34 319
rect 32 318 33 319
rect 31 318 32 319
rect 30 318 31 319
rect 29 318 30 319
rect 28 318 29 319
rect 27 318 28 319
rect 26 318 27 319
rect 25 318 26 319
rect 24 318 25 319
rect 23 318 24 319
rect 22 318 23 319
rect 21 318 22 319
rect 20 318 21 319
rect 19 318 20 319
rect 18 318 19 319
rect 145 319 146 320
rect 144 319 145 320
rect 143 319 144 320
rect 142 319 143 320
rect 141 319 142 320
rect 140 319 141 320
rect 139 319 140 320
rect 138 319 139 320
rect 137 319 138 320
rect 136 319 137 320
rect 135 319 136 320
rect 134 319 135 320
rect 133 319 134 320
rect 132 319 133 320
rect 131 319 132 320
rect 130 319 131 320
rect 129 319 130 320
rect 85 319 86 320
rect 84 319 85 320
rect 83 319 84 320
rect 82 319 83 320
rect 81 319 82 320
rect 80 319 81 320
rect 79 319 80 320
rect 78 319 79 320
rect 77 319 78 320
rect 76 319 77 320
rect 75 319 76 320
rect 74 319 75 320
rect 73 319 74 320
rect 72 319 73 320
rect 71 319 72 320
rect 70 319 71 320
rect 57 319 58 320
rect 56 319 57 320
rect 55 319 56 320
rect 54 319 55 320
rect 53 319 54 320
rect 52 319 53 320
rect 51 319 52 320
rect 50 319 51 320
rect 49 319 50 320
rect 48 319 49 320
rect 47 319 48 320
rect 46 319 47 320
rect 45 319 46 320
rect 44 319 45 320
rect 43 319 44 320
rect 33 319 34 320
rect 32 319 33 320
rect 31 319 32 320
rect 30 319 31 320
rect 29 319 30 320
rect 28 319 29 320
rect 27 319 28 320
rect 26 319 27 320
rect 25 319 26 320
rect 24 319 25 320
rect 23 319 24 320
rect 22 319 23 320
rect 21 319 22 320
rect 20 319 21 320
rect 19 319 20 320
rect 18 319 19 320
rect 145 320 146 321
rect 144 320 145 321
rect 143 320 144 321
rect 142 320 143 321
rect 141 320 142 321
rect 140 320 141 321
rect 139 320 140 321
rect 138 320 139 321
rect 137 320 138 321
rect 136 320 137 321
rect 135 320 136 321
rect 134 320 135 321
rect 133 320 134 321
rect 132 320 133 321
rect 131 320 132 321
rect 130 320 131 321
rect 129 320 130 321
rect 85 320 86 321
rect 84 320 85 321
rect 83 320 84 321
rect 82 320 83 321
rect 81 320 82 321
rect 80 320 81 321
rect 79 320 80 321
rect 78 320 79 321
rect 77 320 78 321
rect 76 320 77 321
rect 75 320 76 321
rect 74 320 75 321
rect 73 320 74 321
rect 72 320 73 321
rect 71 320 72 321
rect 70 320 71 321
rect 69 320 70 321
rect 58 320 59 321
rect 57 320 58 321
rect 56 320 57 321
rect 55 320 56 321
rect 54 320 55 321
rect 53 320 54 321
rect 52 320 53 321
rect 51 320 52 321
rect 50 320 51 321
rect 49 320 50 321
rect 48 320 49 321
rect 47 320 48 321
rect 46 320 47 321
rect 45 320 46 321
rect 44 320 45 321
rect 43 320 44 321
rect 33 320 34 321
rect 32 320 33 321
rect 31 320 32 321
rect 30 320 31 321
rect 29 320 30 321
rect 28 320 29 321
rect 27 320 28 321
rect 26 320 27 321
rect 25 320 26 321
rect 24 320 25 321
rect 23 320 24 321
rect 22 320 23 321
rect 21 320 22 321
rect 20 320 21 321
rect 19 320 20 321
rect 18 320 19 321
rect 146 321 147 322
rect 145 321 146 322
rect 144 321 145 322
rect 143 321 144 322
rect 142 321 143 322
rect 141 321 142 322
rect 133 321 134 322
rect 132 321 133 322
rect 131 321 132 322
rect 130 321 131 322
rect 129 321 130 322
rect 128 321 129 322
rect 85 321 86 322
rect 84 321 85 322
rect 83 321 84 322
rect 82 321 83 322
rect 81 321 82 322
rect 80 321 81 322
rect 79 321 80 322
rect 78 321 79 322
rect 77 321 78 322
rect 76 321 77 322
rect 75 321 76 322
rect 74 321 75 322
rect 73 321 74 322
rect 72 321 73 322
rect 71 321 72 322
rect 70 321 71 322
rect 69 321 70 322
rect 68 321 69 322
rect 59 321 60 322
rect 58 321 59 322
rect 57 321 58 322
rect 56 321 57 322
rect 55 321 56 322
rect 54 321 55 322
rect 53 321 54 322
rect 52 321 53 322
rect 51 321 52 322
rect 50 321 51 322
rect 49 321 50 322
rect 48 321 49 322
rect 47 321 48 322
rect 46 321 47 322
rect 45 321 46 322
rect 44 321 45 322
rect 43 321 44 322
rect 33 321 34 322
rect 32 321 33 322
rect 31 321 32 322
rect 30 321 31 322
rect 29 321 30 322
rect 28 321 29 322
rect 27 321 28 322
rect 26 321 27 322
rect 25 321 26 322
rect 24 321 25 322
rect 23 321 24 322
rect 22 321 23 322
rect 21 321 22 322
rect 20 321 21 322
rect 19 321 20 322
rect 18 321 19 322
rect 146 322 147 323
rect 145 322 146 323
rect 144 322 145 323
rect 143 322 144 323
rect 142 322 143 323
rect 132 322 133 323
rect 131 322 132 323
rect 130 322 131 323
rect 129 322 130 323
rect 128 322 129 323
rect 84 322 85 323
rect 83 322 84 323
rect 82 322 83 323
rect 81 322 82 323
rect 80 322 81 323
rect 79 322 80 323
rect 78 322 79 323
rect 77 322 78 323
rect 76 322 77 323
rect 75 322 76 323
rect 74 322 75 323
rect 73 322 74 323
rect 72 322 73 323
rect 71 322 72 323
rect 70 322 71 323
rect 69 322 70 323
rect 68 322 69 323
rect 67 322 68 323
rect 60 322 61 323
rect 59 322 60 323
rect 58 322 59 323
rect 57 322 58 323
rect 56 322 57 323
rect 55 322 56 323
rect 54 322 55 323
rect 53 322 54 323
rect 52 322 53 323
rect 51 322 52 323
rect 50 322 51 323
rect 49 322 50 323
rect 48 322 49 323
rect 47 322 48 323
rect 46 322 47 323
rect 45 322 46 323
rect 44 322 45 323
rect 43 322 44 323
rect 33 322 34 323
rect 32 322 33 323
rect 31 322 32 323
rect 30 322 31 323
rect 29 322 30 323
rect 28 322 29 323
rect 27 322 28 323
rect 26 322 27 323
rect 25 322 26 323
rect 24 322 25 323
rect 23 322 24 323
rect 22 322 23 323
rect 21 322 22 323
rect 20 322 21 323
rect 19 322 20 323
rect 18 322 19 323
rect 146 323 147 324
rect 145 323 146 324
rect 144 323 145 324
rect 143 323 144 324
rect 142 323 143 324
rect 132 323 133 324
rect 131 323 132 324
rect 130 323 131 324
rect 129 323 130 324
rect 128 323 129 324
rect 84 323 85 324
rect 83 323 84 324
rect 82 323 83 324
rect 81 323 82 324
rect 80 323 81 324
rect 79 323 80 324
rect 78 323 79 324
rect 77 323 78 324
rect 76 323 77 324
rect 75 323 76 324
rect 74 323 75 324
rect 73 323 74 324
rect 72 323 73 324
rect 71 323 72 324
rect 70 323 71 324
rect 69 323 70 324
rect 68 323 69 324
rect 67 323 68 324
rect 66 323 67 324
rect 65 323 66 324
rect 64 323 65 324
rect 63 323 64 324
rect 62 323 63 324
rect 61 323 62 324
rect 60 323 61 324
rect 59 323 60 324
rect 58 323 59 324
rect 57 323 58 324
rect 56 323 57 324
rect 55 323 56 324
rect 54 323 55 324
rect 53 323 54 324
rect 52 323 53 324
rect 51 323 52 324
rect 50 323 51 324
rect 49 323 50 324
rect 48 323 49 324
rect 47 323 48 324
rect 46 323 47 324
rect 45 323 46 324
rect 44 323 45 324
rect 43 323 44 324
rect 33 323 34 324
rect 32 323 33 324
rect 31 323 32 324
rect 30 323 31 324
rect 29 323 30 324
rect 28 323 29 324
rect 27 323 28 324
rect 26 323 27 324
rect 25 323 26 324
rect 24 323 25 324
rect 23 323 24 324
rect 22 323 23 324
rect 21 323 22 324
rect 20 323 21 324
rect 19 323 20 324
rect 18 323 19 324
rect 146 324 147 325
rect 145 324 146 325
rect 144 324 145 325
rect 143 324 144 325
rect 131 324 132 325
rect 130 324 131 325
rect 129 324 130 325
rect 128 324 129 325
rect 84 324 85 325
rect 83 324 84 325
rect 82 324 83 325
rect 81 324 82 325
rect 80 324 81 325
rect 79 324 80 325
rect 78 324 79 325
rect 77 324 78 325
rect 76 324 77 325
rect 75 324 76 325
rect 74 324 75 325
rect 73 324 74 325
rect 72 324 73 325
rect 71 324 72 325
rect 70 324 71 325
rect 69 324 70 325
rect 68 324 69 325
rect 67 324 68 325
rect 66 324 67 325
rect 65 324 66 325
rect 64 324 65 325
rect 63 324 64 325
rect 62 324 63 325
rect 61 324 62 325
rect 60 324 61 325
rect 59 324 60 325
rect 58 324 59 325
rect 57 324 58 325
rect 56 324 57 325
rect 55 324 56 325
rect 54 324 55 325
rect 53 324 54 325
rect 52 324 53 325
rect 51 324 52 325
rect 50 324 51 325
rect 49 324 50 325
rect 48 324 49 325
rect 47 324 48 325
rect 46 324 47 325
rect 45 324 46 325
rect 44 324 45 325
rect 43 324 44 325
rect 33 324 34 325
rect 32 324 33 325
rect 31 324 32 325
rect 30 324 31 325
rect 29 324 30 325
rect 28 324 29 325
rect 27 324 28 325
rect 26 324 27 325
rect 25 324 26 325
rect 24 324 25 325
rect 23 324 24 325
rect 22 324 23 325
rect 21 324 22 325
rect 20 324 21 325
rect 19 324 20 325
rect 18 324 19 325
rect 146 325 147 326
rect 145 325 146 326
rect 144 325 145 326
rect 143 325 144 326
rect 131 325 132 326
rect 130 325 131 326
rect 129 325 130 326
rect 128 325 129 326
rect 84 325 85 326
rect 83 325 84 326
rect 82 325 83 326
rect 81 325 82 326
rect 80 325 81 326
rect 79 325 80 326
rect 78 325 79 326
rect 77 325 78 326
rect 76 325 77 326
rect 75 325 76 326
rect 74 325 75 326
rect 73 325 74 326
rect 72 325 73 326
rect 71 325 72 326
rect 70 325 71 326
rect 69 325 70 326
rect 68 325 69 326
rect 67 325 68 326
rect 66 325 67 326
rect 65 325 66 326
rect 64 325 65 326
rect 63 325 64 326
rect 62 325 63 326
rect 61 325 62 326
rect 60 325 61 326
rect 59 325 60 326
rect 58 325 59 326
rect 57 325 58 326
rect 56 325 57 326
rect 55 325 56 326
rect 54 325 55 326
rect 53 325 54 326
rect 52 325 53 326
rect 51 325 52 326
rect 50 325 51 326
rect 49 325 50 326
rect 48 325 49 326
rect 47 325 48 326
rect 46 325 47 326
rect 45 325 46 326
rect 44 325 45 326
rect 43 325 44 326
rect 33 325 34 326
rect 32 325 33 326
rect 31 325 32 326
rect 30 325 31 326
rect 29 325 30 326
rect 28 325 29 326
rect 27 325 28 326
rect 26 325 27 326
rect 25 325 26 326
rect 24 325 25 326
rect 23 325 24 326
rect 22 325 23 326
rect 21 325 22 326
rect 20 325 21 326
rect 19 325 20 326
rect 18 325 19 326
rect 146 326 147 327
rect 145 326 146 327
rect 144 326 145 327
rect 143 326 144 327
rect 142 326 143 327
rect 132 326 133 327
rect 131 326 132 327
rect 130 326 131 327
rect 129 326 130 327
rect 128 326 129 327
rect 83 326 84 327
rect 82 326 83 327
rect 81 326 82 327
rect 80 326 81 327
rect 79 326 80 327
rect 78 326 79 327
rect 77 326 78 327
rect 76 326 77 327
rect 75 326 76 327
rect 74 326 75 327
rect 73 326 74 327
rect 72 326 73 327
rect 71 326 72 327
rect 70 326 71 327
rect 69 326 70 327
rect 68 326 69 327
rect 67 326 68 327
rect 66 326 67 327
rect 65 326 66 327
rect 64 326 65 327
rect 63 326 64 327
rect 62 326 63 327
rect 61 326 62 327
rect 60 326 61 327
rect 59 326 60 327
rect 58 326 59 327
rect 57 326 58 327
rect 56 326 57 327
rect 55 326 56 327
rect 54 326 55 327
rect 53 326 54 327
rect 52 326 53 327
rect 51 326 52 327
rect 50 326 51 327
rect 49 326 50 327
rect 48 326 49 327
rect 47 326 48 327
rect 46 326 47 327
rect 45 326 46 327
rect 44 326 45 327
rect 43 326 44 327
rect 33 326 34 327
rect 32 326 33 327
rect 31 326 32 327
rect 30 326 31 327
rect 29 326 30 327
rect 28 326 29 327
rect 27 326 28 327
rect 26 326 27 327
rect 25 326 26 327
rect 24 326 25 327
rect 23 326 24 327
rect 22 326 23 327
rect 21 326 22 327
rect 20 326 21 327
rect 19 326 20 327
rect 18 326 19 327
rect 146 327 147 328
rect 145 327 146 328
rect 144 327 145 328
rect 143 327 144 328
rect 142 327 143 328
rect 132 327 133 328
rect 131 327 132 328
rect 130 327 131 328
rect 129 327 130 328
rect 128 327 129 328
rect 83 327 84 328
rect 82 327 83 328
rect 81 327 82 328
rect 80 327 81 328
rect 79 327 80 328
rect 78 327 79 328
rect 77 327 78 328
rect 76 327 77 328
rect 75 327 76 328
rect 74 327 75 328
rect 73 327 74 328
rect 72 327 73 328
rect 71 327 72 328
rect 70 327 71 328
rect 69 327 70 328
rect 68 327 69 328
rect 67 327 68 328
rect 66 327 67 328
rect 65 327 66 328
rect 64 327 65 328
rect 63 327 64 328
rect 62 327 63 328
rect 61 327 62 328
rect 60 327 61 328
rect 59 327 60 328
rect 58 327 59 328
rect 57 327 58 328
rect 56 327 57 328
rect 55 327 56 328
rect 54 327 55 328
rect 53 327 54 328
rect 52 327 53 328
rect 51 327 52 328
rect 50 327 51 328
rect 49 327 50 328
rect 48 327 49 328
rect 47 327 48 328
rect 46 327 47 328
rect 45 327 46 328
rect 44 327 45 328
rect 33 327 34 328
rect 32 327 33 328
rect 31 327 32 328
rect 30 327 31 328
rect 29 327 30 328
rect 28 327 29 328
rect 27 327 28 328
rect 26 327 27 328
rect 25 327 26 328
rect 24 327 25 328
rect 23 327 24 328
rect 22 327 23 328
rect 21 327 22 328
rect 20 327 21 328
rect 19 327 20 328
rect 18 327 19 328
rect 146 328 147 329
rect 145 328 146 329
rect 144 328 145 329
rect 143 328 144 329
rect 142 328 143 329
rect 141 328 142 329
rect 133 328 134 329
rect 132 328 133 329
rect 131 328 132 329
rect 130 328 131 329
rect 129 328 130 329
rect 128 328 129 329
rect 83 328 84 329
rect 82 328 83 329
rect 81 328 82 329
rect 80 328 81 329
rect 79 328 80 329
rect 78 328 79 329
rect 77 328 78 329
rect 76 328 77 329
rect 75 328 76 329
rect 74 328 75 329
rect 73 328 74 329
rect 72 328 73 329
rect 71 328 72 329
rect 70 328 71 329
rect 69 328 70 329
rect 68 328 69 329
rect 67 328 68 329
rect 66 328 67 329
rect 65 328 66 329
rect 64 328 65 329
rect 63 328 64 329
rect 62 328 63 329
rect 61 328 62 329
rect 60 328 61 329
rect 59 328 60 329
rect 58 328 59 329
rect 57 328 58 329
rect 56 328 57 329
rect 55 328 56 329
rect 54 328 55 329
rect 53 328 54 329
rect 52 328 53 329
rect 51 328 52 329
rect 50 328 51 329
rect 49 328 50 329
rect 48 328 49 329
rect 47 328 48 329
rect 46 328 47 329
rect 45 328 46 329
rect 44 328 45 329
rect 33 328 34 329
rect 32 328 33 329
rect 31 328 32 329
rect 30 328 31 329
rect 29 328 30 329
rect 28 328 29 329
rect 27 328 28 329
rect 26 328 27 329
rect 25 328 26 329
rect 24 328 25 329
rect 23 328 24 329
rect 22 328 23 329
rect 21 328 22 329
rect 20 328 21 329
rect 19 328 20 329
rect 18 328 19 329
rect 145 329 146 330
rect 144 329 145 330
rect 143 329 144 330
rect 142 329 143 330
rect 141 329 142 330
rect 140 329 141 330
rect 139 329 140 330
rect 138 329 139 330
rect 137 329 138 330
rect 136 329 137 330
rect 135 329 136 330
rect 134 329 135 330
rect 133 329 134 330
rect 132 329 133 330
rect 131 329 132 330
rect 130 329 131 330
rect 129 329 130 330
rect 82 329 83 330
rect 81 329 82 330
rect 80 329 81 330
rect 79 329 80 330
rect 78 329 79 330
rect 77 329 78 330
rect 76 329 77 330
rect 75 329 76 330
rect 74 329 75 330
rect 73 329 74 330
rect 72 329 73 330
rect 71 329 72 330
rect 70 329 71 330
rect 69 329 70 330
rect 68 329 69 330
rect 67 329 68 330
rect 66 329 67 330
rect 65 329 66 330
rect 64 329 65 330
rect 63 329 64 330
rect 62 329 63 330
rect 61 329 62 330
rect 60 329 61 330
rect 59 329 60 330
rect 58 329 59 330
rect 57 329 58 330
rect 56 329 57 330
rect 55 329 56 330
rect 54 329 55 330
rect 53 329 54 330
rect 52 329 53 330
rect 51 329 52 330
rect 50 329 51 330
rect 49 329 50 330
rect 48 329 49 330
rect 47 329 48 330
rect 46 329 47 330
rect 45 329 46 330
rect 44 329 45 330
rect 33 329 34 330
rect 32 329 33 330
rect 31 329 32 330
rect 30 329 31 330
rect 29 329 30 330
rect 28 329 29 330
rect 27 329 28 330
rect 26 329 27 330
rect 25 329 26 330
rect 24 329 25 330
rect 23 329 24 330
rect 22 329 23 330
rect 21 329 22 330
rect 20 329 21 330
rect 19 329 20 330
rect 18 329 19 330
rect 145 330 146 331
rect 144 330 145 331
rect 143 330 144 331
rect 142 330 143 331
rect 141 330 142 331
rect 140 330 141 331
rect 139 330 140 331
rect 138 330 139 331
rect 137 330 138 331
rect 136 330 137 331
rect 135 330 136 331
rect 134 330 135 331
rect 133 330 134 331
rect 132 330 133 331
rect 131 330 132 331
rect 130 330 131 331
rect 129 330 130 331
rect 82 330 83 331
rect 81 330 82 331
rect 80 330 81 331
rect 79 330 80 331
rect 78 330 79 331
rect 77 330 78 331
rect 76 330 77 331
rect 75 330 76 331
rect 74 330 75 331
rect 73 330 74 331
rect 72 330 73 331
rect 71 330 72 331
rect 70 330 71 331
rect 69 330 70 331
rect 68 330 69 331
rect 67 330 68 331
rect 66 330 67 331
rect 65 330 66 331
rect 64 330 65 331
rect 63 330 64 331
rect 62 330 63 331
rect 61 330 62 331
rect 60 330 61 331
rect 59 330 60 331
rect 58 330 59 331
rect 57 330 58 331
rect 56 330 57 331
rect 55 330 56 331
rect 54 330 55 331
rect 53 330 54 331
rect 52 330 53 331
rect 51 330 52 331
rect 50 330 51 331
rect 49 330 50 331
rect 48 330 49 331
rect 47 330 48 331
rect 46 330 47 331
rect 45 330 46 331
rect 44 330 45 331
rect 33 330 34 331
rect 32 330 33 331
rect 31 330 32 331
rect 30 330 31 331
rect 29 330 30 331
rect 28 330 29 331
rect 27 330 28 331
rect 26 330 27 331
rect 25 330 26 331
rect 24 330 25 331
rect 23 330 24 331
rect 22 330 23 331
rect 21 330 22 331
rect 20 330 21 331
rect 19 330 20 331
rect 18 330 19 331
rect 144 331 145 332
rect 143 331 144 332
rect 142 331 143 332
rect 141 331 142 332
rect 140 331 141 332
rect 139 331 140 332
rect 138 331 139 332
rect 137 331 138 332
rect 136 331 137 332
rect 135 331 136 332
rect 134 331 135 332
rect 133 331 134 332
rect 132 331 133 332
rect 131 331 132 332
rect 130 331 131 332
rect 81 331 82 332
rect 80 331 81 332
rect 79 331 80 332
rect 78 331 79 332
rect 77 331 78 332
rect 76 331 77 332
rect 75 331 76 332
rect 74 331 75 332
rect 73 331 74 332
rect 72 331 73 332
rect 71 331 72 332
rect 70 331 71 332
rect 69 331 70 332
rect 68 331 69 332
rect 67 331 68 332
rect 66 331 67 332
rect 65 331 66 332
rect 64 331 65 332
rect 63 331 64 332
rect 62 331 63 332
rect 61 331 62 332
rect 60 331 61 332
rect 59 331 60 332
rect 58 331 59 332
rect 57 331 58 332
rect 56 331 57 332
rect 55 331 56 332
rect 54 331 55 332
rect 53 331 54 332
rect 52 331 53 332
rect 51 331 52 332
rect 50 331 51 332
rect 49 331 50 332
rect 48 331 49 332
rect 47 331 48 332
rect 46 331 47 332
rect 45 331 46 332
rect 33 331 34 332
rect 32 331 33 332
rect 31 331 32 332
rect 30 331 31 332
rect 29 331 30 332
rect 28 331 29 332
rect 27 331 28 332
rect 26 331 27 332
rect 25 331 26 332
rect 24 331 25 332
rect 23 331 24 332
rect 22 331 23 332
rect 21 331 22 332
rect 20 331 21 332
rect 19 331 20 332
rect 18 331 19 332
rect 143 332 144 333
rect 142 332 143 333
rect 141 332 142 333
rect 140 332 141 333
rect 139 332 140 333
rect 138 332 139 333
rect 137 332 138 333
rect 136 332 137 333
rect 135 332 136 333
rect 134 332 135 333
rect 133 332 134 333
rect 132 332 133 333
rect 131 332 132 333
rect 81 332 82 333
rect 80 332 81 333
rect 79 332 80 333
rect 78 332 79 333
rect 77 332 78 333
rect 76 332 77 333
rect 75 332 76 333
rect 74 332 75 333
rect 73 332 74 333
rect 72 332 73 333
rect 71 332 72 333
rect 70 332 71 333
rect 69 332 70 333
rect 68 332 69 333
rect 67 332 68 333
rect 66 332 67 333
rect 65 332 66 333
rect 64 332 65 333
rect 63 332 64 333
rect 62 332 63 333
rect 61 332 62 333
rect 60 332 61 333
rect 59 332 60 333
rect 58 332 59 333
rect 57 332 58 333
rect 56 332 57 333
rect 55 332 56 333
rect 54 332 55 333
rect 53 332 54 333
rect 52 332 53 333
rect 51 332 52 333
rect 50 332 51 333
rect 49 332 50 333
rect 48 332 49 333
rect 47 332 48 333
rect 46 332 47 333
rect 45 332 46 333
rect 33 332 34 333
rect 32 332 33 333
rect 31 332 32 333
rect 30 332 31 333
rect 29 332 30 333
rect 28 332 29 333
rect 27 332 28 333
rect 26 332 27 333
rect 25 332 26 333
rect 24 332 25 333
rect 23 332 24 333
rect 22 332 23 333
rect 21 332 22 333
rect 20 332 21 333
rect 19 332 20 333
rect 18 332 19 333
rect 142 333 143 334
rect 141 333 142 334
rect 140 333 141 334
rect 139 333 140 334
rect 138 333 139 334
rect 137 333 138 334
rect 136 333 137 334
rect 135 333 136 334
rect 134 333 135 334
rect 133 333 134 334
rect 132 333 133 334
rect 80 333 81 334
rect 79 333 80 334
rect 78 333 79 334
rect 77 333 78 334
rect 76 333 77 334
rect 75 333 76 334
rect 74 333 75 334
rect 73 333 74 334
rect 72 333 73 334
rect 71 333 72 334
rect 70 333 71 334
rect 69 333 70 334
rect 68 333 69 334
rect 67 333 68 334
rect 66 333 67 334
rect 65 333 66 334
rect 64 333 65 334
rect 63 333 64 334
rect 62 333 63 334
rect 61 333 62 334
rect 60 333 61 334
rect 59 333 60 334
rect 58 333 59 334
rect 57 333 58 334
rect 56 333 57 334
rect 55 333 56 334
rect 54 333 55 334
rect 53 333 54 334
rect 52 333 53 334
rect 51 333 52 334
rect 50 333 51 334
rect 49 333 50 334
rect 48 333 49 334
rect 47 333 48 334
rect 46 333 47 334
rect 33 333 34 334
rect 32 333 33 334
rect 31 333 32 334
rect 30 333 31 334
rect 29 333 30 334
rect 28 333 29 334
rect 27 333 28 334
rect 26 333 27 334
rect 25 333 26 334
rect 24 333 25 334
rect 23 333 24 334
rect 22 333 23 334
rect 21 333 22 334
rect 20 333 21 334
rect 19 333 20 334
rect 18 333 19 334
rect 139 334 140 335
rect 138 334 139 335
rect 137 334 138 335
rect 136 334 137 335
rect 135 334 136 335
rect 134 334 135 335
rect 79 334 80 335
rect 78 334 79 335
rect 77 334 78 335
rect 76 334 77 335
rect 75 334 76 335
rect 74 334 75 335
rect 73 334 74 335
rect 72 334 73 335
rect 71 334 72 335
rect 70 334 71 335
rect 69 334 70 335
rect 68 334 69 335
rect 67 334 68 335
rect 66 334 67 335
rect 65 334 66 335
rect 64 334 65 335
rect 63 334 64 335
rect 62 334 63 335
rect 61 334 62 335
rect 60 334 61 335
rect 59 334 60 335
rect 58 334 59 335
rect 57 334 58 335
rect 56 334 57 335
rect 55 334 56 335
rect 54 334 55 335
rect 53 334 54 335
rect 52 334 53 335
rect 51 334 52 335
rect 50 334 51 335
rect 49 334 50 335
rect 48 334 49 335
rect 47 334 48 335
rect 46 334 47 335
rect 33 334 34 335
rect 32 334 33 335
rect 31 334 32 335
rect 30 334 31 335
rect 29 334 30 335
rect 28 334 29 335
rect 27 334 28 335
rect 26 334 27 335
rect 25 334 26 335
rect 24 334 25 335
rect 23 334 24 335
rect 22 334 23 335
rect 21 334 22 335
rect 20 334 21 335
rect 19 334 20 335
rect 18 334 19 335
rect 79 335 80 336
rect 78 335 79 336
rect 77 335 78 336
rect 76 335 77 336
rect 75 335 76 336
rect 74 335 75 336
rect 73 335 74 336
rect 72 335 73 336
rect 71 335 72 336
rect 70 335 71 336
rect 69 335 70 336
rect 68 335 69 336
rect 67 335 68 336
rect 66 335 67 336
rect 65 335 66 336
rect 64 335 65 336
rect 63 335 64 336
rect 62 335 63 336
rect 61 335 62 336
rect 60 335 61 336
rect 59 335 60 336
rect 58 335 59 336
rect 57 335 58 336
rect 56 335 57 336
rect 55 335 56 336
rect 54 335 55 336
rect 53 335 54 336
rect 52 335 53 336
rect 51 335 52 336
rect 50 335 51 336
rect 49 335 50 336
rect 48 335 49 336
rect 47 335 48 336
rect 33 335 34 336
rect 32 335 33 336
rect 31 335 32 336
rect 30 335 31 336
rect 29 335 30 336
rect 28 335 29 336
rect 27 335 28 336
rect 26 335 27 336
rect 25 335 26 336
rect 24 335 25 336
rect 23 335 24 336
rect 22 335 23 336
rect 21 335 22 336
rect 20 335 21 336
rect 19 335 20 336
rect 18 335 19 336
rect 78 336 79 337
rect 77 336 78 337
rect 76 336 77 337
rect 75 336 76 337
rect 74 336 75 337
rect 73 336 74 337
rect 72 336 73 337
rect 71 336 72 337
rect 70 336 71 337
rect 69 336 70 337
rect 68 336 69 337
rect 67 336 68 337
rect 66 336 67 337
rect 65 336 66 337
rect 64 336 65 337
rect 63 336 64 337
rect 62 336 63 337
rect 61 336 62 337
rect 60 336 61 337
rect 59 336 60 337
rect 58 336 59 337
rect 57 336 58 337
rect 56 336 57 337
rect 55 336 56 337
rect 54 336 55 337
rect 53 336 54 337
rect 52 336 53 337
rect 51 336 52 337
rect 50 336 51 337
rect 49 336 50 337
rect 48 336 49 337
rect 33 336 34 337
rect 32 336 33 337
rect 31 336 32 337
rect 30 336 31 337
rect 29 336 30 337
rect 28 336 29 337
rect 27 336 28 337
rect 26 336 27 337
rect 25 336 26 337
rect 24 336 25 337
rect 23 336 24 337
rect 22 336 23 337
rect 21 336 22 337
rect 20 336 21 337
rect 19 336 20 337
rect 18 336 19 337
rect 77 337 78 338
rect 76 337 77 338
rect 75 337 76 338
rect 74 337 75 338
rect 73 337 74 338
rect 72 337 73 338
rect 71 337 72 338
rect 70 337 71 338
rect 69 337 70 338
rect 68 337 69 338
rect 67 337 68 338
rect 66 337 67 338
rect 65 337 66 338
rect 64 337 65 338
rect 63 337 64 338
rect 62 337 63 338
rect 61 337 62 338
rect 60 337 61 338
rect 59 337 60 338
rect 58 337 59 338
rect 57 337 58 338
rect 56 337 57 338
rect 55 337 56 338
rect 54 337 55 338
rect 53 337 54 338
rect 52 337 53 338
rect 51 337 52 338
rect 50 337 51 338
rect 49 337 50 338
rect 48 337 49 338
rect 33 337 34 338
rect 32 337 33 338
rect 31 337 32 338
rect 30 337 31 338
rect 29 337 30 338
rect 28 337 29 338
rect 27 337 28 338
rect 26 337 27 338
rect 25 337 26 338
rect 24 337 25 338
rect 23 337 24 338
rect 22 337 23 338
rect 21 337 22 338
rect 20 337 21 338
rect 19 337 20 338
rect 18 337 19 338
rect 140 338 141 339
rect 139 338 140 339
rect 138 338 139 339
rect 137 338 138 339
rect 136 338 137 339
rect 135 338 136 339
rect 134 338 135 339
rect 75 338 76 339
rect 74 338 75 339
rect 73 338 74 339
rect 72 338 73 339
rect 71 338 72 339
rect 70 338 71 339
rect 69 338 70 339
rect 68 338 69 339
rect 67 338 68 339
rect 66 338 67 339
rect 65 338 66 339
rect 64 338 65 339
rect 63 338 64 339
rect 62 338 63 339
rect 61 338 62 339
rect 60 338 61 339
rect 59 338 60 339
rect 58 338 59 339
rect 57 338 58 339
rect 56 338 57 339
rect 55 338 56 339
rect 54 338 55 339
rect 53 338 54 339
rect 52 338 53 339
rect 51 338 52 339
rect 50 338 51 339
rect 33 338 34 339
rect 32 338 33 339
rect 31 338 32 339
rect 30 338 31 339
rect 29 338 30 339
rect 28 338 29 339
rect 27 338 28 339
rect 26 338 27 339
rect 25 338 26 339
rect 24 338 25 339
rect 23 338 24 339
rect 22 338 23 339
rect 21 338 22 339
rect 20 338 21 339
rect 19 338 20 339
rect 18 338 19 339
rect 143 339 144 340
rect 142 339 143 340
rect 141 339 142 340
rect 140 339 141 340
rect 139 339 140 340
rect 138 339 139 340
rect 137 339 138 340
rect 136 339 137 340
rect 135 339 136 340
rect 134 339 135 340
rect 133 339 134 340
rect 132 339 133 340
rect 74 339 75 340
rect 73 339 74 340
rect 72 339 73 340
rect 71 339 72 340
rect 70 339 71 340
rect 69 339 70 340
rect 68 339 69 340
rect 67 339 68 340
rect 66 339 67 340
rect 65 339 66 340
rect 64 339 65 340
rect 63 339 64 340
rect 62 339 63 340
rect 61 339 62 340
rect 60 339 61 340
rect 59 339 60 340
rect 58 339 59 340
rect 57 339 58 340
rect 56 339 57 340
rect 55 339 56 340
rect 54 339 55 340
rect 53 339 54 340
rect 52 339 53 340
rect 51 339 52 340
rect 33 339 34 340
rect 32 339 33 340
rect 31 339 32 340
rect 30 339 31 340
rect 29 339 30 340
rect 28 339 29 340
rect 27 339 28 340
rect 26 339 27 340
rect 25 339 26 340
rect 24 339 25 340
rect 23 339 24 340
rect 22 339 23 340
rect 21 339 22 340
rect 20 339 21 340
rect 19 339 20 340
rect 18 339 19 340
rect 144 340 145 341
rect 143 340 144 341
rect 142 340 143 341
rect 141 340 142 341
rect 140 340 141 341
rect 139 340 140 341
rect 138 340 139 341
rect 137 340 138 341
rect 136 340 137 341
rect 135 340 136 341
rect 134 340 135 341
rect 133 340 134 341
rect 132 340 133 341
rect 131 340 132 341
rect 72 340 73 341
rect 71 340 72 341
rect 70 340 71 341
rect 69 340 70 341
rect 68 340 69 341
rect 67 340 68 341
rect 66 340 67 341
rect 65 340 66 341
rect 64 340 65 341
rect 63 340 64 341
rect 62 340 63 341
rect 61 340 62 341
rect 60 340 61 341
rect 59 340 60 341
rect 58 340 59 341
rect 57 340 58 341
rect 56 340 57 341
rect 55 340 56 341
rect 54 340 55 341
rect 53 340 54 341
rect 52 340 53 341
rect 145 341 146 342
rect 144 341 145 342
rect 143 341 144 342
rect 142 341 143 342
rect 141 341 142 342
rect 140 341 141 342
rect 139 341 140 342
rect 138 341 139 342
rect 137 341 138 342
rect 136 341 137 342
rect 135 341 136 342
rect 134 341 135 342
rect 133 341 134 342
rect 132 341 133 342
rect 131 341 132 342
rect 130 341 131 342
rect 70 341 71 342
rect 69 341 70 342
rect 68 341 69 342
rect 67 341 68 342
rect 66 341 67 342
rect 65 341 66 342
rect 64 341 65 342
rect 63 341 64 342
rect 62 341 63 342
rect 61 341 62 342
rect 60 341 61 342
rect 59 341 60 342
rect 58 341 59 342
rect 57 341 58 342
rect 56 341 57 342
rect 55 341 56 342
rect 145 342 146 343
rect 144 342 145 343
rect 143 342 144 343
rect 142 342 143 343
rect 141 342 142 343
rect 140 342 141 343
rect 139 342 140 343
rect 138 342 139 343
rect 137 342 138 343
rect 136 342 137 343
rect 135 342 136 343
rect 134 342 135 343
rect 133 342 134 343
rect 132 342 133 343
rect 131 342 132 343
rect 130 342 131 343
rect 129 342 130 343
rect 65 342 66 343
rect 64 342 65 343
rect 63 342 64 343
rect 62 342 63 343
rect 61 342 62 343
rect 60 342 61 343
rect 59 342 60 343
rect 58 342 59 343
rect 146 343 147 344
rect 145 343 146 344
rect 144 343 145 344
rect 143 343 144 344
rect 142 343 143 344
rect 141 343 142 344
rect 140 343 141 344
rect 139 343 140 344
rect 138 343 139 344
rect 137 343 138 344
rect 136 343 137 344
rect 135 343 136 344
rect 134 343 135 344
rect 133 343 134 344
rect 132 343 133 344
rect 131 343 132 344
rect 130 343 131 344
rect 129 343 130 344
rect 146 344 147 345
rect 145 344 146 345
rect 144 344 145 345
rect 143 344 144 345
rect 142 344 143 345
rect 141 344 142 345
rect 133 344 134 345
rect 132 344 133 345
rect 131 344 132 345
rect 130 344 131 345
rect 129 344 130 345
rect 128 344 129 345
rect 146 345 147 346
rect 145 345 146 346
rect 144 345 145 346
rect 143 345 144 346
rect 142 345 143 346
rect 132 345 133 346
rect 131 345 132 346
rect 130 345 131 346
rect 129 345 130 346
rect 128 345 129 346
rect 146 346 147 347
rect 145 346 146 347
rect 144 346 145 347
rect 143 346 144 347
rect 142 346 143 347
rect 132 346 133 347
rect 131 346 132 347
rect 130 346 131 347
rect 129 346 130 347
rect 128 346 129 347
rect 146 347 147 348
rect 145 347 146 348
rect 144 347 145 348
rect 143 347 144 348
rect 131 347 132 348
rect 130 347 131 348
rect 129 347 130 348
rect 128 347 129 348
rect 145 348 146 349
rect 144 348 145 349
rect 143 348 144 349
rect 131 348 132 349
rect 130 348 131 349
rect 129 348 130 349
rect 128 348 129 349
rect 145 349 146 350
rect 144 349 145 350
rect 143 349 144 350
rect 142 349 143 350
rect 132 349 133 350
rect 131 349 132 350
rect 130 349 131 350
rect 129 349 130 350
rect 144 350 145 351
rect 143 350 144 351
rect 142 350 143 351
rect 141 350 142 351
rect 132 350 133 351
rect 131 350 132 351
rect 130 350 131 351
rect 129 350 130 351
rect 144 351 145 352
rect 143 351 144 352
rect 142 351 143 352
rect 141 351 142 352
rect 140 351 141 352
rect 139 351 140 352
rect 134 351 135 352
rect 133 351 134 352
rect 132 351 133 352
rect 131 351 132 352
rect 130 351 131 352
rect 146 352 147 353
rect 145 352 146 353
rect 144 352 145 353
rect 143 352 144 353
rect 142 352 143 353
rect 141 352 142 353
rect 140 352 141 353
rect 139 352 140 353
rect 138 352 139 353
rect 137 352 138 353
rect 136 352 137 353
rect 135 352 136 353
rect 134 352 135 353
rect 133 352 134 353
rect 132 352 133 353
rect 131 352 132 353
rect 130 352 131 353
rect 129 352 130 353
rect 128 352 129 353
rect 127 352 128 353
rect 126 352 127 353
rect 125 352 126 353
rect 124 352 125 353
rect 123 352 124 353
rect 122 352 123 353
rect 121 352 122 353
rect 120 352 121 353
rect 119 352 120 353
rect 57 352 58 353
rect 56 352 57 353
rect 55 352 56 353
rect 54 352 55 353
rect 53 352 54 353
rect 52 352 53 353
rect 51 352 52 353
rect 50 352 51 353
rect 49 352 50 353
rect 48 352 49 353
rect 47 352 48 353
rect 46 352 47 353
rect 146 353 147 354
rect 145 353 146 354
rect 144 353 145 354
rect 143 353 144 354
rect 142 353 143 354
rect 141 353 142 354
rect 140 353 141 354
rect 139 353 140 354
rect 138 353 139 354
rect 137 353 138 354
rect 136 353 137 354
rect 135 353 136 354
rect 134 353 135 354
rect 133 353 134 354
rect 132 353 133 354
rect 131 353 132 354
rect 130 353 131 354
rect 129 353 130 354
rect 128 353 129 354
rect 127 353 128 354
rect 126 353 127 354
rect 125 353 126 354
rect 124 353 125 354
rect 123 353 124 354
rect 122 353 123 354
rect 121 353 122 354
rect 120 353 121 354
rect 119 353 120 354
rect 65 353 66 354
rect 64 353 65 354
rect 63 353 64 354
rect 62 353 63 354
rect 61 353 62 354
rect 60 353 61 354
rect 59 353 60 354
rect 58 353 59 354
rect 57 353 58 354
rect 56 353 57 354
rect 55 353 56 354
rect 54 353 55 354
rect 53 353 54 354
rect 52 353 53 354
rect 51 353 52 354
rect 50 353 51 354
rect 49 353 50 354
rect 48 353 49 354
rect 47 353 48 354
rect 46 353 47 354
rect 45 353 46 354
rect 44 353 45 354
rect 43 353 44 354
rect 42 353 43 354
rect 41 353 42 354
rect 40 353 41 354
rect 39 353 40 354
rect 146 354 147 355
rect 145 354 146 355
rect 144 354 145 355
rect 143 354 144 355
rect 142 354 143 355
rect 141 354 142 355
rect 140 354 141 355
rect 139 354 140 355
rect 138 354 139 355
rect 137 354 138 355
rect 136 354 137 355
rect 135 354 136 355
rect 134 354 135 355
rect 133 354 134 355
rect 132 354 133 355
rect 131 354 132 355
rect 130 354 131 355
rect 129 354 130 355
rect 128 354 129 355
rect 127 354 128 355
rect 126 354 127 355
rect 125 354 126 355
rect 124 354 125 355
rect 123 354 124 355
rect 122 354 123 355
rect 121 354 122 355
rect 120 354 121 355
rect 119 354 120 355
rect 69 354 70 355
rect 68 354 69 355
rect 67 354 68 355
rect 66 354 67 355
rect 65 354 66 355
rect 64 354 65 355
rect 63 354 64 355
rect 62 354 63 355
rect 61 354 62 355
rect 60 354 61 355
rect 59 354 60 355
rect 58 354 59 355
rect 57 354 58 355
rect 56 354 57 355
rect 55 354 56 355
rect 54 354 55 355
rect 53 354 54 355
rect 52 354 53 355
rect 51 354 52 355
rect 50 354 51 355
rect 49 354 50 355
rect 48 354 49 355
rect 47 354 48 355
rect 46 354 47 355
rect 45 354 46 355
rect 44 354 45 355
rect 43 354 44 355
rect 42 354 43 355
rect 41 354 42 355
rect 40 354 41 355
rect 39 354 40 355
rect 38 354 39 355
rect 37 354 38 355
rect 36 354 37 355
rect 35 354 36 355
rect 146 355 147 356
rect 145 355 146 356
rect 144 355 145 356
rect 143 355 144 356
rect 142 355 143 356
rect 141 355 142 356
rect 140 355 141 356
rect 139 355 140 356
rect 138 355 139 356
rect 137 355 138 356
rect 136 355 137 356
rect 135 355 136 356
rect 134 355 135 356
rect 133 355 134 356
rect 132 355 133 356
rect 131 355 132 356
rect 130 355 131 356
rect 129 355 130 356
rect 128 355 129 356
rect 127 355 128 356
rect 126 355 127 356
rect 125 355 126 356
rect 124 355 125 356
rect 123 355 124 356
rect 122 355 123 356
rect 121 355 122 356
rect 120 355 121 356
rect 119 355 120 356
rect 71 355 72 356
rect 70 355 71 356
rect 69 355 70 356
rect 68 355 69 356
rect 67 355 68 356
rect 66 355 67 356
rect 65 355 66 356
rect 64 355 65 356
rect 63 355 64 356
rect 62 355 63 356
rect 61 355 62 356
rect 60 355 61 356
rect 59 355 60 356
rect 58 355 59 356
rect 57 355 58 356
rect 56 355 57 356
rect 55 355 56 356
rect 54 355 55 356
rect 53 355 54 356
rect 52 355 53 356
rect 51 355 52 356
rect 50 355 51 356
rect 49 355 50 356
rect 48 355 49 356
rect 47 355 48 356
rect 46 355 47 356
rect 45 355 46 356
rect 44 355 45 356
rect 43 355 44 356
rect 42 355 43 356
rect 41 355 42 356
rect 40 355 41 356
rect 39 355 40 356
rect 38 355 39 356
rect 37 355 38 356
rect 36 355 37 356
rect 35 355 36 356
rect 34 355 35 356
rect 33 355 34 356
rect 32 355 33 356
rect 146 356 147 357
rect 145 356 146 357
rect 144 356 145 357
rect 143 356 144 357
rect 142 356 143 357
rect 141 356 142 357
rect 140 356 141 357
rect 139 356 140 357
rect 138 356 139 357
rect 137 356 138 357
rect 136 356 137 357
rect 135 356 136 357
rect 134 356 135 357
rect 133 356 134 357
rect 132 356 133 357
rect 131 356 132 357
rect 130 356 131 357
rect 129 356 130 357
rect 128 356 129 357
rect 127 356 128 357
rect 126 356 127 357
rect 125 356 126 357
rect 124 356 125 357
rect 123 356 124 357
rect 122 356 123 357
rect 121 356 122 357
rect 120 356 121 357
rect 119 356 120 357
rect 73 356 74 357
rect 72 356 73 357
rect 71 356 72 357
rect 70 356 71 357
rect 69 356 70 357
rect 68 356 69 357
rect 67 356 68 357
rect 66 356 67 357
rect 65 356 66 357
rect 64 356 65 357
rect 63 356 64 357
rect 62 356 63 357
rect 61 356 62 357
rect 60 356 61 357
rect 59 356 60 357
rect 58 356 59 357
rect 57 356 58 357
rect 56 356 57 357
rect 55 356 56 357
rect 54 356 55 357
rect 53 356 54 357
rect 52 356 53 357
rect 51 356 52 357
rect 50 356 51 357
rect 49 356 50 357
rect 48 356 49 357
rect 47 356 48 357
rect 46 356 47 357
rect 45 356 46 357
rect 44 356 45 357
rect 43 356 44 357
rect 42 356 43 357
rect 41 356 42 357
rect 40 356 41 357
rect 39 356 40 357
rect 38 356 39 357
rect 37 356 38 357
rect 36 356 37 357
rect 35 356 36 357
rect 34 356 35 357
rect 33 356 34 357
rect 32 356 33 357
rect 31 356 32 357
rect 30 356 31 357
rect 75 357 76 358
rect 74 357 75 358
rect 73 357 74 358
rect 72 357 73 358
rect 71 357 72 358
rect 70 357 71 358
rect 69 357 70 358
rect 68 357 69 358
rect 67 357 68 358
rect 66 357 67 358
rect 65 357 66 358
rect 64 357 65 358
rect 63 357 64 358
rect 62 357 63 358
rect 61 357 62 358
rect 60 357 61 358
rect 59 357 60 358
rect 58 357 59 358
rect 57 357 58 358
rect 56 357 57 358
rect 55 357 56 358
rect 54 357 55 358
rect 53 357 54 358
rect 52 357 53 358
rect 51 357 52 358
rect 50 357 51 358
rect 49 357 50 358
rect 48 357 49 358
rect 47 357 48 358
rect 46 357 47 358
rect 45 357 46 358
rect 44 357 45 358
rect 43 357 44 358
rect 42 357 43 358
rect 41 357 42 358
rect 40 357 41 358
rect 39 357 40 358
rect 38 357 39 358
rect 37 357 38 358
rect 36 357 37 358
rect 35 357 36 358
rect 34 357 35 358
rect 33 357 34 358
rect 32 357 33 358
rect 31 357 32 358
rect 30 357 31 358
rect 29 357 30 358
rect 28 357 29 358
rect 77 358 78 359
rect 76 358 77 359
rect 75 358 76 359
rect 74 358 75 359
rect 73 358 74 359
rect 72 358 73 359
rect 71 358 72 359
rect 70 358 71 359
rect 69 358 70 359
rect 68 358 69 359
rect 67 358 68 359
rect 66 358 67 359
rect 65 358 66 359
rect 64 358 65 359
rect 63 358 64 359
rect 62 358 63 359
rect 61 358 62 359
rect 60 358 61 359
rect 59 358 60 359
rect 58 358 59 359
rect 57 358 58 359
rect 56 358 57 359
rect 55 358 56 359
rect 54 358 55 359
rect 53 358 54 359
rect 52 358 53 359
rect 51 358 52 359
rect 50 358 51 359
rect 49 358 50 359
rect 48 358 49 359
rect 47 358 48 359
rect 46 358 47 359
rect 45 358 46 359
rect 44 358 45 359
rect 43 358 44 359
rect 42 358 43 359
rect 41 358 42 359
rect 40 358 41 359
rect 39 358 40 359
rect 38 358 39 359
rect 37 358 38 359
rect 36 358 37 359
rect 35 358 36 359
rect 34 358 35 359
rect 33 358 34 359
rect 32 358 33 359
rect 31 358 32 359
rect 30 358 31 359
rect 29 358 30 359
rect 28 358 29 359
rect 27 358 28 359
rect 78 359 79 360
rect 77 359 78 360
rect 76 359 77 360
rect 75 359 76 360
rect 74 359 75 360
rect 73 359 74 360
rect 72 359 73 360
rect 71 359 72 360
rect 70 359 71 360
rect 69 359 70 360
rect 68 359 69 360
rect 67 359 68 360
rect 66 359 67 360
rect 65 359 66 360
rect 64 359 65 360
rect 63 359 64 360
rect 62 359 63 360
rect 61 359 62 360
rect 60 359 61 360
rect 59 359 60 360
rect 58 359 59 360
rect 57 359 58 360
rect 56 359 57 360
rect 55 359 56 360
rect 54 359 55 360
rect 53 359 54 360
rect 52 359 53 360
rect 51 359 52 360
rect 50 359 51 360
rect 49 359 50 360
rect 48 359 49 360
rect 47 359 48 360
rect 46 359 47 360
rect 45 359 46 360
rect 44 359 45 360
rect 43 359 44 360
rect 42 359 43 360
rect 41 359 42 360
rect 40 359 41 360
rect 39 359 40 360
rect 38 359 39 360
rect 37 359 38 360
rect 36 359 37 360
rect 35 359 36 360
rect 34 359 35 360
rect 33 359 34 360
rect 32 359 33 360
rect 31 359 32 360
rect 30 359 31 360
rect 29 359 30 360
rect 28 359 29 360
rect 27 359 28 360
rect 26 359 27 360
rect 79 360 80 361
rect 78 360 79 361
rect 77 360 78 361
rect 76 360 77 361
rect 75 360 76 361
rect 74 360 75 361
rect 73 360 74 361
rect 72 360 73 361
rect 71 360 72 361
rect 70 360 71 361
rect 69 360 70 361
rect 68 360 69 361
rect 67 360 68 361
rect 66 360 67 361
rect 65 360 66 361
rect 64 360 65 361
rect 63 360 64 361
rect 62 360 63 361
rect 61 360 62 361
rect 60 360 61 361
rect 59 360 60 361
rect 58 360 59 361
rect 57 360 58 361
rect 56 360 57 361
rect 55 360 56 361
rect 54 360 55 361
rect 53 360 54 361
rect 52 360 53 361
rect 51 360 52 361
rect 50 360 51 361
rect 49 360 50 361
rect 48 360 49 361
rect 47 360 48 361
rect 46 360 47 361
rect 45 360 46 361
rect 44 360 45 361
rect 43 360 44 361
rect 42 360 43 361
rect 41 360 42 361
rect 40 360 41 361
rect 39 360 40 361
rect 38 360 39 361
rect 37 360 38 361
rect 36 360 37 361
rect 35 360 36 361
rect 34 360 35 361
rect 33 360 34 361
rect 32 360 33 361
rect 31 360 32 361
rect 30 360 31 361
rect 29 360 30 361
rect 28 360 29 361
rect 27 360 28 361
rect 26 360 27 361
rect 25 360 26 361
rect 24 360 25 361
rect 80 361 81 362
rect 79 361 80 362
rect 78 361 79 362
rect 77 361 78 362
rect 76 361 77 362
rect 75 361 76 362
rect 74 361 75 362
rect 73 361 74 362
rect 72 361 73 362
rect 71 361 72 362
rect 70 361 71 362
rect 69 361 70 362
rect 68 361 69 362
rect 67 361 68 362
rect 66 361 67 362
rect 65 361 66 362
rect 64 361 65 362
rect 63 361 64 362
rect 62 361 63 362
rect 61 361 62 362
rect 60 361 61 362
rect 59 361 60 362
rect 58 361 59 362
rect 57 361 58 362
rect 56 361 57 362
rect 55 361 56 362
rect 54 361 55 362
rect 53 361 54 362
rect 52 361 53 362
rect 51 361 52 362
rect 50 361 51 362
rect 49 361 50 362
rect 48 361 49 362
rect 47 361 48 362
rect 46 361 47 362
rect 45 361 46 362
rect 44 361 45 362
rect 43 361 44 362
rect 42 361 43 362
rect 41 361 42 362
rect 40 361 41 362
rect 39 361 40 362
rect 38 361 39 362
rect 37 361 38 362
rect 36 361 37 362
rect 35 361 36 362
rect 34 361 35 362
rect 33 361 34 362
rect 32 361 33 362
rect 31 361 32 362
rect 30 361 31 362
rect 29 361 30 362
rect 28 361 29 362
rect 27 361 28 362
rect 26 361 27 362
rect 25 361 26 362
rect 24 361 25 362
rect 23 361 24 362
rect 81 362 82 363
rect 80 362 81 363
rect 79 362 80 363
rect 78 362 79 363
rect 77 362 78 363
rect 76 362 77 363
rect 75 362 76 363
rect 74 362 75 363
rect 73 362 74 363
rect 72 362 73 363
rect 71 362 72 363
rect 70 362 71 363
rect 69 362 70 363
rect 68 362 69 363
rect 67 362 68 363
rect 66 362 67 363
rect 65 362 66 363
rect 64 362 65 363
rect 63 362 64 363
rect 62 362 63 363
rect 61 362 62 363
rect 60 362 61 363
rect 59 362 60 363
rect 58 362 59 363
rect 57 362 58 363
rect 56 362 57 363
rect 55 362 56 363
rect 54 362 55 363
rect 53 362 54 363
rect 52 362 53 363
rect 51 362 52 363
rect 50 362 51 363
rect 49 362 50 363
rect 48 362 49 363
rect 47 362 48 363
rect 46 362 47 363
rect 45 362 46 363
rect 44 362 45 363
rect 43 362 44 363
rect 42 362 43 363
rect 41 362 42 363
rect 40 362 41 363
rect 39 362 40 363
rect 38 362 39 363
rect 37 362 38 363
rect 36 362 37 363
rect 35 362 36 363
rect 34 362 35 363
rect 33 362 34 363
rect 32 362 33 363
rect 31 362 32 363
rect 30 362 31 363
rect 29 362 30 363
rect 28 362 29 363
rect 27 362 28 363
rect 26 362 27 363
rect 25 362 26 363
rect 24 362 25 363
rect 23 362 24 363
rect 22 362 23 363
rect 146 363 147 364
rect 145 363 146 364
rect 144 363 145 364
rect 143 363 144 364
rect 142 363 143 364
rect 141 363 142 364
rect 140 363 141 364
rect 139 363 140 364
rect 138 363 139 364
rect 137 363 138 364
rect 136 363 137 364
rect 135 363 136 364
rect 134 363 135 364
rect 133 363 134 364
rect 132 363 133 364
rect 131 363 132 364
rect 130 363 131 364
rect 129 363 130 364
rect 128 363 129 364
rect 127 363 128 364
rect 126 363 127 364
rect 125 363 126 364
rect 124 363 125 364
rect 123 363 124 364
rect 122 363 123 364
rect 121 363 122 364
rect 81 363 82 364
rect 80 363 81 364
rect 79 363 80 364
rect 78 363 79 364
rect 77 363 78 364
rect 76 363 77 364
rect 75 363 76 364
rect 74 363 75 364
rect 73 363 74 364
rect 72 363 73 364
rect 71 363 72 364
rect 70 363 71 364
rect 69 363 70 364
rect 68 363 69 364
rect 67 363 68 364
rect 66 363 67 364
rect 65 363 66 364
rect 64 363 65 364
rect 63 363 64 364
rect 62 363 63 364
rect 61 363 62 364
rect 60 363 61 364
rect 59 363 60 364
rect 58 363 59 364
rect 57 363 58 364
rect 56 363 57 364
rect 55 363 56 364
rect 54 363 55 364
rect 53 363 54 364
rect 52 363 53 364
rect 51 363 52 364
rect 50 363 51 364
rect 49 363 50 364
rect 48 363 49 364
rect 47 363 48 364
rect 46 363 47 364
rect 45 363 46 364
rect 44 363 45 364
rect 43 363 44 364
rect 42 363 43 364
rect 41 363 42 364
rect 40 363 41 364
rect 39 363 40 364
rect 38 363 39 364
rect 37 363 38 364
rect 36 363 37 364
rect 35 363 36 364
rect 34 363 35 364
rect 33 363 34 364
rect 32 363 33 364
rect 31 363 32 364
rect 30 363 31 364
rect 29 363 30 364
rect 28 363 29 364
rect 27 363 28 364
rect 26 363 27 364
rect 25 363 26 364
rect 24 363 25 364
rect 23 363 24 364
rect 22 363 23 364
rect 146 364 147 365
rect 145 364 146 365
rect 144 364 145 365
rect 143 364 144 365
rect 142 364 143 365
rect 141 364 142 365
rect 140 364 141 365
rect 139 364 140 365
rect 138 364 139 365
rect 137 364 138 365
rect 136 364 137 365
rect 135 364 136 365
rect 134 364 135 365
rect 133 364 134 365
rect 132 364 133 365
rect 131 364 132 365
rect 130 364 131 365
rect 129 364 130 365
rect 128 364 129 365
rect 127 364 128 365
rect 126 364 127 365
rect 125 364 126 365
rect 124 364 125 365
rect 123 364 124 365
rect 122 364 123 365
rect 121 364 122 365
rect 82 364 83 365
rect 81 364 82 365
rect 80 364 81 365
rect 79 364 80 365
rect 78 364 79 365
rect 77 364 78 365
rect 76 364 77 365
rect 75 364 76 365
rect 74 364 75 365
rect 73 364 74 365
rect 72 364 73 365
rect 71 364 72 365
rect 70 364 71 365
rect 69 364 70 365
rect 68 364 69 365
rect 67 364 68 365
rect 66 364 67 365
rect 65 364 66 365
rect 64 364 65 365
rect 63 364 64 365
rect 62 364 63 365
rect 61 364 62 365
rect 60 364 61 365
rect 59 364 60 365
rect 58 364 59 365
rect 57 364 58 365
rect 56 364 57 365
rect 55 364 56 365
rect 54 364 55 365
rect 53 364 54 365
rect 52 364 53 365
rect 51 364 52 365
rect 50 364 51 365
rect 49 364 50 365
rect 48 364 49 365
rect 47 364 48 365
rect 46 364 47 365
rect 45 364 46 365
rect 44 364 45 365
rect 43 364 44 365
rect 42 364 43 365
rect 41 364 42 365
rect 40 364 41 365
rect 39 364 40 365
rect 38 364 39 365
rect 37 364 38 365
rect 36 364 37 365
rect 35 364 36 365
rect 34 364 35 365
rect 33 364 34 365
rect 32 364 33 365
rect 31 364 32 365
rect 30 364 31 365
rect 29 364 30 365
rect 28 364 29 365
rect 27 364 28 365
rect 26 364 27 365
rect 25 364 26 365
rect 24 364 25 365
rect 23 364 24 365
rect 22 364 23 365
rect 21 364 22 365
rect 146 365 147 366
rect 145 365 146 366
rect 144 365 145 366
rect 143 365 144 366
rect 142 365 143 366
rect 141 365 142 366
rect 140 365 141 366
rect 139 365 140 366
rect 138 365 139 366
rect 137 365 138 366
rect 136 365 137 366
rect 135 365 136 366
rect 134 365 135 366
rect 133 365 134 366
rect 132 365 133 366
rect 131 365 132 366
rect 130 365 131 366
rect 129 365 130 366
rect 128 365 129 366
rect 127 365 128 366
rect 126 365 127 366
rect 125 365 126 366
rect 124 365 125 366
rect 123 365 124 366
rect 122 365 123 366
rect 121 365 122 366
rect 82 365 83 366
rect 81 365 82 366
rect 80 365 81 366
rect 79 365 80 366
rect 78 365 79 366
rect 77 365 78 366
rect 76 365 77 366
rect 75 365 76 366
rect 74 365 75 366
rect 73 365 74 366
rect 72 365 73 366
rect 71 365 72 366
rect 70 365 71 366
rect 69 365 70 366
rect 68 365 69 366
rect 67 365 68 366
rect 66 365 67 366
rect 65 365 66 366
rect 64 365 65 366
rect 63 365 64 366
rect 62 365 63 366
rect 61 365 62 366
rect 60 365 61 366
rect 59 365 60 366
rect 58 365 59 366
rect 57 365 58 366
rect 56 365 57 366
rect 55 365 56 366
rect 54 365 55 366
rect 53 365 54 366
rect 52 365 53 366
rect 51 365 52 366
rect 50 365 51 366
rect 49 365 50 366
rect 48 365 49 366
rect 47 365 48 366
rect 46 365 47 366
rect 45 365 46 366
rect 44 365 45 366
rect 43 365 44 366
rect 42 365 43 366
rect 41 365 42 366
rect 40 365 41 366
rect 39 365 40 366
rect 38 365 39 366
rect 37 365 38 366
rect 36 365 37 366
rect 35 365 36 366
rect 34 365 35 366
rect 33 365 34 366
rect 32 365 33 366
rect 31 365 32 366
rect 30 365 31 366
rect 29 365 30 366
rect 28 365 29 366
rect 27 365 28 366
rect 26 365 27 366
rect 25 365 26 366
rect 24 365 25 366
rect 23 365 24 366
rect 22 365 23 366
rect 21 365 22 366
rect 20 365 21 366
rect 146 366 147 367
rect 145 366 146 367
rect 144 366 145 367
rect 143 366 144 367
rect 142 366 143 367
rect 141 366 142 367
rect 140 366 141 367
rect 139 366 140 367
rect 138 366 139 367
rect 137 366 138 367
rect 136 366 137 367
rect 135 366 136 367
rect 134 366 135 367
rect 133 366 134 367
rect 132 366 133 367
rect 131 366 132 367
rect 130 366 131 367
rect 129 366 130 367
rect 128 366 129 367
rect 127 366 128 367
rect 126 366 127 367
rect 125 366 126 367
rect 124 366 125 367
rect 123 366 124 367
rect 122 366 123 367
rect 121 366 122 367
rect 83 366 84 367
rect 82 366 83 367
rect 81 366 82 367
rect 80 366 81 367
rect 79 366 80 367
rect 78 366 79 367
rect 77 366 78 367
rect 76 366 77 367
rect 75 366 76 367
rect 74 366 75 367
rect 73 366 74 367
rect 72 366 73 367
rect 71 366 72 367
rect 70 366 71 367
rect 69 366 70 367
rect 68 366 69 367
rect 67 366 68 367
rect 66 366 67 367
rect 65 366 66 367
rect 64 366 65 367
rect 63 366 64 367
rect 62 366 63 367
rect 61 366 62 367
rect 60 366 61 367
rect 59 366 60 367
rect 58 366 59 367
rect 57 366 58 367
rect 56 366 57 367
rect 55 366 56 367
rect 54 366 55 367
rect 53 366 54 367
rect 52 366 53 367
rect 51 366 52 367
rect 50 366 51 367
rect 49 366 50 367
rect 48 366 49 367
rect 47 366 48 367
rect 46 366 47 367
rect 45 366 46 367
rect 44 366 45 367
rect 43 366 44 367
rect 42 366 43 367
rect 41 366 42 367
rect 40 366 41 367
rect 39 366 40 367
rect 38 366 39 367
rect 37 366 38 367
rect 36 366 37 367
rect 35 366 36 367
rect 34 366 35 367
rect 33 366 34 367
rect 32 366 33 367
rect 31 366 32 367
rect 30 366 31 367
rect 29 366 30 367
rect 28 366 29 367
rect 27 366 28 367
rect 26 366 27 367
rect 25 366 26 367
rect 24 366 25 367
rect 23 366 24 367
rect 22 366 23 367
rect 21 366 22 367
rect 20 366 21 367
rect 146 367 147 368
rect 145 367 146 368
rect 144 367 145 368
rect 143 367 144 368
rect 142 367 143 368
rect 141 367 142 368
rect 140 367 141 368
rect 139 367 140 368
rect 138 367 139 368
rect 137 367 138 368
rect 136 367 137 368
rect 135 367 136 368
rect 134 367 135 368
rect 133 367 134 368
rect 132 367 133 368
rect 131 367 132 368
rect 130 367 131 368
rect 129 367 130 368
rect 128 367 129 368
rect 127 367 128 368
rect 126 367 127 368
rect 125 367 126 368
rect 124 367 125 368
rect 123 367 124 368
rect 122 367 123 368
rect 121 367 122 368
rect 83 367 84 368
rect 82 367 83 368
rect 81 367 82 368
rect 80 367 81 368
rect 79 367 80 368
rect 78 367 79 368
rect 77 367 78 368
rect 76 367 77 368
rect 75 367 76 368
rect 74 367 75 368
rect 73 367 74 368
rect 72 367 73 368
rect 71 367 72 368
rect 70 367 71 368
rect 69 367 70 368
rect 68 367 69 368
rect 67 367 68 368
rect 66 367 67 368
rect 65 367 66 368
rect 64 367 65 368
rect 63 367 64 368
rect 62 367 63 368
rect 61 367 62 368
rect 60 367 61 368
rect 59 367 60 368
rect 58 367 59 368
rect 57 367 58 368
rect 56 367 57 368
rect 55 367 56 368
rect 54 367 55 368
rect 53 367 54 368
rect 52 367 53 368
rect 51 367 52 368
rect 50 367 51 368
rect 49 367 50 368
rect 48 367 49 368
rect 47 367 48 368
rect 46 367 47 368
rect 45 367 46 368
rect 44 367 45 368
rect 43 367 44 368
rect 42 367 43 368
rect 41 367 42 368
rect 40 367 41 368
rect 39 367 40 368
rect 38 367 39 368
rect 37 367 38 368
rect 36 367 37 368
rect 35 367 36 368
rect 34 367 35 368
rect 33 367 34 368
rect 32 367 33 368
rect 31 367 32 368
rect 30 367 31 368
rect 29 367 30 368
rect 28 367 29 368
rect 27 367 28 368
rect 26 367 27 368
rect 25 367 26 368
rect 24 367 25 368
rect 23 367 24 368
rect 22 367 23 368
rect 21 367 22 368
rect 20 367 21 368
rect 19 367 20 368
rect 134 368 135 369
rect 133 368 134 369
rect 132 368 133 369
rect 84 368 85 369
rect 83 368 84 369
rect 82 368 83 369
rect 81 368 82 369
rect 80 368 81 369
rect 79 368 80 369
rect 78 368 79 369
rect 77 368 78 369
rect 76 368 77 369
rect 75 368 76 369
rect 74 368 75 369
rect 73 368 74 369
rect 72 368 73 369
rect 71 368 72 369
rect 70 368 71 369
rect 69 368 70 369
rect 68 368 69 369
rect 67 368 68 369
rect 66 368 67 369
rect 65 368 66 369
rect 64 368 65 369
rect 63 368 64 369
rect 62 368 63 369
rect 61 368 62 369
rect 60 368 61 369
rect 59 368 60 369
rect 58 368 59 369
rect 57 368 58 369
rect 56 368 57 369
rect 55 368 56 369
rect 54 368 55 369
rect 53 368 54 369
rect 52 368 53 369
rect 51 368 52 369
rect 50 368 51 369
rect 49 368 50 369
rect 48 368 49 369
rect 47 368 48 369
rect 46 368 47 369
rect 45 368 46 369
rect 44 368 45 369
rect 43 368 44 369
rect 42 368 43 369
rect 41 368 42 369
rect 40 368 41 369
rect 39 368 40 369
rect 38 368 39 369
rect 37 368 38 369
rect 36 368 37 369
rect 35 368 36 369
rect 34 368 35 369
rect 33 368 34 369
rect 32 368 33 369
rect 31 368 32 369
rect 30 368 31 369
rect 29 368 30 369
rect 28 368 29 369
rect 27 368 28 369
rect 26 368 27 369
rect 25 368 26 369
rect 24 368 25 369
rect 23 368 24 369
rect 22 368 23 369
rect 21 368 22 369
rect 20 368 21 369
rect 19 368 20 369
rect 135 369 136 370
rect 134 369 135 370
rect 133 369 134 370
rect 132 369 133 370
rect 84 369 85 370
rect 83 369 84 370
rect 82 369 83 370
rect 81 369 82 370
rect 80 369 81 370
rect 79 369 80 370
rect 78 369 79 370
rect 77 369 78 370
rect 76 369 77 370
rect 75 369 76 370
rect 74 369 75 370
rect 73 369 74 370
rect 72 369 73 370
rect 71 369 72 370
rect 70 369 71 370
rect 69 369 70 370
rect 68 369 69 370
rect 67 369 68 370
rect 66 369 67 370
rect 65 369 66 370
rect 64 369 65 370
rect 63 369 64 370
rect 62 369 63 370
rect 61 369 62 370
rect 60 369 61 370
rect 59 369 60 370
rect 58 369 59 370
rect 57 369 58 370
rect 56 369 57 370
rect 55 369 56 370
rect 54 369 55 370
rect 53 369 54 370
rect 52 369 53 370
rect 51 369 52 370
rect 50 369 51 370
rect 49 369 50 370
rect 48 369 49 370
rect 47 369 48 370
rect 46 369 47 370
rect 45 369 46 370
rect 44 369 45 370
rect 43 369 44 370
rect 42 369 43 370
rect 41 369 42 370
rect 40 369 41 370
rect 39 369 40 370
rect 38 369 39 370
rect 37 369 38 370
rect 36 369 37 370
rect 35 369 36 370
rect 34 369 35 370
rect 33 369 34 370
rect 32 369 33 370
rect 31 369 32 370
rect 30 369 31 370
rect 29 369 30 370
rect 28 369 29 370
rect 27 369 28 370
rect 26 369 27 370
rect 25 369 26 370
rect 24 369 25 370
rect 23 369 24 370
rect 22 369 23 370
rect 21 369 22 370
rect 20 369 21 370
rect 19 369 20 370
rect 136 370 137 371
rect 135 370 136 371
rect 134 370 135 371
rect 133 370 134 371
rect 132 370 133 371
rect 131 370 132 371
rect 130 370 131 371
rect 84 370 85 371
rect 83 370 84 371
rect 82 370 83 371
rect 81 370 82 371
rect 80 370 81 371
rect 79 370 80 371
rect 78 370 79 371
rect 77 370 78 371
rect 76 370 77 371
rect 75 370 76 371
rect 74 370 75 371
rect 73 370 74 371
rect 72 370 73 371
rect 71 370 72 371
rect 70 370 71 371
rect 69 370 70 371
rect 68 370 69 371
rect 67 370 68 371
rect 66 370 67 371
rect 65 370 66 371
rect 64 370 65 371
rect 63 370 64 371
rect 62 370 63 371
rect 61 370 62 371
rect 60 370 61 371
rect 59 370 60 371
rect 58 370 59 371
rect 57 370 58 371
rect 56 370 57 371
rect 55 370 56 371
rect 54 370 55 371
rect 53 370 54 371
rect 52 370 53 371
rect 51 370 52 371
rect 50 370 51 371
rect 49 370 50 371
rect 48 370 49 371
rect 47 370 48 371
rect 46 370 47 371
rect 45 370 46 371
rect 44 370 45 371
rect 43 370 44 371
rect 42 370 43 371
rect 41 370 42 371
rect 40 370 41 371
rect 39 370 40 371
rect 38 370 39 371
rect 37 370 38 371
rect 36 370 37 371
rect 35 370 36 371
rect 34 370 35 371
rect 33 370 34 371
rect 32 370 33 371
rect 31 370 32 371
rect 30 370 31 371
rect 29 370 30 371
rect 28 370 29 371
rect 27 370 28 371
rect 26 370 27 371
rect 25 370 26 371
rect 24 370 25 371
rect 23 370 24 371
rect 22 370 23 371
rect 21 370 22 371
rect 20 370 21 371
rect 19 370 20 371
rect 18 370 19 371
rect 138 371 139 372
rect 137 371 138 372
rect 136 371 137 372
rect 135 371 136 372
rect 134 371 135 372
rect 133 371 134 372
rect 132 371 133 372
rect 131 371 132 372
rect 130 371 131 372
rect 129 371 130 372
rect 84 371 85 372
rect 83 371 84 372
rect 82 371 83 372
rect 81 371 82 372
rect 80 371 81 372
rect 79 371 80 372
rect 78 371 79 372
rect 77 371 78 372
rect 76 371 77 372
rect 75 371 76 372
rect 74 371 75 372
rect 73 371 74 372
rect 72 371 73 372
rect 71 371 72 372
rect 70 371 71 372
rect 69 371 70 372
rect 68 371 69 372
rect 67 371 68 372
rect 66 371 67 372
rect 65 371 66 372
rect 64 371 65 372
rect 63 371 64 372
rect 62 371 63 372
rect 61 371 62 372
rect 60 371 61 372
rect 59 371 60 372
rect 58 371 59 372
rect 57 371 58 372
rect 56 371 57 372
rect 55 371 56 372
rect 54 371 55 372
rect 53 371 54 372
rect 52 371 53 372
rect 51 371 52 372
rect 50 371 51 372
rect 49 371 50 372
rect 48 371 49 372
rect 47 371 48 372
rect 46 371 47 372
rect 45 371 46 372
rect 44 371 45 372
rect 43 371 44 372
rect 42 371 43 372
rect 41 371 42 372
rect 40 371 41 372
rect 39 371 40 372
rect 38 371 39 372
rect 37 371 38 372
rect 36 371 37 372
rect 35 371 36 372
rect 34 371 35 372
rect 33 371 34 372
rect 32 371 33 372
rect 31 371 32 372
rect 30 371 31 372
rect 29 371 30 372
rect 28 371 29 372
rect 27 371 28 372
rect 26 371 27 372
rect 25 371 26 372
rect 24 371 25 372
rect 23 371 24 372
rect 22 371 23 372
rect 21 371 22 372
rect 20 371 21 372
rect 19 371 20 372
rect 18 371 19 372
rect 139 372 140 373
rect 138 372 139 373
rect 137 372 138 373
rect 136 372 137 373
rect 135 372 136 373
rect 134 372 135 373
rect 133 372 134 373
rect 132 372 133 373
rect 131 372 132 373
rect 130 372 131 373
rect 129 372 130 373
rect 128 372 129 373
rect 127 372 128 373
rect 85 372 86 373
rect 84 372 85 373
rect 83 372 84 373
rect 82 372 83 373
rect 81 372 82 373
rect 80 372 81 373
rect 79 372 80 373
rect 78 372 79 373
rect 77 372 78 373
rect 76 372 77 373
rect 75 372 76 373
rect 74 372 75 373
rect 73 372 74 373
rect 72 372 73 373
rect 71 372 72 373
rect 70 372 71 373
rect 69 372 70 373
rect 68 372 69 373
rect 67 372 68 373
rect 66 372 67 373
rect 65 372 66 373
rect 64 372 65 373
rect 63 372 64 373
rect 62 372 63 373
rect 41 372 42 373
rect 40 372 41 373
rect 39 372 40 373
rect 38 372 39 373
rect 37 372 38 373
rect 36 372 37 373
rect 35 372 36 373
rect 34 372 35 373
rect 33 372 34 373
rect 32 372 33 373
rect 31 372 32 373
rect 30 372 31 373
rect 29 372 30 373
rect 28 372 29 373
rect 27 372 28 373
rect 26 372 27 373
rect 25 372 26 373
rect 24 372 25 373
rect 23 372 24 373
rect 22 372 23 373
rect 21 372 22 373
rect 20 372 21 373
rect 19 372 20 373
rect 18 372 19 373
rect 141 373 142 374
rect 140 373 141 374
rect 139 373 140 374
rect 138 373 139 374
rect 137 373 138 374
rect 136 373 137 374
rect 135 373 136 374
rect 134 373 135 374
rect 133 373 134 374
rect 132 373 133 374
rect 131 373 132 374
rect 130 373 131 374
rect 129 373 130 374
rect 128 373 129 374
rect 127 373 128 374
rect 126 373 127 374
rect 85 373 86 374
rect 84 373 85 374
rect 83 373 84 374
rect 82 373 83 374
rect 81 373 82 374
rect 80 373 81 374
rect 79 373 80 374
rect 78 373 79 374
rect 77 373 78 374
rect 76 373 77 374
rect 75 373 76 374
rect 74 373 75 374
rect 73 373 74 374
rect 72 373 73 374
rect 71 373 72 374
rect 70 373 71 374
rect 69 373 70 374
rect 68 373 69 374
rect 67 373 68 374
rect 36 373 37 374
rect 35 373 36 374
rect 34 373 35 374
rect 33 373 34 374
rect 32 373 33 374
rect 31 373 32 374
rect 30 373 31 374
rect 29 373 30 374
rect 28 373 29 374
rect 27 373 28 374
rect 26 373 27 374
rect 25 373 26 374
rect 24 373 25 374
rect 23 373 24 374
rect 22 373 23 374
rect 21 373 22 374
rect 20 373 21 374
rect 19 373 20 374
rect 18 373 19 374
rect 142 374 143 375
rect 141 374 142 375
rect 140 374 141 375
rect 139 374 140 375
rect 138 374 139 375
rect 137 374 138 375
rect 136 374 137 375
rect 135 374 136 375
rect 134 374 135 375
rect 133 374 134 375
rect 132 374 133 375
rect 131 374 132 375
rect 130 374 131 375
rect 129 374 130 375
rect 128 374 129 375
rect 127 374 128 375
rect 126 374 127 375
rect 125 374 126 375
rect 124 374 125 375
rect 85 374 86 375
rect 84 374 85 375
rect 83 374 84 375
rect 82 374 83 375
rect 81 374 82 375
rect 80 374 81 375
rect 79 374 80 375
rect 78 374 79 375
rect 77 374 78 375
rect 76 374 77 375
rect 75 374 76 375
rect 74 374 75 375
rect 73 374 74 375
rect 72 374 73 375
rect 71 374 72 375
rect 70 374 71 375
rect 69 374 70 375
rect 33 374 34 375
rect 32 374 33 375
rect 31 374 32 375
rect 30 374 31 375
rect 29 374 30 375
rect 28 374 29 375
rect 27 374 28 375
rect 26 374 27 375
rect 25 374 26 375
rect 24 374 25 375
rect 23 374 24 375
rect 22 374 23 375
rect 21 374 22 375
rect 20 374 21 375
rect 19 374 20 375
rect 18 374 19 375
rect 17 374 18 375
rect 144 375 145 376
rect 143 375 144 376
rect 142 375 143 376
rect 141 375 142 376
rect 140 375 141 376
rect 139 375 140 376
rect 138 375 139 376
rect 137 375 138 376
rect 136 375 137 376
rect 135 375 136 376
rect 131 375 132 376
rect 130 375 131 376
rect 129 375 130 376
rect 128 375 129 376
rect 127 375 128 376
rect 126 375 127 376
rect 125 375 126 376
rect 124 375 125 376
rect 123 375 124 376
rect 85 375 86 376
rect 84 375 85 376
rect 83 375 84 376
rect 82 375 83 376
rect 81 375 82 376
rect 80 375 81 376
rect 79 375 80 376
rect 78 375 79 376
rect 77 375 78 376
rect 76 375 77 376
rect 75 375 76 376
rect 74 375 75 376
rect 73 375 74 376
rect 72 375 73 376
rect 71 375 72 376
rect 70 375 71 376
rect 32 375 33 376
rect 31 375 32 376
rect 30 375 31 376
rect 29 375 30 376
rect 28 375 29 376
rect 27 375 28 376
rect 26 375 27 376
rect 25 375 26 376
rect 24 375 25 376
rect 23 375 24 376
rect 22 375 23 376
rect 21 375 22 376
rect 20 375 21 376
rect 19 375 20 376
rect 18 375 19 376
rect 17 375 18 376
rect 145 376 146 377
rect 144 376 145 377
rect 143 376 144 377
rect 142 376 143 377
rect 141 376 142 377
rect 140 376 141 377
rect 139 376 140 377
rect 138 376 139 377
rect 137 376 138 377
rect 136 376 137 377
rect 130 376 131 377
rect 129 376 130 377
rect 128 376 129 377
rect 127 376 128 377
rect 126 376 127 377
rect 125 376 126 377
rect 124 376 125 377
rect 123 376 124 377
rect 122 376 123 377
rect 121 376 122 377
rect 85 376 86 377
rect 84 376 85 377
rect 83 376 84 377
rect 82 376 83 377
rect 81 376 82 377
rect 80 376 81 377
rect 79 376 80 377
rect 78 376 79 377
rect 77 376 78 377
rect 76 376 77 377
rect 75 376 76 377
rect 74 376 75 377
rect 73 376 74 377
rect 72 376 73 377
rect 71 376 72 377
rect 31 376 32 377
rect 30 376 31 377
rect 29 376 30 377
rect 28 376 29 377
rect 27 376 28 377
rect 26 376 27 377
rect 25 376 26 377
rect 24 376 25 377
rect 23 376 24 377
rect 22 376 23 377
rect 21 376 22 377
rect 20 376 21 377
rect 19 376 20 377
rect 18 376 19 377
rect 17 376 18 377
rect 146 377 147 378
rect 145 377 146 378
rect 144 377 145 378
rect 143 377 144 378
rect 142 377 143 378
rect 141 377 142 378
rect 140 377 141 378
rect 139 377 140 378
rect 138 377 139 378
rect 128 377 129 378
rect 127 377 128 378
rect 126 377 127 378
rect 125 377 126 378
rect 124 377 125 378
rect 123 377 124 378
rect 122 377 123 378
rect 121 377 122 378
rect 85 377 86 378
rect 84 377 85 378
rect 83 377 84 378
rect 82 377 83 378
rect 81 377 82 378
rect 80 377 81 378
rect 79 377 80 378
rect 78 377 79 378
rect 77 377 78 378
rect 76 377 77 378
rect 75 377 76 378
rect 74 377 75 378
rect 73 377 74 378
rect 72 377 73 378
rect 71 377 72 378
rect 31 377 32 378
rect 30 377 31 378
rect 29 377 30 378
rect 28 377 29 378
rect 27 377 28 378
rect 26 377 27 378
rect 25 377 26 378
rect 24 377 25 378
rect 23 377 24 378
rect 22 377 23 378
rect 21 377 22 378
rect 20 377 21 378
rect 19 377 20 378
rect 18 377 19 378
rect 17 377 18 378
rect 146 378 147 379
rect 145 378 146 379
rect 144 378 145 379
rect 143 378 144 379
rect 142 378 143 379
rect 141 378 142 379
rect 140 378 141 379
rect 139 378 140 379
rect 127 378 128 379
rect 126 378 127 379
rect 125 378 126 379
rect 124 378 125 379
rect 123 378 124 379
rect 122 378 123 379
rect 121 378 122 379
rect 85 378 86 379
rect 84 378 85 379
rect 83 378 84 379
rect 82 378 83 379
rect 81 378 82 379
rect 80 378 81 379
rect 79 378 80 379
rect 78 378 79 379
rect 77 378 78 379
rect 76 378 77 379
rect 75 378 76 379
rect 74 378 75 379
rect 73 378 74 379
rect 72 378 73 379
rect 71 378 72 379
rect 31 378 32 379
rect 30 378 31 379
rect 29 378 30 379
rect 28 378 29 379
rect 27 378 28 379
rect 26 378 27 379
rect 25 378 26 379
rect 24 378 25 379
rect 23 378 24 379
rect 22 378 23 379
rect 21 378 22 379
rect 20 378 21 379
rect 19 378 20 379
rect 18 378 19 379
rect 17 378 18 379
rect 146 379 147 380
rect 145 379 146 380
rect 144 379 145 380
rect 143 379 144 380
rect 142 379 143 380
rect 141 379 142 380
rect 140 379 141 380
rect 125 379 126 380
rect 124 379 125 380
rect 123 379 124 380
rect 122 379 123 380
rect 121 379 122 380
rect 85 379 86 380
rect 84 379 85 380
rect 83 379 84 380
rect 82 379 83 380
rect 81 379 82 380
rect 80 379 81 380
rect 79 379 80 380
rect 78 379 79 380
rect 77 379 78 380
rect 76 379 77 380
rect 75 379 76 380
rect 74 379 75 380
rect 73 379 74 380
rect 72 379 73 380
rect 71 379 72 380
rect 31 379 32 380
rect 30 379 31 380
rect 29 379 30 380
rect 28 379 29 380
rect 27 379 28 380
rect 26 379 27 380
rect 25 379 26 380
rect 24 379 25 380
rect 23 379 24 380
rect 22 379 23 380
rect 21 379 22 380
rect 20 379 21 380
rect 19 379 20 380
rect 18 379 19 380
rect 17 379 18 380
rect 146 380 147 381
rect 145 380 146 381
rect 144 380 145 381
rect 143 380 144 381
rect 142 380 143 381
rect 124 380 125 381
rect 123 380 124 381
rect 122 380 123 381
rect 121 380 122 381
rect 85 380 86 381
rect 84 380 85 381
rect 83 380 84 381
rect 82 380 83 381
rect 81 380 82 381
rect 80 380 81 381
rect 79 380 80 381
rect 78 380 79 381
rect 77 380 78 381
rect 76 380 77 381
rect 75 380 76 381
rect 74 380 75 381
rect 73 380 74 381
rect 72 380 73 381
rect 71 380 72 381
rect 70 380 71 381
rect 32 380 33 381
rect 31 380 32 381
rect 30 380 31 381
rect 29 380 30 381
rect 28 380 29 381
rect 27 380 28 381
rect 26 380 27 381
rect 25 380 26 381
rect 24 380 25 381
rect 23 380 24 381
rect 22 380 23 381
rect 21 380 22 381
rect 20 380 21 381
rect 19 380 20 381
rect 18 380 19 381
rect 17 380 18 381
rect 146 381 147 382
rect 145 381 146 382
rect 144 381 145 382
rect 143 381 144 382
rect 123 381 124 382
rect 122 381 123 382
rect 121 381 122 382
rect 85 381 86 382
rect 84 381 85 382
rect 83 381 84 382
rect 82 381 83 382
rect 81 381 82 382
rect 80 381 81 382
rect 79 381 80 382
rect 78 381 79 382
rect 77 381 78 382
rect 76 381 77 382
rect 75 381 76 382
rect 74 381 75 382
rect 73 381 74 382
rect 72 381 73 382
rect 71 381 72 382
rect 70 381 71 382
rect 69 381 70 382
rect 33 381 34 382
rect 32 381 33 382
rect 31 381 32 382
rect 30 381 31 382
rect 29 381 30 382
rect 28 381 29 382
rect 27 381 28 382
rect 26 381 27 382
rect 25 381 26 382
rect 24 381 25 382
rect 23 381 24 382
rect 22 381 23 382
rect 21 381 22 382
rect 20 381 21 382
rect 19 381 20 382
rect 18 381 19 382
rect 17 381 18 382
rect 146 382 147 383
rect 145 382 146 383
rect 121 382 122 383
rect 85 382 86 383
rect 84 382 85 383
rect 83 382 84 383
rect 82 382 83 383
rect 81 382 82 383
rect 80 382 81 383
rect 79 382 80 383
rect 78 382 79 383
rect 77 382 78 383
rect 76 382 77 383
rect 75 382 76 383
rect 74 382 75 383
rect 73 382 74 383
rect 72 382 73 383
rect 71 382 72 383
rect 70 382 71 383
rect 69 382 70 383
rect 68 382 69 383
rect 67 382 68 383
rect 66 382 67 383
rect 35 382 36 383
rect 34 382 35 383
rect 33 382 34 383
rect 32 382 33 383
rect 31 382 32 383
rect 30 382 31 383
rect 29 382 30 383
rect 28 382 29 383
rect 27 382 28 383
rect 26 382 27 383
rect 25 382 26 383
rect 24 382 25 383
rect 23 382 24 383
rect 22 382 23 383
rect 21 382 22 383
rect 20 382 21 383
rect 19 382 20 383
rect 18 382 19 383
rect 17 382 18 383
rect 146 383 147 384
rect 84 383 85 384
rect 83 383 84 384
rect 82 383 83 384
rect 81 383 82 384
rect 80 383 81 384
rect 79 383 80 384
rect 78 383 79 384
rect 77 383 78 384
rect 76 383 77 384
rect 75 383 76 384
rect 74 383 75 384
rect 73 383 74 384
rect 72 383 73 384
rect 71 383 72 384
rect 70 383 71 384
rect 69 383 70 384
rect 68 383 69 384
rect 67 383 68 384
rect 66 383 67 384
rect 65 383 66 384
rect 64 383 65 384
rect 63 383 64 384
rect 62 383 63 384
rect 39 383 40 384
rect 38 383 39 384
rect 37 383 38 384
rect 36 383 37 384
rect 35 383 36 384
rect 34 383 35 384
rect 33 383 34 384
rect 32 383 33 384
rect 31 383 32 384
rect 30 383 31 384
rect 29 383 30 384
rect 28 383 29 384
rect 27 383 28 384
rect 26 383 27 384
rect 25 383 26 384
rect 24 383 25 384
rect 23 383 24 384
rect 22 383 23 384
rect 21 383 22 384
rect 20 383 21 384
rect 19 383 20 384
rect 18 383 19 384
rect 17 383 18 384
rect 84 384 85 385
rect 83 384 84 385
rect 82 384 83 385
rect 81 384 82 385
rect 80 384 81 385
rect 79 384 80 385
rect 78 384 79 385
rect 77 384 78 385
rect 76 384 77 385
rect 75 384 76 385
rect 74 384 75 385
rect 73 384 74 385
rect 72 384 73 385
rect 71 384 72 385
rect 70 384 71 385
rect 69 384 70 385
rect 68 384 69 385
rect 67 384 68 385
rect 66 384 67 385
rect 65 384 66 385
rect 64 384 65 385
rect 63 384 64 385
rect 62 384 63 385
rect 61 384 62 385
rect 60 384 61 385
rect 59 384 60 385
rect 58 384 59 385
rect 57 384 58 385
rect 56 384 57 385
rect 55 384 56 385
rect 54 384 55 385
rect 53 384 54 385
rect 52 384 53 385
rect 51 384 52 385
rect 50 384 51 385
rect 49 384 50 385
rect 48 384 49 385
rect 47 384 48 385
rect 46 384 47 385
rect 45 384 46 385
rect 44 384 45 385
rect 43 384 44 385
rect 42 384 43 385
rect 41 384 42 385
rect 40 384 41 385
rect 39 384 40 385
rect 38 384 39 385
rect 37 384 38 385
rect 36 384 37 385
rect 35 384 36 385
rect 34 384 35 385
rect 33 384 34 385
rect 32 384 33 385
rect 31 384 32 385
rect 30 384 31 385
rect 29 384 30 385
rect 28 384 29 385
rect 27 384 28 385
rect 26 384 27 385
rect 25 384 26 385
rect 24 384 25 385
rect 23 384 24 385
rect 22 384 23 385
rect 21 384 22 385
rect 20 384 21 385
rect 19 384 20 385
rect 18 384 19 385
rect 138 385 139 386
rect 137 385 138 386
rect 136 385 137 386
rect 84 385 85 386
rect 83 385 84 386
rect 82 385 83 386
rect 81 385 82 386
rect 80 385 81 386
rect 79 385 80 386
rect 78 385 79 386
rect 77 385 78 386
rect 76 385 77 386
rect 75 385 76 386
rect 74 385 75 386
rect 73 385 74 386
rect 72 385 73 386
rect 71 385 72 386
rect 70 385 71 386
rect 69 385 70 386
rect 68 385 69 386
rect 67 385 68 386
rect 66 385 67 386
rect 65 385 66 386
rect 64 385 65 386
rect 63 385 64 386
rect 62 385 63 386
rect 61 385 62 386
rect 60 385 61 386
rect 59 385 60 386
rect 58 385 59 386
rect 57 385 58 386
rect 56 385 57 386
rect 55 385 56 386
rect 54 385 55 386
rect 53 385 54 386
rect 52 385 53 386
rect 51 385 52 386
rect 50 385 51 386
rect 49 385 50 386
rect 48 385 49 386
rect 47 385 48 386
rect 46 385 47 386
rect 45 385 46 386
rect 44 385 45 386
rect 43 385 44 386
rect 42 385 43 386
rect 41 385 42 386
rect 40 385 41 386
rect 39 385 40 386
rect 38 385 39 386
rect 37 385 38 386
rect 36 385 37 386
rect 35 385 36 386
rect 34 385 35 386
rect 33 385 34 386
rect 32 385 33 386
rect 31 385 32 386
rect 30 385 31 386
rect 29 385 30 386
rect 28 385 29 386
rect 27 385 28 386
rect 26 385 27 386
rect 25 385 26 386
rect 24 385 25 386
rect 23 385 24 386
rect 22 385 23 386
rect 21 385 22 386
rect 20 385 21 386
rect 19 385 20 386
rect 18 385 19 386
rect 141 386 142 387
rect 140 386 141 387
rect 139 386 140 387
rect 138 386 139 387
rect 137 386 138 387
rect 136 386 137 387
rect 135 386 136 387
rect 134 386 135 387
rect 133 386 134 387
rect 84 386 85 387
rect 83 386 84 387
rect 82 386 83 387
rect 81 386 82 387
rect 80 386 81 387
rect 79 386 80 387
rect 78 386 79 387
rect 77 386 78 387
rect 76 386 77 387
rect 75 386 76 387
rect 74 386 75 387
rect 73 386 74 387
rect 72 386 73 387
rect 71 386 72 387
rect 70 386 71 387
rect 69 386 70 387
rect 68 386 69 387
rect 67 386 68 387
rect 66 386 67 387
rect 65 386 66 387
rect 64 386 65 387
rect 63 386 64 387
rect 62 386 63 387
rect 61 386 62 387
rect 60 386 61 387
rect 59 386 60 387
rect 58 386 59 387
rect 57 386 58 387
rect 56 386 57 387
rect 55 386 56 387
rect 54 386 55 387
rect 53 386 54 387
rect 52 386 53 387
rect 51 386 52 387
rect 50 386 51 387
rect 49 386 50 387
rect 48 386 49 387
rect 47 386 48 387
rect 46 386 47 387
rect 45 386 46 387
rect 44 386 45 387
rect 43 386 44 387
rect 42 386 43 387
rect 41 386 42 387
rect 40 386 41 387
rect 39 386 40 387
rect 38 386 39 387
rect 37 386 38 387
rect 36 386 37 387
rect 35 386 36 387
rect 34 386 35 387
rect 33 386 34 387
rect 32 386 33 387
rect 31 386 32 387
rect 30 386 31 387
rect 29 386 30 387
rect 28 386 29 387
rect 27 386 28 387
rect 26 386 27 387
rect 25 386 26 387
rect 24 386 25 387
rect 23 386 24 387
rect 22 386 23 387
rect 21 386 22 387
rect 20 386 21 387
rect 19 386 20 387
rect 18 386 19 387
rect 143 387 144 388
rect 142 387 143 388
rect 141 387 142 388
rect 140 387 141 388
rect 139 387 140 388
rect 138 387 139 388
rect 137 387 138 388
rect 136 387 137 388
rect 135 387 136 388
rect 134 387 135 388
rect 133 387 134 388
rect 132 387 133 388
rect 131 387 132 388
rect 83 387 84 388
rect 82 387 83 388
rect 81 387 82 388
rect 80 387 81 388
rect 79 387 80 388
rect 78 387 79 388
rect 77 387 78 388
rect 76 387 77 388
rect 75 387 76 388
rect 74 387 75 388
rect 73 387 74 388
rect 72 387 73 388
rect 71 387 72 388
rect 70 387 71 388
rect 69 387 70 388
rect 68 387 69 388
rect 67 387 68 388
rect 66 387 67 388
rect 65 387 66 388
rect 64 387 65 388
rect 63 387 64 388
rect 62 387 63 388
rect 61 387 62 388
rect 60 387 61 388
rect 59 387 60 388
rect 58 387 59 388
rect 57 387 58 388
rect 56 387 57 388
rect 55 387 56 388
rect 54 387 55 388
rect 53 387 54 388
rect 52 387 53 388
rect 51 387 52 388
rect 50 387 51 388
rect 49 387 50 388
rect 48 387 49 388
rect 47 387 48 388
rect 46 387 47 388
rect 45 387 46 388
rect 44 387 45 388
rect 43 387 44 388
rect 42 387 43 388
rect 41 387 42 388
rect 40 387 41 388
rect 39 387 40 388
rect 38 387 39 388
rect 37 387 38 388
rect 36 387 37 388
rect 35 387 36 388
rect 34 387 35 388
rect 33 387 34 388
rect 32 387 33 388
rect 31 387 32 388
rect 30 387 31 388
rect 29 387 30 388
rect 28 387 29 388
rect 27 387 28 388
rect 26 387 27 388
rect 25 387 26 388
rect 24 387 25 388
rect 23 387 24 388
rect 22 387 23 388
rect 21 387 22 388
rect 20 387 21 388
rect 19 387 20 388
rect 18 387 19 388
rect 144 388 145 389
rect 143 388 144 389
rect 142 388 143 389
rect 141 388 142 389
rect 140 388 141 389
rect 139 388 140 389
rect 138 388 139 389
rect 137 388 138 389
rect 136 388 137 389
rect 135 388 136 389
rect 134 388 135 389
rect 133 388 134 389
rect 132 388 133 389
rect 131 388 132 389
rect 130 388 131 389
rect 83 388 84 389
rect 82 388 83 389
rect 81 388 82 389
rect 80 388 81 389
rect 79 388 80 389
rect 78 388 79 389
rect 77 388 78 389
rect 76 388 77 389
rect 75 388 76 389
rect 74 388 75 389
rect 73 388 74 389
rect 72 388 73 389
rect 71 388 72 389
rect 70 388 71 389
rect 69 388 70 389
rect 68 388 69 389
rect 67 388 68 389
rect 66 388 67 389
rect 65 388 66 389
rect 64 388 65 389
rect 63 388 64 389
rect 62 388 63 389
rect 61 388 62 389
rect 60 388 61 389
rect 59 388 60 389
rect 58 388 59 389
rect 57 388 58 389
rect 56 388 57 389
rect 55 388 56 389
rect 54 388 55 389
rect 53 388 54 389
rect 52 388 53 389
rect 51 388 52 389
rect 50 388 51 389
rect 49 388 50 389
rect 48 388 49 389
rect 47 388 48 389
rect 46 388 47 389
rect 45 388 46 389
rect 44 388 45 389
rect 43 388 44 389
rect 42 388 43 389
rect 41 388 42 389
rect 40 388 41 389
rect 39 388 40 389
rect 38 388 39 389
rect 37 388 38 389
rect 36 388 37 389
rect 35 388 36 389
rect 34 388 35 389
rect 33 388 34 389
rect 32 388 33 389
rect 31 388 32 389
rect 30 388 31 389
rect 29 388 30 389
rect 28 388 29 389
rect 27 388 28 389
rect 26 388 27 389
rect 25 388 26 389
rect 24 388 25 389
rect 23 388 24 389
rect 22 388 23 389
rect 21 388 22 389
rect 20 388 21 389
rect 19 388 20 389
rect 145 389 146 390
rect 144 389 145 390
rect 143 389 144 390
rect 142 389 143 390
rect 141 389 142 390
rect 140 389 141 390
rect 139 389 140 390
rect 138 389 139 390
rect 137 389 138 390
rect 136 389 137 390
rect 135 389 136 390
rect 134 389 135 390
rect 133 389 134 390
rect 132 389 133 390
rect 131 389 132 390
rect 130 389 131 390
rect 129 389 130 390
rect 83 389 84 390
rect 82 389 83 390
rect 81 389 82 390
rect 80 389 81 390
rect 79 389 80 390
rect 78 389 79 390
rect 77 389 78 390
rect 76 389 77 390
rect 75 389 76 390
rect 74 389 75 390
rect 73 389 74 390
rect 72 389 73 390
rect 71 389 72 390
rect 70 389 71 390
rect 69 389 70 390
rect 68 389 69 390
rect 67 389 68 390
rect 66 389 67 390
rect 65 389 66 390
rect 64 389 65 390
rect 63 389 64 390
rect 62 389 63 390
rect 61 389 62 390
rect 60 389 61 390
rect 59 389 60 390
rect 58 389 59 390
rect 57 389 58 390
rect 56 389 57 390
rect 55 389 56 390
rect 54 389 55 390
rect 53 389 54 390
rect 52 389 53 390
rect 51 389 52 390
rect 50 389 51 390
rect 49 389 50 390
rect 48 389 49 390
rect 47 389 48 390
rect 46 389 47 390
rect 45 389 46 390
rect 44 389 45 390
rect 43 389 44 390
rect 42 389 43 390
rect 41 389 42 390
rect 40 389 41 390
rect 39 389 40 390
rect 38 389 39 390
rect 37 389 38 390
rect 36 389 37 390
rect 35 389 36 390
rect 34 389 35 390
rect 33 389 34 390
rect 32 389 33 390
rect 31 389 32 390
rect 30 389 31 390
rect 29 389 30 390
rect 28 389 29 390
rect 27 389 28 390
rect 26 389 27 390
rect 25 389 26 390
rect 24 389 25 390
rect 23 389 24 390
rect 22 389 23 390
rect 21 389 22 390
rect 20 389 21 390
rect 19 389 20 390
rect 145 390 146 391
rect 144 390 145 391
rect 143 390 144 391
rect 142 390 143 391
rect 141 390 142 391
rect 140 390 141 391
rect 139 390 140 391
rect 138 390 139 391
rect 137 390 138 391
rect 136 390 137 391
rect 135 390 136 391
rect 134 390 135 391
rect 133 390 134 391
rect 132 390 133 391
rect 131 390 132 391
rect 130 390 131 391
rect 129 390 130 391
rect 82 390 83 391
rect 81 390 82 391
rect 80 390 81 391
rect 79 390 80 391
rect 78 390 79 391
rect 77 390 78 391
rect 76 390 77 391
rect 75 390 76 391
rect 74 390 75 391
rect 73 390 74 391
rect 72 390 73 391
rect 71 390 72 391
rect 70 390 71 391
rect 69 390 70 391
rect 68 390 69 391
rect 67 390 68 391
rect 66 390 67 391
rect 65 390 66 391
rect 64 390 65 391
rect 63 390 64 391
rect 62 390 63 391
rect 61 390 62 391
rect 60 390 61 391
rect 59 390 60 391
rect 58 390 59 391
rect 57 390 58 391
rect 56 390 57 391
rect 55 390 56 391
rect 54 390 55 391
rect 53 390 54 391
rect 52 390 53 391
rect 51 390 52 391
rect 50 390 51 391
rect 49 390 50 391
rect 48 390 49 391
rect 47 390 48 391
rect 46 390 47 391
rect 45 390 46 391
rect 44 390 45 391
rect 43 390 44 391
rect 42 390 43 391
rect 41 390 42 391
rect 40 390 41 391
rect 39 390 40 391
rect 38 390 39 391
rect 37 390 38 391
rect 36 390 37 391
rect 35 390 36 391
rect 34 390 35 391
rect 33 390 34 391
rect 32 390 33 391
rect 31 390 32 391
rect 30 390 31 391
rect 29 390 30 391
rect 28 390 29 391
rect 27 390 28 391
rect 26 390 27 391
rect 25 390 26 391
rect 24 390 25 391
rect 23 390 24 391
rect 22 390 23 391
rect 21 390 22 391
rect 20 390 21 391
rect 19 390 20 391
rect 145 391 146 392
rect 144 391 145 392
rect 143 391 144 392
rect 142 391 143 392
rect 141 391 142 392
rect 140 391 141 392
rect 134 391 135 392
rect 133 391 134 392
rect 132 391 133 392
rect 131 391 132 392
rect 130 391 131 392
rect 129 391 130 392
rect 81 391 82 392
rect 80 391 81 392
rect 79 391 80 392
rect 78 391 79 392
rect 77 391 78 392
rect 76 391 77 392
rect 75 391 76 392
rect 74 391 75 392
rect 73 391 74 392
rect 72 391 73 392
rect 71 391 72 392
rect 70 391 71 392
rect 69 391 70 392
rect 68 391 69 392
rect 67 391 68 392
rect 66 391 67 392
rect 65 391 66 392
rect 64 391 65 392
rect 63 391 64 392
rect 62 391 63 392
rect 61 391 62 392
rect 60 391 61 392
rect 59 391 60 392
rect 58 391 59 392
rect 57 391 58 392
rect 56 391 57 392
rect 55 391 56 392
rect 54 391 55 392
rect 53 391 54 392
rect 52 391 53 392
rect 51 391 52 392
rect 50 391 51 392
rect 49 391 50 392
rect 48 391 49 392
rect 47 391 48 392
rect 46 391 47 392
rect 45 391 46 392
rect 44 391 45 392
rect 43 391 44 392
rect 42 391 43 392
rect 41 391 42 392
rect 40 391 41 392
rect 39 391 40 392
rect 38 391 39 392
rect 37 391 38 392
rect 36 391 37 392
rect 35 391 36 392
rect 34 391 35 392
rect 33 391 34 392
rect 32 391 33 392
rect 31 391 32 392
rect 30 391 31 392
rect 29 391 30 392
rect 28 391 29 392
rect 27 391 28 392
rect 26 391 27 392
rect 25 391 26 392
rect 24 391 25 392
rect 23 391 24 392
rect 22 391 23 392
rect 21 391 22 392
rect 20 391 21 392
rect 146 392 147 393
rect 145 392 146 393
rect 144 392 145 393
rect 143 392 144 393
rect 142 392 143 393
rect 132 392 133 393
rect 131 392 132 393
rect 130 392 131 393
rect 129 392 130 393
rect 128 392 129 393
rect 81 392 82 393
rect 80 392 81 393
rect 79 392 80 393
rect 78 392 79 393
rect 77 392 78 393
rect 76 392 77 393
rect 75 392 76 393
rect 74 392 75 393
rect 73 392 74 393
rect 72 392 73 393
rect 71 392 72 393
rect 70 392 71 393
rect 69 392 70 393
rect 68 392 69 393
rect 67 392 68 393
rect 66 392 67 393
rect 65 392 66 393
rect 64 392 65 393
rect 63 392 64 393
rect 62 392 63 393
rect 61 392 62 393
rect 60 392 61 393
rect 59 392 60 393
rect 58 392 59 393
rect 57 392 58 393
rect 56 392 57 393
rect 55 392 56 393
rect 54 392 55 393
rect 53 392 54 393
rect 52 392 53 393
rect 51 392 52 393
rect 50 392 51 393
rect 49 392 50 393
rect 48 392 49 393
rect 47 392 48 393
rect 46 392 47 393
rect 45 392 46 393
rect 44 392 45 393
rect 43 392 44 393
rect 42 392 43 393
rect 41 392 42 393
rect 40 392 41 393
rect 39 392 40 393
rect 38 392 39 393
rect 37 392 38 393
rect 36 392 37 393
rect 35 392 36 393
rect 34 392 35 393
rect 33 392 34 393
rect 32 392 33 393
rect 31 392 32 393
rect 30 392 31 393
rect 29 392 30 393
rect 28 392 29 393
rect 27 392 28 393
rect 26 392 27 393
rect 25 392 26 393
rect 24 392 25 393
rect 23 392 24 393
rect 22 392 23 393
rect 21 392 22 393
rect 146 393 147 394
rect 145 393 146 394
rect 144 393 145 394
rect 143 393 144 394
rect 142 393 143 394
rect 132 393 133 394
rect 131 393 132 394
rect 130 393 131 394
rect 129 393 130 394
rect 128 393 129 394
rect 80 393 81 394
rect 79 393 80 394
rect 78 393 79 394
rect 77 393 78 394
rect 76 393 77 394
rect 75 393 76 394
rect 74 393 75 394
rect 73 393 74 394
rect 72 393 73 394
rect 71 393 72 394
rect 70 393 71 394
rect 69 393 70 394
rect 68 393 69 394
rect 67 393 68 394
rect 66 393 67 394
rect 65 393 66 394
rect 64 393 65 394
rect 63 393 64 394
rect 62 393 63 394
rect 61 393 62 394
rect 60 393 61 394
rect 59 393 60 394
rect 58 393 59 394
rect 57 393 58 394
rect 56 393 57 394
rect 55 393 56 394
rect 54 393 55 394
rect 53 393 54 394
rect 52 393 53 394
rect 51 393 52 394
rect 50 393 51 394
rect 49 393 50 394
rect 48 393 49 394
rect 47 393 48 394
rect 46 393 47 394
rect 45 393 46 394
rect 44 393 45 394
rect 43 393 44 394
rect 42 393 43 394
rect 41 393 42 394
rect 40 393 41 394
rect 39 393 40 394
rect 38 393 39 394
rect 37 393 38 394
rect 36 393 37 394
rect 35 393 36 394
rect 34 393 35 394
rect 33 393 34 394
rect 32 393 33 394
rect 31 393 32 394
rect 30 393 31 394
rect 29 393 30 394
rect 28 393 29 394
rect 27 393 28 394
rect 26 393 27 394
rect 25 393 26 394
rect 24 393 25 394
rect 23 393 24 394
rect 22 393 23 394
rect 21 393 22 394
rect 146 394 147 395
rect 145 394 146 395
rect 144 394 145 395
rect 143 394 144 395
rect 131 394 132 395
rect 130 394 131 395
rect 129 394 130 395
rect 128 394 129 395
rect 79 394 80 395
rect 78 394 79 395
rect 77 394 78 395
rect 76 394 77 395
rect 75 394 76 395
rect 74 394 75 395
rect 73 394 74 395
rect 72 394 73 395
rect 71 394 72 395
rect 70 394 71 395
rect 69 394 70 395
rect 68 394 69 395
rect 67 394 68 395
rect 66 394 67 395
rect 65 394 66 395
rect 64 394 65 395
rect 63 394 64 395
rect 62 394 63 395
rect 61 394 62 395
rect 60 394 61 395
rect 59 394 60 395
rect 58 394 59 395
rect 57 394 58 395
rect 56 394 57 395
rect 55 394 56 395
rect 54 394 55 395
rect 53 394 54 395
rect 52 394 53 395
rect 51 394 52 395
rect 50 394 51 395
rect 49 394 50 395
rect 48 394 49 395
rect 47 394 48 395
rect 46 394 47 395
rect 45 394 46 395
rect 44 394 45 395
rect 43 394 44 395
rect 42 394 43 395
rect 41 394 42 395
rect 40 394 41 395
rect 39 394 40 395
rect 38 394 39 395
rect 37 394 38 395
rect 36 394 37 395
rect 35 394 36 395
rect 34 394 35 395
rect 33 394 34 395
rect 32 394 33 395
rect 31 394 32 395
rect 30 394 31 395
rect 29 394 30 395
rect 28 394 29 395
rect 27 394 28 395
rect 26 394 27 395
rect 25 394 26 395
rect 24 394 25 395
rect 23 394 24 395
rect 22 394 23 395
rect 146 395 147 396
rect 145 395 146 396
rect 144 395 145 396
rect 143 395 144 396
rect 131 395 132 396
rect 130 395 131 396
rect 129 395 130 396
rect 128 395 129 396
rect 78 395 79 396
rect 77 395 78 396
rect 76 395 77 396
rect 75 395 76 396
rect 74 395 75 396
rect 73 395 74 396
rect 72 395 73 396
rect 71 395 72 396
rect 70 395 71 396
rect 69 395 70 396
rect 68 395 69 396
rect 67 395 68 396
rect 66 395 67 396
rect 65 395 66 396
rect 64 395 65 396
rect 63 395 64 396
rect 62 395 63 396
rect 61 395 62 396
rect 60 395 61 396
rect 59 395 60 396
rect 58 395 59 396
rect 57 395 58 396
rect 56 395 57 396
rect 55 395 56 396
rect 54 395 55 396
rect 53 395 54 396
rect 52 395 53 396
rect 51 395 52 396
rect 50 395 51 396
rect 49 395 50 396
rect 48 395 49 396
rect 47 395 48 396
rect 46 395 47 396
rect 45 395 46 396
rect 44 395 45 396
rect 43 395 44 396
rect 42 395 43 396
rect 41 395 42 396
rect 40 395 41 396
rect 39 395 40 396
rect 38 395 39 396
rect 37 395 38 396
rect 36 395 37 396
rect 35 395 36 396
rect 34 395 35 396
rect 33 395 34 396
rect 32 395 33 396
rect 31 395 32 396
rect 30 395 31 396
rect 29 395 30 396
rect 28 395 29 396
rect 27 395 28 396
rect 26 395 27 396
rect 25 395 26 396
rect 24 395 25 396
rect 23 395 24 396
rect 146 396 147 397
rect 145 396 146 397
rect 144 396 145 397
rect 143 396 144 397
rect 131 396 132 397
rect 130 396 131 397
rect 129 396 130 397
rect 128 396 129 397
rect 77 396 78 397
rect 76 396 77 397
rect 75 396 76 397
rect 74 396 75 397
rect 73 396 74 397
rect 72 396 73 397
rect 71 396 72 397
rect 70 396 71 397
rect 69 396 70 397
rect 68 396 69 397
rect 67 396 68 397
rect 66 396 67 397
rect 65 396 66 397
rect 64 396 65 397
rect 63 396 64 397
rect 62 396 63 397
rect 61 396 62 397
rect 60 396 61 397
rect 59 396 60 397
rect 58 396 59 397
rect 57 396 58 397
rect 56 396 57 397
rect 55 396 56 397
rect 54 396 55 397
rect 53 396 54 397
rect 52 396 53 397
rect 51 396 52 397
rect 50 396 51 397
rect 49 396 50 397
rect 48 396 49 397
rect 47 396 48 397
rect 46 396 47 397
rect 45 396 46 397
rect 44 396 45 397
rect 43 396 44 397
rect 42 396 43 397
rect 41 396 42 397
rect 40 396 41 397
rect 39 396 40 397
rect 38 396 39 397
rect 37 396 38 397
rect 36 396 37 397
rect 35 396 36 397
rect 34 396 35 397
rect 33 396 34 397
rect 32 396 33 397
rect 31 396 32 397
rect 30 396 31 397
rect 29 396 30 397
rect 28 396 29 397
rect 27 396 28 397
rect 26 396 27 397
rect 25 396 26 397
rect 24 396 25 397
rect 146 397 147 398
rect 145 397 146 398
rect 144 397 145 398
rect 143 397 144 398
rect 142 397 143 398
rect 132 397 133 398
rect 131 397 132 398
rect 130 397 131 398
rect 129 397 130 398
rect 128 397 129 398
rect 76 397 77 398
rect 75 397 76 398
rect 74 397 75 398
rect 73 397 74 398
rect 72 397 73 398
rect 71 397 72 398
rect 70 397 71 398
rect 69 397 70 398
rect 68 397 69 398
rect 67 397 68 398
rect 66 397 67 398
rect 65 397 66 398
rect 64 397 65 398
rect 63 397 64 398
rect 62 397 63 398
rect 61 397 62 398
rect 60 397 61 398
rect 59 397 60 398
rect 58 397 59 398
rect 57 397 58 398
rect 56 397 57 398
rect 55 397 56 398
rect 54 397 55 398
rect 53 397 54 398
rect 52 397 53 398
rect 51 397 52 398
rect 50 397 51 398
rect 49 397 50 398
rect 48 397 49 398
rect 47 397 48 398
rect 46 397 47 398
rect 45 397 46 398
rect 44 397 45 398
rect 43 397 44 398
rect 42 397 43 398
rect 41 397 42 398
rect 40 397 41 398
rect 39 397 40 398
rect 38 397 39 398
rect 37 397 38 398
rect 36 397 37 398
rect 35 397 36 398
rect 34 397 35 398
rect 33 397 34 398
rect 32 397 33 398
rect 31 397 32 398
rect 30 397 31 398
rect 29 397 30 398
rect 28 397 29 398
rect 27 397 28 398
rect 26 397 27 398
rect 25 397 26 398
rect 146 398 147 399
rect 145 398 146 399
rect 144 398 145 399
rect 143 398 144 399
rect 142 398 143 399
rect 141 398 142 399
rect 133 398 134 399
rect 132 398 133 399
rect 131 398 132 399
rect 130 398 131 399
rect 129 398 130 399
rect 128 398 129 399
rect 74 398 75 399
rect 73 398 74 399
rect 72 398 73 399
rect 71 398 72 399
rect 70 398 71 399
rect 69 398 70 399
rect 68 398 69 399
rect 67 398 68 399
rect 66 398 67 399
rect 65 398 66 399
rect 64 398 65 399
rect 63 398 64 399
rect 62 398 63 399
rect 61 398 62 399
rect 60 398 61 399
rect 59 398 60 399
rect 58 398 59 399
rect 57 398 58 399
rect 56 398 57 399
rect 55 398 56 399
rect 54 398 55 399
rect 53 398 54 399
rect 52 398 53 399
rect 51 398 52 399
rect 50 398 51 399
rect 49 398 50 399
rect 48 398 49 399
rect 47 398 48 399
rect 46 398 47 399
rect 45 398 46 399
rect 44 398 45 399
rect 43 398 44 399
rect 42 398 43 399
rect 41 398 42 399
rect 40 398 41 399
rect 39 398 40 399
rect 38 398 39 399
rect 37 398 38 399
rect 36 398 37 399
rect 35 398 36 399
rect 34 398 35 399
rect 33 398 34 399
rect 32 398 33 399
rect 31 398 32 399
rect 30 398 31 399
rect 29 398 30 399
rect 28 398 29 399
rect 27 398 28 399
rect 145 399 146 400
rect 144 399 145 400
rect 143 399 144 400
rect 142 399 143 400
rect 141 399 142 400
rect 140 399 141 400
rect 139 399 140 400
rect 135 399 136 400
rect 134 399 135 400
rect 133 399 134 400
rect 132 399 133 400
rect 131 399 132 400
rect 130 399 131 400
rect 129 399 130 400
rect 72 399 73 400
rect 71 399 72 400
rect 70 399 71 400
rect 69 399 70 400
rect 68 399 69 400
rect 67 399 68 400
rect 66 399 67 400
rect 65 399 66 400
rect 64 399 65 400
rect 63 399 64 400
rect 62 399 63 400
rect 61 399 62 400
rect 60 399 61 400
rect 59 399 60 400
rect 58 399 59 400
rect 57 399 58 400
rect 56 399 57 400
rect 55 399 56 400
rect 54 399 55 400
rect 53 399 54 400
rect 52 399 53 400
rect 51 399 52 400
rect 50 399 51 400
rect 49 399 50 400
rect 48 399 49 400
rect 47 399 48 400
rect 46 399 47 400
rect 45 399 46 400
rect 44 399 45 400
rect 43 399 44 400
rect 42 399 43 400
rect 41 399 42 400
rect 40 399 41 400
rect 39 399 40 400
rect 38 399 39 400
rect 37 399 38 400
rect 36 399 37 400
rect 35 399 36 400
rect 34 399 35 400
rect 33 399 34 400
rect 32 399 33 400
rect 31 399 32 400
rect 30 399 31 400
rect 29 399 30 400
rect 145 400 146 401
rect 144 400 145 401
rect 143 400 144 401
rect 142 400 143 401
rect 141 400 142 401
rect 140 400 141 401
rect 139 400 140 401
rect 138 400 139 401
rect 137 400 138 401
rect 136 400 137 401
rect 135 400 136 401
rect 134 400 135 401
rect 133 400 134 401
rect 132 400 133 401
rect 131 400 132 401
rect 130 400 131 401
rect 129 400 130 401
rect 70 400 71 401
rect 69 400 70 401
rect 68 400 69 401
rect 67 400 68 401
rect 66 400 67 401
rect 65 400 66 401
rect 64 400 65 401
rect 63 400 64 401
rect 62 400 63 401
rect 61 400 62 401
rect 60 400 61 401
rect 59 400 60 401
rect 58 400 59 401
rect 57 400 58 401
rect 56 400 57 401
rect 55 400 56 401
rect 54 400 55 401
rect 53 400 54 401
rect 52 400 53 401
rect 51 400 52 401
rect 50 400 51 401
rect 49 400 50 401
rect 48 400 49 401
rect 47 400 48 401
rect 46 400 47 401
rect 45 400 46 401
rect 44 400 45 401
rect 43 400 44 401
rect 42 400 43 401
rect 41 400 42 401
rect 40 400 41 401
rect 39 400 40 401
rect 38 400 39 401
rect 37 400 38 401
rect 36 400 37 401
rect 35 400 36 401
rect 34 400 35 401
rect 33 400 34 401
rect 32 400 33 401
rect 31 400 32 401
rect 144 401 145 402
rect 143 401 144 402
rect 142 401 143 402
rect 141 401 142 402
rect 140 401 141 402
rect 139 401 140 402
rect 138 401 139 402
rect 137 401 138 402
rect 136 401 137 402
rect 135 401 136 402
rect 134 401 135 402
rect 133 401 134 402
rect 132 401 133 402
rect 131 401 132 402
rect 130 401 131 402
rect 68 401 69 402
rect 67 401 68 402
rect 66 401 67 402
rect 65 401 66 402
rect 64 401 65 402
rect 63 401 64 402
rect 62 401 63 402
rect 61 401 62 402
rect 60 401 61 402
rect 59 401 60 402
rect 58 401 59 402
rect 57 401 58 402
rect 56 401 57 402
rect 55 401 56 402
rect 54 401 55 402
rect 53 401 54 402
rect 52 401 53 402
rect 51 401 52 402
rect 50 401 51 402
rect 49 401 50 402
rect 48 401 49 402
rect 47 401 48 402
rect 46 401 47 402
rect 45 401 46 402
rect 44 401 45 402
rect 43 401 44 402
rect 42 401 43 402
rect 41 401 42 402
rect 40 401 41 402
rect 39 401 40 402
rect 38 401 39 402
rect 37 401 38 402
rect 36 401 37 402
rect 35 401 36 402
rect 34 401 35 402
rect 33 401 34 402
rect 143 402 144 403
rect 142 402 143 403
rect 141 402 142 403
rect 140 402 141 403
rect 139 402 140 403
rect 138 402 139 403
rect 137 402 138 403
rect 136 402 137 403
rect 135 402 136 403
rect 134 402 135 403
rect 133 402 134 403
rect 132 402 133 403
rect 131 402 132 403
rect 130 402 131 403
rect 64 402 65 403
rect 63 402 64 403
rect 62 402 63 403
rect 61 402 62 403
rect 60 402 61 403
rect 59 402 60 403
rect 58 402 59 403
rect 57 402 58 403
rect 56 402 57 403
rect 55 402 56 403
rect 54 402 55 403
rect 53 402 54 403
rect 52 402 53 403
rect 51 402 52 403
rect 50 402 51 403
rect 49 402 50 403
rect 48 402 49 403
rect 47 402 48 403
rect 46 402 47 403
rect 45 402 46 403
rect 44 402 45 403
rect 43 402 44 403
rect 42 402 43 403
rect 41 402 42 403
rect 40 402 41 403
rect 39 402 40 403
rect 38 402 39 403
rect 37 402 38 403
rect 142 403 143 404
rect 141 403 142 404
rect 140 403 141 404
rect 139 403 140 404
rect 138 403 139 404
rect 137 403 138 404
rect 136 403 137 404
rect 135 403 136 404
rect 134 403 135 404
rect 133 403 134 404
rect 132 403 133 404
rect 57 403 58 404
rect 56 403 57 404
rect 55 403 56 404
rect 54 403 55 404
rect 53 403 54 404
rect 52 403 53 404
rect 51 403 52 404
rect 50 403 51 404
rect 49 403 50 404
rect 48 403 49 404
rect 47 403 48 404
rect 46 403 47 404
rect 45 403 46 404
rect 44 403 45 404
rect 140 404 141 405
rect 139 404 140 405
rect 138 404 139 405
rect 137 404 138 405
rect 136 404 137 405
rect 135 404 136 405
rect 134 404 135 405
rect 133 404 134 405
rect 140 408 141 409
rect 139 408 140 409
rect 138 408 139 409
rect 137 408 138 409
rect 136 408 137 409
rect 135 408 136 409
rect 134 408 135 409
rect 142 409 143 410
rect 141 409 142 410
rect 140 409 141 410
rect 139 409 140 410
rect 138 409 139 410
rect 137 409 138 410
rect 136 409 137 410
rect 135 409 136 410
rect 134 409 135 410
rect 133 409 134 410
rect 132 409 133 410
rect 143 410 144 411
rect 142 410 143 411
rect 141 410 142 411
rect 140 410 141 411
rect 139 410 140 411
rect 138 410 139 411
rect 137 410 138 411
rect 136 410 137 411
rect 135 410 136 411
rect 134 410 135 411
rect 133 410 134 411
rect 132 410 133 411
rect 131 410 132 411
rect 144 411 145 412
rect 143 411 144 412
rect 142 411 143 412
rect 141 411 142 412
rect 140 411 141 412
rect 139 411 140 412
rect 138 411 139 412
rect 137 411 138 412
rect 136 411 137 412
rect 135 411 136 412
rect 134 411 135 412
rect 133 411 134 412
rect 132 411 133 412
rect 131 411 132 412
rect 130 411 131 412
rect 84 411 85 412
rect 83 411 84 412
rect 82 411 83 412
rect 81 411 82 412
rect 80 411 81 412
rect 79 411 80 412
rect 78 411 79 412
rect 77 411 78 412
rect 76 411 77 412
rect 75 411 76 412
rect 74 411 75 412
rect 145 412 146 413
rect 144 412 145 413
rect 143 412 144 413
rect 142 412 143 413
rect 141 412 142 413
rect 140 412 141 413
rect 139 412 140 413
rect 138 412 139 413
rect 137 412 138 413
rect 136 412 137 413
rect 135 412 136 413
rect 134 412 135 413
rect 133 412 134 413
rect 132 412 133 413
rect 131 412 132 413
rect 130 412 131 413
rect 129 412 130 413
rect 84 412 85 413
rect 83 412 84 413
rect 82 412 83 413
rect 81 412 82 413
rect 80 412 81 413
rect 79 412 80 413
rect 78 412 79 413
rect 77 412 78 413
rect 76 412 77 413
rect 75 412 76 413
rect 74 412 75 413
rect 73 412 74 413
rect 72 412 73 413
rect 71 412 72 413
rect 70 412 71 413
rect 145 413 146 414
rect 144 413 145 414
rect 143 413 144 414
rect 142 413 143 414
rect 141 413 142 414
rect 140 413 141 414
rect 139 413 140 414
rect 138 413 139 414
rect 137 413 138 414
rect 136 413 137 414
rect 135 413 136 414
rect 134 413 135 414
rect 133 413 134 414
rect 132 413 133 414
rect 131 413 132 414
rect 130 413 131 414
rect 129 413 130 414
rect 84 413 85 414
rect 83 413 84 414
rect 82 413 83 414
rect 81 413 82 414
rect 80 413 81 414
rect 79 413 80 414
rect 78 413 79 414
rect 77 413 78 414
rect 76 413 77 414
rect 75 413 76 414
rect 74 413 75 414
rect 73 413 74 414
rect 72 413 73 414
rect 71 413 72 414
rect 70 413 71 414
rect 69 413 70 414
rect 68 413 69 414
rect 67 413 68 414
rect 146 414 147 415
rect 145 414 146 415
rect 144 414 145 415
rect 143 414 144 415
rect 142 414 143 415
rect 141 414 142 415
rect 133 414 134 415
rect 132 414 133 415
rect 131 414 132 415
rect 130 414 131 415
rect 129 414 130 415
rect 128 414 129 415
rect 84 414 85 415
rect 83 414 84 415
rect 82 414 83 415
rect 81 414 82 415
rect 80 414 81 415
rect 79 414 80 415
rect 78 414 79 415
rect 77 414 78 415
rect 76 414 77 415
rect 75 414 76 415
rect 74 414 75 415
rect 73 414 74 415
rect 72 414 73 415
rect 71 414 72 415
rect 70 414 71 415
rect 69 414 70 415
rect 68 414 69 415
rect 67 414 68 415
rect 66 414 67 415
rect 37 414 38 415
rect 36 414 37 415
rect 35 414 36 415
rect 34 414 35 415
rect 33 414 34 415
rect 32 414 33 415
rect 31 414 32 415
rect 30 414 31 415
rect 29 414 30 415
rect 28 414 29 415
rect 27 414 28 415
rect 26 414 27 415
rect 25 414 26 415
rect 24 414 25 415
rect 23 414 24 415
rect 22 414 23 415
rect 146 415 147 416
rect 145 415 146 416
rect 144 415 145 416
rect 143 415 144 416
rect 142 415 143 416
rect 132 415 133 416
rect 131 415 132 416
rect 130 415 131 416
rect 129 415 130 416
rect 128 415 129 416
rect 84 415 85 416
rect 83 415 84 416
rect 82 415 83 416
rect 81 415 82 416
rect 80 415 81 416
rect 79 415 80 416
rect 78 415 79 416
rect 77 415 78 416
rect 76 415 77 416
rect 75 415 76 416
rect 74 415 75 416
rect 73 415 74 416
rect 72 415 73 416
rect 71 415 72 416
rect 70 415 71 416
rect 69 415 70 416
rect 68 415 69 416
rect 67 415 68 416
rect 66 415 67 416
rect 65 415 66 416
rect 64 415 65 416
rect 36 415 37 416
rect 35 415 36 416
rect 34 415 35 416
rect 33 415 34 416
rect 32 415 33 416
rect 31 415 32 416
rect 30 415 31 416
rect 29 415 30 416
rect 28 415 29 416
rect 27 415 28 416
rect 26 415 27 416
rect 25 415 26 416
rect 24 415 25 416
rect 23 415 24 416
rect 22 415 23 416
rect 21 415 22 416
rect 146 416 147 417
rect 145 416 146 417
rect 144 416 145 417
rect 143 416 144 417
rect 142 416 143 417
rect 132 416 133 417
rect 131 416 132 417
rect 130 416 131 417
rect 129 416 130 417
rect 128 416 129 417
rect 84 416 85 417
rect 83 416 84 417
rect 82 416 83 417
rect 81 416 82 417
rect 80 416 81 417
rect 79 416 80 417
rect 78 416 79 417
rect 77 416 78 417
rect 76 416 77 417
rect 75 416 76 417
rect 74 416 75 417
rect 73 416 74 417
rect 72 416 73 417
rect 71 416 72 417
rect 70 416 71 417
rect 69 416 70 417
rect 68 416 69 417
rect 67 416 68 417
rect 66 416 67 417
rect 65 416 66 417
rect 64 416 65 417
rect 63 416 64 417
rect 36 416 37 417
rect 35 416 36 417
rect 34 416 35 417
rect 33 416 34 417
rect 32 416 33 417
rect 31 416 32 417
rect 30 416 31 417
rect 29 416 30 417
rect 28 416 29 417
rect 27 416 28 417
rect 26 416 27 417
rect 25 416 26 417
rect 24 416 25 417
rect 23 416 24 417
rect 22 416 23 417
rect 21 416 22 417
rect 146 417 147 418
rect 145 417 146 418
rect 144 417 145 418
rect 143 417 144 418
rect 131 417 132 418
rect 130 417 131 418
rect 129 417 130 418
rect 128 417 129 418
rect 84 417 85 418
rect 83 417 84 418
rect 82 417 83 418
rect 81 417 82 418
rect 80 417 81 418
rect 79 417 80 418
rect 78 417 79 418
rect 77 417 78 418
rect 76 417 77 418
rect 75 417 76 418
rect 74 417 75 418
rect 73 417 74 418
rect 72 417 73 418
rect 71 417 72 418
rect 70 417 71 418
rect 69 417 70 418
rect 68 417 69 418
rect 67 417 68 418
rect 66 417 67 418
rect 65 417 66 418
rect 64 417 65 418
rect 63 417 64 418
rect 62 417 63 418
rect 61 417 62 418
rect 35 417 36 418
rect 34 417 35 418
rect 33 417 34 418
rect 32 417 33 418
rect 31 417 32 418
rect 30 417 31 418
rect 29 417 30 418
rect 28 417 29 418
rect 27 417 28 418
rect 26 417 27 418
rect 25 417 26 418
rect 24 417 25 418
rect 23 417 24 418
rect 22 417 23 418
rect 21 417 22 418
rect 146 418 147 419
rect 145 418 146 419
rect 144 418 145 419
rect 143 418 144 419
rect 131 418 132 419
rect 130 418 131 419
rect 129 418 130 419
rect 128 418 129 419
rect 84 418 85 419
rect 83 418 84 419
rect 82 418 83 419
rect 81 418 82 419
rect 80 418 81 419
rect 79 418 80 419
rect 78 418 79 419
rect 77 418 78 419
rect 76 418 77 419
rect 75 418 76 419
rect 74 418 75 419
rect 73 418 74 419
rect 72 418 73 419
rect 71 418 72 419
rect 70 418 71 419
rect 69 418 70 419
rect 68 418 69 419
rect 67 418 68 419
rect 66 418 67 419
rect 65 418 66 419
rect 64 418 65 419
rect 63 418 64 419
rect 62 418 63 419
rect 61 418 62 419
rect 60 418 61 419
rect 35 418 36 419
rect 34 418 35 419
rect 33 418 34 419
rect 32 418 33 419
rect 31 418 32 419
rect 30 418 31 419
rect 29 418 30 419
rect 28 418 29 419
rect 27 418 28 419
rect 26 418 27 419
rect 25 418 26 419
rect 24 418 25 419
rect 23 418 24 419
rect 22 418 23 419
rect 21 418 22 419
rect 20 418 21 419
rect 146 419 147 420
rect 145 419 146 420
rect 144 419 145 420
rect 143 419 144 420
rect 142 419 143 420
rect 132 419 133 420
rect 131 419 132 420
rect 130 419 131 420
rect 129 419 130 420
rect 128 419 129 420
rect 84 419 85 420
rect 83 419 84 420
rect 82 419 83 420
rect 81 419 82 420
rect 80 419 81 420
rect 79 419 80 420
rect 78 419 79 420
rect 77 419 78 420
rect 76 419 77 420
rect 75 419 76 420
rect 74 419 75 420
rect 73 419 74 420
rect 72 419 73 420
rect 71 419 72 420
rect 70 419 71 420
rect 69 419 70 420
rect 68 419 69 420
rect 67 419 68 420
rect 66 419 67 420
rect 65 419 66 420
rect 64 419 65 420
rect 63 419 64 420
rect 62 419 63 420
rect 61 419 62 420
rect 60 419 61 420
rect 59 419 60 420
rect 34 419 35 420
rect 33 419 34 420
rect 32 419 33 420
rect 31 419 32 420
rect 30 419 31 420
rect 29 419 30 420
rect 28 419 29 420
rect 27 419 28 420
rect 26 419 27 420
rect 25 419 26 420
rect 24 419 25 420
rect 23 419 24 420
rect 22 419 23 420
rect 21 419 22 420
rect 20 419 21 420
rect 146 420 147 421
rect 145 420 146 421
rect 144 420 145 421
rect 143 420 144 421
rect 142 420 143 421
rect 132 420 133 421
rect 131 420 132 421
rect 130 420 131 421
rect 129 420 130 421
rect 128 420 129 421
rect 84 420 85 421
rect 83 420 84 421
rect 82 420 83 421
rect 81 420 82 421
rect 80 420 81 421
rect 79 420 80 421
rect 78 420 79 421
rect 77 420 78 421
rect 76 420 77 421
rect 75 420 76 421
rect 74 420 75 421
rect 73 420 74 421
rect 72 420 73 421
rect 71 420 72 421
rect 70 420 71 421
rect 69 420 70 421
rect 68 420 69 421
rect 67 420 68 421
rect 66 420 67 421
rect 65 420 66 421
rect 64 420 65 421
rect 63 420 64 421
rect 62 420 63 421
rect 61 420 62 421
rect 60 420 61 421
rect 59 420 60 421
rect 58 420 59 421
rect 34 420 35 421
rect 33 420 34 421
rect 32 420 33 421
rect 31 420 32 421
rect 30 420 31 421
rect 29 420 30 421
rect 28 420 29 421
rect 27 420 28 421
rect 26 420 27 421
rect 25 420 26 421
rect 24 420 25 421
rect 23 420 24 421
rect 22 420 23 421
rect 21 420 22 421
rect 20 420 21 421
rect 19 420 20 421
rect 146 421 147 422
rect 145 421 146 422
rect 144 421 145 422
rect 143 421 144 422
rect 142 421 143 422
rect 141 421 142 422
rect 133 421 134 422
rect 132 421 133 422
rect 131 421 132 422
rect 130 421 131 422
rect 129 421 130 422
rect 128 421 129 422
rect 84 421 85 422
rect 83 421 84 422
rect 82 421 83 422
rect 81 421 82 422
rect 80 421 81 422
rect 79 421 80 422
rect 78 421 79 422
rect 77 421 78 422
rect 76 421 77 422
rect 75 421 76 422
rect 74 421 75 422
rect 73 421 74 422
rect 72 421 73 422
rect 71 421 72 422
rect 70 421 71 422
rect 69 421 70 422
rect 68 421 69 422
rect 67 421 68 422
rect 66 421 67 422
rect 65 421 66 422
rect 64 421 65 422
rect 63 421 64 422
rect 62 421 63 422
rect 61 421 62 422
rect 60 421 61 422
rect 59 421 60 422
rect 58 421 59 422
rect 33 421 34 422
rect 32 421 33 422
rect 31 421 32 422
rect 30 421 31 422
rect 29 421 30 422
rect 28 421 29 422
rect 27 421 28 422
rect 26 421 27 422
rect 25 421 26 422
rect 24 421 25 422
rect 23 421 24 422
rect 22 421 23 422
rect 21 421 22 422
rect 20 421 21 422
rect 19 421 20 422
rect 145 422 146 423
rect 144 422 145 423
rect 143 422 144 423
rect 142 422 143 423
rect 141 422 142 423
rect 140 422 141 423
rect 139 422 140 423
rect 138 422 139 423
rect 137 422 138 423
rect 136 422 137 423
rect 135 422 136 423
rect 134 422 135 423
rect 133 422 134 423
rect 132 422 133 423
rect 131 422 132 423
rect 130 422 131 423
rect 129 422 130 423
rect 84 422 85 423
rect 83 422 84 423
rect 82 422 83 423
rect 81 422 82 423
rect 80 422 81 423
rect 79 422 80 423
rect 78 422 79 423
rect 77 422 78 423
rect 76 422 77 423
rect 75 422 76 423
rect 74 422 75 423
rect 73 422 74 423
rect 72 422 73 423
rect 71 422 72 423
rect 70 422 71 423
rect 69 422 70 423
rect 68 422 69 423
rect 67 422 68 423
rect 66 422 67 423
rect 65 422 66 423
rect 64 422 65 423
rect 63 422 64 423
rect 62 422 63 423
rect 61 422 62 423
rect 60 422 61 423
rect 59 422 60 423
rect 58 422 59 423
rect 57 422 58 423
rect 33 422 34 423
rect 32 422 33 423
rect 31 422 32 423
rect 30 422 31 423
rect 29 422 30 423
rect 28 422 29 423
rect 27 422 28 423
rect 26 422 27 423
rect 25 422 26 423
rect 24 422 25 423
rect 23 422 24 423
rect 22 422 23 423
rect 21 422 22 423
rect 20 422 21 423
rect 19 422 20 423
rect 145 423 146 424
rect 144 423 145 424
rect 143 423 144 424
rect 142 423 143 424
rect 141 423 142 424
rect 140 423 141 424
rect 139 423 140 424
rect 138 423 139 424
rect 137 423 138 424
rect 136 423 137 424
rect 135 423 136 424
rect 134 423 135 424
rect 133 423 134 424
rect 132 423 133 424
rect 131 423 132 424
rect 130 423 131 424
rect 129 423 130 424
rect 84 423 85 424
rect 83 423 84 424
rect 82 423 83 424
rect 81 423 82 424
rect 80 423 81 424
rect 79 423 80 424
rect 78 423 79 424
rect 77 423 78 424
rect 76 423 77 424
rect 75 423 76 424
rect 74 423 75 424
rect 73 423 74 424
rect 72 423 73 424
rect 71 423 72 424
rect 70 423 71 424
rect 69 423 70 424
rect 68 423 69 424
rect 67 423 68 424
rect 66 423 67 424
rect 65 423 66 424
rect 64 423 65 424
rect 63 423 64 424
rect 62 423 63 424
rect 61 423 62 424
rect 60 423 61 424
rect 59 423 60 424
rect 58 423 59 424
rect 57 423 58 424
rect 56 423 57 424
rect 33 423 34 424
rect 32 423 33 424
rect 31 423 32 424
rect 30 423 31 424
rect 29 423 30 424
rect 28 423 29 424
rect 27 423 28 424
rect 26 423 27 424
rect 25 423 26 424
rect 24 423 25 424
rect 23 423 24 424
rect 22 423 23 424
rect 21 423 22 424
rect 20 423 21 424
rect 19 423 20 424
rect 18 423 19 424
rect 144 424 145 425
rect 143 424 144 425
rect 142 424 143 425
rect 141 424 142 425
rect 140 424 141 425
rect 139 424 140 425
rect 138 424 139 425
rect 137 424 138 425
rect 136 424 137 425
rect 135 424 136 425
rect 134 424 135 425
rect 133 424 134 425
rect 132 424 133 425
rect 131 424 132 425
rect 130 424 131 425
rect 84 424 85 425
rect 83 424 84 425
rect 82 424 83 425
rect 81 424 82 425
rect 80 424 81 425
rect 79 424 80 425
rect 78 424 79 425
rect 77 424 78 425
rect 76 424 77 425
rect 75 424 76 425
rect 74 424 75 425
rect 73 424 74 425
rect 72 424 73 425
rect 71 424 72 425
rect 70 424 71 425
rect 69 424 70 425
rect 68 424 69 425
rect 67 424 68 425
rect 66 424 67 425
rect 65 424 66 425
rect 64 424 65 425
rect 63 424 64 425
rect 62 424 63 425
rect 61 424 62 425
rect 60 424 61 425
rect 59 424 60 425
rect 58 424 59 425
rect 57 424 58 425
rect 56 424 57 425
rect 55 424 56 425
rect 33 424 34 425
rect 32 424 33 425
rect 31 424 32 425
rect 30 424 31 425
rect 29 424 30 425
rect 28 424 29 425
rect 27 424 28 425
rect 26 424 27 425
rect 25 424 26 425
rect 24 424 25 425
rect 23 424 24 425
rect 22 424 23 425
rect 21 424 22 425
rect 20 424 21 425
rect 19 424 20 425
rect 18 424 19 425
rect 143 425 144 426
rect 142 425 143 426
rect 141 425 142 426
rect 140 425 141 426
rect 139 425 140 426
rect 138 425 139 426
rect 137 425 138 426
rect 136 425 137 426
rect 135 425 136 426
rect 134 425 135 426
rect 133 425 134 426
rect 132 425 133 426
rect 131 425 132 426
rect 84 425 85 426
rect 83 425 84 426
rect 82 425 83 426
rect 81 425 82 426
rect 80 425 81 426
rect 79 425 80 426
rect 78 425 79 426
rect 77 425 78 426
rect 76 425 77 426
rect 75 425 76 426
rect 74 425 75 426
rect 73 425 74 426
rect 72 425 73 426
rect 71 425 72 426
rect 70 425 71 426
rect 69 425 70 426
rect 68 425 69 426
rect 67 425 68 426
rect 66 425 67 426
rect 65 425 66 426
rect 64 425 65 426
rect 63 425 64 426
rect 62 425 63 426
rect 61 425 62 426
rect 60 425 61 426
rect 59 425 60 426
rect 58 425 59 426
rect 57 425 58 426
rect 56 425 57 426
rect 55 425 56 426
rect 54 425 55 426
rect 32 425 33 426
rect 31 425 32 426
rect 30 425 31 426
rect 29 425 30 426
rect 28 425 29 426
rect 27 425 28 426
rect 26 425 27 426
rect 25 425 26 426
rect 24 425 25 426
rect 23 425 24 426
rect 22 425 23 426
rect 21 425 22 426
rect 20 425 21 426
rect 19 425 20 426
rect 18 425 19 426
rect 142 426 143 427
rect 141 426 142 427
rect 140 426 141 427
rect 139 426 140 427
rect 138 426 139 427
rect 137 426 138 427
rect 136 426 137 427
rect 135 426 136 427
rect 134 426 135 427
rect 133 426 134 427
rect 132 426 133 427
rect 84 426 85 427
rect 83 426 84 427
rect 82 426 83 427
rect 81 426 82 427
rect 80 426 81 427
rect 79 426 80 427
rect 78 426 79 427
rect 77 426 78 427
rect 76 426 77 427
rect 75 426 76 427
rect 74 426 75 427
rect 73 426 74 427
rect 72 426 73 427
rect 71 426 72 427
rect 70 426 71 427
rect 69 426 70 427
rect 68 426 69 427
rect 67 426 68 427
rect 66 426 67 427
rect 65 426 66 427
rect 64 426 65 427
rect 63 426 64 427
rect 62 426 63 427
rect 61 426 62 427
rect 60 426 61 427
rect 59 426 60 427
rect 58 426 59 427
rect 57 426 58 427
rect 56 426 57 427
rect 55 426 56 427
rect 54 426 55 427
rect 53 426 54 427
rect 32 426 33 427
rect 31 426 32 427
rect 30 426 31 427
rect 29 426 30 427
rect 28 426 29 427
rect 27 426 28 427
rect 26 426 27 427
rect 25 426 26 427
rect 24 426 25 427
rect 23 426 24 427
rect 22 426 23 427
rect 21 426 22 427
rect 20 426 21 427
rect 19 426 20 427
rect 18 426 19 427
rect 139 427 140 428
rect 138 427 139 428
rect 137 427 138 428
rect 136 427 137 428
rect 135 427 136 428
rect 134 427 135 428
rect 84 427 85 428
rect 83 427 84 428
rect 82 427 83 428
rect 81 427 82 428
rect 80 427 81 428
rect 79 427 80 428
rect 78 427 79 428
rect 77 427 78 428
rect 76 427 77 428
rect 75 427 76 428
rect 74 427 75 428
rect 73 427 74 428
rect 72 427 73 428
rect 71 427 72 428
rect 70 427 71 428
rect 69 427 70 428
rect 68 427 69 428
rect 67 427 68 428
rect 66 427 67 428
rect 65 427 66 428
rect 64 427 65 428
rect 63 427 64 428
rect 62 427 63 428
rect 61 427 62 428
rect 60 427 61 428
rect 59 427 60 428
rect 58 427 59 428
rect 57 427 58 428
rect 56 427 57 428
rect 55 427 56 428
rect 54 427 55 428
rect 53 427 54 428
rect 32 427 33 428
rect 31 427 32 428
rect 30 427 31 428
rect 29 427 30 428
rect 28 427 29 428
rect 27 427 28 428
rect 26 427 27 428
rect 25 427 26 428
rect 24 427 25 428
rect 23 427 24 428
rect 22 427 23 428
rect 21 427 22 428
rect 20 427 21 428
rect 19 427 20 428
rect 18 427 19 428
rect 84 428 85 429
rect 83 428 84 429
rect 82 428 83 429
rect 81 428 82 429
rect 80 428 81 429
rect 79 428 80 429
rect 78 428 79 429
rect 77 428 78 429
rect 76 428 77 429
rect 75 428 76 429
rect 74 428 75 429
rect 73 428 74 429
rect 72 428 73 429
rect 71 428 72 429
rect 70 428 71 429
rect 69 428 70 429
rect 68 428 69 429
rect 67 428 68 429
rect 66 428 67 429
rect 65 428 66 429
rect 64 428 65 429
rect 63 428 64 429
rect 62 428 63 429
rect 61 428 62 429
rect 60 428 61 429
rect 59 428 60 429
rect 58 428 59 429
rect 57 428 58 429
rect 56 428 57 429
rect 55 428 56 429
rect 54 428 55 429
rect 53 428 54 429
rect 52 428 53 429
rect 32 428 33 429
rect 31 428 32 429
rect 30 428 31 429
rect 29 428 30 429
rect 28 428 29 429
rect 27 428 28 429
rect 26 428 27 429
rect 25 428 26 429
rect 24 428 25 429
rect 23 428 24 429
rect 22 428 23 429
rect 21 428 22 429
rect 20 428 21 429
rect 19 428 20 429
rect 18 428 19 429
rect 84 429 85 430
rect 83 429 84 430
rect 82 429 83 430
rect 81 429 82 430
rect 80 429 81 430
rect 79 429 80 430
rect 78 429 79 430
rect 77 429 78 430
rect 76 429 77 430
rect 75 429 76 430
rect 74 429 75 430
rect 73 429 74 430
rect 72 429 73 430
rect 71 429 72 430
rect 70 429 71 430
rect 69 429 70 430
rect 68 429 69 430
rect 67 429 68 430
rect 66 429 67 430
rect 65 429 66 430
rect 64 429 65 430
rect 63 429 64 430
rect 62 429 63 430
rect 61 429 62 430
rect 60 429 61 430
rect 59 429 60 430
rect 58 429 59 430
rect 57 429 58 430
rect 56 429 57 430
rect 55 429 56 430
rect 54 429 55 430
rect 53 429 54 430
rect 52 429 53 430
rect 51 429 52 430
rect 32 429 33 430
rect 31 429 32 430
rect 30 429 31 430
rect 29 429 30 430
rect 28 429 29 430
rect 27 429 28 430
rect 26 429 27 430
rect 25 429 26 430
rect 24 429 25 430
rect 23 429 24 430
rect 22 429 23 430
rect 21 429 22 430
rect 20 429 21 430
rect 19 429 20 430
rect 18 429 19 430
rect 17 429 18 430
rect 84 430 85 431
rect 83 430 84 431
rect 82 430 83 431
rect 81 430 82 431
rect 80 430 81 431
rect 79 430 80 431
rect 78 430 79 431
rect 77 430 78 431
rect 76 430 77 431
rect 75 430 76 431
rect 74 430 75 431
rect 73 430 74 431
rect 72 430 73 431
rect 71 430 72 431
rect 70 430 71 431
rect 69 430 70 431
rect 68 430 69 431
rect 67 430 68 431
rect 66 430 67 431
rect 65 430 66 431
rect 64 430 65 431
rect 63 430 64 431
rect 62 430 63 431
rect 61 430 62 431
rect 60 430 61 431
rect 59 430 60 431
rect 58 430 59 431
rect 57 430 58 431
rect 56 430 57 431
rect 55 430 56 431
rect 54 430 55 431
rect 53 430 54 431
rect 52 430 53 431
rect 51 430 52 431
rect 50 430 51 431
rect 32 430 33 431
rect 31 430 32 431
rect 30 430 31 431
rect 29 430 30 431
rect 28 430 29 431
rect 27 430 28 431
rect 26 430 27 431
rect 25 430 26 431
rect 24 430 25 431
rect 23 430 24 431
rect 22 430 23 431
rect 21 430 22 431
rect 20 430 21 431
rect 19 430 20 431
rect 18 430 19 431
rect 17 430 18 431
rect 84 431 85 432
rect 83 431 84 432
rect 82 431 83 432
rect 81 431 82 432
rect 80 431 81 432
rect 79 431 80 432
rect 78 431 79 432
rect 77 431 78 432
rect 76 431 77 432
rect 75 431 76 432
rect 74 431 75 432
rect 73 431 74 432
rect 72 431 73 432
rect 71 431 72 432
rect 70 431 71 432
rect 69 431 70 432
rect 68 431 69 432
rect 67 431 68 432
rect 66 431 67 432
rect 65 431 66 432
rect 64 431 65 432
rect 63 431 64 432
rect 62 431 63 432
rect 61 431 62 432
rect 60 431 61 432
rect 59 431 60 432
rect 58 431 59 432
rect 57 431 58 432
rect 56 431 57 432
rect 55 431 56 432
rect 54 431 55 432
rect 53 431 54 432
rect 52 431 53 432
rect 51 431 52 432
rect 50 431 51 432
rect 49 431 50 432
rect 32 431 33 432
rect 31 431 32 432
rect 30 431 31 432
rect 29 431 30 432
rect 28 431 29 432
rect 27 431 28 432
rect 26 431 27 432
rect 25 431 26 432
rect 24 431 25 432
rect 23 431 24 432
rect 22 431 23 432
rect 21 431 22 432
rect 20 431 21 432
rect 19 431 20 432
rect 18 431 19 432
rect 17 431 18 432
rect 146 432 147 433
rect 145 432 146 433
rect 144 432 145 433
rect 143 432 144 433
rect 142 432 143 433
rect 141 432 142 433
rect 140 432 141 433
rect 139 432 140 433
rect 138 432 139 433
rect 137 432 138 433
rect 136 432 137 433
rect 135 432 136 433
rect 134 432 135 433
rect 133 432 134 433
rect 132 432 133 433
rect 131 432 132 433
rect 130 432 131 433
rect 129 432 130 433
rect 128 432 129 433
rect 127 432 128 433
rect 126 432 127 433
rect 125 432 126 433
rect 124 432 125 433
rect 123 432 124 433
rect 122 432 123 433
rect 121 432 122 433
rect 120 432 121 433
rect 119 432 120 433
rect 84 432 85 433
rect 83 432 84 433
rect 82 432 83 433
rect 81 432 82 433
rect 80 432 81 433
rect 79 432 80 433
rect 78 432 79 433
rect 77 432 78 433
rect 76 432 77 433
rect 75 432 76 433
rect 74 432 75 433
rect 73 432 74 433
rect 72 432 73 433
rect 71 432 72 433
rect 70 432 71 433
rect 69 432 70 433
rect 67 432 68 433
rect 66 432 67 433
rect 65 432 66 433
rect 64 432 65 433
rect 63 432 64 433
rect 62 432 63 433
rect 61 432 62 433
rect 60 432 61 433
rect 59 432 60 433
rect 58 432 59 433
rect 57 432 58 433
rect 56 432 57 433
rect 55 432 56 433
rect 54 432 55 433
rect 53 432 54 433
rect 52 432 53 433
rect 51 432 52 433
rect 50 432 51 433
rect 49 432 50 433
rect 32 432 33 433
rect 31 432 32 433
rect 30 432 31 433
rect 29 432 30 433
rect 28 432 29 433
rect 27 432 28 433
rect 26 432 27 433
rect 25 432 26 433
rect 24 432 25 433
rect 23 432 24 433
rect 22 432 23 433
rect 21 432 22 433
rect 20 432 21 433
rect 19 432 20 433
rect 18 432 19 433
rect 17 432 18 433
rect 146 433 147 434
rect 145 433 146 434
rect 144 433 145 434
rect 143 433 144 434
rect 142 433 143 434
rect 141 433 142 434
rect 140 433 141 434
rect 139 433 140 434
rect 138 433 139 434
rect 137 433 138 434
rect 136 433 137 434
rect 135 433 136 434
rect 134 433 135 434
rect 133 433 134 434
rect 132 433 133 434
rect 131 433 132 434
rect 130 433 131 434
rect 129 433 130 434
rect 128 433 129 434
rect 127 433 128 434
rect 126 433 127 434
rect 125 433 126 434
rect 124 433 125 434
rect 123 433 124 434
rect 122 433 123 434
rect 121 433 122 434
rect 120 433 121 434
rect 119 433 120 434
rect 84 433 85 434
rect 83 433 84 434
rect 82 433 83 434
rect 81 433 82 434
rect 80 433 81 434
rect 79 433 80 434
rect 78 433 79 434
rect 77 433 78 434
rect 76 433 77 434
rect 75 433 76 434
rect 74 433 75 434
rect 73 433 74 434
rect 72 433 73 434
rect 71 433 72 434
rect 70 433 71 434
rect 69 433 70 434
rect 66 433 67 434
rect 65 433 66 434
rect 64 433 65 434
rect 63 433 64 434
rect 62 433 63 434
rect 61 433 62 434
rect 60 433 61 434
rect 59 433 60 434
rect 58 433 59 434
rect 57 433 58 434
rect 56 433 57 434
rect 55 433 56 434
rect 54 433 55 434
rect 53 433 54 434
rect 52 433 53 434
rect 51 433 52 434
rect 50 433 51 434
rect 49 433 50 434
rect 48 433 49 434
rect 32 433 33 434
rect 31 433 32 434
rect 30 433 31 434
rect 29 433 30 434
rect 28 433 29 434
rect 27 433 28 434
rect 26 433 27 434
rect 25 433 26 434
rect 24 433 25 434
rect 23 433 24 434
rect 22 433 23 434
rect 21 433 22 434
rect 20 433 21 434
rect 19 433 20 434
rect 18 433 19 434
rect 17 433 18 434
rect 146 434 147 435
rect 145 434 146 435
rect 144 434 145 435
rect 143 434 144 435
rect 142 434 143 435
rect 141 434 142 435
rect 140 434 141 435
rect 139 434 140 435
rect 138 434 139 435
rect 137 434 138 435
rect 136 434 137 435
rect 135 434 136 435
rect 134 434 135 435
rect 133 434 134 435
rect 132 434 133 435
rect 131 434 132 435
rect 130 434 131 435
rect 129 434 130 435
rect 128 434 129 435
rect 127 434 128 435
rect 126 434 127 435
rect 125 434 126 435
rect 124 434 125 435
rect 123 434 124 435
rect 122 434 123 435
rect 121 434 122 435
rect 120 434 121 435
rect 119 434 120 435
rect 84 434 85 435
rect 83 434 84 435
rect 82 434 83 435
rect 81 434 82 435
rect 80 434 81 435
rect 79 434 80 435
rect 78 434 79 435
rect 77 434 78 435
rect 76 434 77 435
rect 75 434 76 435
rect 74 434 75 435
rect 73 434 74 435
rect 72 434 73 435
rect 71 434 72 435
rect 70 434 71 435
rect 69 434 70 435
rect 65 434 66 435
rect 64 434 65 435
rect 63 434 64 435
rect 62 434 63 435
rect 61 434 62 435
rect 60 434 61 435
rect 59 434 60 435
rect 58 434 59 435
rect 57 434 58 435
rect 56 434 57 435
rect 55 434 56 435
rect 54 434 55 435
rect 53 434 54 435
rect 52 434 53 435
rect 51 434 52 435
rect 50 434 51 435
rect 49 434 50 435
rect 48 434 49 435
rect 47 434 48 435
rect 33 434 34 435
rect 32 434 33 435
rect 31 434 32 435
rect 30 434 31 435
rect 29 434 30 435
rect 28 434 29 435
rect 27 434 28 435
rect 26 434 27 435
rect 25 434 26 435
rect 24 434 25 435
rect 23 434 24 435
rect 22 434 23 435
rect 21 434 22 435
rect 20 434 21 435
rect 19 434 20 435
rect 18 434 19 435
rect 17 434 18 435
rect 146 435 147 436
rect 145 435 146 436
rect 144 435 145 436
rect 143 435 144 436
rect 142 435 143 436
rect 141 435 142 436
rect 140 435 141 436
rect 139 435 140 436
rect 138 435 139 436
rect 137 435 138 436
rect 136 435 137 436
rect 135 435 136 436
rect 134 435 135 436
rect 133 435 134 436
rect 132 435 133 436
rect 131 435 132 436
rect 130 435 131 436
rect 129 435 130 436
rect 128 435 129 436
rect 127 435 128 436
rect 126 435 127 436
rect 125 435 126 436
rect 124 435 125 436
rect 123 435 124 436
rect 122 435 123 436
rect 121 435 122 436
rect 120 435 121 436
rect 119 435 120 436
rect 84 435 85 436
rect 83 435 84 436
rect 82 435 83 436
rect 81 435 82 436
rect 80 435 81 436
rect 79 435 80 436
rect 78 435 79 436
rect 77 435 78 436
rect 76 435 77 436
rect 75 435 76 436
rect 74 435 75 436
rect 73 435 74 436
rect 72 435 73 436
rect 71 435 72 436
rect 70 435 71 436
rect 69 435 70 436
rect 64 435 65 436
rect 63 435 64 436
rect 62 435 63 436
rect 61 435 62 436
rect 60 435 61 436
rect 59 435 60 436
rect 58 435 59 436
rect 57 435 58 436
rect 56 435 57 436
rect 55 435 56 436
rect 54 435 55 436
rect 53 435 54 436
rect 52 435 53 436
rect 51 435 52 436
rect 50 435 51 436
rect 49 435 50 436
rect 48 435 49 436
rect 47 435 48 436
rect 46 435 47 436
rect 33 435 34 436
rect 32 435 33 436
rect 31 435 32 436
rect 30 435 31 436
rect 29 435 30 436
rect 28 435 29 436
rect 27 435 28 436
rect 26 435 27 436
rect 25 435 26 436
rect 24 435 25 436
rect 23 435 24 436
rect 22 435 23 436
rect 21 435 22 436
rect 20 435 21 436
rect 19 435 20 436
rect 18 435 19 436
rect 17 435 18 436
rect 146 436 147 437
rect 145 436 146 437
rect 144 436 145 437
rect 143 436 144 437
rect 142 436 143 437
rect 141 436 142 437
rect 140 436 141 437
rect 139 436 140 437
rect 138 436 139 437
rect 137 436 138 437
rect 136 436 137 437
rect 135 436 136 437
rect 134 436 135 437
rect 133 436 134 437
rect 132 436 133 437
rect 131 436 132 437
rect 130 436 131 437
rect 129 436 130 437
rect 128 436 129 437
rect 127 436 128 437
rect 126 436 127 437
rect 125 436 126 437
rect 124 436 125 437
rect 123 436 124 437
rect 122 436 123 437
rect 121 436 122 437
rect 120 436 121 437
rect 119 436 120 437
rect 84 436 85 437
rect 83 436 84 437
rect 82 436 83 437
rect 81 436 82 437
rect 80 436 81 437
rect 79 436 80 437
rect 78 436 79 437
rect 77 436 78 437
rect 76 436 77 437
rect 75 436 76 437
rect 74 436 75 437
rect 73 436 74 437
rect 72 436 73 437
rect 71 436 72 437
rect 70 436 71 437
rect 69 436 70 437
rect 63 436 64 437
rect 62 436 63 437
rect 61 436 62 437
rect 60 436 61 437
rect 59 436 60 437
rect 58 436 59 437
rect 57 436 58 437
rect 56 436 57 437
rect 55 436 56 437
rect 54 436 55 437
rect 53 436 54 437
rect 52 436 53 437
rect 51 436 52 437
rect 50 436 51 437
rect 49 436 50 437
rect 48 436 49 437
rect 47 436 48 437
rect 46 436 47 437
rect 45 436 46 437
rect 44 436 45 437
rect 34 436 35 437
rect 33 436 34 437
rect 32 436 33 437
rect 31 436 32 437
rect 30 436 31 437
rect 29 436 30 437
rect 28 436 29 437
rect 27 436 28 437
rect 26 436 27 437
rect 25 436 26 437
rect 24 436 25 437
rect 23 436 24 437
rect 22 436 23 437
rect 21 436 22 437
rect 20 436 21 437
rect 19 436 20 437
rect 18 436 19 437
rect 17 436 18 437
rect 146 437 147 438
rect 145 437 146 438
rect 144 437 145 438
rect 143 437 144 438
rect 142 437 143 438
rect 141 437 142 438
rect 140 437 141 438
rect 139 437 140 438
rect 138 437 139 438
rect 137 437 138 438
rect 136 437 137 438
rect 135 437 136 438
rect 134 437 135 438
rect 133 437 134 438
rect 132 437 133 438
rect 131 437 132 438
rect 130 437 131 438
rect 129 437 130 438
rect 128 437 129 438
rect 127 437 128 438
rect 126 437 127 438
rect 125 437 126 438
rect 124 437 125 438
rect 123 437 124 438
rect 122 437 123 438
rect 121 437 122 438
rect 120 437 121 438
rect 119 437 120 438
rect 84 437 85 438
rect 83 437 84 438
rect 82 437 83 438
rect 81 437 82 438
rect 80 437 81 438
rect 79 437 80 438
rect 78 437 79 438
rect 77 437 78 438
rect 76 437 77 438
rect 75 437 76 438
rect 74 437 75 438
rect 73 437 74 438
rect 72 437 73 438
rect 71 437 72 438
rect 70 437 71 438
rect 69 437 70 438
rect 62 437 63 438
rect 61 437 62 438
rect 60 437 61 438
rect 59 437 60 438
rect 58 437 59 438
rect 57 437 58 438
rect 56 437 57 438
rect 55 437 56 438
rect 54 437 55 438
rect 53 437 54 438
rect 52 437 53 438
rect 51 437 52 438
rect 50 437 51 438
rect 49 437 50 438
rect 48 437 49 438
rect 47 437 48 438
rect 46 437 47 438
rect 45 437 46 438
rect 44 437 45 438
rect 43 437 44 438
rect 42 437 43 438
rect 36 437 37 438
rect 35 437 36 438
rect 34 437 35 438
rect 33 437 34 438
rect 32 437 33 438
rect 31 437 32 438
rect 30 437 31 438
rect 29 437 30 438
rect 28 437 29 438
rect 27 437 28 438
rect 26 437 27 438
rect 25 437 26 438
rect 24 437 25 438
rect 23 437 24 438
rect 22 437 23 438
rect 21 437 22 438
rect 20 437 21 438
rect 19 437 20 438
rect 18 437 19 438
rect 17 437 18 438
rect 138 438 139 439
rect 137 438 138 439
rect 136 438 137 439
rect 84 438 85 439
rect 83 438 84 439
rect 82 438 83 439
rect 81 438 82 439
rect 80 438 81 439
rect 79 438 80 439
rect 78 438 79 439
rect 77 438 78 439
rect 76 438 77 439
rect 75 438 76 439
rect 74 438 75 439
rect 73 438 74 439
rect 72 438 73 439
rect 71 438 72 439
rect 70 438 71 439
rect 69 438 70 439
rect 62 438 63 439
rect 61 438 62 439
rect 60 438 61 439
rect 59 438 60 439
rect 58 438 59 439
rect 57 438 58 439
rect 56 438 57 439
rect 55 438 56 439
rect 54 438 55 439
rect 53 438 54 439
rect 52 438 53 439
rect 51 438 52 439
rect 50 438 51 439
rect 49 438 50 439
rect 48 438 49 439
rect 47 438 48 439
rect 46 438 47 439
rect 45 438 46 439
rect 44 438 45 439
rect 43 438 44 439
rect 42 438 43 439
rect 41 438 42 439
rect 40 438 41 439
rect 39 438 40 439
rect 38 438 39 439
rect 37 438 38 439
rect 36 438 37 439
rect 35 438 36 439
rect 34 438 35 439
rect 33 438 34 439
rect 32 438 33 439
rect 31 438 32 439
rect 30 438 31 439
rect 29 438 30 439
rect 28 438 29 439
rect 27 438 28 439
rect 26 438 27 439
rect 25 438 26 439
rect 24 438 25 439
rect 23 438 24 439
rect 22 438 23 439
rect 21 438 22 439
rect 20 438 21 439
rect 19 438 20 439
rect 18 438 19 439
rect 17 438 18 439
rect 139 439 140 440
rect 138 439 139 440
rect 137 439 138 440
rect 136 439 137 440
rect 135 439 136 440
rect 134 439 135 440
rect 84 439 85 440
rect 83 439 84 440
rect 82 439 83 440
rect 81 439 82 440
rect 80 439 81 440
rect 79 439 80 440
rect 78 439 79 440
rect 77 439 78 440
rect 76 439 77 440
rect 75 439 76 440
rect 74 439 75 440
rect 73 439 74 440
rect 72 439 73 440
rect 71 439 72 440
rect 70 439 71 440
rect 69 439 70 440
rect 61 439 62 440
rect 60 439 61 440
rect 59 439 60 440
rect 58 439 59 440
rect 57 439 58 440
rect 56 439 57 440
rect 55 439 56 440
rect 54 439 55 440
rect 53 439 54 440
rect 52 439 53 440
rect 51 439 52 440
rect 50 439 51 440
rect 49 439 50 440
rect 48 439 49 440
rect 47 439 48 440
rect 46 439 47 440
rect 45 439 46 440
rect 44 439 45 440
rect 43 439 44 440
rect 42 439 43 440
rect 41 439 42 440
rect 40 439 41 440
rect 39 439 40 440
rect 38 439 39 440
rect 37 439 38 440
rect 36 439 37 440
rect 35 439 36 440
rect 34 439 35 440
rect 33 439 34 440
rect 32 439 33 440
rect 31 439 32 440
rect 30 439 31 440
rect 29 439 30 440
rect 28 439 29 440
rect 27 439 28 440
rect 26 439 27 440
rect 25 439 26 440
rect 24 439 25 440
rect 23 439 24 440
rect 22 439 23 440
rect 21 439 22 440
rect 20 439 21 440
rect 19 439 20 440
rect 18 439 19 440
rect 17 439 18 440
rect 141 440 142 441
rect 140 440 141 441
rect 139 440 140 441
rect 138 440 139 441
rect 137 440 138 441
rect 136 440 137 441
rect 135 440 136 441
rect 134 440 135 441
rect 133 440 134 441
rect 84 440 85 441
rect 83 440 84 441
rect 82 440 83 441
rect 81 440 82 441
rect 80 440 81 441
rect 79 440 80 441
rect 78 440 79 441
rect 77 440 78 441
rect 76 440 77 441
rect 75 440 76 441
rect 74 440 75 441
rect 73 440 74 441
rect 72 440 73 441
rect 71 440 72 441
rect 70 440 71 441
rect 69 440 70 441
rect 60 440 61 441
rect 59 440 60 441
rect 58 440 59 441
rect 57 440 58 441
rect 56 440 57 441
rect 55 440 56 441
rect 54 440 55 441
rect 53 440 54 441
rect 52 440 53 441
rect 51 440 52 441
rect 50 440 51 441
rect 49 440 50 441
rect 48 440 49 441
rect 47 440 48 441
rect 46 440 47 441
rect 45 440 46 441
rect 44 440 45 441
rect 43 440 44 441
rect 42 440 43 441
rect 41 440 42 441
rect 40 440 41 441
rect 39 440 40 441
rect 38 440 39 441
rect 37 440 38 441
rect 36 440 37 441
rect 35 440 36 441
rect 34 440 35 441
rect 33 440 34 441
rect 32 440 33 441
rect 31 440 32 441
rect 30 440 31 441
rect 29 440 30 441
rect 28 440 29 441
rect 27 440 28 441
rect 26 440 27 441
rect 25 440 26 441
rect 24 440 25 441
rect 23 440 24 441
rect 22 440 23 441
rect 21 440 22 441
rect 20 440 21 441
rect 19 440 20 441
rect 18 440 19 441
rect 17 440 18 441
rect 142 441 143 442
rect 141 441 142 442
rect 140 441 141 442
rect 139 441 140 442
rect 138 441 139 442
rect 137 441 138 442
rect 136 441 137 442
rect 135 441 136 442
rect 134 441 135 442
rect 133 441 134 442
rect 132 441 133 442
rect 131 441 132 442
rect 84 441 85 442
rect 83 441 84 442
rect 82 441 83 442
rect 81 441 82 442
rect 80 441 81 442
rect 79 441 80 442
rect 78 441 79 442
rect 77 441 78 442
rect 76 441 77 442
rect 75 441 76 442
rect 74 441 75 442
rect 73 441 74 442
rect 72 441 73 442
rect 71 441 72 442
rect 70 441 71 442
rect 69 441 70 442
rect 59 441 60 442
rect 58 441 59 442
rect 57 441 58 442
rect 56 441 57 442
rect 55 441 56 442
rect 54 441 55 442
rect 53 441 54 442
rect 52 441 53 442
rect 51 441 52 442
rect 50 441 51 442
rect 49 441 50 442
rect 48 441 49 442
rect 47 441 48 442
rect 46 441 47 442
rect 45 441 46 442
rect 44 441 45 442
rect 43 441 44 442
rect 42 441 43 442
rect 41 441 42 442
rect 40 441 41 442
rect 39 441 40 442
rect 38 441 39 442
rect 37 441 38 442
rect 36 441 37 442
rect 35 441 36 442
rect 34 441 35 442
rect 33 441 34 442
rect 32 441 33 442
rect 31 441 32 442
rect 30 441 31 442
rect 29 441 30 442
rect 28 441 29 442
rect 27 441 28 442
rect 26 441 27 442
rect 25 441 26 442
rect 24 441 25 442
rect 23 441 24 442
rect 22 441 23 442
rect 21 441 22 442
rect 20 441 21 442
rect 19 441 20 442
rect 18 441 19 442
rect 144 442 145 443
rect 143 442 144 443
rect 142 442 143 443
rect 141 442 142 443
rect 140 442 141 443
rect 139 442 140 443
rect 138 442 139 443
rect 137 442 138 443
rect 136 442 137 443
rect 135 442 136 443
rect 134 442 135 443
rect 133 442 134 443
rect 132 442 133 443
rect 131 442 132 443
rect 130 442 131 443
rect 84 442 85 443
rect 83 442 84 443
rect 82 442 83 443
rect 81 442 82 443
rect 80 442 81 443
rect 79 442 80 443
rect 78 442 79 443
rect 77 442 78 443
rect 76 442 77 443
rect 75 442 76 443
rect 74 442 75 443
rect 73 442 74 443
rect 72 442 73 443
rect 71 442 72 443
rect 70 442 71 443
rect 69 442 70 443
rect 59 442 60 443
rect 58 442 59 443
rect 57 442 58 443
rect 56 442 57 443
rect 55 442 56 443
rect 54 442 55 443
rect 53 442 54 443
rect 52 442 53 443
rect 51 442 52 443
rect 50 442 51 443
rect 49 442 50 443
rect 48 442 49 443
rect 47 442 48 443
rect 46 442 47 443
rect 45 442 46 443
rect 44 442 45 443
rect 43 442 44 443
rect 42 442 43 443
rect 41 442 42 443
rect 40 442 41 443
rect 39 442 40 443
rect 38 442 39 443
rect 37 442 38 443
rect 36 442 37 443
rect 35 442 36 443
rect 34 442 35 443
rect 33 442 34 443
rect 32 442 33 443
rect 31 442 32 443
rect 30 442 31 443
rect 29 442 30 443
rect 28 442 29 443
rect 27 442 28 443
rect 26 442 27 443
rect 25 442 26 443
rect 24 442 25 443
rect 23 442 24 443
rect 22 442 23 443
rect 21 442 22 443
rect 20 442 21 443
rect 19 442 20 443
rect 18 442 19 443
rect 145 443 146 444
rect 144 443 145 444
rect 143 443 144 444
rect 142 443 143 444
rect 141 443 142 444
rect 140 443 141 444
rect 139 443 140 444
rect 138 443 139 444
rect 137 443 138 444
rect 136 443 137 444
rect 135 443 136 444
rect 134 443 135 444
rect 133 443 134 444
rect 132 443 133 444
rect 131 443 132 444
rect 130 443 131 444
rect 129 443 130 444
rect 128 443 129 444
rect 84 443 85 444
rect 83 443 84 444
rect 82 443 83 444
rect 81 443 82 444
rect 80 443 81 444
rect 79 443 80 444
rect 78 443 79 444
rect 77 443 78 444
rect 76 443 77 444
rect 75 443 76 444
rect 74 443 75 444
rect 73 443 74 444
rect 72 443 73 444
rect 71 443 72 444
rect 70 443 71 444
rect 69 443 70 444
rect 58 443 59 444
rect 57 443 58 444
rect 56 443 57 444
rect 55 443 56 444
rect 54 443 55 444
rect 53 443 54 444
rect 52 443 53 444
rect 51 443 52 444
rect 50 443 51 444
rect 49 443 50 444
rect 48 443 49 444
rect 47 443 48 444
rect 46 443 47 444
rect 45 443 46 444
rect 44 443 45 444
rect 43 443 44 444
rect 42 443 43 444
rect 41 443 42 444
rect 40 443 41 444
rect 39 443 40 444
rect 38 443 39 444
rect 37 443 38 444
rect 36 443 37 444
rect 35 443 36 444
rect 34 443 35 444
rect 33 443 34 444
rect 32 443 33 444
rect 31 443 32 444
rect 30 443 31 444
rect 29 443 30 444
rect 28 443 29 444
rect 27 443 28 444
rect 26 443 27 444
rect 25 443 26 444
rect 24 443 25 444
rect 23 443 24 444
rect 22 443 23 444
rect 21 443 22 444
rect 20 443 21 444
rect 19 443 20 444
rect 18 443 19 444
rect 146 444 147 445
rect 145 444 146 445
rect 144 444 145 445
rect 143 444 144 445
rect 142 444 143 445
rect 141 444 142 445
rect 140 444 141 445
rect 139 444 140 445
rect 138 444 139 445
rect 135 444 136 445
rect 134 444 135 445
rect 133 444 134 445
rect 132 444 133 445
rect 131 444 132 445
rect 130 444 131 445
rect 129 444 130 445
rect 128 444 129 445
rect 84 444 85 445
rect 83 444 84 445
rect 82 444 83 445
rect 81 444 82 445
rect 80 444 81 445
rect 79 444 80 445
rect 78 444 79 445
rect 77 444 78 445
rect 76 444 77 445
rect 75 444 76 445
rect 74 444 75 445
rect 73 444 74 445
rect 72 444 73 445
rect 71 444 72 445
rect 70 444 71 445
rect 69 444 70 445
rect 58 444 59 445
rect 57 444 58 445
rect 56 444 57 445
rect 55 444 56 445
rect 54 444 55 445
rect 53 444 54 445
rect 52 444 53 445
rect 51 444 52 445
rect 50 444 51 445
rect 49 444 50 445
rect 48 444 49 445
rect 47 444 48 445
rect 46 444 47 445
rect 45 444 46 445
rect 44 444 45 445
rect 43 444 44 445
rect 42 444 43 445
rect 41 444 42 445
rect 40 444 41 445
rect 39 444 40 445
rect 38 444 39 445
rect 37 444 38 445
rect 36 444 37 445
rect 35 444 36 445
rect 34 444 35 445
rect 33 444 34 445
rect 32 444 33 445
rect 31 444 32 445
rect 30 444 31 445
rect 29 444 30 445
rect 28 444 29 445
rect 27 444 28 445
rect 26 444 27 445
rect 25 444 26 445
rect 24 444 25 445
rect 23 444 24 445
rect 22 444 23 445
rect 21 444 22 445
rect 20 444 21 445
rect 19 444 20 445
rect 18 444 19 445
rect 146 445 147 446
rect 145 445 146 446
rect 144 445 145 446
rect 143 445 144 446
rect 142 445 143 446
rect 141 445 142 446
rect 140 445 141 446
rect 133 445 134 446
rect 132 445 133 446
rect 131 445 132 446
rect 130 445 131 446
rect 129 445 130 446
rect 128 445 129 446
rect 84 445 85 446
rect 83 445 84 446
rect 82 445 83 446
rect 81 445 82 446
rect 80 445 81 446
rect 79 445 80 446
rect 78 445 79 446
rect 77 445 78 446
rect 76 445 77 446
rect 75 445 76 446
rect 74 445 75 446
rect 73 445 74 446
rect 72 445 73 446
rect 71 445 72 446
rect 70 445 71 446
rect 69 445 70 446
rect 57 445 58 446
rect 56 445 57 446
rect 55 445 56 446
rect 54 445 55 446
rect 53 445 54 446
rect 52 445 53 446
rect 51 445 52 446
rect 50 445 51 446
rect 49 445 50 446
rect 48 445 49 446
rect 47 445 48 446
rect 46 445 47 446
rect 45 445 46 446
rect 44 445 45 446
rect 43 445 44 446
rect 42 445 43 446
rect 41 445 42 446
rect 40 445 41 446
rect 39 445 40 446
rect 38 445 39 446
rect 37 445 38 446
rect 36 445 37 446
rect 35 445 36 446
rect 34 445 35 446
rect 33 445 34 446
rect 32 445 33 446
rect 31 445 32 446
rect 30 445 31 446
rect 29 445 30 446
rect 28 445 29 446
rect 27 445 28 446
rect 26 445 27 446
rect 25 445 26 446
rect 24 445 25 446
rect 23 445 24 446
rect 22 445 23 446
rect 21 445 22 446
rect 20 445 21 446
rect 19 445 20 446
rect 146 446 147 447
rect 145 446 146 447
rect 144 446 145 447
rect 143 446 144 447
rect 142 446 143 447
rect 141 446 142 447
rect 132 446 133 447
rect 131 446 132 447
rect 130 446 131 447
rect 129 446 130 447
rect 128 446 129 447
rect 84 446 85 447
rect 83 446 84 447
rect 82 446 83 447
rect 81 446 82 447
rect 80 446 81 447
rect 79 446 80 447
rect 78 446 79 447
rect 77 446 78 447
rect 76 446 77 447
rect 75 446 76 447
rect 74 446 75 447
rect 73 446 74 447
rect 72 446 73 447
rect 71 446 72 447
rect 70 446 71 447
rect 69 446 70 447
rect 56 446 57 447
rect 55 446 56 447
rect 54 446 55 447
rect 53 446 54 447
rect 52 446 53 447
rect 51 446 52 447
rect 50 446 51 447
rect 49 446 50 447
rect 48 446 49 447
rect 47 446 48 447
rect 46 446 47 447
rect 45 446 46 447
rect 44 446 45 447
rect 43 446 44 447
rect 42 446 43 447
rect 41 446 42 447
rect 40 446 41 447
rect 39 446 40 447
rect 38 446 39 447
rect 37 446 38 447
rect 36 446 37 447
rect 35 446 36 447
rect 34 446 35 447
rect 33 446 34 447
rect 32 446 33 447
rect 31 446 32 447
rect 30 446 31 447
rect 29 446 30 447
rect 28 446 29 447
rect 27 446 28 447
rect 26 446 27 447
rect 25 446 26 447
rect 24 446 25 447
rect 23 446 24 447
rect 22 446 23 447
rect 21 446 22 447
rect 20 446 21 447
rect 19 446 20 447
rect 146 447 147 448
rect 145 447 146 448
rect 144 447 145 448
rect 143 447 144 448
rect 142 447 143 448
rect 131 447 132 448
rect 130 447 131 448
rect 129 447 130 448
rect 128 447 129 448
rect 84 447 85 448
rect 83 447 84 448
rect 82 447 83 448
rect 81 447 82 448
rect 80 447 81 448
rect 79 447 80 448
rect 78 447 79 448
rect 77 447 78 448
rect 76 447 77 448
rect 75 447 76 448
rect 74 447 75 448
rect 73 447 74 448
rect 72 447 73 448
rect 71 447 72 448
rect 70 447 71 448
rect 69 447 70 448
rect 55 447 56 448
rect 54 447 55 448
rect 53 447 54 448
rect 52 447 53 448
rect 51 447 52 448
rect 50 447 51 448
rect 49 447 50 448
rect 48 447 49 448
rect 47 447 48 448
rect 46 447 47 448
rect 45 447 46 448
rect 44 447 45 448
rect 43 447 44 448
rect 42 447 43 448
rect 41 447 42 448
rect 40 447 41 448
rect 39 447 40 448
rect 38 447 39 448
rect 37 447 38 448
rect 36 447 37 448
rect 35 447 36 448
rect 34 447 35 448
rect 33 447 34 448
rect 32 447 33 448
rect 31 447 32 448
rect 30 447 31 448
rect 29 447 30 448
rect 28 447 29 448
rect 27 447 28 448
rect 26 447 27 448
rect 25 447 26 448
rect 24 447 25 448
rect 23 447 24 448
rect 22 447 23 448
rect 21 447 22 448
rect 20 447 21 448
rect 146 448 147 449
rect 145 448 146 449
rect 144 448 145 449
rect 129 448 130 449
rect 128 448 129 449
rect 84 448 85 449
rect 83 448 84 449
rect 82 448 83 449
rect 81 448 82 449
rect 80 448 81 449
rect 79 448 80 449
rect 78 448 79 449
rect 77 448 78 449
rect 76 448 77 449
rect 75 448 76 449
rect 74 448 75 449
rect 73 448 74 449
rect 72 448 73 449
rect 71 448 72 449
rect 70 448 71 449
rect 69 448 70 449
rect 55 448 56 449
rect 54 448 55 449
rect 53 448 54 449
rect 52 448 53 449
rect 51 448 52 449
rect 50 448 51 449
rect 49 448 50 449
rect 48 448 49 449
rect 47 448 48 449
rect 46 448 47 449
rect 45 448 46 449
rect 44 448 45 449
rect 43 448 44 449
rect 42 448 43 449
rect 41 448 42 449
rect 40 448 41 449
rect 39 448 40 449
rect 38 448 39 449
rect 37 448 38 449
rect 36 448 37 449
rect 35 448 36 449
rect 34 448 35 449
rect 33 448 34 449
rect 32 448 33 449
rect 31 448 32 449
rect 30 448 31 449
rect 29 448 30 449
rect 28 448 29 449
rect 27 448 28 449
rect 26 448 27 449
rect 25 448 26 449
rect 24 448 25 449
rect 23 448 24 449
rect 22 448 23 449
rect 21 448 22 449
rect 20 448 21 449
rect 146 449 147 450
rect 145 449 146 450
rect 128 449 129 450
rect 84 449 85 450
rect 83 449 84 450
rect 82 449 83 450
rect 81 449 82 450
rect 80 449 81 450
rect 79 449 80 450
rect 78 449 79 450
rect 77 449 78 450
rect 76 449 77 450
rect 75 449 76 450
rect 74 449 75 450
rect 73 449 74 450
rect 72 449 73 450
rect 71 449 72 450
rect 70 449 71 450
rect 69 449 70 450
rect 54 449 55 450
rect 53 449 54 450
rect 52 449 53 450
rect 51 449 52 450
rect 50 449 51 450
rect 49 449 50 450
rect 48 449 49 450
rect 47 449 48 450
rect 46 449 47 450
rect 45 449 46 450
rect 44 449 45 450
rect 43 449 44 450
rect 42 449 43 450
rect 41 449 42 450
rect 40 449 41 450
rect 39 449 40 450
rect 38 449 39 450
rect 37 449 38 450
rect 36 449 37 450
rect 35 449 36 450
rect 34 449 35 450
rect 33 449 34 450
rect 32 449 33 450
rect 31 449 32 450
rect 30 449 31 450
rect 29 449 30 450
rect 28 449 29 450
rect 27 449 28 450
rect 26 449 27 450
rect 25 449 26 450
rect 24 449 25 450
rect 23 449 24 450
rect 22 449 23 450
rect 21 449 22 450
rect 84 450 85 451
rect 83 450 84 451
rect 82 450 83 451
rect 81 450 82 451
rect 80 450 81 451
rect 79 450 80 451
rect 78 450 79 451
rect 77 450 78 451
rect 76 450 77 451
rect 75 450 76 451
rect 74 450 75 451
rect 73 450 74 451
rect 72 450 73 451
rect 71 450 72 451
rect 70 450 71 451
rect 69 450 70 451
rect 53 450 54 451
rect 52 450 53 451
rect 51 450 52 451
rect 50 450 51 451
rect 49 450 50 451
rect 48 450 49 451
rect 47 450 48 451
rect 46 450 47 451
rect 45 450 46 451
rect 44 450 45 451
rect 43 450 44 451
rect 42 450 43 451
rect 41 450 42 451
rect 40 450 41 451
rect 39 450 40 451
rect 38 450 39 451
rect 37 450 38 451
rect 36 450 37 451
rect 35 450 36 451
rect 34 450 35 451
rect 33 450 34 451
rect 32 450 33 451
rect 31 450 32 451
rect 30 450 31 451
rect 29 450 30 451
rect 28 450 29 451
rect 27 450 28 451
rect 26 450 27 451
rect 25 450 26 451
rect 24 450 25 451
rect 23 450 24 451
rect 22 450 23 451
rect 21 450 22 451
rect 84 451 85 452
rect 83 451 84 452
rect 82 451 83 452
rect 81 451 82 452
rect 80 451 81 452
rect 79 451 80 452
rect 78 451 79 452
rect 77 451 78 452
rect 76 451 77 452
rect 75 451 76 452
rect 74 451 75 452
rect 73 451 74 452
rect 72 451 73 452
rect 71 451 72 452
rect 70 451 71 452
rect 69 451 70 452
rect 52 451 53 452
rect 51 451 52 452
rect 50 451 51 452
rect 49 451 50 452
rect 48 451 49 452
rect 47 451 48 452
rect 46 451 47 452
rect 45 451 46 452
rect 44 451 45 452
rect 43 451 44 452
rect 42 451 43 452
rect 41 451 42 452
rect 40 451 41 452
rect 39 451 40 452
rect 38 451 39 452
rect 37 451 38 452
rect 36 451 37 452
rect 35 451 36 452
rect 34 451 35 452
rect 33 451 34 452
rect 32 451 33 452
rect 31 451 32 452
rect 30 451 31 452
rect 29 451 30 452
rect 28 451 29 452
rect 27 451 28 452
rect 26 451 27 452
rect 25 451 26 452
rect 24 451 25 452
rect 23 451 24 452
rect 22 451 23 452
rect 84 452 85 453
rect 83 452 84 453
rect 82 452 83 453
rect 81 452 82 453
rect 80 452 81 453
rect 79 452 80 453
rect 78 452 79 453
rect 77 452 78 453
rect 76 452 77 453
rect 75 452 76 453
rect 74 452 75 453
rect 73 452 74 453
rect 72 452 73 453
rect 71 452 72 453
rect 70 452 71 453
rect 69 452 70 453
rect 51 452 52 453
rect 50 452 51 453
rect 49 452 50 453
rect 48 452 49 453
rect 47 452 48 453
rect 46 452 47 453
rect 45 452 46 453
rect 44 452 45 453
rect 43 452 44 453
rect 42 452 43 453
rect 41 452 42 453
rect 40 452 41 453
rect 39 452 40 453
rect 38 452 39 453
rect 37 452 38 453
rect 36 452 37 453
rect 35 452 36 453
rect 34 452 35 453
rect 33 452 34 453
rect 32 452 33 453
rect 31 452 32 453
rect 30 452 31 453
rect 29 452 30 453
rect 28 452 29 453
rect 27 452 28 453
rect 26 452 27 453
rect 25 452 26 453
rect 24 452 25 453
rect 23 452 24 453
rect 84 453 85 454
rect 83 453 84 454
rect 82 453 83 454
rect 81 453 82 454
rect 80 453 81 454
rect 79 453 80 454
rect 78 453 79 454
rect 77 453 78 454
rect 76 453 77 454
rect 75 453 76 454
rect 74 453 75 454
rect 73 453 74 454
rect 72 453 73 454
rect 71 453 72 454
rect 70 453 71 454
rect 69 453 70 454
rect 50 453 51 454
rect 49 453 50 454
rect 48 453 49 454
rect 47 453 48 454
rect 46 453 47 454
rect 45 453 46 454
rect 44 453 45 454
rect 43 453 44 454
rect 42 453 43 454
rect 41 453 42 454
rect 40 453 41 454
rect 39 453 40 454
rect 38 453 39 454
rect 37 453 38 454
rect 36 453 37 454
rect 35 453 36 454
rect 34 453 35 454
rect 33 453 34 454
rect 32 453 33 454
rect 31 453 32 454
rect 30 453 31 454
rect 29 453 30 454
rect 28 453 29 454
rect 27 453 28 454
rect 26 453 27 454
rect 25 453 26 454
rect 24 453 25 454
rect 84 454 85 455
rect 83 454 84 455
rect 82 454 83 455
rect 81 454 82 455
rect 80 454 81 455
rect 79 454 80 455
rect 78 454 79 455
rect 77 454 78 455
rect 76 454 77 455
rect 75 454 76 455
rect 74 454 75 455
rect 73 454 74 455
rect 72 454 73 455
rect 71 454 72 455
rect 70 454 71 455
rect 69 454 70 455
rect 48 454 49 455
rect 47 454 48 455
rect 46 454 47 455
rect 45 454 46 455
rect 44 454 45 455
rect 43 454 44 455
rect 42 454 43 455
rect 41 454 42 455
rect 40 454 41 455
rect 39 454 40 455
rect 38 454 39 455
rect 37 454 38 455
rect 36 454 37 455
rect 35 454 36 455
rect 34 454 35 455
rect 33 454 34 455
rect 32 454 33 455
rect 31 454 32 455
rect 30 454 31 455
rect 29 454 30 455
rect 28 454 29 455
rect 27 454 28 455
rect 26 454 27 455
rect 25 454 26 455
rect 84 455 85 456
rect 83 455 84 456
rect 82 455 83 456
rect 81 455 82 456
rect 80 455 81 456
rect 79 455 80 456
rect 78 455 79 456
rect 77 455 78 456
rect 76 455 77 456
rect 75 455 76 456
rect 74 455 75 456
rect 73 455 74 456
rect 72 455 73 456
rect 71 455 72 456
rect 70 455 71 456
rect 69 455 70 456
rect 46 455 47 456
rect 45 455 46 456
rect 44 455 45 456
rect 43 455 44 456
rect 42 455 43 456
rect 41 455 42 456
rect 40 455 41 456
rect 39 455 40 456
rect 38 455 39 456
rect 37 455 38 456
rect 36 455 37 456
rect 35 455 36 456
rect 34 455 35 456
rect 33 455 34 456
rect 32 455 33 456
rect 31 455 32 456
rect 30 455 31 456
rect 29 455 30 456
rect 28 455 29 456
rect 27 455 28 456
rect 84 456 85 457
rect 83 456 84 457
rect 82 456 83 457
rect 81 456 82 457
rect 80 456 81 457
rect 79 456 80 457
rect 78 456 79 457
rect 77 456 78 457
rect 76 456 77 457
rect 75 456 76 457
rect 74 456 75 457
rect 73 456 74 457
rect 72 456 73 457
rect 71 456 72 457
rect 70 456 71 457
rect 69 456 70 457
rect 44 456 45 457
rect 43 456 44 457
rect 42 456 43 457
rect 41 456 42 457
rect 40 456 41 457
rect 39 456 40 457
rect 38 456 39 457
rect 37 456 38 457
rect 36 456 37 457
rect 35 456 36 457
rect 34 456 35 457
rect 33 456 34 457
rect 32 456 33 457
rect 31 456 32 457
rect 30 456 31 457
rect 29 456 30 457
rect 84 457 85 458
rect 83 457 84 458
rect 82 457 83 458
rect 81 457 82 458
rect 80 457 81 458
rect 79 457 80 458
rect 78 457 79 458
rect 77 457 78 458
rect 76 457 77 458
rect 75 457 76 458
rect 74 457 75 458
rect 73 457 74 458
rect 72 457 73 458
rect 71 457 72 458
rect 70 457 71 458
rect 69 457 70 458
rect 39 457 40 458
rect 38 457 39 458
rect 37 457 38 458
rect 36 457 37 458
rect 35 457 36 458
rect 34 457 35 458
<< end >>
