magic
tech scmos
timestamp 1701862152
<< checkpaint >>
rect 13 71 87 79
rect -7 39 87 71
rect -7 30 67 39
<< nwell >>
rect -6 77 86 136
<< ntransistor >>
rect 19 7 21 17
rect 29 7 31 17
rect 39 7 41 17
<< ptransistor >>
rect 9 93 11 123
rect 19 93 21 123
rect 29 93 31 123
rect 39 93 41 123
rect 59 89 61 119
rect 69 89 71 119
<< ndiffusion >>
rect 18 7 19 17
rect 21 7 22 17
rect 28 7 29 17
rect 31 7 32 17
rect 38 7 39 17
rect 41 7 42 17
<< pdiffusion >>
rect 8 93 9 123
rect 11 93 12 123
rect 18 93 19 123
rect 21 93 22 123
rect 28 93 29 123
rect 31 117 39 123
rect 31 93 32 117
rect 38 93 39 117
rect 41 94 42 123
rect 41 93 44 94
rect 58 89 59 119
rect 61 117 69 119
rect 61 91 62 117
rect 68 91 69 117
rect 61 89 69 91
rect 71 89 72 119
<< ndcontact >>
rect 11 7 18 17
rect 22 7 28 17
rect 32 7 38 17
rect 42 7 48 17
<< pdcontact >>
rect 2 93 8 123
rect 12 93 18 123
rect 22 93 28 123
rect 32 93 38 117
rect 42 94 48 123
rect 52 89 58 119
rect 62 91 68 117
rect 72 89 78 119
<< psubstratepcontact >>
rect -3 -3 83 3
<< nsubstratencontact >>
rect -3 127 83 133
<< polysilicon >>
rect 9 123 11 125
rect 19 123 21 125
rect 29 123 31 125
rect 39 123 41 125
rect 59 119 61 121
rect 69 119 71 121
rect 9 92 11 93
rect 19 92 21 93
rect 9 90 21 92
rect 19 64 21 90
rect 18 58 21 64
rect 19 17 21 58
rect 29 92 31 93
rect 39 92 41 93
rect 29 90 41 92
rect 29 17 31 90
rect 59 85 61 89
rect 69 85 71 89
rect 48 83 71 85
rect 48 28 51 83
rect 39 25 51 28
rect 39 17 41 25
rect 19 5 21 7
rect 29 5 31 7
rect 39 5 41 7
<< polycontact >>
rect 12 58 18 64
rect 42 58 48 64
rect 31 45 37 51
<< metal1 >>
rect -3 133 83 134
rect -3 126 83 127
rect 12 123 18 126
rect 28 120 42 123
rect 2 90 8 93
rect 22 90 28 93
rect 2 87 28 90
rect 52 120 78 123
rect 52 119 58 120
rect 32 91 38 93
rect 32 89 52 91
rect 72 119 78 120
rect 32 88 58 89
rect 62 58 66 91
rect 62 23 66 51
rect 24 20 66 23
rect 24 17 27 20
rect 48 7 51 20
rect 11 4 18 7
rect 32 4 38 7
rect -3 3 83 4
rect -3 -4 83 -3
<< m2contact >>
rect 11 51 18 58
rect 31 51 38 58
rect 41 51 48 58
rect 60 51 67 58
<< metal2 >>
rect 33 58 37 67
rect 63 58 67 67
rect 13 43 17 51
rect 43 43 47 51
<< m1p >>
rect -3 126 83 134
rect -3 -4 83 4
<< m2p >>
rect 33 59 37 67
rect 63 59 67 67
rect 13 43 17 50
rect 43 43 47 50
<< labels >>
rlabel metal2 15 44 15 44 1 A
port 1 n signal input
rlabel metal2 35 65 35 65 1 B
port 2 n signal input
rlabel metal2 45 44 45 44 7 C
port 3 n signal input
rlabel metal2 65 65 65 65 1 Y
port 4 n signal output
rlabel metal1 -3 126 83 134 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -3 -4 83 4 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 80 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
