magic
tech scmos
magscale 1 3
timestamp 1554524574
<< checkpaint >>
rect -60 -60 152 152
<< genericcontact >>
rect 7 79 13 85
rect 19 79 25 85
rect 31 79 37 85
rect 43 79 49 85
rect 55 79 61 85
rect 67 79 73 85
rect 79 79 85 85
rect 7 67 13 73
rect 19 67 25 73
rect 31 67 37 73
rect 43 67 49 73
rect 55 67 61 73
rect 67 67 73 73
rect 79 67 85 73
rect 7 55 13 61
rect 19 55 25 61
rect 31 55 37 61
rect 43 55 49 61
rect 55 55 61 61
rect 67 55 73 61
rect 79 55 85 61
rect 7 43 13 49
rect 19 43 25 49
rect 31 43 37 49
rect 43 43 49 49
rect 55 43 61 49
rect 67 43 73 49
rect 79 43 85 49
rect 7 31 13 37
rect 19 31 25 37
rect 31 31 37 37
rect 43 31 49 37
rect 55 31 61 37
rect 67 31 73 37
rect 79 31 85 37
rect 7 19 13 25
rect 19 19 25 25
rect 31 19 37 25
rect 43 19 49 25
rect 55 19 61 25
rect 67 19 73 25
rect 79 19 85 25
rect 7 7 13 13
rect 19 7 25 13
rect 31 7 37 13
rect 43 7 49 13
rect 55 7 61 13
rect 67 7 73 13
rect 79 7 85 13
<< metal1 >>
rect 0 0 92 92
<< pseudo_rpoly2 >>
rect 1 1 91 91
<< end >>
