/* Verilog module written by vlog2Verilog (qflow) */

module fxp_sqrt_top(
    input ap_clk,
    output ap_done,
    output ap_idle,
    output ap_ready,
    output [27:0] ap_return,
    input ap_rst,
    input ap_start,
    input [23:0] in_val
);

wire vdd = 1'b1;
wire gnd = 1'b0;

wire _1677_ ;
wire _1257_ ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _1486_ ;
wire _1066_ ;
wire _397_ ;
wire ap_done ;
wire _1295_ ;
wire _941__bF$buf0 ;
wire _941__bF$buf1 ;
wire _941__bF$buf2 ;
wire _941__bF$buf3 ;
wire _941__bF$buf4 ;
wire _941__bF$buf5 ;
wire _941__bF$buf6 ;
wire _941__bF$buf7 ;
wire _941__bF$buf8 ;
wire _703_ ;
wire _1389_ ;
wire _19_ ;
wire _1601_ ;
wire _932_ ;
wire _512_ ;
wire _1198_ ;
wire _1410_ ;
wire _741_ ;
wire _321_ ;
wire _57_ ;
wire _970_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire _1504_ ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _1733_ ;
wire _1313_ ;
wire _644_ ;
wire _224_ ;
wire _1542_ ;
wire _1122_ ;
wire _873_ ;
wire _453_ ;
wire _929_ ;
wire _509_ ;
wire _1771_ ;
wire _1351_ ;
wire _682_ ;
wire _262_ ;
wire _1407_ ;
wire _738_ ;
wire _318_ ;
wire _1580_ ;
wire _1160_ ;
wire _491_ ;
wire _1636_ ;
wire _1216_ ;
wire _967_ ;
wire _547_ ;
wire _127_ ;
wire _1445_ ;
wire _1025_ ;
wire _776_ ;
wire _356_ ;
wire _1674_ ;
wire _1254_ ;
wire _585_ ;
wire _165_ ;
wire _1483_ ;
wire _1063_ ;
wire _394_ ;
wire _1539_ ;
wire _1119_ ;
wire _1292_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6  ;
wire _1768_ ;
wire _1348_ ;
wire _679_ ;
wire _259_ ;
wire _1577_ ;
wire _1157_ ;
wire _488_ ;
wire _700_ ;
wire _1386_ ;
wire _297_ ;
wire _16_ ;
wire _1195_ ;
wire _54_ ;
wire _603_ ;
wire _1289_ ;
wire _1501_ ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _1098_ ;
wire _1730_ ;
wire _1310_ ;
wire _641_ ;
wire _221_ ;
wire _870_ ;
wire _450_ ;
wire _926_ ;
wire _506_ ;
wire _1404_ ;
wire _735_ ;
wire _315_ ;
wire _1633_ ;
wire _1213_ ;
wire _964_ ;
wire _544_ ;
wire _124_ ;
wire _1442_ ;
wire _1022_ ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _1671_ ;
wire _1251_ ;
wire _582_ ;
wire _162_ ;
wire _1727_ ;
wire _1307_ ;
wire _638_ ;
wire _218_ ;
wire _1480_ ;
wire _1060_ ;
wire _391_ ;
wire _1536_ ;
wire _1116_ ;
wire _867_ ;
wire _447_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3  ;
wire _1765_ ;
wire _1345_ ;
wire _676_ ;
wire _256_ ;
wire _1574_ ;
wire _1154_ ;
wire _485_ ;
wire _1383_ ;
wire _294_ ;
wire _13_ ;
wire _1439_ ;
wire _1019_ ;
wire _1192_ ;
wire [27:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3  ;
wire _1668_ ;
wire _1248_ ;
wire _999_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _1477_ ;
wire _1057_ ;
wire _388_ ;
wire _600_ ;
wire _1286_ ;
wire _197_ ;
wire _1095_ ;
wire _7_ ;
wire _923_ ;
wire _503_ ;
wire _1189_ ;
wire _1401_ ;
wire _732_ ;
wire _312_ ;
wire _48_ ;
wire _1630_ ;
wire _1210_ ;
wire _961_ ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _1724_ ;
wire _1304_ ;
wire _635_ ;
wire _215_ ;
wire _1533_ ;
wire _1113_ ;
wire _864_ ;
wire _444_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0  ;
wire _1762_ ;
wire _1342_ ;
wire _673_ ;
wire _253_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_reg  ;
wire _729_ ;
wire _309_ ;
wire _1571_ ;
wire _1151_ ;
wire _482_ ;
wire _1627_ ;
wire _1207_ ;
wire _958_ ;
wire _538_ ;
wire _118_ ;
wire _1380_ ;
wire _291_ ;
wire _10_ ;
wire _1436_ ;
wire _1016_ ;
wire _767_ ;
wire _347_ ;
wire _1665_ ;
wire _1245_ ;
wire _996_ ;
wire _576_ ;
wire _156_ ;
wire _1474_ ;
wire _1054_ ;
wire _385_ ;
wire _1283_ ;
wire _194_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0  ;
wire _1759_ ;
wire _1339_ ;
wire _1092_ ;
wire _1568_ ;
wire _1148_ ;
wire _899_ ;
wire _479_ ;
wire _1377_ ;
wire _288_ ;
wire _4_ ;
wire _920_ ;
wire _500_ ;
wire _1186_ ;
wire _45_ ;
wire ap_idle ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _1089_ ;
wire _1721_ ;
wire _1301_ ;
wire _632_ ;
wire _212_ ;
wire _1530_ ;
wire _1110_ ;
wire _861_ ;
wire _441_ ;
wire _917_ ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire _1624_ ;
wire _1204_ ;
wire _955_ ;
wire _535_ ;
wire _115_ ;
wire _1433_ ;
wire _1013_ ;
wire _764_ ;
wire _344_ ;
wire _1662_ ;
wire _1242_ ;
wire _993_ ;
wire _573_ ;
wire _153_ ;
wire _1718_ ;
wire _629_ ;
wire _209_ ;
wire _1471_ ;
wire _1051_ ;
wire _382_ ;
wire _1527_ ;
wire _1107_ ;
wire _858_ ;
wire _438_ ;
wire _1280_ ;
wire _191_ ;
wire _1756_ ;
wire _1336_ ;
wire _667_ ;
wire _247_ ;
wire _1565_ ;
wire _1145_ ;
wire _896_ ;
wire _476_ ;
wire _1374_ ;
wire _285_ ;
wire _1_ ;
wire _1183_ ;
wire _1659_ ;
wire _1239_ ;
wire _42_ ;
wire _1468_ ;
wire _1048_ ;
wire _799_ ;
wire _379_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2  ;
wire _1697_ ;
wire _1277_ ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire _1086_ ;
wire _914_ ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _1621_ ;
wire _1201_ ;
wire _952_ ;
wire _532_ ;
wire _112_ ;
wire _1430_ ;
wire _1010_ ;
wire _761_ ;
wire _341_ ;
wire _817_ ;
wire _77_ ;
wire _990_ ;
wire _570_ ;
wire _150_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4  ;
wire _1715_ ;
wire _626_ ;
wire _206_ ;
wire _1524_ ;
wire _1104_ ;
wire _855_ ;
wire _435_ ;
wire _1753_ ;
wire _1333_ ;
wire _664_ ;
wire _244_ ;
wire _1562_ ;
wire _1142_ ;
wire _893_ ;
wire _473_ ;
wire _1618_ ;
wire _949_ ;
wire _529_ ;
wire _109_ ;
wire _1371_ ;
wire _282_ ;
wire _1427_ ;
wire _1007_ ;
wire _758_ ;
wire _338_ ;
wire _1180_ ;
wire _1656_ ;
wire _1236_ ;
wire _987_ ;
wire _567_ ;
wire _147_ ;
wire _1465_ ;
wire _1045_ ;
wire _796_ ;
wire _376_ ;
wire _1694_ ;
wire _1274_ ;
wire _185_ ;
wire _1083_ ;
wire _1559_ ;
wire _1139_ ;
wire _1368_ ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire _1597_ ;
wire _1177_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_int  ;
wire _467__bF$buf0 ;
wire _467__bF$buf1 ;
wire _467__bF$buf2 ;
wire _467__bF$buf3 ;
wire _467__bF$buf4 ;
wire _467__bF$buf5 ;
wire _467__bF$buf6 ;
wire _720_ ;
wire _300_ ;
wire _36_ ;
wire [28:0] q_1_loc_fu_40 ;
wire _814_ ;
wire _74_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1  ;
wire _1027__bF$buf0 ;
wire _1027__bF$buf1 ;
wire _1027__bF$buf2 ;
wire _1027__bF$buf3 ;
wire _1027__bF$buf4 ;
wire _1027__bF$buf5 ;
wire _1712_ ;
wire _623_ ;
wire _203_ ;
wire _1521_ ;
wire _1101_ ;
wire _852_ ;
wire _432_ ;
wire _908_ ;
wire _1750_ ;
wire _1330_ ;
wire _661_ ;
wire _241_ ;
wire _717_ ;
wire _890_ ;
wire _470_ ;
wire _1615_ ;
wire _946_ ;
wire _526_ ;
wire _106_ ;
wire _1424_ ;
wire _1004_ ;
wire _755_ ;
wire _335_ ;
wire _1653_ ;
wire _1233_ ;
wire _984_ ;
wire _564_ ;
wire _144_ ;
wire _1709_ ;
wire _1462_ ;
wire _1042_ ;
wire _793_ ;
wire _373_ ;
wire _1046__bF$buf0 ;
wire _1046__bF$buf1 ;
wire _1046__bF$buf2 ;
wire _1046__bF$buf3 ;
wire _1046__bF$buf4 ;
wire _1046__bF$buf5 ;
wire _1046__bF$buf6 ;
wire _1046__bF$buf7 ;
wire _1518_ ;
wire _849_ ;
wire _429_ ;
wire _1691_ ;
wire _1271_ ;
wire _182_ ;
wire _1050__bF$buf0 ;
wire _1050__bF$buf1 ;
wire _1050__bF$buf2 ;
wire _1050__bF$buf3 ;
wire _1050__bF$buf4 ;
wire _1050__bF$buf5 ;
wire _1747_ ;
wire _1327_ ;
wire _658_ ;
wire _238_ ;
wire _1080_ ;
wire _1556_ ;
wire _1136_ ;
wire _887_ ;
wire _467_ ;
wire _1365_ ;
wire _696_ ;
wire _276_ ;
wire _1594_ ;
wire _1174_ ;
wire _33_ ;
wire _1459_ ;
wire _1039_ ;
wire _1688_ ;
wire _1268_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire _1497_ ;
wire _1077_ ;
wire _620_ ;
wire _200_ ;
wire _905_ ;
wire _714_ ;
wire _1612_ ;
wire _943_ ;
wire _523_ ;
wire _103_ ;
wire _1421_ ;
wire _1001_ ;
wire _752_ ;
wire _332_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5  ;
wire _808_ ;
wire _68_ ;
wire _1650_ ;
wire _1230_ ;
wire _981_ ;
wire _561_ ;
wire _141_ ;
wire _1706_ ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _1515_ ;
wire _846_ ;
wire _426_ ;
wire _1744_ ;
wire _1324_ ;
wire _655_ ;
wire _235_ ;
wire _1553_ ;
wire _1133_ ;
wire _884_ ;
wire _464_ ;
wire _1609_ ;
wire _1362_ ;
wire _693_ ;
wire _273_ ;
wire _1418_ ;
wire _749_ ;
wire _329_ ;
wire _1591_ ;
wire _1171_ ;
wire _1647_ ;
wire _1227_ ;
wire _978_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _1456_ ;
wire _1036_ ;
wire _787_ ;
wire _367_ ;
wire _1685_ ;
wire _1265_ ;
wire _596_ ;
wire _176_ ;
wire _1494_ ;
wire _1074_ ;
wire [27:0] _1779_ ;
wire _1359_ ;
wire _902_ ;
wire _1588_ ;
wire _1168_ ;
wire _499_ ;
wire _711_ ;
wire _1397_ ;
wire _27_ ;
wire _940_ ;
wire _520_ ;
wire _100_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2  ;
wire _805_ ;
wire _65_ ;
wire _1703_ ;
wire _614_ ;
wire _1512_ ;
wire _843_ ;
wire _423_ ;
wire _1741_ ;
wire _1321_ ;
wire _652_ ;
wire _232_ ;
wire _708_ ;
wire _1550_ ;
wire _1130_ ;
wire _881_ ;
wire _461_ ;
wire _1606_ ;
wire _937_ ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _1415_ ;
wire _746_ ;
wire _326_ ;
wire _1644_ ;
wire _1224_ ;
wire _975_ ;
wire _555_ ;
wire _135_ ;
wire _1453_ ;
wire _1033_ ;
wire _784_ ;
wire _364_ ;
wire _1509_ ;
wire _1682_ ;
wire _1262_ ;
wire _593_ ;
wire _173_ ;
wire _1738_ ;
wire _1318_ ;
wire _649_ ;
wire _229_ ;
wire _1491_ ;
wire _1071_ ;
wire _1547_ ;
wire _1127_ ;
wire _878_ ;
wire _458_ ;
wire _1776_ ;
wire _1356_ ;
wire _687_ ;
wire _267_ ;
wire ap_CS_fsm_state1_bF$buf0 ;
wire ap_CS_fsm_state1_bF$buf1 ;
wire ap_CS_fsm_state1_bF$buf2 ;
wire ap_CS_fsm_state1_bF$buf3 ;
wire ap_CS_fsm_state1_bF$buf4 ;
wire ap_CS_fsm_state1_bF$buf5 ;
wire ap_CS_fsm_state1_bF$buf6 ;
wire _1585_ ;
wire _1165_ ;
wire _496_ ;
wire _1394_ ;
wire _24_ ;
wire _1679_ ;
wire _1259_ ;
wire _802_ ;
wire _62_ ;
wire _1488_ ;
wire _1068_ ;
wire _399_ ;
wire _1700_ ;
wire _611_ ;
wire _1297_ ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire _1603_ ;
wire _934_ ;
wire _514_ ;
wire _1412_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _1641_ ;
wire _1221_ ;
wire _972_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _1450_ ;
wire _1030_ ;
wire _781_ ;
wire _361_ ;
wire _1506_ ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire _1735_ ;
wire _1315_ ;
wire _646_ ;
wire _226_ ;
wire _1544_ ;
wire _1124_ ;
wire _875_ ;
wire _455_ ;
wire _1773_ ;
wire _1353_ ;
wire _684_ ;
wire _264_ ;
wire _1409_ ;
wire _1582_ ;
wire _1162_ ;
wire _493_ ;
wire _1063__bF$buf0 ;
wire _1063__bF$buf1 ;
wire _1063__bF$buf2 ;
wire _1063__bF$buf3 ;
wire _1063__bF$buf4 ;
wire _1638_ ;
wire _1218_ ;
wire _969_ ;
wire _549_ ;
wire _129_ ;
wire _1391_ ;
wire _21_ ;
wire _1447_ ;
wire _1027_ ;
wire _778_ ;
wire _358_ ;
wire _1676_ ;
wire _1256_ ;
wire _587_ ;
wire _167_ ;
wire _1485_ ;
wire _1065_ ;
wire _396_ ;
wire _1294_ ;
wire _1579_ ;
wire _1159_ ;
wire _702_ ;
wire _1388_ ;
wire _299_ ;
wire _18_ ;
wire _1600_ ;
wire _931_ ;
wire _511_ ;
wire _1197_ ;
wire _740_ ;
wire _320_ ;
wire _56_ ;
wire ap_clk_bF$buf10 ;
wire ap_clk_bF$buf11 ;
wire ap_clk_bF$buf12 ;
wire _605_ ;
wire _1503_ ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire _1732_ ;
wire _1312_ ;
wire _643_ ;
wire _223_ ;
wire _1541_ ;
wire _1121_ ;
wire _872_ ;
wire _452_ ;
wire _928_ ;
wire _508_ ;
wire _1770_ ;
wire _1350_ ;
wire _681_ ;
wire _261_ ;
wire _1406_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _1635_ ;
wire _1215_ ;
wire _966_ ;
wire _546_ ;
wire _126_ ;
wire _1444_ ;
wire _1024_ ;
wire _775_ ;
wire _355_ ;
wire _1673_ ;
wire _1253_ ;
wire _584_ ;
wire _164_ ;
wire _1729_ ;
wire _1309_ ;
wire _1482_ ;
wire _1062_ ;
wire _393_ ;
wire _1538_ ;
wire _1118_ ;
wire _869_ ;
wire _449_ ;
wire _1291_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5  ;
wire _1767_ ;
wire _1347_ ;
wire _678_ ;
wire _258_ ;
wire [30:0] s_5_loc_fu_48 ;
wire _1576_ ;
wire _1156_ ;
wire _487_ ;
wire _1385_ ;
wire _296_ ;
wire _15_ ;
wire _1194_ ;
wire _53_ ;
wire _1479_ ;
wire _1059_ ;
wire _602_ ;
wire _1288_ ;
wire _199_ ;
wire _1500_ ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _1097_ ;
wire _640_ ;
wire _220_ ;
wire _9_ ;
wire _925_ ;
wire _505_ ;
wire _1403_ ;
wire _734_ ;
wire _314_ ;
wire [30:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out  ;
wire _1632_ ;
wire _1212_ ;
wire _963_ ;
wire _543_ ;
wire _123_ ;
wire _1441_ ;
wire _1021_ ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire _1670_ ;
wire _1250_ ;
wire _581_ ;
wire _161_ ;
wire _1726_ ;
wire _1306_ ;
wire _637_ ;
wire _217_ ;
wire _390_ ;
wire _1535_ ;
wire _1115_ ;
wire _866_ ;
wire _446_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2  ;
wire _1764_ ;
wire _1344_ ;
wire _675_ ;
wire _255_ ;
wire _1573_ ;
wire _1153_ ;
wire _484_ ;
wire _1629_ ;
wire _1209_ ;
wire _1382_ ;
wire _293_ ;
wire _12_ ;
wire _1438_ ;
wire _1018_ ;
wire _769_ ;
wire _349_ ;
wire _1191_ ;
wire _1667_ ;
wire _1247_ ;
wire _998_ ;
wire _578_ ;
wire _158_ ;
wire [0:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3  ;
wire _50_ ;
wire _1476_ ;
wire _1056_ ;
wire _387_ ;
wire _1285_ ;
wire _196_ ;
wire _1094_ ;
wire _1379_ ;
wire _6_ ;
wire _922_ ;
wire _502_ ;
wire _1188_ ;
wire _1400_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _960_ ;
wire _540_ ;
wire _120_ ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire _1723_ ;
wire _1303_ ;
wire _634_ ;
wire _214_ ;
wire _1532_ ;
wire _1112_ ;
wire _863_ ;
wire _443_ ;
wire _919_ ;
wire _1761_ ;
wire _1341_ ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _1570_ ;
wire _1150_ ;
wire _481_ ;
wire _1626_ ;
wire _1206_ ;
wire _957_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _1435_ ;
wire _1015_ ;
wire _766_ ;
wire _346_ ;
wire _1664_ ;
wire _1244_ ;
wire _995_ ;
wire _575_ ;
wire _155_ ;
wire _1473_ ;
wire _1053_ ;
wire _384_ ;
wire _1529_ ;
wire _1109_ ;
wire _1282_ ;
wire _193_ ;
wire _1758_ ;
wire _1338_ ;
wire _669_ ;
wire _249_ ;
wire _1091_ ;
wire _1567_ ;
wire _1147_ ;
wire _898_ ;
wire _478_ ;
wire _1376_ ;
wire _287_ ;
wire _3_ ;
wire _1185_ ;
wire _44_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4  ;
wire _1699_ ;
wire _1279_ ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _1088_ ;
wire _1720_ ;
wire _1300_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _916_ ;
wire _725_ ;
wire _305_ ;
wire ap_ready ;
wire _1623_ ;
wire _1203_ ;
wire _954_ ;
wire _534_ ;
wire _114_ ;
wire _1432_ ;
wire _1012_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _1661_ ;
wire _1241_ ;
wire _992_ ;
wire _572_ ;
wire _152_ ;
wire _1717_ ;
wire _628_ ;
wire _208_ ;
wire _1470_ ;
wire _1050_ ;
wire _381_ ;
wire _1526_ ;
wire _1106_ ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _1755_ ;
wire _1335_ ;
wire _666_ ;
wire _246_ ;
wire ap_clk_bF$buf0 ;
wire ap_clk_bF$buf1 ;
wire ap_clk_bF$buf2 ;
wire ap_clk_bF$buf3 ;
wire ap_clk_bF$buf4 ;
wire ap_clk_bF$buf5 ;
wire ap_clk_bF$buf6 ;
wire ap_clk_bF$buf7 ;
wire ap_clk_bF$buf8 ;
wire ap_clk_bF$buf9 ;
wire _1564_ ;
wire _1144_ ;
wire _895_ ;
wire _475_ ;
wire _1373_ ;
wire _284_ ;
wire _0_ ;
wire _1429_ ;
wire _1009_ ;
wire _1182_ ;
wire _1658_ ;
wire _1238_ ;
wire _989_ ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _1467_ ;
wire _1047_ ;
wire _798_ ;
wire _378_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1  ;
wire _1696_ ;
wire _1276_ ;
wire _187_ ;
wire _1085_ ;
wire _913_ ;
wire _1599_ ;
wire _1179_ ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _1620_ ;
wire _1200_ ;
wire _951_ ;
wire _531_ ;
wire _111_ ;
wire _760_ ;
wire _340_ ;
wire _436__bF$buf0 ;
wire _436__bF$buf1 ;
wire _436__bF$buf2 ;
wire _436__bF$buf3 ;
wire _436__bF$buf4 ;
wire _436__bF$buf5 ;
wire _436__bF$buf6 ;
wire _816_ ;
wire _76_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3  ;
wire _1714_ ;
wire _625_ ;
wire _205_ ;
wire [27:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90  ;
wire _1523_ ;
wire _1103_ ;
wire _854_ ;
wire _434_ ;
wire _1752_ ;
wire _1332_ ;
wire _663_ ;
wire _243_ ;
wire _719_ ;
wire _1561_ ;
wire _1141_ ;
wire _892_ ;
wire _472_ ;
wire _1617_ ;
wire _948_ ;
wire _528_ ;
wire _108_ ;
wire _1370_ ;
wire _281_ ;
wire _1426_ ;
wire _1006_ ;
wire _757_ ;
wire _337_ ;
wire _1655_ ;
wire _1235_ ;
wire _986_ ;
wire _566_ ;
wire _146_ ;
wire _1464_ ;
wire _1044_ ;
wire _948__bF$buf0 ;
wire _948__bF$buf1 ;
wire _948__bF$buf2 ;
wire _948__bF$buf3 ;
wire _948__bF$buf4 ;
wire _795_ ;
wire _375_ ;
wire _1693_ ;
wire _1273_ ;
wire _184_ ;
wire _1749_ ;
wire _1329_ ;
wire _1082_ ;
wire _1558_ ;
wire _1138_ ;
wire _889_ ;
wire _469_ ;
wire _1367_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire _1596_ ;
wire _1176_ ;
wire _35_ ;
wire _813_ ;
wire _73_ ;
wire _1499_ ;
wire _1079_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0  ;
wire _1711_ ;
wire _622_ ;
wire _202_ ;
wire _1520_ ;
wire _1100_ ;
wire [27:0] p_v_loc_fu_44 ;
wire _851_ ;
wire _431_ ;
wire _1034__bF$buf0 ;
wire _1034__bF$buf1 ;
wire _1034__bF$buf2 ;
wire _1034__bF$buf3 ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire _716_ ;
wire _1614_ ;
wire _945_ ;
wire _525_ ;
wire _105_ ;
wire _1423_ ;
wire _1003_ ;
wire _754_ ;
wire _334_ ;
wire _1652_ ;
wire _1232_ ;
wire _983_ ;
wire _563_ ;
wire _143_ ;
wire _1708_ ;
wire _619_ ;
wire _1461_ ;
wire _1041_ ;
wire _792_ ;
wire _372_ ;
wire _1517_ ;
wire _848_ ;
wire _428_ ;
wire _1690_ ;
wire _1270_ ;
wire _181_ ;
wire _1746_ ;
wire _1326_ ;
wire _657_ ;
wire _237_ ;
wire _1555_ ;
wire _1135_ ;
wire _886_ ;
wire _466_ ;
wire _1364_ ;
wire _695_ ;
wire _275_ ;
wire _955__bF$buf0 ;
wire _955__bF$buf1 ;
wire _955__bF$buf2 ;
wire _955__bF$buf3 ;
wire _955__bF$buf4 ;
wire _1593_ ;
wire _1173_ ;
wire _151__bF$buf0 ;
wire _151__bF$buf1 ;
wire _151__bF$buf2 ;
wire _151__bF$buf3 ;
wire _151__bF$buf4 ;
wire _151__bF$buf5 ;
wire _151__bF$buf6 ;
wire _1649_ ;
wire _1229_ ;
wire _32_ ;
wire _1458_ ;
wire _1038_ ;
wire _789_ ;
wire _369_ ;
wire _1022__bF$buf0 ;
wire _1022__bF$buf1 ;
wire _1022__bF$buf2 ;
wire _1022__bF$buf3 ;
wire _1022__bF$buf4 ;
wire _1022__bF$buf5 ;
wire _1022__bF$buf6 ;
wire _1687_ ;
wire _1267_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire _1496_ ;
wire _1076_ ;
wire _904_ ;
wire _713_ ;
wire _1399_ ;
wire _29_ ;
wire _1611_ ;
wire _942_ ;
wire _522_ ;
wire _102_ ;
wire _1420_ ;
wire _1000_ ;
wire _751_ ;
wire _331_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4  ;
wire _807_ ;
wire _67_ ;
wire _980_ ;
wire _560_ ;
wire _140_ ;
wire _1705_ ;
wire _616_ ;
wire _1514_ ;
wire _845_ ;
wire _425_ ;
wire _1743_ ;
wire _1323_ ;
wire _654_ ;
wire _234_ ;
wire _1552_ ;
wire _1132_ ;
wire _883_ ;
wire _463_ ;
wire [23:0] in_val ;
wire _1608_ ;
wire _939_ ;
wire _519_ ;
wire _1361_ ;
wire _692_ ;
wire _272_ ;
wire _1417_ ;
wire _748_ ;
wire _328_ ;
wire _1590_ ;
wire _1170_ ;
wire _1646_ ;
wire _1226_ ;
wire _977_ ;
wire _557_ ;
wire _137_ ;
wire _1455_ ;
wire _1035_ ;
wire _786_ ;
wire _366_ ;
wire _1684_ ;
wire _1264_ ;
wire _595_ ;
wire _175_ ;
wire _1493_ ;
wire _1073_ ;
wire _1549_ ;
wire _1129_ ;
wire _1778_ ;
wire _1358_ ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _1587_ ;
wire _1167_ ;
wire _498_ ;
wire _710_ ;
wire _1396_ ;
wire _26_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1  ;
wire _804_ ;
wire _64_ ;
wire _1702_ ;
wire _613_ ;
wire _1299_ ;
wire _1511_ ;
wire _842_ ;
wire _422_ ;
wire _1740_ ;
wire _1320_ ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _1605_ ;
wire _936_ ;
wire _516_ ;
wire _1414_ ;
wire _745_ ;
wire _325_ ;
wire _1643_ ;
wire _1223_ ;
wire _974_ ;
wire _554_ ;
wire _134_ ;
wire _1452_ ;
wire _1032_ ;
wire _783_ ;
wire _363_ ;
wire _1508_ ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _1681_ ;
wire _1261_ ;
wire [30:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_1_fu_177_p2  ;
wire _592_ ;
wire _172_ ;
wire _1737_ ;
wire _1317_ ;
wire _648_ ;
wire _228_ ;
wire _1490_ ;
wire _1070_ ;
wire _1546_ ;
wire _1126_ ;
wire _877_ ;
wire _457_ ;
wire _1775_ ;
wire _1355_ ;
wire _686_ ;
wire _266_ ;
wire _1584_ ;
wire _1164_ ;
wire _495_ ;
wire _1393_ ;
wire _23_ ;
wire _1449_ ;
wire _1029_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.flow_control_loop_pipe_sequential_init_U.ap_done_cache  ;
wire [4:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60  ;
wire _1678_ ;
wire _1258_ ;
wire _589_ ;
wire _169_ ;
wire _801_ ;
wire _61_ ;
wire _1487_ ;
wire _1067_ ;
wire _398_ ;
wire _610_ ;
wire _1296_ ;
wire _704_ ;
wire _1602_ ;
wire _933_ ;
wire _513_ ;
wire _1199_ ;
wire _1411_ ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _1640_ ;
wire _1220_ ;
wire _971_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire _780_ ;
wire _360_ ;
wire _1505_ ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _1734_ ;
wire _1314_ ;
wire _645_ ;
wire _225_ ;
wire _1543_ ;
wire _1123_ ;
wire _874_ ;
wire _454_ ;
wire _1772_ ;
wire _1352_ ;
wire _683_ ;
wire _263_ ;
wire _1408_ ;
wire _739_ ;
wire _319_ ;
wire _1581_ ;
wire _1161_ ;
wire _492_ ;
wire _1637_ ;
wire _1217_ ;
wire ap_clk ;
wire _968_ ;
wire _548_ ;
wire _128_ ;
wire _1390_ ;
wire _20_ ;
wire _1446_ ;
wire _1026_ ;
wire _777_ ;
wire _357_ ;
wire grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58_ap_start_reg ;
wire _1675_ ;
wire _1255_ ;
wire _586_ ;
wire _166_ ;
wire _1484_ ;
wire _1064_ ;
wire _395_ ;
wire _1293_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7  ;
wire _1769_ ;
wire _1349_ ;
wire _1578_ ;
wire _1158_ ;
wire _489_ ;
wire _701_ ;
wire _1387_ ;
wire _298_ ;
wire _17_ ;
wire _930_ ;
wire _510_ ;
wire _1196_ ;
wire _55_ ;
wire _604_ ;
wire _1502_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _1099_ ;
wire _1731_ ;
wire _1311_ ;
wire _642_ ;
wire _222_ ;
wire _1540_ ;
wire _1120_ ;
wire _871_ ;
wire _451_ ;
wire _927_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire _1405_ ;
wire _736_ ;
wire _316_ ;
wire _1634_ ;
wire _1214_ ;
wire _965_ ;
wire _545_ ;
wire _125_ ;
wire _1443_ ;
wire _1023_ ;
wire _774_ ;
wire _354_ ;
wire _1672_ ;
wire _1252_ ;
wire _583_ ;
wire _163_ ;
wire _1728_ ;
wire _1308_ ;
wire _639_ ;
wire _219_ ;
wire _1481_ ;
wire _1061_ ;
wire _392_ ;
wire _1537_ ;
wire _1117_ ;
wire _868_ ;
wire _448_ ;
wire _1290_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4  ;
wire _1766_ ;
wire _1346_ ;
wire _677_ ;
wire _257_ ;
wire _1575_ ;
wire _1155_ ;
wire _486_ ;
wire _1384_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.flow_control_loop_pipe_sequential_init_U.ap_loop_init_int  ;
wire _295_ ;
wire _14_ ;
wire _1193_ ;
wire _1669_ ;
wire _1249_ ;
wire _52_ ;
wire _1478_ ;
wire _1058_ ;
wire _389_ ;
wire _601_ ;
wire [28:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72  ;
wire _1287_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _1096_ ;
wire _8_ ;
wire _924_ ;
wire _504_ ;
wire _1402_ ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _1631_ ;
wire _1211_ ;
wire _962_ ;
wire _542_ ;
wire _122_ ;
wire _1440_ ;
wire _1020_ ;
wire _771_ ;
wire _351_ ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire _580_ ;
wire _160_ ;
wire _1725_ ;
wire _1305_ ;
wire _636_ ;
wire _216_ ;
wire _1534_ ;
wire _1114_ ;
wire _865_ ;
wire _445_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1  ;
wire _1763_ ;
wire _1343_ ;
wire _674_ ;
wire _254_ ;
wire _1572_ ;
wire _1152_ ;
wire _483_ ;
wire _1628_ ;
wire _1208_ ;
wire _959_ ;
wire _539_ ;
wire _119_ ;
wire _1381_ ;
wire _292_ ;
wire _11_ ;
wire _1437_ ;
wire _1017_ ;
wire _768_ ;
wire _348_ ;
wire _1190_ ;
wire _1666_ ;
wire _1246_ ;
wire _997_ ;
wire _577_ ;
wire _157_ ;
wire _1475_ ;
wire _1055_ ;
wire _386_ ;
wire _1284_ ;
wire _195_ ;
wire _1093_ ;
wire _1569_ ;
wire _1149_ ;
wire _1378_ ;
wire _289_ ;
wire _5_ ;
wire _921_ ;
wire _501_ ;
wire _1187_ ;
wire _730_ ;
wire _310_ ;
wire _46_ ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _1722_ ;
wire _1302_ ;
wire _633_ ;
wire _213_ ;
wire _1531_ ;
wire _1111_ ;
wire _1064__bF$buf0 ;
wire _1064__bF$buf1 ;
wire _1064__bF$buf2 ;
wire _862_ ;
wire _1064__bF$buf3 ;
wire _442_ ;
wire _1064__bF$buf4 ;
wire _1064__bF$buf5 ;
wire _918_ ;
wire _1760_ ;
wire _1340_ ;
wire _671_ ;
wire _251_ ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire _1625_ ;
wire _1205_ ;
wire _956_ ;
wire _536_ ;
wire _116_ ;
wire _1434_ ;
wire _1014_ ;
wire _765_ ;
wire _345_ ;
wire _1663_ ;
wire _1243_ ;
wire _994_ ;
wire _574_ ;
wire _154_ ;
wire _1719_ ;
wire _1472_ ;
wire _1052_ ;
wire _383_ ;
wire _1528_ ;
wire _1108_ ;
wire _859_ ;
wire _439_ ;
wire _1281_ ;
wire _192_ ;
wire _1757_ ;
wire _1337_ ;
wire _668_ ;
wire _248_ ;
wire _1090_ ;
wire _1566_ ;
wire _1146_ ;
wire _897_ ;
wire _477_ ;
wire _1375_ ;
wire _286_ ;
wire _2_ ;
wire _1184_ ;
wire _43_ ;
wire _1469_ ;
wire _1049_ ;
wire _1052__bF$buf0 ;
wire _1052__bF$buf1 ;
wire _1052__bF$buf2 ;
wire _1052__bF$buf3 ;
wire _1052__bF$buf4 ;
wire _1052__bF$buf5 ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3  ;
wire _1698_ ;
wire _1278_ ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire _1087_ ;
wire _630_ ;
wire _210_ ;
wire _915_ ;
wire _724_ ;
wire _304_ ;
wire _1622_ ;
wire _1202_ ;
wire _953_ ;
wire _533_ ;
wire _113_ ;
wire _1431_ ;
wire _1011_ ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _1660_ ;
wire _1240_ ;
wire _991_ ;
wire _571_ ;
wire _151_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5  ;
wire _1716_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire _1525_ ;
wire _1105_ ;
wire _856_ ;
wire _436_ ;
wire _1754_ ;
wire _1334_ ;
wire _665_ ;
wire _245_ ;
wire _1563_ ;
wire _1143_ ;
wire _894_ ;
wire _474_ ;
wire _1619_ ;
wire _1372_ ;
wire _283_ ;
wire _1428_ ;
wire _1008_ ;
wire _759_ ;
wire _339_ ;
wire _1181_ ;
wire _1657_ ;
wire _1237_ ;
wire _988_ ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _1466_ ;
wire _1046_ ;
wire _797_ ;
wire _377_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0  ;
wire _1695_ ;
wire _1275_ ;
wire _186_ ;
wire _1084_ ;
wire _1369_ ;
wire _912_ ;
wire _1598_ ;
wire _1178_ ;
wire _721_ ;
wire _301_ ;
wire ap_CS_fsm_state1 ;
wire ap_CS_fsm_state2 ;
wire _37_ ;
wire _950_ ;
wire _530_ ;
wire _110_ ;
wire _815_ ;
wire _75_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2  ;
wire _1713_ ;
wire _624_ ;
wire _204_ ;
wire _1522_ ;
wire _1102_ ;
wire _853_ ;
wire _433_ ;
wire _909_ ;
wire _1751_ ;
wire _1331_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _1560_ ;
wire _1140_ ;
wire _891_ ;
wire _471_ ;
wire _1616_ ;
wire ap_start ;
wire _947_ ;
wire _527_ ;
wire _107_ ;
wire _280_ ;
wire _1425_ ;
wire _1005_ ;
wire _756_ ;
wire _336_ ;
wire _1654_ ;
wire _1234_ ;
wire _985_ ;
wire _565_ ;
wire _145_ ;
wire _1463_ ;
wire _1043_ ;
wire _794_ ;
wire _374_ ;
wire [27:0] ap_return ;
wire _1519_ ;
wire _1692_ ;
wire _1272_ ;
wire _183_ ;
wire _1748_ ;
wire _1328_ ;
wire _659_ ;
wire _239_ ;
wire _1081_ ;
wire _1557_ ;
wire _1137_ ;
wire _888_ ;
wire _468_ ;
wire _1366_ ;
wire _697_ ;
wire _277_ ;
wire _1595_ ;
wire _1175_ ;
wire _34_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done  ;
wire _1689_ ;
wire _1269_ ;
wire _812_ ;
wire _72_ ;
wire _1498_ ;
wire _1078_ ;
wire _1710_ ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire [30:0] \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64  ;
wire _1613_ ;
wire _944_ ;
wire _524_ ;
wire _104_ ;
wire _1422_ ;
wire _1002_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _1651_ ;
wire _1231_ ;
wire _982_ ;
wire _562_ ;
wire _142_ ;
wire _1707_ ;
wire _618_ ;
wire _1460_ ;
wire _1040_ ;
wire _791_ ;
wire _371_ ;
wire _1516_ ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _1745_ ;
wire _1325_ ;
wire _656_ ;
wire _236_ ;
wire _1554_ ;
wire _1134_ ;
wire _885_ ;
wire _465_ ;
wire _1363_ ;
wire _694_ ;
wire _274_ ;
wire _1419_ ;
wire _1592_ ;
wire _1172_ ;
wire _1648_ ;
wire _1228_ ;
wire _979_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _1457_ ;
wire _1037_ ;
wire _788_ ;
wire _368_ ;
wire _1686_ ;
wire _1266_ ;
wire _597_ ;
wire _177_ ;
wire _1495_ ;
wire _1075_ ;
wire _903_ ;
wire _1589_ ;
wire _1169_ ;
wire _712_ ;
wire _1398_ ;
wire _28_ ;
wire _1610_ ;
wire _941_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3  ;
wire _806_ ;
wire _66_ ;
wire _1704_ ;
wire _615_ ;
wire _1513_ ;
wire _844_ ;
wire _424_ ;
wire _1742_ ;
wire _1322_ ;
wire _653_ ;
wire _233_ ;
wire _709_ ;
wire _1551_ ;
wire _1131_ ;
wire _882_ ;
wire _462_ ;
wire _1607_ ;
wire _938_ ;
wire _518_ ;
wire _1360_ ;
wire _691_ ;
wire _271_ ;
wire _1416_ ;
wire _747_ ;
wire _327_ ;
wire _1645_ ;
wire _1225_ ;
wire _976_ ;
wire _556_ ;
wire _136_ ;
wire _1454_ ;
wire _1034_ ;
wire _785_ ;
wire _365_ ;
wire _1683_ ;
wire _1263_ ;
wire _594_ ;
wire _174_ ;
wire _1739_ ;
wire _1319_ ;
wire _1492_ ;
wire _1072_ ;
wire _1548_ ;
wire _1128_ ;
wire _879_ ;
wire _459_ ;
wire _1777_ ;
wire _1357_ ;
wire _688_ ;
wire _268_ ;
wire ap_rst ;
wire _339__bF$buf0 ;
wire _339__bF$buf1 ;
wire _339__bF$buf2 ;
wire _339__bF$buf3 ;
wire _339__bF$buf4 ;
wire _339__bF$buf5 ;
wire _339__bF$buf6 ;
wire _900_ ;
wire _1586_ ;
wire _1166_ ;
wire _497_ ;
wire _1395_ ;
wire _25_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0  ;
wire _803_ ;
wire _63_ ;
wire _1489_ ;
wire _1069_ ;
wire _1701_ ;
wire _612_ ;
wire _1298_ ;
wire _1510_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_enable_reg_pp0_iter1  ;
wire _706_ ;
wire _1604_ ;
wire _935_ ;
wire _515_ ;
wire _1413_ ;
wire _744_ ;
wire _324_ ;
wire _1087__bF$buf0 ;
wire _1087__bF$buf1 ;
wire _1087__bF$buf2 ;
wire _1087__bF$buf3 ;
wire _1087__bF$buf4 ;
wire _1642_ ;
wire _1222_ ;
wire _973_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _1451_ ;
wire _1031_ ;
wire \grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init  ;
wire _782_ ;
wire _362_ ;
wire _1507_ ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _1680_ ;
wire _1260_ ;
wire _591_ ;
wire _171_ ;
wire _1736_ ;
wire _1316_ ;
wire _647_ ;
wire _227_ ;
wire _1545_ ;
wire _1125_ ;
wire _876_ ;
wire _456_ ;
wire _1774_ ;
wire _1354_ ;
wire _685_ ;
wire _265_ ;
wire _1583_ ;
wire _1163_ ;
wire _494_ ;
wire _1639_ ;
wire _1219_ ;
wire _1392_ ;
wire _22_ ;
wire _1448_ ;
wire _1028_ ;
wire _779_ ;
wire _359_ ;

BUFX2 BUFX2_insert144 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 )
);

BUFX2 BUFX2_insert143 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 )
);

BUFX2 BUFX2_insert142 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 )
);

BUFX2 BUFX2_insert141 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 )
);

BUFX2 BUFX2_insert140 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 )
);

BUFX2 BUFX2_insert139 (
    .A(_1034_),
    .Y(_1034__bF$buf0)
);

BUFX2 BUFX2_insert138 (
    .A(_1034_),
    .Y(_1034__bF$buf1)
);

BUFX2 BUFX2_insert137 (
    .A(_1034_),
    .Y(_1034__bF$buf2)
);

BUFX2 BUFX2_insert136 (
    .A(_1034_),
    .Y(_1034__bF$buf3)
);

BUFX2 BUFX2_insert135 (
    .A(_941_),
    .Y(_941__bF$buf0)
);

BUFX2 BUFX2_insert134 (
    .A(_941_),
    .Y(_941__bF$buf1)
);

BUFX2 BUFX2_insert133 (
    .A(_941_),
    .Y(_941__bF$buf2)
);

BUFX2 BUFX2_insert132 (
    .A(_941_),
    .Y(_941__bF$buf3)
);

BUFX2 BUFX2_insert131 (
    .A(_941_),
    .Y(_941__bF$buf4)
);

BUFX2 BUFX2_insert130 (
    .A(_941_),
    .Y(_941__bF$buf5)
);

BUFX2 BUFX2_insert129 (
    .A(_941_),
    .Y(_941__bF$buf6)
);

BUFX2 BUFX2_insert128 (
    .A(_941_),
    .Y(_941__bF$buf7)
);

BUFX2 BUFX2_insert127 (
    .A(_941_),
    .Y(_941__bF$buf8)
);

BUFX2 BUFX2_insert126 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf0)
);

BUFX2 BUFX2_insert125 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf1)
);

BUFX2 BUFX2_insert124 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf2)
);

BUFX2 BUFX2_insert123 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf3)
);

BUFX2 BUFX2_insert122 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf4)
);

BUFX2 BUFX2_insert121 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf5)
);

BUFX2 BUFX2_insert120 (
    .A(ap_CS_fsm_state1),
    .Y(ap_CS_fsm_state1_bF$buf6)
);

BUFX2 BUFX2_insert119 (
    .A(_1046_),
    .Y(_1046__bF$buf0)
);

BUFX2 BUFX2_insert118 (
    .A(_1046_),
    .Y(_1046__bF$buf1)
);

BUFX2 BUFX2_insert117 (
    .A(_1046_),
    .Y(_1046__bF$buf2)
);

BUFX2 BUFX2_insert116 (
    .A(_1046_),
    .Y(_1046__bF$buf3)
);

BUFX2 BUFX2_insert115 (
    .A(_1046_),
    .Y(_1046__bF$buf4)
);

BUFX2 BUFX2_insert114 (
    .A(_1046_),
    .Y(_1046__bF$buf5)
);

BUFX2 BUFX2_insert113 (
    .A(_1046_),
    .Y(_1046__bF$buf6)
);

BUFX2 BUFX2_insert112 (
    .A(_1046_),
    .Y(_1046__bF$buf7)
);

BUFX2 BUFX2_insert111 (
    .A(_339_),
    .Y(_339__bF$buf0)
);

BUFX2 BUFX2_insert110 (
    .A(_339_),
    .Y(_339__bF$buf1)
);

BUFX2 BUFX2_insert109 (
    .A(_339_),
    .Y(_339__bF$buf2)
);

BUFX2 BUFX2_insert108 (
    .A(_339_),
    .Y(_339__bF$buf3)
);

BUFX2 BUFX2_insert107 (
    .A(_339_),
    .Y(_339__bF$buf4)
);

BUFX2 BUFX2_insert106 (
    .A(_339_),
    .Y(_339__bF$buf5)
);

BUFX2 BUFX2_insert105 (
    .A(_339_),
    .Y(_339__bF$buf6)
);

BUFX2 BUFX2_insert104 (
    .A(_436_),
    .Y(_436__bF$buf0)
);

BUFX2 BUFX2_insert103 (
    .A(_436_),
    .Y(_436__bF$buf1)
);

BUFX2 BUFX2_insert102 (
    .A(_436_),
    .Y(_436__bF$buf2)
);

BUFX2 BUFX2_insert101 (
    .A(_436_),
    .Y(_436__bF$buf3)
);

BUFX2 BUFX2_insert100 (
    .A(_436_),
    .Y(_436__bF$buf4)
);

BUFX2 BUFX2_insert99 (
    .A(_436_),
    .Y(_436__bF$buf5)
);

BUFX2 BUFX2_insert98 (
    .A(_436_),
    .Y(_436__bF$buf6)
);

BUFX2 BUFX2_insert97 (
    .A(_151_),
    .Y(_151__bF$buf0)
);

BUFX2 BUFX2_insert96 (
    .A(_151_),
    .Y(_151__bF$buf1)
);

BUFX2 BUFX2_insert95 (
    .A(_151_),
    .Y(_151__bF$buf2)
);

BUFX2 BUFX2_insert94 (
    .A(_151_),
    .Y(_151__bF$buf3)
);

BUFX2 BUFX2_insert93 (
    .A(_151_),
    .Y(_151__bF$buf4)
);

BUFX2 BUFX2_insert92 (
    .A(_151_),
    .Y(_151__bF$buf5)
);

BUFX2 BUFX2_insert91 (
    .A(_151_),
    .Y(_151__bF$buf6)
);

BUFX2 BUFX2_insert90 (
    .A(_1087_),
    .Y(_1087__bF$buf0)
);

BUFX2 BUFX2_insert89 (
    .A(_1087_),
    .Y(_1087__bF$buf1)
);

BUFX2 BUFX2_insert88 (
    .A(_1087_),
    .Y(_1087__bF$buf2)
);

BUFX2 BUFX2_insert87 (
    .A(_1087_),
    .Y(_1087__bF$buf3)
);

BUFX2 BUFX2_insert86 (
    .A(_1087_),
    .Y(_1087__bF$buf4)
);

BUFX2 BUFX2_insert85 (
    .A(_1052_),
    .Y(_1052__bF$buf0)
);

BUFX2 BUFX2_insert84 (
    .A(_1052_),
    .Y(_1052__bF$buf1)
);

BUFX2 BUFX2_insert83 (
    .A(_1052_),
    .Y(_1052__bF$buf2)
);

BUFX2 BUFX2_insert82 (
    .A(_1052_),
    .Y(_1052__bF$buf3)
);

BUFX2 BUFX2_insert81 (
    .A(_1052_),
    .Y(_1052__bF$buf4)
);

BUFX2 BUFX2_insert80 (
    .A(_1052_),
    .Y(_1052__bF$buf5)
);

BUFX2 BUFX2_insert79 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 )
);

BUFX2 BUFX2_insert78 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 )
);

BUFX2 BUFX2_insert77 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 )
);

BUFX2 BUFX2_insert76 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 )
);

BUFX2 BUFX2_insert75 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 )
);

BUFX2 BUFX2_insert74 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 )
);

BUFX2 BUFX2_insert73 (
    .A(_1064_),
    .Y(_1064__bF$buf0)
);

BUFX2 BUFX2_insert72 (
    .A(_1064_),
    .Y(_1064__bF$buf1)
);

BUFX2 BUFX2_insert71 (
    .A(_1064_),
    .Y(_1064__bF$buf2)
);

BUFX2 BUFX2_insert70 (
    .A(_1064_),
    .Y(_1064__bF$buf3)
);

BUFX2 BUFX2_insert69 (
    .A(_1064_),
    .Y(_1064__bF$buf4)
);

BUFX2 BUFX2_insert68 (
    .A(_1064_),
    .Y(_1064__bF$buf5)
);

CLKBUF1 CLKBUF1_insert67 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert66 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert65 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert64 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert63 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf4)
);

CLKBUF1 CLKBUF1_insert62 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf5)
);

CLKBUF1 CLKBUF1_insert61 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf6)
);

CLKBUF1 CLKBUF1_insert60 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf7)
);

CLKBUF1 CLKBUF1_insert59 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf8)
);

CLKBUF1 CLKBUF1_insert58 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf9)
);

CLKBUF1 CLKBUF1_insert57 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf10)
);

CLKBUF1 CLKBUF1_insert56 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf11)
);

CLKBUF1 CLKBUF1_insert55 (
    .A(ap_clk),
    .Y(ap_clk_bF$buf12)
);

BUFX2 BUFX2_insert54 (
    .A(_948_),
    .Y(_948__bF$buf0)
);

BUFX2 BUFX2_insert53 (
    .A(_948_),
    .Y(_948__bF$buf1)
);

BUFX2 BUFX2_insert52 (
    .A(_948_),
    .Y(_948__bF$buf2)
);

BUFX2 BUFX2_insert51 (
    .A(_948_),
    .Y(_948__bF$buf3)
);

BUFX2 BUFX2_insert50 (
    .A(_948_),
    .Y(_948__bF$buf4)
);

BUFX2 BUFX2_insert49 (
    .A(_1050_),
    .Y(_1050__bF$buf0)
);

BUFX2 BUFX2_insert48 (
    .A(_1050_),
    .Y(_1050__bF$buf1)
);

BUFX2 BUFX2_insert47 (
    .A(_1050_),
    .Y(_1050__bF$buf2)
);

BUFX2 BUFX2_insert46 (
    .A(_1050_),
    .Y(_1050__bF$buf3)
);

BUFX2 BUFX2_insert45 (
    .A(_1050_),
    .Y(_1050__bF$buf4)
);

BUFX2 BUFX2_insert44 (
    .A(_1050_),
    .Y(_1050__bF$buf5)
);

BUFX2 BUFX2_insert43 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 )
);

BUFX2 BUFX2_insert42 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 )
);

BUFX2 BUFX2_insert41 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 )
);

BUFX2 BUFX2_insert40 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 )
);

BUFX2 BUFX2_insert39 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 )
);

BUFX2 BUFX2_insert38 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 ),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 )
);

BUFX2 BUFX2_insert37 (
    .A(_1027_),
    .Y(_1027__bF$buf0)
);

BUFX2 BUFX2_insert36 (
    .A(_1027_),
    .Y(_1027__bF$buf1)
);

BUFX2 BUFX2_insert35 (
    .A(_1027_),
    .Y(_1027__bF$buf2)
);

BUFX2 BUFX2_insert34 (
    .A(_1027_),
    .Y(_1027__bF$buf3)
);

BUFX2 BUFX2_insert33 (
    .A(_1027_),
    .Y(_1027__bF$buf4)
);

BUFX2 BUFX2_insert32 (
    .A(_1027_),
    .Y(_1027__bF$buf5)
);

BUFX2 BUFX2_insert31 (
    .A(_467_),
    .Y(_467__bF$buf0)
);

BUFX2 BUFX2_insert30 (
    .A(_467_),
    .Y(_467__bF$buf1)
);

BUFX2 BUFX2_insert29 (
    .A(_467_),
    .Y(_467__bF$buf2)
);

BUFX2 BUFX2_insert28 (
    .A(_467_),
    .Y(_467__bF$buf3)
);

BUFX2 BUFX2_insert27 (
    .A(_467_),
    .Y(_467__bF$buf4)
);

BUFX2 BUFX2_insert26 (
    .A(_467_),
    .Y(_467__bF$buf5)
);

BUFX2 BUFX2_insert25 (
    .A(_467_),
    .Y(_467__bF$buf6)
);

BUFX2 BUFX2_insert24 (
    .A(_955_),
    .Y(_955__bF$buf0)
);

BUFX2 BUFX2_insert23 (
    .A(_955_),
    .Y(_955__bF$buf1)
);

BUFX2 BUFX2_insert22 (
    .A(_955_),
    .Y(_955__bF$buf2)
);

BUFX2 BUFX2_insert21 (
    .A(_955_),
    .Y(_955__bF$buf3)
);

BUFX2 BUFX2_insert20 (
    .A(_955_),
    .Y(_955__bF$buf4)
);

BUFX2 BUFX2_insert19 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 )
);

BUFX2 BUFX2_insert18 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 )
);

BUFX2 BUFX2_insert17 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 )
);

BUFX2 BUFX2_insert16 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 )
);

BUFX2 BUFX2_insert15 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 )
);

BUFX2 BUFX2_insert14 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 )
);

BUFX2 BUFX2_insert13 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 )
);

BUFX2 BUFX2_insert12 (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 )
);

BUFX2 BUFX2_insert11 (
    .A(_1022_),
    .Y(_1022__bF$buf0)
);

BUFX2 BUFX2_insert10 (
    .A(_1022_),
    .Y(_1022__bF$buf1)
);

BUFX2 BUFX2_insert9 (
    .A(_1022_),
    .Y(_1022__bF$buf2)
);

BUFX2 BUFX2_insert8 (
    .A(_1022_),
    .Y(_1022__bF$buf3)
);

BUFX2 BUFX2_insert7 (
    .A(_1022_),
    .Y(_1022__bF$buf4)
);

BUFX2 BUFX2_insert6 (
    .A(_1022_),
    .Y(_1022__bF$buf5)
);

BUFX2 BUFX2_insert5 (
    .A(_1022_),
    .Y(_1022__bF$buf6)
);

BUFX2 BUFX2_insert4 (
    .A(_1063_),
    .Y(_1063__bF$buf0)
);

BUFX2 BUFX2_insert3 (
    .A(_1063_),
    .Y(_1063__bF$buf1)
);

BUFX2 BUFX2_insert2 (
    .A(_1063_),
    .Y(_1063__bF$buf2)
);

BUFX2 BUFX2_insert1 (
    .A(_1063_),
    .Y(_1063__bF$buf3)
);

BUFX2 BUFX2_insert0 (
    .A(_1063_),
    .Y(_1063__bF$buf4)
);

INVX1 _1780_ (
    .A(p_v_loc_fu_44[0]),
    .Y(_116_)
);

INVX1 _1781_ (
    .A(s_5_loc_fu_48[30]),
    .Y(_117_)
);

NOR2X1 _1782_ (
    .A(s_5_loc_fu_48[1]),
    .B(s_5_loc_fu_48[0]),
    .Y(_118_)
);

NOR2X1 _1783_ (
    .A(s_5_loc_fu_48[3]),
    .B(s_5_loc_fu_48[2]),
    .Y(_119_)
);

NOR2X1 _1784_ (
    .A(s_5_loc_fu_48[5]),
    .B(s_5_loc_fu_48[4]),
    .Y(_120_)
);

NAND3X1 _1785_ (
    .A(_118_),
    .B(_119_),
    .C(_120_),
    .Y(_121_)
);

INVX1 _1786_ (
    .A(s_5_loc_fu_48[11]),
    .Y(_122_)
);

INVX1 _1787_ (
    .A(s_5_loc_fu_48[10]),
    .Y(_123_)
);

NOR2X1 _1788_ (
    .A(s_5_loc_fu_48[13]),
    .B(s_5_loc_fu_48[12]),
    .Y(_124_)
);

NAND3X1 _1789_ (
    .A(_122_),
    .B(_123_),
    .C(_124_),
    .Y(_125_)
);

INVX1 _1790_ (
    .A(s_5_loc_fu_48[9]),
    .Y(_126_)
);

INVX1 _1791_ (
    .A(s_5_loc_fu_48[8]),
    .Y(_127_)
);

NOR2X1 _1792_ (
    .A(s_5_loc_fu_48[7]),
    .B(s_5_loc_fu_48[6]),
    .Y(_128_)
);

NAND3X1 _1793_ (
    .A(_126_),
    .B(_127_),
    .C(_128_),
    .Y(_129_)
);

NOR3X1 _1794_ (
    .A(_125_),
    .B(_129_),
    .C(_121_),
    .Y(_130_)
);

INVX1 _1795_ (
    .A(s_5_loc_fu_48[19]),
    .Y(_131_)
);

INVX1 _1796_ (
    .A(s_5_loc_fu_48[18]),
    .Y(_132_)
);

NOR2X1 _1797_ (
    .A(s_5_loc_fu_48[21]),
    .B(s_5_loc_fu_48[20]),
    .Y(_133_)
);

NAND3X1 _1798_ (
    .A(_131_),
    .B(_132_),
    .C(_133_),
    .Y(_134_)
);

INVX1 _1799_ (
    .A(s_5_loc_fu_48[17]),
    .Y(_135_)
);

INVX1 _1800_ (
    .A(s_5_loc_fu_48[16]),
    .Y(_136_)
);

NOR2X1 _1801_ (
    .A(s_5_loc_fu_48[15]),
    .B(s_5_loc_fu_48[14]),
    .Y(_137_)
);

NAND3X1 _1802_ (
    .A(_135_),
    .B(_136_),
    .C(_137_),
    .Y(_138_)
);

NOR2X1 _1803_ (
    .A(_134_),
    .B(_138_),
    .Y(_139_)
);

INVX1 _1804_ (
    .A(s_5_loc_fu_48[27]),
    .Y(_140_)
);

INVX1 _1805_ (
    .A(s_5_loc_fu_48[26]),
    .Y(_141_)
);

NOR2X1 _1806_ (
    .A(s_5_loc_fu_48[29]),
    .B(s_5_loc_fu_48[28]),
    .Y(_142_)
);

NAND3X1 _1807_ (
    .A(_140_),
    .B(_141_),
    .C(_142_),
    .Y(_143_)
);

INVX1 _1808_ (
    .A(s_5_loc_fu_48[23]),
    .Y(_144_)
);

INVX1 _1809_ (
    .A(s_5_loc_fu_48[22]),
    .Y(_145_)
);

NOR2X1 _1810_ (
    .A(s_5_loc_fu_48[25]),
    .B(s_5_loc_fu_48[24]),
    .Y(_146_)
);

NAND3X1 _1811_ (
    .A(_144_),
    .B(_145_),
    .C(_146_),
    .Y(_147_)
);

NOR2X1 _1812_ (
    .A(_143_),
    .B(_147_),
    .Y(_148_)
);

NAND3X1 _1813_ (
    .A(_139_),
    .B(_148_),
    .C(_130_),
    .Y(_149_)
);

NAND2X1 _1814_ (
    .A(_117_),
    .B(_149_),
    .Y(_150_)
);

INVX8 _1815_ (
    .A(_150_),
    .Y(_151_)
);

NAND2X1 _1816_ (
    .A(q_1_loc_fu_40[0]),
    .B(q_1_loc_fu_40[1]),
    .Y(_152_)
);

INVX1 _1817_ (
    .A(q_1_loc_fu_40[0]),
    .Y(_153_)
);

INVX1 _1818_ (
    .A(q_1_loc_fu_40[1]),
    .Y(_154_)
);

NAND2X1 _1819_ (
    .A(_153_),
    .B(_154_),
    .Y(_155_)
);

NAND3X1 _1820_ (
    .A(_152_),
    .B(_155_),
    .C(_151__bF$buf6),
    .Y(_156_)
);

OAI21X1 _1821_ (
    .A(_116_),
    .B(_151__bF$buf5),
    .C(_156_),
    .Y(_1779_[0])
);

INVX1 _1822_ (
    .A(p_v_loc_fu_44[1]),
    .Y(_157_)
);

INVX1 _1823_ (
    .A(q_1_loc_fu_40[2]),
    .Y(_158_)
);

AOI21X1 _1824_ (
    .A(q_1_loc_fu_40[0]),
    .B(q_1_loc_fu_40[1]),
    .C(_158_),
    .Y(_159_)
);

NOR2X1 _1825_ (
    .A(q_1_loc_fu_40[2]),
    .B(_152_),
    .Y(_160_)
);

OAI21X1 _1826_ (
    .A(_159_),
    .B(_160_),
    .C(_151__bF$buf4),
    .Y(_161_)
);

OAI21X1 _1827_ (
    .A(_157_),
    .B(_151__bF$buf3),
    .C(_161_),
    .Y(_1779_[1])
);

INVX1 _1828_ (
    .A(p_v_loc_fu_44[2]),
    .Y(_162_)
);

NAND2X1 _1829_ (
    .A(q_1_loc_fu_40[2]),
    .B(q_1_loc_fu_40[3]),
    .Y(_163_)
);

NOR2X1 _1830_ (
    .A(_152_),
    .B(_163_),
    .Y(_164_)
);

INVX2 _1831_ (
    .A(_164_),
    .Y(_165_)
);

INVX1 _1832_ (
    .A(q_1_loc_fu_40[3]),
    .Y(_166_)
);

OAI21X1 _1833_ (
    .A(_158_),
    .B(_152_),
    .C(_166_),
    .Y(_167_)
);

NAND3X1 _1834_ (
    .A(_165_),
    .B(_167_),
    .C(_151__bF$buf2),
    .Y(_168_)
);

OAI21X1 _1835_ (
    .A(_162_),
    .B(_151__bF$buf1),
    .C(_168_),
    .Y(_1779_[2])
);

INVX1 _1836_ (
    .A(p_v_loc_fu_44[3]),
    .Y(_169_)
);

INVX1 _1837_ (
    .A(q_1_loc_fu_40[4]),
    .Y(_170_)
);

NOR2X1 _1838_ (
    .A(_170_),
    .B(_164_),
    .Y(_171_)
);

NOR2X1 _1839_ (
    .A(q_1_loc_fu_40[4]),
    .B(_165_),
    .Y(_172_)
);

OAI21X1 _1840_ (
    .A(_171_),
    .B(_172_),
    .C(_151__bF$buf0),
    .Y(_173_)
);

OAI21X1 _1841_ (
    .A(_169_),
    .B(_151__bF$buf6),
    .C(_173_),
    .Y(_1779_[3])
);

INVX1 _1842_ (
    .A(p_v_loc_fu_44[4]),
    .Y(_174_)
);

NAND2X1 _1843_ (
    .A(q_1_loc_fu_40[4]),
    .B(q_1_loc_fu_40[5]),
    .Y(_175_)
);

NOR2X1 _1844_ (
    .A(_175_),
    .B(_165_),
    .Y(_176_)
);

INVX1 _1845_ (
    .A(_176_),
    .Y(_177_)
);

INVX1 _1846_ (
    .A(q_1_loc_fu_40[5]),
    .Y(_178_)
);

OAI21X1 _1847_ (
    .A(_170_),
    .B(_165_),
    .C(_178_),
    .Y(_179_)
);

NAND3X1 _1848_ (
    .A(_177_),
    .B(_179_),
    .C(_151__bF$buf5),
    .Y(_180_)
);

OAI21X1 _1849_ (
    .A(_174_),
    .B(_151__bF$buf4),
    .C(_180_),
    .Y(_1779_[4])
);

INVX1 _1850_ (
    .A(p_v_loc_fu_44[5]),
    .Y(_181_)
);

NAND2X1 _1851_ (
    .A(q_1_loc_fu_40[6]),
    .B(_176_),
    .Y(_182_)
);

INVX1 _1852_ (
    .A(q_1_loc_fu_40[6]),
    .Y(_183_)
);

OAI21X1 _1853_ (
    .A(_175_),
    .B(_165_),
    .C(_183_),
    .Y(_184_)
);

NAND3X1 _1854_ (
    .A(_182_),
    .B(_184_),
    .C(_151__bF$buf3),
    .Y(_185_)
);

OAI21X1 _1855_ (
    .A(_181_),
    .B(_151__bF$buf2),
    .C(_185_),
    .Y(_1779_[5])
);

INVX1 _1856_ (
    .A(p_v_loc_fu_44[6]),
    .Y(_186_)
);

INVX1 _1857_ (
    .A(q_1_loc_fu_40[7]),
    .Y(_187_)
);

AOI21X1 _1858_ (
    .A(_176_),
    .B(q_1_loc_fu_40[6]),
    .C(_187_),
    .Y(_188_)
);

NOR2X1 _1859_ (
    .A(q_1_loc_fu_40[7]),
    .B(_182_),
    .Y(_189_)
);

OAI21X1 _1860_ (
    .A(_188_),
    .B(_189_),
    .C(_151__bF$buf1),
    .Y(_190_)
);

OAI21X1 _1861_ (
    .A(_186_),
    .B(_151__bF$buf0),
    .C(_190_),
    .Y(_1779_[6])
);

INVX1 _1862_ (
    .A(p_v_loc_fu_44[7]),
    .Y(_191_)
);

INVX1 _1863_ (
    .A(q_1_loc_fu_40[8]),
    .Y(_192_)
);

NAND2X1 _1864_ (
    .A(q_1_loc_fu_40[6]),
    .B(q_1_loc_fu_40[7]),
    .Y(_193_)
);

NOR2X1 _1865_ (
    .A(_175_),
    .B(_193_),
    .Y(_194_)
);

AND2X2 _1866_ (
    .A(_164_),
    .B(_194_),
    .Y(_195_)
);

NOR2X1 _1867_ (
    .A(_192_),
    .B(_195_),
    .Y(_196_)
);

NAND2X1 _1868_ (
    .A(_164_),
    .B(_194_),
    .Y(_197_)
);

NOR2X1 _1869_ (
    .A(q_1_loc_fu_40[8]),
    .B(_197_),
    .Y(_198_)
);

OAI21X1 _1870_ (
    .A(_196_),
    .B(_198_),
    .C(_151__bF$buf6),
    .Y(_199_)
);

OAI21X1 _1871_ (
    .A(_191_),
    .B(_151__bF$buf5),
    .C(_199_),
    .Y(_1779_[7])
);

INVX1 _1872_ (
    .A(p_v_loc_fu_44[8]),
    .Y(_200_)
);

NAND2X1 _1873_ (
    .A(q_1_loc_fu_40[8]),
    .B(q_1_loc_fu_40[9]),
    .Y(_201_)
);

INVX1 _1874_ (
    .A(_201_),
    .Y(_202_)
);

NAND2X1 _1875_ (
    .A(_202_),
    .B(_195_),
    .Y(_203_)
);

INVX1 _1876_ (
    .A(q_1_loc_fu_40[9]),
    .Y(_204_)
);

OAI21X1 _1877_ (
    .A(_192_),
    .B(_197_),
    .C(_204_),
    .Y(_205_)
);

NAND3X1 _1878_ (
    .A(_203_),
    .B(_205_),
    .C(_151__bF$buf4),
    .Y(_206_)
);

OAI21X1 _1879_ (
    .A(_200_),
    .B(_151__bF$buf3),
    .C(_206_),
    .Y(_1779_[8])
);

INVX1 _1880_ (
    .A(p_v_loc_fu_44[9]),
    .Y(_207_)
);

INVX1 _1881_ (
    .A(q_1_loc_fu_40[10]),
    .Y(_208_)
);

AOI21X1 _1882_ (
    .A(_195_),
    .B(_202_),
    .C(_208_),
    .Y(_209_)
);

NOR2X1 _1883_ (
    .A(q_1_loc_fu_40[10]),
    .B(_203_),
    .Y(_210_)
);

OAI21X1 _1884_ (
    .A(_209_),
    .B(_210_),
    .C(_151__bF$buf2),
    .Y(_211_)
);

OAI21X1 _1885_ (
    .A(_207_),
    .B(_151__bF$buf1),
    .C(_211_),
    .Y(_1779_[9])
);

OAI21X1 _1886_ (
    .A(_208_),
    .B(_203_),
    .C(q_1_loc_fu_40[11]),
    .Y(_212_)
);

INVX1 _1887_ (
    .A(q_1_loc_fu_40[11]),
    .Y(_213_)
);

NOR2X1 _1888_ (
    .A(_208_),
    .B(_203_),
    .Y(_214_)
);

NAND2X1 _1889_ (
    .A(_213_),
    .B(_214_),
    .Y(_215_)
);

AND2X2 _1890_ (
    .A(_215_),
    .B(_212_),
    .Y(_216_)
);

NAND2X1 _1891_ (
    .A(p_v_loc_fu_44[10]),
    .B(_150_),
    .Y(_217_)
);

OAI21X1 _1892_ (
    .A(_150_),
    .B(_216_),
    .C(_217_),
    .Y(_1779_[10])
);

INVX1 _1893_ (
    .A(p_v_loc_fu_44[11]),
    .Y(_218_)
);

INVX1 _1894_ (
    .A(q_1_loc_fu_40[12]),
    .Y(_219_)
);

NAND2X1 _1895_ (
    .A(q_1_loc_fu_40[10]),
    .B(q_1_loc_fu_40[11]),
    .Y(_220_)
);

NOR2X1 _1896_ (
    .A(_201_),
    .B(_220_),
    .Y(_221_)
);

NAND2X1 _1897_ (
    .A(_221_),
    .B(_195_),
    .Y(_222_)
);

NAND2X1 _1898_ (
    .A(_219_),
    .B(_222_),
    .Y(_223_)
);

OR2X2 _1899_ (
    .A(_222_),
    .B(_219_),
    .Y(_224_)
);

NAND3X1 _1900_ (
    .A(_223_),
    .B(_224_),
    .C(_151__bF$buf0),
    .Y(_225_)
);

OAI21X1 _1901_ (
    .A(_218_),
    .B(_151__bF$buf6),
    .C(_225_),
    .Y(_1779_[11])
);

INVX1 _1902_ (
    .A(p_v_loc_fu_44[12]),
    .Y(_226_)
);

INVX1 _1903_ (
    .A(q_1_loc_fu_40[13]),
    .Y(_227_)
);

OAI21X1 _1904_ (
    .A(_219_),
    .B(_222_),
    .C(_227_),
    .Y(_228_)
);

INVX1 _1905_ (
    .A(_228_),
    .Y(_229_)
);

NAND2X1 _1906_ (
    .A(q_1_loc_fu_40[12]),
    .B(q_1_loc_fu_40[13]),
    .Y(_230_)
);

OAI21X1 _1907_ (
    .A(_222_),
    .B(_230_),
    .C(_151__bF$buf5),
    .Y(_231_)
);

OAI22X1 _1908_ (
    .A(_226_),
    .B(_151__bF$buf4),
    .C(_229_),
    .D(_231_),
    .Y(_1779_[12])
);

INVX1 _1909_ (
    .A(p_v_loc_fu_44[13]),
    .Y(_232_)
);

INVX1 _1910_ (
    .A(q_1_loc_fu_40[14]),
    .Y(_233_)
);

OAI21X1 _1911_ (
    .A(_230_),
    .B(_222_),
    .C(_233_),
    .Y(_234_)
);

INVX1 _1912_ (
    .A(_230_),
    .Y(_235_)
);

NAND3X1 _1913_ (
    .A(_221_),
    .B(_235_),
    .C(_195_),
    .Y(_236_)
);

NOR2X1 _1914_ (
    .A(_233_),
    .B(_236_),
    .Y(_237_)
);

INVX1 _1915_ (
    .A(_237_),
    .Y(_238_)
);

NAND3X1 _1916_ (
    .A(_234_),
    .B(_238_),
    .C(_151__bF$buf3),
    .Y(_239_)
);

OAI21X1 _1917_ (
    .A(_232_),
    .B(_151__bF$buf2),
    .C(_239_),
    .Y(_1779_[13])
);

INVX1 _1918_ (
    .A(q_1_loc_fu_40[15]),
    .Y(_240_)
);

NOR2X1 _1919_ (
    .A(_240_),
    .B(_237_),
    .Y(_241_)
);

AND2X2 _1920_ (
    .A(_237_),
    .B(_240_),
    .Y(_242_)
);

OAI21X1 _1921_ (
    .A(_241_),
    .B(_242_),
    .C(_151__bF$buf1),
    .Y(_243_)
);

NAND2X1 _1922_ (
    .A(p_v_loc_fu_44[14]),
    .B(_150_),
    .Y(_244_)
);

NAND2X1 _1923_ (
    .A(_244_),
    .B(_243_),
    .Y(_1779_[14])
);

INVX1 _1924_ (
    .A(p_v_loc_fu_44[15]),
    .Y(_245_)
);

INVX1 _1925_ (
    .A(q_1_loc_fu_40[16]),
    .Y(_246_)
);

NAND2X1 _1926_ (
    .A(q_1_loc_fu_40[14]),
    .B(q_1_loc_fu_40[15]),
    .Y(_247_)
);

NOR2X1 _1927_ (
    .A(_230_),
    .B(_247_),
    .Y(_248_)
);

NAND2X1 _1928_ (
    .A(_221_),
    .B(_248_),
    .Y(_249_)
);

NOR2X1 _1929_ (
    .A(_197_),
    .B(_249_),
    .Y(_250_)
);

NOR2X1 _1930_ (
    .A(_246_),
    .B(_250_),
    .Y(_251_)
);

AND2X2 _1931_ (
    .A(_221_),
    .B(_248_),
    .Y(_252_)
);

NAND2X1 _1932_ (
    .A(_195_),
    .B(_252_),
    .Y(_253_)
);

NOR2X1 _1933_ (
    .A(q_1_loc_fu_40[16]),
    .B(_253_),
    .Y(_254_)
);

OAI21X1 _1934_ (
    .A(_251_),
    .B(_254_),
    .C(_151__bF$buf0),
    .Y(_255_)
);

OAI21X1 _1935_ (
    .A(_245_),
    .B(_151__bF$buf6),
    .C(_255_),
    .Y(_1779_[15])
);

INVX1 _1936_ (
    .A(p_v_loc_fu_44[16]),
    .Y(_256_)
);

AOI21X1 _1937_ (
    .A(_250_),
    .B(q_1_loc_fu_40[16]),
    .C(q_1_loc_fu_40[17]),
    .Y(_257_)
);

NAND2X1 _1938_ (
    .A(q_1_loc_fu_40[16]),
    .B(q_1_loc_fu_40[17]),
    .Y(_258_)
);

OAI21X1 _1939_ (
    .A(_253_),
    .B(_258_),
    .C(_151__bF$buf5),
    .Y(_259_)
);

OAI22X1 _1940_ (
    .A(_256_),
    .B(_151__bF$buf4),
    .C(_257_),
    .D(_259_),
    .Y(_1779_[16])
);

INVX1 _1941_ (
    .A(p_v_loc_fu_44[17]),
    .Y(_260_)
);

INVX1 _1942_ (
    .A(q_1_loc_fu_40[18]),
    .Y(_261_)
);

OAI21X1 _1943_ (
    .A(_258_),
    .B(_253_),
    .C(_261_),
    .Y(_262_)
);

NOR2X1 _1944_ (
    .A(_258_),
    .B(_253_),
    .Y(_263_)
);

NAND2X1 _1945_ (
    .A(q_1_loc_fu_40[18]),
    .B(_263_),
    .Y(_264_)
);

NAND3X1 _1946_ (
    .A(_262_),
    .B(_264_),
    .C(_151__bF$buf3),
    .Y(_265_)
);

OAI21X1 _1947_ (
    .A(_260_),
    .B(_151__bF$buf2),
    .C(_265_),
    .Y(_1779_[17])
);

INVX1 _1948_ (
    .A(p_v_loc_fu_44[18]),
    .Y(_266_)
);

INVX1 _1949_ (
    .A(q_1_loc_fu_40[19]),
    .Y(_267_)
);

AOI21X1 _1950_ (
    .A(_263_),
    .B(q_1_loc_fu_40[18]),
    .C(_267_),
    .Y(_268_)
);

INVX1 _1951_ (
    .A(_258_),
    .Y(_269_)
);

NAND2X1 _1952_ (
    .A(_269_),
    .B(_250_),
    .Y(_270_)
);

NOR3X1 _1953_ (
    .A(_261_),
    .B(q_1_loc_fu_40[19]),
    .C(_270_),
    .Y(_271_)
);

OAI21X1 _1954_ (
    .A(_268_),
    .B(_271_),
    .C(_151__bF$buf1),
    .Y(_272_)
);

OAI21X1 _1955_ (
    .A(_266_),
    .B(_151__bF$buf0),
    .C(_272_),
    .Y(_1779_[18])
);

INVX1 _1956_ (
    .A(p_v_loc_fu_44[19]),
    .Y(_273_)
);

NAND2X1 _1957_ (
    .A(q_1_loc_fu_40[18]),
    .B(q_1_loc_fu_40[19]),
    .Y(_274_)
);

NOR2X1 _1958_ (
    .A(_258_),
    .B(_274_),
    .Y(_275_)
);

NAND3X1 _1959_ (
    .A(_275_),
    .B(_195_),
    .C(_252_),
    .Y(_276_)
);

INVX1 _1960_ (
    .A(_276_),
    .Y(_277_)
);

NAND2X1 _1961_ (
    .A(q_1_loc_fu_40[20]),
    .B(_277_),
    .Y(_278_)
);

INVX1 _1962_ (
    .A(q_1_loc_fu_40[20]),
    .Y(_279_)
);

NAND2X1 _1963_ (
    .A(_279_),
    .B(_276_),
    .Y(_280_)
);

NAND3X1 _1964_ (
    .A(_280_),
    .B(_151__bF$buf6),
    .C(_278_),
    .Y(_281_)
);

OAI21X1 _1965_ (
    .A(_273_),
    .B(_151__bF$buf5),
    .C(_281_),
    .Y(_1779_[19])
);

INVX1 _1966_ (
    .A(p_v_loc_fu_44[20]),
    .Y(_282_)
);

INVX1 _1967_ (
    .A(q_1_loc_fu_40[21]),
    .Y(_283_)
);

AOI21X1 _1968_ (
    .A(_277_),
    .B(q_1_loc_fu_40[20]),
    .C(_283_),
    .Y(_284_)
);

NOR3X1 _1969_ (
    .A(_279_),
    .B(q_1_loc_fu_40[21]),
    .C(_276_),
    .Y(_285_)
);

OAI21X1 _1970_ (
    .A(_285_),
    .B(_284_),
    .C(_151__bF$buf4),
    .Y(_286_)
);

OAI21X1 _1971_ (
    .A(_282_),
    .B(_151__bF$buf3),
    .C(_286_),
    .Y(_1779_[20])
);

NAND2X1 _1972_ (
    .A(q_1_loc_fu_40[20]),
    .B(q_1_loc_fu_40[21]),
    .Y(_287_)
);

NOR2X1 _1973_ (
    .A(_287_),
    .B(_276_),
    .Y(_288_)
);

NAND2X1 _1974_ (
    .A(q_1_loc_fu_40[22]),
    .B(_288_),
    .Y(_289_)
);

INVX1 _1975_ (
    .A(q_1_loc_fu_40[22]),
    .Y(_290_)
);

OAI21X1 _1976_ (
    .A(_287_),
    .B(_276_),
    .C(_290_),
    .Y(_291_)
);

NAND2X1 _1977_ (
    .A(_291_),
    .B(_289_),
    .Y(_292_)
);

NAND2X1 _1978_ (
    .A(p_v_loc_fu_44[21]),
    .B(_150_),
    .Y(_293_)
);

OAI21X1 _1979_ (
    .A(_150_),
    .B(_292_),
    .C(_293_),
    .Y(_1779_[21])
);

INVX1 _1980_ (
    .A(q_1_loc_fu_40[23]),
    .Y(_294_)
);

AOI21X1 _1981_ (
    .A(_288_),
    .B(q_1_loc_fu_40[22]),
    .C(_294_),
    .Y(_295_)
);

INVX1 _1982_ (
    .A(_287_),
    .Y(_296_)
);

NAND3X1 _1983_ (
    .A(_275_),
    .B(_296_),
    .C(_250_),
    .Y(_297_)
);

NOR3X1 _1984_ (
    .A(_290_),
    .B(q_1_loc_fu_40[23]),
    .C(_297_),
    .Y(_298_)
);

OAI21X1 _1985_ (
    .A(_298_),
    .B(_295_),
    .C(_151__bF$buf2),
    .Y(_299_)
);

NAND2X1 _1986_ (
    .A(p_v_loc_fu_44[22]),
    .B(_150_),
    .Y(_300_)
);

NAND2X1 _1987_ (
    .A(_300_),
    .B(_299_),
    .Y(_1779_[22])
);

INVX1 _1988_ (
    .A(p_v_loc_fu_44[23]),
    .Y(_301_)
);

NAND2X1 _1989_ (
    .A(q_1_loc_fu_40[22]),
    .B(q_1_loc_fu_40[23]),
    .Y(_302_)
);

NOR2X1 _1990_ (
    .A(_287_),
    .B(_302_),
    .Y(_303_)
);

NAND2X1 _1991_ (
    .A(_275_),
    .B(_303_),
    .Y(_304_)
);

NOR2X1 _1992_ (
    .A(_304_),
    .B(_253_),
    .Y(_305_)
);

NAND2X1 _1993_ (
    .A(q_1_loc_fu_40[24]),
    .B(_305_),
    .Y(_306_)
);

INVX1 _1994_ (
    .A(q_1_loc_fu_40[24]),
    .Y(_307_)
);

OAI21X1 _1995_ (
    .A(_304_),
    .B(_253_),
    .C(_307_),
    .Y(_308_)
);

NAND3X1 _1996_ (
    .A(_308_),
    .B(_306_),
    .C(_151__bF$buf1),
    .Y(_309_)
);

OAI21X1 _1997_ (
    .A(_301_),
    .B(_151__bF$buf0),
    .C(_309_),
    .Y(_1779_[23])
);

INVX1 _1998_ (
    .A(p_v_loc_fu_44[24]),
    .Y(_310_)
);

INVX1 _1999_ (
    .A(q_1_loc_fu_40[25]),
    .Y(_311_)
);

AOI21X1 _2000_ (
    .A(_305_),
    .B(q_1_loc_fu_40[24]),
    .C(_311_),
    .Y(_312_)
);

INVX1 _2001_ (
    .A(_304_),
    .Y(_313_)
);

NAND2X1 _2002_ (
    .A(_313_),
    .B(_250_),
    .Y(_314_)
);

NOR3X1 _2003_ (
    .A(_307_),
    .B(q_1_loc_fu_40[25]),
    .C(_314_),
    .Y(_315_)
);

OAI21X1 _2004_ (
    .A(_312_),
    .B(_315_),
    .C(_151__bF$buf6),
    .Y(_316_)
);

OAI21X1 _2005_ (
    .A(_310_),
    .B(_151__bF$buf5),
    .C(_316_),
    .Y(_1779_[24])
);

INVX1 _2006_ (
    .A(p_v_loc_fu_44[25]),
    .Y(_317_)
);

NAND2X1 _2007_ (
    .A(q_1_loc_fu_40[24]),
    .B(q_1_loc_fu_40[25]),
    .Y(_318_)
);

INVX1 _2008_ (
    .A(_318_),
    .Y(_319_)
);

NAND3X1 _2009_ (
    .A(q_1_loc_fu_40[26]),
    .B(_319_),
    .C(_305_),
    .Y(_320_)
);

INVX1 _2010_ (
    .A(q_1_loc_fu_40[26]),
    .Y(_321_)
);

OAI21X1 _2011_ (
    .A(_318_),
    .B(_314_),
    .C(_321_),
    .Y(_322_)
);

NAND3X1 _2012_ (
    .A(_322_),
    .B(_151__bF$buf4),
    .C(_320_),
    .Y(_323_)
);

OAI21X1 _2013_ (
    .A(_317_),
    .B(_151__bF$buf3),
    .C(_323_),
    .Y(_1779_[25])
);

INVX1 _2014_ (
    .A(p_v_loc_fu_44[26]),
    .Y(_324_)
);

NOR2X1 _2015_ (
    .A(_318_),
    .B(_314_),
    .Y(_325_)
);

AOI21X1 _2016_ (
    .A(_325_),
    .B(q_1_loc_fu_40[26]),
    .C(q_1_loc_fu_40[27]),
    .Y(_326_)
);

INVX1 _2017_ (
    .A(q_1_loc_fu_40[27]),
    .Y(_327_)
);

OAI21X1 _2018_ (
    .A(_327_),
    .B(_320_),
    .C(_151__bF$buf2),
    .Y(_328_)
);

OAI22X1 _2019_ (
    .A(_324_),
    .B(_151__bF$buf1),
    .C(_326_),
    .D(_328_),
    .Y(_1779_[26])
);

INVX1 _2020_ (
    .A(p_v_loc_fu_44[27]),
    .Y(_329_)
);

INVX1 _2021_ (
    .A(q_1_loc_fu_40[28]),
    .Y(_330_)
);

NAND2X1 _2022_ (
    .A(q_1_loc_fu_40[26]),
    .B(q_1_loc_fu_40[27]),
    .Y(_331_)
);

NOR2X1 _2023_ (
    .A(_318_),
    .B(_331_),
    .Y(_332_)
);

AOI21X1 _2024_ (
    .A(_305_),
    .B(_332_),
    .C(_330_),
    .Y(_333_)
);

INVX1 _2025_ (
    .A(_332_),
    .Y(_334_)
);

NOR3X1 _2026_ (
    .A(q_1_loc_fu_40[28]),
    .B(_334_),
    .C(_314_),
    .Y(_335_)
);

OAI21X1 _2027_ (
    .A(_333_),
    .B(_335_),
    .C(_151__bF$buf0),
    .Y(_336_)
);

OAI21X1 _2028_ (
    .A(_329_),
    .B(_151__bF$buf6),
    .C(_336_),
    .Y(_1779_[27])
);

INVX1 _2029_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .Y(_337_)
);

NOR2X1 _2030_ (
    .A(ap_start),
    .B(_337_),
    .Y(_1778_)
);

INVX1 _2031_ (
    .A(s_5_loc_fu_48[0]),
    .Y(_338_)
);

AND2X2 _2032_ (
    .A(ap_CS_fsm_state2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0 ),
    .Y(_339_)
);

NAND2X1 _2033_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_1_fu_177_p2 [0]),
    .B(_339__bF$buf6),
    .Y(_340_)
);

OAI21X1 _2034_ (
    .A(_338_),
    .B(_339__bF$buf5),
    .C(_340_),
    .Y(_3_)
);

INVX1 _2035_ (
    .A(s_5_loc_fu_48[1]),
    .Y(_341_)
);

NAND2X1 _2036_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [1]),
    .B(_339__bF$buf4),
    .Y(_342_)
);

OAI21X1 _2037_ (
    .A(_341_),
    .B(_339__bF$buf3),
    .C(_342_),
    .Y(_4_)
);

INVX1 _2038_ (
    .A(s_5_loc_fu_48[2]),
    .Y(_343_)
);

NAND2X1 _2039_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [2]),
    .B(_339__bF$buf2),
    .Y(_344_)
);

OAI21X1 _2040_ (
    .A(_343_),
    .B(_339__bF$buf1),
    .C(_344_),
    .Y(_5_)
);

INVX1 _2041_ (
    .A(s_5_loc_fu_48[3]),
    .Y(_345_)
);

NAND2X1 _2042_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [3]),
    .B(_339__bF$buf0),
    .Y(_346_)
);

OAI21X1 _2043_ (
    .A(_345_),
    .B(_339__bF$buf6),
    .C(_346_),
    .Y(_6_)
);

INVX1 _2044_ (
    .A(s_5_loc_fu_48[4]),
    .Y(_347_)
);

NAND2X1 _2045_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [4]),
    .B(_339__bF$buf5),
    .Y(_348_)
);

OAI21X1 _2046_ (
    .A(_347_),
    .B(_339__bF$buf4),
    .C(_348_),
    .Y(_7_)
);

INVX1 _2047_ (
    .A(s_5_loc_fu_48[5]),
    .Y(_349_)
);

NAND2X1 _2048_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [5]),
    .B(_339__bF$buf3),
    .Y(_350_)
);

OAI21X1 _2049_ (
    .A(_349_),
    .B(_339__bF$buf2),
    .C(_350_),
    .Y(_8_)
);

INVX1 _2050_ (
    .A(s_5_loc_fu_48[6]),
    .Y(_351_)
);

NAND2X1 _2051_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [6]),
    .B(_339__bF$buf1),
    .Y(_352_)
);

OAI21X1 _2052_ (
    .A(_351_),
    .B(_339__bF$buf0),
    .C(_352_),
    .Y(_9_)
);

INVX1 _2053_ (
    .A(s_5_loc_fu_48[7]),
    .Y(_353_)
);

NAND2X1 _2054_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [7]),
    .B(_339__bF$buf6),
    .Y(_354_)
);

OAI21X1 _2055_ (
    .A(_353_),
    .B(_339__bF$buf5),
    .C(_354_),
    .Y(_10_)
);

NAND2X1 _2056_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [8]),
    .B(_339__bF$buf4),
    .Y(_355_)
);

OAI21X1 _2057_ (
    .A(_127_),
    .B(_339__bF$buf3),
    .C(_355_),
    .Y(_11_)
);

NAND2X1 _2058_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [9]),
    .B(_339__bF$buf2),
    .Y(_356_)
);

OAI21X1 _2059_ (
    .A(_126_),
    .B(_339__bF$buf1),
    .C(_356_),
    .Y(_12_)
);

NAND2X1 _2060_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [10]),
    .B(_339__bF$buf0),
    .Y(_357_)
);

OAI21X1 _2061_ (
    .A(_123_),
    .B(_339__bF$buf6),
    .C(_357_),
    .Y(_13_)
);

NAND2X1 _2062_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [11]),
    .B(_339__bF$buf5),
    .Y(_358_)
);

OAI21X1 _2063_ (
    .A(_122_),
    .B(_339__bF$buf4),
    .C(_358_),
    .Y(_14_)
);

INVX1 _2064_ (
    .A(s_5_loc_fu_48[12]),
    .Y(_359_)
);

NAND2X1 _2065_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [12]),
    .B(_339__bF$buf3),
    .Y(_360_)
);

OAI21X1 _2066_ (
    .A(_359_),
    .B(_339__bF$buf2),
    .C(_360_),
    .Y(_15_)
);

INVX1 _2067_ (
    .A(s_5_loc_fu_48[13]),
    .Y(_361_)
);

NAND2X1 _2068_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [13]),
    .B(_339__bF$buf1),
    .Y(_362_)
);

OAI21X1 _2069_ (
    .A(_361_),
    .B(_339__bF$buf0),
    .C(_362_),
    .Y(_16_)
);

INVX1 _2070_ (
    .A(s_5_loc_fu_48[14]),
    .Y(_363_)
);

NAND2X1 _2071_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [14]),
    .B(_339__bF$buf6),
    .Y(_364_)
);

OAI21X1 _2072_ (
    .A(_363_),
    .B(_339__bF$buf5),
    .C(_364_),
    .Y(_17_)
);

INVX1 _2073_ (
    .A(s_5_loc_fu_48[15]),
    .Y(_365_)
);

NAND2X1 _2074_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [15]),
    .B(_339__bF$buf4),
    .Y(_366_)
);

OAI21X1 _2075_ (
    .A(_365_),
    .B(_339__bF$buf3),
    .C(_366_),
    .Y(_18_)
);

NAND2X1 _2076_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [16]),
    .B(_339__bF$buf2),
    .Y(_367_)
);

OAI21X1 _2077_ (
    .A(_136_),
    .B(_339__bF$buf1),
    .C(_367_),
    .Y(_19_)
);

NAND2X1 _2078_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [17]),
    .B(_339__bF$buf0),
    .Y(_368_)
);

OAI21X1 _2079_ (
    .A(_135_),
    .B(_339__bF$buf6),
    .C(_368_),
    .Y(_20_)
);

NAND2X1 _2080_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [18]),
    .B(_339__bF$buf5),
    .Y(_369_)
);

OAI21X1 _2081_ (
    .A(_132_),
    .B(_339__bF$buf4),
    .C(_369_),
    .Y(_21_)
);

NAND2X1 _2082_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [19]),
    .B(_339__bF$buf3),
    .Y(_370_)
);

OAI21X1 _2083_ (
    .A(_131_),
    .B(_339__bF$buf2),
    .C(_370_),
    .Y(_22_)
);

INVX1 _2084_ (
    .A(s_5_loc_fu_48[20]),
    .Y(_371_)
);

NAND2X1 _2085_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [20]),
    .B(_339__bF$buf1),
    .Y(_372_)
);

OAI21X1 _2086_ (
    .A(_371_),
    .B(_339__bF$buf0),
    .C(_372_),
    .Y(_23_)
);

INVX1 _2087_ (
    .A(s_5_loc_fu_48[21]),
    .Y(_373_)
);

NAND2X1 _2088_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [21]),
    .B(_339__bF$buf6),
    .Y(_374_)
);

OAI21X1 _2089_ (
    .A(_373_),
    .B(_339__bF$buf5),
    .C(_374_),
    .Y(_24_)
);

NAND2X1 _2090_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [22]),
    .B(_339__bF$buf4),
    .Y(_375_)
);

OAI21X1 _2091_ (
    .A(_145_),
    .B(_339__bF$buf3),
    .C(_375_),
    .Y(_25_)
);

NAND2X1 _2092_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [23]),
    .B(_339__bF$buf2),
    .Y(_376_)
);

OAI21X1 _2093_ (
    .A(_144_),
    .B(_339__bF$buf1),
    .C(_376_),
    .Y(_26_)
);

INVX1 _2094_ (
    .A(s_5_loc_fu_48[24]),
    .Y(_377_)
);

NAND2X1 _2095_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [24]),
    .B(_339__bF$buf0),
    .Y(_378_)
);

OAI21X1 _2096_ (
    .A(_377_),
    .B(_339__bF$buf6),
    .C(_378_),
    .Y(_27_)
);

INVX1 _2097_ (
    .A(s_5_loc_fu_48[25]),
    .Y(_379_)
);

NAND2X1 _2098_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [25]),
    .B(_339__bF$buf5),
    .Y(_380_)
);

OAI21X1 _2099_ (
    .A(_379_),
    .B(_339__bF$buf4),
    .C(_380_),
    .Y(_28_)
);

NAND2X1 _2100_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [26]),
    .B(_339__bF$buf3),
    .Y(_381_)
);

OAI21X1 _2101_ (
    .A(_141_),
    .B(_339__bF$buf2),
    .C(_381_),
    .Y(_29_)
);

NAND2X1 _2102_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [27]),
    .B(_339__bF$buf1),
    .Y(_382_)
);

OAI21X1 _2103_ (
    .A(_140_),
    .B(_339__bF$buf0),
    .C(_382_),
    .Y(_30_)
);

INVX1 _2104_ (
    .A(s_5_loc_fu_48[28]),
    .Y(_383_)
);

NAND2X1 _2105_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [28]),
    .B(_339__bF$buf6),
    .Y(_384_)
);

OAI21X1 _2106_ (
    .A(_383_),
    .B(_339__bF$buf5),
    .C(_384_),
    .Y(_31_)
);

INVX1 _2107_ (
    .A(s_5_loc_fu_48[29]),
    .Y(_385_)
);

NAND2X1 _2108_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [29]),
    .B(_339__bF$buf4),
    .Y(_386_)
);

OAI21X1 _2109_ (
    .A(_385_),
    .B(_339__bF$buf3),
    .C(_386_),
    .Y(_32_)
);

NAND2X1 _2110_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [30]),
    .B(_339__bF$buf2),
    .Y(_387_)
);

OAI21X1 _2111_ (
    .A(_117_),
    .B(_339__bF$buf1),
    .C(_387_),
    .Y(_33_)
);

INVX1 _2112_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [4]),
    .Y(_388_)
);

NAND2X1 _2113_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(in_val[0]),
    .Y(_389_)
);

OAI21X1 _2114_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(_388_),
    .C(_389_),
    .Y(_34_)
);

INVX1 _2115_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [5]),
    .Y(_390_)
);

NAND2X1 _2116_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(in_val[1]),
    .Y(_391_)
);

OAI21X1 _2117_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(_390_),
    .C(_391_),
    .Y(_35_)
);

INVX1 _2118_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [6]),
    .Y(_392_)
);

NAND2X1 _2119_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(in_val[2]),
    .Y(_393_)
);

OAI21X1 _2120_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(_392_),
    .C(_393_),
    .Y(_36_)
);

INVX1 _2121_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [7]),
    .Y(_394_)
);

NAND2X1 _2122_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .B(in_val[3]),
    .Y(_395_)
);

OAI21X1 _2123_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(_394_),
    .C(_395_),
    .Y(_37_)
);

INVX1 _2124_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [8]),
    .Y(_396_)
);

NAND2X1 _2125_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(in_val[4]),
    .Y(_397_)
);

OAI21X1 _2126_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(_396_),
    .C(_397_),
    .Y(_38_)
);

INVX1 _2127_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [9]),
    .Y(_398_)
);

NAND2X1 _2128_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(in_val[5]),
    .Y(_399_)
);

OAI21X1 _2129_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(_398_),
    .C(_399_),
    .Y(_39_)
);

INVX1 _2130_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [10]),
    .Y(_400_)
);

NAND2X1 _2131_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(in_val[6]),
    .Y(_401_)
);

OAI21X1 _2132_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .B(_400_),
    .C(_401_),
    .Y(_40_)
);

INVX1 _2133_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [11]),
    .Y(_402_)
);

NAND2X1 _2134_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(in_val[7]),
    .Y(_403_)
);

OAI21X1 _2135_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(_402_),
    .C(_403_),
    .Y(_41_)
);

INVX1 _2136_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [12]),
    .Y(_404_)
);

NAND2X1 _2137_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(in_val[8]),
    .Y(_405_)
);

OAI21X1 _2138_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(_404_),
    .C(_405_),
    .Y(_42_)
);

INVX1 _2139_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [13]),
    .Y(_406_)
);

NAND2X1 _2140_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(in_val[9]),
    .Y(_407_)
);

OAI21X1 _2141_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(_406_),
    .C(_407_),
    .Y(_43_)
);

INVX1 _2142_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [14]),
    .Y(_408_)
);

NAND2X1 _2143_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .B(in_val[10]),
    .Y(_409_)
);

OAI21X1 _2144_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(_408_),
    .C(_409_),
    .Y(_44_)
);

INVX1 _2145_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [15]),
    .Y(_410_)
);

NAND2X1 _2146_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(in_val[11]),
    .Y(_411_)
);

OAI21X1 _2147_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(_410_),
    .C(_411_),
    .Y(_45_)
);

INVX1 _2148_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [16]),
    .Y(_412_)
);

NAND2X1 _2149_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(in_val[12]),
    .Y(_413_)
);

OAI21X1 _2150_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(_412_),
    .C(_413_),
    .Y(_46_)
);

INVX1 _2151_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [17]),
    .Y(_414_)
);

NAND2X1 _2152_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(in_val[13]),
    .Y(_415_)
);

OAI21X1 _2153_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .B(_414_),
    .C(_415_),
    .Y(_47_)
);

INVX1 _2154_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [18]),
    .Y(_416_)
);

NAND2X1 _2155_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(in_val[14]),
    .Y(_417_)
);

OAI21X1 _2156_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(_416_),
    .C(_417_),
    .Y(_48_)
);

INVX1 _2157_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [19]),
    .Y(_418_)
);

NAND2X1 _2158_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(in_val[15]),
    .Y(_419_)
);

OAI21X1 _2159_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(_418_),
    .C(_419_),
    .Y(_49_)
);

INVX1 _2160_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [20]),
    .Y(_420_)
);

NAND2X1 _2161_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(in_val[16]),
    .Y(_421_)
);

OAI21X1 _2162_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(_420_),
    .C(_421_),
    .Y(_50_)
);

INVX1 _2163_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [21]),
    .Y(_422_)
);

NAND2X1 _2164_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .B(in_val[17]),
    .Y(_423_)
);

OAI21X1 _2165_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(_422_),
    .C(_423_),
    .Y(_51_)
);

INVX1 _2166_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [22]),
    .Y(_424_)
);

NAND2X1 _2167_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(in_val[18]),
    .Y(_425_)
);

OAI21X1 _2168_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(_424_),
    .C(_425_),
    .Y(_52_)
);

INVX1 _2169_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [23]),
    .Y(_426_)
);

NAND2X1 _2170_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(in_val[19]),
    .Y(_427_)
);

OAI21X1 _2171_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(_426_),
    .C(_427_),
    .Y(_53_)
);

INVX1 _2172_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [24]),
    .Y(_428_)
);

NAND2X1 _2173_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(in_val[20]),
    .Y(_429_)
);

OAI21X1 _2174_ (
    .A(ap_CS_fsm_state1_bF$buf6),
    .B(_428_),
    .C(_429_),
    .Y(_54_)
);

INVX1 _2175_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [25]),
    .Y(_430_)
);

NAND2X1 _2176_ (
    .A(ap_CS_fsm_state1_bF$buf5),
    .B(in_val[21]),
    .Y(_431_)
);

OAI21X1 _2177_ (
    .A(ap_CS_fsm_state1_bF$buf4),
    .B(_430_),
    .C(_431_),
    .Y(_55_)
);

INVX1 _2178_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [26]),
    .Y(_432_)
);

NAND2X1 _2179_ (
    .A(ap_CS_fsm_state1_bF$buf3),
    .B(in_val[22]),
    .Y(_433_)
);

OAI21X1 _2180_ (
    .A(ap_CS_fsm_state1_bF$buf2),
    .B(_432_),
    .C(_433_),
    .Y(_56_)
);

INVX1 _2181_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [27]),
    .Y(_434_)
);

NAND2X1 _2182_ (
    .A(ap_CS_fsm_state1_bF$buf1),
    .B(in_val[23]),
    .Y(_435_)
);

OAI21X1 _2183_ (
    .A(ap_CS_fsm_state1_bF$buf0),
    .B(_434_),
    .C(_435_),
    .Y(_57_)
);

AND2X2 _2184_ (
    .A(ap_CS_fsm_state2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0 ),
    .Y(_436_)
);

NAND2X1 _2185_ (
    .A(vdd),
    .B(_436__bF$buf6),
    .Y(_437_)
);

OAI21X1 _2186_ (
    .A(_153_),
    .B(_436__bF$buf5),
    .C(_437_),
    .Y(_58_)
);

NAND2X1 _2187_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [0]),
    .B(_436__bF$buf4),
    .Y(_438_)
);

OAI21X1 _2188_ (
    .A(_154_),
    .B(_436__bF$buf3),
    .C(_438_),
    .Y(_59_)
);

NAND2X1 _2189_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [1]),
    .B(_436__bF$buf2),
    .Y(_439_)
);

OAI21X1 _2190_ (
    .A(_158_),
    .B(_436__bF$buf1),
    .C(_439_),
    .Y(_60_)
);

NAND2X1 _2191_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [2]),
    .B(_436__bF$buf0),
    .Y(_440_)
);

OAI21X1 _2192_ (
    .A(_166_),
    .B(_436__bF$buf6),
    .C(_440_),
    .Y(_61_)
);

NAND2X1 _2193_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [3]),
    .B(_436__bF$buf5),
    .Y(_441_)
);

OAI21X1 _2194_ (
    .A(_170_),
    .B(_436__bF$buf4),
    .C(_441_),
    .Y(_62_)
);

NAND2X1 _2195_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [4]),
    .B(_436__bF$buf3),
    .Y(_442_)
);

OAI21X1 _2196_ (
    .A(_178_),
    .B(_436__bF$buf2),
    .C(_442_),
    .Y(_63_)
);

NAND2X1 _2197_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [5]),
    .B(_436__bF$buf1),
    .Y(_443_)
);

OAI21X1 _2198_ (
    .A(_183_),
    .B(_436__bF$buf0),
    .C(_443_),
    .Y(_64_)
);

NAND2X1 _2199_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [6]),
    .B(_436__bF$buf6),
    .Y(_444_)
);

OAI21X1 _2200_ (
    .A(_187_),
    .B(_436__bF$buf5),
    .C(_444_),
    .Y(_65_)
);

NAND2X1 _2201_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [7]),
    .B(_436__bF$buf4),
    .Y(_445_)
);

OAI21X1 _2202_ (
    .A(_192_),
    .B(_436__bF$buf3),
    .C(_445_),
    .Y(_66_)
);

NAND2X1 _2203_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [8]),
    .B(_436__bF$buf2),
    .Y(_446_)
);

OAI21X1 _2204_ (
    .A(_204_),
    .B(_436__bF$buf1),
    .C(_446_),
    .Y(_67_)
);

NAND2X1 _2205_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [9]),
    .B(_436__bF$buf0),
    .Y(_447_)
);

OAI21X1 _2206_ (
    .A(_208_),
    .B(_436__bF$buf6),
    .C(_447_),
    .Y(_68_)
);

NAND2X1 _2207_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [10]),
    .B(_436__bF$buf5),
    .Y(_448_)
);

OAI21X1 _2208_ (
    .A(_213_),
    .B(_436__bF$buf4),
    .C(_448_),
    .Y(_69_)
);

NAND2X1 _2209_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [11]),
    .B(_436__bF$buf3),
    .Y(_449_)
);

OAI21X1 _2210_ (
    .A(_219_),
    .B(_436__bF$buf2),
    .C(_449_),
    .Y(_70_)
);

NAND2X1 _2211_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [12]),
    .B(_436__bF$buf1),
    .Y(_450_)
);

OAI21X1 _2212_ (
    .A(_227_),
    .B(_436__bF$buf0),
    .C(_450_),
    .Y(_71_)
);

NAND2X1 _2213_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [13]),
    .B(_436__bF$buf6),
    .Y(_451_)
);

OAI21X1 _2214_ (
    .A(_233_),
    .B(_436__bF$buf5),
    .C(_451_),
    .Y(_72_)
);

NAND2X1 _2215_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [14]),
    .B(_436__bF$buf4),
    .Y(_452_)
);

OAI21X1 _2216_ (
    .A(_240_),
    .B(_436__bF$buf3),
    .C(_452_),
    .Y(_73_)
);

NAND2X1 _2217_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [15]),
    .B(_436__bF$buf2),
    .Y(_453_)
);

OAI21X1 _2218_ (
    .A(_246_),
    .B(_436__bF$buf1),
    .C(_453_),
    .Y(_74_)
);

INVX1 _2219_ (
    .A(q_1_loc_fu_40[17]),
    .Y(_454_)
);

NAND2X1 _2220_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [16]),
    .B(_436__bF$buf0),
    .Y(_455_)
);

OAI21X1 _2221_ (
    .A(_454_),
    .B(_436__bF$buf6),
    .C(_455_),
    .Y(_75_)
);

NAND2X1 _2222_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [17]),
    .B(_436__bF$buf5),
    .Y(_456_)
);

OAI21X1 _2223_ (
    .A(_261_),
    .B(_436__bF$buf4),
    .C(_456_),
    .Y(_76_)
);

NAND2X1 _2224_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [18]),
    .B(_436__bF$buf3),
    .Y(_457_)
);

OAI21X1 _2225_ (
    .A(_267_),
    .B(_436__bF$buf2),
    .C(_457_),
    .Y(_77_)
);

NAND2X1 _2226_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [19]),
    .B(_436__bF$buf1),
    .Y(_458_)
);

OAI21X1 _2227_ (
    .A(_279_),
    .B(_436__bF$buf0),
    .C(_458_),
    .Y(_78_)
);

NAND2X1 _2228_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [20]),
    .B(_436__bF$buf6),
    .Y(_459_)
);

OAI21X1 _2229_ (
    .A(_283_),
    .B(_436__bF$buf5),
    .C(_459_),
    .Y(_79_)
);

NAND2X1 _2230_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [21]),
    .B(_436__bF$buf4),
    .Y(_460_)
);

OAI21X1 _2231_ (
    .A(_290_),
    .B(_436__bF$buf3),
    .C(_460_),
    .Y(_80_)
);

NAND2X1 _2232_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [22]),
    .B(_436__bF$buf2),
    .Y(_461_)
);

OAI21X1 _2233_ (
    .A(_294_),
    .B(_436__bF$buf1),
    .C(_461_),
    .Y(_81_)
);

NAND2X1 _2234_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [23]),
    .B(_436__bF$buf0),
    .Y(_462_)
);

OAI21X1 _2235_ (
    .A(_307_),
    .B(_436__bF$buf6),
    .C(_462_),
    .Y(_82_)
);

NAND2X1 _2236_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [24]),
    .B(_436__bF$buf5),
    .Y(_463_)
);

OAI21X1 _2237_ (
    .A(_311_),
    .B(_436__bF$buf4),
    .C(_463_),
    .Y(_83_)
);

NAND2X1 _2238_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [25]),
    .B(_436__bF$buf3),
    .Y(_464_)
);

OAI21X1 _2239_ (
    .A(_321_),
    .B(_436__bF$buf2),
    .C(_464_),
    .Y(_84_)
);

NAND2X1 _2240_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [26]),
    .B(_436__bF$buf1),
    .Y(_465_)
);

OAI21X1 _2241_ (
    .A(_327_),
    .B(_436__bF$buf0),
    .C(_465_),
    .Y(_85_)
);

NAND2X1 _2242_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [27]),
    .B(_436__bF$buf6),
    .Y(_466_)
);

OAI21X1 _2243_ (
    .A(_330_),
    .B(_436__bF$buf5),
    .C(_466_),
    .Y(_86_)
);

AND2X2 _2244_ (
    .A(ap_CS_fsm_state2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0 ),
    .Y(_467_)
);

NAND2X1 _2245_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [0]),
    .B(_467__bF$buf6),
    .Y(_468_)
);

OAI21X1 _2246_ (
    .A(_116_),
    .B(_467__bF$buf5),
    .C(_468_),
    .Y(_88_)
);

NAND2X1 _2247_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [1]),
    .B(_467__bF$buf4),
    .Y(_469_)
);

OAI21X1 _2248_ (
    .A(_157_),
    .B(_467__bF$buf3),
    .C(_469_),
    .Y(_89_)
);

NAND2X1 _2249_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [2]),
    .B(_467__bF$buf2),
    .Y(_470_)
);

OAI21X1 _2250_ (
    .A(_162_),
    .B(_467__bF$buf1),
    .C(_470_),
    .Y(_90_)
);

NAND2X1 _2251_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [3]),
    .B(_467__bF$buf0),
    .Y(_471_)
);

OAI21X1 _2252_ (
    .A(_169_),
    .B(_467__bF$buf6),
    .C(_471_),
    .Y(_91_)
);

NAND2X1 _2253_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [4]),
    .B(_467__bF$buf5),
    .Y(_472_)
);

OAI21X1 _2254_ (
    .A(_174_),
    .B(_467__bF$buf4),
    .C(_472_),
    .Y(_92_)
);

NAND2X1 _2255_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [5]),
    .B(_467__bF$buf3),
    .Y(_473_)
);

OAI21X1 _2256_ (
    .A(_181_),
    .B(_467__bF$buf2),
    .C(_473_),
    .Y(_93_)
);

NAND2X1 _2257_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [6]),
    .B(_467__bF$buf1),
    .Y(_474_)
);

OAI21X1 _2258_ (
    .A(_186_),
    .B(_467__bF$buf0),
    .C(_474_),
    .Y(_94_)
);

NAND2X1 _2259_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [7]),
    .B(_467__bF$buf6),
    .Y(_475_)
);

OAI21X1 _2260_ (
    .A(_191_),
    .B(_467__bF$buf5),
    .C(_475_),
    .Y(_95_)
);

NAND2X1 _2261_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [8]),
    .B(_467__bF$buf4),
    .Y(_476_)
);

OAI21X1 _2262_ (
    .A(_200_),
    .B(_467__bF$buf3),
    .C(_476_),
    .Y(_96_)
);

NAND2X1 _2263_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [9]),
    .B(_467__bF$buf2),
    .Y(_477_)
);

OAI21X1 _2264_ (
    .A(_207_),
    .B(_467__bF$buf1),
    .C(_477_),
    .Y(_97_)
);

INVX1 _2265_ (
    .A(p_v_loc_fu_44[10]),
    .Y(_478_)
);

NAND2X1 _2266_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [10]),
    .B(_467__bF$buf0),
    .Y(_479_)
);

OAI21X1 _2267_ (
    .A(_478_),
    .B(_467__bF$buf6),
    .C(_479_),
    .Y(_98_)
);

NAND2X1 _2268_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [11]),
    .B(_467__bF$buf5),
    .Y(_480_)
);

OAI21X1 _2269_ (
    .A(_218_),
    .B(_467__bF$buf4),
    .C(_480_),
    .Y(_99_)
);

NAND2X1 _2270_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [12]),
    .B(_467__bF$buf3),
    .Y(_481_)
);

OAI21X1 _2271_ (
    .A(_226_),
    .B(_467__bF$buf2),
    .C(_481_),
    .Y(_100_)
);

NAND2X1 _2272_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [13]),
    .B(_467__bF$buf1),
    .Y(_482_)
);

OAI21X1 _2273_ (
    .A(_232_),
    .B(_467__bF$buf0),
    .C(_482_),
    .Y(_101_)
);

INVX1 _2274_ (
    .A(p_v_loc_fu_44[14]),
    .Y(_483_)
);

NAND2X1 _2275_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [14]),
    .B(_467__bF$buf6),
    .Y(_484_)
);

OAI21X1 _2276_ (
    .A(_483_),
    .B(_467__bF$buf5),
    .C(_484_),
    .Y(_102_)
);

NAND2X1 _2277_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [15]),
    .B(_467__bF$buf4),
    .Y(_485_)
);

OAI21X1 _2278_ (
    .A(_245_),
    .B(_467__bF$buf3),
    .C(_485_),
    .Y(_103_)
);

NAND2X1 _2279_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [16]),
    .B(_467__bF$buf2),
    .Y(_486_)
);

OAI21X1 _2280_ (
    .A(_256_),
    .B(_467__bF$buf1),
    .C(_486_),
    .Y(_104_)
);

NAND2X1 _2281_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [17]),
    .B(_467__bF$buf0),
    .Y(_487_)
);

OAI21X1 _2282_ (
    .A(_260_),
    .B(_467__bF$buf6),
    .C(_487_),
    .Y(_105_)
);

NAND2X1 _2283_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [18]),
    .B(_467__bF$buf5),
    .Y(_488_)
);

OAI21X1 _2284_ (
    .A(_266_),
    .B(_467__bF$buf4),
    .C(_488_),
    .Y(_106_)
);

NAND2X1 _2285_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [19]),
    .B(_467__bF$buf3),
    .Y(_489_)
);

OAI21X1 _2286_ (
    .A(_273_),
    .B(_467__bF$buf2),
    .C(_489_),
    .Y(_107_)
);

NAND2X1 _2287_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [20]),
    .B(_467__bF$buf1),
    .Y(_490_)
);

OAI21X1 _2288_ (
    .A(_282_),
    .B(_467__bF$buf0),
    .C(_490_),
    .Y(_108_)
);

INVX1 _2289_ (
    .A(p_v_loc_fu_44[21]),
    .Y(_491_)
);

NAND2X1 _2290_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [21]),
    .B(_467__bF$buf6),
    .Y(_492_)
);

OAI21X1 _2291_ (
    .A(_491_),
    .B(_467__bF$buf5),
    .C(_492_),
    .Y(_109_)
);

INVX1 _2292_ (
    .A(p_v_loc_fu_44[22]),
    .Y(_493_)
);

NAND2X1 _2293_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [22]),
    .B(_467__bF$buf4),
    .Y(_494_)
);

OAI21X1 _2294_ (
    .A(_493_),
    .B(_467__bF$buf3),
    .C(_494_),
    .Y(_110_)
);

NAND2X1 _2295_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [23]),
    .B(_467__bF$buf2),
    .Y(_495_)
);

OAI21X1 _2296_ (
    .A(_301_),
    .B(_467__bF$buf1),
    .C(_495_),
    .Y(_111_)
);

NAND2X1 _2297_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [24]),
    .B(_467__bF$buf0),
    .Y(_496_)
);

OAI21X1 _2298_ (
    .A(_310_),
    .B(_467__bF$buf6),
    .C(_496_),
    .Y(_112_)
);

NAND2X1 _2299_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [25]),
    .B(_467__bF$buf5),
    .Y(_497_)
);

OAI21X1 _2300_ (
    .A(_317_),
    .B(_467__bF$buf4),
    .C(_497_),
    .Y(_113_)
);

NAND2X1 _2301_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [26]),
    .B(_467__bF$buf3),
    .Y(_498_)
);

OAI21X1 _2302_ (
    .A(_324_),
    .B(_467__bF$buf2),
    .C(_498_),
    .Y(_114_)
);

NAND2X1 _2303_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [27]),
    .B(_467__bF$buf1),
    .Y(_499_)
);

OAI21X1 _2304_ (
    .A(_329_),
    .B(_467__bF$buf0),
    .C(_499_),
    .Y(_115_)
);

INVX1 _2305_ (
    .A(ap_rst),
    .Y(_500_)
);

NAND2X1 _2306_ (
    .A(ap_start),
    .B(ap_CS_fsm_state1_bF$buf6),
    .Y(_501_)
);

INVX1 _2307_ (
    .A(_501_),
    .Y(_502_)
);

NAND2X1 _2308_ (
    .A(ap_CS_fsm_state2),
    .B(_337_),
    .Y(_503_)
);

NOR2X1 _2309_ (
    .A(_1777_),
    .B(_503_),
    .Y(_504_)
);

OAI21X1 _2310_ (
    .A(_502_),
    .B(_504_),
    .C(_500_),
    .Y(_0_)
);

AOI21X1 _2311_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done ),
    .B(_501_),
    .C(_0_),
    .Y(_1_)
);

NAND3X1 _2312_ (
    .A(ap_CS_fsm_state2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done ),
    .C(_504_),
    .Y(_505_)
);

NOR2X1 _2313_ (
    .A(ap_rst),
    .B(_505_),
    .Y(_2_)
);

INVX1 _2314_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0 ),
    .Y(_506_)
);

NAND2X1 _2315_ (
    .A(grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58_ap_start_reg),
    .B(_506_),
    .Y(_507_)
);

AOI21X1 _2316_ (
    .A(_507_),
    .B(_501_),
    .C(ap_rst),
    .Y(_87_)
);

DFFPOSX1 _2317_ (
    .CLK(ap_clk_bF$buf12),
    .D(_0_),
    .Q(ap_CS_fsm_state1)
);

DFFPOSX1 _2318_ (
    .CLK(ap_clk_bF$buf11),
    .D(_1_),
    .Q(ap_CS_fsm_state2)
);

DFFPOSX1 _2319_ (
    .CLK(ap_clk_bF$buf10),
    .D(_2_),
    .Q(_1777_)
);

DFFPOSX1 _2320_ (
    .CLK(ap_clk_bF$buf9),
    .D(_3_),
    .Q(s_5_loc_fu_48[0])
);

DFFPOSX1 _2321_ (
    .CLK(ap_clk_bF$buf8),
    .D(_4_),
    .Q(s_5_loc_fu_48[1])
);

DFFPOSX1 _2322_ (
    .CLK(ap_clk_bF$buf7),
    .D(_5_),
    .Q(s_5_loc_fu_48[2])
);

DFFPOSX1 _2323_ (
    .CLK(ap_clk_bF$buf6),
    .D(_6_),
    .Q(s_5_loc_fu_48[3])
);

DFFPOSX1 _2324_ (
    .CLK(ap_clk_bF$buf5),
    .D(_7_),
    .Q(s_5_loc_fu_48[4])
);

DFFPOSX1 _2325_ (
    .CLK(ap_clk_bF$buf4),
    .D(_8_),
    .Q(s_5_loc_fu_48[5])
);

DFFPOSX1 _2326_ (
    .CLK(ap_clk_bF$buf3),
    .D(_9_),
    .Q(s_5_loc_fu_48[6])
);

DFFPOSX1 _2327_ (
    .CLK(ap_clk_bF$buf2),
    .D(_10_),
    .Q(s_5_loc_fu_48[7])
);

DFFPOSX1 _2328_ (
    .CLK(ap_clk_bF$buf1),
    .D(_11_),
    .Q(s_5_loc_fu_48[8])
);

DFFPOSX1 _2329_ (
    .CLK(ap_clk_bF$buf0),
    .D(_12_),
    .Q(s_5_loc_fu_48[9])
);

DFFPOSX1 _2330_ (
    .CLK(ap_clk_bF$buf12),
    .D(_13_),
    .Q(s_5_loc_fu_48[10])
);

DFFPOSX1 _2331_ (
    .CLK(ap_clk_bF$buf11),
    .D(_14_),
    .Q(s_5_loc_fu_48[11])
);

DFFPOSX1 _2332_ (
    .CLK(ap_clk_bF$buf10),
    .D(_15_),
    .Q(s_5_loc_fu_48[12])
);

DFFPOSX1 _2333_ (
    .CLK(ap_clk_bF$buf9),
    .D(_16_),
    .Q(s_5_loc_fu_48[13])
);

DFFPOSX1 _2334_ (
    .CLK(ap_clk_bF$buf8),
    .D(_17_),
    .Q(s_5_loc_fu_48[14])
);

DFFPOSX1 _2335_ (
    .CLK(ap_clk_bF$buf7),
    .D(_18_),
    .Q(s_5_loc_fu_48[15])
);

DFFPOSX1 _2336_ (
    .CLK(ap_clk_bF$buf6),
    .D(_19_),
    .Q(s_5_loc_fu_48[16])
);

DFFPOSX1 _2337_ (
    .CLK(ap_clk_bF$buf5),
    .D(_20_),
    .Q(s_5_loc_fu_48[17])
);

DFFPOSX1 _2338_ (
    .CLK(ap_clk_bF$buf4),
    .D(_21_),
    .Q(s_5_loc_fu_48[18])
);

DFFPOSX1 _2339_ (
    .CLK(ap_clk_bF$buf3),
    .D(_22_),
    .Q(s_5_loc_fu_48[19])
);

DFFPOSX1 _2340_ (
    .CLK(ap_clk_bF$buf2),
    .D(_23_),
    .Q(s_5_loc_fu_48[20])
);

DFFPOSX1 _2341_ (
    .CLK(ap_clk_bF$buf1),
    .D(_24_),
    .Q(s_5_loc_fu_48[21])
);

DFFPOSX1 _2342_ (
    .CLK(ap_clk_bF$buf0),
    .D(_25_),
    .Q(s_5_loc_fu_48[22])
);

DFFPOSX1 _2343_ (
    .CLK(ap_clk_bF$buf12),
    .D(_26_),
    .Q(s_5_loc_fu_48[23])
);

DFFPOSX1 _2344_ (
    .CLK(ap_clk_bF$buf11),
    .D(_27_),
    .Q(s_5_loc_fu_48[24])
);

DFFPOSX1 _2345_ (
    .CLK(ap_clk_bF$buf10),
    .D(_28_),
    .Q(s_5_loc_fu_48[25])
);

DFFPOSX1 _2346_ (
    .CLK(ap_clk_bF$buf9),
    .D(_29_),
    .Q(s_5_loc_fu_48[26])
);

DFFPOSX1 _2347_ (
    .CLK(ap_clk_bF$buf8),
    .D(_30_),
    .Q(s_5_loc_fu_48[27])
);

DFFPOSX1 _2348_ (
    .CLK(ap_clk_bF$buf7),
    .D(_31_),
    .Q(s_5_loc_fu_48[28])
);

DFFPOSX1 _2349_ (
    .CLK(ap_clk_bF$buf6),
    .D(_32_),
    .Q(s_5_loc_fu_48[29])
);

DFFPOSX1 _2350_ (
    .CLK(ap_clk_bF$buf5),
    .D(_33_),
    .Q(s_5_loc_fu_48[30])
);

DFFPOSX1 _2351_ (
    .CLK(ap_clk_bF$buf4),
    .D(_34_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [4])
);

DFFPOSX1 _2352_ (
    .CLK(ap_clk_bF$buf3),
    .D(_35_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [5])
);

DFFPOSX1 _2353_ (
    .CLK(ap_clk_bF$buf2),
    .D(_36_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [6])
);

DFFPOSX1 _2354_ (
    .CLK(ap_clk_bF$buf1),
    .D(_37_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [7])
);

DFFPOSX1 _2355_ (
    .CLK(ap_clk_bF$buf0),
    .D(_38_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [8])
);

DFFPOSX1 _2356_ (
    .CLK(ap_clk_bF$buf12),
    .D(_39_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [9])
);

DFFPOSX1 _2357_ (
    .CLK(ap_clk_bF$buf11),
    .D(_40_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [10])
);

DFFPOSX1 _2358_ (
    .CLK(ap_clk_bF$buf10),
    .D(_41_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [11])
);

DFFPOSX1 _2359_ (
    .CLK(ap_clk_bF$buf9),
    .D(_42_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [12])
);

DFFPOSX1 _2360_ (
    .CLK(ap_clk_bF$buf8),
    .D(_43_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [13])
);

DFFPOSX1 _2361_ (
    .CLK(ap_clk_bF$buf7),
    .D(_44_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [14])
);

DFFPOSX1 _2362_ (
    .CLK(ap_clk_bF$buf6),
    .D(_45_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [15])
);

DFFPOSX1 _2363_ (
    .CLK(ap_clk_bF$buf5),
    .D(_46_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [16])
);

DFFPOSX1 _2364_ (
    .CLK(ap_clk_bF$buf4),
    .D(_47_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [17])
);

DFFPOSX1 _2365_ (
    .CLK(ap_clk_bF$buf3),
    .D(_48_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [18])
);

DFFPOSX1 _2366_ (
    .CLK(ap_clk_bF$buf2),
    .D(_49_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [19])
);

DFFPOSX1 _2367_ (
    .CLK(ap_clk_bF$buf1),
    .D(_50_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [20])
);

DFFPOSX1 _2368_ (
    .CLK(ap_clk_bF$buf0),
    .D(_51_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [21])
);

DFFPOSX1 _2369_ (
    .CLK(ap_clk_bF$buf12),
    .D(_52_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [22])
);

DFFPOSX1 _2370_ (
    .CLK(ap_clk_bF$buf11),
    .D(_53_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [23])
);

DFFPOSX1 _2371_ (
    .CLK(ap_clk_bF$buf10),
    .D(_54_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [24])
);

DFFPOSX1 _2372_ (
    .CLK(ap_clk_bF$buf9),
    .D(_55_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [25])
);

DFFPOSX1 _2373_ (
    .CLK(ap_clk_bF$buf8),
    .D(_56_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [26])
);

DFFPOSX1 _2374_ (
    .CLK(ap_clk_bF$buf7),
    .D(_57_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [27])
);

DFFPOSX1 _2375_ (
    .CLK(ap_clk_bF$buf6),
    .D(_58_),
    .Q(q_1_loc_fu_40[0])
);

DFFPOSX1 _2376_ (
    .CLK(ap_clk_bF$buf5),
    .D(_59_),
    .Q(q_1_loc_fu_40[1])
);

DFFPOSX1 _2377_ (
    .CLK(ap_clk_bF$buf4),
    .D(_60_),
    .Q(q_1_loc_fu_40[2])
);

DFFPOSX1 _2378_ (
    .CLK(ap_clk_bF$buf3),
    .D(_61_),
    .Q(q_1_loc_fu_40[3])
);

DFFPOSX1 _2379_ (
    .CLK(ap_clk_bF$buf2),
    .D(_62_),
    .Q(q_1_loc_fu_40[4])
);

DFFPOSX1 _2380_ (
    .CLK(ap_clk_bF$buf1),
    .D(_63_),
    .Q(q_1_loc_fu_40[5])
);

DFFPOSX1 _2381_ (
    .CLK(ap_clk_bF$buf0),
    .D(_64_),
    .Q(q_1_loc_fu_40[6])
);

DFFPOSX1 _2382_ (
    .CLK(ap_clk_bF$buf12),
    .D(_65_),
    .Q(q_1_loc_fu_40[7])
);

DFFPOSX1 _2383_ (
    .CLK(ap_clk_bF$buf11),
    .D(_66_),
    .Q(q_1_loc_fu_40[8])
);

DFFPOSX1 _2384_ (
    .CLK(ap_clk_bF$buf10),
    .D(_67_),
    .Q(q_1_loc_fu_40[9])
);

DFFPOSX1 _2385_ (
    .CLK(ap_clk_bF$buf9),
    .D(_68_),
    .Q(q_1_loc_fu_40[10])
);

DFFPOSX1 _2386_ (
    .CLK(ap_clk_bF$buf8),
    .D(_69_),
    .Q(q_1_loc_fu_40[11])
);

DFFPOSX1 _2387_ (
    .CLK(ap_clk_bF$buf7),
    .D(_70_),
    .Q(q_1_loc_fu_40[12])
);

DFFPOSX1 _2388_ (
    .CLK(ap_clk_bF$buf6),
    .D(_71_),
    .Q(q_1_loc_fu_40[13])
);

DFFPOSX1 _2389_ (
    .CLK(ap_clk_bF$buf5),
    .D(_72_),
    .Q(q_1_loc_fu_40[14])
);

DFFPOSX1 _2390_ (
    .CLK(ap_clk_bF$buf4),
    .D(_73_),
    .Q(q_1_loc_fu_40[15])
);

DFFPOSX1 _2391_ (
    .CLK(ap_clk_bF$buf3),
    .D(_74_),
    .Q(q_1_loc_fu_40[16])
);

DFFPOSX1 _2392_ (
    .CLK(ap_clk_bF$buf2),
    .D(_75_),
    .Q(q_1_loc_fu_40[17])
);

DFFPOSX1 _2393_ (
    .CLK(ap_clk_bF$buf1),
    .D(_76_),
    .Q(q_1_loc_fu_40[18])
);

DFFPOSX1 _2394_ (
    .CLK(ap_clk_bF$buf0),
    .D(_77_),
    .Q(q_1_loc_fu_40[19])
);

DFFPOSX1 _2395_ (
    .CLK(ap_clk_bF$buf12),
    .D(_78_),
    .Q(q_1_loc_fu_40[20])
);

DFFPOSX1 _2396_ (
    .CLK(ap_clk_bF$buf11),
    .D(_79_),
    .Q(q_1_loc_fu_40[21])
);

DFFPOSX1 _2397_ (
    .CLK(ap_clk_bF$buf10),
    .D(_80_),
    .Q(q_1_loc_fu_40[22])
);

DFFPOSX1 _2398_ (
    .CLK(ap_clk_bF$buf9),
    .D(_81_),
    .Q(q_1_loc_fu_40[23])
);

DFFPOSX1 _2399_ (
    .CLK(ap_clk_bF$buf8),
    .D(_82_),
    .Q(q_1_loc_fu_40[24])
);

DFFPOSX1 _2400_ (
    .CLK(ap_clk_bF$buf7),
    .D(_83_),
    .Q(q_1_loc_fu_40[25])
);

DFFPOSX1 _2401_ (
    .CLK(ap_clk_bF$buf6),
    .D(_84_),
    .Q(q_1_loc_fu_40[26])
);

DFFPOSX1 _2402_ (
    .CLK(ap_clk_bF$buf5),
    .D(_85_),
    .Q(q_1_loc_fu_40[27])
);

DFFPOSX1 _2403_ (
    .CLK(ap_clk_bF$buf4),
    .D(_86_),
    .Q(q_1_loc_fu_40[28])
);

DFFPOSX1 _2404_ (
    .CLK(ap_clk_bF$buf3),
    .D(_87_),
    .Q(grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58_ap_start_reg)
);

DFFPOSX1 _2405_ (
    .CLK(ap_clk_bF$buf2),
    .D(_88_),
    .Q(p_v_loc_fu_44[0])
);

DFFPOSX1 _2406_ (
    .CLK(ap_clk_bF$buf1),
    .D(_89_),
    .Q(p_v_loc_fu_44[1])
);

DFFPOSX1 _2407_ (
    .CLK(ap_clk_bF$buf0),
    .D(_90_),
    .Q(p_v_loc_fu_44[2])
);

DFFPOSX1 _2408_ (
    .CLK(ap_clk_bF$buf12),
    .D(_91_),
    .Q(p_v_loc_fu_44[3])
);

DFFPOSX1 _2409_ (
    .CLK(ap_clk_bF$buf11),
    .D(_92_),
    .Q(p_v_loc_fu_44[4])
);

DFFPOSX1 _2410_ (
    .CLK(ap_clk_bF$buf10),
    .D(_93_),
    .Q(p_v_loc_fu_44[5])
);

DFFPOSX1 _2411_ (
    .CLK(ap_clk_bF$buf9),
    .D(_94_),
    .Q(p_v_loc_fu_44[6])
);

DFFPOSX1 _2412_ (
    .CLK(ap_clk_bF$buf8),
    .D(_95_),
    .Q(p_v_loc_fu_44[7])
);

DFFPOSX1 _2413_ (
    .CLK(ap_clk_bF$buf7),
    .D(_96_),
    .Q(p_v_loc_fu_44[8])
);

DFFPOSX1 _2414_ (
    .CLK(ap_clk_bF$buf6),
    .D(_97_),
    .Q(p_v_loc_fu_44[9])
);

DFFPOSX1 _2415_ (
    .CLK(ap_clk_bF$buf5),
    .D(_98_),
    .Q(p_v_loc_fu_44[10])
);

DFFPOSX1 _2416_ (
    .CLK(ap_clk_bF$buf4),
    .D(_99_),
    .Q(p_v_loc_fu_44[11])
);

DFFPOSX1 _2417_ (
    .CLK(ap_clk_bF$buf3),
    .D(_100_),
    .Q(p_v_loc_fu_44[12])
);

DFFPOSX1 _2418_ (
    .CLK(ap_clk_bF$buf2),
    .D(_101_),
    .Q(p_v_loc_fu_44[13])
);

DFFPOSX1 _2419_ (
    .CLK(ap_clk_bF$buf1),
    .D(_102_),
    .Q(p_v_loc_fu_44[14])
);

DFFPOSX1 _2420_ (
    .CLK(ap_clk_bF$buf0),
    .D(_103_),
    .Q(p_v_loc_fu_44[15])
);

DFFPOSX1 _2421_ (
    .CLK(ap_clk_bF$buf12),
    .D(_104_),
    .Q(p_v_loc_fu_44[16])
);

DFFPOSX1 _2422_ (
    .CLK(ap_clk_bF$buf11),
    .D(_105_),
    .Q(p_v_loc_fu_44[17])
);

DFFPOSX1 _2423_ (
    .CLK(ap_clk_bF$buf10),
    .D(_106_),
    .Q(p_v_loc_fu_44[18])
);

DFFPOSX1 _2424_ (
    .CLK(ap_clk_bF$buf9),
    .D(_107_),
    .Q(p_v_loc_fu_44[19])
);

DFFPOSX1 _2425_ (
    .CLK(ap_clk_bF$buf8),
    .D(_108_),
    .Q(p_v_loc_fu_44[20])
);

DFFPOSX1 _2426_ (
    .CLK(ap_clk_bF$buf7),
    .D(_109_),
    .Q(p_v_loc_fu_44[21])
);

DFFPOSX1 _2427_ (
    .CLK(ap_clk_bF$buf6),
    .D(_110_),
    .Q(p_v_loc_fu_44[22])
);

DFFPOSX1 _2428_ (
    .CLK(ap_clk_bF$buf5),
    .D(_111_),
    .Q(p_v_loc_fu_44[23])
);

DFFPOSX1 _2429_ (
    .CLK(ap_clk_bF$buf4),
    .D(_112_),
    .Q(p_v_loc_fu_44[24])
);

DFFPOSX1 _2430_ (
    .CLK(ap_clk_bF$buf3),
    .D(_113_),
    .Q(p_v_loc_fu_44[25])
);

DFFPOSX1 _2431_ (
    .CLK(ap_clk_bF$buf2),
    .D(_114_),
    .Q(p_v_loc_fu_44[26])
);

DFFPOSX1 _2432_ (
    .CLK(ap_clk_bF$buf1),
    .D(_115_),
    .Q(p_v_loc_fu_44[27])
);

INVX1 _2433_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_enable_reg_pp0_iter1 ),
    .Y(_1021_)
);

INVX8 _2434_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .Y(_1022_)
);

NAND2X1 _2435_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_1022__bF$buf6),
    .Y(_1023_)
);

NAND2X1 _2436_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .Y(_1024_)
);

NOR2X1 _2437_ (
    .A(_1024_),
    .B(_1023_),
    .Y(_1025_)
);

NAND2X1 _2438_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(_1025_),
    .Y(_1026_)
);

NOR2X1 _2439_ (
    .A(_1021_),
    .B(_1026_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0 )
);

INVX8 _2440_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .Y(_1027_)
);

NAND2X1 _2441_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [0]),
    .B(_1027__bF$buf5),
    .Y(_1028_)
);

INVX1 _2442_ (
    .A(_1028_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [0])
);

INVX1 _2443_ (
    .A(_1026_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_1_fu_177_p2 [0])
);

INVX2 _2444_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .Y(_1029_)
);

INVX1 _2445_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [0]),
    .Y(_1030_)
);

AOI21X1 _2446_ (
    .A(_1027__bF$buf4),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .Y(_1031_)
);

NAND3X1 _2447_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .C(_1031_),
    .Y(_1032_)
);

OAI21X1 _2448_ (
    .A(_1029_),
    .B(_1032_),
    .C(_1030_),
    .Y(_1033_)
);

INVX4 _2449_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .Y(_1034_)
);

OAI21X1 _2450_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .B(_1034__bF$buf3),
    .C(_1022__bF$buf5),
    .Y(_1035_)
);

NOR2X1 _2451_ (
    .A(_1024_),
    .B(_1035_),
    .Y(_1036_)
);

NAND3X1 _2452_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [0]),
    .C(_1036_),
    .Y(_1037_)
);

NAND2X1 _2453_ (
    .A(_1037_),
    .B(_1033_),
    .Y(_1038_)
);

INVX1 _2454_ (
    .A(_1038_),
    .Y(_1039_)
);

OAI21X1 _2455_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .B(_1026_),
    .C(_1039_),
    .Y(_1040_)
);

NAND3X1 _2456_ (
    .A(_1027__bF$buf3),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_1_fu_177_p2 [0]),
    .C(_1038_),
    .Y(_1041_)
);

NAND2X1 _2457_ (
    .A(_1041_),
    .B(_1040_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [1])
);

OAI21X1 _2458_ (
    .A(_1022__bF$buf4),
    .B(_1024_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .Y(_1042_)
);

AND2X2 _2459_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .Y(_1043_)
);

NAND2X1 _2460_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .B(_1043_),
    .Y(_1044_)
);

OR2X2 _2461_ (
    .A(_1044_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .Y(_1045_)
);

NAND2X1 _2462_ (
    .A(_1042_),
    .B(_1045_),
    .Y(_1046_)
);

INVX1 _2463_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .Y(_1047_)
);

INVX2 _2464_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .Y(_1048_)
);

OAI21X1 _2465_ (
    .A(_1022__bF$buf3),
    .B(_1048_),
    .C(_1047_),
    .Y(_1049_)
);

OAI21X1 _2466_ (
    .A(_1022__bF$buf2),
    .B(_1024_),
    .C(_1049_),
    .Y(_1050_)
);

NOR2X1 _2467_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .Y(_1051_)
);

NOR2X1 _2468_ (
    .A(_1051_),
    .B(_1043_),
    .Y(_1052_)
);

NAND2X1 _2469_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_1034__bF$buf2),
    .Y(_1053_)
);

NAND3X1 _2470_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [0]),
    .C(_1027__bF$buf2),
    .Y(_1054_)
);

NAND2X1 _2471_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .B(_1034__bF$buf1),
    .Y(_1055_)
);

NAND3X1 _2472_ (
    .A(_1022__bF$buf1),
    .B(_1055_),
    .C(_1054_),
    .Y(_1056_)
);

NAND3X1 _2473_ (
    .A(_1052__bF$buf5),
    .B(_1053_),
    .C(_1056_),
    .Y(_1057_)
);

NOR2X1 _2474_ (
    .A(_1050__bF$buf5),
    .B(_1057_),
    .Y(_1058_)
);

NAND3X1 _2475_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [1]),
    .B(_1046__bF$buf7),
    .C(_1058_),
    .Y(_1059_)
);

INVX1 _2476_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [1]),
    .Y(_1060_)
);

OAI21X1 _2477_ (
    .A(_1022__bF$buf0),
    .B(_1024_),
    .C(_1029_),
    .Y(_1061_)
);

OR2X2 _2478_ (
    .A(_1044_),
    .B(_1029_),
    .Y(_1062_)
);

NAND2X1 _2479_ (
    .A(_1061_),
    .B(_1062_),
    .Y(_1063_)
);

AND2X2 _2480_ (
    .A(_1044_),
    .B(_1049_),
    .Y(_1064_)
);

NAND2X1 _2481_ (
    .A(_1023_),
    .B(_1053_),
    .Y(_1065_)
);

AOI22X1 _2482_ (
    .A(_1034__bF$buf0),
    .B(_1027__bF$buf1),
    .C(_1065_),
    .D(_1028_),
    .Y(_1066_)
);

NAND3X1 _2483_ (
    .A(_1052__bF$buf4),
    .B(_1064__bF$buf5),
    .C(_1066_),
    .Y(_1067_)
);

OAI21X1 _2484_ (
    .A(_1063__bF$buf4),
    .B(_1067_),
    .C(_1060_),
    .Y(_1068_)
);

NAND2X1 _2485_ (
    .A(_1068_),
    .B(_1059_),
    .Y(_1069_)
);

OAI21X1 _2486_ (
    .A(_1029_),
    .B(_1032_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [0]),
    .Y(_1070_)
);

INVX1 _2487_ (
    .A(_1070_),
    .Y(_1071_)
);

AOI21X1 _2488_ (
    .A(_1038_),
    .B(_1026_),
    .C(_1071_),
    .Y(_1072_)
);

NAND2X1 _2489_ (
    .A(_1027__bF$buf0),
    .B(_1072_),
    .Y(_1073_)
);

OAI21X1 _2490_ (
    .A(_1027__bF$buf5),
    .B(_1037_),
    .C(_1073_),
    .Y(_1074_)
);

NAND2X1 _2491_ (
    .A(_1069_),
    .B(_1074_),
    .Y(_1075_)
);

OR2X2 _2492_ (
    .A(_1074_),
    .B(_1069_),
    .Y(_1076_)
);

NAND2X1 _2493_ (
    .A(_1075_),
    .B(_1076_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [2])
);

NAND2X1 _2494_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [1]),
    .Y(_1077_)
);

NAND3X1 _2495_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [0]),
    .B(_1034__bF$buf3),
    .C(_1027__bF$buf4),
    .Y(_1078_)
);

NAND3X1 _2496_ (
    .A(_1022__bF$buf6),
    .B(_1077_),
    .C(_1078_),
    .Y(_1079_)
);

NAND3X1 _2497_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .C(_1027__bF$buf3),
    .Y(_1080_)
);

NAND3X1 _2498_ (
    .A(_1052__bF$buf3),
    .B(_1080_),
    .C(_1079_),
    .Y(_1081_)
);

NOR2X1 _2499_ (
    .A(_1050__bF$buf4),
    .B(_1081_),
    .Y(_1082_)
);

NAND3X1 _2500_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [2]),
    .B(_1046__bF$buf6),
    .C(_1082_),
    .Y(_1083_)
);

INVX1 _2501_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [2]),
    .Y(_1084_)
);

NAND2X1 _2502_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .Y(_1085_)
);

NAND2X1 _2503_ (
    .A(_1022__bF$buf5),
    .B(_1048_),
    .Y(_1086_)
);

NAND2X1 _2504_ (
    .A(_1085_),
    .B(_1086_),
    .Y(_1087_)
);

OAI21X1 _2505_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .B(_1034__bF$buf2),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .Y(_1088_)
);

INVX1 _2506_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [0]),
    .Y(_1089_)
);

OAI21X1 _2507_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .B(_1089_),
    .C(_1034__bF$buf1),
    .Y(_1090_)
);

INVX1 _2508_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [1]),
    .Y(_1091_)
);

NAND2X1 _2509_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(_1091_),
    .Y(_1092_)
);

NAND3X1 _2510_ (
    .A(_1022__bF$buf4),
    .B(_1092_),
    .C(_1090_),
    .Y(_1093_)
);

AOI21X1 _2511_ (
    .A(_1093_),
    .B(_1088_),
    .C(_1087__bF$buf4),
    .Y(_1094_)
);

NAND2X1 _2512_ (
    .A(_1064__bF$buf4),
    .B(_1094_),
    .Y(_1095_)
);

OAI21X1 _2513_ (
    .A(_1063__bF$buf3),
    .B(_1095_),
    .C(_1084_),
    .Y(_1096_)
);

NAND2X1 _2514_ (
    .A(_1083_),
    .B(_1096_),
    .Y(_1097_)
);

OAI21X1 _2515_ (
    .A(_1037_),
    .B(_1069_),
    .C(_1059_),
    .Y(_1098_)
);

OAI21X1 _2516_ (
    .A(_1063__bF$buf2),
    .B(_1067_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [1]),
    .Y(_1099_)
);

NOR3X1 _2517_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [1]),
    .B(_1063__bF$buf1),
    .C(_1067_),
    .Y(_1100_)
);

OAI21X1 _2518_ (
    .A(_1072_),
    .B(_1100_),
    .C(_1099_),
    .Y(_1101_)
);

NAND2X1 _2519_ (
    .A(_1027__bF$buf2),
    .B(_1101_),
    .Y(_1102_)
);

OAI21X1 _2520_ (
    .A(_1027__bF$buf1),
    .B(_1098_),
    .C(_1102_),
    .Y(_1103_)
);

AND2X2 _2521_ (
    .A(_1103_),
    .B(_1097_),
    .Y(_1104_)
);

NOR2X1 _2522_ (
    .A(_1097_),
    .B(_1103_),
    .Y(_1105_)
);

NOR2X1 _2523_ (
    .A(_1105_),
    .B(_1104_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [3])
);

NAND3X1 _2524_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(_1055_),
    .C(_1054_),
    .Y(_1106_)
);

MUX2X1 _2525_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [2]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [1]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .Y(_1107_)
);

NAND2X1 _2526_ (
    .A(_1022__bF$buf3),
    .B(_1107_),
    .Y(_1108_)
);

NAND3X1 _2527_ (
    .A(_1052__bF$buf2),
    .B(_1106_),
    .C(_1108_),
    .Y(_1109_)
);

NAND2X1 _2528_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_1051_),
    .Y(_1110_)
);

AOI21X1 _2529_ (
    .A(_1109_),
    .B(_1110_),
    .C(_1050__bF$buf3),
    .Y(_1111_)
);

NAND3X1 _2530_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [3]),
    .B(_1046__bF$buf5),
    .C(_1111_),
    .Y(_1112_)
);

INVX1 _2531_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [3]),
    .Y(_1113_)
);

NAND2X1 _2532_ (
    .A(_1034__bF$buf0),
    .B(_1091_),
    .Y(_1114_)
);

INVX1 _2533_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [2]),
    .Y(_1115_)
);

NAND2X1 _2534_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(_1115_),
    .Y(_1116_)
);

NAND3X1 _2535_ (
    .A(_1022__bF$buf2),
    .B(_1116_),
    .C(_1114_),
    .Y(_1117_)
);

NAND2X1 _2536_ (
    .A(_1034__bF$buf3),
    .B(_1027__bF$buf0),
    .Y(_1118_)
);

OAI21X1 _2537_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .B(_1089_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .Y(_1119_)
);

NAND3X1 _2538_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_1118_),
    .C(_1119_),
    .Y(_1120_)
);

NAND3X1 _2539_ (
    .A(_1052__bF$buf1),
    .B(_1117_),
    .C(_1120_),
    .Y(_1121_)
);

OAI21X1 _2540_ (
    .A(_1043_),
    .B(_1051_),
    .C(_1023_),
    .Y(_1122_)
);

NAND3X1 _2541_ (
    .A(_1064__bF$buf3),
    .B(_1122_),
    .C(_1121_),
    .Y(_1123_)
);

OAI21X1 _2542_ (
    .A(_1063__bF$buf0),
    .B(_1123_),
    .C(_1113_),
    .Y(_1124_)
);

AND2X2 _2543_ (
    .A(_1124_),
    .B(_1112_),
    .Y(_1125_)
);

AOI21X1 _2544_ (
    .A(_1082_),
    .B(_1046__bF$buf4),
    .C(_1084_),
    .Y(_1126_)
);

AOI21X1 _2545_ (
    .A(_1101_),
    .B(_1097_),
    .C(_1126_),
    .Y(_1127_)
);

INVX1 _2546_ (
    .A(_1037_),
    .Y(_1128_)
);

NAND2X1 _2547_ (
    .A(_1128_),
    .B(_1068_),
    .Y(_1129_)
);

AND2X2 _2548_ (
    .A(_1129_),
    .B(_1059_),
    .Y(_1130_)
);

OAI21X1 _2549_ (
    .A(_1097_),
    .B(_1130_),
    .C(_1083_),
    .Y(_1131_)
);

MUX2X1 _2550_ (
    .A(_1131_),
    .B(_1127_),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .Y(_1132_)
);

OR2X2 _2551_ (
    .A(_1132_),
    .B(_1125_),
    .Y(_1133_)
);

NAND2X1 _2552_ (
    .A(_1125_),
    .B(_1132_),
    .Y(_1134_)
);

NAND2X1 _2553_ (
    .A(_1134_),
    .B(_1133_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [4])
);

NAND3X1 _2554_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_1092_),
    .C(_1090_),
    .Y(_1135_)
);

NAND2X1 _2555_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [3]),
    .Y(_1136_)
);

OAI21X1 _2556_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(_1115_),
    .C(_1136_),
    .Y(_1137_)
);

NAND2X1 _2557_ (
    .A(_1022__bF$buf1),
    .B(_1137_),
    .Y(_1138_)
);

NAND3X1 _2558_ (
    .A(_1052__bF$buf0),
    .B(_1138_),
    .C(_1135_),
    .Y(_1139_)
);

OAI21X1 _2559_ (
    .A(_1043_),
    .B(_1051_),
    .C(_1035_),
    .Y(_1140_)
);

NAND3X1 _2560_ (
    .A(_1064__bF$buf2),
    .B(_1140_),
    .C(_1139_),
    .Y(_1141_)
);

OAI21X1 _2561_ (
    .A(_1029_),
    .B(_1141_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [4]),
    .Y(_1142_)
);

INVX1 _2562_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [4]),
    .Y(_1143_)
);

MUX2X1 _2563_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [3]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [2]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .Y(_1144_)
);

NAND2X1 _2564_ (
    .A(_1022__bF$buf0),
    .B(_1144_),
    .Y(_1145_)
);

NAND3X1 _2565_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .B(_1077_),
    .C(_1078_),
    .Y(_1146_)
);

NAND3X1 _2566_ (
    .A(_1052__bF$buf5),
    .B(_1145_),
    .C(_1146_),
    .Y(_1147_)
);

OAI21X1 _2567_ (
    .A(_1034__bF$buf2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .C(_1051_),
    .Y(_1148_)
);

AOI21X1 _2568_ (
    .A(_1147_),
    .B(_1148_),
    .C(_1050__bF$buf2),
    .Y(_1149_)
);

NAND3X1 _2569_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(_1143_),
    .C(_1149_),
    .Y(_1150_)
);

NAND2X1 _2570_ (
    .A(_1150_),
    .B(_1142_),
    .Y(_1151_)
);

INVX1 _2571_ (
    .A(_1151_),
    .Y(_1152_)
);

INVX1 _2572_ (
    .A(_1126_),
    .Y(_1153_)
);

NAND3X1 _2573_ (
    .A(_1084_),
    .B(_1046__bF$buf3),
    .C(_1082_),
    .Y(_1154_)
);

NAND2X1 _2574_ (
    .A(_1112_),
    .B(_1124_),
    .Y(_1155_)
);

AOI21X1 _2575_ (
    .A(_1153_),
    .B(_1154_),
    .C(_1155_),
    .Y(_1156_)
);

OAI21X1 _2576_ (
    .A(_1083_),
    .B(_1155_),
    .C(_1112_),
    .Y(_1157_)
);

AOI21X1 _2577_ (
    .A(_1156_),
    .B(_1098_),
    .C(_1157_),
    .Y(_1158_)
);

OAI21X1 _2578_ (
    .A(_1063__bF$buf4),
    .B(_1123_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [3]),
    .Y(_1159_)
);

AND2X2 _2579_ (
    .A(_1159_),
    .B(_1027__bF$buf5),
    .Y(_1160_)
);

OAI21X1 _2580_ (
    .A(_1125_),
    .B(_1127_),
    .C(_1160_),
    .Y(_1161_)
);

OAI21X1 _2581_ (
    .A(_1027__bF$buf4),
    .B(_1158_),
    .C(_1161_),
    .Y(_1162_)
);

OR2X2 _2582_ (
    .A(_1162_),
    .B(_1152_),
    .Y(_1163_)
);

NAND2X1 _2583_ (
    .A(_1152_),
    .B(_1162_),
    .Y(_1164_)
);

NAND2X1 _2584_ (
    .A(_1164_),
    .B(_1163_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [5])
);

INVX1 _2585_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [5]),
    .Y(_1165_)
);

MUX2X1 _2586_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [4]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [3]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .Y(_1166_)
);

NAND2X1 _2587_ (
    .A(_1022__bF$buf6),
    .B(_1166_),
    .Y(_1167_)
);

NAND2X1 _2588_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(_1107_),
    .Y(_1168_)
);

NAND3X1 _2589_ (
    .A(_1052__bF$buf4),
    .B(_1167_),
    .C(_1168_),
    .Y(_1169_)
);

NAND3X1 _2590_ (
    .A(_1087__bF$buf3),
    .B(_1053_),
    .C(_1056_),
    .Y(_1170_)
);

AOI21X1 _2591_ (
    .A(_1169_),
    .B(_1170_),
    .C(_1050__bF$buf1),
    .Y(_1171_)
);

AOI21X1 _2592_ (
    .A(_1171_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .C(_1165_),
    .Y(_1172_)
);

NAND3X1 _2593_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .B(_1116_),
    .C(_1114_),
    .Y(_1173_)
);

INVX1 _2594_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [3]),
    .Y(_1174_)
);

NAND2X1 _2595_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [4]),
    .Y(_1175_)
);

OAI21X1 _2596_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_1174_),
    .C(_1175_),
    .Y(_1176_)
);

NAND2X1 _2597_ (
    .A(_1022__bF$buf5),
    .B(_1176_),
    .Y(_1177_)
);

NAND3X1 _2598_ (
    .A(_1052__bF$buf3),
    .B(_1173_),
    .C(_1177_),
    .Y(_1178_)
);

NAND2X1 _2599_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .Y(_1179_)
);

NAND3X1 _2600_ (
    .A(_1022__bF$buf4),
    .B(_1118_),
    .C(_1119_),
    .Y(_1180_)
);

NAND3X1 _2601_ (
    .A(_1087__bF$buf2),
    .B(_1179_),
    .C(_1180_),
    .Y(_1181_)
);

NAND3X1 _2602_ (
    .A(_1064__bF$buf1),
    .B(_1178_),
    .C(_1181_),
    .Y(_1182_)
);

NOR3X1 _2603_ (
    .A(_1029_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [5]),
    .C(_1182_),
    .Y(_1183_)
);

NOR3X1 _2604_ (
    .A(_1029_),
    .B(_1143_),
    .C(_1141_),
    .Y(_1184_)
);

NOR2X1 _2605_ (
    .A(_1027__bF$buf3),
    .B(_1184_),
    .Y(_1185_)
);

OAI21X1 _2606_ (
    .A(_1152_),
    .B(_1158_),
    .C(_1185_),
    .Y(_1186_)
);

INVX1 _2607_ (
    .A(_1072_),
    .Y(_1187_)
);

NAND3X1 _2608_ (
    .A(_1069_),
    .B(_1187_),
    .C(_1097_),
    .Y(_1188_)
);

INVX1 _2609_ (
    .A(_1099_),
    .Y(_1189_)
);

AOI21X1 _2610_ (
    .A(_1189_),
    .B(_1154_),
    .C(_1126_),
    .Y(_1190_)
);

NAND3X1 _2611_ (
    .A(_1142_),
    .B(_1150_),
    .C(_1155_),
    .Y(_1191_)
);

AOI21X1 _2612_ (
    .A(_1188_),
    .B(_1190_),
    .C(_1191_),
    .Y(_1192_)
);

OAI21X1 _2613_ (
    .A(_1159_),
    .B(_1151_),
    .C(_1142_),
    .Y(_1193_)
);

NOR2X1 _2614_ (
    .A(_1193_),
    .B(_1192_),
    .Y(_1194_)
);

OAI21X1 _2615_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .B(_1194_),
    .C(_1186_),
    .Y(_1195_)
);

OAI21X1 _2616_ (
    .A(_1172_),
    .B(_1183_),
    .C(_1195_),
    .Y(_1196_)
);

OAI21X1 _2617_ (
    .A(_1029_),
    .B(_1182_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [5]),
    .Y(_1197_)
);

NAND3X1 _2618_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(_1165_),
    .C(_1171_),
    .Y(_1198_)
);

NAND2X1 _2619_ (
    .A(_1198_),
    .B(_1197_),
    .Y(_1199_)
);

OR2X2 _2620_ (
    .A(_1195_),
    .B(_1199_),
    .Y(_1200_)
);

NAND2X1 _2621_ (
    .A(_1196_),
    .B(_1200_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [6])
);

MUX2X1 _2622_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [5]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [4]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .Y(_1201_)
);

MUX2X1 _2623_ (
    .A(_1201_),
    .B(_1144_),
    .S(_1022__bF$buf3),
    .Y(_1202_)
);

NAND2X1 _2624_ (
    .A(_1052__bF$buf2),
    .B(_1202_),
    .Y(_1203_)
);

NAND3X1 _2625_ (
    .A(_1087__bF$buf1),
    .B(_1080_),
    .C(_1079_),
    .Y(_1204_)
);

AOI21X1 _2626_ (
    .A(_1203_),
    .B(_1204_),
    .C(_1050__bF$buf0),
    .Y(_1205_)
);

NAND3X1 _2627_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [6]),
    .B(_1046__bF$buf2),
    .C(_1205_),
    .Y(_1206_)
);

INVX1 _2628_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [6]),
    .Y(_1207_)
);

NAND2X1 _2629_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_1137_),
    .Y(_1208_)
);

INVX1 _2630_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [4]),
    .Y(_1209_)
);

NAND2X1 _2631_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [5]),
    .Y(_1210_)
);

OAI21X1 _2632_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(_1209_),
    .C(_1210_),
    .Y(_1211_)
);

NAND2X1 _2633_ (
    .A(_1022__bF$buf2),
    .B(_1211_),
    .Y(_1212_)
);

NAND3X1 _2634_ (
    .A(_1052__bF$buf1),
    .B(_1208_),
    .C(_1212_),
    .Y(_1213_)
);

NAND3X1 _2635_ (
    .A(_1087__bF$buf0),
    .B(_1088_),
    .C(_1093_),
    .Y(_1214_)
);

NAND3X1 _2636_ (
    .A(_1064__bF$buf0),
    .B(_1213_),
    .C(_1214_),
    .Y(_1215_)
);

OAI21X1 _2637_ (
    .A(_1063__bF$buf3),
    .B(_1215_),
    .C(_1207_),
    .Y(_1216_)
);

NAND2X1 _2638_ (
    .A(_1216_),
    .B(_1206_),
    .Y(_1217_)
);

NAND2X1 _2639_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(_1171_),
    .Y(_1218_)
);

NOR2X1 _2640_ (
    .A(_1165_),
    .B(_1218_),
    .Y(_1219_)
);

AOI21X1 _2641_ (
    .A(_1199_),
    .B(_1184_),
    .C(_1219_),
    .Y(_1220_)
);

AOI22X1 _2642_ (
    .A(_1142_),
    .B(_1150_),
    .C(_1197_),
    .D(_1198_),
    .Y(_1221_)
);

INVX1 _2643_ (
    .A(_1221_),
    .Y(_1222_)
);

OAI21X1 _2644_ (
    .A(_1222_),
    .B(_1158_),
    .C(_1220_),
    .Y(_1223_)
);

NAND2X1 _2645_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .B(_1223_),
    .Y(_1224_)
);

NOR2X1 _2646_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .B(_1172_),
    .Y(_1225_)
);

OAI21X1 _2647_ (
    .A(_1199_),
    .B(_1194_),
    .C(_1225_),
    .Y(_1226_)
);

NAND2X1 _2648_ (
    .A(_1224_),
    .B(_1226_),
    .Y(_1227_)
);

OR2X2 _2649_ (
    .A(_1227_),
    .B(_1217_),
    .Y(_1228_)
);

NAND2X1 _2650_ (
    .A(_1217_),
    .B(_1227_),
    .Y(_1229_)
);

NAND2X1 _2651_ (
    .A(_1229_),
    .B(_1228_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [7])
);

OR2X2 _2652_ (
    .A(_1023_),
    .B(_1048_),
    .Y(_1230_)
);

NAND2X1 _2653_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_1176_),
    .Y(_1231_)
);

INVX1 _2654_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [5]),
    .Y(_1232_)
);

NAND2X1 _2655_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6]),
    .Y(_1233_)
);

OAI21X1 _2656_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(_1232_),
    .C(_1233_),
    .Y(_1234_)
);

NAND2X1 _2657_ (
    .A(_1022__bF$buf1),
    .B(_1234_),
    .Y(_1235_)
);

NAND3X1 _2658_ (
    .A(_1052__bF$buf0),
    .B(_1231_),
    .C(_1235_),
    .Y(_1236_)
);

NAND3X1 _2659_ (
    .A(_1087__bF$buf4),
    .B(_1117_),
    .C(_1120_),
    .Y(_1237_)
);

NAND3X1 _2660_ (
    .A(_1064__bF$buf5),
    .B(_1236_),
    .C(_1237_),
    .Y(_1238_)
);

OAI21X1 _2661_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .B(_1230_),
    .C(_1238_),
    .Y(_1239_)
);

NAND3X1 _2662_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [7]),
    .B(_1046__bF$buf1),
    .C(_1239_),
    .Y(_1240_)
);

INVX1 _2663_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [7]),
    .Y(_1241_)
);

NAND3X1 _2664_ (
    .A(_1087__bF$buf3),
    .B(_1106_),
    .C(_1108_),
    .Y(_1242_)
);

MUX2X1 _2665_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [5]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .Y(_1243_)
);

NAND2X1 _2666_ (
    .A(_1022__bF$buf0),
    .B(_1243_),
    .Y(_1244_)
);

NAND2X1 _2667_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .B(_1166_),
    .Y(_1245_)
);

NAND3X1 _2668_ (
    .A(_1052__bF$buf5),
    .B(_1244_),
    .C(_1245_),
    .Y(_1246_)
);

NAND3X1 _2669_ (
    .A(_1064__bF$buf4),
    .B(_1242_),
    .C(_1246_),
    .Y(_1247_)
);

OAI21X1 _2670_ (
    .A(_1048_),
    .B(_1023_),
    .C(_1050__bF$buf5),
    .Y(_1248_)
);

NAND2X1 _2671_ (
    .A(_1248_),
    .B(_1247_),
    .Y(_1249_)
);

OAI21X1 _2672_ (
    .A(_1063__bF$buf2),
    .B(_1249_),
    .C(_1241_),
    .Y(_1250_)
);

NAND2X1 _2673_ (
    .A(_1240_),
    .B(_1250_),
    .Y(_1251_)
);

AOI21X1 _2674_ (
    .A(_1205_),
    .B(_1046__bF$buf0),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [6]),
    .Y(_1252_)
);

OAI21X1 _2675_ (
    .A(_1063__bF$buf1),
    .B(_1215_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [6]),
    .Y(_1253_)
);

NAND3X1 _2676_ (
    .A(_1207_),
    .B(_1046__bF$buf7),
    .C(_1205_),
    .Y(_1254_)
);

NAND2X1 _2677_ (
    .A(_1253_),
    .B(_1254_),
    .Y(_1255_)
);

NOR2X1 _2678_ (
    .A(_1199_),
    .B(_1255_),
    .Y(_1256_)
);

NAND2X1 _2679_ (
    .A(_1159_),
    .B(_1142_),
    .Y(_1257_)
);

NAND2X1 _2680_ (
    .A(_1150_),
    .B(_1257_),
    .Y(_1258_)
);

NAND3X1 _2681_ (
    .A(_1197_),
    .B(_1198_),
    .C(_1217_),
    .Y(_1259_)
);

INVX1 _2682_ (
    .A(_1253_),
    .Y(_1260_)
);

AOI21X1 _2683_ (
    .A(_1172_),
    .B(_1254_),
    .C(_1260_),
    .Y(_1261_)
);

OAI21X1 _2684_ (
    .A(_1258_),
    .B(_1259_),
    .C(_1261_),
    .Y(_1262_)
);

AOI21X1 _2685_ (
    .A(_1192_),
    .B(_1256_),
    .C(_1262_),
    .Y(_1263_)
);

NAND2X1 _2686_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .B(_1206_),
    .Y(_1264_)
);

OAI21X1 _2687_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .B(_1263_),
    .C(_1264_),
    .Y(_1265_)
);

OAI21X1 _2688_ (
    .A(_1252_),
    .B(_1224_),
    .C(_1265_),
    .Y(_1266_)
);

OR2X2 _2689_ (
    .A(_1266_),
    .B(_1251_),
    .Y(_1267_)
);

NAND3X1 _2690_ (
    .A(_1046__bF$buf6),
    .B(_1248_),
    .C(_1247_),
    .Y(_1268_)
);

NOR2X1 _2691_ (
    .A(_1241_),
    .B(_1268_),
    .Y(_1269_)
);

AND2X2 _2692_ (
    .A(_1268_),
    .B(_1241_),
    .Y(_1270_)
);

OAI21X1 _2693_ (
    .A(_1269_),
    .B(_1270_),
    .C(_1266_),
    .Y(_1271_)
);

NAND2X1 _2694_ (
    .A(_1271_),
    .B(_1267_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [8])
);

NAND2X1 _2695_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .B(_1031_),
    .Y(_1272_)
);

NAND2X1 _2696_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(_1211_),
    .Y(_1273_)
);

INVX1 _2697_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6]),
    .Y(_1274_)
);

NAND2X1 _2698_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [7]),
    .Y(_1275_)
);

OAI21X1 _2699_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(_1274_),
    .C(_1275_),
    .Y(_1276_)
);

NAND2X1 _2700_ (
    .A(_1022__bF$buf6),
    .B(_1276_),
    .Y(_1277_)
);

NAND3X1 _2701_ (
    .A(_1052__bF$buf4),
    .B(_1273_),
    .C(_1277_),
    .Y(_1278_)
);

NAND3X1 _2702_ (
    .A(_1087__bF$buf2),
    .B(_1138_),
    .C(_1135_),
    .Y(_1279_)
);

NAND3X1 _2703_ (
    .A(_1064__bF$buf3),
    .B(_1278_),
    .C(_1279_),
    .Y(_1280_)
);

OAI21X1 _2704_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .B(_1272_),
    .C(_1280_),
    .Y(_1281_)
);

NAND3X1 _2705_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [8]),
    .B(_1046__bF$buf5),
    .C(_1281_),
    .Y(_1282_)
);

INVX1 _2706_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [8]),
    .Y(_1283_)
);

NAND2X1 _2707_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6]),
    .B(_1034__bF$buf1),
    .Y(_1284_)
);

NAND3X1 _2708_ (
    .A(_1022__bF$buf5),
    .B(_1275_),
    .C(_1284_),
    .Y(_1285_)
);

NAND2X1 _2709_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .B(_1201_),
    .Y(_1286_)
);

NAND3X1 _2710_ (
    .A(_1052__bF$buf3),
    .B(_1285_),
    .C(_1286_),
    .Y(_1287_)
);

NAND3X1 _2711_ (
    .A(_1087__bF$buf1),
    .B(_1145_),
    .C(_1146_),
    .Y(_1288_)
);

NAND3X1 _2712_ (
    .A(_1064__bF$buf2),
    .B(_1287_),
    .C(_1288_),
    .Y(_1289_)
);

OAI21X1 _2713_ (
    .A(_1048_),
    .B(_1035_),
    .C(_1050__bF$buf4),
    .Y(_1290_)
);

NAND2X1 _2714_ (
    .A(_1290_),
    .B(_1289_),
    .Y(_1291_)
);

OAI21X1 _2715_ (
    .A(_1063__bF$buf0),
    .B(_1291_),
    .C(_1283_),
    .Y(_1292_)
);

NAND2X1 _2716_ (
    .A(_1292_),
    .B(_1282_),
    .Y(_1293_)
);

INVX1 _2717_ (
    .A(_1154_),
    .Y(_1294_)
);

OAI21X1 _2718_ (
    .A(_1126_),
    .B(_1294_),
    .C(_1125_),
    .Y(_1295_)
);

INVX1 _2719_ (
    .A(_1083_),
    .Y(_1296_)
);

INVX1 _2720_ (
    .A(_1112_),
    .Y(_1297_)
);

AOI21X1 _2721_ (
    .A(_1296_),
    .B(_1124_),
    .C(_1297_),
    .Y(_1298_)
);

OAI21X1 _2722_ (
    .A(_1130_),
    .B(_1295_),
    .C(_1298_),
    .Y(_1299_)
);

NAND3X1 _2723_ (
    .A(_1240_),
    .B(_1250_),
    .C(_1255_),
    .Y(_1300_)
);

NOR2X1 _2724_ (
    .A(_1300_),
    .B(_1222_),
    .Y(_1301_)
);

INVX1 _2725_ (
    .A(_1206_),
    .Y(_1302_)
);

AOI21X1 _2726_ (
    .A(_1302_),
    .B(_1250_),
    .C(_1269_),
    .Y(_1303_)
);

OAI21X1 _2727_ (
    .A(_1300_),
    .B(_1220_),
    .C(_1303_),
    .Y(_1304_)
);

AOI21X1 _2728_ (
    .A(_1299_),
    .B(_1301_),
    .C(_1304_),
    .Y(_1305_)
);

NAND2X1 _2729_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [7]),
    .B(_1268_),
    .Y(_1306_)
);

NAND3X1 _2730_ (
    .A(_1241_),
    .B(_1046__bF$buf4),
    .C(_1239_),
    .Y(_1307_)
);

NAND2X1 _2731_ (
    .A(_1306_),
    .B(_1307_),
    .Y(_1308_)
);

AND2X2 _2732_ (
    .A(_1268_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [7]),
    .Y(_1309_)
);

NOR2X1 _2733_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .B(_1309_),
    .Y(_1310_)
);

OAI21X1 _2734_ (
    .A(_1308_),
    .B(_1263_),
    .C(_1310_),
    .Y(_1311_)
);

OAI21X1 _2735_ (
    .A(_1027__bF$buf2),
    .B(_1305_),
    .C(_1311_),
    .Y(_1312_)
);

OR2X2 _2736_ (
    .A(_1312_),
    .B(_1293_),
    .Y(_1313_)
);

NAND3X1 _2737_ (
    .A(_1046__bF$buf3),
    .B(_1290_),
    .C(_1289_),
    .Y(_1314_)
);

NOR2X1 _2738_ (
    .A(_1283_),
    .B(_1314_),
    .Y(_1315_)
);

INVX1 _2739_ (
    .A(_1292_),
    .Y(_1316_)
);

OAI21X1 _2740_ (
    .A(_1315_),
    .B(_1316_),
    .C(_1312_),
    .Y(_1317_)
);

NAND2X1 _2741_ (
    .A(_1317_),
    .B(_1313_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [9])
);

MUX2X1 _2742_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [7]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .Y(_1318_)
);

NAND2X1 _2743_ (
    .A(_1022__bF$buf4),
    .B(_1318_),
    .Y(_1319_)
);

NAND2X1 _2744_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(_1243_),
    .Y(_1320_)
);

NAND3X1 _2745_ (
    .A(_1052__bF$buf2),
    .B(_1319_),
    .C(_1320_),
    .Y(_1321_)
);

MUX2X1 _2746_ (
    .A(_1166_),
    .B(_1107_),
    .S(_1022__bF$buf3),
    .Y(_1322_)
);

NAND2X1 _2747_ (
    .A(_1087__bF$buf0),
    .B(_1322_),
    .Y(_1323_)
);

NAND3X1 _2748_ (
    .A(_1064__bF$buf1),
    .B(_1321_),
    .C(_1323_),
    .Y(_1324_)
);

NAND2X1 _2749_ (
    .A(_1050__bF$buf3),
    .B(_1057_),
    .Y(_1325_)
);

NAND3X1 _2750_ (
    .A(_1046__bF$buf2),
    .B(_1325_),
    .C(_1324_),
    .Y(_1326_)
);

NAND2X1 _2751_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [9]),
    .B(_1326_),
    .Y(_1327_)
);

INVX1 _2752_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [9]),
    .Y(_1328_)
);

MUX2X1 _2753_ (
    .A(_1318_),
    .B(_1243_),
    .S(_1022__bF$buf2),
    .Y(_1329_)
);

MUX2X1 _2754_ (
    .A(_1322_),
    .B(_1329_),
    .S(_1087__bF$buf4),
    .Y(_1330_)
);

MUX2X1 _2755_ (
    .A(_1330_),
    .B(_1057_),
    .S(_1064__bF$buf0),
    .Y(_1331_)
);

NAND3X1 _2756_ (
    .A(_1328_),
    .B(_1046__bF$buf1),
    .C(_1331_),
    .Y(_1332_)
);

NAND2X1 _2757_ (
    .A(_1332_),
    .B(_1327_),
    .Y(_1333_)
);

INVX1 _2758_ (
    .A(_1333_),
    .Y(_1334_)
);

OAI21X1 _2759_ (
    .A(_1063__bF$buf4),
    .B(_1291_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [8]),
    .Y(_1335_)
);

NOR2X1 _2760_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [8]),
    .B(_1314_),
    .Y(_1336_)
);

OAI21X1 _2761_ (
    .A(_1306_),
    .B(_1336_),
    .C(_1335_),
    .Y(_1337_)
);

OAI21X1 _2762_ (
    .A(_1269_),
    .B(_1270_),
    .C(_1293_),
    .Y(_1338_)
);

NOR2X1 _2763_ (
    .A(_1338_),
    .B(_1263_),
    .Y(_1339_)
);

NOR2X1 _2764_ (
    .A(_1337_),
    .B(_1339_),
    .Y(_1340_)
);

NOR2X1 _2765_ (
    .A(_1027__bF$buf1),
    .B(_1315_),
    .Y(_1341_)
);

OAI21X1 _2766_ (
    .A(_1316_),
    .B(_1305_),
    .C(_1341_),
    .Y(_1342_)
);

OAI21X1 _2767_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .B(_1340_),
    .C(_1342_),
    .Y(_1343_)
);

OR2X2 _2768_ (
    .A(_1343_),
    .B(_1334_),
    .Y(_1344_)
);

NOR2X1 _2769_ (
    .A(_1328_),
    .B(_1326_),
    .Y(_1345_)
);

AOI21X1 _2770_ (
    .A(_1331_),
    .B(_1046__bF$buf0),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [9]),
    .Y(_1346_)
);

OAI21X1 _2771_ (
    .A(_1345_),
    .B(_1346_),
    .C(_1343_),
    .Y(_1347_)
);

AND2X2 _2772_ (
    .A(_1344_),
    .B(_1347_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [10])
);

MUX2X1 _2773_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [7]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .Y(_1348_)
);

MUX2X1 _2774_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [9]),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8]),
    .S(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .Y(_1349_)
);

MUX2X1 _2775_ (
    .A(_1349_),
    .B(_1348_),
    .S(_1022__bF$buf1),
    .Y(_1350_)
);

MUX2X1 _2776_ (
    .A(_1202_),
    .B(_1350_),
    .S(_1087__bF$buf3),
    .Y(_1351_)
);

MUX2X1 _2777_ (
    .A(_1351_),
    .B(_1081_),
    .S(_1064__bF$buf5),
    .Y(_1352_)
);

NAND3X1 _2778_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [10]),
    .B(_1046__bF$buf7),
    .C(_1352_),
    .Y(_1353_)
);

INVX1 _2779_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [10]),
    .Y(_1354_)
);

NAND2X1 _2780_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [9]),
    .Y(_1355_)
);

NAND2X1 _2781_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8]),
    .B(_1034__bF$buf0),
    .Y(_1356_)
);

NAND3X1 _2782_ (
    .A(_1022__bF$buf0),
    .B(_1355_),
    .C(_1356_),
    .Y(_1357_)
);

NAND2X1 _2783_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_1348_),
    .Y(_1358_)
);

NAND3X1 _2784_ (
    .A(_1052__bF$buf1),
    .B(_1357_),
    .C(_1358_),
    .Y(_1359_)
);

NAND2X1 _2785_ (
    .A(_1022__bF$buf6),
    .B(_1201_),
    .Y(_1360_)
);

NAND2X1 _2786_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_1144_),
    .Y(_1361_)
);

NAND3X1 _2787_ (
    .A(_1087__bF$buf2),
    .B(_1360_),
    .C(_1361_),
    .Y(_1362_)
);

NAND3X1 _2788_ (
    .A(_1064__bF$buf4),
    .B(_1359_),
    .C(_1362_),
    .Y(_1363_)
);

NAND2X1 _2789_ (
    .A(_1050__bF$buf2),
    .B(_1081_),
    .Y(_1364_)
);

NAND3X1 _2790_ (
    .A(_1046__bF$buf6),
    .B(_1364_),
    .C(_1363_),
    .Y(_1365_)
);

NAND2X1 _2791_ (
    .A(_1354_),
    .B(_1365_),
    .Y(_1366_)
);

NAND2X1 _2792_ (
    .A(_1366_),
    .B(_1353_),
    .Y(_1367_)
);

INVX1 _2793_ (
    .A(_1367_),
    .Y(_1368_)
);

NAND3X1 _2794_ (
    .A(_1283_),
    .B(_1046__bF$buf5),
    .C(_1281_),
    .Y(_1369_)
);

AOI22X1 _2795_ (
    .A(_1327_),
    .B(_1332_),
    .C(_1335_),
    .D(_1369_),
    .Y(_1370_)
);

INVX1 _2796_ (
    .A(_1370_),
    .Y(_1371_)
);

NAND2X1 _2797_ (
    .A(_1328_),
    .B(_1326_),
    .Y(_1372_)
);

AOI21X1 _2798_ (
    .A(_1315_),
    .B(_1372_),
    .C(_1345_),
    .Y(_1373_)
);

OAI21X1 _2799_ (
    .A(_1371_),
    .B(_1305_),
    .C(_1373_),
    .Y(_1374_)
);

INVX1 _2800_ (
    .A(_1374_),
    .Y(_1375_)
);

AOI21X1 _2801_ (
    .A(_1331_),
    .B(_1046__bF$buf4),
    .C(_1328_),
    .Y(_1376_)
);

NOR2X1 _2802_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .B(_1376_),
    .Y(_1377_)
);

OAI21X1 _2803_ (
    .A(_1333_),
    .B(_1340_),
    .C(_1377_),
    .Y(_1378_)
);

OAI21X1 _2804_ (
    .A(_1027__bF$buf0),
    .B(_1375_),
    .C(_1378_),
    .Y(_1379_)
);

OR2X2 _2805_ (
    .A(_1379_),
    .B(_1368_),
    .Y(_1380_)
);

AOI21X1 _2806_ (
    .A(_1352_),
    .B(_1046__bF$buf3),
    .C(_1354_),
    .Y(_1381_)
);

NOR2X1 _2807_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [10]),
    .B(_1365_),
    .Y(_1382_)
);

OAI21X1 _2808_ (
    .A(_1381_),
    .B(_1382_),
    .C(_1379_),
    .Y(_1383_)
);

AND2X2 _2809_ (
    .A(_1380_),
    .B(_1383_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [11])
);

NAND2X1 _2810_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [10]),
    .Y(_1384_)
);

NAND2X1 _2811_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [9]),
    .B(_1034__bF$buf3),
    .Y(_1385_)
);

NAND3X1 _2812_ (
    .A(_1022__bF$buf5),
    .B(_1384_),
    .C(_1385_),
    .Y(_1386_)
);

NAND2X1 _2813_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .B(_1318_),
    .Y(_1387_)
);

NAND3X1 _2814_ (
    .A(_1052__bF$buf0),
    .B(_1386_),
    .C(_1387_),
    .Y(_1388_)
);

NAND3X1 _2815_ (
    .A(_1087__bF$buf1),
    .B(_1244_),
    .C(_1245_),
    .Y(_1389_)
);

NAND3X1 _2816_ (
    .A(_1064__bF$buf3),
    .B(_1388_),
    .C(_1389_),
    .Y(_1390_)
);

NAND3X1 _2817_ (
    .A(_1050__bF$buf1),
    .B(_1110_),
    .C(_1109_),
    .Y(_1391_)
);

NAND3X1 _2818_ (
    .A(_1046__bF$buf2),
    .B(_1391_),
    .C(_1390_),
    .Y(_1392_)
);

NAND2X1 _2819_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [11]),
    .B(_1392_),
    .Y(_1393_)
);

INVX1 _2820_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [11]),
    .Y(_1394_)
);

NAND3X1 _2821_ (
    .A(_1050__bF$buf0),
    .B(_1122_),
    .C(_1121_),
    .Y(_1395_)
);

INVX1 _2822_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [7]),
    .Y(_1396_)
);

NAND2X1 _2823_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8]),
    .Y(_1397_)
);

OAI21X1 _2824_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_1396_),
    .C(_1397_),
    .Y(_1398_)
);

NAND2X1 _2825_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(_1398_),
    .Y(_1399_)
);

INVX1 _2826_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [9]),
    .Y(_1400_)
);

OAI21X1 _2827_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(_1400_),
    .C(_1384_),
    .Y(_1401_)
);

NAND2X1 _2828_ (
    .A(_1022__bF$buf4),
    .B(_1401_),
    .Y(_1402_)
);

NAND3X1 _2829_ (
    .A(_1052__bF$buf5),
    .B(_1399_),
    .C(_1402_),
    .Y(_1403_)
);

NAND3X1 _2830_ (
    .A(_1087__bF$buf0),
    .B(_1231_),
    .C(_1235_),
    .Y(_1404_)
);

NAND3X1 _2831_ (
    .A(_1064__bF$buf2),
    .B(_1403_),
    .C(_1404_),
    .Y(_1405_)
);

NAND2X1 _2832_ (
    .A(_1395_),
    .B(_1405_),
    .Y(_1406_)
);

NAND3X1 _2833_ (
    .A(_1394_),
    .B(_1046__bF$buf1),
    .C(_1406_),
    .Y(_1407_)
);

NAND3X1 _2834_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [9]),
    .B(_1046__bF$buf0),
    .C(_1331_),
    .Y(_1408_)
);

AOI22X1 _2835_ (
    .A(_1353_),
    .B(_1366_),
    .C(_1372_),
    .D(_1408_),
    .Y(_1409_)
);

NAND3X1 _2836_ (
    .A(_1251_),
    .B(_1293_),
    .C(_1409_),
    .Y(_1410_)
);

NAND2X1 _2837_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [10]),
    .B(_1365_),
    .Y(_1411_)
);

OAI21X1 _2838_ (
    .A(_1327_),
    .B(_1382_),
    .C(_1411_),
    .Y(_1412_)
);

AOI21X1 _2839_ (
    .A(_1337_),
    .B(_1409_),
    .C(_1412_),
    .Y(_1413_)
);

OAI21X1 _2840_ (
    .A(_1410_),
    .B(_1263_),
    .C(_1413_),
    .Y(_1414_)
);

NOR2X1 _2841_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .B(_1414_),
    .Y(_1415_)
);

INVX1 _2842_ (
    .A(_1365_),
    .Y(_1416_)
);

OAI21X1 _2843_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [10]),
    .B(_1416_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .Y(_1417_)
);

AOI21X1 _2844_ (
    .A(_1375_),
    .B(_1353_),
    .C(_1417_),
    .Y(_1418_)
);

NOR2X1 _2845_ (
    .A(_1415_),
    .B(_1418_),
    .Y(_1419_)
);

NAND3X1 _2846_ (
    .A(_1393_),
    .B(_1407_),
    .C(_1419_),
    .Y(_1420_)
);

NAND2X1 _2847_ (
    .A(_1393_),
    .B(_1407_),
    .Y(_1421_)
);

OAI21X1 _2848_ (
    .A(_1415_),
    .B(_1418_),
    .C(_1421_),
    .Y(_1422_)
);

AND2X2 _2849_ (
    .A(_1420_),
    .B(_1422_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [12])
);

NAND3X1 _2850_ (
    .A(_1050__bF$buf5),
    .B(_1140_),
    .C(_1139_),
    .Y(_1423_)
);

INVX1 _2851_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8]),
    .Y(_1424_)
);

OAI21X1 _2852_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .B(_1424_),
    .C(_1355_),
    .Y(_1425_)
);

NAND2X1 _2853_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .B(_1425_),
    .Y(_1426_)
);

INVX1 _2854_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [10]),
    .Y(_1427_)
);

NAND2X1 _2855_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [11]),
    .Y(_1428_)
);

OAI21X1 _2856_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(_1427_),
    .C(_1428_),
    .Y(_1429_)
);

NAND2X1 _2857_ (
    .A(_1022__bF$buf3),
    .B(_1429_),
    .Y(_1430_)
);

NAND3X1 _2858_ (
    .A(_1052__bF$buf4),
    .B(_1426_),
    .C(_1430_),
    .Y(_1431_)
);

NAND3X1 _2859_ (
    .A(_1087__bF$buf4),
    .B(_1273_),
    .C(_1277_),
    .Y(_1432_)
);

NAND3X1 _2860_ (
    .A(_1064__bF$buf1),
    .B(_1431_),
    .C(_1432_),
    .Y(_1433_)
);

NAND2X1 _2861_ (
    .A(_1423_),
    .B(_1433_),
    .Y(_1434_)
);

NAND3X1 _2862_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [12]),
    .B(_1046__bF$buf7),
    .C(_1434_),
    .Y(_1435_)
);

INVX1 _2863_ (
    .A(_1435_),
    .Y(_1436_)
);

INVX1 _2864_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [12]),
    .Y(_1437_)
);

NAND2X1 _2865_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [10]),
    .B(_1034__bF$buf2),
    .Y(_1438_)
);

NAND3X1 _2866_ (
    .A(_1022__bF$buf2),
    .B(_1428_),
    .C(_1438_),
    .Y(_1439_)
);

NAND2X1 _2867_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(_1349_),
    .Y(_1440_)
);

NAND3X1 _2868_ (
    .A(_1052__bF$buf3),
    .B(_1439_),
    .C(_1440_),
    .Y(_1441_)
);

NAND3X1 _2869_ (
    .A(_1087__bF$buf3),
    .B(_1285_),
    .C(_1286_),
    .Y(_1442_)
);

NAND3X1 _2870_ (
    .A(_1064__bF$buf0),
    .B(_1441_),
    .C(_1442_),
    .Y(_1443_)
);

NAND3X1 _2871_ (
    .A(_1050__bF$buf4),
    .B(_1148_),
    .C(_1147_),
    .Y(_1444_)
);

NAND3X1 _2872_ (
    .A(_1046__bF$buf6),
    .B(_1443_),
    .C(_1444_),
    .Y(_1445_)
);

NAND2X1 _2873_ (
    .A(_1437_),
    .B(_1445_),
    .Y(_1446_)
);

INVX1 _2874_ (
    .A(_1446_),
    .Y(_1447_)
);

NAND3X1 _2875_ (
    .A(_1354_),
    .B(_1046__bF$buf5),
    .C(_1352_),
    .Y(_1448_)
);

AOI22X1 _2876_ (
    .A(_1411_),
    .B(_1448_),
    .C(_1407_),
    .D(_1393_),
    .Y(_1449_)
);

NAND2X1 _2877_ (
    .A(_1449_),
    .B(_1370_),
    .Y(_1450_)
);

OAI21X1 _2878_ (
    .A(_1282_),
    .B(_1346_),
    .C(_1408_),
    .Y(_1451_)
);

NAND2X1 _2879_ (
    .A(_1394_),
    .B(_1392_),
    .Y(_1452_)
);

OAI21X1 _2880_ (
    .A(_1394_),
    .B(_1392_),
    .C(_1353_),
    .Y(_1453_)
);

AOI22X1 _2881_ (
    .A(_1452_),
    .B(_1453_),
    .C(_1451_),
    .D(_1449_),
    .Y(_1454_)
);

OAI21X1 _2882_ (
    .A(_1450_),
    .B(_1305_),
    .C(_1454_),
    .Y(_1455_)
);

NAND2X1 _2883_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .B(_1455_),
    .Y(_1456_)
);

INVX1 _2884_ (
    .A(_1414_),
    .Y(_1457_)
);

AOI21X1 _2885_ (
    .A(_1406_),
    .B(_1046__bF$buf4),
    .C(_1394_),
    .Y(_1458_)
);

NOR2X1 _2886_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .B(_1458_),
    .Y(_1459_)
);

OAI21X1 _2887_ (
    .A(_1421_),
    .B(_1457_),
    .C(_1459_),
    .Y(_1460_)
);

NAND2X1 _2888_ (
    .A(_1456_),
    .B(_1460_),
    .Y(_1461_)
);

INVX1 _2889_ (
    .A(_1461_),
    .Y(_1462_)
);

OAI21X1 _2890_ (
    .A(_1436_),
    .B(_1447_),
    .C(_1462_),
    .Y(_1463_)
);

AOI21X1 _2891_ (
    .A(_1434_),
    .B(_1046__bF$buf3),
    .C(_1437_),
    .Y(_1464_)
);

NOR2X1 _2892_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [12]),
    .B(_1445_),
    .Y(_1465_)
);

OAI21X1 _2893_ (
    .A(_1464_),
    .B(_1465_),
    .C(_1461_),
    .Y(_1466_)
);

AND2X2 _2894_ (
    .A(_1463_),
    .B(_1466_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [13])
);

OAI21X1 _2895_ (
    .A(_1087__bF$buf2),
    .B(_1322_),
    .C(_1181_),
    .Y(_1467_)
);

INVX1 _2896_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [11]),
    .Y(_1468_)
);

NAND2X1 _2897_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [12]),
    .Y(_1469_)
);

OAI21X1 _2898_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(_1468_),
    .C(_1469_),
    .Y(_1470_)
);

MUX2X1 _2899_ (
    .A(_1470_),
    .B(_1401_),
    .S(_1022__bF$buf1),
    .Y(_1471_)
);

NAND2X1 _2900_ (
    .A(_1052__bF$buf2),
    .B(_1471_),
    .Y(_1472_)
);

NAND2X1 _2901_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_1234_),
    .Y(_1473_)
);

NAND2X1 _2902_ (
    .A(_1022__bF$buf0),
    .B(_1398_),
    .Y(_1474_)
);

NAND3X1 _2903_ (
    .A(_1087__bF$buf1),
    .B(_1473_),
    .C(_1474_),
    .Y(_1475_)
);

NAND3X1 _2904_ (
    .A(_1064__bF$buf5),
    .B(_1475_),
    .C(_1472_),
    .Y(_1476_)
);

OAI21X1 _2905_ (
    .A(_1064__bF$buf4),
    .B(_1467_),
    .C(_1476_),
    .Y(_1477_)
);

NAND3X1 _2906_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [13]),
    .B(_1046__bF$buf2),
    .C(_1477_),
    .Y(_1478_)
);

INVX2 _2907_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [13]),
    .Y(_1479_)
);

NAND2X1 _2908_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [11]),
    .B(_1034__bF$buf1),
    .Y(_1480_)
);

NAND3X1 _2909_ (
    .A(_1022__bF$buf6),
    .B(_1469_),
    .C(_1480_),
    .Y(_1481_)
);

NAND3X1 _2910_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_1384_),
    .C(_1385_),
    .Y(_1482_)
);

NAND3X1 _2911_ (
    .A(_1052__bF$buf1),
    .B(_1481_),
    .C(_1482_),
    .Y(_1483_)
);

NAND2X1 _2912_ (
    .A(_1087__bF$buf0),
    .B(_1329_),
    .Y(_1484_)
);

NAND3X1 _2913_ (
    .A(_1064__bF$buf3),
    .B(_1483_),
    .C(_1484_),
    .Y(_1485_)
);

NAND3X1 _2914_ (
    .A(_1050__bF$buf3),
    .B(_1170_),
    .C(_1169_),
    .Y(_1486_)
);

NAND3X1 _2915_ (
    .A(_1046__bF$buf1),
    .B(_1486_),
    .C(_1485_),
    .Y(_1487_)
);

NAND2X1 _2916_ (
    .A(_1479_),
    .B(_1487_),
    .Y(_1488_)
);

NAND2X1 _2917_ (
    .A(_1488_),
    .B(_1478_),
    .Y(_1489_)
);

INVX1 _2918_ (
    .A(_1489_),
    .Y(_1490_)
);

NAND2X1 _2919_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [12]),
    .B(_1445_),
    .Y(_1491_)
);

OAI21X1 _2920_ (
    .A(_1393_),
    .B(_1465_),
    .C(_1491_),
    .Y(_1492_)
);

NAND3X1 _2921_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [11]),
    .B(_1046__bF$buf0),
    .C(_1406_),
    .Y(_1493_)
);

AOI22X1 _2922_ (
    .A(_1493_),
    .B(_1452_),
    .C(_1435_),
    .D(_1446_),
    .Y(_1494_)
);

AOI21X1 _2923_ (
    .A(_1414_),
    .B(_1494_),
    .C(_1492_),
    .Y(_1495_)
);

NAND2X1 _2924_ (
    .A(_1027__bF$buf5),
    .B(_1495_),
    .Y(_1496_)
);

NOR2X1 _2925_ (
    .A(_1027__bF$buf4),
    .B(_1447_),
    .Y(_1497_)
);

OAI21X1 _2926_ (
    .A(_1436_),
    .B(_1455_),
    .C(_1497_),
    .Y(_1498_)
);

NAND2X1 _2927_ (
    .A(_1498_),
    .B(_1496_),
    .Y(_1499_)
);

OR2X2 _2928_ (
    .A(_1499_),
    .B(_1490_),
    .Y(_1500_)
);

NAND2X1 _2929_ (
    .A(_1490_),
    .B(_1499_),
    .Y(_1501_)
);

AND2X2 _2930_ (
    .A(_1500_),
    .B(_1501_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [14])
);

NAND3X1 _2931_ (
    .A(_1050__bF$buf2),
    .B(_1213_),
    .C(_1214_),
    .Y(_1502_)
);

INVX1 _2932_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [12]),
    .Y(_1503_)
);

NAND2X1 _2933_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [13]),
    .Y(_1504_)
);

OAI21X1 _2934_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_1503_),
    .C(_1504_),
    .Y(_1505_)
);

MUX2X1 _2935_ (
    .A(_1505_),
    .B(_1429_),
    .S(_1022__bF$buf5),
    .Y(_1506_)
);

NAND2X1 _2936_ (
    .A(_1052__bF$buf0),
    .B(_1506_),
    .Y(_1507_)
);

NAND2X1 _2937_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .B(_1276_),
    .Y(_1508_)
);

NAND2X1 _2938_ (
    .A(_1022__bF$buf4),
    .B(_1425_),
    .Y(_1509_)
);

NAND3X1 _2939_ (
    .A(_1087__bF$buf4),
    .B(_1508_),
    .C(_1509_),
    .Y(_1510_)
);

NAND3X1 _2940_ (
    .A(_1064__bF$buf2),
    .B(_1510_),
    .C(_1507_),
    .Y(_1511_)
);

NAND2X1 _2941_ (
    .A(_1502_),
    .B(_1511_),
    .Y(_1512_)
);

NAND3X1 _2942_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [14]),
    .B(_1046__bF$buf7),
    .C(_1512_),
    .Y(_1513_)
);

INVX1 _2943_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [14]),
    .Y(_1514_)
);

NAND2X1 _2944_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [12]),
    .B(_1034__bF$buf0),
    .Y(_1515_)
);

NAND3X1 _2945_ (
    .A(_1022__bF$buf3),
    .B(_1504_),
    .C(_1515_),
    .Y(_1516_)
);

NAND3X1 _2946_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(_1428_),
    .C(_1438_),
    .Y(_1517_)
);

NAND3X1 _2947_ (
    .A(_1052__bF$buf5),
    .B(_1516_),
    .C(_1517_),
    .Y(_1518_)
);

NAND2X1 _2948_ (
    .A(_1087__bF$buf3),
    .B(_1350_),
    .Y(_1519_)
);

NAND3X1 _2949_ (
    .A(_1064__bF$buf1),
    .B(_1518_),
    .C(_1519_),
    .Y(_1520_)
);

NAND3X1 _2950_ (
    .A(_1050__bF$buf1),
    .B(_1204_),
    .C(_1203_),
    .Y(_1521_)
);

NAND3X1 _2951_ (
    .A(_1046__bF$buf6),
    .B(_1520_),
    .C(_1521_),
    .Y(_1522_)
);

NAND2X1 _2952_ (
    .A(_1514_),
    .B(_1522_),
    .Y(_1523_)
);

NAND2X1 _2953_ (
    .A(_1513_),
    .B(_1523_),
    .Y(_1524_)
);

INVX1 _2954_ (
    .A(_1524_),
    .Y(_1525_)
);

NAND3X1 _2955_ (
    .A(_1437_),
    .B(_1046__bF$buf5),
    .C(_1434_),
    .Y(_1526_)
);

NAND2X1 _2956_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [13]),
    .B(_1487_),
    .Y(_1527_)
);

NAND3X1 _2957_ (
    .A(_1479_),
    .B(_1046__bF$buf4),
    .C(_1477_),
    .Y(_1528_)
);

AOI22X1 _2958_ (
    .A(_1491_),
    .B(_1526_),
    .C(_1528_),
    .D(_1527_),
    .Y(_1529_)
);

AND2X2 _2959_ (
    .A(_1487_),
    .B(_1479_),
    .Y(_1530_)
);

OAI21X1 _2960_ (
    .A(_1435_),
    .B(_1530_),
    .C(_1478_),
    .Y(_1531_)
);

AOI21X1 _2961_ (
    .A(_1455_),
    .B(_1529_),
    .C(_1531_),
    .Y(_1532_)
);

INVX1 _2962_ (
    .A(_1487_),
    .Y(_1533_)
);

OAI21X1 _2963_ (
    .A(_1479_),
    .B(_1533_),
    .C(_1027__bF$buf3),
    .Y(_1534_)
);

INVX1 _2964_ (
    .A(_1534_),
    .Y(_1535_)
);

OAI21X1 _2965_ (
    .A(_1490_),
    .B(_1495_),
    .C(_1535_),
    .Y(_1536_)
);

OAI21X1 _2966_ (
    .A(_1027__bF$buf2),
    .B(_1532_),
    .C(_1536_),
    .Y(_1537_)
);

OR2X2 _2967_ (
    .A(_1537_),
    .B(_1525_),
    .Y(_1538_)
);

AOI21X1 _2968_ (
    .A(_1512_),
    .B(_1046__bF$buf3),
    .C(_1514_),
    .Y(_1539_)
);

NOR2X1 _2969_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [14]),
    .B(_1522_),
    .Y(_1540_)
);

OAI21X1 _2970_ (
    .A(_1539_),
    .B(_1540_),
    .C(_1537_),
    .Y(_1541_)
);

AND2X2 _2971_ (
    .A(_1538_),
    .B(_1541_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [15])
);

INVX1 _2972_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [15]),
    .Y(_1542_)
);

NAND2X1 _2973_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [14]),
    .Y(_1543_)
);

NAND2X1 _2974_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [13]),
    .B(_1034__bF$buf3),
    .Y(_1544_)
);

NAND3X1 _2975_ (
    .A(_1022__bF$buf2),
    .B(_1543_),
    .C(_1544_),
    .Y(_1545_)
);

NAND3X1 _2976_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .B(_1469_),
    .C(_1480_),
    .Y(_1546_)
);

NAND3X1 _2977_ (
    .A(_1052__bF$buf4),
    .B(_1545_),
    .C(_1546_),
    .Y(_1547_)
);

NAND3X1 _2978_ (
    .A(_1087__bF$buf2),
    .B(_1386_),
    .C(_1387_),
    .Y(_1548_)
);

NAND3X1 _2979_ (
    .A(_1064__bF$buf0),
    .B(_1547_),
    .C(_1548_),
    .Y(_1549_)
);

NAND3X1 _2980_ (
    .A(_1050__bF$buf0),
    .B(_1242_),
    .C(_1246_),
    .Y(_1550_)
);

NAND3X1 _2981_ (
    .A(_1046__bF$buf2),
    .B(_1549_),
    .C(_1550_),
    .Y(_1551_)
);

NAND2X1 _2982_ (
    .A(_1025_),
    .B(_1063__bF$buf3),
    .Y(_1552_)
);

AOI21X1 _2983_ (
    .A(_1551_),
    .B(_1552_),
    .C(_1542_),
    .Y(_1553_)
);

NAND2X1 _2984_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(_1470_),
    .Y(_1554_)
);

INVX1 _2985_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [13]),
    .Y(_1555_)
);

OAI21X1 _2986_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .B(_1555_),
    .C(_1543_),
    .Y(_1556_)
);

NAND2X1 _2987_ (
    .A(_1022__bF$buf1),
    .B(_1556_),
    .Y(_1557_)
);

NAND3X1 _2988_ (
    .A(_1052__bF$buf3),
    .B(_1554_),
    .C(_1557_),
    .Y(_1558_)
);

NAND3X1 _2989_ (
    .A(_1087__bF$buf1),
    .B(_1399_),
    .C(_1402_),
    .Y(_1559_)
);

NAND3X1 _2990_ (
    .A(_1064__bF$buf5),
    .B(_1558_),
    .C(_1559_),
    .Y(_1560_)
);

NAND3X1 _2991_ (
    .A(_1050__bF$buf5),
    .B(_1236_),
    .C(_1237_),
    .Y(_1561_)
);

NAND3X1 _2992_ (
    .A(_1046__bF$buf1),
    .B(_1560_),
    .C(_1561_),
    .Y(_1562_)
);

OAI21X1 _2993_ (
    .A(_1047_),
    .B(_1230_),
    .C(_1063__bF$buf2),
    .Y(_1563_)
);

AOI21X1 _2994_ (
    .A(_1562_),
    .B(_1563_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [15]),
    .Y(_1564_)
);

AOI22X1 _2995_ (
    .A(_1523_),
    .B(_1513_),
    .C(_1478_),
    .D(_1488_),
    .Y(_1565_)
);

NAND2X1 _2996_ (
    .A(_1494_),
    .B(_1565_),
    .Y(_1566_)
);

OR2X2 _2997_ (
    .A(_1566_),
    .B(_1410_),
    .Y(_1567_)
);

AND2X2 _2998_ (
    .A(_1314_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [8]),
    .Y(_1568_)
);

AOI21X1 _2999_ (
    .A(_1309_),
    .B(_1369_),
    .C(_1568_),
    .Y(_1569_)
);

OAI21X1 _3000_ (
    .A(_1345_),
    .B(_1346_),
    .C(_1367_),
    .Y(_1570_)
);

AOI21X1 _3001_ (
    .A(_1376_),
    .B(_1448_),
    .C(_1381_),
    .Y(_1571_)
);

OAI21X1 _3002_ (
    .A(_1569_),
    .B(_1570_),
    .C(_1571_),
    .Y(_1572_)
);

AND2X2 _3003_ (
    .A(_1565_),
    .B(_1494_),
    .Y(_1573_)
);

AOI21X1 _3004_ (
    .A(_1458_),
    .B(_1526_),
    .C(_1464_),
    .Y(_1574_)
);

NOR2X1 _3005_ (
    .A(_1479_),
    .B(_1487_),
    .Y(_1575_)
);

NOR2X1 _3006_ (
    .A(_1514_),
    .B(_1522_),
    .Y(_1576_)
);

AOI21X1 _3007_ (
    .A(_1512_),
    .B(_1046__bF$buf0),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [14]),
    .Y(_1577_)
);

OAI22X1 _3008_ (
    .A(_1575_),
    .B(_1530_),
    .C(_1577_),
    .D(_1576_),
    .Y(_1578_)
);

AND2X2 _3009_ (
    .A(_1487_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [13]),
    .Y(_1579_)
);

NAND3X1 _3010_ (
    .A(_1514_),
    .B(_1046__bF$buf7),
    .C(_1512_),
    .Y(_1580_)
);

AOI21X1 _3011_ (
    .A(_1579_),
    .B(_1580_),
    .C(_1539_),
    .Y(_1581_)
);

OAI21X1 _3012_ (
    .A(_1574_),
    .B(_1578_),
    .C(_1581_),
    .Y(_1582_)
);

AOI21X1 _3013_ (
    .A(_1572_),
    .B(_1573_),
    .C(_1582_),
    .Y(_1583_)
);

OAI21X1 _3014_ (
    .A(_1263_),
    .B(_1567_),
    .C(_1583_),
    .Y(_1584_)
);

NOR2X1 _3015_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .B(_1584_),
    .Y(_1585_)
);

NAND2X1 _3016_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .B(_1523_),
    .Y(_1586_)
);

AOI21X1 _3017_ (
    .A(_1532_),
    .B(_1513_),
    .C(_1586_),
    .Y(_1587_)
);

NOR2X1 _3018_ (
    .A(_1585_),
    .B(_1587_),
    .Y(_1588_)
);

OAI21X1 _3019_ (
    .A(_1553_),
    .B(_1564_),
    .C(_1588_),
    .Y(_1589_)
);

NAND3X1 _3020_ (
    .A(_1542_),
    .B(_1563_),
    .C(_1562_),
    .Y(_1590_)
);

NAND3X1 _3021_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [15]),
    .B(_1552_),
    .C(_1551_),
    .Y(_1591_)
);

NAND2X1 _3022_ (
    .A(_1591_),
    .B(_1590_),
    .Y(_1592_)
);

OAI21X1 _3023_ (
    .A(_1585_),
    .B(_1587_),
    .C(_1592_),
    .Y(_1593_)
);

AND2X2 _3024_ (
    .A(_1589_),
    .B(_1593_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [16])
);

INVX1 _3025_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [16]),
    .Y(_1594_)
);

NAND3X1 _3026_ (
    .A(_1050__bF$buf4),
    .B(_1278_),
    .C(_1279_),
    .Y(_1595_)
);

NAND2X1 _3027_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_1505_),
    .Y(_1596_)
);

INVX1 _3028_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [14]),
    .Y(_1597_)
);

NAND2X1 _3029_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [15]),
    .Y(_1598_)
);

OAI21X1 _3030_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(_1597_),
    .C(_1598_),
    .Y(_1599_)
);

NAND2X1 _3031_ (
    .A(_1022__bF$buf0),
    .B(_1599_),
    .Y(_1600_)
);

NAND3X1 _3032_ (
    .A(_1052__bF$buf2),
    .B(_1596_),
    .C(_1600_),
    .Y(_1601_)
);

OAI21X1 _3033_ (
    .A(_1022__bF$buf6),
    .B(_1425_),
    .C(_1439_),
    .Y(_1602_)
);

OAI21X1 _3034_ (
    .A(_1043_),
    .B(_1051_),
    .C(_1602_),
    .Y(_1603_)
);

NAND3X1 _3035_ (
    .A(_1064__bF$buf4),
    .B(_1601_),
    .C(_1603_),
    .Y(_1604_)
);

NAND3X1 _3036_ (
    .A(_1046__bF$buf6),
    .B(_1595_),
    .C(_1604_),
    .Y(_1605_)
);

OAI21X1 _3037_ (
    .A(_1047_),
    .B(_1272_),
    .C(_1063__bF$buf1),
    .Y(_1606_)
);

NAND3X1 _3038_ (
    .A(_1594_),
    .B(_1606_),
    .C(_1605_),
    .Y(_1607_)
);

NAND2X1 _3039_ (
    .A(_1596_),
    .B(_1600_),
    .Y(_1608_)
);

NAND2X1 _3040_ (
    .A(_1052__bF$buf1),
    .B(_1608_),
    .Y(_1609_)
);

NAND3X1 _3041_ (
    .A(_1087__bF$buf0),
    .B(_1439_),
    .C(_1440_),
    .Y(_1610_)
);

NAND3X1 _3042_ (
    .A(_1064__bF$buf3),
    .B(_1610_),
    .C(_1609_),
    .Y(_1611_)
);

NAND3X1 _3043_ (
    .A(_1050__bF$buf3),
    .B(_1287_),
    .C(_1288_),
    .Y(_1612_)
);

NAND3X1 _3044_ (
    .A(_1046__bF$buf5),
    .B(_1612_),
    .C(_1611_),
    .Y(_1613_)
);

NAND2X1 _3045_ (
    .A(_1036_),
    .B(_1063__bF$buf0),
    .Y(_1614_)
);

NAND3X1 _3046_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [16]),
    .B(_1614_),
    .C(_1613_),
    .Y(_1615_)
);

AOI21X1 _3047_ (
    .A(_1551_),
    .B(_1552_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [15]),
    .Y(_1616_)
);

NAND3X1 _3048_ (
    .A(_1155_),
    .B(_1152_),
    .C(_1256_),
    .Y(_1617_)
);

OAI21X1 _3049_ (
    .A(_1197_),
    .B(_1255_),
    .C(_1253_),
    .Y(_1618_)
);

AOI21X1 _3050_ (
    .A(_1256_),
    .B(_1193_),
    .C(_1618_),
    .Y(_1619_)
);

OAI21X1 _3051_ (
    .A(_1127_),
    .B(_1617_),
    .C(_1619_),
    .Y(_1620_)
);

NOR2X1 _3052_ (
    .A(_1410_),
    .B(_1566_),
    .Y(_1621_)
);

NAND2X1 _3053_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [14]),
    .B(_1522_),
    .Y(_1622_)
);

OAI21X1 _3054_ (
    .A(_1527_),
    .B(_1540_),
    .C(_1622_),
    .Y(_1623_)
);

AOI21X1 _3055_ (
    .A(_1492_),
    .B(_1565_),
    .C(_1623_),
    .Y(_1624_)
);

OAI21X1 _3056_ (
    .A(_1566_),
    .B(_1413_),
    .C(_1624_),
    .Y(_1625_)
);

AOI21X1 _3057_ (
    .A(_1620_),
    .B(_1621_),
    .C(_1625_),
    .Y(_1626_)
);

OAI21X1 _3058_ (
    .A(_1616_),
    .B(_1626_),
    .C(_1591_),
    .Y(_1627_)
);

NAND2X1 _3059_ (
    .A(_1027__bF$buf1),
    .B(_1627_),
    .Y(_1628_)
);

NAND2X1 _3060_ (
    .A(_1452_),
    .B(_1453_),
    .Y(_1629_)
);

NOR2X1 _3061_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [11]),
    .B(_1392_),
    .Y(_1630_)
);

OAI22X1 _3062_ (
    .A(_1381_),
    .B(_1382_),
    .C(_1630_),
    .D(_1458_),
    .Y(_1631_)
);

OAI21X1 _3063_ (
    .A(_1631_),
    .B(_1373_),
    .C(_1629_),
    .Y(_1632_)
);

AOI22X1 _3064_ (
    .A(_1622_),
    .B(_1580_),
    .C(_1590_),
    .D(_1591_),
    .Y(_1633_)
);

AND2X2 _3065_ (
    .A(_1633_),
    .B(_1529_),
    .Y(_1634_)
);

OAI22X1 _3066_ (
    .A(_1437_),
    .B(_1445_),
    .C(_1479_),
    .D(_1487_),
    .Y(_1635_)
);

OAI21X1 _3067_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [13]),
    .B(_1533_),
    .C(_1635_),
    .Y(_1636_)
);

AOI21X1 _3068_ (
    .A(_1562_),
    .B(_1563_),
    .C(_1542_),
    .Y(_1637_)
);

OAI22X1 _3069_ (
    .A(_1539_),
    .B(_1540_),
    .C(_1616_),
    .D(_1637_),
    .Y(_1638_)
);

NAND3X1 _3070_ (
    .A(_1542_),
    .B(_1552_),
    .C(_1551_),
    .Y(_1639_)
);

AOI21X1 _3071_ (
    .A(_1576_),
    .B(_1639_),
    .C(_1553_),
    .Y(_1640_)
);

OAI21X1 _3072_ (
    .A(_1636_),
    .B(_1638_),
    .C(_1640_),
    .Y(_1641_)
);

AOI21X1 _3073_ (
    .A(_1632_),
    .B(_1634_),
    .C(_1641_),
    .Y(_1642_)
);

NAND2X1 _3074_ (
    .A(_1529_),
    .B(_1633_),
    .Y(_1643_)
);

OR2X2 _3075_ (
    .A(_1643_),
    .B(_1450_),
    .Y(_1644_)
);

OAI21X1 _3076_ (
    .A(_1644_),
    .B(_1305_),
    .C(_1642_),
    .Y(_1645_)
);

OAI21X1 _3077_ (
    .A(_1027__bF$buf0),
    .B(_1645_),
    .C(_1628_),
    .Y(_1646_)
);

NAND3X1 _3078_ (
    .A(_1607_),
    .B(_1615_),
    .C(_1646_),
    .Y(_1647_)
);

AOI21X1 _3079_ (
    .A(_1613_),
    .B(_1614_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [16]),
    .Y(_1648_)
);

INVX1 _3080_ (
    .A(_1615_),
    .Y(_1649_)
);

INVX1 _3081_ (
    .A(_1646_),
    .Y(_1650_)
);

OAI21X1 _3082_ (
    .A(_1648_),
    .B(_1649_),
    .C(_1650_),
    .Y(_1651_)
);

AND2X2 _3083_ (
    .A(_1651_),
    .B(_1647_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [17])
);

NAND2X1 _3084_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_1556_),
    .Y(_1652_)
);

INVX1 _3085_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [15]),
    .Y(_1653_)
);

NAND2X1 _3086_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [16]),
    .Y(_1654_)
);

OAI21X1 _3087_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(_1653_),
    .C(_1654_),
    .Y(_1655_)
);

NAND2X1 _3088_ (
    .A(_1022__bF$buf5),
    .B(_1655_),
    .Y(_1656_)
);

NAND3X1 _3089_ (
    .A(_1052__bF$buf0),
    .B(_1652_),
    .C(_1656_),
    .Y(_1657_)
);

NAND2X1 _3090_ (
    .A(_1087__bF$buf4),
    .B(_1471_),
    .Y(_1658_)
);

NAND3X1 _3091_ (
    .A(_1064__bF$buf2),
    .B(_1657_),
    .C(_1658_),
    .Y(_1659_)
);

NAND2X1 _3092_ (
    .A(_1321_),
    .B(_1323_),
    .Y(_1660_)
);

NAND2X1 _3093_ (
    .A(_1050__bF$buf2),
    .B(_1660_),
    .Y(_1661_)
);

NAND3X1 _3094_ (
    .A(_1046__bF$buf4),
    .B(_1659_),
    .C(_1661_),
    .Y(_1662_)
);

OAI21X1 _3095_ (
    .A(_1050__bF$buf1),
    .B(_1057_),
    .C(_1063__bF$buf4),
    .Y(_1663_)
);

NAND3X1 _3096_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [17]),
    .B(_1663_),
    .C(_1662_),
    .Y(_1664_)
);

INVX1 _3097_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [17]),
    .Y(_1665_)
);

OAI21X1 _3098_ (
    .A(_1064__bF$buf1),
    .B(_1330_),
    .C(_1659_),
    .Y(_1666_)
);

NAND2X1 _3099_ (
    .A(_1046__bF$buf3),
    .B(_1666_),
    .Y(_1667_)
);

NAND2X1 _3100_ (
    .A(_1063__bF$buf3),
    .B(_1058_),
    .Y(_1668_)
);

NAND3X1 _3101_ (
    .A(_1665_),
    .B(_1668_),
    .C(_1667_),
    .Y(_1669_)
);

NAND2X1 _3102_ (
    .A(_1664_),
    .B(_1669_),
    .Y(_1670_)
);

INVX1 _3103_ (
    .A(_1670_),
    .Y(_1671_)
);

AOI21X1 _3104_ (
    .A(_1637_),
    .B(_1607_),
    .C(_1649_),
    .Y(_1672_)
);

NAND3X1 _3105_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [16]),
    .B(_1606_),
    .C(_1605_),
    .Y(_1673_)
);

NAND3X1 _3106_ (
    .A(_1594_),
    .B(_1614_),
    .C(_1613_),
    .Y(_1674_)
);

AOI21X1 _3107_ (
    .A(_1673_),
    .B(_1674_),
    .C(_1592_),
    .Y(_1675_)
);

NAND2X1 _3108_ (
    .A(_1675_),
    .B(_1584_),
    .Y(_1676_)
);

NAND2X1 _3109_ (
    .A(_1672_),
    .B(_1676_),
    .Y(_1677_)
);

NAND2X1 _3110_ (
    .A(_1027__bF$buf5),
    .B(_1677_),
    .Y(_1678_)
);

NAND2X1 _3111_ (
    .A(_1674_),
    .B(_1645_),
    .Y(_1679_)
);

NAND3X1 _3112_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .B(_1673_),
    .C(_1679_),
    .Y(_1680_)
);

NAND3X1 _3113_ (
    .A(_1671_),
    .B(_1680_),
    .C(_1678_),
    .Y(_1681_)
);

NAND2X1 _3114_ (
    .A(_1680_),
    .B(_1678_),
    .Y(_1682_)
);

NAND2X1 _3115_ (
    .A(_1670_),
    .B(_1682_),
    .Y(_1683_)
);

AND2X2 _3116_ (
    .A(_1683_),
    .B(_1681_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [18])
);

NAND2X1 _3117_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .B(_1599_),
    .Y(_1684_)
);

INVX1 _3118_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [16]),
    .Y(_1685_)
);

NAND2X1 _3119_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [17]),
    .Y(_1686_)
);

OAI21X1 _3120_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_1685_),
    .C(_1686_),
    .Y(_1687_)
);

NAND2X1 _3121_ (
    .A(_1022__bF$buf4),
    .B(_1687_),
    .Y(_1688_)
);

NAND3X1 _3122_ (
    .A(_1052__bF$buf5),
    .B(_1684_),
    .C(_1688_),
    .Y(_1689_)
);

OAI21X1 _3123_ (
    .A(_1043_),
    .B(_1051_),
    .C(_1506_),
    .Y(_1690_)
);

NAND3X1 _3124_ (
    .A(_1064__bF$buf0),
    .B(_1689_),
    .C(_1690_),
    .Y(_1691_)
);

NAND2X1 _3125_ (
    .A(_1359_),
    .B(_1362_),
    .Y(_1692_)
);

AOI21X1 _3126_ (
    .A(_1692_),
    .B(_1050__bF$buf0),
    .C(_1063__bF$buf2),
    .Y(_1693_)
);

NAND2X1 _3127_ (
    .A(_1691_),
    .B(_1693_),
    .Y(_1694_)
);

OAI21X1 _3128_ (
    .A(_1050__bF$buf5),
    .B(_1081_),
    .C(_1063__bF$buf1),
    .Y(_1695_)
);

NAND3X1 _3129_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [18]),
    .B(_1695_),
    .C(_1694_),
    .Y(_1696_)
);

INVX1 _3130_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [18]),
    .Y(_1697_)
);

INVX1 _3131_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [17]),
    .Y(_1698_)
);

NAND2X1 _3132_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(_1698_),
    .Y(_1699_)
);

OAI21X1 _3133_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [16]),
    .C(_1699_),
    .Y(_1700_)
);

OAI21X1 _3134_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(_1700_),
    .C(_1684_),
    .Y(_1701_)
);

NAND2X1 _3135_ (
    .A(_1052__bF$buf4),
    .B(_1701_),
    .Y(_1702_)
);

OR2X2 _3136_ (
    .A(_1506_),
    .B(_1052__bF$buf3),
    .Y(_1703_)
);

NAND3X1 _3137_ (
    .A(_1064__bF$buf5),
    .B(_1702_),
    .C(_1703_),
    .Y(_1704_)
);

NAND2X1 _3138_ (
    .A(_1050__bF$buf4),
    .B(_1351_),
    .Y(_1705_)
);

NAND3X1 _3139_ (
    .A(_1046__bF$buf2),
    .B(_1705_),
    .C(_1704_),
    .Y(_1706_)
);

NAND2X1 _3140_ (
    .A(_1063__bF$buf0),
    .B(_1082_),
    .Y(_1707_)
);

NAND3X1 _3141_ (
    .A(_1697_),
    .B(_1707_),
    .C(_1706_),
    .Y(_1708_)
);

NAND2X1 _3142_ (
    .A(_1708_),
    .B(_1696_),
    .Y(_1709_)
);

NAND3X1 _3143_ (
    .A(_1255_),
    .B(_1221_),
    .C(_1308_),
    .Y(_1710_)
);

OR2X2 _3144_ (
    .A(_1218_),
    .B(_1165_),
    .Y(_1711_)
);

OAI21X1 _3145_ (
    .A(_1172_),
    .B(_1183_),
    .C(_1184_),
    .Y(_1712_)
);

NAND2X1 _3146_ (
    .A(_1711_),
    .B(_1712_),
    .Y(_1713_)
);

AOI21X1 _3147_ (
    .A(_1306_),
    .B(_1307_),
    .C(_1217_),
    .Y(_1714_)
);

OAI21X1 _3148_ (
    .A(_1206_),
    .B(_1270_),
    .C(_1240_),
    .Y(_1715_)
);

AOI21X1 _3149_ (
    .A(_1713_),
    .B(_1714_),
    .C(_1715_),
    .Y(_1716_)
);

OAI21X1 _3150_ (
    .A(_1158_),
    .B(_1710_),
    .C(_1716_),
    .Y(_1717_)
);

NAND3X1 _3151_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [15]),
    .B(_1563_),
    .C(_1562_),
    .Y(_1718_)
);

OAI21X1 _3152_ (
    .A(_1513_),
    .B(_1564_),
    .C(_1718_),
    .Y(_1719_)
);

AOI21X1 _3153_ (
    .A(_1531_),
    .B(_1633_),
    .C(_1719_),
    .Y(_1720_)
);

OAI21X1 _3154_ (
    .A(_1454_),
    .B(_1643_),
    .C(_1720_),
    .Y(_1721_)
);

NOR2X1 _3155_ (
    .A(_1450_),
    .B(_1643_),
    .Y(_1722_)
);

AOI21X1 _3156_ (
    .A(_1717_),
    .B(_1722_),
    .C(_1721_),
    .Y(_1723_)
);

NAND3X1 _3157_ (
    .A(_1665_),
    .B(_1663_),
    .C(_1662_),
    .Y(_1724_)
);

NAND3X1 _3158_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [17]),
    .B(_1668_),
    .C(_1667_),
    .Y(_1725_)
);

AOI22X1 _3159_ (
    .A(_1607_),
    .B(_1615_),
    .C(_1725_),
    .D(_1724_),
    .Y(_1726_)
);

INVX1 _3160_ (
    .A(_1726_),
    .Y(_1727_)
);

AOI21X1 _3161_ (
    .A(_1662_),
    .B(_1663_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [17]),
    .Y(_1728_)
);

OAI21X1 _3162_ (
    .A(_1673_),
    .B(_1728_),
    .C(_1664_),
    .Y(_1729_)
);

INVX1 _3163_ (
    .A(_1729_),
    .Y(_1730_)
);

OAI21X1 _3164_ (
    .A(_1727_),
    .B(_1723_),
    .C(_1730_),
    .Y(_1731_)
);

NAND2X1 _3165_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .B(_1731_),
    .Y(_1732_)
);

NAND2X1 _3166_ (
    .A(_1027__bF$buf4),
    .B(_1725_),
    .Y(_1733_)
);

AOI21X1 _3167_ (
    .A(_1677_),
    .B(_1670_),
    .C(_1733_),
    .Y(_1734_)
);

INVX1 _3168_ (
    .A(_1734_),
    .Y(_1735_)
);

NAND3X1 _3169_ (
    .A(_1709_),
    .B(_1732_),
    .C(_1735_),
    .Y(_1736_)
);

INVX1 _3170_ (
    .A(_1709_),
    .Y(_1737_)
);

INVX1 _3171_ (
    .A(_1732_),
    .Y(_1738_)
);

OAI21X1 _3172_ (
    .A(_1738_),
    .B(_1734_),
    .C(_1737_),
    .Y(_1739_)
);

AND2X2 _3173_ (
    .A(_1736_),
    .B(_1739_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [19])
);

INVX1 _3174_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [19]),
    .Y(_1740_)
);

NAND2X1 _3175_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .B(_1655_),
    .Y(_1741_)
);

NAND2X1 _3176_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [18]),
    .Y(_1742_)
);

OAI21X1 _3177_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(_1698_),
    .C(_1742_),
    .Y(_1743_)
);

NAND2X1 _3178_ (
    .A(_1022__bF$buf3),
    .B(_1743_),
    .Y(_1744_)
);

NAND3X1 _3179_ (
    .A(_1052__bF$buf2),
    .B(_1741_),
    .C(_1744_),
    .Y(_1745_)
);

NAND3X1 _3180_ (
    .A(_1087__bF$buf3),
    .B(_1554_),
    .C(_1557_),
    .Y(_1746_)
);

NAND3X1 _3181_ (
    .A(_1064__bF$buf4),
    .B(_1745_),
    .C(_1746_),
    .Y(_1747_)
);

NAND3X1 _3182_ (
    .A(_1050__bF$buf3),
    .B(_1403_),
    .C(_1404_),
    .Y(_1748_)
);

NAND3X1 _3183_ (
    .A(_1046__bF$buf1),
    .B(_1747_),
    .C(_1748_),
    .Y(_1749_)
);

NAND2X1 _3184_ (
    .A(_1063__bF$buf4),
    .B(_1123_),
    .Y(_1750_)
);

NAND3X1 _3185_ (
    .A(_1740_),
    .B(_1750_),
    .C(_1749_),
    .Y(_1751_)
);

OAI21X1 _3186_ (
    .A(_1046__bF$buf0),
    .B(_1111_),
    .C(_1749_),
    .Y(_1752_)
);

NAND2X1 _3187_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [19]),
    .B(_1752_),
    .Y(_1753_)
);

NAND2X1 _3188_ (
    .A(_1751_),
    .B(_1753_),
    .Y(_1754_)
);

INVX1 _3189_ (
    .A(_1754_),
    .Y(_1755_)
);

AOI22X1 _3190_ (
    .A(_1696_),
    .B(_1708_),
    .C(_1664_),
    .D(_1669_),
    .Y(_1756_)
);

NAND2X1 _3191_ (
    .A(_1756_),
    .B(_1675_),
    .Y(_1757_)
);

INVX1 _3192_ (
    .A(_1757_),
    .Y(_1758_)
);

NAND2X1 _3193_ (
    .A(_1709_),
    .B(_1670_),
    .Y(_1759_)
);

AOI21X1 _3194_ (
    .A(_1706_),
    .B(_1707_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [18]),
    .Y(_1760_)
);

NAND3X1 _3195_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [18]),
    .B(_1707_),
    .C(_1706_),
    .Y(_1761_)
);

OAI21X1 _3196_ (
    .A(_1725_),
    .B(_1760_),
    .C(_1761_),
    .Y(_1762_)
);

INVX1 _3197_ (
    .A(_1762_),
    .Y(_1763_)
);

OAI21X1 _3198_ (
    .A(_1672_),
    .B(_1759_),
    .C(_1763_),
    .Y(_1764_)
);

AOI21X1 _3199_ (
    .A(_1584_),
    .B(_1758_),
    .C(_1764_),
    .Y(_1765_)
);

NAND2X1 _3200_ (
    .A(_1027__bF$buf3),
    .B(_1765_),
    .Y(_1766_)
);

INVX1 _3201_ (
    .A(_1696_),
    .Y(_1767_)
);

AND2X2 _3202_ (
    .A(_1708_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .Y(_1768_)
);

OAI21X1 _3203_ (
    .A(_1767_),
    .B(_1731_),
    .C(_1768_),
    .Y(_1769_)
);

NAND3X1 _3204_ (
    .A(_1755_),
    .B(_1766_),
    .C(_1769_),
    .Y(_575_)
);

OAI21X1 _3205_ (
    .A(_1591_),
    .B(_1648_),
    .C(_1615_),
    .Y(_576_)
);

AOI21X1 _3206_ (
    .A(_576_),
    .B(_1756_),
    .C(_1762_),
    .Y(_577_)
);

OAI21X1 _3207_ (
    .A(_1757_),
    .B(_1626_),
    .C(_577_),
    .Y(_578_)
);

OAI21X1 _3208_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .B(_578_),
    .C(_1769_),
    .Y(_579_)
);

NAND2X1 _3209_ (
    .A(_1754_),
    .B(_579_),
    .Y(_580_)
);

AND2X2 _3210_ (
    .A(_580_),
    .B(_575_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [20])
);

INVX1 _3211_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [20]),
    .Y(_581_)
);

NAND2X1 _3212_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(_1687_),
    .Y(_582_)
);

INVX1 _3213_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [18]),
    .Y(_583_)
);

NAND2X1 _3214_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [19]),
    .Y(_584_)
);

OAI21X1 _3215_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(_583_),
    .C(_584_),
    .Y(_585_)
);

NAND2X1 _3216_ (
    .A(_1022__bF$buf2),
    .B(_585_),
    .Y(_586_)
);

NAND3X1 _3217_ (
    .A(_1052__bF$buf1),
    .B(_582_),
    .C(_586_),
    .Y(_587_)
);

OAI21X1 _3218_ (
    .A(_1052__bF$buf0),
    .B(_1608_),
    .C(_587_),
    .Y(_588_)
);

OAI21X1 _3219_ (
    .A(_1087__bF$buf2),
    .B(_1602_),
    .C(_1442_),
    .Y(_589_)
);

AOI21X1 _3220_ (
    .A(_589_),
    .B(_1050__bF$buf2),
    .C(_1063__bF$buf3),
    .Y(_590_)
);

OAI21X1 _3221_ (
    .A(_1050__bF$buf1),
    .B(_588_),
    .C(_590_),
    .Y(_591_)
);

NAND2X1 _3222_ (
    .A(_1063__bF$buf2),
    .B(_1141_),
    .Y(_592_)
);

NAND3X1 _3223_ (
    .A(_581_),
    .B(_592_),
    .C(_591_),
    .Y(_593_)
);

NAND2X1 _3224_ (
    .A(_1431_),
    .B(_1432_),
    .Y(_594_)
);

MUX2X1 _3225_ (
    .A(_588_),
    .B(_594_),
    .S(_1064__bF$buf3),
    .Y(_595_)
);

NAND2X1 _3226_ (
    .A(_1046__bF$buf7),
    .B(_595_),
    .Y(_596_)
);

NAND2X1 _3227_ (
    .A(_1063__bF$buf1),
    .B(_1149_),
    .Y(_597_)
);

NAND3X1 _3228_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [20]),
    .B(_597_),
    .C(_596_),
    .Y(_598_)
);

NAND3X1 _3229_ (
    .A(_1059_),
    .B(_1083_),
    .C(_1129_),
    .Y(_599_)
);

NAND3X1 _3230_ (
    .A(_1096_),
    .B(_1124_),
    .C(_599_),
    .Y(_600_)
);

AOI21X1 _3231_ (
    .A(_600_),
    .B(_1112_),
    .C(_1710_),
    .Y(_601_)
);

OAI21X1 _3232_ (
    .A(_601_),
    .B(_1304_),
    .C(_1722_),
    .Y(_602_)
);

NAND3X1 _3233_ (
    .A(_1697_),
    .B(_1695_),
    .C(_1694_),
    .Y(_603_)
);

AOI22X1 _3234_ (
    .A(_603_),
    .B(_1761_),
    .C(_1751_),
    .D(_1753_),
    .Y(_604_)
);

NAND2X1 _3235_ (
    .A(_1726_),
    .B(_604_),
    .Y(_605_)
);

AOI21X1 _3236_ (
    .A(_602_),
    .B(_1642_),
    .C(_605_),
    .Y(_606_)
);

NAND3X1 _3237_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [19]),
    .B(_1750_),
    .C(_1749_),
    .Y(_607_)
);

AOI21X1 _3238_ (
    .A(_1749_),
    .B(_1750_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [19]),
    .Y(_608_)
);

OAI21X1 _3239_ (
    .A(_608_),
    .B(_1696_),
    .C(_607_),
    .Y(_609_)
);

AOI21X1 _3240_ (
    .A(_1729_),
    .B(_604_),
    .C(_609_),
    .Y(_610_)
);

INVX1 _3241_ (
    .A(_610_),
    .Y(_611_)
);

OAI21X1 _3242_ (
    .A(_611_),
    .B(_606_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .Y(_612_)
);

AOI21X1 _3243_ (
    .A(_1749_),
    .B(_1750_),
    .C(_1740_),
    .Y(_613_)
);

NOR2X1 _3244_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .B(_613_),
    .Y(_614_)
);

OAI21X1 _3245_ (
    .A(_1754_),
    .B(_1765_),
    .C(_614_),
    .Y(_615_)
);

AND2X2 _3246_ (
    .A(_615_),
    .B(_612_),
    .Y(_616_)
);

NAND3X1 _3247_ (
    .A(_593_),
    .B(_598_),
    .C(_616_),
    .Y(_617_)
);

AOI21X1 _3248_ (
    .A(_596_),
    .B(_597_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [20]),
    .Y(_618_)
);

AOI21X1 _3249_ (
    .A(_591_),
    .B(_592_),
    .C(_581_),
    .Y(_619_)
);

NAND2X1 _3250_ (
    .A(_612_),
    .B(_615_),
    .Y(_620_)
);

OAI21X1 _3251_ (
    .A(_618_),
    .B(_619_),
    .C(_620_),
    .Y(_621_)
);

AND2X2 _3252_ (
    .A(_617_),
    .B(_621_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [21])
);

OAI21X1 _3253_ (
    .A(_1050__bF$buf0),
    .B(_1467_),
    .C(_1063__bF$buf0),
    .Y(_622_)
);

NAND3X1 _3254_ (
    .A(_1050__bF$buf5),
    .B(_1475_),
    .C(_1472_),
    .Y(_623_)
);

NAND2X1 _3255_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_1743_),
    .Y(_624_)
);

INVX1 _3256_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [19]),
    .Y(_625_)
);

NAND2X1 _3257_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [20]),
    .Y(_626_)
);

OAI21X1 _3258_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_625_),
    .C(_626_),
    .Y(_627_)
);

NAND2X1 _3259_ (
    .A(_1022__bF$buf1),
    .B(_627_),
    .Y(_628_)
);

NAND3X1 _3260_ (
    .A(_1052__bF$buf5),
    .B(_624_),
    .C(_628_),
    .Y(_629_)
);

NAND3X1 _3261_ (
    .A(_1087__bF$buf1),
    .B(_1652_),
    .C(_1656_),
    .Y(_630_)
);

NAND3X1 _3262_ (
    .A(_1064__bF$buf2),
    .B(_629_),
    .C(_630_),
    .Y(_631_)
);

NAND3X1 _3263_ (
    .A(_1046__bF$buf6),
    .B(_631_),
    .C(_623_),
    .Y(_632_)
);

NAND3X1 _3264_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [21]),
    .B(_632_),
    .C(_622_),
    .Y(_633_)
);

INVX1 _3265_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [21]),
    .Y(_634_)
);

OAI21X1 _3266_ (
    .A(_1046__bF$buf5),
    .B(_1171_),
    .C(_632_),
    .Y(_635_)
);

NAND2X1 _3267_ (
    .A(_634_),
    .B(_635_),
    .Y(_636_)
);

NAND2X1 _3268_ (
    .A(_633_),
    .B(_636_),
    .Y(_637_)
);

INVX1 _3269_ (
    .A(_637_),
    .Y(_638_)
);

INVX1 _3270_ (
    .A(_608_),
    .Y(_639_)
);

NAND3X1 _3271_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [20]),
    .B(_592_),
    .C(_591_),
    .Y(_640_)
);

NAND3X1 _3272_ (
    .A(_581_),
    .B(_597_),
    .C(_596_),
    .Y(_641_)
);

AOI22X1 _3273_ (
    .A(_641_),
    .B(_640_),
    .C(_607_),
    .D(_639_),
    .Y(_642_)
);

INVX1 _3274_ (
    .A(_642_),
    .Y(_643_)
);

AOI21X1 _3275_ (
    .A(_613_),
    .B(_593_),
    .C(_619_),
    .Y(_644_)
);

OAI21X1 _3276_ (
    .A(_643_),
    .B(_1765_),
    .C(_644_),
    .Y(_645_)
);

NAND2X1 _3277_ (
    .A(_1027__bF$buf2),
    .B(_645_),
    .Y(_646_)
);

OAI21X1 _3278_ (
    .A(_611_),
    .B(_606_),
    .C(_641_),
    .Y(_647_)
);

NAND3X1 _3279_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .B(_640_),
    .C(_647_),
    .Y(_648_)
);

NAND3X1 _3280_ (
    .A(_638_),
    .B(_648_),
    .C(_646_),
    .Y(_649_)
);

OAI21X1 _3281_ (
    .A(_1753_),
    .B(_618_),
    .C(_598_),
    .Y(_650_)
);

AOI21X1 _3282_ (
    .A(_578_),
    .B(_642_),
    .C(_650_),
    .Y(_651_)
);

OAI21X1 _3283_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .B(_651_),
    .C(_648_),
    .Y(_652_)
);

NAND2X1 _3284_ (
    .A(_637_),
    .B(_652_),
    .Y(_653_)
);

AND2X2 _3285_ (
    .A(_653_),
    .B(_649_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [22])
);

INVX1 _3286_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [22]),
    .Y(_654_)
);

NAND2X1 _3287_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_585_),
    .Y(_655_)
);

INVX1 _3288_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [20]),
    .Y(_656_)
);

NAND2X1 _3289_ (
    .A(_1034__bF$buf2),
    .B(_656_),
    .Y(_657_)
);

INVX1 _3290_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [21]),
    .Y(_658_)
);

NAND2X1 _3291_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(_658_),
    .Y(_659_)
);

NAND3X1 _3292_ (
    .A(_1022__bF$buf0),
    .B(_659_),
    .C(_657_),
    .Y(_660_)
);

NAND3X1 _3293_ (
    .A(_1052__bF$buf4),
    .B(_660_),
    .C(_655_),
    .Y(_661_)
);

NAND3X1 _3294_ (
    .A(_1087__bF$buf0),
    .B(_1684_),
    .C(_1688_),
    .Y(_662_)
);

AOI21X1 _3295_ (
    .A(_662_),
    .B(_661_),
    .C(_1050__bF$buf4),
    .Y(_663_)
);

AOI21X1 _3296_ (
    .A(_1507_),
    .B(_1510_),
    .C(_1064__bF$buf1),
    .Y(_664_)
);

OAI21X1 _3297_ (
    .A(_663_),
    .B(_664_),
    .C(_1046__bF$buf4),
    .Y(_665_)
);

NAND2X1 _3298_ (
    .A(_1063__bF$buf4),
    .B(_1215_),
    .Y(_666_)
);

NAND3X1 _3299_ (
    .A(_654_),
    .B(_666_),
    .C(_665_),
    .Y(_667_)
);

AOI21X1 _3300_ (
    .A(_665_),
    .B(_666_),
    .C(_654_),
    .Y(_668_)
);

INVX1 _3301_ (
    .A(_668_),
    .Y(_669_)
);

NAND2X1 _3302_ (
    .A(_667_),
    .B(_669_),
    .Y(_670_)
);

INVX1 _3303_ (
    .A(_670_),
    .Y(_671_)
);

NAND2X1 _3304_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [21]),
    .B(_635_),
    .Y(_672_)
);

INVX1 _3305_ (
    .A(_672_),
    .Y(_673_)
);

NOR2X1 _3306_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .B(_673_),
    .Y(_674_)
);

OAI21X1 _3307_ (
    .A(_638_),
    .B(_651_),
    .C(_674_),
    .Y(_675_)
);

OR2X2 _3308_ (
    .A(_635_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [21]),
    .Y(_676_)
);

AOI22X1 _3309_ (
    .A(_593_),
    .B(_598_),
    .C(_676_),
    .D(_672_),
    .Y(_677_)
);

OAI21X1 _3310_ (
    .A(_611_),
    .B(_606_),
    .C(_677_),
    .Y(_678_)
);

AOI21X1 _3311_ (
    .A(_622_),
    .B(_632_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [21]),
    .Y(_679_)
);

OAI21X1 _3312_ (
    .A(_679_),
    .B(_640_),
    .C(_633_),
    .Y(_680_)
);

INVX1 _3313_ (
    .A(_680_),
    .Y(_681_)
);

NAND2X1 _3314_ (
    .A(_681_),
    .B(_678_),
    .Y(_682_)
);

NAND2X1 _3315_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .B(_682_),
    .Y(_683_)
);

NAND3X1 _3316_ (
    .A(_671_),
    .B(_683_),
    .C(_675_),
    .Y(_684_)
);

INVX1 _3317_ (
    .A(_674_),
    .Y(_685_)
);

AOI21X1 _3318_ (
    .A(_645_),
    .B(_637_),
    .C(_685_),
    .Y(_686_)
);

AOI21X1 _3319_ (
    .A(_678_),
    .B(_681_),
    .C(_1027__bF$buf1),
    .Y(_687_)
);

OAI21X1 _3320_ (
    .A(_687_),
    .B(_686_),
    .C(_670_),
    .Y(_688_)
);

AND2X2 _3321_ (
    .A(_688_),
    .B(_684_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [23])
);

INVX1 _3322_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [23]),
    .Y(_689_)
);

NAND3X1 _3323_ (
    .A(_1087__bF$buf4),
    .B(_1741_),
    .C(_1744_),
    .Y(_690_)
);

NAND2X1 _3324_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf0 ),
    .B(_627_),
    .Y(_691_)
);

NAND2X1 _3325_ (
    .A(_1034__bF$buf1),
    .B(_658_),
    .Y(_692_)
);

INVX1 _3326_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [22]),
    .Y(_693_)
);

NAND2X1 _3327_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .B(_693_),
    .Y(_694_)
);

NAND3X1 _3328_ (
    .A(_1022__bF$buf6),
    .B(_694_),
    .C(_692_),
    .Y(_695_)
);

NAND3X1 _3329_ (
    .A(_1052__bF$buf3),
    .B(_695_),
    .C(_691_),
    .Y(_696_)
);

AOI21X1 _3330_ (
    .A(_690_),
    .B(_696_),
    .C(_1050__bF$buf3),
    .Y(_697_)
);

AOI21X1 _3331_ (
    .A(_1558_),
    .B(_1559_),
    .C(_1064__bF$buf0),
    .Y(_698_)
);

OAI21X1 _3332_ (
    .A(_697_),
    .B(_698_),
    .C(_1046__bF$buf3),
    .Y(_699_)
);

NAND2X1 _3333_ (
    .A(_1063__bF$buf3),
    .B(_1249_),
    .Y(_700_)
);

NAND3X1 _3334_ (
    .A(_689_),
    .B(_699_),
    .C(_700_),
    .Y(_701_)
);

OAI21X1 _3335_ (
    .A(_1046__bF$buf2),
    .B(_1239_),
    .C(_699_),
    .Y(_702_)
);

NAND2X1 _3336_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [23]),
    .B(_702_),
    .Y(_703_)
);

NAND2X1 _3337_ (
    .A(_701_),
    .B(_703_),
    .Y(_704_)
);

INVX1 _3338_ (
    .A(_704_),
    .Y(_705_)
);

NAND3X1 _3339_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [22]),
    .B(_666_),
    .C(_665_),
    .Y(_706_)
);

OAI21X1 _3340_ (
    .A(_1052__bF$buf2),
    .B(_1350_),
    .C(_1507_),
    .Y(_707_)
);

AOI21X1 _3341_ (
    .A(_1050__bF$buf2),
    .B(_707_),
    .C(_663_),
    .Y(_708_)
);

NAND2X1 _3342_ (
    .A(_1046__bF$buf1),
    .B(_708_),
    .Y(_709_)
);

NAND2X1 _3343_ (
    .A(_1063__bF$buf2),
    .B(_1205_),
    .Y(_710_)
);

NAND3X1 _3344_ (
    .A(_654_),
    .B(_710_),
    .C(_709_),
    .Y(_711_)
);

AOI22X1 _3345_ (
    .A(_633_),
    .B(_636_),
    .C(_711_),
    .D(_706_),
    .Y(_712_)
);

AND2X2 _3346_ (
    .A(_712_),
    .B(_642_),
    .Y(_713_)
);

NAND2X1 _3347_ (
    .A(_713_),
    .B(_1758_),
    .Y(_714_)
);

INVX1 _3348_ (
    .A(_706_),
    .Y(_715_)
);

AOI21X1 _3349_ (
    .A(_665_),
    .B(_666_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [22]),
    .Y(_716_)
);

OAI21X1 _3350_ (
    .A(_716_),
    .B(_715_),
    .C(_637_),
    .Y(_717_)
);

AOI21X1 _3351_ (
    .A(_673_),
    .B(_667_),
    .C(_668_),
    .Y(_718_)
);

OAI21X1 _3352_ (
    .A(_644_),
    .B(_717_),
    .C(_718_),
    .Y(_719_)
);

AOI21X1 _3353_ (
    .A(_1764_),
    .B(_713_),
    .C(_719_),
    .Y(_720_)
);

OAI21X1 _3354_ (
    .A(_714_),
    .B(_1626_),
    .C(_720_),
    .Y(_721_)
);

NOR2X1 _3355_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .B(_721_),
    .Y(_722_)
);

INVX1 _3356_ (
    .A(_722_),
    .Y(_723_)
);

OAI21X1 _3357_ (
    .A(_1046__bF$buf0),
    .B(_1215_),
    .C(_709_),
    .Y(_724_)
);

OAI21X1 _3358_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [22]),
    .B(_724_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .Y(_725_)
);

INVX1 _3359_ (
    .A(_725_),
    .Y(_726_)
);

OAI21X1 _3360_ (
    .A(_715_),
    .B(_682_),
    .C(_726_),
    .Y(_727_)
);

NAND3X1 _3361_ (
    .A(_705_),
    .B(_723_),
    .C(_727_),
    .Y(_728_)
);

OAI21X1 _3362_ (
    .A(_605_),
    .B(_1723_),
    .C(_610_),
    .Y(_729_)
);

OAI21X1 _3363_ (
    .A(_634_),
    .B(_635_),
    .C(_640_),
    .Y(_730_)
);

AOI22X1 _3364_ (
    .A(_636_),
    .B(_730_),
    .C(_729_),
    .D(_677_),
    .Y(_731_)
);

AOI21X1 _3365_ (
    .A(_731_),
    .B(_706_),
    .C(_725_),
    .Y(_732_)
);

OAI21X1 _3366_ (
    .A(_722_),
    .B(_732_),
    .C(_704_),
    .Y(_733_)
);

AND2X2 _3367_ (
    .A(_733_),
    .B(_728_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [24])
);

INVX1 _3368_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [24]),
    .Y(_734_)
);

OAI21X1 _3369_ (
    .A(_1022__bF$buf5),
    .B(_1700_),
    .C(_586_),
    .Y(_735_)
);

OAI21X1 _3370_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [20]),
    .C(_659_),
    .Y(_736_)
);

NAND2X1 _3371_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [23]),
    .Y(_737_)
);

OAI21X1 _3372_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(_693_),
    .C(_737_),
    .Y(_738_)
);

NAND2X1 _3373_ (
    .A(_1022__bF$buf4),
    .B(_738_),
    .Y(_739_)
);

OAI21X1 _3374_ (
    .A(_1022__bF$buf3),
    .B(_736_),
    .C(_739_),
    .Y(_740_)
);

MUX2X1 _3375_ (
    .A(_735_),
    .B(_740_),
    .S(_1087__bF$buf3),
    .Y(_741_)
);

AOI21X1 _3376_ (
    .A(_1603_),
    .B(_1601_),
    .C(_1064__bF$buf5),
    .Y(_742_)
);

AOI21X1 _3377_ (
    .A(_1064__bF$buf4),
    .B(_741_),
    .C(_742_),
    .Y(_743_)
);

NAND2X1 _3378_ (
    .A(_1063__bF$buf1),
    .B(_1291_),
    .Y(_744_)
);

OAI21X1 _3379_ (
    .A(_1063__bF$buf0),
    .B(_743_),
    .C(_744_),
    .Y(_745_)
);

NOR2X1 _3380_ (
    .A(_734_),
    .B(_745_),
    .Y(_746_)
);

INVX1 _3381_ (
    .A(_745_),
    .Y(_747_)
);

NOR2X1 _3382_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [24]),
    .B(_747_),
    .Y(_748_)
);

AOI22X1 _3383_ (
    .A(_701_),
    .B(_703_),
    .C(_669_),
    .D(_667_),
    .Y(_749_)
);

NAND2X1 _3384_ (
    .A(_677_),
    .B(_749_),
    .Y(_750_)
);

OR2X2 _3385_ (
    .A(_702_),
    .B(_689_),
    .Y(_751_)
);

AOI21X1 _3386_ (
    .A(_700_),
    .B(_699_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [23]),
    .Y(_752_)
);

OAI21X1 _3387_ (
    .A(_706_),
    .B(_752_),
    .C(_751_),
    .Y(_753_)
);

AOI21X1 _3388_ (
    .A(_680_),
    .B(_749_),
    .C(_753_),
    .Y(_754_)
);

OAI21X1 _3389_ (
    .A(_610_),
    .B(_750_),
    .C(_754_),
    .Y(_755_)
);

NOR2X1 _3390_ (
    .A(_605_),
    .B(_750_),
    .Y(_756_)
);

AOI21X1 _3391_ (
    .A(_1645_),
    .B(_756_),
    .C(_755_),
    .Y(_757_)
);

NOR2X1 _3392_ (
    .A(_1027__bF$buf0),
    .B(_757_),
    .Y(_758_)
);

NAND2X1 _3393_ (
    .A(_1027__bF$buf5),
    .B(_703_),
    .Y(_759_)
);

AOI21X1 _3394_ (
    .A(_721_),
    .B(_705_),
    .C(_759_),
    .Y(_760_)
);

NOR2X1 _3395_ (
    .A(_760_),
    .B(_758_),
    .Y(_761_)
);

OAI21X1 _3396_ (
    .A(_746_),
    .B(_748_),
    .C(_761_),
    .Y(_762_)
);

NAND2X1 _3397_ (
    .A(_734_),
    .B(_747_),
    .Y(_763_)
);

NAND2X1 _3398_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [24]),
    .B(_745_),
    .Y(_764_)
);

NAND2X1 _3399_ (
    .A(_764_),
    .B(_763_),
    .Y(_765_)
);

OAI21X1 _3400_ (
    .A(_760_),
    .B(_758_),
    .C(_765_),
    .Y(_766_)
);

AND2X2 _3401_ (
    .A(_762_),
    .B(_766_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [25])
);

NAND2X1 _3402_ (
    .A(_1063__bF$buf4),
    .B(_1331_),
    .Y(_767_)
);

NAND2X1 _3403_ (
    .A(_624_),
    .B(_628_),
    .Y(_768_)
);

OAI21X1 _3404_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [21]),
    .C(_694_),
    .Y(_769_)
);

INVX1 _3405_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [23]),
    .Y(_770_)
);

NAND2X1 _3406_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [24]),
    .Y(_771_)
);

OAI21X1 _3407_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf7 ),
    .B(_770_),
    .C(_771_),
    .Y(_772_)
);

NAND2X1 _3408_ (
    .A(_1022__bF$buf2),
    .B(_772_),
    .Y(_773_)
);

OAI21X1 _3409_ (
    .A(_1022__bF$buf1),
    .B(_769_),
    .C(_773_),
    .Y(_774_)
);

MUX2X1 _3410_ (
    .A(_774_),
    .B(_768_),
    .S(_1052__bF$buf1),
    .Y(_775_)
);

AOI21X1 _3411_ (
    .A(_1658_),
    .B(_1657_),
    .C(_1064__bF$buf3),
    .Y(_776_)
);

AOI21X1 _3412_ (
    .A(_1064__bF$buf2),
    .B(_775_),
    .C(_776_),
    .Y(_777_)
);

NAND2X1 _3413_ (
    .A(_1046__bF$buf7),
    .B(_777_),
    .Y(_778_)
);

NAND2X1 _3414_ (
    .A(_767_),
    .B(_778_),
    .Y(_779_)
);

NAND2X1 _3415_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [25]),
    .B(_779_),
    .Y(_780_)
);

OR2X2 _3416_ (
    .A(_779_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [25]),
    .Y(_781_)
);

NAND2X1 _3417_ (
    .A(_780_),
    .B(_781_),
    .Y(_782_)
);

INVX1 _3418_ (
    .A(_782_),
    .Y(_783_)
);

NAND2X1 _3419_ (
    .A(_642_),
    .B(_712_),
    .Y(_784_)
);

NOR2X1 _3420_ (
    .A(_1757_),
    .B(_784_),
    .Y(_785_)
);

INVX1 _3421_ (
    .A(_667_),
    .Y(_786_)
);

OAI21X1 _3422_ (
    .A(_672_),
    .B(_786_),
    .C(_669_),
    .Y(_787_)
);

AOI21X1 _3423_ (
    .A(_650_),
    .B(_712_),
    .C(_787_),
    .Y(_788_)
);

OAI21X1 _3424_ (
    .A(_577_),
    .B(_784_),
    .C(_788_),
    .Y(_789_)
);

AOI21X1 _3425_ (
    .A(_1584_),
    .B(_785_),
    .C(_789_),
    .Y(_790_)
);

OAI21X1 _3426_ (
    .A(_746_),
    .B(_748_),
    .C(_705_),
    .Y(_791_)
);

INVX1 _3427_ (
    .A(_703_),
    .Y(_792_)
);

INVX1 _3428_ (
    .A(_764_),
    .Y(_793_)
);

AOI21X1 _3429_ (
    .A(_763_),
    .B(_792_),
    .C(_793_),
    .Y(_794_)
);

OAI21X1 _3430_ (
    .A(_791_),
    .B(_790_),
    .C(_794_),
    .Y(_795_)
);

NAND2X1 _3431_ (
    .A(_1027__bF$buf4),
    .B(_795_),
    .Y(_796_)
);

OAI21X1 _3432_ (
    .A(_734_),
    .B(_745_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .Y(_797_)
);

INVX1 _3433_ (
    .A(_797_),
    .Y(_798_)
);

OAI21X1 _3434_ (
    .A(_748_),
    .B(_757_),
    .C(_798_),
    .Y(_799_)
);

NAND3X1 _3435_ (
    .A(_783_),
    .B(_799_),
    .C(_796_),
    .Y(_800_)
);

INVX1 _3436_ (
    .A(_791_),
    .Y(_801_)
);

INVX1 _3437_ (
    .A(_794_),
    .Y(_802_)
);

AOI21X1 _3438_ (
    .A(_721_),
    .B(_801_),
    .C(_802_),
    .Y(_803_)
);

OAI21X1 _3439_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .B(_803_),
    .C(_799_),
    .Y(_804_)
);

NAND2X1 _3440_ (
    .A(_782_),
    .B(_804_),
    .Y(_805_)
);

AND2X2 _3441_ (
    .A(_805_),
    .B(_800_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [26])
);

OAI21X1 _3442_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf5 ),
    .B(_736_),
    .C(_655_),
    .Y(_806_)
);

INVX1 _3443_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [24]),
    .Y(_807_)
);

NAND2X1 _3444_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf6 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [25]),
    .Y(_808_)
);

OAI21X1 _3445_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf5 ),
    .B(_807_),
    .C(_808_),
    .Y(_809_)
);

OAI22X1 _3446_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf4 ),
    .B(_809_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .D(_738_),
    .Y(_810_)
);

NAND2X1 _3447_ (
    .A(_1086_),
    .B(_810_),
    .Y(_811_)
);

OAI21X1 _3448_ (
    .A(_1052__bF$buf0),
    .B(_806_),
    .C(_811_),
    .Y(_812_)
);

AOI21X1 _3449_ (
    .A(_1690_),
    .B(_1689_),
    .C(_1064__bF$buf1),
    .Y(_813_)
);

AOI21X1 _3450_ (
    .A(_1064__bF$buf0),
    .B(_812_),
    .C(_813_),
    .Y(_814_)
);

NAND2X1 _3451_ (
    .A(_1046__bF$buf6),
    .B(_814_),
    .Y(_815_)
);

NAND2X1 _3452_ (
    .A(_1063__bF$buf3),
    .B(_1352_),
    .Y(_816_)
);

NAND2X1 _3453_ (
    .A(_816_),
    .B(_815_),
    .Y(_817_)
);

NAND2X1 _3454_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [26]),
    .B(_817_),
    .Y(_818_)
);

OR2X2 _3455_ (
    .A(_817_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [26]),
    .Y(_819_)
);

NAND2X1 _3456_ (
    .A(_818_),
    .B(_819_),
    .Y(_820_)
);

AND2X2 _3457_ (
    .A(_604_),
    .B(_1726_),
    .Y(_821_)
);

NAND3X1 _3458_ (
    .A(_677_),
    .B(_749_),
    .C(_821_),
    .Y(_822_)
);

AOI21X1 _3459_ (
    .A(_1642_),
    .B(_602_),
    .C(_822_),
    .Y(_823_)
);

AOI21X1 _3460_ (
    .A(_763_),
    .B(_764_),
    .C(_782_),
    .Y(_824_)
);

OAI21X1 _3461_ (
    .A(_755_),
    .B(_823_),
    .C(_824_),
    .Y(_825_)
);

OAI21X1 _3462_ (
    .A(_734_),
    .B(_745_),
    .C(_780_),
    .Y(_826_)
);

OAI21X1 _3463_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [25]),
    .B(_779_),
    .C(_826_),
    .Y(_827_)
);

NAND2X1 _3464_ (
    .A(_827_),
    .B(_825_),
    .Y(_828_)
);

NAND2X1 _3465_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf4 ),
    .B(_828_),
    .Y(_829_)
);

INVX1 _3466_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [25]),
    .Y(_830_)
);

OAI21X1 _3467_ (
    .A(_830_),
    .B(_779_),
    .C(_1027__bF$buf3),
    .Y(_831_)
);

INVX1 _3468_ (
    .A(_831_),
    .Y(_832_)
);

OAI21X1 _3469_ (
    .A(_783_),
    .B(_803_),
    .C(_832_),
    .Y(_833_)
);

NAND3X1 _3470_ (
    .A(_820_),
    .B(_833_),
    .C(_829_),
    .Y(_834_)
);

INVX1 _3471_ (
    .A(_820_),
    .Y(_835_)
);

AOI21X1 _3472_ (
    .A(_825_),
    .B(_827_),
    .C(_1027__bF$buf2),
    .Y(_836_)
);

AOI21X1 _3473_ (
    .A(_795_),
    .B(_782_),
    .C(_831_),
    .Y(_837_)
);

OAI21X1 _3474_ (
    .A(_836_),
    .B(_837_),
    .C(_835_),
    .Y(_838_)
);

AND2X2 _3475_ (
    .A(_838_),
    .B(_834_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [27])
);

AND2X2 _3476_ (
    .A(_691_),
    .B(_695_),
    .Y(_839_)
);

INVX1 _3477_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [26]),
    .Y(_840_)
);

NAND2X1 _3478_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf4 ),
    .B(_840_),
    .Y(_841_)
);

OAI21X1 _3479_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [25]),
    .C(_841_),
    .Y(_842_)
);

NAND2X1 _3480_ (
    .A(_1022__bF$buf0),
    .B(_842_),
    .Y(_843_)
);

OAI21X1 _3481_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .B(_772_),
    .C(_843_),
    .Y(_844_)
);

AOI22X1 _3482_ (
    .A(_1087__bF$buf2),
    .B(_839_),
    .C(_844_),
    .D(_1086_),
    .Y(_845_)
);

NOR2X1 _3483_ (
    .A(_1050__bF$buf1),
    .B(_845_),
    .Y(_846_)
);

AOI21X1 _3484_ (
    .A(_1745_),
    .B(_1746_),
    .C(_1064__bF$buf5),
    .Y(_847_)
);

OAI21X1 _3485_ (
    .A(_847_),
    .B(_846_),
    .C(_1046__bF$buf5),
    .Y(_848_)
);

OAI21X1 _3486_ (
    .A(_1046__bF$buf4),
    .B(_1406_),
    .C(_848_),
    .Y(_849_)
);

INVX1 _3487_ (
    .A(_849_),
    .Y(_850_)
);

NAND2X1 _3488_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [27]),
    .B(_850_),
    .Y(_851_)
);

INVX1 _3489_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [27]),
    .Y(_852_)
);

NAND2X1 _3490_ (
    .A(_852_),
    .B(_849_),
    .Y(_853_)
);

NAND2X1 _3491_ (
    .A(_853_),
    .B(_851_),
    .Y(_854_)
);

NOR2X1 _3492_ (
    .A(_830_),
    .B(_779_),
    .Y(_855_)
);

INVX1 _3493_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [26]),
    .Y(_856_)
);

NOR2X1 _3494_ (
    .A(_856_),
    .B(_817_),
    .Y(_857_)
);

AOI21X1 _3495_ (
    .A(_820_),
    .B(_855_),
    .C(_857_),
    .Y(_858_)
);

INVX1 _3496_ (
    .A(_818_),
    .Y(_859_)
);

NOR2X1 _3497_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [26]),
    .B(_817_),
    .Y(_860_)
);

OAI21X1 _3498_ (
    .A(_859_),
    .B(_860_),
    .C(_782_),
    .Y(_861_)
);

OAI21X1 _3499_ (
    .A(_794_),
    .B(_861_),
    .C(_858_),
    .Y(_862_)
);

NOR2X1 _3500_ (
    .A(_791_),
    .B(_861_),
    .Y(_863_)
);

AOI21X1 _3501_ (
    .A(_721_),
    .B(_863_),
    .C(_862_),
    .Y(_864_)
);

NAND2X1 _3502_ (
    .A(_1027__bF$buf1),
    .B(_864_),
    .Y(_865_)
);

NOR2X1 _3503_ (
    .A(_1027__bF$buf0),
    .B(_860_),
    .Y(_866_)
);

OAI21X1 _3504_ (
    .A(_859_),
    .B(_828_),
    .C(_866_),
    .Y(_867_)
);

NAND3X1 _3505_ (
    .A(_854_),
    .B(_865_),
    .C(_867_),
    .Y(_868_)
);

INVX1 _3506_ (
    .A(_854_),
    .Y(_869_)
);

INVX1 _3507_ (
    .A(_865_),
    .Y(_870_)
);

NAND3X1 _3508_ (
    .A(_818_),
    .B(_827_),
    .C(_825_),
    .Y(_871_)
);

AND2X2 _3509_ (
    .A(_871_),
    .B(_866_),
    .Y(_872_)
);

OAI21X1 _3510_ (
    .A(_870_),
    .B(_872_),
    .C(_869_),
    .Y(_873_)
);

AND2X2 _3511_ (
    .A(_873_),
    .B(_868_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [28])
);

OAI21X1 _3512_ (
    .A(_1050__bF$buf0),
    .B(_589_),
    .C(_1444_),
    .Y(_874_)
);

NOR2X1 _3513_ (
    .A(_1064__bF$buf4),
    .B(_588_),
    .Y(_875_)
);

NOR2X1 _3514_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [26]),
    .Y(_876_)
);

NOR2X1 _3515_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [27]),
    .B(_1034__bF$buf0),
    .Y(_877_)
);

OAI21X1 _3516_ (
    .A(_876_),
    .B(_877_),
    .C(_1022__bF$buf6),
    .Y(_878_)
);

OAI21X1 _3517_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .B(_809_),
    .C(_878_),
    .Y(_879_)
);

OAI21X1 _3518_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .C(_879_),
    .Y(_880_)
);

OAI21X1 _3519_ (
    .A(_1052__bF$buf5),
    .B(_740_),
    .C(_880_),
    .Y(_881_)
);

NOR2X1 _3520_ (
    .A(_1050__bF$buf5),
    .B(_881_),
    .Y(_882_)
);

OAI21X1 _3521_ (
    .A(_875_),
    .B(_882_),
    .C(_1046__bF$buf3),
    .Y(_883_)
);

OAI21X1 _3522_ (
    .A(_1046__bF$buf2),
    .B(_874_),
    .C(_883_),
    .Y(_884_)
);

NAND2X1 _3523_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [28]),
    .B(_884_),
    .Y(_885_)
);

OR2X2 _3524_ (
    .A(_884_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [28]),
    .Y(_886_)
);

NAND2X1 _3525_ (
    .A(_885_),
    .B(_886_),
    .Y(_887_)
);

OAI21X1 _3526_ (
    .A(_852_),
    .B(_850_),
    .C(_1027__bF$buf5),
    .Y(_888_)
);

INVX1 _3527_ (
    .A(_888_),
    .Y(_889_)
);

OAI21X1 _3528_ (
    .A(_869_),
    .B(_864_),
    .C(_889_),
    .Y(_890_)
);

INVX1 _3529_ (
    .A(_827_),
    .Y(_891_)
);

OAI21X1 _3530_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [27]),
    .B(_850_),
    .C(_859_),
    .Y(_892_)
);

OAI21X1 _3531_ (
    .A(_852_),
    .B(_849_),
    .C(_892_),
    .Y(_893_)
);

NOR2X1 _3532_ (
    .A(_891_),
    .B(_893_),
    .Y(_894_)
);

NAND2X1 _3533_ (
    .A(_852_),
    .B(_850_),
    .Y(_895_)
);

NAND2X1 _3534_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [27]),
    .B(_849_),
    .Y(_896_)
);

AOI21X1 _3535_ (
    .A(_895_),
    .B(_896_),
    .C(_820_),
    .Y(_897_)
);

OAI21X1 _3536_ (
    .A(_893_),
    .B(_897_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf3 ),
    .Y(_898_)
);

AOI21X1 _3537_ (
    .A(_825_),
    .B(_894_),
    .C(_898_),
    .Y(_899_)
);

INVX1 _3538_ (
    .A(_899_),
    .Y(_900_)
);

NAND3X1 _3539_ (
    .A(_887_),
    .B(_890_),
    .C(_900_),
    .Y(_901_)
);

INVX1 _3540_ (
    .A(_887_),
    .Y(_902_)
);

INVX1 _3541_ (
    .A(_862_),
    .Y(_903_)
);

INVX1 _3542_ (
    .A(_863_),
    .Y(_904_)
);

OAI21X1 _3543_ (
    .A(_790_),
    .B(_904_),
    .C(_903_),
    .Y(_905_)
);

AOI21X1 _3544_ (
    .A(_905_),
    .B(_854_),
    .C(_888_),
    .Y(_906_)
);

OAI21X1 _3545_ (
    .A(_899_),
    .B(_906_),
    .C(_902_),
    .Y(_907_)
);

AND2X2 _3546_ (
    .A(_907_),
    .B(_901_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [29])
);

NOR2X1 _3547_ (
    .A(_1052__bF$buf4),
    .B(_774_),
    .Y(_908_)
);

INVX1 _3548_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [27]),
    .Y(_909_)
);

NAND2X1 _3549_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf1 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [28]),
    .Y(_910_)
);

OAI21X1 _3550_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_0_bF$buf0 ),
    .B(_909_),
    .C(_910_),
    .Y(_911_)
);

NAND2X1 _3551_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf2 ),
    .B(_842_),
    .Y(_912_)
);

OAI21X1 _3552_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60_1_bF$buf1 ),
    .B(_911_),
    .C(_912_),
    .Y(_913_)
);

AOI21X1 _3553_ (
    .A(_1052__bF$buf3),
    .B(_913_),
    .C(_908_),
    .Y(_914_)
);

NOR2X1 _3554_ (
    .A(_1050__bF$buf4),
    .B(_914_),
    .Y(_915_)
);

AOI21X1 _3555_ (
    .A(_629_),
    .B(_630_),
    .C(_1064__bF$buf3),
    .Y(_916_)
);

OAI21X1 _3556_ (
    .A(_916_),
    .B(_915_),
    .C(_1046__bF$buf1),
    .Y(_917_)
);

OAI21X1 _3557_ (
    .A(_1046__bF$buf0),
    .B(_1477_),
    .C(_917_),
    .Y(_918_)
);

NAND2X1 _3558_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [29]),
    .B(_918_),
    .Y(_919_)
);

OR2X2 _3559_ (
    .A(_918_),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [29]),
    .Y(_920_)
);

NAND2X1 _3560_ (
    .A(_919_),
    .B(_920_),
    .Y(_921_)
);

INVX1 _3561_ (
    .A(_921_),
    .Y(_922_)
);

NAND2X1 _3562_ (
    .A(_854_),
    .B(_887_),
    .Y(_923_)
);

INVX1 _3563_ (
    .A(_896_),
    .Y(_924_)
);

INVX1 _3564_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [28]),
    .Y(_925_)
);

OAI21X1 _3565_ (
    .A(_925_),
    .B(_884_),
    .C(_1027__bF$buf4),
    .Y(_926_)
);

AOI21X1 _3566_ (
    .A(_887_),
    .B(_924_),
    .C(_926_),
    .Y(_927_)
);

OAI21X1 _3567_ (
    .A(_923_),
    .B(_864_),
    .C(_927_),
    .Y(_928_)
);

INVX1 _3568_ (
    .A(_885_),
    .Y(_929_)
);

AOI22X1 _3569_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf2 ),
    .B(_929_),
    .C(_899_),
    .D(_886_),
    .Y(_930_)
);

NAND3X1 _3570_ (
    .A(_922_),
    .B(_928_),
    .C(_930_),
    .Y(_931_)
);

NAND2X1 _3571_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf1 ),
    .B(_929_),
    .Y(_932_)
);

NAND2X1 _3572_ (
    .A(_824_),
    .B(_897_),
    .Y(_933_)
);

AOI21X1 _3573_ (
    .A(_897_),
    .B(_891_),
    .C(_893_),
    .Y(_934_)
);

OAI21X1 _3574_ (
    .A(_933_),
    .B(_757_),
    .C(_934_),
    .Y(_935_)
);

NAND3X1 _3575_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf0 ),
    .B(_886_),
    .C(_935_),
    .Y(_936_)
);

NAND3X1 _3576_ (
    .A(_932_),
    .B(_936_),
    .C(_928_),
    .Y(_937_)
);

NAND2X1 _3577_ (
    .A(_921_),
    .B(_937_),
    .Y(_938_)
);

AND2X2 _3578_ (
    .A(_938_),
    .B(_931_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [30])
);

INVX1 _3579_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_reg ),
    .Y(_939_)
);

OAI21X1 _3580_ (
    .A(_1021_),
    .B(_1026_),
    .C(_939_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_int )
);

NOR2X1 _3581_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_enable_reg_pp0_iter1 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .Y(_940_)
);

INVX8 _3582_ (
    .A(_940_),
    .Y(_941_)
);

NOR2X1 _3583_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 ),
    .B(_1021_),
    .Y(_942_)
);

NAND3X1 _3584_ (
    .A(_868_),
    .B(_942_),
    .C(_873_),
    .Y(_943_)
);

OAI21X1 _3585_ (
    .A(_925_),
    .B(_941__bF$buf8),
    .C(_943_),
    .Y(_508_)
);

INVX1 _3586_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [29]),
    .Y(_944_)
);

NAND3X1 _3587_ (
    .A(_901_),
    .B(_942_),
    .C(_907_),
    .Y(_945_)
);

OAI21X1 _3588_ (
    .A(_944_),
    .B(_941__bF$buf7),
    .C(_945_),
    .Y(_509_)
);

NAND2X1 _3589_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3_bF$buf5 ),
    .B(_940_),
    .Y(_946_)
);

NAND3X1 _3590_ (
    .A(_931_),
    .B(_942_),
    .C(_938_),
    .Y(_947_)
);

NAND2X1 _3591_ (
    .A(_946_),
    .B(_947_),
    .Y(_510_)
);

INVX8 _3592_ (
    .A(_942_),
    .Y(_948_)
);

OAI21X1 _3593_ (
    .A(_1089_),
    .B(_941__bF$buf6),
    .C(_948__bF$buf4),
    .Y(_511_)
);

OAI22X1 _3594_ (
    .A(_1091_),
    .B(_941__bF$buf5),
    .C(_1028_),
    .D(_948__bF$buf3),
    .Y(_512_)
);

OAI22X1 _3595_ (
    .A(_1115_),
    .B(_941__bF$buf4),
    .C(_1091_),
    .D(_948__bF$buf2),
    .Y(_513_)
);

OAI22X1 _3596_ (
    .A(_1174_),
    .B(_941__bF$buf3),
    .C(_1115_),
    .D(_948__bF$buf1),
    .Y(_514_)
);

OAI22X1 _3597_ (
    .A(_1209_),
    .B(_941__bF$buf2),
    .C(_1174_),
    .D(_948__bF$buf0),
    .Y(_515_)
);

OAI22X1 _3598_ (
    .A(_1232_),
    .B(_941__bF$buf1),
    .C(_1209_),
    .D(_948__bF$buf4),
    .Y(_516_)
);

OAI22X1 _3599_ (
    .A(_1274_),
    .B(_941__bF$buf0),
    .C(_1232_),
    .D(_948__bF$buf3),
    .Y(_517_)
);

OAI22X1 _3600_ (
    .A(_1396_),
    .B(_941__bF$buf8),
    .C(_1274_),
    .D(_948__bF$buf2),
    .Y(_518_)
);

OAI22X1 _3601_ (
    .A(_1424_),
    .B(_941__bF$buf7),
    .C(_1396_),
    .D(_948__bF$buf1),
    .Y(_519_)
);

OAI22X1 _3602_ (
    .A(_1400_),
    .B(_941__bF$buf6),
    .C(_1424_),
    .D(_948__bF$buf0),
    .Y(_520_)
);

OAI22X1 _3603_ (
    .A(_1427_),
    .B(_941__bF$buf5),
    .C(_1400_),
    .D(_948__bF$buf4),
    .Y(_521_)
);

OAI22X1 _3604_ (
    .A(_1468_),
    .B(_941__bF$buf4),
    .C(_1427_),
    .D(_948__bF$buf3),
    .Y(_522_)
);

OAI22X1 _3605_ (
    .A(_1503_),
    .B(_941__bF$buf3),
    .C(_1468_),
    .D(_948__bF$buf2),
    .Y(_523_)
);

OAI22X1 _3606_ (
    .A(_1555_),
    .B(_941__bF$buf2),
    .C(_1503_),
    .D(_948__bF$buf1),
    .Y(_524_)
);

OAI22X1 _3607_ (
    .A(_1597_),
    .B(_941__bF$buf1),
    .C(_1555_),
    .D(_948__bF$buf0),
    .Y(_525_)
);

OAI22X1 _3608_ (
    .A(_1653_),
    .B(_941__bF$buf0),
    .C(_1597_),
    .D(_948__bF$buf4),
    .Y(_526_)
);

OAI22X1 _3609_ (
    .A(_1685_),
    .B(_941__bF$buf8),
    .C(_1653_),
    .D(_948__bF$buf3),
    .Y(_527_)
);

OAI22X1 _3610_ (
    .A(_1698_),
    .B(_941__bF$buf7),
    .C(_1685_),
    .D(_948__bF$buf2),
    .Y(_528_)
);

OAI22X1 _3611_ (
    .A(_583_),
    .B(_941__bF$buf6),
    .C(_1698_),
    .D(_948__bF$buf1),
    .Y(_529_)
);

OAI22X1 _3612_ (
    .A(_625_),
    .B(_941__bF$buf5),
    .C(_583_),
    .D(_948__bF$buf0),
    .Y(_530_)
);

OAI22X1 _3613_ (
    .A(_656_),
    .B(_941__bF$buf4),
    .C(_625_),
    .D(_948__bF$buf4),
    .Y(_531_)
);

OAI22X1 _3614_ (
    .A(_658_),
    .B(_941__bF$buf3),
    .C(_656_),
    .D(_948__bF$buf3),
    .Y(_532_)
);

OAI22X1 _3615_ (
    .A(_693_),
    .B(_941__bF$buf2),
    .C(_658_),
    .D(_948__bF$buf2),
    .Y(_533_)
);

OAI22X1 _3616_ (
    .A(_770_),
    .B(_941__bF$buf1),
    .C(_693_),
    .D(_948__bF$buf1),
    .Y(_534_)
);

OAI22X1 _3617_ (
    .A(_807_),
    .B(_941__bF$buf0),
    .C(_770_),
    .D(_948__bF$buf0),
    .Y(_535_)
);

INVX1 _3618_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [25]),
    .Y(_949_)
);

OAI22X1 _3619_ (
    .A(_949_),
    .B(_941__bF$buf8),
    .C(_807_),
    .D(_948__bF$buf4),
    .Y(_536_)
);

OAI22X1 _3620_ (
    .A(_840_),
    .B(_941__bF$buf7),
    .C(_949_),
    .D(_948__bF$buf3),
    .Y(_537_)
);

OAI22X1 _3621_ (
    .A(_909_),
    .B(_941__bF$buf6),
    .C(_840_),
    .D(_948__bF$buf2),
    .Y(_538_)
);

NAND2X1 _3622_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [28]),
    .B(_940_),
    .Y(_950_)
);

OAI21X1 _3623_ (
    .A(_909_),
    .B(_948__bF$buf1),
    .C(_950_),
    .Y(_539_)
);

MUX2X1 _3624_ (
    .A(_948__bF$buf0),
    .B(_941__bF$buf5),
    .S(_1034__bF$buf3),
    .Y(_540_)
);

NAND2X1 _3625_ (
    .A(_942_),
    .B(_1065_),
    .Y(_951_)
);

OAI21X1 _3626_ (
    .A(_1022__bF$buf5),
    .B(_941__bF$buf4),
    .C(_951_),
    .Y(_541_)
);

INVX1 _3627_ (
    .A(_1179_),
    .Y(_952_)
);

NAND2X1 _3628_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_enable_reg_pp0_iter1 ),
    .B(_952_),
    .Y(_953_)
);

NOR2X1 _3629_ (
    .A(_1048_),
    .B(_953_),
    .Y(_954_)
);

INVX8 _3630_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 ),
    .Y(_955_)
);

INVX1 _3631_ (
    .A(_953_),
    .Y(_956_)
);

OAI21X1 _3632_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2]),
    .B(_956_),
    .C(_955__bF$buf4),
    .Y(_957_)
);

NOR2X1 _3633_ (
    .A(_954_),
    .B(_957_),
    .Y(_542_)
);

NOR2X1 _3634_ (
    .A(_1024_),
    .B(_953_),
    .Y(_958_)
);

OAI21X1 _3635_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3]),
    .B(_954_),
    .C(_955__bF$buf3),
    .Y(_959_)
);

OR2X2 _3636_ (
    .A(_959_),
    .B(_958_),
    .Y(_960_)
);

INVX1 _3637_ (
    .A(_960_),
    .Y(_543_)
);

OAI21X1 _3638_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(_958_),
    .C(_955__bF$buf2),
    .Y(_961_)
);

AOI21X1 _3639_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4]),
    .B(_958_),
    .C(_961_),
    .Y(_544_)
);

INVX1 _3640_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_condition_exit_pp0_iter1_stage0 ),
    .Y(_962_)
);

AOI22X1 _3641_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 ),
    .B(gnd),
    .C(_940_),
    .D(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [0]),
    .Y(_963_)
);

OAI21X1 _3642_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 ),
    .B(_962_),
    .C(_963_),
    .Y(_547_)
);

NAND2X1 _3643_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [1]),
    .B(_940_),
    .Y(_964_)
);

MUX2X1 _3644_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [1]),
    .B(gnd),
    .S(_955__bF$buf1),
    .Y(_965_)
);

OAI21X1 _3645_ (
    .A(_940_),
    .B(_965_),
    .C(_964_),
    .Y(_548_)
);

NOR2X1 _3646_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [2]),
    .Y(_966_)
);

OAI21X1 _3647_ (
    .A(_955__bF$buf0),
    .B(gnd),
    .C(_941__bF$buf3),
    .Y(_967_)
);

OAI22X1 _3648_ (
    .A(_1084_),
    .B(_941__bF$buf2),
    .C(_967_),
    .D(_966_),
    .Y(_549_)
);

NOR2X1 _3649_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [3]),
    .Y(_968_)
);

OAI21X1 _3650_ (
    .A(_955__bF$buf4),
    .B(gnd),
    .C(_941__bF$buf1),
    .Y(_969_)
);

OAI22X1 _3651_ (
    .A(_1113_),
    .B(_941__bF$buf0),
    .C(_969_),
    .D(_968_),
    .Y(_550_)
);

NOR2X1 _3652_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [4]),
    .Y(_970_)
);

OAI21X1 _3653_ (
    .A(_955__bF$buf3),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [4]),
    .C(_941__bF$buf8),
    .Y(_971_)
);

OAI22X1 _3654_ (
    .A(_1143_),
    .B(_941__bF$buf7),
    .C(_971_),
    .D(_970_),
    .Y(_551_)
);

NOR2X1 _3655_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [5]),
    .Y(_972_)
);

OAI21X1 _3656_ (
    .A(_955__bF$buf2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [5]),
    .C(_941__bF$buf6),
    .Y(_973_)
);

OAI22X1 _3657_ (
    .A(_1165_),
    .B(_941__bF$buf5),
    .C(_973_),
    .D(_972_),
    .Y(_552_)
);

NOR2X1 _3658_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [6]),
    .Y(_974_)
);

OAI21X1 _3659_ (
    .A(_955__bF$buf1),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [6]),
    .C(_941__bF$buf4),
    .Y(_975_)
);

OAI22X1 _3660_ (
    .A(_1207_),
    .B(_941__bF$buf3),
    .C(_975_),
    .D(_974_),
    .Y(_553_)
);

NOR2X1 _3661_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [7]),
    .Y(_976_)
);

OAI21X1 _3662_ (
    .A(_955__bF$buf0),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [7]),
    .C(_941__bF$buf2),
    .Y(_977_)
);

OAI22X1 _3663_ (
    .A(_1241_),
    .B(_941__bF$buf1),
    .C(_977_),
    .D(_976_),
    .Y(_554_)
);

NOR2X1 _3664_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [8]),
    .Y(_978_)
);

OAI21X1 _3665_ (
    .A(_955__bF$buf4),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [8]),
    .C(_941__bF$buf0),
    .Y(_979_)
);

OAI22X1 _3666_ (
    .A(_1283_),
    .B(_941__bF$buf8),
    .C(_979_),
    .D(_978_),
    .Y(_555_)
);

NOR2X1 _3667_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 ),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_5_out [9]),
    .Y(_980_)
);

OAI21X1 _3668_ (
    .A(_955__bF$buf3),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [9]),
    .C(_941__bF$buf7),
    .Y(_981_)
);

OAI22X1 _3669_ (
    .A(_1328_),
    .B(_941__bF$buf6),
    .C(_981_),
    .D(_980_),
    .Y(_556_)
);

AOI21X1 _3670_ (
    .A(_1344_),
    .B(_1347_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 ),
    .Y(_982_)
);

OAI21X1 _3671_ (
    .A(_955__bF$buf2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [10]),
    .C(_941__bF$buf5),
    .Y(_983_)
);

OAI22X1 _3672_ (
    .A(_1354_),
    .B(_941__bF$buf4),
    .C(_983_),
    .D(_982_),
    .Y(_557_)
);

AOI21X1 _3673_ (
    .A(_1380_),
    .B(_1383_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 ),
    .Y(_984_)
);

OAI21X1 _3674_ (
    .A(_955__bF$buf1),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [11]),
    .C(_941__bF$buf3),
    .Y(_985_)
);

OAI22X1 _3675_ (
    .A(_1394_),
    .B(_941__bF$buf2),
    .C(_985_),
    .D(_984_),
    .Y(_558_)
);

AOI21X1 _3676_ (
    .A(_1420_),
    .B(_1422_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .Y(_986_)
);

OAI21X1 _3677_ (
    .A(_955__bF$buf0),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [12]),
    .C(_941__bF$buf1),
    .Y(_987_)
);

OAI22X1 _3678_ (
    .A(_1437_),
    .B(_941__bF$buf0),
    .C(_987_),
    .D(_986_),
    .Y(_559_)
);

AOI21X1 _3679_ (
    .A(_1463_),
    .B(_1466_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 ),
    .Y(_988_)
);

OAI21X1 _3680_ (
    .A(_955__bF$buf4),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [13]),
    .C(_941__bF$buf8),
    .Y(_989_)
);

OAI22X1 _3681_ (
    .A(_1479_),
    .B(_941__bF$buf7),
    .C(_989_),
    .D(_988_),
    .Y(_560_)
);

AOI21X1 _3682_ (
    .A(_1500_),
    .B(_1501_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 ),
    .Y(_990_)
);

OAI21X1 _3683_ (
    .A(_955__bF$buf3),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [14]),
    .C(_941__bF$buf6),
    .Y(_991_)
);

OAI22X1 _3684_ (
    .A(_1514_),
    .B(_941__bF$buf5),
    .C(_991_),
    .D(_990_),
    .Y(_561_)
);

AOI21X1 _3685_ (
    .A(_1538_),
    .B(_1541_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 ),
    .Y(_992_)
);

OAI21X1 _3686_ (
    .A(_955__bF$buf2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [15]),
    .C(_941__bF$buf4),
    .Y(_993_)
);

OAI22X1 _3687_ (
    .A(_1542_),
    .B(_941__bF$buf3),
    .C(_993_),
    .D(_992_),
    .Y(_562_)
);

AOI21X1 _3688_ (
    .A(_1589_),
    .B(_1593_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 ),
    .Y(_994_)
);

OAI21X1 _3689_ (
    .A(_955__bF$buf1),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [16]),
    .C(_941__bF$buf2),
    .Y(_995_)
);

OAI22X1 _3690_ (
    .A(_1594_),
    .B(_941__bF$buf1),
    .C(_995_),
    .D(_994_),
    .Y(_563_)
);

AOI21X1 _3691_ (
    .A(_1651_),
    .B(_1647_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .Y(_996_)
);

OAI21X1 _3692_ (
    .A(_955__bF$buf0),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [17]),
    .C(_941__bF$buf0),
    .Y(_997_)
);

OAI22X1 _3693_ (
    .A(_1665_),
    .B(_941__bF$buf8),
    .C(_997_),
    .D(_996_),
    .Y(_564_)
);

AOI21X1 _3694_ (
    .A(_1683_),
    .B(_1681_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 ),
    .Y(_998_)
);

OAI21X1 _3695_ (
    .A(_955__bF$buf4),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [18]),
    .C(_941__bF$buf7),
    .Y(_999_)
);

OAI22X1 _3696_ (
    .A(_1697_),
    .B(_941__bF$buf6),
    .C(_999_),
    .D(_998_),
    .Y(_565_)
);

AOI21X1 _3697_ (
    .A(_1736_),
    .B(_1739_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 ),
    .Y(_1000_)
);

OAI21X1 _3698_ (
    .A(_955__bF$buf3),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [19]),
    .C(_941__bF$buf5),
    .Y(_1001_)
);

OAI22X1 _3699_ (
    .A(_1740_),
    .B(_941__bF$buf4),
    .C(_1001_),
    .D(_1000_),
    .Y(_566_)
);

AOI21X1 _3700_ (
    .A(_580_),
    .B(_575_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 ),
    .Y(_1002_)
);

OAI21X1 _3701_ (
    .A(_955__bF$buf2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [20]),
    .C(_941__bF$buf3),
    .Y(_1003_)
);

OAI22X1 _3702_ (
    .A(_581_),
    .B(_941__bF$buf2),
    .C(_1003_),
    .D(_1002_),
    .Y(_567_)
);

AOI21X1 _3703_ (
    .A(_617_),
    .B(_621_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 ),
    .Y(_1004_)
);

OAI21X1 _3704_ (
    .A(_955__bF$buf1),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [21]),
    .C(_941__bF$buf1),
    .Y(_1005_)
);

OAI22X1 _3705_ (
    .A(_634_),
    .B(_941__bF$buf0),
    .C(_1005_),
    .D(_1004_),
    .Y(_568_)
);

AOI21X1 _3706_ (
    .A(_653_),
    .B(_649_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .Y(_1006_)
);

OAI21X1 _3707_ (
    .A(_955__bF$buf0),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [22]),
    .C(_941__bF$buf8),
    .Y(_1007_)
);

OAI22X1 _3708_ (
    .A(_654_),
    .B(_941__bF$buf7),
    .C(_1007_),
    .D(_1006_),
    .Y(_569_)
);

AOI21X1 _3709_ (
    .A(_688_),
    .B(_684_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf3 ),
    .Y(_1008_)
);

OAI21X1 _3710_ (
    .A(_955__bF$buf4),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [23]),
    .C(_941__bF$buf6),
    .Y(_1009_)
);

OAI22X1 _3711_ (
    .A(_689_),
    .B(_941__bF$buf5),
    .C(_1009_),
    .D(_1008_),
    .Y(_570_)
);

NAND2X1 _3712_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [24]),
    .B(_940_),
    .Y(_1010_)
);

AOI21X1 _3713_ (
    .A(_733_),
    .B(_728_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf2 ),
    .Y(_1011_)
);

OAI21X1 _3714_ (
    .A(_955__bF$buf3),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [24]),
    .C(_941__bF$buf4),
    .Y(_1012_)
);

OAI21X1 _3715_ (
    .A(_1012_),
    .B(_1011_),
    .C(_1010_),
    .Y(_571_)
);

AOI21X1 _3716_ (
    .A(_762_),
    .B(_766_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf1 ),
    .Y(_1013_)
);

OAI21X1 _3717_ (
    .A(_955__bF$buf2),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [25]),
    .C(_941__bF$buf3),
    .Y(_1014_)
);

OAI22X1 _3718_ (
    .A(_830_),
    .B(_941__bF$buf2),
    .C(_1014_),
    .D(_1013_),
    .Y(_572_)
);

AOI21X1 _3719_ (
    .A(_805_),
    .B(_800_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf0 ),
    .Y(_1015_)
);

OAI21X1 _3720_ (
    .A(_955__bF$buf1),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [26]),
    .C(_941__bF$buf1),
    .Y(_1016_)
);

OAI22X1 _3721_ (
    .A(_856_),
    .B(_941__bF$buf0),
    .C(_1016_),
    .D(_1015_),
    .Y(_573_)
);

AOI21X1 _3722_ (
    .A(_838_),
    .B(_834_),
    .C(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init_bF$buf4 ),
    .Y(_1017_)
);

OAI21X1 _3723_ (
    .A(_955__bF$buf0),
    .B(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.zext_ln90 [27]),
    .C(_941__bF$buf8),
    .Y(_1018_)
);

OAI22X1 _3724_ (
    .A(_852_),
    .B(_941__bF$buf7),
    .C(_1018_),
    .D(_1017_),
    .Y(_574_)
);

OAI21X1 _3725_ (
    .A(_1021_),
    .B(_1026_),
    .C(grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58_ap_start_reg),
    .Y(_1019_)
);

NOR2X1 _3726_ (
    .A(ap_rst),
    .B(_1019_),
    .Y(_545_)
);

NOR2X1 _3727_ (
    .A(vdd),
    .B(ap_rst),
    .Y(_1020_)
);

AND2X2 _3728_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_int ),
    .B(_1020_),
    .Y(_546_)
);

BUFX2 _3729_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [1]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [1])
);

BUFX2 _3730_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [2]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [2])
);

BUFX2 _3731_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [3]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [3])
);

BUFX2 _3732_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [4]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [4])
);

BUFX2 _3733_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [5]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [5])
);

BUFX2 _3734_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [6])
);

BUFX2 _3735_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [7]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [7])
);

BUFX2 _3736_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [8])
);

BUFX2 _3737_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [9]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [9])
);

BUFX2 _3738_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [10]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [10])
);

BUFX2 _3739_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [11]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [11])
);

BUFX2 _3740_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [12]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [12])
);

BUFX2 _3741_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [13]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [13])
);

BUFX2 _3742_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [14]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [14])
);

BUFX2 _3743_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [15]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [15])
);

BUFX2 _3744_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [16]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [16])
);

BUFX2 _3745_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [17]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [17])
);

BUFX2 _3746_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [18]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [18])
);

BUFX2 _3747_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [19]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [19])
);

BUFX2 _3748_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [20]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [20])
);

BUFX2 _3749_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [21]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [21])
);

BUFX2 _3750_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [22]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [22])
);

BUFX2 _3751_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [23]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [23])
);

BUFX2 _3752_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [24]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [24])
);

BUFX2 _3753_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [25]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [25])
);

BUFX2 _3754_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [26]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [26])
);

BUFX2 _3755_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [27]),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.empty_8_fu_220_p3 [27])
);

DFFPOSX1 _3756_ (
    .CLK(ap_clk_bF$buf0),
    .D(_508_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [28])
);

DFFPOSX1 _3757_ (
    .CLK(ap_clk_bF$buf12),
    .D(_509_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [29])
);

DFFPOSX1 _3758_ (
    .CLK(ap_clk_bF$buf11),
    .D(_510_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.tmp_fu_139_p3 )
);

DFFPOSX1 _3759_ (
    .CLK(ap_clk_bF$buf10),
    .D(_511_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [0])
);

DFFPOSX1 _3760_ (
    .CLK(ap_clk_bF$buf9),
    .D(_512_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [1])
);

DFFPOSX1 _3761_ (
    .CLK(ap_clk_bF$buf8),
    .D(_513_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [2])
);

DFFPOSX1 _3762_ (
    .CLK(ap_clk_bF$buf7),
    .D(_514_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [3])
);

DFFPOSX1 _3763_ (
    .CLK(ap_clk_bF$buf6),
    .D(_515_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [4])
);

DFFPOSX1 _3764_ (
    .CLK(ap_clk_bF$buf5),
    .D(_516_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [5])
);

DFFPOSX1 _3765_ (
    .CLK(ap_clk_bF$buf4),
    .D(_517_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [6])
);

DFFPOSX1 _3766_ (
    .CLK(ap_clk_bF$buf3),
    .D(_518_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [7])
);

DFFPOSX1 _3767_ (
    .CLK(ap_clk_bF$buf2),
    .D(_519_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [8])
);

DFFPOSX1 _3768_ (
    .CLK(ap_clk_bF$buf1),
    .D(_520_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [9])
);

DFFPOSX1 _3769_ (
    .CLK(ap_clk_bF$buf0),
    .D(_521_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [10])
);

DFFPOSX1 _3770_ (
    .CLK(ap_clk_bF$buf12),
    .D(_522_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [11])
);

DFFPOSX1 _3771_ (
    .CLK(ap_clk_bF$buf11),
    .D(_523_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [12])
);

DFFPOSX1 _3772_ (
    .CLK(ap_clk_bF$buf10),
    .D(_524_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [13])
);

DFFPOSX1 _3773_ (
    .CLK(ap_clk_bF$buf9),
    .D(_525_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [14])
);

DFFPOSX1 _3774_ (
    .CLK(ap_clk_bF$buf8),
    .D(_526_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [15])
);

DFFPOSX1 _3775_ (
    .CLK(ap_clk_bF$buf7),
    .D(_527_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [16])
);

DFFPOSX1 _3776_ (
    .CLK(ap_clk_bF$buf6),
    .D(_528_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [17])
);

DFFPOSX1 _3777_ (
    .CLK(ap_clk_bF$buf5),
    .D(_529_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [18])
);

DFFPOSX1 _3778_ (
    .CLK(ap_clk_bF$buf4),
    .D(_530_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [19])
);

DFFPOSX1 _3779_ (
    .CLK(ap_clk_bF$buf3),
    .D(_531_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [20])
);

DFFPOSX1 _3780_ (
    .CLK(ap_clk_bF$buf2),
    .D(_532_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [21])
);

DFFPOSX1 _3781_ (
    .CLK(ap_clk_bF$buf1),
    .D(_533_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [22])
);

DFFPOSX1 _3782_ (
    .CLK(ap_clk_bF$buf0),
    .D(_534_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [23])
);

DFFPOSX1 _3783_ (
    .CLK(ap_clk_bF$buf12),
    .D(_535_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [24])
);

DFFPOSX1 _3784_ (
    .CLK(ap_clk_bF$buf11),
    .D(_536_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [25])
);

DFFPOSX1 _3785_ (
    .CLK(ap_clk_bF$buf10),
    .D(_537_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [26])
);

DFFPOSX1 _3786_ (
    .CLK(ap_clk_bF$buf9),
    .D(_538_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [27])
);

DFFPOSX1 _3787_ (
    .CLK(ap_clk_bF$buf8),
    .D(_539_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.q6_fu_72 [28])
);

DFFPOSX1 _3788_ (
    .CLK(ap_clk_bF$buf7),
    .D(_540_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [0])
);

DFFPOSX1 _3789_ (
    .CLK(ap_clk_bF$buf6),
    .D(_541_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [1])
);

DFFPOSX1 _3790_ (
    .CLK(ap_clk_bF$buf5),
    .D(_542_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [2])
);

DFFPOSX1 _3791_ (
    .CLK(ap_clk_bF$buf4),
    .D(_543_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [3])
);

DFFPOSX1 _3792_ (
    .CLK(ap_clk_bF$buf3),
    .D(_544_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.i1_fu_60 [4])
);

DFFPOSX1 _3793_ (
    .CLK(ap_clk_bF$buf2),
    .D(_545_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_enable_reg_pp0_iter1 )
);

DFFPOSX1 _3794_ (
    .CLK(ap_clk_bF$buf1),
    .D(_546_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_reg )
);

DFFPOSX1 _3795_ (
    .CLK(ap_clk_bF$buf0),
    .D(_547_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [0])
);

DFFPOSX1 _3796_ (
    .CLK(ap_clk_bF$buf12),
    .D(_548_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [1])
);

DFFPOSX1 _3797_ (
    .CLK(ap_clk_bF$buf11),
    .D(_549_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [2])
);

DFFPOSX1 _3798_ (
    .CLK(ap_clk_bF$buf10),
    .D(_550_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [3])
);

DFFPOSX1 _3799_ (
    .CLK(ap_clk_bF$buf9),
    .D(_551_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [4])
);

DFFPOSX1 _3800_ (
    .CLK(ap_clk_bF$buf8),
    .D(_552_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [5])
);

DFFPOSX1 _3801_ (
    .CLK(ap_clk_bF$buf7),
    .D(_553_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [6])
);

DFFPOSX1 _3802_ (
    .CLK(ap_clk_bF$buf6),
    .D(_554_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [7])
);

DFFPOSX1 _3803_ (
    .CLK(ap_clk_bF$buf5),
    .D(_555_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [8])
);

DFFPOSX1 _3804_ (
    .CLK(ap_clk_bF$buf4),
    .D(_556_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [9])
);

DFFPOSX1 _3805_ (
    .CLK(ap_clk_bF$buf3),
    .D(_557_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [10])
);

DFFPOSX1 _3806_ (
    .CLK(ap_clk_bF$buf2),
    .D(_558_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [11])
);

DFFPOSX1 _3807_ (
    .CLK(ap_clk_bF$buf1),
    .D(_559_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [12])
);

DFFPOSX1 _3808_ (
    .CLK(ap_clk_bF$buf0),
    .D(_560_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [13])
);

DFFPOSX1 _3809_ (
    .CLK(ap_clk_bF$buf12),
    .D(_561_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [14])
);

DFFPOSX1 _3810_ (
    .CLK(ap_clk_bF$buf11),
    .D(_562_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [15])
);

DFFPOSX1 _3811_ (
    .CLK(ap_clk_bF$buf10),
    .D(_563_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [16])
);

DFFPOSX1 _3812_ (
    .CLK(ap_clk_bF$buf9),
    .D(_564_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [17])
);

DFFPOSX1 _3813_ (
    .CLK(ap_clk_bF$buf8),
    .D(_565_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [18])
);

DFFPOSX1 _3814_ (
    .CLK(ap_clk_bF$buf7),
    .D(_566_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [19])
);

DFFPOSX1 _3815_ (
    .CLK(ap_clk_bF$buf6),
    .D(_567_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [20])
);

DFFPOSX1 _3816_ (
    .CLK(ap_clk_bF$buf5),
    .D(_568_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [21])
);

DFFPOSX1 _3817_ (
    .CLK(ap_clk_bF$buf4),
    .D(_569_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [22])
);

DFFPOSX1 _3818_ (
    .CLK(ap_clk_bF$buf3),
    .D(_570_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [23])
);

DFFPOSX1 _3819_ (
    .CLK(ap_clk_bF$buf2),
    .D(_571_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [24])
);

DFFPOSX1 _3820_ (
    .CLK(ap_clk_bF$buf1),
    .D(_572_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [25])
);

DFFPOSX1 _3821_ (
    .CLK(ap_clk_bF$buf0),
    .D(_573_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [26])
);

DFFPOSX1 _3822_ (
    .CLK(ap_clk_bF$buf12),
    .D(_574_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.s_22_fu_64 [27])
);

INVX1 _3823_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_int ),
    .Y(_1772_)
);

INVX1 _3824_ (
    .A(grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58_ap_start_reg),
    .Y(_1773_)
);

NAND2X1 _3825_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.flow_control_loop_pipe_sequential_init_U.ap_done_cache ),
    .B(_1773_),
    .Y(_1774_)
);

NAND2X1 _3826_ (
    .A(_1772_),
    .B(_1774_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done )
);

INVX1 _3827_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.flow_control_loop_pipe_sequential_init_U.ap_loop_init_int ),
    .Y(_1775_)
);

NOR2X1 _3828_ (
    .A(_1773_),
    .B(_1775_),
    .Y(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_loop_init )
);

AOI21X1 _3829_ (
    .A(_1774_),
    .B(_1772_),
    .C(ap_rst),
    .Y(_1770_)
);

NOR2X1 _3830_ (
    .A(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.ap_done_int ),
    .B(ap_rst),
    .Y(_1776_)
);

OAI21X1 _3831_ (
    .A(_1775_),
    .B(grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58_ap_start_reg),
    .C(_1776_),
    .Y(_1771_)
);

DFFPOSX1 _3832_ (
    .CLK(ap_clk_bF$buf11),
    .D(_1770_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.flow_control_loop_pipe_sequential_init_U.ap_done_cache )
);

DFFPOSX1 _3833_ (
    .CLK(ap_clk_bF$buf10),
    .D(_1771_),
    .Q(\grp_fxp_sqrt_top_Pipeline_VITIS_LOOP_104_1_fu_58.flow_control_loop_pipe_sequential_init_U.ap_loop_init_int )
);

BUFX2 _3834_ (
    .A(_1777_),
    .Y(ap_done)
);

BUFX2 _3835_ (
    .A(_1778_),
    .Y(ap_idle)
);

BUFX2 _3836_ (
    .A(_1777_),
    .Y(ap_ready)
);

BUFX2 _3837_ (
    .A(_1779_[0]),
    .Y(ap_return[0])
);

BUFX2 _3838_ (
    .A(_1779_[1]),
    .Y(ap_return[1])
);

BUFX2 _3839_ (
    .A(_1779_[10]),
    .Y(ap_return[10])
);

BUFX2 _3840_ (
    .A(_1779_[11]),
    .Y(ap_return[11])
);

BUFX2 _3841_ (
    .A(_1779_[12]),
    .Y(ap_return[12])
);

BUFX2 _3842_ (
    .A(_1779_[13]),
    .Y(ap_return[13])
);

BUFX2 _3843_ (
    .A(_1779_[14]),
    .Y(ap_return[14])
);

BUFX2 _3844_ (
    .A(_1779_[15]),
    .Y(ap_return[15])
);

BUFX2 _3845_ (
    .A(_1779_[16]),
    .Y(ap_return[16])
);

BUFX2 _3846_ (
    .A(_1779_[17]),
    .Y(ap_return[17])
);

BUFX2 _3847_ (
    .A(_1779_[18]),
    .Y(ap_return[18])
);

BUFX2 _3848_ (
    .A(_1779_[19]),
    .Y(ap_return[19])
);

BUFX2 _3849_ (
    .A(_1779_[2]),
    .Y(ap_return[2])
);

BUFX2 _3850_ (
    .A(_1779_[20]),
    .Y(ap_return[20])
);

BUFX2 _3851_ (
    .A(_1779_[21]),
    .Y(ap_return[21])
);

BUFX2 _3852_ (
    .A(_1779_[22]),
    .Y(ap_return[22])
);

BUFX2 _3853_ (
    .A(_1779_[23]),
    .Y(ap_return[23])
);

BUFX2 _3854_ (
    .A(_1779_[24]),
    .Y(ap_return[24])
);

BUFX2 _3855_ (
    .A(_1779_[25]),
    .Y(ap_return[25])
);

BUFX2 _3856_ (
    .A(_1779_[26]),
    .Y(ap_return[26])
);

BUFX2 _3857_ (
    .A(_1779_[27]),
    .Y(ap_return[27])
);

BUFX2 _3858_ (
    .A(_1779_[3]),
    .Y(ap_return[3])
);

BUFX2 _3859_ (
    .A(_1779_[4]),
    .Y(ap_return[4])
);

BUFX2 _3860_ (
    .A(_1779_[5]),
    .Y(ap_return[5])
);

BUFX2 _3861_ (
    .A(_1779_[6]),
    .Y(ap_return[6])
);

BUFX2 _3862_ (
    .A(_1779_[7]),
    .Y(ap_return[7])
);

BUFX2 _3863_ (
    .A(_1779_[8]),
    .Y(ap_return[8])
);

BUFX2 _3864_ (
    .A(_1779_[9]),
    .Y(ap_return[9])
);

endmodule
