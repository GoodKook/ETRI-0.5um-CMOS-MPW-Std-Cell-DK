magic
tech scmos
magscale 1 2
timestamp 1727735982
<< error_s >>
rect 122 1149 1219 1161
rect 760 1101 762 1141
rect 610 1089 612 1101
rect 864 1061 868 1141
rect 760 909 762 941
rect 864 909 868 949
rect 119 889 1172 901
rect 0 834 1172 846
rect 0 594 1109 606
rect 0 534 510 546
rect 800 534 975 546
rect 108 294 800 306
rect 865 294 983 306
rect 43 234 1237 246
rect 81 -6 1307 6
<< metal1 >>
rect -97 1163 -37 1214
rect -97 1147 42 1163
rect -97 848 -37 1147
rect 1387 903 1447 1201
rect 1252 887 1447 903
rect -97 832 24 848
rect -97 548 -37 832
rect 1387 608 1447 887
rect 1160 592 1447 608
rect -97 532 21 548
rect -97 248 -37 532
rect 1387 308 1447 592
rect 949 292 1447 308
rect -97 232 28 248
rect -97 -47 -37 232
rect 1387 8 1447 292
rect 1292 -8 1447 8
rect 1387 -57 1447 -8
use AND2X1  AND2X1_0
timestamp 1727692839
transform 1 0 0 0 1 0
box -13 -8 112 252
use AND2X2  AND2X2_0
timestamp 1727694586
transform 1 0 92 0 1 0
box -12 -8 112 252
use AOI21X1  AOI21X1_0
timestamp 1727693469
transform 1 0 184 0 1 0
box -12 -8 112 252
use AOI22X1  AOI22X1_0
timestamp 1727694220
transform 1 0 276 0 1 0
box -14 -8 132 252
use BUFX2  BUFX2_0
timestamp 1727694371
transform 1 0 388 0 1 0
box -12 -8 92 252
use BUFX4  BUFX4_0
timestamp 1727694467
transform 1 0 460 0 1 0
box -13 -8 114 252
use CLKBUF1  CLKBUF1_0
timestamp 1727732147
transform 1 0 552 0 1 0
box -12 -8 212 252
use CLKBUF2  CLKBUF2_0
timestamp 1727732269
transform 1 0 738 0 1 0
box -12 -8 292 252
use CLKBUF3  CLKBUF3_0
timestamp 1727732429
transform 1 0 1005 0 1 0
box -12 -8 374 252
use DFFNEGX1  DFFNEGX1_0
timestamp 1727732648
transform 1 0 0 0 1 300
box -13 -8 252 252
use DFFPOSX1  DFFPOSX1_0
timestamp 1727732734
transform 1 0 230 0 1 300
box -13 -8 253 252
use DFFSR  DFFSR_0
timestamp 1727696105
transform 1 0 470 0 1 300
box -12 -8 492 252
use FAX1  FAX1_0
timestamp 1727136778
transform 1 0 191 0 1 895
box -13 -8 313 272
use FILL  FILL_0
timestamp 1727732812
transform 1 0 957 0 1 300
box -12 -8 32 252
use HAX1  HAX1_0
timestamp 1727136778
transform 1 0 500 0 1 895
box -13 -8 213 272
use INVX1  INVX1_0
timestamp 1727732874
transform 1 0 0 0 1 600
box -12 -8 72 252
use INVX2  INVX2_0
timestamp 1727732939
transform 1 0 46 0 1 600
box -12 -8 72 252
use INVX4  INVX4_0
timestamp 1727733003
transform 1 0 92 0 1 600
box -12 -8 92 252
use INVX8  INVX8_0
timestamp 1727733069
transform 1 0 157 0 1 600
box -12 -8 133 252
use LATCH  LATCH_0
timestamp 1727136778
transform 1 0 41 0 1 895
box -12 -8 153 272
use MUX2X1  MUX2X1_0
timestamp 1727733471
transform 1 0 262 0 1 600
box -12 -8 131 252
use NAND2X1  NAND2X1_0
timestamp 1727733579
transform 1 0 383 0 1 600
box -12 -8 92 252
use NAND3X1  NAND3X1_0
timestamp 1727733736
transform 1 0 449 0 1 600
box -12 -8 112 252
use NOR2X1  NOR2X1_0
timestamp 1727734357
transform 1 0 536 0 1 600
box -12 -8 92 252
use NOR3X1  NOR3X1_0
timestamp 1727734009
transform 1 0 602 0 1 600
box -12 -8 192 253
use OAI21X1  OAI21X1_0
timestamp 1727734141
transform 1 0 776 0 1 600
box -12 -8 112 252
use OAI22X1  OAI22X1_0
timestamp 1727734691
transform 1 0 867 0 1 600
box -12 -8 132 252
use OR2X1  OR2X1_0
timestamp 1727734834
transform 1 0 976 0 1 600
box -13 -8 112 252
use OR2X2  OR2X2_0
timestamp 1727735028
transform 1 0 1067 0 1 600
box -12 -8 112 252
use TBUFX1  TBUFX1_0
timestamp 1727136778
transform 1 0 710 0 1 895
box -14 -8 113 272
use TBUFX2  TBUFX2_0
timestamp 1727136778
transform 1 0 820 0 1 895
box -13 -8 153 272
use XNOR2X1  XNOR2X1_0
timestamp 1727423980
transform 1 0 970 0 1 895
box -12 -8 152 272
use XOR2X1  XOR2X1_0
timestamp 1727424219
transform 1 0 1118 0 1 895
box -12 -8 151 272
<< labels >>
rlabel metal1 -73 921 -73 921 0 vdd
port 1 nsew power bidirectional abutment
rlabel metal1 1414 905 1414 905 0 gnd
port 2 nsew ground bidirectional abutment
<< end >>
