magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -56 -56 254 84
<< diffusion >>
rect 5 5 193 23
<< metal1 >>
rect 4 4 194 24
<< end >>
