** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1_TB.sch
**.subckt inverter_x1_TB
Vdd VDD GND 5
R1 VDD Vout 1mega m=1
Vin Vin GND 0
x1 Vin Vout VDD GND inverter_x1
**** begin user architecture code



* ngspice commands
.include ~/ETRI050_DesignKit/devel/tech/05cmos_model_240201.lib
.dc vin 0 5 0.01
.save all



**** end user architecture code
**.ends

* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1.sym # of pins=4
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1.sym
.include ../inverter_x1.spice
.GLOBAL VDD
.GLOBAL GND
.end
