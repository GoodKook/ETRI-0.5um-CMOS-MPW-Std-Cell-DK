magic
tech scmos
magscale 1 6
timestamp 1569139307
<< checkpaint >>
rect -146 -140 450 1376
<< ntransistor >>
rect 52 0 66 1200
rect 238 0 252 1200
<< ndiffusion >>
rect 0 0 52 1200
rect 66 0 238 1200
rect 252 0 304 1200
<< polysilicon >>
rect 41 1220 77 1256
rect 227 1220 263 1256
rect 52 1200 66 1220
rect 238 1200 252 1220
rect 52 -20 66 0
rect 238 -20 252 0
<< metal1 >>
rect 41 1220 77 1256
rect 227 1220 263 1256
rect -24 0 76 1200
rect 92 0 212 1200
rect 228 0 328 1200
<< metal2 >>
rect -24 0 76 1200
rect 98 0 206 1200
rect 228 0 328 1200
<< metal3 >>
rect -26 0 78 1200
rect 226 0 330 1200
use CONT  CONT_0
timestamp 1569139307
transform 1 0 245 0 1 1238
box -6 -6 6 6
use CONT  CONT_1
timestamp 1569139307
transform 1 0 59 0 1 1238
box -6 -6 6 6
use CONT  CONT_2
array 0 0 0 0 28 36
timestamp 1569139307
transform 1 0 278 0 1 96
box -6 -6 6 6
use CONT  CONT_3
array 0 0 0 0 28 36
timestamp 1569139307
transform 1 0 26 0 1 96
box -6 -6 6 6
use CONT  CONT_4
array 0 0 0 0 28 36
timestamp 1569139307
transform 1 0 152 0 1 96
box -6 -6 6 6
use VIA1  VIA1_0
array 0 1 64 0 32 36
timestamp 1569139307
transform 1 0 120 0 1 24
box -8 -8 8 8
use VIA1  VIA1_1
array 0 1 60 0 32 36
timestamp 1569139307
transform 1 0 248 0 1 24
box -8 -8 8 8
use VIA1  VIA1_2
array 0 1 60 0 32 36
timestamp 1569139307
transform 1 0 -4 0 1 24
box -8 -8 8 8
<< end >>
