magic
tech scmos
magscale 1 30
timestamp 1741135076
<< checkpaint >>
rect -1237 8506 15389 36025
rect -1100 8445 13695 8506
rect -1100 8350 12430 8445
rect -1100 -3460 11590 8350
<< nwell >>
rect 0 30150 12195 32010
rect 0 20350 12200 28350
rect 100 9150 12100 16950
<< psubstratepdiff >>
rect 100 32550 12100 34210
<< nsubstratendiff >>
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
<< metal3 >>
rect 100 32550 12100 34210
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 6600 0 1 9150
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 600 0 1 9150
box -35 0 5035 25060
use pad80_CDNS_704676826050  pad80_CDNS_704676826050_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 1850 0 1 0
box 0 0 8500 8500
<< end >>
