magic
tech scmos
timestamp 1723010178
<< checkpaint >>
rect -20 -20 110 110
use pdiode_CDNS_7230122529126  pdiode_CDNS_7230122529126_0
timestamp 1723012252
transform 1 0 0 0 1 0
box 0 0 90 90
<< end >>
