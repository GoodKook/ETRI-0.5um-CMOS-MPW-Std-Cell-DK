magic
tech scmos
magscale 1 2
timestamp 1702308645
<< nwell >>
rect -13 153 74 272
<< ntransistor >>
rect 18 14 22 34
rect 38 14 42 34
<< ptransistor >>
rect 18 166 22 246
rect 32 166 36 246
<< ndiffusion >>
rect 16 14 18 34
rect 22 14 24 34
rect 36 14 38 34
rect 42 14 44 34
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 32 246
rect 36 166 38 246
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 34
rect 44 14 56 34
<< pdcontact >>
rect 4 166 16 246
rect 38 166 50 246
<< psubstratepcontact >>
rect -7 -6 67 6
<< nsubstratencontact >>
rect -7 254 67 266
<< polysilicon >>
rect 18 246 22 250
rect 32 246 36 250
rect 18 117 22 166
rect 32 164 36 166
rect 32 160 42 164
rect 17 105 22 117
rect 18 34 22 105
rect 38 117 42 160
rect 38 105 43 117
rect 38 34 42 105
rect 18 10 22 14
rect 38 10 42 14
<< polycontact >>
rect 5 105 17 117
rect 43 105 55 117
<< metal1 >>
rect -7 266 67 268
rect -7 252 67 254
rect 4 246 16 252
rect 26 166 38 174
rect 3 123 17 137
rect 5 117 17 123
rect 26 117 34 166
rect 43 123 57 137
rect 43 117 55 123
rect 23 103 37 117
rect 26 34 34 103
rect 4 8 16 14
rect 44 8 56 14
rect -7 6 67 8
rect -7 -8 67 -6
<< m1p >>
rect -7 252 67 268
rect 3 123 17 137
rect 43 123 57 137
rect 23 103 37 117
rect -7 -8 67 8
<< labels >>
rlabel nsubstratencontact 30 260 30 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 30 0 30 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 10 127 10 127 0 A
port 1 nsew signal input
rlabel metal1 50 127 50 127 0 B
port 2 nsew signal input
rlabel metal1 30 111 30 111 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
