magic
tech scmos
magscale 1 2
timestamp 1702508443
<< nwell >>
rect -13 154 213 272
<< ntransistor >>
rect 23 14 27 54
rect 33 14 37 54
rect 73 14 77 34
rect 93 14 97 54
rect 113 14 117 54
rect 133 14 137 54
rect 173 14 177 34
<< ptransistor >>
rect 23 206 27 246
rect 43 206 47 246
rect 83 206 87 246
rect 103 206 107 246
rect 123 166 127 246
rect 133 166 137 246
rect 173 206 177 246
<< ndiffusion >>
rect 21 14 23 54
rect 27 14 33 54
rect 37 14 39 54
rect 79 48 93 54
rect 63 33 73 34
rect 71 14 73 33
rect 77 14 79 34
rect 91 14 93 48
rect 97 14 99 54
rect 111 14 113 54
rect 117 26 119 54
rect 131 26 133 54
rect 117 14 133 26
rect 137 50 143 54
rect 137 46 151 50
rect 137 18 139 46
rect 137 14 151 18
rect 171 14 173 34
rect 177 14 179 34
<< pdiffusion >>
rect 21 206 23 246
rect 27 214 29 246
rect 41 214 43 246
rect 27 206 43 214
rect 47 206 49 246
rect 81 206 83 246
rect 87 206 89 246
rect 101 206 103 246
rect 107 206 109 246
rect 121 166 123 246
rect 127 166 133 246
rect 137 166 139 246
rect 171 206 173 246
rect 177 206 179 246
<< ndcontact >>
rect 9 14 21 54
rect 39 14 51 54
rect 59 14 71 33
rect 79 14 91 48
rect 99 14 111 54
rect 119 26 131 54
rect 139 18 151 46
rect 159 14 171 34
rect 179 14 191 34
<< pdcontact >>
rect 9 206 21 246
rect 29 214 41 246
rect 49 206 61 246
rect 69 206 81 246
rect 89 206 101 246
rect 109 166 121 246
rect 139 166 151 246
rect 159 206 171 246
rect 179 206 191 246
<< psubstratepcontact >>
rect -6 -6 206 6
<< nsubstratencontact >>
rect -6 254 206 266
<< polysilicon >>
rect 23 246 27 250
rect 43 246 47 250
rect 83 246 87 250
rect 103 246 107 250
rect 123 246 127 250
rect 133 246 137 250
rect 173 246 177 250
rect 23 116 27 206
rect 23 54 27 103
rect 43 99 47 206
rect 83 204 87 206
rect 103 204 107 206
rect 83 200 107 204
rect 42 68 46 87
rect 33 63 46 68
rect 83 66 87 200
rect 173 204 177 206
rect 159 200 177 204
rect 123 162 127 166
rect 113 158 127 162
rect 113 104 117 158
rect 133 152 137 166
rect 133 147 141 152
rect 33 54 37 63
rect 77 60 97 66
rect 93 54 97 60
rect 113 54 117 92
rect 137 83 141 147
rect 159 71 163 200
rect 133 54 137 71
rect 161 59 163 71
rect 73 34 77 54
rect 159 40 163 59
rect 159 36 177 40
rect 173 34 177 36
rect 23 10 27 14
rect 33 10 37 14
rect 73 10 77 14
rect 93 10 97 14
rect 113 10 117 14
rect 133 10 137 14
rect 173 10 177 14
<< polycontact >>
rect 19 103 31 116
rect 42 87 54 99
rect 105 92 117 104
rect 65 54 77 66
rect 129 71 141 83
rect 149 59 161 71
<< metal1 >>
rect -6 266 206 268
rect -6 252 206 254
rect 29 246 41 252
rect 89 246 101 252
rect 139 246 151 252
rect 29 210 41 214
rect 11 204 21 206
rect 49 204 57 206
rect 11 198 57 204
rect 47 119 53 198
rect 69 117 77 206
rect 159 246 171 252
rect 181 200 187 206
rect 171 194 187 200
rect 111 153 117 166
rect 111 147 133 153
rect 19 81 28 103
rect 54 92 105 97
rect 54 91 117 92
rect 124 95 133 147
rect 171 117 177 194
rect 158 103 177 117
rect 124 89 157 95
rect 19 74 129 81
rect 151 71 157 89
rect 53 54 65 66
rect 119 59 149 65
rect 119 54 131 59
rect 59 33 73 34
rect 139 46 151 50
rect 111 18 139 20
rect 171 48 177 103
rect 171 42 187 48
rect 181 34 187 42
rect 111 14 151 18
rect 9 8 21 14
rect 79 8 91 14
rect 159 8 171 14
rect -6 6 206 8
rect -6 -8 206 -6
<< m2contact >>
rect 5 103 19 117
rect 46 105 60 119
rect 66 103 80 117
rect 103 104 117 117
rect 103 103 105 104
rect 105 103 117 104
rect 144 103 158 117
rect 39 54 53 68
rect 59 34 73 48
<< metal2 >>
rect 66 117 74 134
rect 106 117 114 134
rect 6 86 14 103
rect 46 68 53 105
rect 69 48 77 103
rect 146 86 154 103
rect 73 34 77 48
<< m1p >>
rect -6 252 206 268
rect -6 -8 206 8
<< m2p >>
rect 66 119 74 134
rect 106 119 114 134
rect 6 86 14 101
rect 146 86 154 101
<< labels >>
rlabel metal2 10 90 10 90 7 A
port 1 n signal input
rlabel metal2 110 131 110 131 3 B
port 2 n signal input
rlabel metal2 150 90 150 90 3 YS
port 3 n signal output
rlabel metal2 70 131 70 131 7 YC
port 4 n signal output
rlabel metal1 -6 252 206 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 206 8 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 200 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
