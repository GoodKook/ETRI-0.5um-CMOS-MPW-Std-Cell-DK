magic
tech scmos
magscale 1 3
timestamp 1555589239
<< checkpaint >>
rect -50 -50 300 300
<< ndiffusion >>
rect 75 75 175 175
<< psubstratepdiff >>
rect 10 220 240 240
rect 10 30 30 220
rect 220 30 240 220
rect 10 10 240 30
<< metal1 >>
rect 10 220 240 240
rect 10 30 30 220
rect 75 75 175 175
rect 220 30 240 220
rect 10 10 240 30
use ntap_CDNS_7046768260512  ntap_CDNS_7046768260512_0
timestamp 1555589239
transform 1 0 71 0 1 71
box 4 4 104 104
use ptap_CDNS_7046768260511  ptap_CDNS_7046768260511_0
timestamp 1555589239
transform 1 0 216 0 1 26
box 4 4 24 194
use ptap_CDNS_7046768260511  ptap_CDNS_7046768260511_1
timestamp 1555589239
transform 0 1 26 1 0 216
box 4 4 24 194
use ptap_CDNS_7046768260511  ptap_CDNS_7046768260511_2
timestamp 1555589239
transform 0 1 26 1 0 6
box 4 4 24 194
use ptap_CDNS_7046768260511  ptap_CDNS_7046768260511_3
timestamp 1555589239
transform 1 0 6 0 1 26
box 4 4 24 194
<< end >>
