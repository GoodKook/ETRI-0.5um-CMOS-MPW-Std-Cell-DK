magic
tech scmos
magscale 1 3
timestamp 1725348157
<< checkpaint >>
rect -44 432 158 438
rect -58 425 164 432
rect 278 425 454 435
rect -58 158 454 425
rect -58 -36 459 158
rect -55 -38 459 -36
<< nwell >>
rect 110 110 300 300
<< psubstratepdiff >>
rect 45 345 365 365
rect 45 65 65 345
rect 195 195 215 215
rect 345 65 365 345
rect 45 45 365 65
<< nsubstratendiff >>
rect 130 260 280 280
rect 130 150 150 260
rect 260 150 280 260
rect 130 130 280 150
<< genericcontact >>
rect 70 345 340 365
rect 45 75 65 340
rect 150 260 260 280
rect 130 150 150 260
rect 195 195 215 215
rect 260 150 280 260
rect 150 130 260 150
rect 345 70 365 340
rect 70 45 340 65
<< metal1 >>
rect 45 345 365 365
rect 45 65 65 345
rect 130 260 280 280
rect 130 150 150 260
rect 194 194 216 216
rect 260 150 280 260
rect 130 130 280 150
rect 345 65 365 345
rect 45 45 365 65
<< labels >>
rlabel metal1 194 194 216 216 0 EMITTER
port 1 nsew
rlabel metal1 130 260 280 280 0 BASE
port 2 nsew
rlabel metal1 45 345 365 365 0 COLLECTOR
port 3 nsew
<< end >>
