magic
tech scmos
magscale 1 2
timestamp 1702508443
<< nwell >>
rect -12 154 72 272
<< ntransistor >>
rect 18 14 22 34
rect 38 14 42 54
<< ptransistor >>
rect 18 206 22 246
rect 38 166 42 246
<< ndiffusion >>
rect 16 14 18 34
rect 22 14 24 34
rect 36 14 38 54
rect 42 14 44 54
<< pdiffusion >>
rect 16 206 18 246
rect 22 206 24 246
rect 36 178 38 246
rect 24 166 38 178
rect 42 166 44 246
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 54
rect 44 14 56 54
<< pdcontact >>
rect 4 206 16 246
rect 24 178 36 246
rect 44 166 56 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 18 34 22 206
rect 38 160 42 166
rect 38 54 42 60
rect 18 10 22 14
rect 38 10 42 14
<< polycontact >>
rect 6 117 18 129
rect 30 148 42 160
rect 30 60 42 72
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 24 246 36 252
rect 4 160 12 206
rect 4 154 30 160
rect 30 72 36 148
rect 48 117 56 166
rect 4 60 30 66
rect 4 34 12 60
rect 48 54 56 103
rect 24 8 36 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m2contact >>
rect 6 103 20 117
rect 42 103 56 117
<< metal2 >>
rect 46 117 54 134
rect 6 86 14 103
<< m1p >>
rect -6 252 66 268
rect -6 -8 66 8
<< m2p >>
rect 46 119 54 134
rect 6 86 14 101
<< labels >>
rlabel metal2 10 90 10 90 1 A
port 1 n signal input
rlabel metal2 50 130 50 130 5 Y
port 2 n signal output
rlabel metal1 -6 252 66 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 66 8 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
