magic
tech scmos
magscale 1 6
timestamp 1537935238
<< checkpaint >>
rect -184 -162 544 766
<< ntransistor >>
rect 103 480 113 604
rect 221 480 231 604
<< ptransistor >>
rect -17 0 -7 124
rect 43 0 53 124
rect 103 0 113 124
rect 221 0 231 124
rect 281 0 291 124
rect 341 0 351 124
<< ndiffusion >>
rect 60 562 103 604
rect 60 550 72 562
rect 84 550 103 562
rect 60 506 103 550
rect 60 494 72 506
rect 84 494 103 506
rect 60 480 103 494
rect 113 562 156 604
rect 113 550 132 562
rect 144 550 156 562
rect 113 506 156 550
rect 113 494 132 506
rect 144 494 156 506
rect 113 480 156 494
rect 178 562 221 604
rect 178 550 190 562
rect 202 550 221 562
rect 178 506 221 550
rect 178 494 190 506
rect 202 494 221 506
rect 178 480 221 494
rect 231 562 274 604
rect 231 550 250 562
rect 262 550 274 562
rect 231 506 274 550
rect 231 494 250 506
rect 262 494 274 506
rect 231 480 274 494
<< ndcontact >>
rect 72 550 84 562
rect 72 494 84 506
rect 132 550 144 562
rect 132 494 144 506
rect 190 550 202 562
rect 190 494 202 506
rect 250 550 262 562
rect 250 494 262 506
<< psubstratepdiff >>
rect -60 110 -17 124
rect -60 98 -48 110
rect -36 98 -17 110
rect -60 54 -17 98
rect -60 42 -48 54
rect -36 42 -17 54
rect -60 0 -17 42
rect -7 110 43 124
rect -7 98 12 110
rect 24 98 43 110
rect -7 54 43 98
rect -7 42 12 54
rect 24 42 43 54
rect -7 0 43 42
rect 53 110 103 124
rect 53 98 72 110
rect 84 98 103 110
rect 53 54 103 98
rect 53 42 72 54
rect 84 42 103 54
rect 53 0 103 42
rect 113 110 156 124
rect 113 98 132 110
rect 144 98 156 110
rect 113 54 156 98
rect 113 42 132 54
rect 144 42 156 54
rect 113 0 156 42
rect 176 110 221 124
rect 176 98 190 110
rect 202 98 221 110
rect 176 54 221 98
rect 176 42 190 54
rect 202 42 221 54
rect 176 0 221 42
rect 231 110 281 124
rect 231 98 250 110
rect 262 98 281 110
rect 231 54 281 98
rect 231 42 250 54
rect 262 42 281 54
rect 231 0 281 42
rect 291 110 341 124
rect 291 98 310 110
rect 322 98 341 110
rect 291 54 341 98
rect 291 42 310 54
rect 322 42 341 54
rect 291 0 341 42
rect 351 110 394 124
rect 351 98 370 110
rect 382 98 394 110
rect 351 54 394 98
rect 351 42 370 54
rect 382 42 394 54
rect 351 0 394 42
<< psubstratepcontact >>
rect -48 98 -36 110
rect -48 42 -36 54
rect 12 98 24 110
rect 12 42 24 54
rect 72 98 84 110
rect 72 42 84 54
rect 132 98 144 110
rect 132 42 144 54
rect 190 98 202 110
rect 190 42 202 54
rect 250 98 262 110
rect 250 42 262 54
rect 310 98 322 110
rect 310 42 322 54
rect 370 98 382 110
rect 370 42 382 54
<< polysilicon >>
rect 103 604 113 614
rect 221 604 231 614
rect 103 456 113 480
rect 221 456 231 480
rect -17 124 -7 148
rect 43 124 53 148
rect 103 124 113 148
rect 221 124 231 148
rect 281 124 291 148
rect 341 124 351 148
rect -17 -10 -7 0
rect 43 -10 53 0
rect 103 -10 113 0
rect 221 -10 231 0
rect 281 -10 291 0
rect 341 -10 351 0
<< metal1 >>
rect 116 622 276 646
rect 58 562 100 606
rect 58 550 72 562
rect 84 550 100 562
rect 58 506 100 550
rect 58 494 72 506
rect 84 494 100 506
rect 58 478 100 494
rect 116 562 156 622
rect 116 550 132 562
rect 144 550 156 562
rect 116 506 156 550
rect 116 494 132 506
rect 144 494 156 506
rect 116 478 156 494
rect 176 562 218 606
rect 176 550 190 562
rect 202 550 218 562
rect 176 506 218 550
rect 176 494 190 506
rect 202 494 218 506
rect 176 478 218 494
rect 234 562 276 622
rect 234 550 250 562
rect 262 550 276 562
rect 234 506 276 550
rect 234 494 250 506
rect 262 494 276 506
rect 234 478 276 494
rect 62 418 154 462
rect 180 418 272 458
rect -30 146 154 186
rect 179 146 364 186
rect 356 126 398 128
rect -64 110 -20 126
rect -64 98 -48 110
rect -36 98 -20 110
rect -64 54 -20 98
rect -64 42 -48 54
rect -36 42 -20 54
rect -64 -2 -20 42
rect -4 110 40 126
rect -4 98 12 110
rect 24 98 40 110
rect -4 54 40 98
rect -4 42 12 54
rect 24 42 40 54
rect -4 -18 40 42
rect 56 110 100 126
rect 56 98 72 110
rect 84 98 100 110
rect 56 54 100 98
rect 56 42 72 54
rect 84 42 100 54
rect 56 -2 100 42
rect 116 110 158 126
rect 116 98 132 110
rect 144 98 158 110
rect 116 54 158 98
rect 116 42 132 54
rect 144 42 158 54
rect 116 -18 158 42
rect 176 110 218 126
rect 176 98 190 110
rect 202 98 218 110
rect 176 54 218 98
rect 176 42 190 54
rect 202 42 218 54
rect 176 -2 218 42
rect 234 110 276 126
rect 234 98 250 110
rect 262 98 276 110
rect 234 54 276 98
rect 234 42 250 54
rect 262 42 276 54
rect 234 -18 276 42
rect 294 110 338 126
rect 294 98 310 110
rect 322 98 338 110
rect 294 54 338 98
rect 294 42 310 54
rect 322 42 338 54
rect 294 -2 338 42
rect 354 110 398 126
rect 354 98 370 110
rect 382 98 398 110
rect 354 54 398 98
rect 354 42 370 54
rect 382 42 398 54
rect 354 -18 398 42
rect -4 -42 398 -18
<< metal2 >>
rect 58 478 98 606
rect 176 478 216 606
rect 236 519 276 606
rect 236 478 424 519
rect 62 418 154 458
rect 180 418 272 458
rect 116 186 154 418
rect 232 186 272 418
rect -30 146 154 186
rect 179 146 364 186
rect 384 126 424 478
rect -62 -2 -22 126
rect 58 -2 98 126
rect 176 -2 424 126
<< metal3 >>
rect 58 478 98 606
rect 176 478 216 606
rect -62 -2 -22 126
rect 58 -2 98 126
rect 176 -2 218 126
rect 296 -2 336 126
use CONT  CONT_0
timestamp 1537935238
transform 1 0 138 0 1 528
box -6 -6 6 6
use CONT  CONT_1
timestamp 1537935238
transform -1 0 256 0 -1 76
box -6 -6 6 6
use CONT  CONT_2
timestamp 1537935238
transform 1 0 138 0 1 584
box -6 -6 6 6
use CONT  CONT_3
timestamp 1537935238
transform -1 0 256 0 -1 20
box -6 -6 6 6
use CONT  CONT_4
timestamp 1537935238
transform -1 0 138 0 -1 76
box -6 -6 6 6
use CONT  CONT_5
timestamp 1537935238
transform -1 0 138 0 -1 20
box -6 -6 6 6
use CONT  CONT_6
timestamp 1537935238
transform -1 0 18 0 -1 20
box -6 -6 6 6
use CONT  CONT_7
timestamp 1537935238
transform -1 0 18 0 -1 76
box -6 -6 6 6
use CONT  CONT_8
timestamp 1537935238
transform -1 0 376 0 -1 76
box -6 -6 6 6
use CONT  CONT_9
timestamp 1537935238
transform -1 0 376 0 -1 20
box -6 -6 6 6
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_0
timestamp 1537935238
transform -1 0 126 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_1
timestamp 1537935238
transform 1 0 268 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_2
timestamp 1537935238
transform 1 0 208 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_3
timestamp 1537935238
transform -1 0 244 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_4
timestamp 1537935238
transform 1 0 90 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_5
timestamp 1537935238
transform 1 0 -30 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_6
timestamp 1537935238
transform 1 0 30 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_7
timestamp 1537935238
transform 1 0 328 0 1 146
box 0 0 36 36
use VIA1  VIA1_0
timestamp 1537935238
transform 1 0 199 0 1 166
box -8 -8 8 8
use VIA1  VIA1_1
timestamp 1537935238
transform 1 0 78 0 1 528
box -8 -8 8 8
use VIA1  VIA1_2
timestamp 1537935238
transform 1 0 78 0 1 584
box -8 -8 8 8
use VIA1  VIA1_3
timestamp 1537935238
transform 1 0 200 0 1 438
box -8 -8 8 8
use VIA1  VIA1_4
timestamp 1537935238
transform -1 0 316 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_5
timestamp 1537935238
transform 1 0 134 0 1 438
box -8 -8 8 8
use VIA1  VIA1_6
timestamp 1537935238
transform 1 0 134 0 1 166
box -8 -8 8 8
use VIA1  VIA1_7
timestamp 1537935238
transform 1 0 256 0 1 166
box -8 -8 8 8
use VIA1  VIA1_8
timestamp 1537935238
transform 1 0 252 0 1 438
box -8 -8 8 8
use VIA1  VIA1_9
timestamp 1537935238
transform 1 0 316 0 1 166
box -8 -8 8 8
use VIA1  VIA1_10
timestamp 1537935238
transform 1 0 78 0 1 166
box -8 -8 8 8
use VIA1  VIA1_11
timestamp 1537935238
transform 1 0 82 0 1 438
box -8 -8 8 8
use VIA1  VIA1_12
timestamp 1537935238
transform -1 0 196 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_13
timestamp 1537935238
transform -1 0 196 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_14
timestamp 1537935238
transform -1 0 78 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_15
timestamp 1537935238
transform -1 0 78 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_16
timestamp 1537935238
transform -1 0 -42 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_17
timestamp 1537935238
transform 1 0 196 0 1 528
box -8 -8 8 8
use VIA1  VIA1_18
timestamp 1537935238
transform 1 0 18 0 1 166
box -8 -8 8 8
use VIA1  VIA1_19
timestamp 1537935238
transform -1 0 -42 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_20
timestamp 1537935238
transform -1 0 316 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_21
timestamp 1537935238
transform 1 0 196 0 1 584
box -8 -8 8 8
use VIA1  VIA1_22
timestamp 1537935238
transform 1 0 256 0 1 528
box -8 -8 8 8
use VIA1  VIA1_23
timestamp 1537935238
transform 1 0 256 0 1 584
box -8 -8 8 8
use VIA2  VIA2_0
timestamp 1537935238
transform 1 0 78 0 1 500
box -8 -8 8 8
use VIA2  VIA2_1
timestamp 1537935238
transform 1 0 78 0 1 556
box -8 -8 8 8
use VIA2  VIA2_2
timestamp 1537935238
transform 1 0 196 0 1 556
box -8 -8 8 8
use VIA2  VIA2_3
timestamp 1537935238
transform -1 0 78 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_4
timestamp 1537935238
transform -1 0 78 0 -1 104
box -8 -8 8 8
use VIA2  VIA2_5
timestamp 1537935238
transform -1 0 -42 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_6
timestamp 1537935238
transform -1 0 -42 0 -1 104
box -8 -8 8 8
use VIA2  VIA2_7
timestamp 1537935238
transform 1 0 196 0 1 500
box -8 -8 8 8
<< end >>
