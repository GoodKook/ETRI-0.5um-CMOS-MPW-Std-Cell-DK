magic
tech scmos
magscale 1 6
timestamp 1555589239
<< checkpaint >>
rect -122 -162 546 766
<< ntransistor >>
rect 103 480 113 604
rect 221 480 231 604
rect 339 480 349 604
<< ptransistor >>
rect 43 0 53 124
rect 103 0 113 124
rect 163 0 173 124
rect 223 0 233 124
rect 283 0 293 124
rect 343 0 353 124
<< ndiffusion >>
rect 60 562 103 604
rect 60 550 72 562
rect 84 550 103 562
rect 60 506 103 550
rect 60 494 72 506
rect 84 494 103 506
rect 60 480 103 494
rect 113 562 156 604
rect 113 550 132 562
rect 144 550 156 562
rect 113 506 156 550
rect 113 494 132 506
rect 144 494 156 506
rect 113 480 156 494
rect 178 562 221 604
rect 178 550 190 562
rect 202 550 221 562
rect 178 506 221 550
rect 178 494 190 506
rect 202 494 221 506
rect 178 480 221 494
rect 231 562 274 604
rect 231 550 250 562
rect 262 550 274 562
rect 231 506 274 550
rect 231 494 250 506
rect 262 494 274 506
rect 231 480 274 494
rect 296 562 339 604
rect 296 550 308 562
rect 320 550 339 562
rect 296 506 339 550
rect 296 494 308 506
rect 320 494 339 506
rect 296 480 339 494
rect 349 562 392 604
rect 349 550 368 562
rect 380 550 392 562
rect 349 506 392 550
rect 349 494 368 506
rect 380 494 392 506
rect 349 480 392 494
<< ndcontact >>
rect 72 550 84 562
rect 72 494 84 506
rect 132 550 144 562
rect 132 494 144 506
rect 190 550 202 562
rect 190 494 202 506
rect 250 550 262 562
rect 250 494 262 506
rect 308 550 320 562
rect 308 494 320 506
rect 368 550 380 562
rect 368 494 380 506
<< psubstratepdiff >>
rect 0 110 43 124
rect 0 98 12 110
rect 24 98 43 110
rect 0 54 43 98
rect 0 42 12 54
rect 24 42 43 54
rect 0 0 43 42
rect 53 110 103 124
rect 53 98 72 110
rect 84 98 103 110
rect 53 54 103 98
rect 53 42 72 54
rect 84 42 103 54
rect 53 0 103 42
rect 113 110 163 124
rect 113 98 132 110
rect 144 98 163 110
rect 113 54 163 98
rect 113 42 132 54
rect 144 42 163 54
rect 113 0 163 42
rect 173 110 223 124
rect 173 98 192 110
rect 204 98 223 110
rect 173 54 223 98
rect 173 42 192 54
rect 204 42 223 54
rect 173 0 223 42
rect 233 110 283 124
rect 233 98 252 110
rect 264 98 283 110
rect 233 54 283 98
rect 233 42 252 54
rect 264 42 283 54
rect 233 0 283 42
rect 293 110 343 124
rect 293 98 312 110
rect 324 98 343 110
rect 293 54 343 98
rect 293 42 312 54
rect 324 42 343 54
rect 293 0 343 42
rect 353 110 396 124
rect 353 98 372 110
rect 384 98 396 110
rect 353 54 396 98
rect 353 42 372 54
rect 384 42 396 54
rect 353 0 396 42
<< psubstratepcontact >>
rect 12 98 24 110
rect 12 42 24 54
rect 72 98 84 110
rect 72 42 84 54
rect 132 98 144 110
rect 132 42 144 54
rect 192 98 204 110
rect 192 42 204 54
rect 252 98 264 110
rect 252 42 264 54
rect 312 98 324 110
rect 312 42 324 54
rect 372 98 384 110
rect 372 42 384 54
<< polysilicon >>
rect 103 604 113 614
rect 221 604 231 614
rect 339 604 349 614
rect 103 456 113 480
rect 221 456 231 480
rect 339 456 349 480
rect 43 124 53 148
rect 103 124 113 148
rect 163 124 173 148
rect 223 124 233 148
rect 283 124 293 148
rect 343 124 353 148
rect 43 -10 53 0
rect 103 -10 113 0
rect 163 -10 173 0
rect 223 -10 233 0
rect 283 -10 293 0
rect 343 -10 353 0
<< metal1 >>
rect 116 622 394 646
rect 58 562 100 606
rect 58 550 72 562
rect 84 550 100 562
rect 58 506 100 550
rect 58 494 72 506
rect 84 494 100 506
rect 58 478 100 494
rect 116 562 158 622
rect 116 550 132 562
rect 144 550 158 562
rect 116 506 158 550
rect 116 494 132 506
rect 144 494 158 506
rect 116 478 158 494
rect 176 562 218 606
rect 176 550 190 562
rect 202 550 218 562
rect 176 506 218 550
rect 176 494 190 506
rect 202 494 218 506
rect 176 478 218 494
rect 234 562 276 622
rect 234 550 250 562
rect 262 550 276 562
rect 234 506 276 550
rect 234 494 250 506
rect 262 494 276 506
rect 234 478 276 494
rect 294 562 336 606
rect 294 550 308 562
rect 320 550 336 562
rect 294 506 336 550
rect 294 494 308 506
rect 320 494 336 506
rect 294 478 336 494
rect 352 562 394 622
rect 352 550 368 562
rect 380 550 394 562
rect 352 506 394 550
rect 352 494 368 506
rect 380 494 394 506
rect 352 478 394 494
rect 90 418 362 462
rect 30 146 366 186
rect -2 110 40 126
rect -2 98 12 110
rect 24 98 40 110
rect -2 54 40 98
rect -2 42 12 54
rect 24 42 40 54
rect -2 -18 40 42
rect 56 110 100 126
rect 56 98 72 110
rect 84 98 100 110
rect 56 54 100 98
rect 56 42 72 54
rect 84 42 100 54
rect 56 -2 100 42
rect 116 110 158 126
rect 116 98 132 110
rect 144 98 158 110
rect 116 54 158 98
rect 116 42 132 54
rect 144 42 158 54
rect 116 -2 158 42
rect 176 110 220 126
rect 176 98 192 110
rect 204 98 220 110
rect 176 54 220 98
rect 176 42 192 54
rect 204 42 220 54
rect 176 -2 220 42
rect 236 110 278 126
rect 236 98 252 110
rect 264 98 278 110
rect 236 54 278 98
rect 236 42 252 54
rect 264 42 278 54
rect 236 -2 278 42
rect 296 110 340 126
rect 296 98 312 110
rect 324 98 340 110
rect 296 54 340 98
rect 296 42 312 54
rect 324 42 340 54
rect 296 -2 340 42
rect 356 110 398 126
rect 356 98 372 110
rect 384 98 398 110
rect 356 54 398 98
rect 356 42 372 54
rect 384 42 398 54
rect 116 -18 160 -2
rect 236 -18 280 -2
rect 356 -18 398 42
rect -2 -42 398 -18
<< metal2 >>
rect 58 478 98 606
rect 176 478 216 606
rect 294 478 334 606
rect 354 478 426 606
rect 90 418 362 458
rect 184 186 212 418
rect 30 146 366 186
rect 386 126 426 478
rect 58 -2 98 126
rect 178 -2 218 126
rect 298 -2 338 126
rect 358 -2 426 126
<< metal3 >>
rect 58 478 98 606
rect 176 478 216 606
rect 294 478 334 606
rect 58 -2 98 126
rect 178 -2 218 126
rect 298 -2 338 126
use CONT  CONT_0
timestamp 1555589239
transform -1 0 18 0 -1 76
box -6 -6 6 6
use CONT  CONT_1
timestamp 1555589239
transform 1 0 138 0 1 528
box -6 -6 6 6
use CONT  CONT_2
timestamp 1555589239
transform -1 0 18 0 -1 20
box -6 -6 6 6
use CONT  CONT_3
timestamp 1555589239
transform 1 0 138 0 1 584
box -6 -6 6 6
use CONT  CONT_4
timestamp 1555589239
transform -1 0 258 0 -1 76
box -6 -6 6 6
use CONT  CONT_5
timestamp 1555589239
transform -1 0 258 0 -1 20
box -6 -6 6 6
use CONT  CONT_6
timestamp 1555589239
transform -1 0 138 0 -1 20
box -6 -6 6 6
use CONT  CONT_7
timestamp 1555589239
transform -1 0 138 0 -1 76
box -6 -6 6 6
use CONT  CONT_8
timestamp 1555589239
transform 1 0 256 0 1 528
box -6 -6 6 6
use CONT  CONT_9
timestamp 1555589239
transform 1 0 256 0 1 584
box -6 -6 6 6
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_0
timestamp 1555589239
transform 1 0 90 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_1
timestamp 1555589239
transform -1 0 126 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_2
timestamp 1555589239
transform 1 0 30 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_3
timestamp 1555589239
transform 1 0 210 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_4
timestamp 1555589239
transform 1 0 150 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_5
timestamp 1555589239
transform 1 0 330 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_6
timestamp 1555589239
transform 1 0 270 0 1 146
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_7
timestamp 1555589239
transform -1 0 244 0 -1 458
box 0 0 36 36
use poly1cont_CDNS_704676826053  poly1cont_CDNS_704676826053_8
timestamp 1555589239
transform -1 0 362 0 -1 458
box 0 0 36 36
use VIA1  VIA1_0
timestamp 1555589239
transform 1 0 78 0 1 528
box -8 -8 8 8
use VIA1  VIA1_1
timestamp 1555589239
transform 1 0 78 0 1 584
box -8 -8 8 8
use VIA1  VIA1_2
timestamp 1555589239
transform 1 0 138 0 1 166
box -8 -8 8 8
use VIA1  VIA1_3
timestamp 1555589239
transform 1 0 258 0 1 166
box -8 -8 8 8
use VIA1  VIA1_4
timestamp 1555589239
transform -1 0 78 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_5
timestamp 1555589239
transform 1 0 78 0 1 166
box -8 -8 8 8
use VIA1  VIA1_6
timestamp 1555589239
transform 1 0 146 0 1 438
box -8 -8 8 8
use VIA1  VIA1_7
timestamp 1555589239
transform -1 0 78 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_8
timestamp 1555589239
transform 1 0 182 0 1 438
box -8 -8 8 8
use VIA1  VIA1_9
timestamp 1555589239
transform 1 0 266 0 1 438
box -8 -8 8 8
use VIA1  VIA1_10
timestamp 1555589239
transform 1 0 302 0 1 438
box -8 -8 8 8
use VIA1  VIA1_11
timestamp 1555589239
transform 1 0 198 0 1 166
box -8 -8 8 8
use VIA1  VIA1_12
timestamp 1555589239
transform 1 0 320 0 1 166
box -8 -8 8 8
use VIA1  VIA1_13
timestamp 1555589239
transform -1 0 198 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_14
timestamp 1555589239
transform -1 0 198 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_15
timestamp 1555589239
transform -1 0 378 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_16
timestamp 1555589239
transform -1 0 378 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_17
timestamp 1555589239
transform -1 0 318 0 -1 76
box -8 -8 8 8
use VIA1  VIA1_18
timestamp 1555589239
transform -1 0 318 0 -1 20
box -8 -8 8 8
use VIA1  VIA1_19
timestamp 1555589239
transform 1 0 196 0 1 528
box -8 -8 8 8
use VIA1  VIA1_20
timestamp 1555589239
transform 1 0 196 0 1 584
box -8 -8 8 8
use VIA1  VIA1_21
timestamp 1555589239
transform 1 0 314 0 1 528
box -8 -8 8 8
use VIA1  VIA1_22
timestamp 1555589239
transform 1 0 314 0 1 584
box -8 -8 8 8
use VIA1  VIA1_23
timestamp 1555589239
transform 1 0 374 0 1 528
box -8 -8 8 8
use VIA1  VIA1_24
timestamp 1555589239
transform 1 0 374 0 1 584
box -8 -8 8 8
use VIA2  VIA2_0
timestamp 1555589239
transform 1 0 78 0 1 500
box -8 -8 8 8
use VIA2  VIA2_1
timestamp 1555589239
transform -1 0 78 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_2
timestamp 1555589239
transform 1 0 78 0 1 556
box -8 -8 8 8
use VIA2  VIA2_3
timestamp 1555589239
transform -1 0 78 0 -1 104
box -8 -8 8 8
use VIA2  VIA2_4
timestamp 1555589239
transform 1 0 314 0 1 500
box -8 -8 8 8
use VIA2  VIA2_5
timestamp 1555589239
transform 1 0 196 0 1 500
box -8 -8 8 8
use VIA2  VIA2_6
timestamp 1555589239
transform -1 0 198 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_7
timestamp 1555589239
transform -1 0 198 0 -1 104
box -8 -8 8 8
use VIA2  VIA2_8
timestamp 1555589239
transform -1 0 318 0 -1 48
box -8 -8 8 8
use VIA2  VIA2_9
timestamp 1555589239
transform -1 0 318 0 -1 104
box -8 -8 8 8
use VIA2  VIA2_10
timestamp 1555589239
transform 1 0 196 0 1 556
box -8 -8 8 8
use VIA2  VIA2_11
timestamp 1555589239
transform 1 0 314 0 1 556
box -8 -8 8 8
<< end >>
