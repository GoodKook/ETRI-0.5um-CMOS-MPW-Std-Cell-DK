#--------------------------------------------------
# LEF file for Route & Via Rile
#  Ported from osu050 by GoodKook@gmail.com
#

VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;

UNITS
  DATABASE MICRONS 1000 ;
END UNITS

USEMINSPACING OBS ON ;
USEMINSPACING PIN OFF ;
CLEARANCEMEASURE EUCLIDEAN ;

MANUFACTURINGGRID 0.15 ;

LAYER nwell
  TYPE	MASTERSLICE ;
END nwell

LAYER nactive
  TYPE	MASTERSLICE ;
END nactive

LAYER pactive
  TYPE	MASTERSLICE ;
END pactive

LAYER poly
  TYPE	MASTERSLICE ;
END poly

LAYER cc
  TYPE	CUT ;
  SPACING	0.9 ;
END cc

LAYER metal1
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH	    0.9 ;   # ETRI050 Rule: WIDTH=0.8
  SPACING	1.05 ;  # ETRI050 Rule: SPACING=1.0
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 3.2e-05 ;
END metal1

LAYER via1
  TYPE	CUT ;
  SPACING	0.9 ;
END via1

LAYER metal2
  TYPE		ROUTING ;
  DIRECTION	VERTICAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.05 ;  # ETRI050 Rule: WIDTH=1.0
  SPACING	1.05 ;  # ETRI050 Rule: SPACING=1.0
  RESISTANCE	RPERSQ 0.09 ;
  CAPACITANCE	CPERSQDIST 1.6e-05 ;
END metal2

LAYER via2
  TYPE	CUT ;
  SPACING	0.9 ;
END via2

LAYER metal3
  TYPE		ROUTING ;
  DIRECTION	HORIZONTAL ;
  PITCH		3.0 ;
  OFFSET	1.5 ;
  WIDTH		1.2 ;   # ETRI050 Rule: WIDTH=1.2
  SPACING	1.05 ;  # ETRI050 Rule: SPACING=1.0
  RESISTANCE	RPERSQ 0.05 ;
  CAPACITANCE	CPERSQDIST 1e-05 ;
END metal3

SPACING
  SAMENET cc   via1	0.900 ;
  SAMENET via1 via2	0.900 ;
END SPACING

VIA M2_M1 DEFAULT
  LAYER metal1 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via1 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M2_M1

VIA M3_M2 DEFAULT
  LAYER metal2 ;
    RECT -1.050 -1.050 1.050 1.050 ;
  LAYER via2 ;
    RECT -0.450 -0.450 0.450 0.450 ;
  LAYER metal3 ;
    RECT -1.050 -1.050 1.050 1.050 ;
END M3_M2


VIARULE viagen21 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via1 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
    WIDTH 2.1 TO 210 ;
    OVERHANG 0.0 ;
    METALOVERHANG 0 ;
  LAYER via2 ;
#    RECT -1.05 -1.05 1.05 1.05 ;
    RECT -0.450 -0.450 0.450 0.450 ;
    SPACING 0.9 BY 0.9 ;
END viagen32

VIARULE TURN1 GENERATE
  LAYER metal1 ;
    DIRECTION HORIZONTAL ;
  LAYER metal1 ;
    DIRECTION VERTICAL ;
END TURN1

VIARULE TURN2 GENERATE
  LAYER metal2 ;
    DIRECTION HORIZONTAL ;
  LAYER metal2 ;
    DIRECTION VERTICAL ;
END TURN2

VIARULE TURN3 GENERATE
  LAYER metal3 ;
    DIRECTION HORIZONTAL ;
  LAYER metal3 ;
    DIRECTION VERTICAL ;
END TURN3

SITE  corner
    CLASS	PAD ;
    SYMMETRY	R90 Y ;
    SIZE	300.000 BY 300.000 ;
END  corner

SITE  IO
    CLASS	PAD ;
    SYMMETRY	Y ;
    SIZE	90.000 BY 300.000 ;
END  IO

SITE  core
    CLASS	CORE ;
    SYMMETRY	Y ;
    SIZE	3.000 BY 30.000 ;
END  core

# =====================================================================
#  Core MACROS
# =====================================================================
MACRO AND2X1
  CLASS CORE ;
  FOREIGN AND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 30.900 2.400 37.500 ;
        RECT 3.600 30.900 5.400 36.900 ;
        RECT 6.600 30.900 8.400 37.500 ;
        RECT 9.600 30.900 11.400 36.900 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 3.600 10.800 4.500 30.900 ;
        RECT 9.900 20.850 11.100 30.900 ;
        RECT 6.450 14.550 7.800 15.150 ;
        RECT 5.700 12.750 7.800 14.550 ;
        RECT 0.600 9.600 9.000 10.800 ;
        RECT 0.600 2.100 2.400 9.600 ;
        RECT 7.200 9.000 9.000 9.600 ;
        RECT 5.100 1.500 6.900 8.100 ;
        RECT 9.900 6.000 11.100 18.150 ;
        RECT 8.100 5.100 11.100 6.000 ;
        RECT 8.100 2.100 9.900 5.100 ;
  END
END AND2X1
MACRO AND2X2
  CLASS CORE ;
  FOREIGN AND2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 30.900 2.400 37.500 ;
        RECT 3.600 30.900 5.400 36.900 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.600 10.800 4.500 30.900 ;
        RECT 6.600 24.900 8.400 37.500 ;
        RECT 9.600 24.900 11.400 36.900 ;
        RECT 9.900 20.850 11.100 24.900 ;
        RECT 6.450 14.550 7.800 15.150 ;
        RECT 5.700 12.750 7.800 14.550 ;
        RECT 0.600 9.900 9.000 10.800 ;
        RECT 0.600 2.100 2.400 9.900 ;
        RECT 7.200 9.000 9.000 9.900 ;
        RECT 9.900 8.100 11.100 18.150 ;
        RECT 5.100 1.500 6.900 8.100 ;
        RECT 8.100 6.000 11.100 8.100 ;
        RECT 8.100 2.100 9.900 6.000 ;
  END
END AND2X2
MACRO AOI21X1
  CLASS CORE ;
  FOREIGN AOI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
        RECT 3.600 26.700 5.400 37.800 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT 1.500 1.200 3.300 8.100 ;
        RECT 9.000 1.200 10.800 5.100 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 25.800 2.400 36.900 ;
        RECT 6.600 25.800 8.400 36.900 ;
        RECT 0.600 24.900 8.400 25.800 ;
        RECT 9.600 24.900 11.400 36.900 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 6.600 15.750 8.400 18.150 ;
        RECT 9.750 17.850 10.950 24.900 ;
        RECT 3.750 12.750 5.550 15.150 ;
        RECT 9.750 8.100 10.950 15.150 ;
        RECT 6.000 7.050 10.950 8.100 ;
        RECT 6.000 2.100 7.800 7.050 ;
  END
END AOI21X1
MACRO AOI22X1
  CLASS CORE ;
  FOREIGN AOI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 26.250 2.400 36.900 ;
        RECT 3.600 27.150 5.400 37.500 ;
        RECT 6.600 36.000 14.400 36.900 ;
        RECT 6.600 26.250 8.400 36.000 ;
        RECT 0.600 25.350 8.400 26.250 ;
        RECT 9.600 24.150 11.400 35.100 ;
        RECT 12.600 24.900 14.400 36.000 ;
        RECT 6.900 23.250 11.400 24.150 ;
        RECT 6.900 20.850 8.100 23.250 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 14.550 5.550 15.150 ;
        RECT 3.900 12.750 5.700 14.550 ;
        RECT 6.600 8.100 7.500 18.150 ;
        RECT 12.450 15.300 14.250 18.150 ;
        RECT 9.450 14.100 11.100 15.150 ;
        RECT 8.700 12.300 11.100 14.100 ;
        RECT 1.200 1.500 3.000 8.100 ;
        RECT 5.700 2.100 7.500 8.100 ;
        RECT 10.200 1.500 12.000 8.100 ;
  END
END AOI22X1
MACRO BUFX2
  CLASS CORE ;
  FOREIGN BUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 9.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 30.900 2.400 36.900 ;
        RECT 0.600 24.150 1.800 30.900 ;
        RECT 3.600 26.700 5.400 37.500 ;
        RECT 6.600 25.050 8.400 36.900 ;
        RECT 0.600 23.100 6.300 24.150 ;
        RECT 4.500 22.350 6.300 23.100 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 4.500 10.800 5.550 22.350 ;
        RECT 7.200 20.850 8.400 25.050 ;
        RECT 4.500 10.200 6.300 10.800 ;
        RECT 0.600 9.000 6.300 10.200 ;
        RECT 0.600 5.100 1.800 9.000 ;
        RECT 7.200 8.100 8.400 18.150 ;
        RECT 0.600 2.100 2.400 5.100 ;
        RECT 3.600 1.500 5.400 8.100 ;
        RECT 6.600 2.100 8.400 8.100 ;
  END
END BUFX2
MACRO BUFX4
  CLASS CORE ;
  FOREIGN BUFX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 27.900 2.400 36.900 ;
        RECT 0.600 24.300 1.800 27.900 ;
        RECT 3.600 25.200 5.400 37.500 ;
        RECT 6.600 25.200 8.400 36.900 ;
        RECT 0.600 23.400 5.550 24.300 ;
        RECT 4.500 23.250 5.550 23.400 ;
        RECT 7.350 24.000 8.400 25.200 ;
        RECT 9.600 24.900 11.400 37.500 ;
        RECT 4.500 21.450 6.300 23.250 ;
        RECT 7.350 23.100 11.100 24.000 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 4.650 10.800 5.550 21.450 ;
        RECT 9.900 20.850 11.100 23.100 ;
        RECT 4.650 9.900 6.450 10.800 ;
        RECT 9.900 10.200 11.100 18.150 ;
        RECT 0.600 9.000 6.450 9.900 ;
        RECT 7.350 9.000 11.100 10.200 ;
        RECT 0.600 6.600 1.800 9.000 ;
        RECT 7.350 8.100 8.400 9.000 ;
        RECT 0.600 2.100 2.400 6.600 ;
        RECT 3.600 1.500 5.400 8.100 ;
        RECT 6.600 2.100 8.400 8.100 ;
        RECT 9.600 1.500 11.400 8.100 ;
  END
END BUFX4
MACRO CLKBUF1
  CLASS CORE ;
  FOREIGN CLKBUF1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 27.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.450 18.450 26.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 27.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 27.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.000 5.400 36.900 ;
        RECT 6.600 24.900 8.400 37.500 ;
        RECT 9.600 24.000 11.400 36.900 ;
        RECT 12.600 24.900 14.400 37.500 ;
        RECT 15.600 24.000 17.400 36.900 ;
        RECT 18.600 24.900 20.400 37.500 ;
        RECT 21.600 24.000 23.400 36.900 ;
        RECT 24.600 24.900 26.400 37.500 ;
        RECT 3.600 22.800 6.900 24.000 ;
        RECT 9.600 22.800 13.500 24.000 ;
        RECT 15.600 22.800 19.500 24.000 ;
        RECT 21.600 22.800 26.100 24.000 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 5.700 17.400 6.900 22.800 ;
        RECT 8.700 17.400 10.500 18.000 ;
        RECT 5.700 16.200 10.500 17.400 ;
        RECT 12.300 17.400 13.500 22.800 ;
        RECT 14.700 17.400 16.500 18.000 ;
        RECT 12.300 16.200 16.500 17.400 ;
        RECT 18.300 17.400 19.500 22.800 ;
        RECT 24.750 20.850 26.100 22.800 ;
        RECT 20.700 17.400 22.500 18.000 ;
        RECT 18.300 16.200 22.500 17.400 ;
        RECT 5.700 10.200 6.900 16.200 ;
        RECT 12.300 10.200 13.500 16.200 ;
        RECT 18.300 10.200 19.500 16.200 ;
        RECT 24.750 10.200 26.100 18.150 ;
        RECT 3.600 9.000 6.900 10.200 ;
        RECT 9.600 9.000 13.500 10.200 ;
        RECT 15.600 9.000 19.500 10.200 ;
        RECT 21.600 9.000 26.100 10.200 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 9.000 ;
        RECT 6.600 1.500 8.400 8.100 ;
        RECT 9.600 2.100 11.400 9.000 ;
        RECT 12.600 1.500 14.400 8.100 ;
        RECT 15.600 2.100 17.400 9.000 ;
        RECT 18.600 1.500 20.400 8.100 ;
        RECT 21.600 2.100 23.400 9.000 ;
        RECT 24.600 1.500 26.400 8.100 ;
  END
END CLKBUF1
MACRO CLKBUF2
  CLASS CORE ;
  FOREIGN CLKBUF2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 39.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 36.450 18.450 38.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 39.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 39.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.000 5.400 36.900 ;
        RECT 6.600 24.900 8.400 37.500 ;
        RECT 9.600 24.000 11.400 36.900 ;
        RECT 12.600 24.900 14.400 37.500 ;
        RECT 15.600 24.000 17.400 36.900 ;
        RECT 18.600 24.900 20.400 37.500 ;
        RECT 21.600 24.000 23.400 36.900 ;
        RECT 24.600 24.900 26.400 37.500 ;
        RECT 27.600 24.000 29.400 36.900 ;
        RECT 30.600 24.900 32.400 37.500 ;
        RECT 33.600 24.000 35.400 36.900 ;
        RECT 36.600 24.900 38.400 37.500 ;
        RECT 3.600 22.800 6.900 24.000 ;
        RECT 9.600 22.800 13.500 24.000 ;
        RECT 15.600 22.800 19.500 24.000 ;
        RECT 21.600 22.800 25.800 24.000 ;
        RECT 27.600 22.800 30.900 24.000 ;
        RECT 33.600 22.800 38.100 24.000 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 5.700 17.700 6.900 22.800 ;
        RECT 8.700 17.700 10.500 18.300 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 5.700 16.500 10.500 17.700 ;
        RECT 12.300 17.700 13.500 22.800 ;
        RECT 14.700 17.700 16.500 18.300 ;
        RECT 12.300 16.500 16.500 17.700 ;
        RECT 18.300 17.700 19.500 22.800 ;
        RECT 20.700 17.700 22.500 18.300 ;
        RECT 18.300 16.500 22.500 17.700 ;
        RECT 24.600 17.700 25.800 22.800 ;
        RECT 26.700 17.700 28.500 18.300 ;
        RECT 24.600 16.500 28.500 17.700 ;
        RECT 29.700 17.700 30.900 22.800 ;
        RECT 36.900 20.850 38.100 22.800 ;
        RECT 32.700 17.700 34.500 18.300 ;
        RECT 29.700 16.500 34.500 17.700 ;
        RECT 5.700 10.200 6.900 16.500 ;
        RECT 12.300 10.200 13.500 16.500 ;
        RECT 18.300 10.200 19.500 16.500 ;
        RECT 24.600 10.200 25.800 16.500 ;
        RECT 29.700 10.200 30.900 16.500 ;
        RECT 36.900 10.200 38.100 18.150 ;
        RECT 3.600 9.000 6.900 10.200 ;
        RECT 9.600 9.000 13.500 10.200 ;
        RECT 15.600 9.000 19.500 10.200 ;
        RECT 21.600 9.000 25.800 10.200 ;
        RECT 27.600 9.000 30.900 10.200 ;
        RECT 33.600 9.000 38.100 10.200 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 9.000 ;
        RECT 6.600 1.500 8.400 8.100 ;
        RECT 9.600 2.100 11.400 9.000 ;
        RECT 12.600 1.500 14.400 8.100 ;
        RECT 15.600 2.100 17.400 9.000 ;
        RECT 18.600 1.500 20.400 8.100 ;
        RECT 21.600 2.100 23.400 9.000 ;
        RECT 24.600 1.500 26.400 8.100 ;
        RECT 27.600 2.100 29.400 9.000 ;
        RECT 30.600 1.500 32.400 8.100 ;
        RECT 33.600 2.100 35.400 9.000 ;
        RECT 36.600 1.500 38.400 8.100 ;
  END
END CLKBUF2
MACRO CLKBUF3
  CLASS CORE ;
  FOREIGN CLKBUF3 ;
  ORIGIN 0.000 0.000 ;
  SIZE 51.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 45.450 18.450 47.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 51.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 51.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.000 5.400 36.900 ;
        RECT 6.600 24.900 8.400 37.500 ;
        RECT 9.600 24.000 11.400 36.900 ;
        RECT 12.600 24.900 14.400 37.500 ;
        RECT 15.600 24.000 17.400 36.900 ;
        RECT 18.600 24.900 20.400 37.500 ;
        RECT 21.600 24.000 23.400 36.900 ;
        RECT 24.600 24.900 26.400 37.500 ;
        RECT 27.600 24.000 29.400 36.900 ;
        RECT 30.600 24.900 32.400 37.500 ;
        RECT 33.600 24.000 35.400 36.900 ;
        RECT 36.600 24.900 38.400 37.500 ;
        RECT 39.600 24.000 41.400 36.900 ;
        RECT 42.600 24.900 44.400 37.500 ;
        RECT 45.600 24.900 47.400 36.900 ;
        RECT 48.600 24.900 50.400 37.500 ;
        RECT 3.600 22.800 7.050 24.000 ;
        RECT 9.600 22.800 13.500 24.000 ;
        RECT 15.600 22.800 19.500 24.000 ;
        RECT 21.600 22.800 25.800 24.000 ;
        RECT 27.600 22.800 30.900 24.000 ;
        RECT 33.600 22.800 37.500 24.000 ;
        RECT 39.600 22.800 43.500 24.000 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 5.850 17.400 7.050 22.800 ;
        RECT 8.700 17.400 10.500 18.000 ;
        RECT 5.850 16.200 10.500 17.400 ;
        RECT 12.300 17.400 13.500 22.800 ;
        RECT 14.700 17.400 16.500 18.000 ;
        RECT 12.300 16.200 16.500 17.400 ;
        RECT 18.300 17.400 19.500 22.800 ;
        RECT 20.700 17.400 22.500 18.000 ;
        RECT 18.300 16.200 22.500 17.400 ;
        RECT 24.600 17.400 25.800 22.800 ;
        RECT 26.700 17.400 28.500 18.000 ;
        RECT 24.600 16.200 28.500 17.400 ;
        RECT 29.700 17.400 30.900 22.800 ;
        RECT 32.700 17.400 34.500 18.000 ;
        RECT 29.700 16.200 34.500 17.400 ;
        RECT 36.300 17.400 37.500 22.800 ;
        RECT 38.700 17.400 40.500 18.000 ;
        RECT 36.300 16.200 40.500 17.400 ;
        RECT 5.850 10.200 7.050 16.200 ;
        RECT 12.300 10.200 13.500 16.200 ;
        RECT 18.300 10.200 19.500 16.200 ;
        RECT 24.600 10.200 25.800 16.200 ;
        RECT 29.700 10.200 30.900 16.200 ;
        RECT 36.300 10.200 37.500 16.200 ;
        RECT 42.300 16.050 43.500 22.800 ;
        RECT 45.900 20.850 47.400 24.900 ;
        RECT 42.300 14.850 46.500 16.050 ;
        RECT 42.300 10.200 43.500 14.850 ;
        RECT 44.700 14.250 46.500 14.850 ;
        RECT 47.850 10.200 48.900 20.550 ;
        RECT 3.600 9.000 7.050 10.200 ;
        RECT 9.600 9.000 13.500 10.200 ;
        RECT 15.600 9.000 19.500 10.200 ;
        RECT 21.600 9.000 25.800 10.200 ;
        RECT 27.600 9.000 30.900 10.200 ;
        RECT 33.600 9.000 37.500 10.200 ;
        RECT 39.600 9.000 43.500 10.200 ;
        RECT 45.600 9.000 48.900 10.200 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 9.000 ;
        RECT 6.600 1.500 8.400 8.100 ;
        RECT 9.600 2.100 11.400 9.000 ;
        RECT 12.600 1.500 14.400 8.100 ;
        RECT 15.600 2.100 17.400 9.000 ;
        RECT 18.600 1.500 20.400 8.100 ;
        RECT 21.600 2.100 23.400 9.000 ;
        RECT 24.600 1.500 26.400 8.100 ;
        RECT 27.600 2.100 29.400 9.000 ;
        RECT 30.600 1.500 32.400 8.100 ;
        RECT 33.600 2.100 35.400 9.000 ;
        RECT 36.600 1.500 38.400 8.100 ;
        RECT 39.600 2.100 41.400 9.000 ;
        RECT 42.600 1.500 44.400 8.100 ;
        RECT 45.600 2.100 47.400 9.000 ;
        RECT 48.600 1.500 50.400 8.100 ;
  END
END CLKBUF3
MACRO DFFNEGX1
  CLASS CORE ;
  FOREIGN DFFNEGX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 33.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.450 18.450 32.550 20.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 33.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 33.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.300 24.300 2.100 36.900 ;
        RECT 3.300 25.350 5.100 37.500 ;
        RECT 8.100 32.100 9.900 36.900 ;
        RECT 6.000 30.900 9.900 32.100 ;
        RECT 12.900 30.900 14.700 37.500 ;
        RECT 15.900 30.900 17.700 36.900 ;
        RECT 18.900 30.900 20.700 37.500 ;
        RECT 23.400 30.900 25.200 36.900 ;
        RECT 6.000 28.800 8.100 30.900 ;
        RECT 15.900 30.000 16.800 30.900 ;
        RECT 9.000 27.300 10.800 30.000 ;
        RECT 12.000 29.100 18.600 30.000 ;
        RECT 12.000 28.200 13.800 29.100 ;
        RECT 16.800 28.200 18.600 29.100 ;
        RECT 23.100 28.800 25.200 30.900 ;
        RECT 9.000 25.200 11.100 27.300 ;
        RECT 24.000 27.000 25.800 27.600 ;
        RECT 18.900 25.800 25.800 27.000 ;
        RECT 18.900 25.200 20.700 25.800 ;
        RECT 18.900 24.300 19.800 25.200 ;
        RECT 27.900 24.900 29.700 37.500 ;
        RECT 30.900 24.900 32.700 36.900 ;
        RECT 0.300 23.400 19.800 24.300 ;
        RECT 0.300 8.100 1.200 23.400 ;
        RECT 7.200 23.100 19.800 23.400 ;
        RECT 7.200 22.500 9.000 23.100 ;
        RECT 30.900 22.800 32.100 24.900 ;
        RECT 26.400 21.000 32.100 22.800 ;
        RECT 30.450 20.850 32.100 21.000 ;
        RECT 2.700 18.450 3.150 20.550 ;
        RECT 6.450 19.200 8.250 19.650 ;
        RECT 6.450 18.450 12.150 19.200 ;
        RECT 2.700 18.150 3.450 18.450 ;
        RECT 6.450 18.150 12.450 18.450 ;
        RECT 2.700 12.000 3.900 18.150 ;
        RECT 6.450 17.850 14.550 18.150 ;
        RECT 5.850 15.000 7.950 15.900 ;
        RECT 5.850 14.100 15.600 15.000 ;
        RECT 5.850 13.800 7.950 14.100 ;
        RECT 13.800 13.200 15.600 14.100 ;
        RECT 23.100 14.400 25.200 14.700 ;
        RECT 2.100 11.400 3.900 12.000 ;
        RECT 8.700 11.400 10.800 13.200 ;
        RECT 23.100 12.600 29.400 14.400 ;
        RECT 2.100 10.200 22.500 11.400 ;
        RECT 7.200 8.400 9.000 10.200 ;
        RECT 20.700 9.600 22.500 10.200 ;
        RECT 26.400 10.650 28.200 11.250 ;
        RECT 30.900 10.650 32.100 18.150 ;
        RECT 26.400 9.450 32.100 10.650 ;
        RECT 30.900 8.100 32.100 9.450 ;
        RECT 0.300 2.100 2.100 8.100 ;
        RECT 3.300 1.500 5.100 8.100 ;
        RECT 6.300 5.100 8.400 7.200 ;
        RECT 12.000 6.900 13.800 7.800 ;
        RECT 12.000 6.000 16.800 6.900 ;
        RECT 15.900 5.100 16.800 6.000 ;
        RECT 6.300 4.050 9.900 5.100 ;
        RECT 8.100 2.100 9.900 4.050 ;
        RECT 12.600 1.500 14.400 5.100 ;
        RECT 15.900 2.100 17.700 5.100 ;
        RECT 18.900 1.500 20.700 5.100 ;
        RECT 23.100 4.200 25.200 7.200 ;
        RECT 23.400 2.100 25.200 4.200 ;
        RECT 27.900 1.500 29.700 8.100 ;
        RECT 30.900 2.100 32.700 8.100 ;
      LAYER via1 ;
        RECT 8.700 11.100 10.800 13.200 ;
        RECT 23.100 5.100 25.200 7.200 ;
      LAYER metal2 ;
        RECT 6.000 28.800 8.100 30.900 ;
        RECT 23.100 28.800 25.200 30.900 ;
        RECT 6.450 15.900 7.500 28.800 ;
        RECT 9.000 25.200 11.100 27.300 ;
        RECT 23.100 27.000 24.300 28.800 ;
        RECT 23.100 25.800 24.000 27.000 ;
        RECT 5.850 13.800 7.950 15.900 ;
        RECT 6.450 7.200 7.500 13.800 ;
        RECT 9.450 13.200 10.800 25.200 ;
        RECT 8.700 11.100 10.800 13.200 ;
        RECT 23.100 14.700 24.300 25.800 ;
        RECT 23.100 12.600 25.200 14.700 ;
        RECT 23.100 7.200 24.300 12.600 ;
        RECT 6.300 5.100 8.400 7.200 ;
        RECT 23.100 5.100 25.200 7.200 ;
  END
END DFFNEGX1
MACRO DFFPOSX1
  CLASS CORE ;
  FOREIGN DFFPOSX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 36.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 18.450 17.550 20.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.450 18.450 32.550 20.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 36.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 36.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.650 26.700 3.450 36.900 ;
        RECT 1.050 24.900 3.450 26.700 ;
        RECT 4.650 24.900 6.450 37.500 ;
        RECT 10.050 31.800 11.850 36.900 ;
        RECT 7.950 30.900 11.850 31.800 ;
        RECT 14.850 30.900 16.650 37.500 ;
        RECT 17.850 30.900 19.650 36.900 ;
        RECT 20.850 30.900 22.650 37.500 ;
        RECT 25.350 30.900 27.150 36.900 ;
        RECT 7.950 28.800 10.050 30.900 ;
        RECT 17.850 30.000 18.750 30.900 ;
        RECT 13.950 29.100 20.550 30.000 ;
        RECT 13.950 28.200 15.750 29.100 ;
        RECT 18.750 28.200 20.550 29.100 ;
        RECT 25.050 28.800 27.150 30.900 ;
        RECT 7.950 27.000 10.050 27.900 ;
        RECT 22.350 27.300 24.150 27.900 ;
        RECT 7.950 25.800 17.550 27.000 ;
        RECT 15.750 25.200 17.550 25.800 ;
        RECT 18.450 26.400 24.150 27.300 ;
        RECT 1.050 24.000 1.950 24.900 ;
        RECT 18.450 24.300 19.350 26.400 ;
        RECT 22.350 26.100 24.150 26.400 ;
        RECT 25.050 26.100 28.050 27.900 ;
        RECT 25.050 25.200 26.250 26.100 ;
        RECT 10.950 24.000 19.350 24.300 ;
        RECT 1.050 23.400 19.350 24.000 ;
        RECT 21.450 24.300 26.250 25.200 ;
        RECT 30.150 24.900 31.950 37.500 ;
        RECT 1.050 22.800 12.750 23.400 ;
        RECT 1.050 8.100 1.950 22.800 ;
        RECT 10.950 22.500 12.750 22.800 ;
        RECT 7.350 18.450 15.150 19.500 ;
        RECT 3.450 15.750 5.250 18.150 ;
        RECT 7.350 17.700 9.150 18.450 ;
        RECT 4.050 12.900 5.250 15.750 ;
        RECT 9.600 12.900 11.400 13.500 ;
        RECT 4.050 11.700 11.400 12.900 ;
        RECT 21.450 11.700 22.350 24.300 ;
        RECT 33.150 20.550 34.950 36.900 ;
        RECT 28.200 18.450 30.150 20.250 ;
        RECT 32.850 18.450 34.950 20.550 ;
        RECT 25.050 13.500 27.150 14.400 ;
        RECT 30.450 13.500 32.250 14.250 ;
        RECT 25.050 12.450 32.250 13.500 ;
        RECT 25.050 12.300 27.150 12.450 ;
        RECT 10.350 10.500 22.350 11.700 ;
        RECT 10.350 8.700 11.400 10.500 ;
        RECT 20.550 9.900 22.350 10.500 ;
        RECT 27.750 11.100 29.550 11.550 ;
        RECT 33.150 11.100 34.950 18.450 ;
        RECT 27.750 9.750 34.950 11.100 ;
        RECT 1.050 6.300 3.450 8.100 ;
        RECT 1.650 2.100 3.450 6.300 ;
        RECT 4.650 1.500 6.450 8.100 ;
        RECT 7.350 5.700 9.450 7.200 ;
        RECT 10.350 6.900 12.150 8.700 ;
        RECT 13.350 6.900 15.150 7.800 ;
        RECT 13.350 6.000 18.150 6.900 ;
        RECT 7.350 5.100 11.250 5.700 ;
        RECT 17.250 5.100 18.150 6.000 ;
        RECT 24.750 5.100 27.150 7.200 ;
        RECT 7.650 4.200 11.250 5.100 ;
        RECT 9.450 2.100 11.250 4.200 ;
        RECT 13.950 1.500 15.750 5.100 ;
        RECT 17.250 2.100 19.050 5.100 ;
        RECT 20.250 2.100 22.050 5.100 ;
        RECT 24.750 2.100 26.550 5.100 ;
        RECT 20.250 1.500 21.450 2.100 ;
        RECT 29.850 1.500 31.650 8.100 ;
        RECT 33.150 2.100 34.950 9.750 ;
      LAYER via1 ;
        RECT 25.050 5.100 27.150 7.200 ;
      LAYER metal2 ;
        RECT 7.950 25.800 10.050 30.900 ;
        RECT 25.050 28.800 27.150 30.900 ;
        RECT 8.250 22.950 9.450 25.800 ;
        RECT 7.650 21.750 9.450 22.950 ;
        RECT 7.650 7.200 8.850 21.750 ;
        RECT 25.050 14.400 26.250 28.800 ;
        RECT 25.050 12.300 27.150 14.400 ;
        RECT 25.050 7.200 26.250 12.300 ;
        RECT 7.350 5.100 9.450 7.200 ;
        RECT 25.050 5.100 27.150 7.200 ;
  END
END DFFPOSX1
MACRO DFFSR
  CLASS CORE ;
  FOREIGN DFFSR ;
  ORIGIN 0.000 0.000 ;
  SIZE 69.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 27.450 12.450 29.550 14.550 ;
    END
  END D
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END S
  PIN R
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END R
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 33.450 12.450 35.550 14.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 63.450 18.450 65.550 20.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 69.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 69.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 30.900 3.000 37.500 ;
        RECT 4.200 31.800 6.000 36.900 ;
        RECT 3.900 30.900 6.000 31.800 ;
        RECT 7.200 30.900 9.000 37.500 ;
        RECT 3.900 30.000 4.800 30.900 ;
        RECT 1.200 29.100 4.800 30.000 ;
        RECT 1.200 13.050 2.400 29.100 ;
        RECT 5.700 27.900 7.500 28.200 ;
        RECT 10.200 27.900 12.000 36.900 ;
        RECT 13.200 30.900 15.000 37.500 ;
        RECT 16.800 34.050 18.600 36.900 ;
        RECT 16.800 31.950 18.900 34.050 ;
        RECT 19.800 33.900 21.600 36.900 ;
        RECT 19.800 31.800 21.900 33.900 ;
        RECT 22.800 30.900 24.600 36.900 ;
        RECT 25.800 30.900 27.600 37.500 ;
        RECT 22.200 28.800 24.300 30.900 ;
        RECT 29.850 29.550 31.650 36.900 ;
        RECT 32.850 30.900 34.650 37.500 ;
        RECT 35.850 30.900 37.650 36.900 ;
        RECT 38.850 33.900 40.650 36.900 ;
        RECT 41.850 33.900 43.650 36.900 ;
        RECT 44.850 33.900 46.650 36.900 ;
        RECT 38.850 31.800 40.950 33.900 ;
        RECT 41.850 31.800 43.950 33.900 ;
        RECT 44.850 31.800 46.950 33.900 ;
        RECT 47.850 30.900 49.650 37.500 ;
        RECT 53.850 36.900 55.500 37.500 ;
        RECT 50.850 30.900 52.650 36.900 ;
        RECT 53.850 30.900 55.650 36.900 ;
        RECT 56.850 30.900 58.650 36.900 ;
        RECT 59.850 30.900 61.650 37.500 ;
        RECT 5.700 26.850 24.900 27.900 ;
        RECT 29.850 27.450 32.550 29.550 ;
        RECT 35.850 28.800 38.850 30.900 ;
        RECT 41.850 30.000 43.950 30.900 ;
        RECT 41.850 28.800 49.950 30.000 ;
        RECT 35.850 27.000 38.550 28.800 ;
        RECT 48.150 28.200 49.950 28.800 ;
        RECT 50.850 28.050 51.900 30.900 ;
        RECT 57.450 30.000 58.650 30.900 ;
        RECT 57.450 29.100 61.350 30.000 ;
        RECT 63.000 29.100 64.800 36.900 ;
        RECT 66.000 30.900 67.800 37.500 ;
        RECT 54.750 28.050 56.550 28.800 ;
        RECT 5.700 26.400 7.500 26.850 ;
        RECT 23.850 26.100 24.900 26.850 ;
        RECT 39.450 26.100 41.550 27.150 ;
        RECT 9.000 25.200 10.800 25.800 ;
        RECT 18.900 25.200 21.000 25.800 ;
        RECT 9.000 24.000 21.000 25.200 ;
        RECT 23.850 25.050 41.550 26.100 ;
        RECT 44.850 26.100 46.950 27.150 ;
        RECT 50.850 27.000 56.550 28.050 ;
        RECT 60.450 26.100 61.350 29.100 ;
        RECT 44.850 25.050 61.350 26.100 ;
        RECT 18.900 23.700 21.000 24.000 ;
        RECT 23.850 23.100 59.550 24.150 ;
        RECT 23.850 22.350 24.900 23.100 ;
        RECT 57.750 22.350 59.550 23.100 ;
        RECT 13.950 21.300 24.900 22.350 ;
        RECT 35.550 22.050 37.650 22.200 ;
        RECT 3.600 15.450 5.400 18.150 ;
        RECT 10.200 17.700 11.550 18.150 ;
        RECT 13.950 17.700 15.000 21.300 ;
        RECT 21.900 19.350 23.700 19.950 ;
        RECT 30.450 19.350 32.550 20.850 ;
        RECT 33.750 20.250 37.650 22.050 ;
        RECT 35.550 20.100 37.650 20.250 ;
        RECT 21.900 19.200 32.550 19.350 ;
        RECT 42.750 19.200 44.550 21.600 ;
        RECT 21.900 18.150 44.550 19.200 ;
        RECT 47.250 20.250 52.650 22.050 ;
        RECT 10.200 16.650 15.000 17.700 ;
        RECT 47.250 17.250 48.150 20.250 ;
        RECT 10.200 15.900 12.600 16.650 ;
        RECT 16.950 16.200 48.150 17.250 ;
        RECT 4.350 15.000 5.400 15.450 ;
        RECT 16.950 15.000 18.000 16.200 ;
        RECT 4.350 13.950 18.000 15.000 ;
        RECT 18.900 13.050 20.700 14.850 ;
        RECT 1.200 11.700 18.000 13.050 ;
        RECT 1.200 8.100 2.400 11.700 ;
        RECT 15.900 10.950 18.000 11.700 ;
        RECT 5.400 10.200 7.200 10.800 ;
        RECT 5.400 9.000 13.800 10.200 ;
        RECT 12.300 8.100 13.800 9.000 ;
        RECT 18.900 9.900 19.800 13.050 ;
        RECT 27.450 11.100 29.100 12.150 ;
        RECT 18.900 8.850 26.100 9.900 ;
        RECT 27.300 9.300 29.100 11.100 ;
        RECT 33.750 9.300 35.550 12.150 ;
        RECT 51.750 11.400 59.550 13.200 ;
        RECT 21.300 8.100 23.100 8.850 ;
        RECT 25.200 8.100 26.100 8.850 ;
        RECT 40.950 8.100 47.550 9.900 ;
        RECT 51.750 8.100 53.250 11.400 ;
        RECT 60.450 8.100 61.350 25.050 ;
        RECT 63.450 20.850 64.800 29.100 ;
        RECT 1.200 2.100 3.000 8.100 ;
        RECT 6.600 1.500 8.400 8.100 ;
        RECT 12.000 2.100 13.800 8.100 ;
        RECT 16.200 5.100 18.300 7.200 ;
        RECT 19.200 5.100 21.300 7.200 ;
        RECT 22.200 5.100 24.300 7.200 ;
        RECT 25.200 7.050 27.900 8.100 ;
        RECT 26.100 6.150 27.900 7.050 ;
        RECT 29.850 6.000 32.550 8.100 ;
        RECT 16.200 2.100 18.000 5.100 ;
        RECT 19.200 2.100 21.000 5.100 ;
        RECT 22.200 2.100 24.000 5.100 ;
        RECT 25.200 1.500 27.000 5.100 ;
        RECT 29.850 2.100 31.650 6.000 ;
        RECT 35.850 5.100 37.950 7.200 ;
        RECT 38.850 5.100 40.950 7.200 ;
        RECT 41.850 5.100 43.950 7.200 ;
        RECT 44.850 5.100 46.950 7.200 ;
        RECT 48.900 6.900 53.250 8.100 ;
        RECT 32.850 1.500 34.650 5.100 ;
        RECT 35.850 2.100 37.650 5.100 ;
        RECT 38.850 2.100 40.650 5.100 ;
        RECT 41.850 2.100 43.650 5.100 ;
        RECT 44.850 2.100 46.650 5.100 ;
        RECT 48.900 2.100 50.700 6.900 ;
        RECT 54.150 1.500 55.950 8.100 ;
        RECT 59.550 2.100 61.350 8.100 ;
        RECT 63.450 5.100 64.800 18.150 ;
        RECT 63.000 2.100 64.800 5.100 ;
        RECT 66.000 1.500 67.800 5.100 ;
      LAYER via1 ;
        RECT 30.450 27.450 32.550 29.550 ;
        RECT 36.750 28.800 38.850 30.900 ;
        RECT 39.450 25.050 41.550 27.150 ;
        RECT 30.450 18.750 32.550 20.850 ;
        RECT 30.450 6.000 32.550 8.100 ;
      LAYER metal2 ;
        RECT 15.900 31.950 18.900 34.050 ;
        RECT 15.900 13.050 17.400 31.950 ;
        RECT 19.800 31.800 21.900 33.900 ;
        RECT 38.850 31.800 40.950 33.900 ;
        RECT 19.800 25.800 21.000 31.800 ;
        RECT 18.900 23.700 21.000 25.800 ;
        RECT 15.900 10.950 18.000 13.050 ;
        RECT 16.200 7.200 17.550 10.950 ;
        RECT 19.800 7.200 21.000 23.700 ;
        RECT 22.200 28.800 24.300 30.900 ;
        RECT 22.200 7.200 23.400 28.800 ;
        RECT 30.450 27.450 32.550 29.550 ;
        RECT 36.750 28.800 38.850 30.900 ;
        RECT 30.900 20.850 31.950 27.450 ;
        RECT 36.750 22.200 37.950 28.800 ;
        RECT 39.750 27.150 40.950 31.800 ;
        RECT 41.850 28.800 43.950 33.900 ;
        RECT 39.450 25.050 41.550 27.150 ;
        RECT 30.450 18.750 32.550 20.850 ;
        RECT 35.550 20.100 37.950 22.200 ;
        RECT 30.900 8.100 31.950 18.750 ;
        RECT 16.200 5.100 18.300 7.200 ;
        RECT 19.200 5.100 21.300 7.200 ;
        RECT 22.200 5.100 24.300 7.200 ;
        RECT 30.450 6.000 32.550 8.100 ;
        RECT 36.750 7.200 37.950 20.100 ;
        RECT 39.750 7.200 40.950 25.050 ;
        RECT 42.750 7.200 43.950 28.800 ;
        RECT 35.850 5.100 37.950 7.200 ;
        RECT 38.850 5.100 40.950 7.200 ;
        RECT 41.850 5.100 43.950 7.200 ;
        RECT 44.850 31.800 46.950 33.900 ;
        RECT 44.850 27.150 46.200 31.800 ;
        RECT 44.850 25.050 46.950 27.150 ;
        RECT 44.850 7.200 46.200 25.050 ;
        RECT 44.850 5.100 46.950 7.200 ;
  END
END DFFSR
MACRO FAX1
  CLASS CORE ;
  FOREIGN FAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 45.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 30.450 15.450 32.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END C
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 36.450 15.450 38.550 17.550 ;
    END
  END YS
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 42.450 15.450 44.550 17.550 ;
    END
  END YC
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 45.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 45.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 25.800 3.000 36.900 ;
        RECT 4.200 26.700 6.000 37.500 ;
        RECT 7.200 25.800 9.000 36.900 ;
        RECT 1.200 24.900 9.000 25.800 ;
        RECT 10.200 26.100 12.000 36.900 ;
        RECT 10.200 24.750 12.900 26.100 ;
        RECT 14.700 24.900 16.500 37.500 ;
        RECT 17.700 27.000 19.500 36.900 ;
        RECT 20.700 27.900 22.500 37.500 ;
        RECT 23.700 27.000 25.500 36.900 ;
        RECT 17.700 26.400 25.500 27.000 ;
        RECT 17.700 26.100 24.900 26.400 ;
        RECT 17.700 24.900 19.500 26.100 ;
        RECT 10.800 24.000 12.900 24.750 ;
        RECT 21.900 24.000 24.000 24.300 ;
        RECT 26.700 24.000 28.650 36.900 ;
        RECT 21.900 22.200 25.800 24.000 ;
        RECT 26.700 22.800 28.800 24.000 ;
        RECT 26.700 21.900 32.100 22.800 ;
        RECT 33.000 22.500 34.800 37.500 ;
        RECT 36.000 32.250 37.800 36.900 ;
        RECT 35.700 30.900 37.800 32.250 ;
        RECT 39.000 30.900 40.800 37.500 ;
        RECT 42.000 32.850 43.800 36.900 ;
        RECT 42.000 30.900 44.100 32.850 ;
        RECT 35.700 23.400 36.600 30.900 ;
        RECT 37.500 26.400 39.600 26.550 ;
        RECT 37.500 24.600 41.400 26.400 ;
        RECT 37.500 24.450 39.600 24.600 ;
        RECT 35.700 22.500 38.100 23.400 ;
        RECT 31.200 21.150 32.100 21.900 ;
        RECT 31.200 20.250 35.700 21.150 ;
        RECT 33.900 19.350 35.700 20.250 ;
        RECT 3.450 17.550 5.100 18.150 ;
        RECT 20.100 17.550 21.900 18.150 ;
        RECT 26.550 17.550 28.350 18.150 ;
        RECT 36.900 17.850 38.100 22.500 ;
        RECT 42.900 17.850 44.100 30.900 ;
        RECT 3.300 15.750 5.100 17.550 ;
        RECT 8.850 16.350 28.350 17.550 ;
        RECT 8.850 15.750 11.100 16.350 ;
        RECT 26.550 16.200 28.350 16.350 ;
        RECT 3.450 10.800 5.100 15.750 ;
        RECT 30.450 14.400 32.100 15.150 ;
        RECT 28.500 13.500 32.100 14.400 ;
        RECT 6.300 12.600 32.100 13.500 ;
        RECT 6.300 12.450 13.500 12.600 ;
        RECT 6.300 11.700 8.100 12.450 ;
        RECT 11.700 11.700 13.500 12.450 ;
        RECT 17.700 11.700 19.500 12.600 ;
        RECT 14.700 10.800 16.500 11.400 ;
        RECT 32.400 10.800 34.200 11.550 ;
        RECT 3.450 9.900 34.200 10.800 ;
        RECT 14.700 9.600 16.500 9.900 ;
        RECT 32.400 9.600 34.200 9.900 ;
        RECT 1.200 7.200 9.000 8.100 ;
        RECT 1.200 2.100 3.000 7.200 ;
        RECT 4.200 1.500 6.000 6.300 ;
        RECT 7.200 2.100 9.000 7.200 ;
        RECT 10.200 6.900 12.300 9.000 ;
        RECT 10.200 2.100 12.000 6.900 ;
        RECT 14.700 1.500 16.500 7.500 ;
        RECT 17.700 6.900 25.500 7.800 ;
        RECT 17.700 2.100 19.500 6.900 ;
        RECT 20.700 1.500 22.500 6.000 ;
        RECT 23.700 2.100 25.500 6.900 ;
        RECT 26.700 6.600 28.800 8.700 ;
        RECT 26.700 2.100 28.650 6.600 ;
        RECT 33.000 2.100 34.800 7.800 ;
        RECT 36.900 7.200 38.100 15.150 ;
        RECT 36.300 6.000 38.100 7.200 ;
        RECT 36.300 5.100 37.200 6.000 ;
        RECT 42.900 5.100 44.100 15.150 ;
        RECT 36.000 2.100 37.800 5.100 ;
        RECT 33.000 1.500 34.200 2.100 ;
        RECT 39.000 1.500 40.800 5.100 ;
        RECT 42.000 2.100 44.100 5.100 ;
      LAYER metal2 ;
        RECT 10.800 25.800 12.900 26.100 ;
        RECT 37.500 25.800 39.600 26.550 ;
        RECT 10.800 24.900 39.600 25.800 ;
        RECT 10.800 24.000 12.900 24.900 ;
        RECT 11.250 9.000 12.150 24.000 ;
        RECT 21.900 22.200 24.000 24.900 ;
        RECT 37.500 24.450 39.600 24.900 ;
        RECT 26.700 21.900 28.800 24.000 ;
        RECT 10.200 6.900 12.300 9.000 ;
        RECT 27.300 8.700 28.200 21.900 ;
        RECT 26.700 6.600 28.800 8.700 ;
  END
END FAX1
MACRO FILL
  CLASS CORE ;
  FOREIGN FILL ;
  ORIGIN 0.000 0.000 ;
  SIZE 3.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 3.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 3.900 1.200 ;
    END
  END gnd
END FILL
MACRO HAX1
  CLASS CORE ;
  FOREIGN HAX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 30.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.450 17.550 17.550 ;
    END
  END B
  PIN YS
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 24.450 18.450 26.550 20.550 ;
    END
  END YS
  PIN YC
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END YC
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 30.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 30.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.350 30.900 3.150 36.900 ;
        RECT 4.350 31.500 6.150 37.500 ;
        RECT 1.650 30.600 3.150 30.900 ;
        RECT 7.350 30.900 9.150 36.900 ;
        RECT 10.350 30.900 12.150 36.900 ;
        RECT 13.350 30.900 15.150 37.500 ;
        RECT 7.350 30.600 8.550 30.900 ;
        RECT 1.650 29.700 8.550 30.600 ;
        RECT 7.050 20.550 7.950 29.700 ;
        RECT 10.350 20.550 11.550 30.900 ;
        RECT 16.350 24.900 18.150 36.900 ;
        RECT 20.850 24.900 22.650 37.500 ;
        RECT 23.850 30.900 25.650 37.500 ;
        RECT 26.850 30.900 28.650 36.900 ;
        RECT 27.150 30.000 28.050 30.900 ;
        RECT 24.900 29.100 28.050 30.000 ;
        RECT 16.650 24.000 17.550 24.900 ;
        RECT 16.650 23.100 24.000 24.000 ;
        RECT 22.200 22.200 24.000 23.100 ;
        RECT 6.450 18.450 8.550 20.550 ;
        RECT 9.750 18.450 12.150 20.550 ;
        RECT 16.950 18.300 18.750 20.100 ;
        RECT 3.450 17.550 5.100 18.150 ;
        RECT 16.950 17.850 18.150 18.300 ;
        RECT 17.550 17.550 18.150 17.850 ;
        RECT 3.450 15.750 5.250 17.550 ;
        RECT 6.450 16.800 8.250 17.100 ;
        RECT 6.450 15.750 15.150 16.800 ;
        RECT 4.050 12.300 4.950 15.750 ;
        RECT 6.450 15.300 8.250 15.750 ;
        RECT 17.850 15.450 18.150 17.550 ;
        RECT 19.350 12.300 21.150 13.200 ;
        RECT 4.050 11.400 21.150 12.300 ;
        RECT 22.650 10.650 23.550 22.200 ;
        RECT 24.900 20.850 26.100 29.100 ;
        RECT 5.850 9.900 7.950 10.200 ;
        RECT 5.850 8.100 11.550 9.900 ;
        RECT 22.200 9.750 24.000 10.650 ;
        RECT 17.850 8.850 24.000 9.750 ;
        RECT 1.350 1.500 3.150 8.100 ;
        RECT 5.850 2.100 7.650 8.100 ;
        RECT 8.850 4.950 10.950 7.200 ;
        RECT 8.850 2.100 10.650 4.950 ;
        RECT 11.850 1.500 13.650 7.200 ;
        RECT 14.850 3.000 16.650 8.100 ;
        RECT 17.850 3.900 19.650 8.850 ;
        RECT 20.850 3.000 22.650 7.500 ;
        RECT 24.900 7.200 26.100 18.150 ;
        RECT 24.900 6.300 28.050 7.200 ;
        RECT 27.150 5.100 28.050 6.300 ;
        RECT 14.850 2.100 22.650 3.000 ;
        RECT 23.850 1.500 25.650 5.100 ;
        RECT 26.850 2.100 28.650 5.100 ;
      LAYER via1 ;
        RECT 8.850 5.100 10.950 7.200 ;
      LAYER metal2 ;
        RECT 6.450 18.450 8.550 20.550 ;
        RECT 9.750 18.450 11.850 20.550 ;
        RECT 7.050 10.200 7.950 18.450 ;
        RECT 5.850 8.100 7.950 10.200 ;
        RECT 9.750 7.200 10.950 18.450 ;
        RECT 8.850 5.100 10.950 7.200 ;
  END
END HAX1
MACRO INVX1
  CLASS CORE ;
  FOREIGN INVX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 6.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 6.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 30.900 2.400 37.500 ;
        RECT 3.600 30.900 5.400 36.900 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 17.850 5.100 30.900 ;
        RECT 3.900 5.100 5.100 15.150 ;
        RECT 0.600 1.500 2.400 5.100 ;
        RECT 3.600 2.100 5.400 5.100 ;
  END
END INVX1
MACRO INVX2
  CLASS CORE ;
  FOREIGN INVX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 6.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 6.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 6.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.900 5.400 36.900 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 17.850 5.100 24.900 ;
        RECT 3.900 8.100 5.100 15.150 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 8.100 ;
  END
END INVX2
MACRO INVX4
  CLASS CORE ;
  FOREIGN INVX4 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 9.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.900 5.400 36.900 ;
        RECT 6.600 24.900 8.400 37.500 ;
        RECT 3.900 22.650 5.100 24.900 ;
        RECT 3.900 21.450 8.100 22.650 ;
        RECT 6.900 20.850 8.100 21.450 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 6.900 10.950 8.100 18.150 ;
        RECT 3.900 9.750 8.100 10.950 ;
        RECT 3.900 8.100 5.100 9.750 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 8.100 ;
        RECT 6.600 1.500 8.400 8.100 ;
  END
END INVX4
MACRO INVX8
  CLASS CORE ;
  FOREIGN INVX8 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END A
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.000 5.400 36.900 ;
        RECT 6.600 24.900 8.400 37.500 ;
        RECT 9.600 24.900 11.400 36.900 ;
        RECT 12.600 24.900 14.400 37.500 ;
        RECT 9.600 24.000 11.100 24.900 ;
        RECT 3.600 23.100 11.100 24.000 ;
        RECT 9.900 20.850 11.100 23.100 ;
        RECT 3.600 15.750 5.400 18.150 ;
        RECT 9.900 10.200 11.100 18.150 ;
        RECT 3.600 9.000 11.100 10.200 ;
        RECT 3.600 8.100 4.800 9.000 ;
        RECT 9.600 8.100 11.100 9.000 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 8.100 ;
        RECT 6.600 1.500 8.400 8.100 ;
        RECT 9.600 2.100 11.400 8.100 ;
        RECT 12.600 1.500 14.400 8.100 ;
  END
END INVX8
MACRO LATCH
  CLASS CORE ;
  FOREIGN LATCH ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END D
  PIN CLK
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END CLK
  PIN Q
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.450 18.450 20.550 20.550 ;
    END
  END Q
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 21.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 21.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 24.900 3.000 36.900 ;
        RECT 4.200 24.900 6.000 37.500 ;
        RECT 9.300 30.900 11.250 36.900 ;
        RECT 9.600 28.800 11.700 30.900 ;
        RECT 1.200 24.000 2.400 24.900 ;
        RECT 9.600 24.000 11.700 25.200 ;
        RECT 15.000 24.900 16.800 37.500 ;
        RECT 18.000 25.950 19.800 36.900 ;
        RECT 18.000 24.900 20.100 25.950 ;
        RECT 1.200 23.100 8.700 24.000 ;
        RECT 9.600 23.100 17.400 24.000 ;
        RECT 1.200 21.300 2.550 23.100 ;
        RECT 0.450 19.200 2.550 21.300 ;
        RECT 7.500 22.200 8.700 23.100 ;
        RECT 15.600 22.200 17.400 23.100 ;
        RECT 7.500 20.400 9.900 22.200 ;
        RECT 18.900 20.850 20.100 24.900 ;
        RECT 6.750 18.450 12.150 19.050 ;
        RECT 6.750 18.150 12.450 18.450 ;
        RECT 3.450 17.550 5.100 18.150 ;
        RECT 3.150 15.750 5.100 17.550 ;
        RECT 1.050 8.100 3.150 10.200 ;
        RECT 4.050 9.900 5.100 15.750 ;
        RECT 6.750 14.400 7.800 18.150 ;
        RECT 18.900 14.850 20.100 18.150 ;
        RECT 6.000 12.600 7.800 14.400 ;
        RECT 10.800 13.050 12.600 14.850 ;
        RECT 14.100 13.050 20.100 14.850 ;
        RECT 10.800 9.900 11.700 13.050 ;
        RECT 4.050 9.000 11.700 9.900 ;
        RECT 8.550 8.100 11.700 9.000 ;
        RECT 18.900 8.100 20.100 13.050 ;
        RECT 1.200 2.100 3.000 8.100 ;
        RECT 4.200 1.500 6.000 8.100 ;
        RECT 9.600 5.100 11.700 7.200 ;
        RECT 9.300 2.100 11.400 5.100 ;
        RECT 15.000 1.500 16.800 8.100 ;
        RECT 18.000 6.750 20.100 8.100 ;
        RECT 18.000 2.100 19.800 6.750 ;
      LAYER metal2 ;
        RECT 9.600 28.800 11.700 30.900 ;
        RECT 9.600 25.200 10.800 28.800 ;
        RECT 9.600 23.100 11.700 25.200 ;
        RECT 0.450 19.200 2.550 21.300 ;
        RECT 1.200 10.200 2.400 19.200 ;
        RECT 1.050 8.100 3.150 10.200 ;
        RECT 9.600 7.200 10.800 23.100 ;
        RECT 9.600 5.100 11.700 7.200 ;
  END
END LATCH
MACRO MUX2X1
  CLASS CORE ;
  FOREIGN MUX2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 15.450 14.550 17.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN S
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END S
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 15.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 15.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 29.850 2.400 35.700 ;
        RECT 0.600 29.700 1.800 29.850 ;
        RECT 0.600 24.600 1.500 29.700 ;
        RECT 3.600 25.500 5.400 37.500 ;
        RECT 8.100 26.400 9.900 36.900 ;
        RECT 8.100 25.500 11.100 26.400 ;
        RECT 0.600 23.700 8.400 24.600 ;
        RECT 0.600 15.750 2.400 18.150 ;
        RECT 7.200 16.500 8.400 23.700 ;
        RECT 9.900 20.850 11.100 25.500 ;
        RECT 12.600 24.900 14.400 37.500 ;
        RECT 3.600 12.750 5.400 15.150 ;
        RECT 6.600 14.700 8.400 16.500 ;
        RECT 7.050 10.500 8.400 14.700 ;
        RECT 0.600 9.600 8.400 10.500 ;
        RECT 0.600 6.300 1.500 9.600 ;
        RECT 9.900 8.700 11.100 18.150 ;
        RECT 12.600 13.050 14.400 15.150 ;
        RECT 0.600 3.300 2.400 6.300 ;
        RECT 3.600 3.900 5.400 8.700 ;
        RECT 8.100 7.050 11.100 8.700 ;
        RECT 3.600 1.500 4.800 3.900 ;
        RECT 8.100 3.300 9.900 7.050 ;
        RECT 12.600 3.300 14.400 9.300 ;
        RECT 12.600 1.500 13.800 3.300 ;
  END
END MUX2X1
MACRO NAND2X1
  CLASS CORE ;
  FOREIGN NAND2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 9.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 9.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 30.900 2.400 37.500 ;
        RECT 3.600 30.900 5.400 36.900 ;
        RECT 6.600 30.900 8.400 37.500 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 17.850 5.100 30.900 ;
        RECT 6.450 15.750 8.250 18.150 ;
        RECT 3.900 9.000 5.100 15.150 ;
        RECT 3.900 8.100 7.950 9.000 ;
        RECT 1.050 2.100 2.850 8.100 ;
        RECT 6.150 2.100 7.950 8.100 ;
        RECT 1.050 1.500 2.250 2.100 ;
  END
END NAND2X1
MACRO NAND3X1
  CLASS CORE ;
  FOREIGN NAND3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 37.800 12.900 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -0.900 -1.200 12.900 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 30.900 2.400 37.500 ;
        RECT 3.600 30.900 5.400 36.900 ;
        RECT 6.600 31.500 8.400 37.500 ;
        RECT 3.900 30.600 5.400 30.900 ;
        RECT 9.600 30.900 11.400 36.900 ;
        RECT 9.600 30.600 11.100 30.900 ;
        RECT 3.900 29.700 11.100 30.600 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 6.750 16.200 8.550 18.150 ;
        RECT 9.900 17.850 11.100 29.700 ;
        RECT 3.900 15.000 5.550 15.150 ;
        RECT 3.900 13.200 6.300 15.000 ;
        RECT 9.900 11.400 11.100 15.150 ;
        RECT 0.600 1.500 2.400 11.100 ;
        RECT 7.200 10.500 11.100 11.400 ;
        RECT 7.200 2.100 9.000 10.500 ;
  END
END NAND3X1
MACRO NOR2X1
  CLASS CORE ;
  FOREIGN NOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 9.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 10.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 10.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 5.700 26.100 7.500 36.900 ;
        RECT 3.900 24.900 7.500 26.100 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 17.850 5.100 24.900 ;
        RECT 6.450 15.750 8.250 18.150 ;
        RECT 3.900 5.100 5.100 15.150 ;
        RECT 0.600 1.500 2.400 5.100 ;
        RECT 3.600 2.100 5.400 5.100 ;
        RECT 6.600 1.500 8.400 5.100 ;
  END
END NOR2X1
MACRO NOR3X1
  CLASS CORE ;
  FOREIGN NOR3X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 24.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 18.450 5.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 15.450 8.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 15.450 17.550 17.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 25.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 25.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 27.000 2.400 36.900 ;
        RECT 3.600 27.900 5.400 37.500 ;
        RECT 6.600 36.000 14.400 36.900 ;
        RECT 6.600 27.000 8.400 36.000 ;
        RECT 0.600 26.100 8.400 27.000 ;
        RECT 9.600 27.300 11.400 35.100 ;
        RECT 12.600 28.200 14.400 36.000 ;
        RECT 15.600 36.000 23.400 36.900 ;
        RECT 15.600 27.300 17.400 36.000 ;
        RECT 9.600 26.400 17.400 27.300 ;
        RECT 18.600 27.300 20.400 35.100 ;
        RECT 18.600 22.500 19.800 27.300 ;
        RECT 21.600 26.700 23.400 36.000 ;
        RECT 15.900 21.450 19.800 22.500 ;
        RECT 3.750 15.750 5.550 18.150 ;
        RECT 12.450 15.750 14.250 18.150 ;
        RECT 15.900 17.850 17.100 21.450 ;
        RECT 6.900 14.850 8.550 15.150 ;
        RECT 6.900 13.050 9.300 14.850 ;
        RECT 15.900 7.050 17.100 15.150 ;
        RECT 7.200 6.000 17.100 7.050 ;
        RECT 7.200 5.100 8.100 6.000 ;
        RECT 14.400 5.100 15.300 6.000 ;
        RECT 3.450 1.500 5.400 5.100 ;
        RECT 6.600 2.100 8.400 5.100 ;
        RECT 9.600 1.500 11.400 5.100 ;
        RECT 12.600 2.100 15.300 5.100 ;
  END
END NOR3X1
MACRO OAI21X1
  CLASS CORE ;
  FOREIGN OAI21X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END C
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 13.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 13.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.050 24.900 2.850 37.500 ;
        RECT 6.150 26.100 7.950 36.900 ;
        RECT 9.150 30.900 10.950 37.500 ;
        RECT 6.150 24.900 8.100 26.100 ;
        RECT 6.900 20.850 8.100 24.900 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 4.050 14.550 5.550 15.150 ;
        RECT 4.050 12.750 5.850 14.550 ;
        RECT 6.900 10.350 8.100 18.150 ;
        RECT 9.450 12.750 11.250 15.150 ;
        RECT 6.900 9.450 10.800 10.350 ;
        RECT 0.600 7.650 8.400 8.550 ;
        RECT 0.600 2.100 2.400 7.650 ;
        RECT 3.600 1.500 5.400 6.750 ;
        RECT 6.600 2.100 8.400 7.650 ;
        RECT 9.600 8.100 10.800 9.450 ;
        RECT 9.600 2.100 11.400 8.100 ;
  END
END OAI21X1
MACRO OAI22X1
  CLASS CORE ;
  FOREIGN OAI22X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN C
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END C
  PIN D
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 15.450 11.550 17.550 ;
    END
  END D
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 16.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 16.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 5.100 24.900 8.400 36.900 ;
        RECT 11.100 24.900 12.900 37.500 ;
        RECT 6.900 20.850 8.100 24.900 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 14.550 5.550 15.150 ;
        RECT 3.900 12.750 5.700 14.550 ;
        RECT 6.900 11.700 8.100 18.150 ;
        RECT 12.450 15.750 14.250 18.150 ;
        RECT 9.450 14.550 10.800 15.150 ;
        RECT 9.000 12.750 10.800 14.550 ;
        RECT 6.900 10.650 10.800 11.700 ;
        RECT 0.600 7.650 8.400 8.550 ;
        RECT 9.900 8.100 10.800 10.650 ;
        RECT 0.600 2.100 2.400 7.650 ;
        RECT 3.600 1.500 5.400 6.750 ;
        RECT 6.600 3.000 8.400 7.650 ;
        RECT 9.600 3.900 11.400 8.100 ;
        RECT 12.600 3.000 14.400 8.100 ;
        RECT 6.600 2.100 14.400 3.000 ;
  END
END OAI22X1
MACRO OR2X1
  CLASS CORE ;
  FOREIGN OR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 13.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 13.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.000 2.400 36.900 ;
        RECT 5.100 24.900 6.900 37.500 ;
        RECT 8.700 30.900 10.500 36.900 ;
        RECT 8.700 30.000 11.100 30.900 ;
        RECT 0.600 23.100 9.000 24.000 ;
        RECT 7.200 22.200 9.000 23.100 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 14.700 5.550 15.150 ;
        RECT 3.900 12.900 6.300 14.700 ;
        RECT 7.500 10.050 8.550 22.200 ;
        RECT 9.900 20.850 11.100 30.000 ;
        RECT 6.900 9.300 8.700 10.050 ;
        RECT 3.900 8.250 8.700 9.300 ;
        RECT 3.900 5.100 4.800 8.250 ;
        RECT 9.900 5.100 11.100 18.150 ;
        RECT 0.600 1.500 2.400 5.100 ;
        RECT 3.600 2.100 5.400 5.100 ;
        RECT 6.600 1.500 8.400 5.100 ;
        RECT 9.600 2.100 11.400 5.100 ;
  END
END OR2X1
MACRO OR2X2
  CLASS CORE ;
  FOREIGN OR2X2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 12.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 3.450 15.450 5.550 17.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 13.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 13.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 36.900 ;
        RECT 5.100 24.900 6.900 37.500 ;
        RECT 8.100 27.300 9.900 36.900 ;
        RECT 8.100 24.900 11.100 27.300 ;
        RECT 0.600 23.400 1.800 24.900 ;
        RECT 0.600 22.200 9.000 23.400 ;
        RECT 7.200 21.600 9.000 22.200 ;
        RECT 0.750 15.750 2.550 18.150 ;
        RECT 3.900 14.550 5.550 15.150 ;
        RECT 3.900 12.750 6.300 14.550 ;
        RECT 7.200 10.800 8.550 21.600 ;
        RECT 9.900 20.850 11.100 24.900 ;
        RECT 7.200 10.050 9.000 10.800 ;
        RECT 3.900 9.000 9.000 10.050 ;
        RECT 3.900 5.100 4.800 9.000 ;
        RECT 9.900 8.100 11.100 18.150 ;
        RECT 0.600 2.100 2.400 5.100 ;
        RECT 3.600 2.100 5.400 5.100 ;
        RECT 0.600 1.500 1.800 2.100 ;
        RECT 6.600 1.500 8.400 7.500 ;
        RECT 9.600 2.100 11.400 8.100 ;
  END
END OR2X2
MACRO TBUFX1
  CLASS CORE ;
  FOREIGN TBUFX1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 15.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 12.450 18.450 14.550 20.550 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 6.450 18.450 8.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 16.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 16.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 1.200 30.900 3.000 37.500 ;
        RECT 4.200 30.900 6.000 36.900 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 0.900 15.750 3.300 17.550 ;
        RECT 4.350 12.000 5.550 30.900 ;
        RECT 7.500 26.850 9.300 36.900 ;
        RECT 6.900 24.900 9.300 26.850 ;
        RECT 12.000 24.900 13.800 37.500 ;
        RECT 6.900 20.850 8.100 24.900 ;
        RECT 6.900 14.400 8.100 18.150 ;
        RECT 12.450 17.550 14.100 18.150 ;
        RECT 12.300 15.750 14.100 17.550 ;
        RECT 6.900 13.050 8.850 14.400 ;
        RECT 4.350 10.200 6.900 12.000 ;
        RECT 4.350 5.100 6.000 10.200 ;
        RECT 7.800 8.100 8.850 13.050 ;
        RECT 1.200 1.500 3.000 5.100 ;
        RECT 4.200 2.100 6.000 5.100 ;
        RECT 7.500 2.100 9.300 8.100 ;
        RECT 12.000 1.500 13.800 8.100 ;
  END
END TBUFX1
MACRO TBUFX2
  CLASS CORE ;
  FOREIGN TBUFX2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 21.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 18.450 18.450 20.550 20.550 ;
    END
  END A
  PIN EN
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END EN
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 22.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 22.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 24.900 2.400 37.500 ;
        RECT 3.600 24.900 5.400 36.900 ;
        RECT 6.600 36.000 14.400 36.900 ;
        RECT 6.600 24.900 8.400 36.000 ;
        RECT 9.600 24.900 11.400 35.100 ;
        RECT 12.600 26.100 14.400 36.000 ;
        RECT 15.600 27.000 17.400 37.500 ;
        RECT 18.600 26.100 20.400 36.900 ;
        RECT 12.600 24.900 20.400 26.100 ;
        RECT 4.500 22.200 5.400 24.900 ;
        RECT 4.500 20.400 6.300 22.200 ;
        RECT 9.900 20.850 11.100 24.900 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 4.500 8.100 5.400 20.400 ;
        RECT 9.900 8.100 11.100 18.150 ;
        RECT 18.450 17.550 20.100 18.150 ;
        RECT 18.300 15.750 20.100 17.550 ;
        RECT 12.600 8.100 19.800 9.000 ;
        RECT 0.600 1.500 2.400 8.100 ;
        RECT 3.600 2.100 5.400 8.100 ;
        RECT 6.600 3.000 8.400 8.100 ;
        RECT 9.600 3.900 11.400 8.100 ;
        RECT 12.600 3.000 14.400 8.100 ;
        RECT 6.600 2.100 14.400 3.000 ;
        RECT 15.600 1.500 17.400 7.200 ;
        RECT 18.600 2.100 20.400 8.100 ;
  END
END TBUFX2
MACRO XNOR2X1
  CLASS CORE ;
  FOREIGN XNOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 18.450 17.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
    PORT
      LAYER metal1 ;
        RECT 8.850 18.450 9.150 19.800 ;
        RECT 8.850 18.150 9.450 18.450 ;
        RECT 8.850 8.850 9.750 18.150 ;
        RECT 8.850 8.550 9.450 8.850 ;
        RECT 8.850 7.500 9.150 8.550 ;
        RECT 7.950 6.450 9.150 7.500 ;
        RECT 9.450 6.450 11.550 8.550 ;
        RECT 7.950 6.150 9.450 6.450 ;
        RECT 7.950 2.100 9.750 6.150 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 19.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 19.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 25.950 2.400 36.900 ;
        RECT 3.600 27.000 5.550 37.500 ;
        RECT 8.100 25.950 9.900 36.900 ;
        RECT 12.450 27.000 14.400 37.500 ;
        RECT 15.600 26.100 17.400 36.900 ;
        RECT 0.600 24.600 5.400 25.950 ;
        RECT 8.100 24.900 11.100 25.950 ;
        RECT 3.300 23.850 5.400 24.600 ;
        RECT 3.300 22.950 8.550 23.850 ;
        RECT 6.750 21.000 8.550 22.950 ;
        RECT 9.900 20.850 11.100 24.900 ;
        RECT 12.450 24.900 17.400 26.100 ;
        RECT 12.450 24.000 14.550 24.900 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 4.950 18.000 6.750 19.800 ;
        RECT 0.900 15.750 2.700 17.550 ;
        RECT 5.400 15.900 7.500 18.000 ;
        RECT 15.450 17.550 17.100 18.150 ;
        RECT 1.650 15.000 2.700 15.750 ;
        RECT 10.650 15.150 12.450 16.950 ;
        RECT 15.300 15.750 17.100 17.550 ;
        RECT 1.650 13.650 7.500 15.000 ;
        RECT 5.400 12.900 7.500 13.650 ;
        RECT 10.650 13.050 12.750 15.150 ;
        RECT 6.150 12.000 7.350 12.900 ;
        RECT 3.150 10.500 5.250 11.100 ;
        RECT 0.600 9.000 5.250 10.500 ;
        RECT 6.150 10.200 7.950 12.000 ;
        RECT 12.900 9.000 15.000 11.550 ;
        RECT 0.600 8.100 2.250 9.000 ;
        RECT 12.900 8.100 17.400 9.000 ;
        RECT 0.600 2.100 2.400 8.100 ;
        RECT 3.600 1.500 5.400 7.200 ;
        RECT 12.450 1.500 14.250 7.200 ;
        RECT 15.600 2.100 17.400 8.100 ;
      LAYER via1 ;
        RECT 3.150 9.000 5.250 11.100 ;
        RECT 12.900 9.450 15.000 11.550 ;
      LAYER metal2 ;
        RECT 3.300 23.850 5.400 25.950 ;
        RECT 12.450 24.000 14.550 26.100 ;
        RECT 3.450 11.100 4.350 23.850 ;
        RECT 5.400 17.250 7.500 18.000 ;
        RECT 13.500 17.250 14.550 24.000 ;
        RECT 5.400 16.200 14.550 17.250 ;
        RECT 5.400 15.900 7.500 16.200 ;
        RECT 5.400 14.850 7.500 15.000 ;
        RECT 10.650 14.850 12.750 15.150 ;
        RECT 5.400 13.350 12.750 14.850 ;
        RECT 5.400 12.900 7.500 13.350 ;
        RECT 10.650 13.050 12.750 13.350 ;
        RECT 13.650 11.550 14.550 16.200 ;
        RECT 3.150 9.000 5.250 11.100 ;
        RECT 12.900 9.450 15.000 11.550 ;
  END
END XNOR2X1
MACRO XOR2X1
  CLASS CORE ;
  FOREIGN XOR2X1 ;
  ORIGIN 0.000 0.000 ;
  SIZE 18.000 BY 39.000 ;
  SYMMETRY X Y ;
  SITE core ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 0.450 18.450 2.550 20.550 ;
    END
  END A
  PIN B
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 15.450 18.450 17.550 20.550 ;
    END
  END B
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER metal1 ;
        RECT 9.450 18.450 11.550 20.550 ;
    END
    PORT
      LAYER metal1 ;
        RECT 8.850 18.150 9.450 18.450 ;
        RECT 8.850 17.550 11.100 18.150 ;
        RECT 8.850 8.850 9.900 17.550 ;
        RECT 8.850 8.550 9.450 8.850 ;
        RECT 8.850 8.100 9.150 8.550 ;
        RECT 8.100 6.450 9.150 8.100 ;
        RECT 9.450 6.450 11.550 8.550 ;
        RECT 8.100 6.150 9.450 6.450 ;
        RECT 8.100 2.100 9.900 6.150 ;
    END
  END Y
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 37.800 19.050 40.200 ;
    END
  END vdd
  PIN gnd
    DIRECTION INOUT ;
    USE GROUND ;
    SHAPE ABUTMENT ;
    PORT
      LAYER metal1 ;
        RECT -1.050 -1.200 19.050 1.200 ;
    END
  END gnd
  OBS
      LAYER metal1 ;
        RECT 0.600 25.800 2.400 36.900 ;
        RECT 3.600 27.000 5.400 37.500 ;
        RECT 0.600 24.900 5.250 25.800 ;
        RECT 8.100 24.900 9.900 36.900 ;
        RECT 12.600 27.000 14.400 37.500 ;
        RECT 15.600 26.100 17.400 36.900 ;
        RECT 3.150 22.800 5.250 24.900 ;
        RECT 8.850 23.400 9.900 24.900 ;
        RECT 12.600 24.900 17.400 26.100 ;
        RECT 12.600 24.000 14.700 24.900 ;
        RECT 8.850 22.350 11.100 23.400 ;
        RECT 6.300 21.150 8.400 21.450 ;
        RECT 4.500 19.350 8.400 21.150 ;
        RECT 9.450 20.850 11.100 22.350 ;
        RECT 0.900 17.550 2.550 18.150 ;
        RECT 6.150 17.550 7.950 18.150 ;
        RECT 15.450 17.550 17.100 18.150 ;
        RECT 0.900 16.350 7.950 17.550 ;
        RECT 0.900 15.750 2.700 16.350 ;
        RECT 10.950 14.850 12.750 16.650 ;
        RECT 15.300 15.750 17.100 17.550 ;
        RECT 6.150 13.050 7.950 14.850 ;
        RECT 5.850 10.950 7.950 13.050 ;
        RECT 10.800 12.750 12.900 14.850 ;
        RECT 1.350 9.900 7.950 10.950 ;
        RECT 1.350 8.100 2.400 9.900 ;
        RECT 12.600 9.150 14.700 10.200 ;
        RECT 12.600 8.100 17.400 9.150 ;
        RECT 0.600 2.100 2.400 8.100 ;
        RECT 3.600 1.500 5.400 7.200 ;
        RECT 12.600 1.500 14.400 7.200 ;
        RECT 15.600 2.100 17.400 8.100 ;
      LAYER via1 ;
        RECT 6.300 19.350 8.400 21.450 ;
      LAYER metal2 ;
        RECT 3.150 22.800 5.250 24.900 ;
        RECT 12.600 24.000 14.700 26.100 ;
        RECT 3.900 13.050 4.800 22.800 ;
        RECT 6.300 19.350 8.400 21.450 ;
        RECT 7.500 17.700 8.400 19.350 ;
        RECT 13.800 17.700 14.700 24.000 ;
        RECT 7.500 16.800 14.700 17.700 ;
        RECT 10.800 13.950 12.900 14.850 ;
        RECT 7.050 13.050 12.900 13.950 ;
        RECT 3.900 12.900 12.900 13.050 ;
        RECT 3.900 12.000 7.950 12.900 ;
        RECT 10.800 12.750 12.900 12.900 ;
        RECT 5.850 10.950 7.950 12.000 ;
        RECT 13.800 10.200 14.700 16.800 ;
        RECT 12.600 8.100 14.700 10.200 ;
  END
END XOR2X1
END LIBRARY
