magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -56 -56 84 174
<< diffusion >>
rect 5 5 23 113
<< genericcontact >>
rect 11 98 17 104
rect 11 70 17 76
rect 11 42 17 48
rect 11 14 17 20
<< metal1 >>
rect 4 4 24 114
<< end >>
