magic
tech scmos
magscale 1 2
timestamp 1727503886
<< nwell >>
rect -6 152 246 272
<< ntransistor >>
rect 25 14 29 54
rect 45 14 49 34
rect 55 14 59 34
rect 77 14 81 34
rect 87 14 91 34
rect 109 14 113 34
rect 153 14 157 34
rect 161 14 165 34
rect 183 14 187 34
rect 193 14 197 34
rect 215 14 219 54
<< ptransistor >>
rect 25 166 29 246
rect 45 206 49 246
rect 61 206 65 246
rect 81 206 85 246
rect 93 206 97 246
rect 113 206 117 246
rect 157 206 161 246
rect 165 206 169 246
rect 185 226 189 246
rect 193 226 197 246
rect 215 166 219 246
<< ndiffusion >>
rect 23 14 25 54
rect 29 34 39 54
rect 202 34 215 54
rect 29 14 31 34
rect 43 14 45 34
rect 49 14 55 34
rect 59 14 63 34
rect 75 14 77 34
rect 81 14 87 34
rect 91 14 93 34
rect 105 14 109 34
rect 113 14 115 34
rect 151 14 153 34
rect 157 14 161 34
rect 165 14 167 34
rect 179 14 183 34
rect 187 14 193 34
rect 197 14 199 34
rect 211 14 215 34
rect 219 14 221 54
<< pdiffusion >>
rect 23 166 25 246
rect 29 206 31 246
rect 43 206 45 246
rect 49 206 61 246
rect 65 206 67 246
rect 79 206 81 246
rect 85 206 93 246
rect 97 206 99 246
rect 111 206 113 246
rect 117 206 119 246
rect 155 206 157 246
rect 161 206 165 246
rect 169 226 171 246
rect 183 226 185 246
rect 189 226 193 246
rect 197 226 201 246
rect 213 226 215 246
rect 169 206 180 226
rect 29 166 38 206
rect 206 166 215 226
rect 219 166 221 246
<< ndcontact >>
rect 11 14 23 54
rect 31 14 43 34
rect 63 14 75 34
rect 93 14 105 34
rect 115 14 127 34
rect 139 14 151 34
rect 167 14 179 34
rect 199 14 211 34
rect 221 14 233 54
<< pdcontact >>
rect 11 166 23 246
rect 31 206 43 246
rect 67 206 79 246
rect 99 206 111 246
rect 119 206 131 246
rect 143 206 155 246
rect 171 226 183 246
rect 201 226 213 246
rect 221 166 233 246
<< psubstratepcontact >>
rect 0 -6 240 6
<< nsubstratencontact >>
rect 0 254 240 266
<< polysilicon >>
rect 25 246 29 250
rect 45 246 49 250
rect 61 246 65 250
rect 81 246 85 250
rect 93 246 97 250
rect 113 246 117 250
rect 157 246 161 250
rect 165 246 169 250
rect 185 246 189 250
rect 193 246 197 250
rect 215 246 219 250
rect 25 103 29 166
rect 45 106 49 206
rect 61 138 65 206
rect 81 162 85 206
rect 93 200 97 206
rect 85 150 88 162
rect 61 133 68 138
rect 25 54 29 91
rect 45 34 49 94
rect 64 90 68 133
rect 84 70 88 150
rect 55 66 88 70
rect 55 34 59 66
rect 79 46 81 58
rect 93 52 97 188
rect 113 180 117 206
rect 157 202 161 206
rect 125 200 161 202
rect 137 198 161 200
rect 77 34 81 46
rect 87 40 89 42
rect 87 38 101 40
rect 87 34 91 38
rect 109 34 113 168
rect 125 42 129 188
rect 165 174 169 206
rect 185 186 189 226
rect 193 200 197 226
rect 193 196 201 200
rect 141 51 145 66
rect 163 59 167 174
rect 197 167 201 196
rect 193 161 201 167
rect 193 115 197 161
rect 215 154 219 166
rect 217 142 219 154
rect 163 55 187 59
rect 141 46 165 51
rect 125 38 157 42
rect 153 34 157 38
rect 161 34 165 46
rect 183 34 187 55
rect 193 34 197 103
rect 215 54 219 142
rect 25 10 29 14
rect 45 10 49 14
rect 55 10 59 14
rect 77 10 81 14
rect 87 10 91 14
rect 109 10 113 14
rect 153 10 157 14
rect 161 10 165 14
rect 183 10 187 14
rect 193 10 197 14
rect 215 10 219 14
<< polycontact >>
rect 93 188 105 200
rect 73 150 85 162
rect 24 91 36 103
rect 44 94 56 106
rect 64 78 76 90
rect 67 46 79 58
rect 105 168 117 180
rect 125 188 137 200
rect 89 40 101 52
rect 153 174 165 186
rect 177 174 189 186
rect 137 66 149 78
rect 205 142 217 154
rect 191 103 203 115
<< metal1 >>
rect 0 266 240 268
rect 0 252 240 254
rect 31 246 43 252
rect 99 246 111 252
rect 143 246 155 252
rect 201 246 213 252
rect 67 200 75 206
rect 119 200 131 206
rect 57 186 75 200
rect 105 193 125 200
rect 171 192 183 226
rect 67 180 75 186
rect 67 172 105 180
rect 123 176 153 182
rect 11 160 17 166
rect 123 162 129 176
rect 171 168 177 186
rect 11 152 73 160
rect 11 54 17 152
rect 85 156 129 162
rect 143 162 177 168
rect 56 103 83 106
rect 56 98 97 103
rect 30 86 36 91
rect 30 78 64 86
rect 143 78 149 162
rect 197 154 211 162
rect 225 117 233 166
rect 217 103 233 117
rect 69 70 137 78
rect 69 58 76 70
rect 225 54 233 103
rect 101 40 122 47
rect 50 34 57 40
rect 115 34 122 40
rect 172 40 183 48
rect 172 34 179 40
rect 50 28 63 34
rect 31 8 43 14
rect 93 8 105 14
rect 139 8 151 14
rect 199 8 211 14
rect 0 6 240 8
rect 0 -8 240 -6
<< m2contact >>
rect 43 186 57 200
rect 183 192 197 206
rect 23 103 37 117
rect 83 103 97 117
rect 183 154 197 168
rect 203 103 217 117
rect 43 40 57 54
rect 183 40 197 54
<< metal2 >>
rect 23 117 37 137
rect 48 54 56 186
rect 183 168 191 192
rect 83 117 97 137
rect 183 54 191 154
rect 203 83 217 103
<< m2p >>
rect 23 123 37 137
rect 83 123 97 137
rect 203 83 217 97
<< labels >>
rlabel metal2 83 123 97 137 0 D
port 0 nsew signal input
rlabel metal2 23 123 37 137 0 CLK
port 1 nsew clock input
rlabel metal2 203 83 217 97 0 Q
port 2 nsew signal output
rlabel metal1 0 266 240 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 254 240 266 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 252 240 254 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 0 6 240 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -6 240 6 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 0 -8 240 -6 0 gnd
port 4 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 240 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
