magic
tech scmos
magscale 1 2
timestamp 1700733945
<< checkpaint >>
rect -46 214 66 306
rect -46 -46 66 46
<< nwell >>
rect -13 154 33 272
<< psubstratepcontact >>
rect -6 -6 26 6
<< nsubstratencontact >>
rect -6 254 26 266
<< metal1 >>
rect -6 266 26 268
rect -6 252 26 254
rect -6 6 26 8
rect -6 -8 26 -6
<< m1p >>
rect -6 252 26 268
rect -6 -8 26 8
<< labels >>
rlabel nsubstratencontact 10 260 10 260 0 vdd
port 1 nsew power bidirectional abutment
rlabel psubstratepcontact 10 0 10 0 0 gnd
port 2 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 20 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
