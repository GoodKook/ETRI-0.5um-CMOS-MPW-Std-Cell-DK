VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 729.000 BY 699.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 684.300 726.300 686.700 ;
        RECT 717.300 614.700 726.300 684.300 ;
        RECT 0.600 612.300 726.300 614.700 ;
        RECT 717.300 542.700 726.300 612.300 ;
        RECT 0.600 540.300 726.300 542.700 ;
        RECT 717.300 470.700 726.300 540.300 ;
        RECT 0.600 468.300 726.300 470.700 ;
        RECT 717.300 398.700 726.300 468.300 ;
        RECT 0.600 396.300 726.300 398.700 ;
        RECT 717.300 326.700 726.300 396.300 ;
        RECT 0.600 324.300 726.300 326.700 ;
        RECT 717.300 254.700 726.300 324.300 ;
        RECT 0.600 252.300 726.300 254.700 ;
        RECT 717.300 182.700 726.300 252.300 ;
        RECT 0.600 180.300 726.300 182.700 ;
        RECT 717.300 110.700 726.300 180.300 ;
        RECT 0.600 108.300 726.300 110.700 ;
        RECT 717.300 38.700 726.300 108.300 ;
        RECT 0.600 36.300 726.300 38.700 ;
        RECT 717.300 0.300 726.300 36.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.300 650.700 -0.300 686.700 ;
        RECT -9.300 648.300 716.400 650.700 ;
        RECT -9.300 578.700 -0.300 648.300 ;
        RECT -9.300 576.300 716.400 578.700 ;
        RECT -9.300 506.700 -0.300 576.300 ;
        RECT -9.300 504.300 716.400 506.700 ;
        RECT -9.300 434.700 -0.300 504.300 ;
        RECT -9.300 432.300 716.400 434.700 ;
        RECT -9.300 362.700 -0.300 432.300 ;
        RECT -9.300 360.300 716.400 362.700 ;
        RECT -9.300 290.700 -0.300 360.300 ;
        RECT -9.300 288.300 716.400 290.700 ;
        RECT -9.300 218.700 -0.300 288.300 ;
        RECT -9.300 216.300 716.400 218.700 ;
        RECT -9.300 146.700 -0.300 216.300 ;
        RECT -9.300 144.300 716.400 146.700 ;
        RECT -9.300 74.700 -0.300 144.300 ;
        RECT -9.300 72.300 716.400 74.700 ;
        RECT -9.300 2.700 -0.300 72.300 ;
        RECT -9.300 0.300 716.400 2.700 ;
    END
  END vdd
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 214.950 207.450 217.050 208.050 ;
        RECT 212.550 206.550 217.050 207.450 ;
        RECT 212.550 195.450 213.450 206.550 ;
        RECT 214.950 205.950 217.050 206.550 ;
        RECT 214.950 195.450 217.050 196.050 ;
        RECT 212.550 194.550 217.050 195.450 ;
        RECT 214.950 193.950 217.050 194.550 ;
        RECT 145.950 28.950 148.050 31.050 ;
        RECT 146.550 19.050 147.450 28.950 ;
        RECT 145.950 16.950 148.050 19.050 ;
      LAYER metal2 ;
        RECT 208.950 451.950 211.050 454.050 ;
        RECT 209.400 448.050 210.450 451.950 ;
        RECT 217.950 448.950 220.050 451.050 ;
        RECT 218.400 448.050 219.450 448.950 ;
        RECT 208.950 445.950 211.050 448.050 ;
        RECT 217.950 445.950 220.050 448.050 ;
        RECT 209.400 399.450 210.450 445.950 ;
        RECT 209.400 398.400 213.450 399.450 ;
        RECT 208.950 376.950 211.050 379.050 ;
        RECT 209.400 376.050 210.450 376.950 ;
        RECT 212.400 376.050 213.450 398.400 ;
        RECT 208.950 373.950 211.050 376.050 ;
        RECT 211.950 373.950 214.050 376.050 ;
        RECT 238.950 373.950 241.050 376.050 ;
        RECT 239.400 244.050 240.450 373.950 ;
        RECT 229.950 241.950 232.050 244.050 ;
        RECT 238.950 241.950 241.050 244.050 ;
        RECT 230.400 214.050 231.450 241.950 ;
        RECT 214.950 211.950 217.050 214.050 ;
        RECT 229.950 211.950 232.050 214.050 ;
        RECT 215.400 208.050 216.450 211.950 ;
        RECT 214.950 205.950 217.050 208.050 ;
        RECT 214.950 193.950 217.050 196.050 ;
        RECT 215.400 183.450 216.450 193.950 ;
        RECT 215.400 182.400 219.450 183.450 ;
        RECT 218.400 163.050 219.450 182.400 ;
        RECT 211.950 160.950 214.050 163.050 ;
        RECT 217.950 160.950 220.050 163.050 ;
        RECT 220.950 160.950 223.050 163.050 ;
        RECT 221.400 130.050 222.450 160.950 ;
        RECT 220.950 127.950 223.050 130.050 ;
        RECT 199.950 124.950 202.050 127.050 ;
        RECT 200.400 108.450 201.450 124.950 ;
        RECT 200.400 107.400 204.450 108.450 ;
        RECT 203.400 103.050 204.450 107.400 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 202.950 100.950 205.050 103.050 ;
        RECT 191.400 67.050 192.450 100.950 ;
        RECT 145.950 64.950 148.050 67.050 ;
        RECT 190.950 64.950 193.050 67.050 ;
        RECT 146.400 31.050 147.450 64.950 ;
        RECT 145.950 28.950 148.050 31.050 ;
        RECT 145.950 16.950 148.050 19.050 ;
        RECT 146.400 13.050 147.450 16.950 ;
        RECT 145.950 10.950 148.050 13.050 ;
        RECT 220.950 10.950 223.050 13.050 ;
        RECT 221.400 -3.600 222.450 10.950 ;
      LAYER metal3 ;
        RECT 208.950 447.600 211.050 448.050 ;
        RECT 217.950 447.600 220.050 448.050 ;
        RECT 208.950 446.400 220.050 447.600 ;
        RECT 208.950 445.950 211.050 446.400 ;
        RECT 217.950 445.950 220.050 446.400 ;
        RECT 208.950 375.600 211.050 376.050 ;
        RECT 211.950 375.600 214.050 376.050 ;
        RECT 238.950 375.600 241.050 376.050 ;
        RECT 208.950 374.400 241.050 375.600 ;
        RECT 208.950 373.950 211.050 374.400 ;
        RECT 211.950 373.950 214.050 374.400 ;
        RECT 238.950 373.950 241.050 374.400 ;
        RECT 229.950 243.600 232.050 244.050 ;
        RECT 238.950 243.600 241.050 244.050 ;
        RECT 229.950 242.400 241.050 243.600 ;
        RECT 229.950 241.950 232.050 242.400 ;
        RECT 238.950 241.950 241.050 242.400 ;
        RECT 214.950 213.600 217.050 214.050 ;
        RECT 229.950 213.600 232.050 214.050 ;
        RECT 214.950 212.400 232.050 213.600 ;
        RECT 214.950 211.950 217.050 212.400 ;
        RECT 229.950 211.950 232.050 212.400 ;
        RECT 211.950 162.600 214.050 163.050 ;
        RECT 217.950 162.600 220.050 163.050 ;
        RECT 220.950 162.600 223.050 163.050 ;
        RECT 211.950 161.400 223.050 162.600 ;
        RECT 211.950 160.950 214.050 161.400 ;
        RECT 217.950 160.950 220.050 161.400 ;
        RECT 220.950 160.950 223.050 161.400 ;
        RECT 220.950 129.600 223.050 130.050 ;
        RECT 209.400 128.400 223.050 129.600 ;
        RECT 199.950 126.600 202.050 127.050 ;
        RECT 209.400 126.600 210.600 128.400 ;
        RECT 220.950 127.950 223.050 128.400 ;
        RECT 199.950 125.400 210.600 126.600 ;
        RECT 199.950 124.950 202.050 125.400 ;
        RECT 190.950 102.600 193.050 103.050 ;
        RECT 202.950 102.600 205.050 103.050 ;
        RECT 190.950 101.400 205.050 102.600 ;
        RECT 190.950 100.950 193.050 101.400 ;
        RECT 202.950 100.950 205.050 101.400 ;
        RECT 145.950 66.600 148.050 67.050 ;
        RECT 190.950 66.600 193.050 67.050 ;
        RECT 145.950 65.400 193.050 66.600 ;
        RECT 145.950 64.950 148.050 65.400 ;
        RECT 190.950 64.950 193.050 65.400 ;
        RECT 145.950 12.600 148.050 13.050 ;
        RECT 220.950 12.600 223.050 13.050 ;
        RECT 145.950 11.400 223.050 12.600 ;
        RECT 145.950 10.950 148.050 11.400 ;
        RECT 220.950 10.950 223.050 11.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 334.950 94.950 337.050 97.050 ;
        RECT 331.950 84.450 334.050 85.050 ;
        RECT 335.550 84.450 336.450 94.950 ;
        RECT 331.950 83.550 336.450 84.450 ;
        RECT 331.950 82.950 334.050 83.550 ;
      LAYER metal2 ;
        RECT 175.950 493.950 178.050 496.050 ;
        RECT 274.950 493.950 277.050 496.050 ;
        RECT 176.400 490.050 177.450 493.950 ;
        RECT 275.400 490.050 276.450 493.950 ;
        RECT 142.950 487.950 145.050 490.050 ;
        RECT 157.950 487.950 160.050 490.050 ;
        RECT 175.950 487.950 178.050 490.050 ;
        RECT 274.950 487.950 277.050 490.050 ;
        RECT 130.950 484.950 133.050 487.050 ;
        RECT 283.950 481.950 286.050 484.050 ;
        RECT 284.400 468.450 285.450 481.950 ;
        RECT 284.400 467.400 288.450 468.450 ;
        RECT 127.950 448.950 130.050 451.050 ;
        RECT 229.950 448.950 232.050 451.050 ;
        RECT 128.400 427.050 129.450 448.950 ;
        RECT 230.400 448.050 231.450 448.950 ;
        RECT 229.950 445.950 232.050 448.050 ;
        RECT 235.950 445.950 238.050 448.050 ;
        RECT 236.400 427.050 237.450 445.950 ;
        RECT 287.400 427.050 288.450 467.400 ;
        RECT 127.950 424.950 130.050 427.050 ;
        RECT 133.950 424.950 136.050 427.050 ;
        RECT 235.950 424.950 238.050 427.050 ;
        RECT 286.950 424.950 289.050 427.050 ;
        RECT 134.400 418.050 135.450 424.950 ;
        RECT 133.950 415.950 136.050 418.050 ;
        RECT 236.400 352.050 237.450 424.950 ;
        RECT 220.950 349.950 223.050 352.050 ;
        RECT 235.950 349.950 238.050 352.050 ;
        RECT 221.400 333.450 222.450 349.950 ;
        RECT 218.400 332.400 222.450 333.450 ;
        RECT 218.400 289.050 219.450 332.400 ;
        RECT 208.950 286.950 211.050 289.050 ;
        RECT 217.950 286.950 220.050 289.050 ;
        RECT 209.400 211.050 210.450 286.950 ;
        RECT 187.950 208.950 190.050 211.050 ;
        RECT 208.950 208.950 211.050 211.050 ;
        RECT 211.950 208.950 214.050 211.050 ;
        RECT 232.950 208.950 235.050 211.050 ;
        RECT 188.400 202.050 189.450 208.950 ;
        RECT 187.950 199.950 190.050 202.050 ;
        RECT 212.400 169.050 213.450 208.950 ;
        RECT 233.400 202.050 234.450 208.950 ;
        RECT 232.950 199.950 235.050 202.050 ;
        RECT 211.950 166.950 214.050 169.050 ;
        RECT 223.950 163.950 226.050 166.050 ;
        RECT 224.400 148.050 225.450 163.950 ;
        RECT 223.950 145.950 226.050 148.050 ;
        RECT 262.950 145.950 265.050 148.050 ;
        RECT 263.400 130.050 264.450 145.950 ;
        RECT 235.950 127.950 238.050 130.050 ;
        RECT 262.950 127.950 265.050 130.050 ;
        RECT 280.950 127.950 283.050 130.050 ;
        RECT 281.400 103.050 282.450 127.950 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 335.400 97.050 336.450 100.950 ;
        RECT 334.950 94.950 337.050 97.050 ;
        RECT 331.950 82.950 334.050 85.050 ;
        RECT 332.400 58.050 333.450 82.950 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 314.400 51.450 315.450 55.950 ;
        RECT 314.400 50.400 318.450 51.450 ;
        RECT 317.400 10.050 318.450 50.400 ;
        RECT 262.950 7.950 265.050 10.050 ;
        RECT 316.950 7.950 319.050 10.050 ;
        RECT 263.400 -3.600 264.450 7.950 ;
      LAYER metal3 ;
        RECT 175.950 495.600 178.050 496.050 ;
        RECT 274.950 495.600 277.050 496.050 ;
        RECT 175.950 494.400 277.050 495.600 ;
        RECT 175.950 493.950 178.050 494.400 ;
        RECT 274.950 493.950 277.050 494.400 ;
        RECT 142.950 489.600 145.050 490.050 ;
        RECT 157.950 489.600 160.050 490.050 ;
        RECT 175.950 489.600 178.050 490.050 ;
        RECT 134.400 488.400 178.050 489.600 ;
        RECT 130.950 486.600 133.050 487.050 ;
        RECT 134.400 486.600 135.600 488.400 ;
        RECT 142.950 487.950 145.050 488.400 ;
        RECT 157.950 487.950 160.050 488.400 ;
        RECT 175.950 487.950 178.050 488.400 ;
        RECT 274.950 487.950 277.050 490.050 ;
        RECT 130.950 485.400 135.600 486.600 ;
        RECT 275.400 486.600 276.600 487.950 ;
        RECT 275.400 485.400 285.600 486.600 ;
        RECT 130.950 484.950 133.050 485.400 ;
        RECT 284.400 484.050 285.600 485.400 ;
        RECT 283.950 481.950 286.050 484.050 ;
        RECT 229.950 447.600 232.050 448.050 ;
        RECT 235.950 447.600 238.050 448.050 ;
        RECT 229.950 446.400 238.050 447.600 ;
        RECT 229.950 445.950 232.050 446.400 ;
        RECT 235.950 445.950 238.050 446.400 ;
        RECT 127.950 426.600 130.050 427.050 ;
        RECT 133.950 426.600 136.050 427.050 ;
        RECT 235.950 426.600 238.050 427.050 ;
        RECT 286.950 426.600 289.050 427.050 ;
        RECT 127.950 425.400 289.050 426.600 ;
        RECT 127.950 424.950 130.050 425.400 ;
        RECT 133.950 424.950 136.050 425.400 ;
        RECT 235.950 424.950 238.050 425.400 ;
        RECT 286.950 424.950 289.050 425.400 ;
        RECT 220.950 351.600 223.050 352.050 ;
        RECT 235.950 351.600 238.050 352.050 ;
        RECT 220.950 350.400 238.050 351.600 ;
        RECT 220.950 349.950 223.050 350.400 ;
        RECT 235.950 349.950 238.050 350.400 ;
        RECT 208.950 288.600 211.050 289.050 ;
        RECT 217.950 288.600 220.050 289.050 ;
        RECT 208.950 287.400 220.050 288.600 ;
        RECT 208.950 286.950 211.050 287.400 ;
        RECT 217.950 286.950 220.050 287.400 ;
        RECT 187.950 210.600 190.050 211.050 ;
        RECT 208.950 210.600 211.050 211.050 ;
        RECT 211.950 210.600 214.050 211.050 ;
        RECT 232.950 210.600 235.050 211.050 ;
        RECT 187.950 209.400 235.050 210.600 ;
        RECT 187.950 208.950 190.050 209.400 ;
        RECT 208.950 208.950 211.050 209.400 ;
        RECT 211.950 208.950 214.050 209.400 ;
        RECT 232.950 208.950 235.050 209.400 ;
        RECT 211.950 166.950 214.050 169.050 ;
        RECT 212.400 165.600 213.600 166.950 ;
        RECT 223.950 165.600 226.050 166.050 ;
        RECT 212.400 164.400 226.050 165.600 ;
        RECT 223.950 163.950 226.050 164.400 ;
        RECT 223.950 147.600 226.050 148.050 ;
        RECT 262.950 147.600 265.050 148.050 ;
        RECT 223.950 146.400 265.050 147.600 ;
        RECT 223.950 145.950 226.050 146.400 ;
        RECT 262.950 145.950 265.050 146.400 ;
        RECT 235.950 129.600 238.050 130.050 ;
        RECT 262.950 129.600 265.050 130.050 ;
        RECT 280.950 129.600 283.050 130.050 ;
        RECT 235.950 128.400 283.050 129.600 ;
        RECT 235.950 127.950 238.050 128.400 ;
        RECT 262.950 127.950 265.050 128.400 ;
        RECT 280.950 127.950 283.050 128.400 ;
        RECT 280.950 102.600 283.050 103.050 ;
        RECT 334.950 102.600 337.050 103.050 ;
        RECT 280.950 101.400 337.050 102.600 ;
        RECT 280.950 100.950 283.050 101.400 ;
        RECT 334.950 100.950 337.050 101.400 ;
        RECT 313.950 57.600 316.050 58.050 ;
        RECT 331.950 57.600 334.050 58.050 ;
        RECT 313.950 56.400 334.050 57.600 ;
        RECT 313.950 55.950 316.050 56.400 ;
        RECT 331.950 55.950 334.050 56.400 ;
        RECT 262.950 9.600 265.050 10.050 ;
        RECT 316.950 9.600 319.050 10.050 ;
        RECT 262.950 8.400 319.050 9.600 ;
        RECT 262.950 7.950 265.050 8.400 ;
        RECT 316.950 7.950 319.050 8.400 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 256.950 495.450 259.050 496.050 ;
        RECT 265.950 495.450 268.050 496.050 ;
        RECT 256.950 494.550 268.050 495.450 ;
        RECT 256.950 493.950 259.050 494.550 ;
        RECT 265.950 493.950 268.050 494.550 ;
      LAYER metal2 ;
        RECT 268.950 505.950 271.050 508.050 ;
        RECT 295.950 505.950 298.050 508.050 ;
        RECT 256.950 502.950 259.050 505.050 ;
        RECT 169.950 499.950 172.050 502.050 ;
        RECT 170.400 496.050 171.450 499.950 ;
        RECT 257.400 496.050 258.450 502.950 ;
        RECT 124.950 493.950 127.050 496.050 ;
        RECT 169.950 493.950 172.050 496.050 ;
        RECT 256.950 493.950 259.050 496.050 ;
        RECT 265.950 495.450 268.050 496.050 ;
        RECT 269.400 495.450 270.450 505.950 ;
        RECT 265.950 494.400 270.450 495.450 ;
        RECT 265.950 493.950 268.050 494.400 ;
        RECT 125.400 487.050 126.450 493.950 ;
        RECT 170.400 490.050 171.450 493.950 ;
        RECT 296.400 490.050 297.450 505.950 ;
        RECT 169.950 487.950 172.050 490.050 ;
        RECT 283.950 487.950 286.050 490.050 ;
        RECT 295.950 487.950 298.050 490.050 ;
        RECT 124.950 484.950 127.050 487.050 ;
        RECT 304.950 481.950 307.050 484.050 ;
        RECT 305.400 471.450 306.450 481.950 ;
        RECT 302.400 470.400 306.450 471.450 ;
        RECT 196.950 448.950 199.050 451.050 ;
        RECT 197.400 424.050 198.450 448.950 ;
        RECT 302.400 445.050 303.450 470.400 ;
        RECT 241.950 442.950 244.050 445.050 ;
        RECT 301.950 442.950 304.050 445.050 ;
        RECT 242.400 424.050 243.450 442.950 ;
        RECT 196.950 421.950 199.050 424.050 ;
        RECT 241.950 421.950 244.050 424.050 ;
        RECT 121.950 415.950 124.050 418.050 ;
        RECT 142.950 415.950 145.050 418.050 ;
        RECT 143.400 391.050 144.450 415.950 ;
        RECT 197.400 400.050 198.450 421.950 ;
        RECT 163.950 397.950 166.050 400.050 ;
        RECT 196.950 397.950 199.050 400.050 ;
        RECT 164.400 391.050 165.450 397.950 ;
        RECT 142.950 388.950 145.050 391.050 ;
        RECT 163.950 388.950 166.050 391.050 ;
        RECT 164.400 346.050 165.450 388.950 ;
        RECT 148.950 343.950 151.050 346.050 ;
        RECT 163.950 343.950 166.050 346.050 ;
        RECT 187.950 343.950 190.050 346.050 ;
        RECT 188.400 334.050 189.450 343.950 ;
        RECT 172.950 331.950 175.050 334.050 ;
        RECT 187.950 331.950 190.050 334.050 ;
        RECT 173.400 313.050 174.450 331.950 ;
        RECT 172.950 310.950 175.050 313.050 ;
        RECT 193.950 301.950 196.050 304.050 ;
        RECT 194.400 277.050 195.450 301.950 ;
        RECT 193.950 274.950 196.050 277.050 ;
        RECT 256.950 274.950 259.050 277.050 ;
        RECT 257.400 271.050 258.450 274.950 ;
        RECT 256.950 268.950 259.050 271.050 ;
        RECT 268.950 268.950 271.050 271.050 ;
        RECT 269.400 264.450 270.450 268.950 ;
        RECT 269.400 263.400 273.450 264.450 ;
        RECT 272.400 241.050 273.450 263.400 ;
        RECT 271.950 238.950 274.050 241.050 ;
        RECT 274.950 232.950 277.050 235.050 ;
        RECT 275.400 211.050 276.450 232.950 ;
        RECT 259.950 208.950 262.050 211.050 ;
        RECT 274.950 208.950 277.050 211.050 ;
        RECT 277.950 208.950 280.050 211.050 ;
        RECT 260.400 202.050 261.450 208.950 ;
        RECT 124.950 199.950 127.050 202.050 ;
        RECT 259.950 199.950 262.050 202.050 ;
        RECT 124.950 193.950 127.050 196.050 ;
        RECT 125.400 175.050 126.450 193.950 ;
        RECT 278.400 184.050 279.450 208.950 ;
        RECT 277.950 181.950 280.050 184.050 ;
        RECT 301.950 181.950 304.050 184.050 ;
        RECT 124.950 172.950 127.050 175.050 ;
        RECT 133.950 172.950 136.050 175.050 ;
        RECT 134.400 160.050 135.450 172.950 ;
        RECT 196.950 160.950 199.050 163.050 ;
        RECT 197.400 160.050 198.450 160.950 ;
        RECT 133.950 157.950 136.050 160.050 ;
        RECT 196.950 157.950 199.050 160.050 ;
        RECT 208.950 157.950 211.050 160.050 ;
        RECT 209.400 136.050 210.450 157.950 ;
        RECT 302.400 154.050 303.450 181.950 ;
        RECT 244.950 151.950 247.050 154.050 ;
        RECT 283.950 151.950 286.050 154.050 ;
        RECT 301.950 151.950 304.050 154.050 ;
        RECT 245.400 136.050 246.450 151.950 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 217.950 133.950 220.050 136.050 ;
        RECT 244.950 133.950 247.050 136.050 ;
        RECT 218.400 100.050 219.450 133.950 ;
        RECT 284.400 130.050 285.450 151.950 ;
        RECT 283.950 127.950 286.050 130.050 ;
        RECT 217.950 97.950 220.050 100.050 ;
        RECT 226.950 97.950 229.050 100.050 ;
        RECT 227.400 82.050 228.450 97.950 ;
        RECT 226.950 79.950 229.050 82.050 ;
        RECT 247.950 79.950 250.050 82.050 ;
        RECT 248.400 61.050 249.450 79.950 ;
        RECT 247.950 58.950 250.050 61.050 ;
        RECT 271.950 49.950 274.050 52.050 ;
        RECT 272.400 19.050 273.450 49.950 ;
        RECT 271.950 16.950 274.050 19.050 ;
        RECT 283.950 16.950 286.050 19.050 ;
        RECT 284.400 -3.600 285.450 16.950 ;
      LAYER metal3 ;
        RECT 268.950 507.600 271.050 508.050 ;
        RECT 295.950 507.600 298.050 508.050 ;
        RECT 268.950 506.400 298.050 507.600 ;
        RECT 268.950 505.950 271.050 506.400 ;
        RECT 295.950 505.950 298.050 506.400 ;
        RECT 256.950 504.600 259.050 505.050 ;
        RECT 209.400 503.400 259.050 504.600 ;
        RECT 169.950 501.600 172.050 502.050 ;
        RECT 209.400 501.600 210.600 503.400 ;
        RECT 256.950 502.950 259.050 503.400 ;
        RECT 169.950 500.400 210.600 501.600 ;
        RECT 169.950 499.950 172.050 500.400 ;
        RECT 124.950 495.600 127.050 496.050 ;
        RECT 169.950 495.600 172.050 496.050 ;
        RECT 124.950 494.400 172.050 495.600 ;
        RECT 124.950 493.950 127.050 494.400 ;
        RECT 169.950 493.950 172.050 494.400 ;
        RECT 283.950 489.600 286.050 490.050 ;
        RECT 295.950 489.600 298.050 490.050 ;
        RECT 283.950 488.400 298.050 489.600 ;
        RECT 283.950 487.950 286.050 488.400 ;
        RECT 287.400 486.600 288.600 488.400 ;
        RECT 295.950 487.950 298.050 488.400 ;
        RECT 287.400 485.400 306.600 486.600 ;
        RECT 305.400 484.050 306.600 485.400 ;
        RECT 304.950 481.950 307.050 484.050 ;
        RECT 241.950 444.600 244.050 445.050 ;
        RECT 301.950 444.600 304.050 445.050 ;
        RECT 241.950 443.400 304.050 444.600 ;
        RECT 241.950 442.950 244.050 443.400 ;
        RECT 301.950 442.950 304.050 443.400 ;
        RECT 196.950 423.600 199.050 424.050 ;
        RECT 241.950 423.600 244.050 424.050 ;
        RECT 196.950 422.400 244.050 423.600 ;
        RECT 196.950 421.950 199.050 422.400 ;
        RECT 241.950 421.950 244.050 422.400 ;
        RECT 121.950 417.600 124.050 418.050 ;
        RECT 142.950 417.600 145.050 418.050 ;
        RECT 121.950 416.400 145.050 417.600 ;
        RECT 121.950 415.950 124.050 416.400 ;
        RECT 142.950 415.950 145.050 416.400 ;
        RECT 163.950 399.600 166.050 400.050 ;
        RECT 196.950 399.600 199.050 400.050 ;
        RECT 163.950 398.400 199.050 399.600 ;
        RECT 163.950 397.950 166.050 398.400 ;
        RECT 196.950 397.950 199.050 398.400 ;
        RECT 142.950 390.600 145.050 391.050 ;
        RECT 163.950 390.600 166.050 391.050 ;
        RECT 142.950 389.400 166.050 390.600 ;
        RECT 142.950 388.950 145.050 389.400 ;
        RECT 163.950 388.950 166.050 389.400 ;
        RECT 148.950 345.600 151.050 346.050 ;
        RECT 163.950 345.600 166.050 346.050 ;
        RECT 187.950 345.600 190.050 346.050 ;
        RECT 148.950 344.400 190.050 345.600 ;
        RECT 148.950 343.950 151.050 344.400 ;
        RECT 163.950 343.950 166.050 344.400 ;
        RECT 187.950 343.950 190.050 344.400 ;
        RECT 172.950 333.600 175.050 334.050 ;
        RECT 187.950 333.600 190.050 334.050 ;
        RECT 172.950 332.400 190.050 333.600 ;
        RECT 172.950 331.950 175.050 332.400 ;
        RECT 187.950 331.950 190.050 332.400 ;
        RECT 172.950 312.600 175.050 313.050 ;
        RECT 167.400 311.400 175.050 312.600 ;
        RECT 167.400 303.600 168.600 311.400 ;
        RECT 172.950 310.950 175.050 311.400 ;
        RECT 193.950 303.600 196.050 304.050 ;
        RECT 167.400 302.400 196.050 303.600 ;
        RECT 193.950 301.950 196.050 302.400 ;
        RECT 193.950 276.600 196.050 277.050 ;
        RECT 256.950 276.600 259.050 277.050 ;
        RECT 193.950 275.400 259.050 276.600 ;
        RECT 193.950 274.950 196.050 275.400 ;
        RECT 256.950 274.950 259.050 275.400 ;
        RECT 256.950 270.600 259.050 271.050 ;
        RECT 268.950 270.600 271.050 271.050 ;
        RECT 256.950 269.400 271.050 270.600 ;
        RECT 256.950 268.950 259.050 269.400 ;
        RECT 268.950 268.950 271.050 269.400 ;
        RECT 271.950 238.950 274.050 241.050 ;
        RECT 272.400 234.600 273.600 238.950 ;
        RECT 274.950 234.600 277.050 235.050 ;
        RECT 272.400 233.400 277.050 234.600 ;
        RECT 274.950 232.950 277.050 233.400 ;
        RECT 259.950 210.600 262.050 211.050 ;
        RECT 274.950 210.600 277.050 211.050 ;
        RECT 277.950 210.600 280.050 211.050 ;
        RECT 259.950 209.400 280.050 210.600 ;
        RECT 259.950 208.950 262.050 209.400 ;
        RECT 274.950 208.950 277.050 209.400 ;
        RECT 277.950 208.950 280.050 209.400 ;
        RECT 124.950 199.950 127.050 202.050 ;
        RECT 125.400 196.050 126.600 199.950 ;
        RECT 124.950 193.950 127.050 196.050 ;
        RECT 277.950 183.600 280.050 184.050 ;
        RECT 301.950 183.600 304.050 184.050 ;
        RECT 277.950 182.400 304.050 183.600 ;
        RECT 277.950 181.950 280.050 182.400 ;
        RECT 301.950 181.950 304.050 182.400 ;
        RECT 124.950 174.600 127.050 175.050 ;
        RECT 133.950 174.600 136.050 175.050 ;
        RECT 124.950 173.400 136.050 174.600 ;
        RECT 124.950 172.950 127.050 173.400 ;
        RECT 133.950 172.950 136.050 173.400 ;
        RECT 133.950 159.600 136.050 160.050 ;
        RECT 196.950 159.600 199.050 160.050 ;
        RECT 208.950 159.600 211.050 160.050 ;
        RECT 133.950 158.400 211.050 159.600 ;
        RECT 133.950 157.950 136.050 158.400 ;
        RECT 196.950 157.950 199.050 158.400 ;
        RECT 208.950 157.950 211.050 158.400 ;
        RECT 244.950 153.600 247.050 154.050 ;
        RECT 283.950 153.600 286.050 154.050 ;
        RECT 301.950 153.600 304.050 154.050 ;
        RECT 244.950 152.400 304.050 153.600 ;
        RECT 244.950 151.950 247.050 152.400 ;
        RECT 283.950 151.950 286.050 152.400 ;
        RECT 301.950 151.950 304.050 152.400 ;
        RECT 224.400 137.400 240.600 138.600 ;
        RECT 208.950 135.600 211.050 136.050 ;
        RECT 217.950 135.600 220.050 136.050 ;
        RECT 224.400 135.600 225.600 137.400 ;
        RECT 208.950 134.400 225.600 135.600 ;
        RECT 239.400 135.600 240.600 137.400 ;
        RECT 244.950 135.600 247.050 136.050 ;
        RECT 239.400 134.400 247.050 135.600 ;
        RECT 208.950 133.950 211.050 134.400 ;
        RECT 217.950 133.950 220.050 134.400 ;
        RECT 244.950 133.950 247.050 134.400 ;
        RECT 217.950 99.600 220.050 100.050 ;
        RECT 226.950 99.600 229.050 100.050 ;
        RECT 217.950 98.400 229.050 99.600 ;
        RECT 217.950 97.950 220.050 98.400 ;
        RECT 226.950 97.950 229.050 98.400 ;
        RECT 226.950 81.600 229.050 82.050 ;
        RECT 247.950 81.600 250.050 82.050 ;
        RECT 226.950 80.400 250.050 81.600 ;
        RECT 226.950 79.950 229.050 80.400 ;
        RECT 247.950 79.950 250.050 80.400 ;
        RECT 247.950 60.600 250.050 61.050 ;
        RECT 247.950 59.400 270.600 60.600 ;
        RECT 247.950 58.950 250.050 59.400 ;
        RECT 269.400 57.600 270.600 59.400 ;
        RECT 269.400 56.400 273.600 57.600 ;
        RECT 272.400 52.050 273.600 56.400 ;
        RECT 271.950 49.950 274.050 52.050 ;
        RECT 271.950 18.600 274.050 19.050 ;
        RECT 283.950 18.600 286.050 19.050 ;
        RECT 271.950 17.400 286.050 18.600 ;
        RECT 271.950 16.950 274.050 17.400 ;
        RECT 283.950 16.950 286.050 17.400 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal2 ;
        RECT 49.950 490.950 52.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 118.950 490.950 121.050 493.050 ;
        RECT 50.400 487.050 51.450 490.950 ;
        RECT 59.400 490.050 60.450 490.950 ;
        RECT 58.950 487.950 61.050 490.050 ;
        RECT 49.950 484.950 52.050 487.050 ;
        RECT 119.400 481.050 120.450 490.950 ;
        RECT 109.950 478.950 112.050 481.050 ;
        RECT 118.950 478.950 121.050 481.050 ;
        RECT 110.400 427.050 111.450 478.950 ;
        RECT 91.950 424.950 94.050 427.050 ;
        RECT 109.950 424.950 112.050 427.050 ;
        RECT 92.400 418.050 93.450 424.950 ;
        RECT 91.950 415.950 94.050 418.050 ;
        RECT 110.400 417.450 111.450 424.950 ;
        RECT 107.400 416.400 111.450 417.450 ;
        RECT 107.400 388.050 108.450 416.400 ;
        RECT 106.950 385.950 109.050 388.050 ;
        RECT 103.950 376.950 106.050 379.050 ;
        RECT 104.400 354.450 105.450 376.950 ;
        RECT 101.400 353.400 105.450 354.450 ;
        RECT 101.400 343.050 102.450 353.400 ;
        RECT 100.950 340.950 103.050 343.050 ;
        RECT 100.950 331.950 103.050 334.050 ;
        RECT 101.400 289.050 102.450 331.950 ;
        RECT 100.950 286.950 103.050 289.050 ;
        RECT 115.950 286.950 118.050 289.050 ;
        RECT 116.400 267.450 117.450 286.950 ;
        RECT 116.400 266.400 120.450 267.450 ;
        RECT 119.400 241.050 120.450 266.400 ;
        RECT 118.950 238.950 121.050 241.050 ;
        RECT 106.950 235.950 109.050 238.050 ;
        RECT 107.400 208.050 108.450 235.950 ;
        RECT 58.950 205.950 61.050 208.050 ;
        RECT 106.950 205.950 109.050 208.050 ;
        RECT 59.400 202.050 60.450 205.950 ;
        RECT 49.950 199.950 52.050 202.050 ;
        RECT 58.950 199.950 61.050 202.050 ;
        RECT 55.950 193.950 58.050 196.050 ;
        RECT 56.400 178.050 57.450 193.950 ;
        RECT 55.950 175.950 58.050 178.050 ;
        RECT 88.950 175.950 91.050 178.050 ;
        RECT 89.400 127.050 90.450 175.950 ;
        RECT 88.950 124.950 91.050 127.050 ;
        RECT 94.950 118.950 97.050 121.050 ;
        RECT 95.400 97.050 96.450 118.950 ;
        RECT 94.950 94.950 97.050 97.050 ;
        RECT 40.950 85.950 43.050 88.050 ;
        RECT 76.950 85.950 79.050 88.050 ;
        RECT 41.400 58.050 42.450 85.950 ;
        RECT 77.400 76.050 78.450 85.950 ;
        RECT 76.950 73.950 79.050 76.050 ;
        RECT 91.950 73.950 94.050 76.050 ;
        RECT 160.950 73.950 163.050 76.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 92.400 31.050 93.450 73.950 ;
        RECT 161.400 58.050 162.450 73.950 ;
        RECT 160.950 55.950 163.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 298.950 55.950 301.050 58.050 ;
        RECT 91.950 28.950 94.050 31.050 ;
        RECT 127.950 28.950 130.050 31.050 ;
        RECT 128.400 7.050 129.450 28.950 ;
        RECT 280.950 16.950 283.050 19.050 ;
        RECT 281.400 7.050 282.450 16.950 ;
        RECT 290.400 7.050 291.450 55.950 ;
        RECT 127.950 4.950 130.050 7.050 ;
        RECT 280.950 4.950 283.050 7.050 ;
        RECT 289.950 4.950 292.050 7.050 ;
        RECT 290.400 -3.600 291.450 4.950 ;
      LAYER metal3 ;
        RECT 49.950 492.600 52.050 493.050 ;
        RECT 58.950 492.600 61.050 493.050 ;
        RECT 118.950 492.600 121.050 493.050 ;
        RECT 49.950 491.400 121.050 492.600 ;
        RECT 49.950 490.950 52.050 491.400 ;
        RECT 58.950 490.950 61.050 491.400 ;
        RECT 118.950 490.950 121.050 491.400 ;
        RECT 109.950 480.600 112.050 481.050 ;
        RECT 118.950 480.600 121.050 481.050 ;
        RECT 109.950 479.400 121.050 480.600 ;
        RECT 109.950 478.950 112.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 91.950 426.600 94.050 427.050 ;
        RECT 109.950 426.600 112.050 427.050 ;
        RECT 91.950 425.400 112.050 426.600 ;
        RECT 91.950 424.950 94.050 425.400 ;
        RECT 109.950 424.950 112.050 425.400 ;
        RECT 106.950 385.950 109.050 388.050 ;
        RECT 103.950 378.600 106.050 379.050 ;
        RECT 107.400 378.600 108.600 385.950 ;
        RECT 103.950 377.400 108.600 378.600 ;
        RECT 103.950 376.950 106.050 377.400 ;
        RECT 100.950 340.950 103.050 343.050 ;
        RECT 101.400 334.050 102.600 340.950 ;
        RECT 100.950 331.950 103.050 334.050 ;
        RECT 100.950 288.600 103.050 289.050 ;
        RECT 115.950 288.600 118.050 289.050 ;
        RECT 100.950 287.400 118.050 288.600 ;
        RECT 100.950 286.950 103.050 287.400 ;
        RECT 115.950 286.950 118.050 287.400 ;
        RECT 118.950 240.600 121.050 241.050 ;
        RECT 116.400 239.400 121.050 240.600 ;
        RECT 106.950 237.600 109.050 238.050 ;
        RECT 116.400 237.600 117.600 239.400 ;
        RECT 118.950 238.950 121.050 239.400 ;
        RECT 106.950 236.400 117.600 237.600 ;
        RECT 106.950 235.950 109.050 236.400 ;
        RECT 58.950 207.600 61.050 208.050 ;
        RECT 106.950 207.600 109.050 208.050 ;
        RECT 50.400 206.400 109.050 207.600 ;
        RECT 50.400 202.050 51.600 206.400 ;
        RECT 58.950 205.950 61.050 206.400 ;
        RECT 106.950 205.950 109.050 206.400 ;
        RECT 49.950 199.950 52.050 202.050 ;
        RECT 58.950 201.600 61.050 202.050 ;
        RECT 56.400 200.400 61.050 201.600 ;
        RECT 56.400 196.050 57.600 200.400 ;
        RECT 58.950 199.950 61.050 200.400 ;
        RECT 55.950 193.950 58.050 196.050 ;
        RECT 55.950 177.600 58.050 178.050 ;
        RECT 88.950 177.600 91.050 178.050 ;
        RECT 55.950 176.400 91.050 177.600 ;
        RECT 55.950 175.950 58.050 176.400 ;
        RECT 88.950 175.950 91.050 176.400 ;
        RECT 88.950 126.600 91.050 127.050 ;
        RECT 88.950 125.400 96.600 126.600 ;
        RECT 88.950 124.950 91.050 125.400 ;
        RECT 95.400 121.050 96.600 125.400 ;
        RECT 94.950 118.950 97.050 121.050 ;
        RECT 94.950 96.600 97.050 97.050 ;
        RECT 89.400 95.400 97.050 96.600 ;
        RECT 89.400 93.600 90.600 95.400 ;
        RECT 94.950 94.950 97.050 95.400 ;
        RECT 77.400 92.400 90.600 93.600 ;
        RECT 77.400 88.050 78.600 92.400 ;
        RECT 40.950 87.600 43.050 88.050 ;
        RECT 76.950 87.600 79.050 88.050 ;
        RECT 40.950 86.400 79.050 87.600 ;
        RECT 40.950 85.950 43.050 86.400 ;
        RECT 76.950 85.950 79.050 86.400 ;
        RECT 76.950 75.600 79.050 76.050 ;
        RECT 91.950 75.600 94.050 76.050 ;
        RECT 160.950 75.600 163.050 76.050 ;
        RECT 76.950 74.400 163.050 75.600 ;
        RECT 76.950 73.950 79.050 74.400 ;
        RECT 91.950 73.950 94.050 74.400 ;
        RECT 160.950 73.950 163.050 74.400 ;
        RECT 289.950 57.600 292.050 58.050 ;
        RECT 298.950 57.600 301.050 58.050 ;
        RECT 289.950 56.400 301.050 57.600 ;
        RECT 289.950 55.950 292.050 56.400 ;
        RECT 298.950 55.950 301.050 56.400 ;
        RECT 91.950 30.600 94.050 31.050 ;
        RECT 127.950 30.600 130.050 31.050 ;
        RECT 91.950 29.400 130.050 30.600 ;
        RECT 91.950 28.950 94.050 29.400 ;
        RECT 127.950 28.950 130.050 29.400 ;
        RECT 127.950 6.600 130.050 7.050 ;
        RECT 280.950 6.600 283.050 7.050 ;
        RECT 289.950 6.600 292.050 7.050 ;
        RECT 127.950 5.400 292.050 6.600 ;
        RECT 127.950 4.950 130.050 5.400 ;
        RECT 280.950 4.950 283.050 5.400 ;
        RECT 289.950 4.950 292.050 5.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal2 ;
        RECT 10.950 313.950 13.050 316.050 ;
        RECT 11.400 313.050 12.450 313.950 ;
        RECT 10.950 310.950 13.050 313.050 ;
        RECT 46.950 307.950 49.050 310.050 ;
        RECT 47.400 286.050 48.450 307.950 ;
        RECT 46.950 283.950 49.050 286.050 ;
        RECT 91.950 283.950 94.050 286.050 ;
        RECT 92.400 268.050 93.450 283.950 ;
        RECT 91.950 265.950 94.050 268.050 ;
        RECT 103.950 265.950 106.050 268.050 ;
        RECT 104.400 243.450 105.450 265.950 ;
        RECT 101.400 242.400 105.450 243.450 ;
        RECT 101.400 168.450 102.450 242.400 ;
        RECT 101.400 167.400 105.450 168.450 ;
        RECT 104.400 133.050 105.450 167.400 ;
        RECT 61.950 130.950 64.050 133.050 ;
        RECT 103.950 130.950 106.050 133.050 ;
        RECT 62.400 106.050 63.450 130.950 ;
        RECT 61.950 103.950 64.050 106.050 ;
        RECT 91.950 103.950 94.050 106.050 ;
        RECT 92.400 100.050 93.450 103.950 ;
        RECT 91.950 97.950 94.050 100.050 ;
        RECT 124.950 97.950 127.050 100.050 ;
        RECT 92.400 97.050 93.450 97.950 ;
        RECT 91.950 94.950 94.050 97.050 ;
        RECT 125.400 60.450 126.450 97.950 ;
        RECT 122.400 59.400 126.450 60.450 ;
        RECT 122.400 52.050 123.450 59.400 ;
        RECT 121.950 49.950 124.050 52.050 ;
        RECT 148.950 46.950 151.050 49.050 ;
        RECT 149.400 28.050 150.450 46.950 ;
        RECT 148.950 25.950 151.050 28.050 ;
        RECT 196.950 25.950 199.050 28.050 ;
        RECT 197.400 4.050 198.450 25.950 ;
        RECT 286.950 22.950 289.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 296.400 4.050 297.450 22.950 ;
        RECT 196.950 1.950 199.050 4.050 ;
        RECT 295.950 1.950 298.050 4.050 ;
        RECT 296.400 -3.600 297.450 1.950 ;
      LAYER metal3 ;
        RECT 10.950 315.600 13.050 316.050 ;
        RECT 10.950 314.400 48.600 315.600 ;
        RECT 10.950 313.950 13.050 314.400 ;
        RECT 47.400 310.050 48.600 314.400 ;
        RECT 46.950 307.950 49.050 310.050 ;
        RECT 46.950 285.600 49.050 286.050 ;
        RECT 91.950 285.600 94.050 286.050 ;
        RECT 46.950 284.400 94.050 285.600 ;
        RECT 46.950 283.950 49.050 284.400 ;
        RECT 91.950 283.950 94.050 284.400 ;
        RECT 91.950 267.600 94.050 268.050 ;
        RECT 103.950 267.600 106.050 268.050 ;
        RECT 91.950 266.400 106.050 267.600 ;
        RECT 91.950 265.950 94.050 266.400 ;
        RECT 103.950 265.950 106.050 266.400 ;
        RECT 61.950 132.600 64.050 133.050 ;
        RECT 103.950 132.600 106.050 133.050 ;
        RECT 61.950 131.400 106.050 132.600 ;
        RECT 61.950 130.950 64.050 131.400 ;
        RECT 103.950 130.950 106.050 131.400 ;
        RECT 61.950 105.600 64.050 106.050 ;
        RECT 91.950 105.600 94.050 106.050 ;
        RECT 61.950 104.400 94.050 105.600 ;
        RECT 61.950 103.950 64.050 104.400 ;
        RECT 91.950 103.950 94.050 104.400 ;
        RECT 91.950 99.600 94.050 100.050 ;
        RECT 124.950 99.600 127.050 100.050 ;
        RECT 91.950 98.400 127.050 99.600 ;
        RECT 91.950 97.950 94.050 98.400 ;
        RECT 124.950 97.950 127.050 98.400 ;
        RECT 121.950 51.600 124.050 52.050 ;
        RECT 121.950 50.400 144.600 51.600 ;
        RECT 121.950 49.950 124.050 50.400 ;
        RECT 143.400 48.600 144.600 50.400 ;
        RECT 148.950 48.600 151.050 49.050 ;
        RECT 143.400 47.400 151.050 48.600 ;
        RECT 148.950 46.950 151.050 47.400 ;
        RECT 148.950 27.600 151.050 28.050 ;
        RECT 196.950 27.600 199.050 28.050 ;
        RECT 148.950 26.400 199.050 27.600 ;
        RECT 148.950 25.950 151.050 26.400 ;
        RECT 196.950 25.950 199.050 26.400 ;
        RECT 286.950 24.600 289.050 25.050 ;
        RECT 295.950 24.600 298.050 25.050 ;
        RECT 286.950 23.400 298.050 24.600 ;
        RECT 286.950 22.950 289.050 23.400 ;
        RECT 295.950 22.950 298.050 23.400 ;
        RECT 196.950 3.600 199.050 4.050 ;
        RECT 295.950 3.600 298.050 4.050 ;
        RECT 196.950 2.400 298.050 3.600 ;
        RECT 196.950 1.950 199.050 2.400 ;
        RECT 295.950 1.950 298.050 2.400 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal1 ;
        RECT 313.950 58.950 316.050 61.050 ;
        RECT 314.550 49.050 315.450 58.950 ;
        RECT 313.950 46.950 316.050 49.050 ;
      LAYER metal2 ;
        RECT 76.950 240.450 79.050 241.050 ;
        RECT 76.950 239.400 81.450 240.450 ;
        RECT 76.950 238.950 79.050 239.400 ;
        RECT 80.400 234.450 81.450 239.400 ;
        RECT 77.400 233.400 81.450 234.450 ;
        RECT 77.400 199.050 78.450 233.400 ;
        RECT 76.950 196.950 79.050 199.050 ;
        RECT 73.950 190.950 76.050 193.050 ;
        RECT 74.400 160.050 75.450 190.950 ;
        RECT 73.950 157.950 76.050 160.050 ;
        RECT 79.950 157.950 82.050 160.050 ;
        RECT 70.950 121.950 73.050 124.050 ;
        RECT 71.400 112.050 72.450 121.950 ;
        RECT 80.400 112.050 81.450 157.950 ;
        RECT 70.950 109.950 73.050 112.050 ;
        RECT 79.950 109.950 82.050 112.050 ;
        RECT 82.950 109.950 85.050 112.050 ;
        RECT 115.950 109.950 118.050 112.050 ;
        RECT 83.400 85.050 84.450 109.950 ;
        RECT 116.400 99.450 117.450 109.950 ;
        RECT 116.400 98.400 120.450 99.450 ;
        RECT 119.400 97.050 120.450 98.400 ;
        RECT 118.950 94.950 121.050 97.050 ;
        RECT 82.950 82.950 85.050 85.050 ;
        RECT 313.950 82.950 316.050 85.050 ;
        RECT 314.400 61.050 315.450 82.950 ;
        RECT 313.950 58.950 316.050 61.050 ;
        RECT 313.950 46.950 316.050 49.050 ;
        RECT 314.400 31.050 315.450 46.950 ;
        RECT 313.950 28.950 316.050 31.050 ;
        RECT 322.950 28.950 325.050 31.050 ;
        RECT 314.400 25.050 315.450 28.950 ;
        RECT 313.950 22.950 316.050 25.050 ;
        RECT 323.400 4.050 324.450 28.950 ;
        RECT 316.950 1.950 319.050 4.050 ;
        RECT 322.950 1.950 325.050 4.050 ;
        RECT 317.400 -3.600 318.450 1.950 ;
      LAYER metal3 ;
        RECT 76.950 196.950 79.050 199.050 ;
        RECT 73.950 192.600 76.050 193.050 ;
        RECT 77.400 192.600 78.600 196.950 ;
        RECT 73.950 191.400 78.600 192.600 ;
        RECT 73.950 190.950 76.050 191.400 ;
        RECT 73.950 159.600 76.050 160.050 ;
        RECT 79.950 159.600 82.050 160.050 ;
        RECT 73.950 158.400 82.050 159.600 ;
        RECT 73.950 157.950 76.050 158.400 ;
        RECT 79.950 157.950 82.050 158.400 ;
        RECT 70.950 111.600 73.050 112.050 ;
        RECT 79.950 111.600 82.050 112.050 ;
        RECT 82.950 111.600 85.050 112.050 ;
        RECT 115.950 111.600 118.050 112.050 ;
        RECT 70.950 110.400 118.050 111.600 ;
        RECT 70.950 109.950 73.050 110.400 ;
        RECT 79.950 109.950 82.050 110.400 ;
        RECT 82.950 109.950 85.050 110.400 ;
        RECT 115.950 109.950 118.050 110.400 ;
        RECT 82.950 84.600 85.050 85.050 ;
        RECT 313.950 84.600 316.050 85.050 ;
        RECT 82.950 83.400 316.050 84.600 ;
        RECT 82.950 82.950 85.050 83.400 ;
        RECT 313.950 82.950 316.050 83.400 ;
        RECT 313.950 30.600 316.050 31.050 ;
        RECT 322.950 30.600 325.050 31.050 ;
        RECT 313.950 29.400 325.050 30.600 ;
        RECT 313.950 28.950 316.050 29.400 ;
        RECT 322.950 28.950 325.050 29.400 ;
        RECT 316.950 3.600 319.050 4.050 ;
        RECT 322.950 3.600 325.050 4.050 ;
        RECT 316.950 2.400 325.050 3.600 ;
        RECT 316.950 1.950 319.050 2.400 ;
        RECT 322.950 1.950 325.050 2.400 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 13.950 514.950 16.050 517.050 ;
        RECT 14.400 490.050 15.450 514.950 ;
        RECT 13.950 487.950 16.050 490.050 ;
        RECT 13.950 481.950 16.050 484.050 ;
      LAYER metal3 ;
        RECT -3.600 531.600 -2.400 534.600 ;
        RECT -6.600 530.400 -2.400 531.600 ;
        RECT -6.600 516.600 -5.400 530.400 ;
        RECT 13.950 516.600 16.050 517.050 ;
        RECT -6.600 515.400 16.050 516.600 ;
        RECT 13.950 514.950 16.050 515.400 ;
        RECT 13.950 487.950 16.050 490.050 ;
        RECT 14.400 484.050 15.600 487.950 ;
        RECT 13.950 481.950 16.050 484.050 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 611.400 673.050 612.450 693.450 ;
        RECT 610.950 670.950 613.050 673.050 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal2 ;
        RECT 55.950 523.950 58.050 526.050 ;
        RECT 56.400 520.050 57.450 523.950 ;
        RECT 61.950 520.950 64.050 523.050 ;
        RECT 100.950 520.950 103.050 523.050 ;
        RECT 62.400 520.050 63.450 520.950 ;
        RECT 101.400 520.050 102.450 520.950 ;
        RECT 55.950 517.950 58.050 520.050 ;
        RECT 61.950 517.950 64.050 520.050 ;
        RECT 100.950 517.950 103.050 520.050 ;
      LAYER metal3 ;
        RECT -3.600 525.600 -2.400 528.600 ;
        RECT 55.950 525.600 58.050 526.050 ;
        RECT -3.600 524.400 58.050 525.600 ;
        RECT 55.950 523.950 58.050 524.400 ;
        RECT 55.950 519.600 58.050 520.050 ;
        RECT 61.950 519.600 64.050 520.050 ;
        RECT 100.950 519.600 103.050 520.050 ;
        RECT 55.950 518.400 103.050 519.600 ;
        RECT 55.950 517.950 58.050 518.400 ;
        RECT 61.950 517.950 64.050 518.400 ;
        RECT 100.950 517.950 103.050 518.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal2 ;
        RECT 1.950 520.950 4.050 523.050 ;
        RECT 187.950 520.950 190.050 523.050 ;
        RECT 193.950 520.950 196.050 523.050 ;
        RECT 2.400 514.050 3.450 520.950 ;
        RECT 188.400 514.050 189.450 520.950 ;
        RECT 1.950 511.950 4.050 514.050 ;
        RECT 187.950 511.950 190.050 514.050 ;
      LAYER metal3 ;
        RECT 1.950 522.600 4.050 523.050 ;
        RECT -3.600 521.400 4.050 522.600 ;
        RECT 1.950 520.950 4.050 521.400 ;
        RECT 187.950 522.600 190.050 523.050 ;
        RECT 193.950 522.600 196.050 523.050 ;
        RECT 187.950 521.400 196.050 522.600 ;
        RECT 187.950 520.950 190.050 521.400 ;
        RECT 193.950 520.950 196.050 521.400 ;
        RECT 1.950 513.600 4.050 514.050 ;
        RECT 187.950 513.600 190.050 514.050 ;
        RECT 1.950 512.400 190.050 513.600 ;
        RECT 1.950 511.950 4.050 512.400 ;
        RECT 187.950 511.950 190.050 512.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal2 ;
        RECT 55.950 448.950 58.050 451.050 ;
        RECT 85.950 448.950 88.050 451.050 ;
        RECT 100.950 448.950 103.050 451.050 ;
        RECT 56.400 445.050 57.450 448.950 ;
        RECT 55.950 442.950 58.050 445.050 ;
      LAYER metal3 ;
        RECT 55.950 450.600 58.050 451.050 ;
        RECT 85.950 450.600 88.050 451.050 ;
        RECT 100.950 450.600 103.050 451.050 ;
        RECT -3.600 444.600 -2.400 450.600 ;
        RECT 55.950 449.400 103.050 450.600 ;
        RECT 55.950 448.950 58.050 449.400 ;
        RECT 85.950 448.950 88.050 449.400 ;
        RECT 100.950 448.950 103.050 449.400 ;
        RECT 55.950 444.600 58.050 445.050 ;
        RECT -3.600 443.400 58.050 444.600 ;
        RECT 55.950 442.950 58.050 443.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal2 ;
        RECT 157.950 421.950 160.050 424.050 ;
        RECT 169.950 421.950 172.050 424.050 ;
        RECT 158.400 418.050 159.450 421.950 ;
        RECT 157.950 415.950 160.050 418.050 ;
        RECT 170.400 403.050 171.450 421.950 ;
        RECT 169.950 400.950 172.050 403.050 ;
        RECT 220.950 400.950 223.050 403.050 ;
        RECT 221.400 385.050 222.450 400.950 ;
        RECT 220.950 382.950 223.050 385.050 ;
        RECT 226.950 376.950 229.050 379.050 ;
      LAYER metal3 ;
        RECT 157.950 423.600 160.050 424.050 ;
        RECT 169.950 423.600 172.050 424.050 ;
        RECT 157.950 422.400 172.050 423.600 ;
        RECT 157.950 421.950 160.050 422.400 ;
        RECT 169.950 421.950 172.050 422.400 ;
        RECT -3.600 402.600 -2.400 414.600 ;
        RECT 169.950 402.600 172.050 403.050 ;
        RECT 220.950 402.600 223.050 403.050 ;
        RECT -3.600 401.400 223.050 402.600 ;
        RECT 169.950 400.950 172.050 401.400 ;
        RECT 220.950 400.950 223.050 401.400 ;
        RECT 220.950 382.950 223.050 385.050 ;
        RECT 221.400 378.600 222.600 382.950 ;
        RECT 226.950 378.600 229.050 379.050 ;
        RECT 221.400 377.400 229.050 378.600 ;
        RECT 226.950 376.950 229.050 377.400 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 635.400 688.050 636.450 693.450 ;
        RECT 619.950 685.950 622.050 688.050 ;
        RECT 634.950 685.950 637.050 688.050 ;
        RECT 620.400 676.050 621.450 685.950 ;
        RECT 544.950 673.950 547.050 676.050 ;
        RECT 619.950 673.950 622.050 676.050 ;
        RECT 545.400 589.050 546.450 673.950 ;
        RECT 355.950 586.950 358.050 589.050 ;
        RECT 544.950 586.950 547.050 589.050 ;
        RECT 356.400 556.050 357.450 586.950 ;
        RECT 319.950 553.950 322.050 556.050 ;
        RECT 355.950 553.950 358.050 556.050 ;
      LAYER metal3 ;
        RECT 619.950 687.600 622.050 688.050 ;
        RECT 634.950 687.600 637.050 688.050 ;
        RECT 619.950 686.400 637.050 687.600 ;
        RECT 619.950 685.950 622.050 686.400 ;
        RECT 634.950 685.950 637.050 686.400 ;
        RECT 544.950 675.600 547.050 676.050 ;
        RECT 619.950 675.600 622.050 676.050 ;
        RECT 544.950 674.400 622.050 675.600 ;
        RECT 544.950 673.950 547.050 674.400 ;
        RECT 619.950 673.950 622.050 674.400 ;
        RECT 355.950 588.600 358.050 589.050 ;
        RECT 544.950 588.600 547.050 589.050 ;
        RECT 355.950 587.400 547.050 588.600 ;
        RECT 355.950 586.950 358.050 587.400 ;
        RECT 544.950 586.950 547.050 587.400 ;
        RECT 319.950 555.600 322.050 556.050 ;
        RECT 355.950 555.600 358.050 556.050 ;
        RECT 319.950 554.400 358.050 555.600 ;
        RECT 319.950 553.950 322.050 554.400 ;
        RECT 355.950 553.950 358.050 554.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal2 ;
        RECT 629.400 682.050 630.450 693.450 ;
        RECT 592.950 679.950 595.050 682.050 ;
        RECT 628.950 679.950 631.050 682.050 ;
        RECT 593.400 658.050 594.450 679.950 ;
        RECT 367.950 655.950 370.050 658.050 ;
        RECT 592.950 655.950 595.050 658.050 ;
        RECT 364.950 627.450 367.050 628.050 ;
        RECT 368.400 627.450 369.450 655.950 ;
        RECT 364.950 626.400 369.450 627.450 ;
        RECT 364.950 625.950 367.050 626.400 ;
      LAYER metal3 ;
        RECT 592.950 681.600 595.050 682.050 ;
        RECT 628.950 681.600 631.050 682.050 ;
        RECT 592.950 680.400 631.050 681.600 ;
        RECT 592.950 679.950 595.050 680.400 ;
        RECT 628.950 679.950 631.050 680.400 ;
        RECT 367.950 657.600 370.050 658.050 ;
        RECT 592.950 657.600 595.050 658.050 ;
        RECT 367.950 656.400 595.050 657.600 ;
        RECT 367.950 655.950 370.050 656.400 ;
        RECT 592.950 655.950 595.050 656.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal2 ;
        RECT 623.400 685.050 624.450 693.450 ;
        RECT 604.950 682.950 607.050 685.050 ;
        RECT 622.950 682.950 625.050 685.050 ;
        RECT 605.400 661.050 606.450 682.950 ;
        RECT 361.950 658.950 364.050 661.050 ;
        RECT 604.950 658.950 607.050 661.050 ;
        RECT 362.400 601.050 363.450 658.950 ;
        RECT 361.950 598.950 364.050 601.050 ;
      LAYER metal3 ;
        RECT 604.950 684.600 607.050 685.050 ;
        RECT 622.950 684.600 625.050 685.050 ;
        RECT 604.950 683.400 625.050 684.600 ;
        RECT 604.950 682.950 607.050 683.400 ;
        RECT 622.950 682.950 625.050 683.400 ;
        RECT 361.950 660.600 364.050 661.050 ;
        RECT 604.950 660.600 607.050 661.050 ;
        RECT 361.950 659.400 607.050 660.600 ;
        RECT 361.950 658.950 364.050 659.400 ;
        RECT 604.950 658.950 607.050 659.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal2 ;
        RECT 617.400 688.050 618.450 693.450 ;
        RECT 607.950 685.950 610.050 688.050 ;
        RECT 616.950 685.950 619.050 688.050 ;
        RECT 608.400 664.050 609.450 685.950 ;
        RECT 568.950 661.950 571.050 664.050 ;
        RECT 607.950 661.950 610.050 664.050 ;
        RECT 569.400 553.050 570.450 661.950 ;
        RECT 568.950 550.950 571.050 553.050 ;
        RECT 610.950 550.950 613.050 553.050 ;
        RECT 611.400 517.050 612.450 550.950 ;
        RECT 574.950 514.950 577.050 517.050 ;
        RECT 610.950 514.950 613.050 517.050 ;
        RECT 575.400 483.450 576.450 514.950 ;
        RECT 577.950 483.450 580.050 484.050 ;
        RECT 575.400 482.400 580.050 483.450 ;
        RECT 577.950 481.950 580.050 482.400 ;
      LAYER metal3 ;
        RECT 607.950 687.600 610.050 688.050 ;
        RECT 616.950 687.600 619.050 688.050 ;
        RECT 607.950 686.400 619.050 687.600 ;
        RECT 607.950 685.950 610.050 686.400 ;
        RECT 616.950 685.950 619.050 686.400 ;
        RECT 568.950 663.600 571.050 664.050 ;
        RECT 607.950 663.600 610.050 664.050 ;
        RECT 568.950 662.400 610.050 663.600 ;
        RECT 568.950 661.950 571.050 662.400 ;
        RECT 607.950 661.950 610.050 662.400 ;
        RECT 568.950 552.600 571.050 553.050 ;
        RECT 610.950 552.600 613.050 553.050 ;
        RECT 568.950 551.400 613.050 552.600 ;
        RECT 568.950 550.950 571.050 551.400 ;
        RECT 610.950 550.950 613.050 551.400 ;
        RECT 574.950 516.600 577.050 517.050 ;
        RECT 610.950 516.600 613.050 517.050 ;
        RECT 574.950 515.400 613.050 516.600 ;
        RECT 574.950 514.950 577.050 515.400 ;
        RECT 610.950 514.950 613.050 515.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal2 ;
        RECT 715.950 196.950 718.050 199.050 ;
        RECT 712.950 192.450 715.050 193.050 ;
        RECT 716.400 192.450 717.450 196.950 ;
        RECT 712.950 191.400 717.450 192.450 ;
        RECT 712.950 190.950 715.050 191.400 ;
      LAYER metal3 ;
        RECT 715.950 198.600 718.050 199.050 ;
        RECT 715.950 197.400 723.600 198.600 ;
        RECT 715.950 196.950 718.050 197.400 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal2 ;
        RECT 697.950 550.950 700.050 553.050 ;
        RECT 698.400 550.050 699.450 550.950 ;
        RECT 697.950 547.950 700.050 550.050 ;
      LAYER metal3 ;
        RECT 697.950 549.600 700.050 550.050 ;
        RECT 722.400 549.600 723.600 552.600 ;
        RECT 697.950 548.400 723.600 549.600 ;
        RECT 697.950 547.950 700.050 548.400 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal2 ;
        RECT 700.950 550.950 703.050 553.050 ;
      LAYER metal3 ;
        RECT 722.400 555.600 723.600 558.600 ;
        RECT 719.400 554.400 723.600 555.600 ;
        RECT 700.950 552.600 703.050 553.050 ;
        RECT 719.400 552.600 720.600 554.400 ;
        RECT 700.950 551.400 720.600 552.600 ;
        RECT 700.950 550.950 703.050 551.400 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 697.950 603.450 700.050 604.050 ;
        RECT 695.400 602.400 700.050 603.450 ;
        RECT 695.400 595.050 696.450 602.400 ;
        RECT 697.950 601.950 700.050 602.400 ;
        RECT 694.950 592.950 697.050 595.050 ;
      LAYER metal3 ;
        RECT 694.950 594.600 697.050 595.050 ;
        RECT 694.950 593.400 723.600 594.600 ;
        RECT 694.950 592.950 697.050 593.400 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 695.400 692.400 699.450 693.450 ;
        RECT 698.400 673.050 699.450 692.400 ;
        RECT 697.950 670.950 700.050 673.050 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal2 ;
        RECT 683.400 692.400 687.450 693.450 ;
        RECT 686.400 594.450 687.450 692.400 ;
        RECT 683.400 593.400 687.450 594.450 ;
        RECT 683.400 555.450 684.450 593.400 ;
        RECT 685.950 555.450 688.050 556.050 ;
        RECT 683.400 554.400 688.050 555.450 ;
        RECT 685.950 553.950 688.050 554.400 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 647.400 688.050 648.450 693.450 ;
        RECT 646.950 685.950 649.050 688.050 ;
        RECT 652.950 685.950 655.050 688.050 ;
        RECT 653.400 634.050 654.450 685.950 ;
        RECT 652.950 631.950 655.050 634.050 ;
        RECT 640.950 625.950 643.050 628.050 ;
      LAYER metal3 ;
        RECT 646.950 687.600 649.050 688.050 ;
        RECT 652.950 687.600 655.050 688.050 ;
        RECT 646.950 686.400 655.050 687.600 ;
        RECT 646.950 685.950 649.050 686.400 ;
        RECT 652.950 685.950 655.050 686.400 ;
        RECT 652.950 633.600 655.050 634.050 ;
        RECT 644.400 632.400 655.050 633.600 ;
        RECT 640.950 627.600 643.050 628.050 ;
        RECT 644.400 627.600 645.600 632.400 ;
        RECT 652.950 631.950 655.050 632.400 ;
        RECT 640.950 626.400 645.600 627.600 ;
        RECT 640.950 625.950 643.050 626.400 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal1 ;
        RECT 649.950 603.450 652.050 604.050 ;
        RECT 649.950 602.550 654.450 603.450 ;
        RECT 649.950 601.950 652.050 602.550 ;
        RECT 653.550 595.050 654.450 602.550 ;
        RECT 652.950 592.950 655.050 595.050 ;
      LAYER metal2 ;
        RECT 638.400 692.400 642.450 693.450 ;
        RECT 638.400 624.450 639.450 692.400 ;
        RECT 638.400 623.400 642.450 624.450 ;
        RECT 641.400 613.050 642.450 623.400 ;
        RECT 640.950 610.950 643.050 613.050 ;
        RECT 649.950 610.950 652.050 613.050 ;
        RECT 650.400 604.050 651.450 610.950 ;
        RECT 649.950 601.950 652.050 604.050 ;
        RECT 652.950 592.950 655.050 595.050 ;
        RECT 653.400 541.050 654.450 592.950 ;
        RECT 625.950 538.950 628.050 541.050 ;
        RECT 652.950 538.950 655.050 541.050 ;
        RECT 626.400 487.050 627.450 538.950 ;
        RECT 625.950 484.950 628.050 487.050 ;
        RECT 613.950 481.950 616.050 484.050 ;
      LAYER metal3 ;
        RECT 640.950 612.600 643.050 613.050 ;
        RECT 649.950 612.600 652.050 613.050 ;
        RECT 640.950 611.400 652.050 612.600 ;
        RECT 640.950 610.950 643.050 611.400 ;
        RECT 649.950 610.950 652.050 611.400 ;
        RECT 625.950 540.600 628.050 541.050 ;
        RECT 652.950 540.600 655.050 541.050 ;
        RECT 625.950 539.400 655.050 540.600 ;
        RECT 625.950 538.950 628.050 539.400 ;
        RECT 652.950 538.950 655.050 539.400 ;
        RECT 625.950 484.950 628.050 487.050 ;
        RECT 613.950 483.600 616.050 484.050 ;
        RECT 626.400 483.600 627.600 484.950 ;
        RECT 613.950 482.400 627.600 483.600 ;
        RECT 613.950 481.950 616.050 482.400 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal2 ;
        RECT 599.400 692.400 603.450 693.450 ;
        RECT 599.400 669.450 600.450 692.400 ;
        RECT 601.950 669.450 604.050 670.050 ;
        RECT 599.400 668.400 604.050 669.450 ;
        RECT 601.950 667.950 604.050 668.400 ;
        RECT 602.400 625.050 603.450 667.950 ;
        RECT 565.950 622.950 568.050 625.050 ;
        RECT 601.950 622.950 604.050 625.050 ;
        RECT 370.950 595.950 373.050 598.050 ;
        RECT 371.400 586.050 372.450 595.950 ;
        RECT 566.400 586.050 567.450 622.950 ;
        RECT 370.950 583.950 373.050 586.050 ;
        RECT 565.950 583.950 568.050 586.050 ;
        RECT 371.400 562.050 372.450 583.950 ;
        RECT 349.950 559.950 352.050 562.050 ;
        RECT 370.950 559.950 373.050 562.050 ;
        RECT 350.400 559.050 351.450 559.950 ;
        RECT 349.950 556.950 352.050 559.050 ;
        RECT 566.400 553.050 567.450 583.950 ;
        RECT 553.950 550.950 556.050 553.050 ;
        RECT 565.950 550.950 568.050 553.050 ;
        RECT 554.400 523.050 555.450 550.950 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 689.400 523.050 690.450 523.950 ;
        RECT 532.950 520.950 535.050 523.050 ;
        RECT 553.950 520.950 556.050 523.050 ;
        RECT 688.950 520.950 691.050 523.050 ;
        RECT 533.400 483.450 534.450 520.950 ;
        RECT 530.400 482.400 534.450 483.450 ;
        RECT 530.400 454.050 531.450 482.400 ;
        RECT 523.950 451.950 526.050 454.050 ;
        RECT 529.950 451.950 532.050 454.050 ;
        RECT 524.400 417.450 525.450 451.950 ;
        RECT 524.400 416.400 528.450 417.450 ;
        RECT 527.400 379.050 528.450 416.400 ;
        RECT 607.950 379.950 610.050 382.050 ;
        RECT 608.400 379.050 609.450 379.950 ;
        RECT 514.950 376.950 517.050 379.050 ;
        RECT 526.950 376.950 529.050 379.050 ;
        RECT 607.950 376.950 610.050 379.050 ;
        RECT 352.950 307.950 355.050 310.050 ;
        RECT 353.400 277.050 354.450 307.950 ;
        RECT 515.400 304.050 516.450 376.950 ;
        RECT 514.950 301.950 517.050 304.050 ;
        RECT 523.950 301.950 526.050 304.050 ;
        RECT 352.950 274.950 355.050 277.050 ;
        RECT 370.950 274.950 373.050 277.050 ;
        RECT 371.400 261.450 372.450 274.950 ;
        RECT 524.400 265.050 525.450 301.950 ;
        RECT 517.950 262.950 520.050 265.050 ;
        RECT 523.950 262.950 526.050 265.050 ;
        RECT 371.400 260.400 375.450 261.450 ;
        RECT 374.400 226.050 375.450 260.400 ;
        RECT 518.400 226.050 519.450 262.950 ;
        RECT 373.950 223.950 376.050 226.050 ;
        RECT 511.950 223.950 514.050 226.050 ;
        RECT 517.950 223.950 520.050 226.050 ;
        RECT 512.400 166.050 513.450 223.950 ;
        RECT 511.950 163.950 514.050 166.050 ;
        RECT 523.950 163.950 526.050 166.050 ;
        RECT 553.950 163.950 556.050 166.050 ;
      LAYER metal3 ;
        RECT 565.950 624.600 568.050 625.050 ;
        RECT 601.950 624.600 604.050 625.050 ;
        RECT 565.950 623.400 604.050 624.600 ;
        RECT 565.950 622.950 568.050 623.400 ;
        RECT 601.950 622.950 604.050 623.400 ;
        RECT 370.950 585.600 373.050 586.050 ;
        RECT 565.950 585.600 568.050 586.050 ;
        RECT 370.950 584.400 568.050 585.600 ;
        RECT 370.950 583.950 373.050 584.400 ;
        RECT 565.950 583.950 568.050 584.400 ;
        RECT 349.950 561.600 352.050 562.050 ;
        RECT 370.950 561.600 373.050 562.050 ;
        RECT 349.950 560.400 373.050 561.600 ;
        RECT 349.950 559.950 352.050 560.400 ;
        RECT 370.950 559.950 373.050 560.400 ;
        RECT 553.950 552.600 556.050 553.050 ;
        RECT 565.950 552.600 568.050 553.050 ;
        RECT 553.950 551.400 568.050 552.600 ;
        RECT 553.950 550.950 556.050 551.400 ;
        RECT 565.950 550.950 568.050 551.400 ;
        RECT 532.950 522.600 535.050 523.050 ;
        RECT 553.950 522.600 556.050 523.050 ;
        RECT 688.950 522.600 691.050 523.050 ;
        RECT 532.950 521.400 691.050 522.600 ;
        RECT 532.950 520.950 535.050 521.400 ;
        RECT 553.950 520.950 556.050 521.400 ;
        RECT 688.950 520.950 691.050 521.400 ;
        RECT 523.950 453.600 526.050 454.050 ;
        RECT 529.950 453.600 532.050 454.050 ;
        RECT 523.950 452.400 532.050 453.600 ;
        RECT 523.950 451.950 526.050 452.400 ;
        RECT 529.950 451.950 532.050 452.400 ;
        RECT 514.950 378.600 517.050 379.050 ;
        RECT 526.950 378.600 529.050 379.050 ;
        RECT 607.950 378.600 610.050 379.050 ;
        RECT 514.950 377.400 610.050 378.600 ;
        RECT 514.950 376.950 517.050 377.400 ;
        RECT 526.950 376.950 529.050 377.400 ;
        RECT 607.950 376.950 610.050 377.400 ;
        RECT 514.950 303.600 517.050 304.050 ;
        RECT 523.950 303.600 526.050 304.050 ;
        RECT 514.950 302.400 526.050 303.600 ;
        RECT 514.950 301.950 517.050 302.400 ;
        RECT 523.950 301.950 526.050 302.400 ;
        RECT 352.950 276.600 355.050 277.050 ;
        RECT 370.950 276.600 373.050 277.050 ;
        RECT 352.950 275.400 373.050 276.600 ;
        RECT 352.950 274.950 355.050 275.400 ;
        RECT 370.950 274.950 373.050 275.400 ;
        RECT 517.950 264.600 520.050 265.050 ;
        RECT 523.950 264.600 526.050 265.050 ;
        RECT 517.950 263.400 526.050 264.600 ;
        RECT 517.950 262.950 520.050 263.400 ;
        RECT 523.950 262.950 526.050 263.400 ;
        RECT 373.950 225.600 376.050 226.050 ;
        RECT 511.950 225.600 514.050 226.050 ;
        RECT 517.950 225.600 520.050 226.050 ;
        RECT 373.950 224.400 520.050 225.600 ;
        RECT 373.950 223.950 376.050 224.400 ;
        RECT 511.950 223.950 514.050 224.400 ;
        RECT 517.950 223.950 520.050 224.400 ;
        RECT 511.950 165.600 514.050 166.050 ;
        RECT 523.950 165.600 526.050 166.050 ;
        RECT 553.950 165.600 556.050 166.050 ;
        RECT 511.950 164.400 556.050 165.600 ;
        RECT 511.950 163.950 514.050 164.400 ;
        RECT 523.950 163.950 526.050 164.400 ;
        RECT 553.950 163.950 556.050 164.400 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 5.700 680.400 7.500 683.250 ;
        RECT 9.000 679.050 10.800 683.250 ;
        RECT 5.100 677.400 10.800 679.050 ;
        RECT 13.200 677.400 15.000 683.250 ;
        RECT 5.100 670.950 6.300 677.400 ;
        RECT 23.100 675.000 24.900 683.250 ;
        RECT 8.100 672.150 9.900 673.950 ;
        RECT 4.950 668.850 7.050 670.950 ;
        RECT 7.950 670.050 10.050 672.150 ;
        RECT 10.950 671.850 13.050 673.950 ;
        RECT 14.100 672.150 15.900 673.950 ;
        RECT 20.400 673.350 24.900 675.000 ;
        RECT 28.500 674.400 30.300 683.250 ;
        RECT 32.700 674.400 34.500 683.250 ;
        RECT 38.100 675.000 39.900 683.250 ;
        RECT 53.100 675.000 54.900 683.250 ;
        RECT 38.100 673.350 42.600 675.000 ;
        RECT 11.100 670.050 12.900 671.850 ;
        RECT 13.950 670.050 16.050 672.150 ;
        RECT 20.400 669.150 21.600 673.350 ;
        RECT 41.400 669.150 42.600 673.350 ;
        RECT 50.400 673.350 54.900 675.000 ;
        RECT 58.500 674.400 60.300 683.250 ;
        RECT 63.000 677.400 64.800 683.250 ;
        RECT 67.200 679.050 69.000 683.250 ;
        RECT 70.500 680.400 72.300 683.250 ;
        RECT 67.200 677.400 72.900 679.050 ;
        RECT 50.400 669.150 51.600 673.350 ;
        RECT 62.100 672.150 63.900 673.950 ;
        RECT 61.950 670.050 64.050 672.150 ;
        RECT 64.950 671.850 67.050 673.950 ;
        RECT 68.100 672.150 69.900 673.950 ;
        RECT 65.100 670.050 66.900 671.850 ;
        RECT 67.950 670.050 70.050 672.150 ;
        RECT 71.700 670.950 72.900 677.400 ;
        RECT 77.550 678.300 79.350 683.250 ;
        RECT 80.550 679.200 82.350 683.250 ;
        RECT 83.550 678.300 85.350 683.250 ;
        RECT 77.550 676.950 85.350 678.300 ;
        RECT 86.550 677.400 88.350 683.250 ;
        RECT 92.550 678.300 94.350 683.250 ;
        RECT 95.550 679.200 97.350 683.250 ;
        RECT 98.550 678.300 100.350 683.250 ;
        RECT 73.950 673.950 76.050 676.050 ;
        RECT 86.550 675.300 87.750 677.400 ;
        RECT 92.550 676.950 100.350 678.300 ;
        RECT 101.550 677.400 103.350 683.250 ;
        RECT 101.550 675.300 102.750 677.400 ;
        RECT 84.000 674.250 87.750 675.300 ;
        RECT 99.000 674.250 102.750 675.300 ;
        RECT 113.100 675.000 114.900 683.250 ;
        RECT 5.100 663.600 6.300 668.850 ;
        RECT 19.950 667.050 22.050 669.150 ;
        RECT 4.650 651.750 6.450 663.600 ;
        RECT 7.650 662.700 15.450 663.600 ;
        RECT 7.650 651.750 9.450 662.700 ;
        RECT 10.650 651.750 12.450 661.800 ;
        RECT 13.650 651.750 15.450 662.700 ;
        RECT 20.250 658.800 21.300 667.050 ;
        RECT 22.950 665.850 25.050 667.950 ;
        RECT 28.950 665.850 31.050 667.950 ;
        RECT 31.950 665.850 34.050 667.950 ;
        RECT 37.950 665.850 40.050 667.950 ;
        RECT 40.950 667.050 43.050 669.150 ;
        RECT 49.950 667.050 52.050 669.150 ;
        RECT 70.950 668.850 73.050 670.950 ;
        RECT 22.950 664.050 24.750 665.850 ;
        RECT 25.950 662.850 28.050 664.950 ;
        RECT 29.100 664.050 30.900 665.850 ;
        RECT 32.100 664.050 33.900 665.850 ;
        RECT 34.950 662.850 37.050 664.950 ;
        RECT 38.250 664.050 40.050 665.850 ;
        RECT 26.100 661.050 27.900 662.850 ;
        RECT 35.100 661.050 36.900 662.850 ;
        RECT 41.700 658.800 42.750 667.050 ;
        RECT 20.250 657.900 27.300 658.800 ;
        RECT 20.250 657.600 21.450 657.900 ;
        RECT 19.650 651.750 21.450 657.600 ;
        RECT 25.650 657.600 27.300 657.900 ;
        RECT 35.700 657.900 42.750 658.800 ;
        RECT 35.700 657.600 37.350 657.900 ;
        RECT 22.650 651.750 24.450 657.000 ;
        RECT 25.650 651.750 27.450 657.600 ;
        RECT 28.650 651.750 30.450 657.600 ;
        RECT 32.550 651.750 34.350 657.600 ;
        RECT 35.550 651.750 37.350 657.600 ;
        RECT 41.550 657.600 42.750 657.900 ;
        RECT 50.250 658.800 51.300 667.050 ;
        RECT 52.950 665.850 55.050 667.950 ;
        RECT 58.950 665.850 61.050 667.950 ;
        RECT 52.950 664.050 54.750 665.850 ;
        RECT 55.950 662.850 58.050 664.950 ;
        RECT 59.100 664.050 60.900 665.850 ;
        RECT 71.700 663.600 72.900 668.850 ;
        RECT 74.550 667.050 75.450 673.950 ;
        RECT 80.100 672.150 81.900 673.950 ;
        RECT 76.950 668.850 79.050 670.950 ;
        RECT 79.950 670.050 82.050 672.150 ;
        RECT 83.850 670.950 85.050 674.250 ;
        RECT 95.100 672.150 96.900 673.950 ;
        RECT 82.950 668.850 85.050 670.950 ;
        RECT 91.950 668.850 94.050 670.950 ;
        RECT 94.950 670.050 97.050 672.150 ;
        RECT 98.850 670.950 100.050 674.250 ;
        RECT 97.950 668.850 100.050 670.950 ;
        RECT 110.400 673.350 114.900 675.000 ;
        RECT 118.500 674.400 120.300 683.250 ;
        RECT 122.700 674.400 124.500 683.250 ;
        RECT 128.100 675.000 129.900 683.250 ;
        RECT 137.850 677.400 139.650 683.250 ;
        RECT 142.350 676.200 144.150 683.250 ;
        RECT 140.550 675.300 144.150 676.200 ;
        RECT 128.100 673.350 132.600 675.000 ;
        RECT 110.400 669.150 111.600 673.350 ;
        RECT 131.400 669.150 132.600 673.350 ;
        RECT 137.100 669.150 138.900 670.950 ;
        RECT 77.100 667.050 78.900 668.850 ;
        RECT 73.950 664.950 76.050 667.050 ;
        RECT 82.950 663.600 84.150 668.850 ;
        RECT 85.950 665.850 88.050 667.950 ;
        RECT 92.100 667.050 93.900 668.850 ;
        RECT 85.950 664.050 87.750 665.850 ;
        RECT 97.950 663.600 99.150 668.850 ;
        RECT 100.950 665.850 103.050 667.950 ;
        RECT 109.950 667.050 112.050 669.150 ;
        RECT 100.950 664.050 102.750 665.850 ;
        RECT 56.100 661.050 57.900 662.850 ;
        RECT 62.550 662.700 70.350 663.600 ;
        RECT 50.250 657.900 57.300 658.800 ;
        RECT 50.250 657.600 51.450 657.900 ;
        RECT 38.550 651.750 40.350 657.000 ;
        RECT 41.550 651.750 43.350 657.600 ;
        RECT 49.650 651.750 51.450 657.600 ;
        RECT 55.650 657.600 57.300 657.900 ;
        RECT 52.650 651.750 54.450 657.000 ;
        RECT 55.650 651.750 57.450 657.600 ;
        RECT 58.650 651.750 60.450 657.600 ;
        RECT 62.550 651.750 64.350 662.700 ;
        RECT 65.550 651.750 67.350 661.800 ;
        RECT 68.550 651.750 70.350 662.700 ;
        RECT 71.550 651.750 73.350 663.600 ;
        RECT 78.300 651.750 80.100 663.600 ;
        RECT 82.500 651.750 84.300 663.600 ;
        RECT 85.800 651.750 87.600 657.600 ;
        RECT 93.300 651.750 95.100 663.600 ;
        RECT 97.500 651.750 99.300 663.600 ;
        RECT 110.250 658.800 111.300 667.050 ;
        RECT 112.950 665.850 115.050 667.950 ;
        RECT 118.950 665.850 121.050 667.950 ;
        RECT 121.950 665.850 124.050 667.950 ;
        RECT 127.950 665.850 130.050 667.950 ;
        RECT 130.950 667.050 133.050 669.150 ;
        RECT 136.950 667.050 139.050 669.150 ;
        RECT 140.550 667.950 141.750 675.300 ;
        RECT 149.700 674.400 151.500 683.250 ;
        RECT 155.100 675.000 156.900 683.250 ;
        RECT 165.000 677.400 166.800 683.250 ;
        RECT 169.200 679.050 171.000 683.250 ;
        RECT 172.500 680.400 174.300 683.250 ;
        RECT 169.200 677.400 174.900 679.050 ;
        RECT 155.100 673.350 159.600 675.000 ;
        RECT 143.100 669.150 144.900 670.950 ;
        RECT 158.400 669.150 159.600 673.350 ;
        RECT 164.100 672.150 165.900 673.950 ;
        RECT 163.950 670.050 166.050 672.150 ;
        RECT 166.950 671.850 169.050 673.950 ;
        RECT 170.100 672.150 171.900 673.950 ;
        RECT 167.100 670.050 168.900 671.850 ;
        RECT 169.950 670.050 172.050 672.150 ;
        RECT 173.700 670.950 174.900 677.400 ;
        RECT 182.850 676.200 184.650 683.250 ;
        RECT 187.350 677.400 189.150 683.250 ;
        RECT 193.650 680.400 195.450 683.250 ;
        RECT 196.650 680.400 198.450 683.250 ;
        RECT 199.650 680.400 201.450 683.250 ;
        RECT 182.850 675.300 186.450 676.200 ;
        RECT 112.950 664.050 114.750 665.850 ;
        RECT 115.950 662.850 118.050 664.950 ;
        RECT 119.100 664.050 120.900 665.850 ;
        RECT 122.100 664.050 123.900 665.850 ;
        RECT 124.950 662.850 127.050 664.950 ;
        RECT 128.250 664.050 130.050 665.850 ;
        RECT 116.100 661.050 117.900 662.850 ;
        RECT 125.100 661.050 126.900 662.850 ;
        RECT 131.700 658.800 132.750 667.050 ;
        RECT 139.950 665.850 142.050 667.950 ;
        RECT 142.950 667.050 145.050 669.150 ;
        RECT 148.950 665.850 151.050 667.950 ;
        RECT 154.950 665.850 157.050 667.950 ;
        RECT 157.950 667.050 160.050 669.150 ;
        RECT 172.950 668.850 175.050 670.950 ;
        RECT 182.100 669.150 183.900 670.950 ;
        RECT 110.250 657.900 117.300 658.800 ;
        RECT 110.250 657.600 111.450 657.900 ;
        RECT 100.800 651.750 102.600 657.600 ;
        RECT 109.650 651.750 111.450 657.600 ;
        RECT 115.650 657.600 117.300 657.900 ;
        RECT 125.700 657.900 132.750 658.800 ;
        RECT 125.700 657.600 127.350 657.900 ;
        RECT 112.650 651.750 114.450 657.000 ;
        RECT 115.650 651.750 117.450 657.600 ;
        RECT 118.650 651.750 120.450 657.600 ;
        RECT 122.550 651.750 124.350 657.600 ;
        RECT 125.550 651.750 127.350 657.600 ;
        RECT 131.550 657.600 132.750 657.900 ;
        RECT 140.550 657.600 141.750 665.850 ;
        RECT 149.100 664.050 150.900 665.850 ;
        RECT 151.950 662.850 154.050 664.950 ;
        RECT 155.250 664.050 157.050 665.850 ;
        RECT 152.100 661.050 153.900 662.850 ;
        RECT 158.700 658.800 159.750 667.050 ;
        RECT 173.700 663.600 174.900 668.850 ;
        RECT 181.950 667.050 184.050 669.150 ;
        RECT 185.250 667.950 186.450 675.300 ;
        RECT 196.950 673.950 198.000 680.400 ;
        RECT 205.650 677.400 207.450 683.250 ;
        RECT 206.250 675.300 207.450 677.400 ;
        RECT 208.650 678.300 210.450 683.250 ;
        RECT 211.650 679.200 213.450 683.250 ;
        RECT 214.650 678.300 216.450 683.250 ;
        RECT 208.650 676.950 216.450 678.300 ;
        RECT 221.850 676.200 223.650 683.250 ;
        RECT 226.350 677.400 228.150 683.250 ;
        RECT 230.550 680.400 232.350 683.250 ;
        RECT 233.550 680.400 235.350 683.250 ;
        RECT 236.550 680.400 238.350 683.250 ;
        RECT 221.850 675.300 225.450 676.200 ;
        RECT 206.250 674.250 210.000 675.300 ;
        RECT 196.950 671.850 199.050 673.950 ;
        RECT 188.100 669.150 189.900 670.950 ;
        RECT 184.950 665.850 187.050 667.950 ;
        RECT 187.950 667.050 190.050 669.150 ;
        RECT 193.950 668.850 196.050 670.950 ;
        RECT 194.100 667.050 195.900 668.850 ;
        RECT 152.700 657.900 159.750 658.800 ;
        RECT 152.700 657.600 154.350 657.900 ;
        RECT 128.550 651.750 130.350 657.000 ;
        RECT 131.550 651.750 133.350 657.600 ;
        RECT 137.550 651.750 139.350 657.600 ;
        RECT 140.550 651.750 142.350 657.600 ;
        RECT 143.550 651.750 145.350 657.600 ;
        RECT 149.550 651.750 151.350 657.600 ;
        RECT 152.550 651.750 154.350 657.600 ;
        RECT 158.550 657.600 159.750 657.900 ;
        RECT 164.550 662.700 172.350 663.600 ;
        RECT 155.550 651.750 157.350 657.000 ;
        RECT 158.550 651.750 160.350 657.600 ;
        RECT 164.550 651.750 166.350 662.700 ;
        RECT 167.550 651.750 169.350 661.800 ;
        RECT 170.550 651.750 172.350 662.700 ;
        RECT 173.550 651.750 175.350 663.600 ;
        RECT 185.250 657.600 186.450 665.850 ;
        RECT 196.950 664.650 198.000 671.850 ;
        RECT 208.950 670.950 210.150 674.250 ;
        RECT 212.100 672.150 213.900 673.950 ;
        RECT 199.950 668.850 202.050 670.950 ;
        RECT 208.950 668.850 211.050 670.950 ;
        RECT 211.950 670.050 214.050 672.150 ;
        RECT 214.950 668.850 217.050 670.950 ;
        RECT 221.100 669.150 222.900 670.950 ;
        RECT 200.100 667.050 201.900 668.850 ;
        RECT 205.950 665.850 208.050 667.950 ;
        RECT 195.450 663.600 198.000 664.650 ;
        RECT 206.250 664.050 208.050 665.850 ;
        RECT 209.850 663.600 211.050 668.850 ;
        RECT 215.100 667.050 216.900 668.850 ;
        RECT 220.950 667.050 223.050 669.150 ;
        RECT 224.250 667.950 225.450 675.300 ;
        RECT 234.000 673.950 235.050 680.400 ;
        RECT 242.700 674.400 244.500 683.250 ;
        RECT 248.100 675.000 249.900 683.250 ;
        RECT 260.700 680.400 262.500 683.250 ;
        RECT 264.000 679.050 265.800 683.250 ;
        RECT 260.100 677.400 265.800 679.050 ;
        RECT 268.200 677.400 270.000 683.250 ;
        RECT 272.550 680.400 274.350 683.250 ;
        RECT 275.550 680.400 277.350 683.250 ;
        RECT 283.650 680.400 285.450 683.250 ;
        RECT 286.650 680.400 288.450 683.250 ;
        RECT 232.950 671.850 235.050 673.950 ;
        RECT 248.100 673.350 252.600 675.000 ;
        RECT 227.100 669.150 228.900 670.950 ;
        RECT 223.950 665.850 226.050 667.950 ;
        RECT 226.950 667.050 229.050 669.150 ;
        RECT 229.950 668.850 232.050 670.950 ;
        RECT 230.100 667.050 231.900 668.850 ;
        RECT 181.650 651.750 183.450 657.600 ;
        RECT 184.650 651.750 186.450 657.600 ;
        RECT 187.650 651.750 189.450 657.600 ;
        RECT 195.450 651.750 197.250 663.600 ;
        RECT 199.650 651.750 201.450 663.600 ;
        RECT 206.400 651.750 208.200 657.600 ;
        RECT 209.700 651.750 211.500 663.600 ;
        RECT 213.900 651.750 215.700 663.600 ;
        RECT 224.250 657.600 225.450 665.850 ;
        RECT 234.000 664.650 235.050 671.850 ;
        RECT 235.950 668.850 238.050 670.950 ;
        RECT 251.400 669.150 252.600 673.350 ;
        RECT 260.100 670.950 261.300 677.400 ;
        RECT 263.100 672.150 264.900 673.950 ;
        RECT 236.100 667.050 237.900 668.850 ;
        RECT 241.950 665.850 244.050 667.950 ;
        RECT 247.950 665.850 250.050 667.950 ;
        RECT 250.950 667.050 253.050 669.150 ;
        RECT 259.950 668.850 262.050 670.950 ;
        RECT 262.950 670.050 265.050 672.150 ;
        RECT 265.950 671.850 268.050 673.950 ;
        RECT 269.100 672.150 270.900 673.950 ;
        RECT 266.100 670.050 267.900 671.850 ;
        RECT 268.950 670.050 271.050 672.150 ;
        RECT 271.950 671.850 274.050 673.950 ;
        RECT 275.400 672.150 276.600 680.400 ;
        RECT 284.400 672.150 285.600 680.400 ;
        RECT 291.000 677.400 292.800 683.250 ;
        RECT 295.200 679.050 297.000 683.250 ;
        RECT 298.500 680.400 300.300 683.250 ;
        RECT 305.550 680.400 307.350 683.250 ;
        RECT 308.550 680.400 310.350 683.250 ;
        RECT 311.550 680.400 313.350 683.250 ;
        RECT 317.550 680.400 319.350 683.250 ;
        RECT 320.550 680.400 322.350 683.250 ;
        RECT 295.200 677.400 300.900 679.050 ;
        RECT 272.100 670.050 273.900 671.850 ;
        RECT 274.950 670.050 277.050 672.150 ;
        RECT 283.950 670.050 286.050 672.150 ;
        RECT 286.950 671.850 289.050 673.950 ;
        RECT 290.100 672.150 291.900 673.950 ;
        RECT 287.100 670.050 288.900 671.850 ;
        RECT 289.950 670.050 292.050 672.150 ;
        RECT 292.950 671.850 295.050 673.950 ;
        RECT 296.100 672.150 297.900 673.950 ;
        RECT 293.100 670.050 294.900 671.850 ;
        RECT 295.950 670.050 298.050 672.150 ;
        RECT 299.700 670.950 300.900 677.400 ;
        RECT 309.000 673.950 310.050 680.400 ;
        RECT 307.950 671.850 310.050 673.950 ;
        RECT 316.950 671.850 319.050 673.950 ;
        RECT 320.400 672.150 321.600 680.400 ;
        RECT 326.550 678.300 328.350 683.250 ;
        RECT 329.550 679.200 331.350 683.250 ;
        RECT 332.550 678.300 334.350 683.250 ;
        RECT 326.550 676.950 334.350 678.300 ;
        RECT 335.550 677.400 337.350 683.250 ;
        RECT 343.650 682.500 351.450 683.250 ;
        RECT 343.650 677.400 345.450 682.500 ;
        RECT 346.650 677.400 348.450 681.600 ;
        RECT 349.650 678.000 351.450 682.500 ;
        RECT 352.650 678.900 354.450 683.250 ;
        RECT 355.650 678.000 357.450 683.250 ;
        RECT 359.550 680.400 361.350 683.250 ;
        RECT 362.550 680.400 364.350 683.250 ;
        RECT 365.550 680.400 367.350 683.250 ;
        RECT 335.550 675.300 336.750 677.400 ;
        RECT 333.000 674.250 336.750 675.300 ;
        RECT 347.250 675.900 348.150 677.400 ;
        RECT 349.650 677.100 357.450 678.000 ;
        RECT 363.450 676.200 364.350 680.400 ;
        RECT 368.550 677.400 370.350 683.250 ;
        RECT 375.000 677.400 376.800 683.250 ;
        RECT 379.200 679.050 381.000 683.250 ;
        RECT 382.500 680.400 384.300 683.250 ;
        RECT 379.200 677.400 384.900 679.050 ;
        RECT 394.800 677.400 396.600 683.250 ;
        RECT 399.000 677.400 400.800 683.250 ;
        RECT 403.200 677.400 405.000 683.250 ;
        RECT 408.150 677.400 409.950 683.250 ;
        RECT 411.150 680.400 412.950 683.250 ;
        RECT 415.950 681.300 417.750 683.250 ;
        RECT 414.000 680.400 417.750 681.300 ;
        RECT 420.450 680.400 422.250 683.250 ;
        RECT 423.750 680.400 425.550 683.250 ;
        RECT 427.650 680.400 429.450 683.250 ;
        RECT 431.850 680.400 433.650 683.250 ;
        RECT 436.350 680.400 438.150 683.250 ;
        RECT 414.000 679.500 415.050 680.400 ;
        RECT 412.950 677.400 415.050 679.500 ;
        RECT 423.750 678.600 424.800 680.400 ;
        RECT 347.250 674.850 351.600 675.900 ;
        RECT 363.450 675.300 366.750 676.200 ;
        RECT 329.100 672.150 330.900 673.950 ;
        RECT 234.000 663.600 236.550 664.650 ;
        RECT 242.100 664.050 243.900 665.850 ;
        RECT 220.650 651.750 222.450 657.600 ;
        RECT 223.650 651.750 225.450 657.600 ;
        RECT 226.650 651.750 228.450 657.600 ;
        RECT 230.550 651.750 232.350 663.600 ;
        RECT 234.750 651.750 236.550 663.600 ;
        RECT 244.950 662.850 247.050 664.950 ;
        RECT 248.250 664.050 250.050 665.850 ;
        RECT 245.100 661.050 246.900 662.850 ;
        RECT 251.700 658.800 252.750 667.050 ;
        RECT 260.100 663.600 261.300 668.850 ;
        RECT 245.700 657.900 252.750 658.800 ;
        RECT 245.700 657.600 247.350 657.900 ;
        RECT 242.550 651.750 244.350 657.600 ;
        RECT 245.550 651.750 247.350 657.600 ;
        RECT 251.550 657.600 252.750 657.900 ;
        RECT 248.550 651.750 250.350 657.000 ;
        RECT 251.550 651.750 253.350 657.600 ;
        RECT 259.650 651.750 261.450 663.600 ;
        RECT 262.650 662.700 270.450 663.600 ;
        RECT 262.650 651.750 264.450 662.700 ;
        RECT 265.650 651.750 267.450 661.800 ;
        RECT 268.650 651.750 270.450 662.700 ;
        RECT 275.400 657.600 276.600 670.050 ;
        RECT 284.400 657.600 285.600 670.050 ;
        RECT 298.950 668.850 301.050 670.950 ;
        RECT 304.950 668.850 307.050 670.950 ;
        RECT 299.700 663.600 300.900 668.850 ;
        RECT 305.100 667.050 306.900 668.850 ;
        RECT 309.000 664.650 310.050 671.850 ;
        RECT 310.950 668.850 313.050 670.950 ;
        RECT 317.100 670.050 318.900 671.850 ;
        RECT 319.950 670.050 322.050 672.150 ;
        RECT 311.100 667.050 312.900 668.850 ;
        RECT 309.000 663.600 311.550 664.650 ;
        RECT 290.550 662.700 298.350 663.600 ;
        RECT 272.550 651.750 274.350 657.600 ;
        RECT 275.550 651.750 277.350 657.600 ;
        RECT 283.650 651.750 285.450 657.600 ;
        RECT 286.650 651.750 288.450 657.600 ;
        RECT 290.550 651.750 292.350 662.700 ;
        RECT 293.550 651.750 295.350 661.800 ;
        RECT 296.550 651.750 298.350 662.700 ;
        RECT 299.550 651.750 301.350 663.600 ;
        RECT 305.550 651.750 307.350 663.600 ;
        RECT 309.750 651.750 311.550 663.600 ;
        RECT 320.400 657.600 321.600 670.050 ;
        RECT 325.950 668.850 328.050 670.950 ;
        RECT 328.950 670.050 331.050 672.150 ;
        RECT 332.850 670.950 334.050 674.250 ;
        RECT 347.700 672.150 349.500 673.950 ;
        RECT 331.950 668.850 334.050 670.950 ;
        RECT 343.950 668.850 346.050 670.950 ;
        RECT 346.950 670.050 349.050 672.150 ;
        RECT 350.400 670.950 351.600 674.850 ;
        RECT 364.950 674.400 366.750 675.300 ;
        RECT 353.100 672.150 354.900 673.950 ;
        RECT 349.950 668.850 352.050 670.950 ;
        RECT 352.950 670.050 355.050 672.150 ;
        RECT 358.950 671.850 361.050 673.950 ;
        RECT 355.950 668.850 358.050 670.950 ;
        RECT 359.100 670.050 360.900 671.850 ;
        RECT 361.950 668.850 364.050 670.950 ;
        RECT 326.100 667.050 327.900 668.850 ;
        RECT 331.950 663.600 333.150 668.850 ;
        RECT 334.950 665.850 337.050 667.950 ;
        RECT 344.250 667.050 346.050 668.850 ;
        RECT 334.950 664.050 336.750 665.850 ;
        RECT 350.250 663.600 351.450 668.850 ;
        RECT 356.100 667.050 357.900 668.850 ;
        RECT 362.100 667.050 363.900 668.850 ;
        RECT 365.700 666.150 366.600 674.400 ;
        RECT 369.000 672.150 370.050 677.400 ;
        RECT 374.100 672.150 375.900 673.950 ;
        RECT 367.950 670.050 370.050 672.150 ;
        RECT 373.950 670.050 376.050 672.150 ;
        RECT 376.950 671.850 379.050 673.950 ;
        RECT 380.100 672.150 381.900 673.950 ;
        RECT 377.100 670.050 378.900 671.850 ;
        RECT 379.950 670.050 382.050 672.150 ;
        RECT 383.700 670.950 384.900 677.400 ;
        RECT 395.250 672.150 397.050 673.950 ;
        RECT 364.950 666.000 366.750 666.150 ;
        RECT 359.550 664.800 366.750 666.000 ;
        RECT 359.550 663.600 360.750 664.800 ;
        RECT 364.950 664.350 366.750 664.800 ;
        RECT 317.550 651.750 319.350 657.600 ;
        RECT 320.550 651.750 322.350 657.600 ;
        RECT 327.300 651.750 329.100 663.600 ;
        RECT 331.500 651.750 333.300 663.600 ;
        RECT 334.800 651.750 336.600 657.600 ;
        RECT 345.150 651.750 346.950 663.600 ;
        RECT 349.650 651.750 352.950 663.600 ;
        RECT 355.650 651.750 357.450 663.600 ;
        RECT 359.550 651.750 361.350 663.600 ;
        RECT 368.100 663.450 369.450 670.050 ;
        RECT 382.950 668.850 385.050 670.950 ;
        RECT 391.950 668.850 394.050 670.950 ;
        RECT 394.950 670.050 397.050 672.150 ;
        RECT 399.000 670.950 400.050 677.400 ;
        RECT 397.950 668.850 400.050 670.950 ;
        RECT 400.950 672.150 402.750 673.950 ;
        RECT 400.950 670.050 403.050 672.150 ;
        RECT 403.950 668.850 406.050 670.950 ;
        RECT 383.700 663.600 384.900 668.850 ;
        RECT 392.100 667.050 393.900 668.850 ;
        RECT 397.950 665.400 398.850 668.850 ;
        RECT 403.950 667.050 405.750 668.850 ;
        RECT 394.800 664.500 398.850 665.400 ;
        RECT 408.150 664.800 409.050 677.400 ;
        RECT 416.550 676.800 418.350 678.600 ;
        RECT 419.850 677.550 424.800 678.600 ;
        RECT 432.300 679.500 433.350 680.400 ;
        RECT 432.300 678.300 436.050 679.500 ;
        RECT 419.850 676.800 421.650 677.550 ;
        RECT 416.850 675.900 417.900 676.800 ;
        RECT 427.050 676.200 428.850 678.000 ;
        RECT 433.950 677.400 436.050 678.300 ;
        RECT 439.650 677.400 441.450 683.250 ;
        RECT 445.650 680.400 447.450 683.250 ;
        RECT 448.650 680.400 450.450 683.250 ;
        RECT 427.050 675.900 427.950 676.200 ;
        RECT 416.850 675.000 427.950 675.900 ;
        RECT 440.250 675.150 441.450 677.400 ;
        RECT 416.850 673.800 417.900 675.000 ;
        RECT 411.000 672.600 417.900 673.800 ;
        RECT 411.000 671.850 411.900 672.600 ;
        RECT 416.100 672.000 417.900 672.600 ;
        RECT 410.100 670.050 411.900 671.850 ;
        RECT 413.100 670.950 414.900 671.700 ;
        RECT 427.050 670.950 427.950 675.000 ;
        RECT 436.950 673.050 441.450 675.150 ;
        RECT 435.150 671.250 439.050 673.050 ;
        RECT 436.950 670.950 439.050 671.250 ;
        RECT 413.100 669.900 421.050 670.950 ;
        RECT 418.950 668.850 421.050 669.900 ;
        RECT 424.950 668.850 427.950 670.950 ;
        RECT 417.450 665.100 419.250 665.400 ;
        RECT 417.450 664.800 425.850 665.100 ;
        RECT 394.800 663.600 396.600 664.500 ;
        RECT 408.150 664.200 425.850 664.800 ;
        RECT 408.150 663.600 419.250 664.200 ;
        RECT 364.050 651.750 365.850 663.450 ;
        RECT 367.050 662.100 369.450 663.450 ;
        RECT 374.550 662.700 382.350 663.600 ;
        RECT 367.050 651.750 368.850 662.100 ;
        RECT 374.550 651.750 376.350 662.700 ;
        RECT 377.550 651.750 379.350 661.800 ;
        RECT 380.550 651.750 382.350 662.700 ;
        RECT 383.550 651.750 385.350 663.600 ;
        RECT 391.650 652.500 393.450 663.600 ;
        RECT 394.650 653.400 396.450 663.600 ;
        RECT 397.650 662.400 405.450 663.300 ;
        RECT 397.650 652.500 399.450 662.400 ;
        RECT 391.650 651.750 399.450 652.500 ;
        RECT 400.650 651.750 402.450 661.500 ;
        RECT 403.650 651.750 405.450 662.400 ;
        RECT 408.150 651.750 409.950 663.600 ;
        RECT 422.250 662.700 424.050 663.300 ;
        RECT 416.550 661.500 424.050 662.700 ;
        RECT 424.950 662.100 425.850 664.200 ;
        RECT 427.050 664.200 427.950 668.850 ;
        RECT 437.250 665.400 439.050 667.200 ;
        RECT 433.950 664.200 438.150 665.400 ;
        RECT 427.050 663.300 433.050 664.200 ;
        RECT 433.950 663.300 436.050 664.200 ;
        RECT 440.250 663.600 441.450 673.050 ;
        RECT 446.400 672.150 447.600 680.400 ;
        RECT 454.650 677.400 456.450 683.250 ;
        RECT 455.250 675.300 456.450 677.400 ;
        RECT 457.650 678.300 459.450 683.250 ;
        RECT 460.650 679.200 462.450 683.250 ;
        RECT 463.650 678.300 465.450 683.250 ;
        RECT 469.650 680.400 471.450 683.250 ;
        RECT 472.650 680.400 474.450 683.250 ;
        RECT 475.650 680.400 477.450 683.250 ;
        RECT 469.950 678.450 472.050 679.050 ;
        RECT 457.650 676.950 465.450 678.300 ;
        RECT 467.550 677.550 472.050 678.450 ;
        RECT 455.250 674.250 459.000 675.300 ;
        RECT 445.950 670.050 448.050 672.150 ;
        RECT 448.950 671.850 451.050 673.950 ;
        RECT 449.100 670.050 450.900 671.850 ;
        RECT 457.950 670.950 459.150 674.250 ;
        RECT 461.100 672.150 462.900 673.950 ;
        RECT 432.150 662.400 433.050 663.300 ;
        RECT 429.450 662.100 431.250 662.400 ;
        RECT 416.550 660.600 417.750 661.500 ;
        RECT 424.950 661.200 431.250 662.100 ;
        RECT 429.450 660.600 431.250 661.200 ;
        RECT 432.150 660.600 434.850 662.400 ;
        RECT 412.950 658.500 417.750 660.600 ;
        RECT 420.150 658.500 427.050 660.300 ;
        RECT 416.550 657.600 417.750 658.500 ;
        RECT 411.150 651.750 412.950 657.600 ;
        RECT 416.250 651.750 418.050 657.600 ;
        RECT 421.050 651.750 422.850 657.600 ;
        RECT 424.050 651.750 425.850 658.500 ;
        RECT 432.150 657.600 436.050 659.700 ;
        RECT 427.950 651.750 429.750 657.600 ;
        RECT 432.150 651.750 433.950 657.600 ;
        RECT 436.650 651.750 438.450 654.600 ;
        RECT 439.650 651.750 441.450 663.600 ;
        RECT 446.400 657.600 447.600 670.050 ;
        RECT 457.950 668.850 460.050 670.950 ;
        RECT 460.950 670.050 463.050 672.150 ;
        RECT 463.950 668.850 466.050 670.950 ;
        RECT 454.950 665.850 457.050 667.950 ;
        RECT 455.250 664.050 457.050 665.850 ;
        RECT 458.850 663.600 460.050 668.850 ;
        RECT 464.100 667.050 465.900 668.850 ;
        RECT 467.550 667.050 468.450 677.550 ;
        RECT 469.950 676.950 472.050 677.550 ;
        RECT 472.950 673.950 474.000 680.400 ;
        RECT 481.650 677.400 483.450 683.250 ;
        RECT 482.250 675.300 483.450 677.400 ;
        RECT 484.650 678.300 486.450 683.250 ;
        RECT 487.650 679.200 489.450 683.250 ;
        RECT 490.650 678.300 492.450 683.250 ;
        RECT 496.650 680.400 498.450 683.250 ;
        RECT 499.650 680.400 501.450 683.250 ;
        RECT 502.650 680.400 504.450 683.250 ;
        RECT 508.650 680.400 510.450 683.250 ;
        RECT 511.650 680.400 513.450 683.250 ;
        RECT 484.650 676.950 492.450 678.300 ;
        RECT 482.250 674.250 486.000 675.300 ;
        RECT 472.950 671.850 475.050 673.950 ;
        RECT 469.950 668.850 472.050 670.950 ;
        RECT 470.100 667.050 471.900 668.850 ;
        RECT 466.950 664.950 469.050 667.050 ;
        RECT 472.950 664.650 474.000 671.850 ;
        RECT 484.950 670.950 486.150 674.250 ;
        RECT 499.950 673.950 501.000 680.400 ;
        RECT 488.100 672.150 489.900 673.950 ;
        RECT 475.950 668.850 478.050 670.950 ;
        RECT 484.950 668.850 487.050 670.950 ;
        RECT 487.950 670.050 490.050 672.150 ;
        RECT 499.950 671.850 502.050 673.950 ;
        RECT 509.400 672.150 510.600 680.400 ;
        RECT 515.550 677.400 517.350 683.250 ;
        RECT 518.850 680.400 520.650 683.250 ;
        RECT 523.350 680.400 525.150 683.250 ;
        RECT 527.550 680.400 529.350 683.250 ;
        RECT 531.450 680.400 533.250 683.250 ;
        RECT 534.750 680.400 536.550 683.250 ;
        RECT 539.250 681.300 541.050 683.250 ;
        RECT 539.250 680.400 543.000 681.300 ;
        RECT 544.050 680.400 545.850 683.250 ;
        RECT 523.650 679.500 524.700 680.400 ;
        RECT 520.950 678.300 524.700 679.500 ;
        RECT 532.200 678.600 533.250 680.400 ;
        RECT 541.950 679.500 543.000 680.400 ;
        RECT 520.950 677.400 523.050 678.300 ;
        RECT 515.550 675.150 516.750 677.400 ;
        RECT 528.150 676.200 529.950 678.000 ;
        RECT 532.200 677.550 537.150 678.600 ;
        RECT 535.350 676.800 537.150 677.550 ;
        RECT 538.650 676.800 540.450 678.600 ;
        RECT 541.950 677.400 544.050 679.500 ;
        RECT 547.050 677.400 548.850 683.250 ;
        RECT 529.050 675.900 529.950 676.200 ;
        RECT 539.100 675.900 540.150 676.800 ;
        RECT 490.950 668.850 493.050 670.950 ;
        RECT 496.950 668.850 499.050 670.950 ;
        RECT 476.100 667.050 477.900 668.850 ;
        RECT 481.950 665.850 484.050 667.950 ;
        RECT 471.450 663.600 474.000 664.650 ;
        RECT 482.250 664.050 484.050 665.850 ;
        RECT 485.850 663.600 487.050 668.850 ;
        RECT 491.100 667.050 492.900 668.850 ;
        RECT 497.100 667.050 498.900 668.850 ;
        RECT 499.950 664.650 501.000 671.850 ;
        RECT 502.950 668.850 505.050 670.950 ;
        RECT 508.950 670.050 511.050 672.150 ;
        RECT 511.950 671.850 514.050 673.950 ;
        RECT 515.550 673.050 520.050 675.150 ;
        RECT 529.050 675.000 540.150 675.900 ;
        RECT 512.100 670.050 513.900 671.850 ;
        RECT 503.100 667.050 504.900 668.850 ;
        RECT 498.450 663.600 501.000 664.650 ;
        RECT 445.650 651.750 447.450 657.600 ;
        RECT 448.650 651.750 450.450 657.600 ;
        RECT 455.400 651.750 457.200 657.600 ;
        RECT 458.700 651.750 460.500 663.600 ;
        RECT 462.900 651.750 464.700 663.600 ;
        RECT 471.450 651.750 473.250 663.600 ;
        RECT 475.650 651.750 477.450 663.600 ;
        RECT 482.400 651.750 484.200 657.600 ;
        RECT 485.700 651.750 487.500 663.600 ;
        RECT 489.900 651.750 491.700 663.600 ;
        RECT 498.450 651.750 500.250 663.600 ;
        RECT 502.650 651.750 504.450 663.600 ;
        RECT 509.400 657.600 510.600 670.050 ;
        RECT 515.550 663.600 516.750 673.050 ;
        RECT 517.950 671.250 521.850 673.050 ;
        RECT 517.950 670.950 520.050 671.250 ;
        RECT 529.050 670.950 529.950 675.000 ;
        RECT 539.100 673.800 540.150 675.000 ;
        RECT 539.100 672.600 546.000 673.800 ;
        RECT 539.100 672.000 540.900 672.600 ;
        RECT 545.100 671.850 546.000 672.600 ;
        RECT 542.100 670.950 543.900 671.700 ;
        RECT 529.050 668.850 532.050 670.950 ;
        RECT 535.950 669.900 543.900 670.950 ;
        RECT 545.100 670.050 546.900 671.850 ;
        RECT 535.950 668.850 538.050 669.900 ;
        RECT 517.950 665.400 519.750 667.200 ;
        RECT 518.850 664.200 523.050 665.400 ;
        RECT 529.050 664.200 529.950 668.850 ;
        RECT 537.750 665.100 539.550 665.400 ;
        RECT 508.650 651.750 510.450 657.600 ;
        RECT 511.650 651.750 513.450 657.600 ;
        RECT 515.550 651.750 517.350 663.600 ;
        RECT 520.950 663.300 523.050 664.200 ;
        RECT 523.950 663.300 529.950 664.200 ;
        RECT 531.150 664.800 539.550 665.100 ;
        RECT 547.950 664.800 548.850 677.400 ;
        RECT 551.550 678.300 553.350 683.250 ;
        RECT 554.550 679.200 556.350 683.250 ;
        RECT 557.550 678.300 559.350 683.250 ;
        RECT 551.550 676.950 559.350 678.300 ;
        RECT 560.550 677.400 562.350 683.250 ;
        RECT 566.850 677.400 568.650 683.250 ;
        RECT 560.550 675.300 561.750 677.400 ;
        RECT 571.350 676.200 573.150 683.250 ;
        RECT 580.650 677.400 582.450 683.250 ;
        RECT 583.650 677.400 585.450 683.250 ;
        RECT 586.650 677.400 588.450 683.250 ;
        RECT 589.650 677.400 591.450 683.250 ;
        RECT 592.650 677.400 594.450 683.250 ;
        RECT 583.800 676.500 585.600 677.400 ;
        RECT 589.800 676.500 591.600 677.400 ;
        RECT 595.650 676.500 597.450 683.250 ;
        RECT 598.650 677.400 600.450 683.250 ;
        RECT 601.650 677.400 603.450 683.250 ;
        RECT 604.650 677.400 606.450 683.250 ;
        RECT 610.350 677.400 612.150 683.250 ;
        RECT 613.350 677.400 615.150 683.250 ;
        RECT 616.650 680.400 618.450 683.250 ;
        RECT 601.800 676.500 603.600 677.400 ;
        RECT 582.900 676.350 585.600 676.500 ;
        RECT 558.000 674.250 561.750 675.300 ;
        RECT 569.550 675.300 573.150 676.200 ;
        RECT 582.750 675.300 585.600 676.350 ;
        RECT 587.700 675.300 591.600 676.500 ;
        RECT 593.700 675.300 597.450 676.500 ;
        RECT 599.550 675.300 603.600 676.500 ;
        RECT 554.100 672.150 555.900 673.950 ;
        RECT 550.950 668.850 553.050 670.950 ;
        RECT 553.950 670.050 556.050 672.150 ;
        RECT 557.850 670.950 559.050 674.250 ;
        RECT 556.950 668.850 559.050 670.950 ;
        RECT 566.100 669.150 567.900 670.950 ;
        RECT 551.100 667.050 552.900 668.850 ;
        RECT 531.150 664.200 548.850 664.800 ;
        RECT 523.950 662.400 524.850 663.300 ;
        RECT 522.150 660.600 524.850 662.400 ;
        RECT 525.750 662.100 527.550 662.400 ;
        RECT 531.150 662.100 532.050 664.200 ;
        RECT 537.750 663.600 548.850 664.200 ;
        RECT 556.950 663.600 558.150 668.850 ;
        RECT 559.950 665.850 562.050 667.950 ;
        RECT 565.950 667.050 568.050 669.150 ;
        RECT 569.550 667.950 570.750 675.300 ;
        RECT 582.750 672.150 583.800 675.300 ;
        RECT 587.700 674.400 588.900 675.300 ;
        RECT 593.700 674.400 594.900 675.300 ;
        RECT 599.550 674.400 600.750 675.300 ;
        RECT 584.700 672.600 588.900 674.400 ;
        RECT 590.700 672.600 594.900 674.400 ;
        RECT 596.700 672.600 600.750 674.400 ;
        RECT 572.100 669.150 573.900 670.950 ;
        RECT 580.950 670.050 583.800 672.150 ;
        RECT 568.950 665.850 571.050 667.950 ;
        RECT 571.950 667.050 574.050 669.150 ;
        RECT 559.950 664.050 561.750 665.850 ;
        RECT 525.750 661.200 532.050 662.100 ;
        RECT 532.950 662.700 534.750 663.300 ;
        RECT 532.950 661.500 540.450 662.700 ;
        RECT 525.750 660.600 527.550 661.200 ;
        RECT 539.250 660.600 540.450 661.500 ;
        RECT 520.950 657.600 524.850 659.700 ;
        RECT 529.950 658.500 536.850 660.300 ;
        RECT 539.250 658.500 544.050 660.600 ;
        RECT 518.550 651.750 520.350 654.600 ;
        RECT 523.050 651.750 524.850 657.600 ;
        RECT 527.250 651.750 529.050 657.600 ;
        RECT 531.150 651.750 532.950 658.500 ;
        RECT 539.250 657.600 540.450 658.500 ;
        RECT 534.150 651.750 535.950 657.600 ;
        RECT 538.950 651.750 540.750 657.600 ;
        RECT 544.050 651.750 545.850 657.600 ;
        RECT 547.050 651.750 548.850 663.600 ;
        RECT 552.300 651.750 554.100 663.600 ;
        RECT 556.500 651.750 558.300 663.600 ;
        RECT 569.550 657.600 570.750 665.850 ;
        RECT 582.750 665.700 583.800 670.050 ;
        RECT 587.700 665.700 588.900 672.600 ;
        RECT 593.700 665.700 594.900 672.600 ;
        RECT 599.550 665.700 600.750 672.600 ;
        RECT 602.100 672.150 603.900 673.950 ;
        RECT 601.950 670.050 604.050 672.150 ;
        RECT 610.650 670.950 611.850 677.400 ;
        RECT 616.650 676.500 617.850 680.400 ;
        RECT 620.850 677.400 622.650 683.250 ;
        RECT 612.750 675.600 617.850 676.500 ;
        RECT 625.350 676.200 627.150 683.250 ;
        RECT 632.550 680.400 634.350 683.250 ;
        RECT 635.550 680.400 637.350 683.250 ;
        RECT 612.750 674.700 615.000 675.600 ;
        RECT 610.650 668.850 613.050 670.950 ;
        RECT 582.750 664.500 585.450 665.700 ;
        RECT 587.700 664.500 591.450 665.700 ;
        RECT 593.700 664.500 597.450 665.700 ;
        RECT 599.550 664.500 603.450 665.700 ;
        RECT 559.800 651.750 561.600 657.600 ;
        RECT 566.550 651.750 568.350 657.600 ;
        RECT 569.550 651.750 571.350 657.600 ;
        RECT 572.550 651.750 574.350 657.600 ;
        RECT 580.650 651.750 582.450 663.600 ;
        RECT 583.650 651.750 585.450 664.500 ;
        RECT 586.650 651.750 588.450 663.600 ;
        RECT 589.650 651.750 591.450 664.500 ;
        RECT 592.650 651.750 594.450 663.600 ;
        RECT 595.650 651.750 597.450 664.500 ;
        RECT 598.650 651.750 600.450 663.600 ;
        RECT 601.650 651.750 603.450 664.500 ;
        RECT 610.650 663.600 611.850 668.850 ;
        RECT 613.950 666.300 615.000 674.700 ;
        RECT 623.550 675.300 627.150 676.200 ;
        RECT 616.950 668.850 619.050 670.950 ;
        RECT 620.100 669.150 621.900 670.950 ;
        RECT 617.100 667.050 618.900 668.850 ;
        RECT 619.950 667.050 622.050 669.150 ;
        RECT 623.550 667.950 624.750 675.300 ;
        RECT 631.950 671.850 634.050 673.950 ;
        RECT 635.400 672.150 636.600 680.400 ;
        RECT 641.550 678.300 643.350 683.250 ;
        RECT 644.550 679.200 646.350 683.250 ;
        RECT 647.550 678.300 649.350 683.250 ;
        RECT 641.550 676.950 649.350 678.300 ;
        RECT 650.550 677.400 652.350 683.250 ;
        RECT 656.550 677.400 658.350 683.250 ;
        RECT 659.850 680.400 661.650 683.250 ;
        RECT 664.350 680.400 666.150 683.250 ;
        RECT 668.550 680.400 670.350 683.250 ;
        RECT 672.450 680.400 674.250 683.250 ;
        RECT 675.750 680.400 677.550 683.250 ;
        RECT 680.250 681.300 682.050 683.250 ;
        RECT 680.250 680.400 684.000 681.300 ;
        RECT 685.050 680.400 686.850 683.250 ;
        RECT 664.650 679.500 665.700 680.400 ;
        RECT 661.950 678.300 665.700 679.500 ;
        RECT 673.200 678.600 674.250 680.400 ;
        RECT 682.950 679.500 684.000 680.400 ;
        RECT 661.950 677.400 664.050 678.300 ;
        RECT 650.550 675.300 651.750 677.400 ;
        RECT 648.000 674.250 651.750 675.300 ;
        RECT 656.550 675.150 657.750 677.400 ;
        RECT 669.150 676.200 670.950 678.000 ;
        RECT 673.200 677.550 678.150 678.600 ;
        RECT 676.350 676.800 678.150 677.550 ;
        RECT 679.650 676.800 681.450 678.600 ;
        RECT 682.950 677.400 685.050 679.500 ;
        RECT 688.050 677.400 689.850 683.250 ;
        RECT 692.550 680.400 694.350 683.250 ;
        RECT 670.050 675.900 670.950 676.200 ;
        RECT 680.100 675.900 681.150 676.800 ;
        RECT 644.100 672.150 645.900 673.950 ;
        RECT 626.100 669.150 627.900 670.950 ;
        RECT 632.100 670.050 633.900 671.850 ;
        RECT 634.950 670.050 637.050 672.150 ;
        RECT 612.750 665.400 615.000 666.300 ;
        RECT 622.950 665.850 625.050 667.950 ;
        RECT 625.950 667.050 628.050 669.150 ;
        RECT 612.750 664.500 618.450 665.400 ;
        RECT 604.650 651.750 606.450 663.600 ;
        RECT 610.350 651.750 612.150 663.600 ;
        RECT 613.350 651.750 615.150 663.600 ;
        RECT 617.250 657.600 618.450 664.500 ;
        RECT 623.550 657.600 624.750 665.850 ;
        RECT 635.400 657.600 636.600 670.050 ;
        RECT 640.950 668.850 643.050 670.950 ;
        RECT 643.950 670.050 646.050 672.150 ;
        RECT 647.850 670.950 649.050 674.250 ;
        RECT 646.950 668.850 649.050 670.950 ;
        RECT 656.550 673.050 661.050 675.150 ;
        RECT 670.050 675.000 681.150 675.900 ;
        RECT 641.100 667.050 642.900 668.850 ;
        RECT 646.950 663.600 648.150 668.850 ;
        RECT 649.950 665.850 652.050 667.950 ;
        RECT 649.950 664.050 651.750 665.850 ;
        RECT 656.550 663.600 657.750 673.050 ;
        RECT 658.950 671.250 662.850 673.050 ;
        RECT 658.950 670.950 661.050 671.250 ;
        RECT 670.050 670.950 670.950 675.000 ;
        RECT 680.100 673.800 681.150 675.000 ;
        RECT 680.100 672.600 687.000 673.800 ;
        RECT 680.100 672.000 681.900 672.600 ;
        RECT 686.100 671.850 687.000 672.600 ;
        RECT 683.100 670.950 684.900 671.700 ;
        RECT 670.050 668.850 673.050 670.950 ;
        RECT 676.950 669.900 684.900 670.950 ;
        RECT 686.100 670.050 687.900 671.850 ;
        RECT 676.950 668.850 679.050 669.900 ;
        RECT 658.950 665.400 660.750 667.200 ;
        RECT 659.850 664.200 664.050 665.400 ;
        RECT 670.050 664.200 670.950 668.850 ;
        RECT 678.750 665.100 680.550 665.400 ;
        RECT 616.650 651.750 618.450 657.600 ;
        RECT 620.550 651.750 622.350 657.600 ;
        RECT 623.550 651.750 625.350 657.600 ;
        RECT 626.550 651.750 628.350 657.600 ;
        RECT 632.550 651.750 634.350 657.600 ;
        RECT 635.550 651.750 637.350 657.600 ;
        RECT 642.300 651.750 644.100 663.600 ;
        RECT 646.500 651.750 648.300 663.600 ;
        RECT 649.800 651.750 651.600 657.600 ;
        RECT 656.550 651.750 658.350 663.600 ;
        RECT 661.950 663.300 664.050 664.200 ;
        RECT 664.950 663.300 670.950 664.200 ;
        RECT 672.150 664.800 680.550 665.100 ;
        RECT 688.950 664.800 689.850 677.400 ;
        RECT 693.150 676.500 694.350 680.400 ;
        RECT 695.850 677.400 697.650 683.250 ;
        RECT 698.850 677.400 700.650 683.250 ;
        RECT 704.850 677.400 706.650 683.250 ;
        RECT 693.150 675.600 698.250 676.500 ;
        RECT 696.000 674.700 698.250 675.600 ;
        RECT 691.950 668.850 694.050 670.950 ;
        RECT 692.100 667.050 693.900 668.850 ;
        RECT 696.000 666.300 697.050 674.700 ;
        RECT 699.150 670.950 700.350 677.400 ;
        RECT 709.350 676.200 711.150 683.250 ;
        RECT 707.550 675.300 711.150 676.200 ;
        RECT 697.950 668.850 700.350 670.950 ;
        RECT 704.100 669.150 705.900 670.950 ;
        RECT 696.000 665.400 698.250 666.300 ;
        RECT 672.150 664.200 689.850 664.800 ;
        RECT 664.950 662.400 665.850 663.300 ;
        RECT 663.150 660.600 665.850 662.400 ;
        RECT 666.750 662.100 668.550 662.400 ;
        RECT 672.150 662.100 673.050 664.200 ;
        RECT 678.750 663.600 689.850 664.200 ;
        RECT 666.750 661.200 673.050 662.100 ;
        RECT 673.950 662.700 675.750 663.300 ;
        RECT 673.950 661.500 681.450 662.700 ;
        RECT 666.750 660.600 668.550 661.200 ;
        RECT 680.250 660.600 681.450 661.500 ;
        RECT 661.950 657.600 665.850 659.700 ;
        RECT 670.950 658.500 677.850 660.300 ;
        RECT 680.250 658.500 685.050 660.600 ;
        RECT 659.550 651.750 661.350 654.600 ;
        RECT 664.050 651.750 665.850 657.600 ;
        RECT 668.250 651.750 670.050 657.600 ;
        RECT 672.150 651.750 673.950 658.500 ;
        RECT 680.250 657.600 681.450 658.500 ;
        RECT 675.150 651.750 676.950 657.600 ;
        RECT 679.950 651.750 681.750 657.600 ;
        RECT 685.050 651.750 686.850 657.600 ;
        RECT 688.050 651.750 689.850 663.600 ;
        RECT 692.550 664.500 698.250 665.400 ;
        RECT 692.550 657.600 693.750 664.500 ;
        RECT 699.150 663.600 700.350 668.850 ;
        RECT 703.950 667.050 706.050 669.150 ;
        RECT 707.550 667.950 708.750 675.300 ;
        RECT 710.100 669.150 711.900 670.950 ;
        RECT 706.950 665.850 709.050 667.950 ;
        RECT 709.950 667.050 712.050 669.150 ;
        RECT 692.550 651.750 694.350 657.600 ;
        RECT 695.850 651.750 697.650 663.600 ;
        RECT 698.850 651.750 700.650 663.600 ;
        RECT 707.550 657.600 708.750 665.850 ;
        RECT 704.550 651.750 706.350 657.600 ;
        RECT 707.550 651.750 709.350 657.600 ;
        RECT 710.550 651.750 712.350 657.600 ;
        RECT 4.650 641.400 6.450 647.250 ;
        RECT 7.650 641.400 9.450 647.250 ;
        RECT 10.650 641.400 12.450 647.250 ;
        RECT 8.250 633.150 9.450 641.400 ;
        RECT 14.550 636.300 16.350 647.250 ;
        RECT 17.550 637.200 19.350 647.250 ;
        RECT 20.550 636.300 22.350 647.250 ;
        RECT 14.550 635.400 22.350 636.300 ;
        RECT 23.550 635.400 25.350 647.250 ;
        RECT 31.650 641.400 33.450 647.250 ;
        RECT 34.650 641.400 36.450 647.250 ;
        RECT 37.650 641.400 39.450 647.250 ;
        RECT 4.950 629.850 7.050 631.950 ;
        RECT 7.950 631.050 10.050 633.150 ;
        RECT 5.100 628.050 6.900 629.850 ;
        RECT 8.250 623.700 9.450 631.050 ;
        RECT 10.950 629.850 13.050 631.950 ;
        RECT 23.700 630.150 24.900 635.400 ;
        RECT 35.250 633.150 36.450 641.400 ;
        RECT 45.450 635.400 47.250 647.250 ;
        RECT 49.650 635.400 51.450 647.250 ;
        RECT 56.400 641.400 58.200 647.250 ;
        RECT 59.700 635.400 61.500 647.250 ;
        RECT 63.900 635.400 65.700 647.250 ;
        RECT 69.300 635.400 71.100 647.250 ;
        RECT 73.500 635.400 75.300 647.250 ;
        RECT 76.800 641.400 78.600 647.250 ;
        RECT 85.650 641.400 87.450 647.250 ;
        RECT 88.650 641.400 90.450 647.250 ;
        RECT 45.450 634.350 48.000 635.400 ;
        RECT 11.100 628.050 12.900 629.850 ;
        RECT 13.950 626.850 16.050 628.950 ;
        RECT 17.100 627.150 18.900 628.950 ;
        RECT 14.100 625.050 15.900 626.850 ;
        RECT 16.950 625.050 19.050 627.150 ;
        RECT 19.950 626.850 22.050 628.950 ;
        RECT 22.950 628.050 25.050 630.150 ;
        RECT 31.950 629.850 34.050 631.950 ;
        RECT 34.950 631.050 37.050 633.150 ;
        RECT 32.100 628.050 33.900 629.850 ;
        RECT 20.100 625.050 21.900 626.850 ;
        RECT 5.850 622.800 9.450 623.700 ;
        RECT 5.850 615.750 7.650 622.800 ;
        RECT 23.700 621.600 24.900 628.050 ;
        RECT 35.250 623.700 36.450 631.050 ;
        RECT 37.950 629.850 40.050 631.950 ;
        RECT 44.100 630.150 45.900 631.950 ;
        RECT 38.100 628.050 39.900 629.850 ;
        RECT 43.950 628.050 46.050 630.150 ;
        RECT 10.350 615.750 12.150 621.600 ;
        RECT 15.000 615.750 16.800 621.600 ;
        RECT 19.200 619.950 24.900 621.600 ;
        RECT 32.850 622.800 36.450 623.700 ;
        RECT 46.950 627.150 48.000 634.350 ;
        RECT 56.250 633.150 58.050 634.950 ;
        RECT 50.100 630.150 51.900 631.950 ;
        RECT 55.950 631.050 58.050 633.150 ;
        RECT 59.850 630.150 61.050 635.400 ;
        RECT 65.100 630.150 66.900 631.950 ;
        RECT 68.100 630.150 69.900 631.950 ;
        RECT 73.950 630.150 75.150 635.400 ;
        RECT 76.950 633.150 78.750 634.950 ;
        RECT 76.950 631.050 79.050 633.150 ;
        RECT 49.950 628.050 52.050 630.150 ;
        RECT 58.950 628.050 61.050 630.150 ;
        RECT 46.950 625.050 49.050 627.150 ;
        RECT 19.200 615.750 21.000 619.950 ;
        RECT 22.500 615.750 24.300 618.600 ;
        RECT 32.850 615.750 34.650 622.800 ;
        RECT 37.350 615.750 39.150 621.600 ;
        RECT 46.950 618.600 48.000 625.050 ;
        RECT 58.950 624.750 60.150 628.050 ;
        RECT 61.950 626.850 64.050 628.950 ;
        RECT 64.950 628.050 67.050 630.150 ;
        RECT 67.950 628.050 70.050 630.150 ;
        RECT 70.950 626.850 73.050 628.950 ;
        RECT 73.950 628.050 76.050 630.150 ;
        RECT 86.400 628.950 87.600 641.400 ;
        RECT 94.650 635.400 96.450 647.250 ;
        RECT 97.650 636.300 99.450 647.250 ;
        RECT 100.650 637.200 102.450 647.250 ;
        RECT 103.650 636.300 105.450 647.250 ;
        RECT 109.650 641.400 111.450 647.250 ;
        RECT 112.650 641.400 114.450 647.250 ;
        RECT 116.550 641.400 118.350 647.250 ;
        RECT 119.550 641.400 121.350 647.250 ;
        RECT 122.550 642.000 124.350 647.250 ;
        RECT 97.650 635.400 105.450 636.300 ;
        RECT 95.100 630.150 96.300 635.400 ;
        RECT 62.100 625.050 63.900 626.850 ;
        RECT 71.100 625.050 72.900 626.850 ;
        RECT 74.850 624.750 76.050 628.050 ;
        RECT 85.950 626.850 88.050 628.950 ;
        RECT 89.100 627.150 90.900 628.950 ;
        RECT 94.950 628.050 97.050 630.150 ;
        RECT 110.400 628.950 111.600 641.400 ;
        RECT 119.700 641.100 121.350 641.400 ;
        RECT 125.550 641.400 127.350 647.250 ;
        RECT 133.650 646.500 141.450 647.250 ;
        RECT 125.550 641.100 126.750 641.400 ;
        RECT 119.700 640.200 126.750 641.100 ;
        RECT 119.100 636.150 120.900 637.950 ;
        RECT 116.100 633.150 117.900 634.950 ;
        RECT 118.950 634.050 121.050 636.150 ;
        RECT 122.250 633.150 124.050 634.950 ;
        RECT 115.950 631.050 118.050 633.150 ;
        RECT 121.950 631.050 124.050 633.150 ;
        RECT 125.700 631.950 126.750 640.200 ;
        RECT 133.650 635.400 135.450 646.500 ;
        RECT 136.650 635.400 138.450 645.600 ;
        RECT 139.650 636.600 141.450 646.500 ;
        RECT 142.650 637.500 144.450 647.250 ;
        RECT 145.650 636.600 147.450 647.250 ;
        RECT 151.650 641.400 153.450 647.250 ;
        RECT 154.650 642.000 156.450 647.250 ;
        RECT 139.650 635.700 147.450 636.600 ;
        RECT 152.250 641.100 153.450 641.400 ;
        RECT 157.650 641.400 159.450 647.250 ;
        RECT 160.650 641.400 162.450 647.250 ;
        RECT 164.550 641.400 166.350 647.250 ;
        RECT 167.550 641.400 169.350 647.250 ;
        RECT 170.550 642.000 172.350 647.250 ;
        RECT 157.650 641.100 159.300 641.400 ;
        RECT 152.250 640.200 159.300 641.100 ;
        RECT 167.700 641.100 169.350 641.400 ;
        RECT 173.550 641.400 175.350 647.250 ;
        RECT 181.650 641.400 183.450 647.250 ;
        RECT 184.650 641.400 186.450 647.250 ;
        RECT 187.650 641.400 189.450 647.250 ;
        RECT 193.650 641.400 195.450 647.250 ;
        RECT 196.650 642.000 198.450 647.250 ;
        RECT 173.550 641.100 174.750 641.400 ;
        RECT 167.700 640.200 174.750 641.100 ;
        RECT 136.800 634.500 138.600 635.400 ;
        RECT 136.800 633.600 140.850 634.500 ;
        RECT 124.950 629.850 127.050 631.950 ;
        RECT 134.100 630.150 135.900 631.950 ;
        RECT 139.950 630.150 140.850 633.600 ;
        RECT 152.250 631.950 153.300 640.200 ;
        RECT 158.100 636.150 159.900 637.950 ;
        RECT 167.100 636.150 168.900 637.950 ;
        RECT 154.950 633.150 156.750 634.950 ;
        RECT 157.950 634.050 160.050 636.150 ;
        RECT 161.100 633.150 162.900 634.950 ;
        RECT 164.100 633.150 165.900 634.950 ;
        RECT 166.950 634.050 169.050 636.150 ;
        RECT 170.250 633.150 172.050 634.950 ;
        RECT 145.950 630.150 147.750 631.950 ;
        RECT 56.250 623.700 60.000 624.750 ;
        RECT 75.000 623.700 78.750 624.750 ;
        RECT 56.250 621.600 57.450 623.700 ;
        RECT 43.650 615.750 45.450 618.600 ;
        RECT 46.650 615.750 48.450 618.600 ;
        RECT 49.650 615.750 51.450 618.600 ;
        RECT 55.650 615.750 57.450 621.600 ;
        RECT 58.650 620.700 66.450 622.050 ;
        RECT 58.650 615.750 60.450 620.700 ;
        RECT 61.650 615.750 63.450 619.800 ;
        RECT 64.650 615.750 66.450 620.700 ;
        RECT 68.550 620.700 76.350 622.050 ;
        RECT 68.550 615.750 70.350 620.700 ;
        RECT 71.550 615.750 73.350 619.800 ;
        RECT 74.550 615.750 76.350 620.700 ;
        RECT 77.550 621.600 78.750 623.700 ;
        RECT 77.550 615.750 79.350 621.600 ;
        RECT 86.400 618.600 87.600 626.850 ;
        RECT 88.950 625.050 91.050 627.150 ;
        RECT 95.100 621.600 96.300 628.050 ;
        RECT 97.950 626.850 100.050 628.950 ;
        RECT 101.100 627.150 102.900 628.950 ;
        RECT 98.100 625.050 99.900 626.850 ;
        RECT 100.950 625.050 103.050 627.150 ;
        RECT 103.950 626.850 106.050 628.950 ;
        RECT 109.950 626.850 112.050 628.950 ;
        RECT 113.100 627.150 114.900 628.950 ;
        RECT 104.100 625.050 105.900 626.850 ;
        RECT 95.100 619.950 100.800 621.600 ;
        RECT 85.650 615.750 87.450 618.600 ;
        RECT 88.650 615.750 90.450 618.600 ;
        RECT 95.700 615.750 97.500 618.600 ;
        RECT 99.000 615.750 100.800 619.950 ;
        RECT 103.200 615.750 105.000 621.600 ;
        RECT 110.400 618.600 111.600 626.850 ;
        RECT 112.950 625.050 115.050 627.150 ;
        RECT 125.400 625.650 126.600 629.850 ;
        RECT 133.950 628.050 136.050 630.150 ;
        RECT 136.950 626.850 139.050 628.950 ;
        RECT 139.950 628.050 142.050 630.150 ;
        RECT 109.650 615.750 111.450 618.600 ;
        RECT 112.650 615.750 114.450 618.600 ;
        RECT 116.700 615.750 118.500 624.600 ;
        RECT 122.100 624.000 126.600 625.650 ;
        RECT 137.250 625.050 139.050 626.850 ;
        RECT 122.100 615.750 123.900 624.000 ;
        RECT 141.000 621.600 142.050 628.050 ;
        RECT 142.950 626.850 145.050 628.950 ;
        RECT 145.950 628.050 148.050 630.150 ;
        RECT 151.950 629.850 154.050 631.950 ;
        RECT 154.950 631.050 157.050 633.150 ;
        RECT 160.950 631.050 163.050 633.150 ;
        RECT 163.950 631.050 166.050 633.150 ;
        RECT 169.950 631.050 172.050 633.150 ;
        RECT 173.700 631.950 174.750 640.200 ;
        RECT 185.250 633.150 186.450 641.400 ;
        RECT 194.250 641.100 195.450 641.400 ;
        RECT 199.650 641.400 201.450 647.250 ;
        RECT 202.650 641.400 204.450 647.250 ;
        RECT 208.650 641.400 210.450 647.250 ;
        RECT 211.650 641.400 213.450 647.250 ;
        RECT 214.650 641.400 216.450 647.250 ;
        RECT 218.550 641.400 220.350 647.250 ;
        RECT 221.550 641.400 223.350 647.250 ;
        RECT 224.550 642.000 226.350 647.250 ;
        RECT 199.650 641.100 201.300 641.400 ;
        RECT 194.250 640.200 201.300 641.100 ;
        RECT 172.950 629.850 175.050 631.950 ;
        RECT 181.950 629.850 184.050 631.950 ;
        RECT 184.950 631.050 187.050 633.150 ;
        RECT 194.250 631.950 195.300 640.200 ;
        RECT 200.100 636.150 201.900 637.950 ;
        RECT 196.950 633.150 198.750 634.950 ;
        RECT 199.950 634.050 202.050 636.150 ;
        RECT 203.100 633.150 204.900 634.950 ;
        RECT 212.250 633.150 213.450 641.400 ;
        RECT 221.700 641.100 223.350 641.400 ;
        RECT 227.550 641.400 229.350 647.250 ;
        RECT 227.550 641.100 228.750 641.400 ;
        RECT 221.700 640.200 228.750 641.100 ;
        RECT 221.100 636.150 222.900 637.950 ;
        RECT 218.100 633.150 219.900 634.950 ;
        RECT 220.950 634.050 223.050 636.150 ;
        RECT 224.250 633.150 226.050 634.950 ;
        RECT 142.950 625.050 144.750 626.850 ;
        RECT 152.400 625.650 153.600 629.850 ;
        RECT 173.400 625.650 174.600 629.850 ;
        RECT 182.100 628.050 183.900 629.850 ;
        RECT 152.400 624.000 156.900 625.650 ;
        RECT 136.800 615.750 138.600 621.600 ;
        RECT 141.000 615.750 142.800 621.600 ;
        RECT 145.200 615.750 147.000 621.600 ;
        RECT 155.100 615.750 156.900 624.000 ;
        RECT 160.500 615.750 162.300 624.600 ;
        RECT 164.700 615.750 166.500 624.600 ;
        RECT 170.100 624.000 174.600 625.650 ;
        RECT 170.100 615.750 171.900 624.000 ;
        RECT 185.250 623.700 186.450 631.050 ;
        RECT 187.950 629.850 190.050 631.950 ;
        RECT 193.950 629.850 196.050 631.950 ;
        RECT 196.950 631.050 199.050 633.150 ;
        RECT 202.950 631.050 205.050 633.150 ;
        RECT 208.950 629.850 211.050 631.950 ;
        RECT 211.950 631.050 214.050 633.150 ;
        RECT 188.100 628.050 189.900 629.850 ;
        RECT 194.400 625.650 195.600 629.850 ;
        RECT 209.100 628.050 210.900 629.850 ;
        RECT 194.400 624.000 198.900 625.650 ;
        RECT 182.850 622.800 186.450 623.700 ;
        RECT 182.850 615.750 184.650 622.800 ;
        RECT 187.350 615.750 189.150 621.600 ;
        RECT 197.100 615.750 198.900 624.000 ;
        RECT 202.500 615.750 204.300 624.600 ;
        RECT 212.250 623.700 213.450 631.050 ;
        RECT 214.950 629.850 217.050 631.950 ;
        RECT 217.950 631.050 220.050 633.150 ;
        RECT 223.950 631.050 226.050 633.150 ;
        RECT 227.700 631.950 228.750 640.200 ;
        RECT 237.450 635.400 239.250 647.250 ;
        RECT 241.650 635.400 243.450 647.250 ;
        RECT 249.450 635.400 251.250 647.250 ;
        RECT 253.650 635.400 255.450 647.250 ;
        RECT 258.300 635.400 260.100 647.250 ;
        RECT 262.500 635.400 264.300 647.250 ;
        RECT 265.800 641.400 267.600 647.250 ;
        RECT 274.650 641.400 276.450 647.250 ;
        RECT 277.650 641.400 279.450 647.250 ;
        RECT 280.650 641.400 282.450 647.250 ;
        RECT 284.550 641.400 286.350 647.250 ;
        RECT 287.550 641.400 289.350 647.250 ;
        RECT 293.550 641.400 295.350 647.250 ;
        RECT 296.550 641.400 298.350 647.250 ;
        RECT 299.550 642.000 301.350 647.250 ;
        RECT 237.450 634.350 240.000 635.400 ;
        RECT 249.450 634.350 252.000 635.400 ;
        RECT 226.950 629.850 229.050 631.950 ;
        RECT 236.100 630.150 237.900 631.950 ;
        RECT 215.100 628.050 216.900 629.850 ;
        RECT 227.400 625.650 228.600 629.850 ;
        RECT 235.950 628.050 238.050 630.150 ;
        RECT 209.850 622.800 213.450 623.700 ;
        RECT 209.850 615.750 211.650 622.800 ;
        RECT 214.350 615.750 216.150 621.600 ;
        RECT 218.700 615.750 220.500 624.600 ;
        RECT 224.100 624.000 228.600 625.650 ;
        RECT 238.950 627.150 240.000 634.350 ;
        RECT 242.100 630.150 243.900 631.950 ;
        RECT 248.100 630.150 249.900 631.950 ;
        RECT 241.950 628.050 244.050 630.150 ;
        RECT 247.950 628.050 250.050 630.150 ;
        RECT 250.950 627.150 252.000 634.350 ;
        RECT 254.100 630.150 255.900 631.950 ;
        RECT 257.100 630.150 258.900 631.950 ;
        RECT 262.950 630.150 264.150 635.400 ;
        RECT 265.950 633.150 267.750 634.950 ;
        RECT 278.250 633.150 279.450 641.400 ;
        RECT 265.950 631.050 268.050 633.150 ;
        RECT 253.950 628.050 256.050 630.150 ;
        RECT 256.950 628.050 259.050 630.150 ;
        RECT 238.950 625.050 241.050 627.150 ;
        RECT 250.950 625.050 253.050 627.150 ;
        RECT 259.950 626.850 262.050 628.950 ;
        RECT 262.950 628.050 265.050 630.150 ;
        RECT 274.950 629.850 277.050 631.950 ;
        RECT 277.950 631.050 280.050 633.150 ;
        RECT 275.100 628.050 276.900 629.850 ;
        RECT 260.100 625.050 261.900 626.850 ;
        RECT 224.100 615.750 225.900 624.000 ;
        RECT 238.950 618.600 240.000 625.050 ;
        RECT 250.950 618.600 252.000 625.050 ;
        RECT 263.850 624.750 265.050 628.050 ;
        RECT 264.000 623.700 267.750 624.750 ;
        RECT 278.250 623.700 279.450 631.050 ;
        RECT 280.950 629.850 283.050 631.950 ;
        RECT 281.100 628.050 282.900 629.850 ;
        RECT 287.400 628.950 288.600 641.400 ;
        RECT 296.700 641.100 298.350 641.400 ;
        RECT 302.550 641.400 304.350 647.250 ;
        RECT 308.550 641.400 310.350 647.250 ;
        RECT 311.550 641.400 313.350 647.250 ;
        RECT 314.550 642.000 316.350 647.250 ;
        RECT 302.550 641.100 303.750 641.400 ;
        RECT 296.700 640.200 303.750 641.100 ;
        RECT 311.700 641.100 313.350 641.400 ;
        RECT 317.550 641.400 319.350 647.250 ;
        RECT 317.550 641.100 318.750 641.400 ;
        RECT 311.700 640.200 318.750 641.100 ;
        RECT 296.100 636.150 297.900 637.950 ;
        RECT 293.100 633.150 294.900 634.950 ;
        RECT 295.950 634.050 298.050 636.150 ;
        RECT 299.250 633.150 301.050 634.950 ;
        RECT 292.950 631.050 295.050 633.150 ;
        RECT 298.950 631.050 301.050 633.150 ;
        RECT 302.700 631.950 303.750 640.200 ;
        RECT 311.100 636.150 312.900 637.950 ;
        RECT 308.100 633.150 309.900 634.950 ;
        RECT 310.950 634.050 313.050 636.150 ;
        RECT 314.250 633.150 316.050 634.950 ;
        RECT 301.950 629.850 304.050 631.950 ;
        RECT 307.950 631.050 310.050 633.150 ;
        RECT 313.950 631.050 316.050 633.150 ;
        RECT 317.700 631.950 318.750 640.200 ;
        RECT 324.150 635.400 325.950 647.250 ;
        RECT 327.150 641.400 328.950 647.250 ;
        RECT 332.250 641.400 334.050 647.250 ;
        RECT 337.050 641.400 338.850 647.250 ;
        RECT 332.550 640.500 333.750 641.400 ;
        RECT 340.050 640.500 341.850 647.250 ;
        RECT 343.950 641.400 345.750 647.250 ;
        RECT 348.150 641.400 349.950 647.250 ;
        RECT 352.650 644.400 354.450 647.250 ;
        RECT 328.950 638.400 333.750 640.500 ;
        RECT 336.150 638.700 343.050 640.500 ;
        RECT 348.150 639.300 352.050 641.400 ;
        RECT 332.550 637.500 333.750 638.400 ;
        RECT 345.450 637.800 347.250 638.400 ;
        RECT 332.550 636.300 340.050 637.500 ;
        RECT 338.250 635.700 340.050 636.300 ;
        RECT 340.950 636.900 347.250 637.800 ;
        RECT 324.150 634.800 335.250 635.400 ;
        RECT 340.950 634.800 341.850 636.900 ;
        RECT 345.450 636.600 347.250 636.900 ;
        RECT 348.150 636.600 350.850 638.400 ;
        RECT 348.150 635.700 349.050 636.600 ;
        RECT 324.150 634.200 341.850 634.800 ;
        RECT 316.950 629.850 319.050 631.950 ;
        RECT 284.100 627.150 285.900 628.950 ;
        RECT 283.950 625.050 286.050 627.150 ;
        RECT 286.950 626.850 289.050 628.950 ;
        RECT 257.550 620.700 265.350 622.050 ;
        RECT 235.650 615.750 237.450 618.600 ;
        RECT 238.650 615.750 240.450 618.600 ;
        RECT 241.650 615.750 243.450 618.600 ;
        RECT 247.650 615.750 249.450 618.600 ;
        RECT 250.650 615.750 252.450 618.600 ;
        RECT 253.650 615.750 255.450 618.600 ;
        RECT 257.550 615.750 259.350 620.700 ;
        RECT 260.550 615.750 262.350 619.800 ;
        RECT 263.550 615.750 265.350 620.700 ;
        RECT 266.550 621.600 267.750 623.700 ;
        RECT 275.850 622.800 279.450 623.700 ;
        RECT 266.550 615.750 268.350 621.600 ;
        RECT 275.850 615.750 277.650 622.800 ;
        RECT 280.350 615.750 282.150 621.600 ;
        RECT 287.400 618.600 288.600 626.850 ;
        RECT 302.400 625.650 303.600 629.850 ;
        RECT 317.400 625.650 318.600 629.850 ;
        RECT 284.550 615.750 286.350 618.600 ;
        RECT 287.550 615.750 289.350 618.600 ;
        RECT 293.700 615.750 295.500 624.600 ;
        RECT 299.100 624.000 303.600 625.650 ;
        RECT 299.100 615.750 300.900 624.000 ;
        RECT 308.700 615.750 310.500 624.600 ;
        RECT 314.100 624.000 318.600 625.650 ;
        RECT 314.100 615.750 315.900 624.000 ;
        RECT 324.150 621.600 325.050 634.200 ;
        RECT 333.450 633.900 341.850 634.200 ;
        RECT 343.050 634.800 349.050 635.700 ;
        RECT 349.950 634.800 352.050 635.700 ;
        RECT 355.650 635.400 357.450 647.250 ;
        RECT 333.450 633.600 335.250 633.900 ;
        RECT 343.050 630.150 343.950 634.800 ;
        RECT 349.950 633.600 354.150 634.800 ;
        RECT 353.250 631.800 355.050 633.600 ;
        RECT 334.950 629.100 337.050 630.150 ;
        RECT 326.100 627.150 327.900 628.950 ;
        RECT 329.100 628.050 337.050 629.100 ;
        RECT 340.950 628.050 343.950 630.150 ;
        RECT 329.100 627.300 330.900 628.050 ;
        RECT 327.000 626.400 327.900 627.150 ;
        RECT 332.100 626.400 333.900 627.000 ;
        RECT 327.000 625.200 333.900 626.400 ;
        RECT 332.850 624.000 333.900 625.200 ;
        RECT 343.050 624.000 343.950 628.050 ;
        RECT 352.950 627.750 355.050 628.050 ;
        RECT 351.150 625.950 355.050 627.750 ;
        RECT 356.250 625.950 357.450 635.400 ;
        RECT 359.550 641.400 361.350 647.250 ;
        RECT 359.550 634.500 360.750 641.400 ;
        RECT 362.850 635.400 364.650 647.250 ;
        RECT 365.850 635.400 367.650 647.250 ;
        RECT 373.650 641.400 375.450 647.250 ;
        RECT 376.650 641.400 378.450 647.250 ;
        RECT 359.550 633.600 365.250 634.500 ;
        RECT 363.000 632.700 365.250 633.600 ;
        RECT 359.100 630.150 360.900 631.950 ;
        RECT 358.950 628.050 361.050 630.150 ;
        RECT 332.850 623.100 343.950 624.000 ;
        RECT 352.950 623.850 357.450 625.950 ;
        RECT 332.850 622.200 333.900 623.100 ;
        RECT 343.050 622.800 343.950 623.100 ;
        RECT 324.150 615.750 325.950 621.600 ;
        RECT 328.950 619.500 331.050 621.600 ;
        RECT 332.550 620.400 334.350 622.200 ;
        RECT 335.850 621.450 337.650 622.200 ;
        RECT 335.850 620.400 340.800 621.450 ;
        RECT 343.050 621.000 344.850 622.800 ;
        RECT 356.250 621.600 357.450 623.850 ;
        RECT 363.000 624.300 364.050 632.700 ;
        RECT 366.150 630.150 367.350 635.400 ;
        RECT 364.950 628.050 367.350 630.150 ;
        RECT 374.400 628.950 375.600 641.400 ;
        RECT 384.450 635.400 386.250 647.250 ;
        RECT 388.650 635.400 390.450 647.250 ;
        RECT 392.550 635.400 394.350 647.250 ;
        RECT 395.550 644.400 397.350 647.250 ;
        RECT 400.050 641.400 401.850 647.250 ;
        RECT 404.250 641.400 406.050 647.250 ;
        RECT 397.950 639.300 401.850 641.400 ;
        RECT 408.150 640.500 409.950 647.250 ;
        RECT 411.150 641.400 412.950 647.250 ;
        RECT 415.950 641.400 417.750 647.250 ;
        RECT 421.050 641.400 422.850 647.250 ;
        RECT 416.250 640.500 417.450 641.400 ;
        RECT 406.950 638.700 413.850 640.500 ;
        RECT 416.250 638.400 421.050 640.500 ;
        RECT 399.150 636.600 401.850 638.400 ;
        RECT 402.750 637.800 404.550 638.400 ;
        RECT 402.750 636.900 409.050 637.800 ;
        RECT 416.250 637.500 417.450 638.400 ;
        RECT 402.750 636.600 404.550 636.900 ;
        RECT 400.950 635.700 401.850 636.600 ;
        RECT 384.450 634.350 387.000 635.400 ;
        RECT 383.100 630.150 384.900 631.950 ;
        RECT 363.000 623.400 365.250 624.300 ;
        RECT 349.950 620.700 352.050 621.600 ;
        RECT 330.000 618.600 331.050 619.500 ;
        RECT 339.750 618.600 340.800 620.400 ;
        RECT 348.300 619.500 352.050 620.700 ;
        RECT 348.300 618.600 349.350 619.500 ;
        RECT 327.150 615.750 328.950 618.600 ;
        RECT 330.000 617.700 333.750 618.600 ;
        RECT 331.950 615.750 333.750 617.700 ;
        RECT 336.450 615.750 338.250 618.600 ;
        RECT 339.750 615.750 341.550 618.600 ;
        RECT 343.650 615.750 345.450 618.600 ;
        RECT 347.850 615.750 349.650 618.600 ;
        RECT 352.350 615.750 354.150 618.600 ;
        RECT 355.650 615.750 357.450 621.600 ;
        RECT 360.150 622.500 365.250 623.400 ;
        RECT 360.150 618.600 361.350 622.500 ;
        RECT 366.150 621.600 367.350 628.050 ;
        RECT 373.950 626.850 376.050 628.950 ;
        RECT 377.100 627.150 378.900 628.950 ;
        RECT 382.950 628.050 385.050 630.150 ;
        RECT 385.950 627.150 387.000 634.350 ;
        RECT 389.100 630.150 390.900 631.950 ;
        RECT 388.950 628.050 391.050 630.150 ;
        RECT 359.550 615.750 361.350 618.600 ;
        RECT 362.850 615.750 364.650 621.600 ;
        RECT 365.850 615.750 367.650 621.600 ;
        RECT 374.400 618.600 375.600 626.850 ;
        RECT 376.950 625.050 379.050 627.150 ;
        RECT 385.950 625.050 388.050 627.150 ;
        RECT 392.550 625.950 393.750 635.400 ;
        RECT 397.950 634.800 400.050 635.700 ;
        RECT 400.950 634.800 406.950 635.700 ;
        RECT 395.850 633.600 400.050 634.800 ;
        RECT 394.950 631.800 396.750 633.600 ;
        RECT 406.050 630.150 406.950 634.800 ;
        RECT 408.150 634.800 409.050 636.900 ;
        RECT 409.950 636.300 417.450 637.500 ;
        RECT 409.950 635.700 411.750 636.300 ;
        RECT 424.050 635.400 425.850 647.250 ;
        RECT 428.550 641.400 430.350 647.250 ;
        RECT 431.550 641.400 433.350 647.250 ;
        RECT 414.750 634.800 425.850 635.400 ;
        RECT 408.150 634.200 425.850 634.800 ;
        RECT 408.150 633.900 416.550 634.200 ;
        RECT 414.750 633.600 416.550 633.900 ;
        RECT 406.050 628.050 409.050 630.150 ;
        RECT 412.950 629.100 415.050 630.150 ;
        RECT 412.950 628.050 420.900 629.100 ;
        RECT 394.950 627.750 397.050 628.050 ;
        RECT 394.950 625.950 398.850 627.750 ;
        RECT 385.950 618.600 387.000 625.050 ;
        RECT 392.550 623.850 397.050 625.950 ;
        RECT 406.050 624.000 406.950 628.050 ;
        RECT 419.100 627.300 420.900 628.050 ;
        RECT 422.100 627.150 423.900 628.950 ;
        RECT 416.100 626.400 417.900 627.000 ;
        RECT 422.100 626.400 423.000 627.150 ;
        RECT 416.100 625.200 423.000 626.400 ;
        RECT 416.100 624.000 417.150 625.200 ;
        RECT 392.550 621.600 393.750 623.850 ;
        RECT 406.050 623.100 417.150 624.000 ;
        RECT 406.050 622.800 406.950 623.100 ;
        RECT 373.650 615.750 375.450 618.600 ;
        RECT 376.650 615.750 378.450 618.600 ;
        RECT 382.650 615.750 384.450 618.600 ;
        RECT 385.650 615.750 387.450 618.600 ;
        RECT 388.650 615.750 390.450 618.600 ;
        RECT 392.550 615.750 394.350 621.600 ;
        RECT 397.950 620.700 400.050 621.600 ;
        RECT 405.150 621.000 406.950 622.800 ;
        RECT 416.100 622.200 417.150 623.100 ;
        RECT 412.350 621.450 414.150 622.200 ;
        RECT 397.950 619.500 401.700 620.700 ;
        RECT 400.650 618.600 401.700 619.500 ;
        RECT 409.200 620.400 414.150 621.450 ;
        RECT 415.650 620.400 417.450 622.200 ;
        RECT 424.950 621.600 425.850 634.200 ;
        RECT 431.400 628.950 432.600 641.400 ;
        RECT 441.450 635.400 443.250 647.250 ;
        RECT 445.650 635.400 447.450 647.250 ;
        RECT 450.300 635.400 452.100 647.250 ;
        RECT 454.500 635.400 456.300 647.250 ;
        RECT 457.800 641.400 459.600 647.250 ;
        RECT 464.550 641.400 466.350 647.250 ;
        RECT 467.550 641.400 469.350 647.250 ;
        RECT 470.550 641.400 472.350 647.250 ;
        RECT 478.650 641.400 480.450 647.250 ;
        RECT 481.650 641.400 483.450 647.250 ;
        RECT 484.650 641.400 486.450 647.250 ;
        RECT 490.650 641.400 492.450 647.250 ;
        RECT 493.650 641.400 495.450 647.250 ;
        RECT 496.650 641.400 498.450 647.250 ;
        RECT 441.450 634.350 444.000 635.400 ;
        RECT 440.100 630.150 441.900 631.950 ;
        RECT 428.100 627.150 429.900 628.950 ;
        RECT 427.950 625.050 430.050 627.150 ;
        RECT 430.950 626.850 433.050 628.950 ;
        RECT 439.950 628.050 442.050 630.150 ;
        RECT 442.950 627.150 444.000 634.350 ;
        RECT 446.100 630.150 447.900 631.950 ;
        RECT 449.100 630.150 450.900 631.950 ;
        RECT 454.950 630.150 456.150 635.400 ;
        RECT 457.950 633.150 459.750 634.950 ;
        RECT 467.550 633.150 468.750 641.400 ;
        RECT 482.250 633.150 483.450 641.400 ;
        RECT 494.250 633.150 495.450 641.400 ;
        RECT 500.550 635.400 502.350 647.250 ;
        RECT 504.750 635.400 506.550 647.250 ;
        RECT 504.000 634.350 506.550 635.400 ;
        RECT 513.150 635.400 514.950 647.250 ;
        RECT 516.150 641.400 517.950 647.250 ;
        RECT 521.250 641.400 523.050 647.250 ;
        RECT 526.050 641.400 527.850 647.250 ;
        RECT 521.550 640.500 522.750 641.400 ;
        RECT 529.050 640.500 530.850 647.250 ;
        RECT 532.950 641.400 534.750 647.250 ;
        RECT 537.150 641.400 538.950 647.250 ;
        RECT 541.650 644.400 543.450 647.250 ;
        RECT 517.950 638.400 522.750 640.500 ;
        RECT 525.150 638.700 532.050 640.500 ;
        RECT 537.150 639.300 541.050 641.400 ;
        RECT 521.550 637.500 522.750 638.400 ;
        RECT 534.450 637.800 536.250 638.400 ;
        RECT 521.550 636.300 529.050 637.500 ;
        RECT 527.250 635.700 529.050 636.300 ;
        RECT 529.950 636.900 536.250 637.800 ;
        RECT 513.150 634.800 524.250 635.400 ;
        RECT 529.950 634.800 530.850 636.900 ;
        RECT 534.450 636.600 536.250 636.900 ;
        RECT 537.150 636.600 539.850 638.400 ;
        RECT 537.150 635.700 538.050 636.600 ;
        RECT 457.950 631.050 460.050 633.150 ;
        RECT 445.950 628.050 448.050 630.150 ;
        RECT 448.950 628.050 451.050 630.150 ;
        RECT 409.200 618.600 410.250 620.400 ;
        RECT 418.950 619.500 421.050 621.600 ;
        RECT 418.950 618.600 420.000 619.500 ;
        RECT 395.850 615.750 397.650 618.600 ;
        RECT 400.350 615.750 402.150 618.600 ;
        RECT 404.550 615.750 406.350 618.600 ;
        RECT 408.450 615.750 410.250 618.600 ;
        RECT 411.750 615.750 413.550 618.600 ;
        RECT 416.250 617.700 420.000 618.600 ;
        RECT 416.250 615.750 418.050 617.700 ;
        RECT 421.050 615.750 422.850 618.600 ;
        RECT 424.050 615.750 425.850 621.600 ;
        RECT 431.400 618.600 432.600 626.850 ;
        RECT 442.950 625.050 445.050 627.150 ;
        RECT 451.950 626.850 454.050 628.950 ;
        RECT 454.950 628.050 457.050 630.150 ;
        RECT 463.950 629.850 466.050 631.950 ;
        RECT 466.950 631.050 469.050 633.150 ;
        RECT 464.100 628.050 465.900 629.850 ;
        RECT 452.100 625.050 453.900 626.850 ;
        RECT 442.950 618.600 444.000 625.050 ;
        RECT 455.850 624.750 457.050 628.050 ;
        RECT 456.000 623.700 459.750 624.750 ;
        RECT 449.550 620.700 457.350 622.050 ;
        RECT 428.550 615.750 430.350 618.600 ;
        RECT 431.550 615.750 433.350 618.600 ;
        RECT 439.650 615.750 441.450 618.600 ;
        RECT 442.650 615.750 444.450 618.600 ;
        RECT 445.650 615.750 447.450 618.600 ;
        RECT 449.550 615.750 451.350 620.700 ;
        RECT 452.550 615.750 454.350 619.800 ;
        RECT 455.550 615.750 457.350 620.700 ;
        RECT 458.550 621.600 459.750 623.700 ;
        RECT 467.550 623.700 468.750 631.050 ;
        RECT 469.950 629.850 472.050 631.950 ;
        RECT 478.950 629.850 481.050 631.950 ;
        RECT 481.950 631.050 484.050 633.150 ;
        RECT 470.100 628.050 471.900 629.850 ;
        RECT 479.100 628.050 480.900 629.850 ;
        RECT 482.250 623.700 483.450 631.050 ;
        RECT 484.950 629.850 487.050 631.950 ;
        RECT 490.950 629.850 493.050 631.950 ;
        RECT 493.950 631.050 496.050 633.150 ;
        RECT 485.100 628.050 486.900 629.850 ;
        RECT 491.100 628.050 492.900 629.850 ;
        RECT 494.250 623.700 495.450 631.050 ;
        RECT 496.950 629.850 499.050 631.950 ;
        RECT 500.100 630.150 501.900 631.950 ;
        RECT 497.100 628.050 498.900 629.850 ;
        RECT 499.950 628.050 502.050 630.150 ;
        RECT 504.000 627.150 505.050 634.350 ;
        RECT 513.150 634.200 530.850 634.800 ;
        RECT 506.100 630.150 507.900 631.950 ;
        RECT 505.950 628.050 508.050 630.150 ;
        RECT 502.950 625.050 505.050 627.150 ;
        RECT 467.550 622.800 471.150 623.700 ;
        RECT 458.550 615.750 460.350 621.600 ;
        RECT 464.850 615.750 466.650 621.600 ;
        RECT 469.350 615.750 471.150 622.800 ;
        RECT 479.850 622.800 483.450 623.700 ;
        RECT 491.850 622.800 495.450 623.700 ;
        RECT 479.850 615.750 481.650 622.800 ;
        RECT 484.350 615.750 486.150 621.600 ;
        RECT 491.850 615.750 493.650 622.800 ;
        RECT 496.350 615.750 498.150 621.600 ;
        RECT 504.000 618.600 505.050 625.050 ;
        RECT 513.150 621.600 514.050 634.200 ;
        RECT 522.450 633.900 530.850 634.200 ;
        RECT 532.050 634.800 538.050 635.700 ;
        RECT 538.950 634.800 541.050 635.700 ;
        RECT 544.650 635.400 546.450 647.250 ;
        RECT 550.650 641.400 552.450 647.250 ;
        RECT 553.650 641.400 555.450 647.250 ;
        RECT 556.650 641.400 558.450 647.250 ;
        RECT 522.450 633.600 524.250 633.900 ;
        RECT 532.050 630.150 532.950 634.800 ;
        RECT 538.950 633.600 543.150 634.800 ;
        RECT 542.250 631.800 544.050 633.600 ;
        RECT 523.950 629.100 526.050 630.150 ;
        RECT 515.100 627.150 516.900 628.950 ;
        RECT 518.100 628.050 526.050 629.100 ;
        RECT 529.950 628.050 532.950 630.150 ;
        RECT 518.100 627.300 519.900 628.050 ;
        RECT 516.000 626.400 516.900 627.150 ;
        RECT 521.100 626.400 522.900 627.000 ;
        RECT 516.000 625.200 522.900 626.400 ;
        RECT 521.850 624.000 522.900 625.200 ;
        RECT 532.050 624.000 532.950 628.050 ;
        RECT 541.950 627.750 544.050 628.050 ;
        RECT 540.150 625.950 544.050 627.750 ;
        RECT 545.250 625.950 546.450 635.400 ;
        RECT 554.250 633.150 555.450 641.400 ;
        RECT 560.550 635.400 562.350 647.250 ;
        RECT 564.750 635.400 566.550 647.250 ;
        RECT 564.000 634.350 566.550 635.400 ;
        RECT 572.550 635.400 574.350 647.250 ;
        RECT 575.550 644.400 577.350 647.250 ;
        RECT 580.050 641.400 581.850 647.250 ;
        RECT 584.250 641.400 586.050 647.250 ;
        RECT 577.950 639.300 581.850 641.400 ;
        RECT 588.150 640.500 589.950 647.250 ;
        RECT 591.150 641.400 592.950 647.250 ;
        RECT 595.950 641.400 597.750 647.250 ;
        RECT 601.050 641.400 602.850 647.250 ;
        RECT 596.250 640.500 597.450 641.400 ;
        RECT 586.950 638.700 593.850 640.500 ;
        RECT 596.250 638.400 601.050 640.500 ;
        RECT 579.150 636.600 581.850 638.400 ;
        RECT 582.750 637.800 584.550 638.400 ;
        RECT 582.750 636.900 589.050 637.800 ;
        RECT 596.250 637.500 597.450 638.400 ;
        RECT 582.750 636.600 584.550 636.900 ;
        RECT 580.950 635.700 581.850 636.600 ;
        RECT 550.950 629.850 553.050 631.950 ;
        RECT 553.950 631.050 556.050 633.150 ;
        RECT 551.100 628.050 552.900 629.850 ;
        RECT 521.850 623.100 532.950 624.000 ;
        RECT 541.950 623.850 546.450 625.950 ;
        RECT 521.850 622.200 522.900 623.100 ;
        RECT 532.050 622.800 532.950 623.100 ;
        RECT 500.550 615.750 502.350 618.600 ;
        RECT 503.550 615.750 505.350 618.600 ;
        RECT 506.550 615.750 508.350 618.600 ;
        RECT 513.150 615.750 514.950 621.600 ;
        RECT 517.950 619.500 520.050 621.600 ;
        RECT 521.550 620.400 523.350 622.200 ;
        RECT 524.850 621.450 526.650 622.200 ;
        RECT 524.850 620.400 529.800 621.450 ;
        RECT 532.050 621.000 533.850 622.800 ;
        RECT 545.250 621.600 546.450 623.850 ;
        RECT 554.250 623.700 555.450 631.050 ;
        RECT 556.950 629.850 559.050 631.950 ;
        RECT 560.100 630.150 561.900 631.950 ;
        RECT 557.100 628.050 558.900 629.850 ;
        RECT 559.950 628.050 562.050 630.150 ;
        RECT 564.000 627.150 565.050 634.350 ;
        RECT 566.100 630.150 567.900 631.950 ;
        RECT 565.950 628.050 568.050 630.150 ;
        RECT 562.950 625.050 565.050 627.150 ;
        RECT 538.950 620.700 541.050 621.600 ;
        RECT 519.000 618.600 520.050 619.500 ;
        RECT 528.750 618.600 529.800 620.400 ;
        RECT 537.300 619.500 541.050 620.700 ;
        RECT 537.300 618.600 538.350 619.500 ;
        RECT 516.150 615.750 517.950 618.600 ;
        RECT 519.000 617.700 522.750 618.600 ;
        RECT 520.950 615.750 522.750 617.700 ;
        RECT 525.450 615.750 527.250 618.600 ;
        RECT 528.750 615.750 530.550 618.600 ;
        RECT 532.650 615.750 534.450 618.600 ;
        RECT 536.850 615.750 538.650 618.600 ;
        RECT 541.350 615.750 543.150 618.600 ;
        RECT 544.650 615.750 546.450 621.600 ;
        RECT 551.850 622.800 555.450 623.700 ;
        RECT 551.850 615.750 553.650 622.800 ;
        RECT 556.350 615.750 558.150 621.600 ;
        RECT 564.000 618.600 565.050 625.050 ;
        RECT 572.550 625.950 573.750 635.400 ;
        RECT 577.950 634.800 580.050 635.700 ;
        RECT 580.950 634.800 586.950 635.700 ;
        RECT 575.850 633.600 580.050 634.800 ;
        RECT 574.950 631.800 576.750 633.600 ;
        RECT 586.050 630.150 586.950 634.800 ;
        RECT 588.150 634.800 589.050 636.900 ;
        RECT 589.950 636.300 597.450 637.500 ;
        RECT 589.950 635.700 591.750 636.300 ;
        RECT 604.050 635.400 605.850 647.250 ;
        RECT 608.550 635.400 610.350 647.250 ;
        RECT 612.750 635.400 614.550 647.250 ;
        RECT 622.650 635.400 624.450 647.250 ;
        RECT 625.650 636.300 627.450 647.250 ;
        RECT 628.650 637.200 630.450 647.250 ;
        RECT 631.650 636.300 633.450 647.250 ;
        RECT 625.650 635.400 633.450 636.300 ;
        RECT 635.550 641.400 637.350 647.250 ;
        RECT 594.750 634.800 605.850 635.400 ;
        RECT 588.150 634.200 605.850 634.800 ;
        RECT 588.150 633.900 596.550 634.200 ;
        RECT 594.750 633.600 596.550 633.900 ;
        RECT 586.050 628.050 589.050 630.150 ;
        RECT 592.950 629.100 595.050 630.150 ;
        RECT 592.950 628.050 600.900 629.100 ;
        RECT 574.950 627.750 577.050 628.050 ;
        RECT 574.950 625.950 578.850 627.750 ;
        RECT 572.550 623.850 577.050 625.950 ;
        RECT 586.050 624.000 586.950 628.050 ;
        RECT 599.100 627.300 600.900 628.050 ;
        RECT 602.100 627.150 603.900 628.950 ;
        RECT 596.100 626.400 597.900 627.000 ;
        RECT 602.100 626.400 603.000 627.150 ;
        RECT 596.100 625.200 603.000 626.400 ;
        RECT 596.100 624.000 597.150 625.200 ;
        RECT 572.550 621.600 573.750 623.850 ;
        RECT 586.050 623.100 597.150 624.000 ;
        RECT 586.050 622.800 586.950 623.100 ;
        RECT 560.550 615.750 562.350 618.600 ;
        RECT 563.550 615.750 565.350 618.600 ;
        RECT 566.550 615.750 568.350 618.600 ;
        RECT 572.550 615.750 574.350 621.600 ;
        RECT 577.950 620.700 580.050 621.600 ;
        RECT 585.150 621.000 586.950 622.800 ;
        RECT 596.100 622.200 597.150 623.100 ;
        RECT 592.350 621.450 594.150 622.200 ;
        RECT 577.950 619.500 581.700 620.700 ;
        RECT 580.650 618.600 581.700 619.500 ;
        RECT 589.200 620.400 594.150 621.450 ;
        RECT 595.650 620.400 597.450 622.200 ;
        RECT 604.950 621.600 605.850 634.200 ;
        RECT 612.000 634.350 614.550 635.400 ;
        RECT 608.100 630.150 609.900 631.950 ;
        RECT 607.950 628.050 610.050 630.150 ;
        RECT 612.000 627.150 613.050 634.350 ;
        RECT 614.100 630.150 615.900 631.950 ;
        RECT 623.100 630.150 624.300 635.400 ;
        RECT 635.550 634.500 636.750 641.400 ;
        RECT 638.850 635.400 640.650 647.250 ;
        RECT 641.850 635.400 643.650 647.250 ;
        RECT 651.450 635.400 653.250 647.250 ;
        RECT 655.650 635.400 657.450 647.250 ;
        RECT 661.650 635.400 663.450 647.250 ;
        RECT 664.650 636.300 666.450 647.250 ;
        RECT 667.650 637.200 669.450 647.250 ;
        RECT 670.650 636.300 672.450 647.250 ;
        RECT 664.650 635.400 672.450 636.300 ;
        RECT 674.550 635.400 676.350 647.250 ;
        RECT 677.550 644.400 679.350 647.250 ;
        RECT 682.050 641.400 683.850 647.250 ;
        RECT 686.250 641.400 688.050 647.250 ;
        RECT 679.950 639.300 683.850 641.400 ;
        RECT 690.150 640.500 691.950 647.250 ;
        RECT 693.150 641.400 694.950 647.250 ;
        RECT 697.950 641.400 699.750 647.250 ;
        RECT 703.050 641.400 704.850 647.250 ;
        RECT 698.250 640.500 699.450 641.400 ;
        RECT 688.950 638.700 695.850 640.500 ;
        RECT 698.250 638.400 703.050 640.500 ;
        RECT 681.150 636.600 683.850 638.400 ;
        RECT 684.750 637.800 686.550 638.400 ;
        RECT 684.750 636.900 691.050 637.800 ;
        RECT 698.250 637.500 699.450 638.400 ;
        RECT 684.750 636.600 686.550 636.900 ;
        RECT 682.950 635.700 683.850 636.600 ;
        RECT 635.550 633.600 641.250 634.500 ;
        RECT 639.000 632.700 641.250 633.600 ;
        RECT 635.100 630.150 636.900 631.950 ;
        RECT 613.950 628.050 616.050 630.150 ;
        RECT 622.950 628.050 625.050 630.150 ;
        RECT 610.950 625.050 613.050 627.150 ;
        RECT 589.200 618.600 590.250 620.400 ;
        RECT 598.950 619.500 601.050 621.600 ;
        RECT 598.950 618.600 600.000 619.500 ;
        RECT 575.850 615.750 577.650 618.600 ;
        RECT 580.350 615.750 582.150 618.600 ;
        RECT 584.550 615.750 586.350 618.600 ;
        RECT 588.450 615.750 590.250 618.600 ;
        RECT 591.750 615.750 593.550 618.600 ;
        RECT 596.250 617.700 600.000 618.600 ;
        RECT 596.250 615.750 598.050 617.700 ;
        RECT 601.050 615.750 602.850 618.600 ;
        RECT 604.050 615.750 605.850 621.600 ;
        RECT 612.000 618.600 613.050 625.050 ;
        RECT 623.100 621.600 624.300 628.050 ;
        RECT 625.950 626.850 628.050 628.950 ;
        RECT 629.100 627.150 630.900 628.950 ;
        RECT 626.100 625.050 627.900 626.850 ;
        RECT 628.950 625.050 631.050 627.150 ;
        RECT 631.950 626.850 634.050 628.950 ;
        RECT 634.950 628.050 637.050 630.150 ;
        RECT 632.100 625.050 633.900 626.850 ;
        RECT 639.000 624.300 640.050 632.700 ;
        RECT 642.150 630.150 643.350 635.400 ;
        RECT 651.450 634.350 654.000 635.400 ;
        RECT 650.100 630.150 651.900 631.950 ;
        RECT 640.950 628.050 643.350 630.150 ;
        RECT 649.950 628.050 652.050 630.150 ;
        RECT 639.000 623.400 641.250 624.300 ;
        RECT 636.150 622.500 641.250 623.400 ;
        RECT 623.100 619.950 628.800 621.600 ;
        RECT 608.550 615.750 610.350 618.600 ;
        RECT 611.550 615.750 613.350 618.600 ;
        RECT 614.550 615.750 616.350 618.600 ;
        RECT 623.700 615.750 625.500 618.600 ;
        RECT 627.000 615.750 628.800 619.950 ;
        RECT 631.200 615.750 633.000 621.600 ;
        RECT 636.150 618.600 637.350 622.500 ;
        RECT 642.150 621.600 643.350 628.050 ;
        RECT 652.950 627.150 654.000 634.350 ;
        RECT 656.100 630.150 657.900 631.950 ;
        RECT 662.100 630.150 663.300 635.400 ;
        RECT 655.950 628.050 658.050 630.150 ;
        RECT 661.950 628.050 664.050 630.150 ;
        RECT 652.950 625.050 655.050 627.150 ;
        RECT 635.550 615.750 637.350 618.600 ;
        RECT 638.850 615.750 640.650 621.600 ;
        RECT 641.850 615.750 643.650 621.600 ;
        RECT 652.950 618.600 654.000 625.050 ;
        RECT 662.100 621.600 663.300 628.050 ;
        RECT 664.950 626.850 667.050 628.950 ;
        RECT 668.100 627.150 669.900 628.950 ;
        RECT 665.100 625.050 666.900 626.850 ;
        RECT 667.950 625.050 670.050 627.150 ;
        RECT 670.950 626.850 673.050 628.950 ;
        RECT 671.100 625.050 672.900 626.850 ;
        RECT 674.550 625.950 675.750 635.400 ;
        RECT 679.950 634.800 682.050 635.700 ;
        RECT 682.950 634.800 688.950 635.700 ;
        RECT 677.850 633.600 682.050 634.800 ;
        RECT 676.950 631.800 678.750 633.600 ;
        RECT 688.050 630.150 688.950 634.800 ;
        RECT 690.150 634.800 691.050 636.900 ;
        RECT 691.950 636.300 699.450 637.500 ;
        RECT 691.950 635.700 693.750 636.300 ;
        RECT 706.050 635.400 707.850 647.250 ;
        RECT 696.750 634.800 707.850 635.400 ;
        RECT 690.150 634.200 707.850 634.800 ;
        RECT 690.150 633.900 698.550 634.200 ;
        RECT 696.750 633.600 698.550 633.900 ;
        RECT 688.050 628.050 691.050 630.150 ;
        RECT 694.950 629.100 697.050 630.150 ;
        RECT 694.950 628.050 702.900 629.100 ;
        RECT 676.950 627.750 679.050 628.050 ;
        RECT 676.950 625.950 680.850 627.750 ;
        RECT 674.550 623.850 679.050 625.950 ;
        RECT 688.050 624.000 688.950 628.050 ;
        RECT 701.100 627.300 702.900 628.050 ;
        RECT 704.100 627.150 705.900 628.950 ;
        RECT 698.100 626.400 699.900 627.000 ;
        RECT 704.100 626.400 705.000 627.150 ;
        RECT 698.100 625.200 705.000 626.400 ;
        RECT 698.100 624.000 699.150 625.200 ;
        RECT 674.550 621.600 675.750 623.850 ;
        RECT 688.050 623.100 699.150 624.000 ;
        RECT 688.050 622.800 688.950 623.100 ;
        RECT 662.100 619.950 667.800 621.600 ;
        RECT 649.650 615.750 651.450 618.600 ;
        RECT 652.650 615.750 654.450 618.600 ;
        RECT 655.650 615.750 657.450 618.600 ;
        RECT 662.700 615.750 664.500 618.600 ;
        RECT 666.000 615.750 667.800 619.950 ;
        RECT 670.200 615.750 672.000 621.600 ;
        RECT 674.550 615.750 676.350 621.600 ;
        RECT 679.950 620.700 682.050 621.600 ;
        RECT 687.150 621.000 688.950 622.800 ;
        RECT 698.100 622.200 699.150 623.100 ;
        RECT 694.350 621.450 696.150 622.200 ;
        RECT 679.950 619.500 683.700 620.700 ;
        RECT 682.650 618.600 683.700 619.500 ;
        RECT 691.200 620.400 696.150 621.450 ;
        RECT 697.650 620.400 699.450 622.200 ;
        RECT 706.950 621.600 707.850 634.200 ;
        RECT 691.200 618.600 692.250 620.400 ;
        RECT 700.950 619.500 703.050 621.600 ;
        RECT 700.950 618.600 702.000 619.500 ;
        RECT 677.850 615.750 679.650 618.600 ;
        RECT 682.350 615.750 684.150 618.600 ;
        RECT 686.550 615.750 688.350 618.600 ;
        RECT 690.450 615.750 692.250 618.600 ;
        RECT 693.750 615.750 695.550 618.600 ;
        RECT 698.250 617.700 702.000 618.600 ;
        RECT 698.250 615.750 700.050 617.700 ;
        RECT 703.050 615.750 704.850 618.600 ;
        RECT 706.050 615.750 707.850 621.600 ;
        RECT 5.850 604.200 7.650 611.250 ;
        RECT 10.350 605.400 12.150 611.250 ;
        RECT 14.850 605.400 16.650 611.250 ;
        RECT 19.350 604.200 21.150 611.250 ;
        RECT 5.850 603.300 9.450 604.200 ;
        RECT 5.100 597.150 6.900 598.950 ;
        RECT 4.950 595.050 7.050 597.150 ;
        RECT 8.250 595.950 9.450 603.300 ;
        RECT 17.550 603.300 21.150 604.200 ;
        RECT 29.850 604.200 31.650 611.250 ;
        RECT 34.350 605.400 36.150 611.250 ;
        RECT 40.650 605.400 42.450 611.250 ;
        RECT 29.850 603.300 33.450 604.200 ;
        RECT 11.100 597.150 12.900 598.950 ;
        RECT 14.100 597.150 15.900 598.950 ;
        RECT 7.950 593.850 10.050 595.950 ;
        RECT 10.950 595.050 13.050 597.150 ;
        RECT 13.950 595.050 16.050 597.150 ;
        RECT 17.550 595.950 18.750 603.300 ;
        RECT 20.100 597.150 21.900 598.950 ;
        RECT 29.100 597.150 30.900 598.950 ;
        RECT 16.950 593.850 19.050 595.950 ;
        RECT 19.950 595.050 22.050 597.150 ;
        RECT 28.950 595.050 31.050 597.150 ;
        RECT 32.250 595.950 33.450 603.300 ;
        RECT 41.250 603.300 42.450 605.400 ;
        RECT 43.650 606.300 45.450 611.250 ;
        RECT 46.650 607.200 48.450 611.250 ;
        RECT 49.650 606.300 51.450 611.250 ;
        RECT 43.650 604.950 51.450 606.300 ;
        RECT 54.000 605.400 55.800 611.250 ;
        RECT 58.200 607.050 60.000 611.250 ;
        RECT 61.500 608.400 63.300 611.250 ;
        RECT 70.650 608.400 72.450 611.250 ;
        RECT 73.650 608.400 75.450 611.250 ;
        RECT 76.650 608.400 78.450 611.250 ;
        RECT 58.200 605.400 63.900 607.050 ;
        RECT 41.250 602.250 45.000 603.300 ;
        RECT 43.950 598.950 45.150 602.250 ;
        RECT 47.100 600.150 48.900 601.950 ;
        RECT 53.100 600.150 54.900 601.950 ;
        RECT 35.100 597.150 36.900 598.950 ;
        RECT 31.950 593.850 34.050 595.950 ;
        RECT 34.950 595.050 37.050 597.150 ;
        RECT 43.950 596.850 46.050 598.950 ;
        RECT 46.950 598.050 49.050 600.150 ;
        RECT 49.950 596.850 52.050 598.950 ;
        RECT 52.950 598.050 55.050 600.150 ;
        RECT 55.950 599.850 58.050 601.950 ;
        RECT 59.100 600.150 60.900 601.950 ;
        RECT 56.100 598.050 57.900 599.850 ;
        RECT 58.950 598.050 61.050 600.150 ;
        RECT 62.700 598.950 63.900 605.400 ;
        RECT 73.950 601.950 75.000 608.400 ;
        RECT 80.850 605.400 82.650 611.250 ;
        RECT 85.350 604.200 87.150 611.250 ;
        RECT 92.550 606.300 94.350 611.250 ;
        RECT 95.550 607.200 97.350 611.250 ;
        RECT 98.550 606.300 100.350 611.250 ;
        RECT 92.550 604.950 100.350 606.300 ;
        RECT 101.550 605.400 103.350 611.250 ;
        RECT 83.550 603.300 87.150 604.200 ;
        RECT 101.550 603.300 102.750 605.400 ;
        RECT 73.950 599.850 76.050 601.950 ;
        RECT 61.950 596.850 64.050 598.950 ;
        RECT 70.950 596.850 73.050 598.950 ;
        RECT 40.950 593.850 43.050 595.950 ;
        RECT 8.250 585.600 9.450 593.850 ;
        RECT 17.550 585.600 18.750 593.850 ;
        RECT 32.250 585.600 33.450 593.850 ;
        RECT 41.250 592.050 43.050 593.850 ;
        RECT 44.850 591.600 46.050 596.850 ;
        RECT 50.100 595.050 51.900 596.850 ;
        RECT 62.700 591.600 63.900 596.850 ;
        RECT 71.100 595.050 72.900 596.850 ;
        RECT 73.950 592.650 75.000 599.850 ;
        RECT 76.950 596.850 79.050 598.950 ;
        RECT 80.100 597.150 81.900 598.950 ;
        RECT 77.100 595.050 78.900 596.850 ;
        RECT 79.950 595.050 82.050 597.150 ;
        RECT 83.550 595.950 84.750 603.300 ;
        RECT 99.000 602.250 102.750 603.300 ;
        RECT 113.100 603.000 114.900 611.250 ;
        RECT 95.100 600.150 96.900 601.950 ;
        RECT 86.100 597.150 87.900 598.950 ;
        RECT 82.950 593.850 85.050 595.950 ;
        RECT 85.950 595.050 88.050 597.150 ;
        RECT 91.950 596.850 94.050 598.950 ;
        RECT 94.950 598.050 97.050 600.150 ;
        RECT 98.850 598.950 100.050 602.250 ;
        RECT 97.950 596.850 100.050 598.950 ;
        RECT 110.400 601.350 114.900 603.000 ;
        RECT 118.500 602.400 120.300 611.250 ;
        RECT 122.700 602.400 124.500 611.250 ;
        RECT 128.100 603.000 129.900 611.250 ;
        RECT 139.650 605.400 141.450 611.250 ;
        RECT 140.250 603.300 141.450 605.400 ;
        RECT 142.650 606.300 144.450 611.250 ;
        RECT 145.650 607.200 147.450 611.250 ;
        RECT 148.650 606.300 150.450 611.250 ;
        RECT 142.650 604.950 150.450 606.300 ;
        RECT 152.550 606.300 154.350 611.250 ;
        RECT 155.550 607.200 157.350 611.250 ;
        RECT 158.550 606.300 160.350 611.250 ;
        RECT 152.550 604.950 160.350 606.300 ;
        RECT 161.550 605.400 163.350 611.250 ;
        RECT 169.650 608.400 171.450 611.250 ;
        RECT 172.650 608.400 174.450 611.250 ;
        RECT 161.550 603.300 162.750 605.400 ;
        RECT 128.100 601.350 132.600 603.000 ;
        RECT 140.250 602.250 144.000 603.300 ;
        RECT 159.000 602.250 162.750 603.300 ;
        RECT 110.400 597.150 111.600 601.350 ;
        RECT 131.400 597.150 132.600 601.350 ;
        RECT 142.950 598.950 144.150 602.250 ;
        RECT 146.100 600.150 147.900 601.950 ;
        RECT 155.100 600.150 156.900 601.950 ;
        RECT 92.100 595.050 93.900 596.850 ;
        RECT 72.450 591.600 75.000 592.650 ;
        RECT 4.650 579.750 6.450 585.600 ;
        RECT 7.650 579.750 9.450 585.600 ;
        RECT 10.650 579.750 12.450 585.600 ;
        RECT 14.550 579.750 16.350 585.600 ;
        RECT 17.550 579.750 19.350 585.600 ;
        RECT 20.550 579.750 22.350 585.600 ;
        RECT 28.650 579.750 30.450 585.600 ;
        RECT 31.650 579.750 33.450 585.600 ;
        RECT 34.650 579.750 36.450 585.600 ;
        RECT 41.400 579.750 43.200 585.600 ;
        RECT 44.700 579.750 46.500 591.600 ;
        RECT 48.900 579.750 50.700 591.600 ;
        RECT 53.550 590.700 61.350 591.600 ;
        RECT 53.550 579.750 55.350 590.700 ;
        RECT 56.550 579.750 58.350 589.800 ;
        RECT 59.550 579.750 61.350 590.700 ;
        RECT 62.550 579.750 64.350 591.600 ;
        RECT 72.450 579.750 74.250 591.600 ;
        RECT 76.650 579.750 78.450 591.600 ;
        RECT 83.550 585.600 84.750 593.850 ;
        RECT 97.950 591.600 99.150 596.850 ;
        RECT 100.950 593.850 103.050 595.950 ;
        RECT 109.950 595.050 112.050 597.150 ;
        RECT 100.950 592.050 102.750 593.850 ;
        RECT 80.550 579.750 82.350 585.600 ;
        RECT 83.550 579.750 85.350 585.600 ;
        RECT 86.550 579.750 88.350 585.600 ;
        RECT 93.300 579.750 95.100 591.600 ;
        RECT 97.500 579.750 99.300 591.600 ;
        RECT 110.250 586.800 111.300 595.050 ;
        RECT 112.950 593.850 115.050 595.950 ;
        RECT 118.950 593.850 121.050 595.950 ;
        RECT 121.950 593.850 124.050 595.950 ;
        RECT 127.950 593.850 130.050 595.950 ;
        RECT 130.950 595.050 133.050 597.150 ;
        RECT 142.950 596.850 145.050 598.950 ;
        RECT 145.950 598.050 148.050 600.150 ;
        RECT 148.950 596.850 151.050 598.950 ;
        RECT 151.950 596.850 154.050 598.950 ;
        RECT 154.950 598.050 157.050 600.150 ;
        RECT 158.850 598.950 160.050 602.250 ;
        RECT 170.400 600.150 171.600 608.400 ;
        RECT 182.100 603.000 183.900 611.250 ;
        RECT 157.950 596.850 160.050 598.950 ;
        RECT 169.950 598.050 172.050 600.150 ;
        RECT 172.950 599.850 175.050 601.950 ;
        RECT 179.400 601.350 183.900 603.000 ;
        RECT 187.500 602.400 189.300 611.250 ;
        RECT 191.550 608.400 193.350 611.250 ;
        RECT 194.550 608.400 196.350 611.250 ;
        RECT 173.100 598.050 174.900 599.850 ;
        RECT 112.950 592.050 114.750 593.850 ;
        RECT 115.950 590.850 118.050 592.950 ;
        RECT 119.100 592.050 120.900 593.850 ;
        RECT 122.100 592.050 123.900 593.850 ;
        RECT 124.950 590.850 127.050 592.950 ;
        RECT 128.250 592.050 130.050 593.850 ;
        RECT 116.100 589.050 117.900 590.850 ;
        RECT 125.100 589.050 126.900 590.850 ;
        RECT 131.700 586.800 132.750 595.050 ;
        RECT 139.950 593.850 142.050 595.950 ;
        RECT 140.250 592.050 142.050 593.850 ;
        RECT 143.850 591.600 145.050 596.850 ;
        RECT 149.100 595.050 150.900 596.850 ;
        RECT 152.100 595.050 153.900 596.850 ;
        RECT 157.950 591.600 159.150 596.850 ;
        RECT 160.950 593.850 163.050 595.950 ;
        RECT 160.950 592.050 162.750 593.850 ;
        RECT 110.250 585.900 117.300 586.800 ;
        RECT 110.250 585.600 111.450 585.900 ;
        RECT 100.800 579.750 102.600 585.600 ;
        RECT 109.650 579.750 111.450 585.600 ;
        RECT 115.650 585.600 117.300 585.900 ;
        RECT 125.700 585.900 132.750 586.800 ;
        RECT 125.700 585.600 127.350 585.900 ;
        RECT 112.650 579.750 114.450 585.000 ;
        RECT 115.650 579.750 117.450 585.600 ;
        RECT 118.650 579.750 120.450 585.600 ;
        RECT 122.550 579.750 124.350 585.600 ;
        RECT 125.550 579.750 127.350 585.600 ;
        RECT 131.550 585.600 132.750 585.900 ;
        RECT 128.550 579.750 130.350 585.000 ;
        RECT 131.550 579.750 133.350 585.600 ;
        RECT 140.400 579.750 142.200 585.600 ;
        RECT 143.700 579.750 145.500 591.600 ;
        RECT 147.900 579.750 149.700 591.600 ;
        RECT 153.300 579.750 155.100 591.600 ;
        RECT 157.500 579.750 159.300 591.600 ;
        RECT 170.400 585.600 171.600 598.050 ;
        RECT 179.400 597.150 180.600 601.350 ;
        RECT 190.950 599.850 193.050 601.950 ;
        RECT 194.400 600.150 195.600 608.400 ;
        RECT 200.700 602.400 202.500 611.250 ;
        RECT 206.100 603.000 207.900 611.250 ;
        RECT 206.100 601.350 210.600 603.000 ;
        RECT 215.700 602.400 217.500 611.250 ;
        RECT 221.100 603.000 222.900 611.250 ;
        RECT 230.850 605.400 232.650 611.250 ;
        RECT 235.350 604.200 237.150 611.250 ;
        RECT 244.650 608.400 246.450 611.250 ;
        RECT 247.650 608.400 249.450 611.250 ;
        RECT 250.650 608.400 252.450 611.250 ;
        RECT 233.550 603.300 237.150 604.200 ;
        RECT 221.100 601.350 225.600 603.000 ;
        RECT 191.100 598.050 192.900 599.850 ;
        RECT 193.950 598.050 196.050 600.150 ;
        RECT 178.950 595.050 181.050 597.150 ;
        RECT 179.250 586.800 180.300 595.050 ;
        RECT 181.950 593.850 184.050 595.950 ;
        RECT 187.950 593.850 190.050 595.950 ;
        RECT 181.950 592.050 183.750 593.850 ;
        RECT 184.950 590.850 187.050 592.950 ;
        RECT 188.100 592.050 189.900 593.850 ;
        RECT 185.100 589.050 186.900 590.850 ;
        RECT 179.250 585.900 186.300 586.800 ;
        RECT 179.250 585.600 180.450 585.900 ;
        RECT 160.800 579.750 162.600 585.600 ;
        RECT 169.650 579.750 171.450 585.600 ;
        RECT 172.650 579.750 174.450 585.600 ;
        RECT 178.650 579.750 180.450 585.600 ;
        RECT 184.650 585.600 186.300 585.900 ;
        RECT 194.400 585.600 195.600 598.050 ;
        RECT 209.400 597.150 210.600 601.350 ;
        RECT 224.400 597.150 225.600 601.350 ;
        RECT 230.100 597.150 231.900 598.950 ;
        RECT 199.950 593.850 202.050 595.950 ;
        RECT 205.950 593.850 208.050 595.950 ;
        RECT 208.950 595.050 211.050 597.150 ;
        RECT 200.100 592.050 201.900 593.850 ;
        RECT 202.950 590.850 205.050 592.950 ;
        RECT 206.250 592.050 208.050 593.850 ;
        RECT 203.100 589.050 204.900 590.850 ;
        RECT 209.700 586.800 210.750 595.050 ;
        RECT 214.950 593.850 217.050 595.950 ;
        RECT 220.950 593.850 223.050 595.950 ;
        RECT 223.950 595.050 226.050 597.150 ;
        RECT 229.950 595.050 232.050 597.150 ;
        RECT 233.550 595.950 234.750 603.300 ;
        RECT 247.950 601.950 249.000 608.400 ;
        RECT 258.150 606.900 259.950 611.250 ;
        RECT 256.650 605.400 259.950 606.900 ;
        RECT 261.150 605.400 262.950 611.250 ;
        RECT 247.950 599.850 250.050 601.950 ;
        RECT 236.100 597.150 237.900 598.950 ;
        RECT 215.100 592.050 216.900 593.850 ;
        RECT 217.950 590.850 220.050 592.950 ;
        RECT 221.250 592.050 223.050 593.850 ;
        RECT 218.100 589.050 219.900 590.850 ;
        RECT 224.700 586.800 225.750 595.050 ;
        RECT 232.950 593.850 235.050 595.950 ;
        RECT 235.950 595.050 238.050 597.150 ;
        RECT 244.950 596.850 247.050 598.950 ;
        RECT 245.100 595.050 246.900 596.850 ;
        RECT 203.700 585.900 210.750 586.800 ;
        RECT 203.700 585.600 205.350 585.900 ;
        RECT 181.650 579.750 183.450 585.000 ;
        RECT 184.650 579.750 186.450 585.600 ;
        RECT 187.650 579.750 189.450 585.600 ;
        RECT 191.550 579.750 193.350 585.600 ;
        RECT 194.550 579.750 196.350 585.600 ;
        RECT 200.550 579.750 202.350 585.600 ;
        RECT 203.550 579.750 205.350 585.600 ;
        RECT 209.550 585.600 210.750 585.900 ;
        RECT 218.700 585.900 225.750 586.800 ;
        RECT 218.700 585.600 220.350 585.900 ;
        RECT 206.550 579.750 208.350 585.000 ;
        RECT 209.550 579.750 211.350 585.600 ;
        RECT 215.550 579.750 217.350 585.600 ;
        RECT 218.550 579.750 220.350 585.600 ;
        RECT 224.550 585.600 225.750 585.900 ;
        RECT 233.550 585.600 234.750 593.850 ;
        RECT 247.950 592.650 249.000 599.850 ;
        RECT 256.650 598.950 257.850 605.400 ;
        RECT 259.950 603.900 261.750 604.500 ;
        RECT 265.650 603.900 267.450 611.250 ;
        RECT 271.650 605.400 273.450 611.250 ;
        RECT 259.950 602.700 267.450 603.900 ;
        RECT 272.250 603.300 273.450 605.400 ;
        RECT 274.650 606.300 276.450 611.250 ;
        RECT 277.650 607.200 279.450 611.250 ;
        RECT 280.650 606.300 282.450 611.250 ;
        RECT 284.550 608.400 286.350 611.250 ;
        RECT 287.550 608.400 289.350 611.250 ;
        RECT 290.550 608.400 292.350 611.250 ;
        RECT 298.650 608.400 300.450 611.250 ;
        RECT 301.650 608.400 303.450 611.250 ;
        RECT 274.650 604.950 282.450 606.300 ;
        RECT 250.950 596.850 253.050 598.950 ;
        RECT 256.650 596.850 259.050 598.950 ;
        RECT 260.100 597.150 261.900 598.950 ;
        RECT 251.100 595.050 252.900 596.850 ;
        RECT 246.450 591.600 249.000 592.650 ;
        RECT 256.650 591.600 257.850 596.850 ;
        RECT 259.950 595.050 262.050 597.150 ;
        RECT 221.550 579.750 223.350 585.000 ;
        RECT 224.550 579.750 226.350 585.600 ;
        RECT 230.550 579.750 232.350 585.600 ;
        RECT 233.550 579.750 235.350 585.600 ;
        RECT 236.550 579.750 238.350 585.600 ;
        RECT 246.450 579.750 248.250 591.600 ;
        RECT 250.650 579.750 252.450 591.600 ;
        RECT 256.050 579.750 257.850 591.600 ;
        RECT 259.050 579.750 260.850 591.600 ;
        RECT 263.100 585.600 264.300 602.700 ;
        RECT 272.250 602.250 276.000 603.300 ;
        RECT 274.950 598.950 276.150 602.250 ;
        RECT 288.000 601.950 289.050 608.400 ;
        RECT 278.100 600.150 279.900 601.950 ;
        RECT 265.950 596.850 268.050 598.950 ;
        RECT 274.950 596.850 277.050 598.950 ;
        RECT 277.950 598.050 280.050 600.150 ;
        RECT 286.950 599.850 289.050 601.950 ;
        RECT 299.400 600.150 300.600 608.400 ;
        RECT 305.550 606.300 307.350 611.250 ;
        RECT 308.550 607.200 310.350 611.250 ;
        RECT 311.550 606.300 313.350 611.250 ;
        RECT 305.550 604.950 313.350 606.300 ;
        RECT 314.550 605.400 316.350 611.250 ;
        RECT 320.550 608.400 322.350 611.250 ;
        RECT 323.550 608.400 325.350 611.250 ;
        RECT 314.550 603.300 315.750 605.400 ;
        RECT 312.000 602.250 315.750 603.300 ;
        RECT 280.950 596.850 283.050 598.950 ;
        RECT 283.950 596.850 286.050 598.950 ;
        RECT 266.100 595.050 267.900 596.850 ;
        RECT 271.950 593.850 274.050 595.950 ;
        RECT 272.250 592.050 274.050 593.850 ;
        RECT 275.850 591.600 277.050 596.850 ;
        RECT 281.100 595.050 282.900 596.850 ;
        RECT 284.100 595.050 285.900 596.850 ;
        RECT 288.000 592.650 289.050 599.850 ;
        RECT 289.950 596.850 292.050 598.950 ;
        RECT 298.950 598.050 301.050 600.150 ;
        RECT 301.950 599.850 304.050 601.950 ;
        RECT 308.100 600.150 309.900 601.950 ;
        RECT 302.100 598.050 303.900 599.850 ;
        RECT 290.100 595.050 291.900 596.850 ;
        RECT 288.000 591.600 290.550 592.650 ;
        RECT 262.650 579.750 264.450 585.600 ;
        RECT 265.650 579.750 267.450 585.600 ;
        RECT 272.400 579.750 274.200 585.600 ;
        RECT 275.700 579.750 277.500 591.600 ;
        RECT 279.900 579.750 281.700 591.600 ;
        RECT 284.550 579.750 286.350 591.600 ;
        RECT 288.750 579.750 290.550 591.600 ;
        RECT 299.400 585.600 300.600 598.050 ;
        RECT 304.950 596.850 307.050 598.950 ;
        RECT 307.950 598.050 310.050 600.150 ;
        RECT 311.850 598.950 313.050 602.250 ;
        RECT 319.950 599.850 322.050 601.950 ;
        RECT 323.400 600.150 324.600 608.400 ;
        RECT 329.850 605.400 331.650 611.250 ;
        RECT 334.350 604.200 336.150 611.250 ;
        RECT 332.550 603.300 336.150 604.200 ;
        RECT 310.950 596.850 313.050 598.950 ;
        RECT 320.100 598.050 321.900 599.850 ;
        RECT 322.950 598.050 325.050 600.150 ;
        RECT 305.100 595.050 306.900 596.850 ;
        RECT 310.950 591.600 312.150 596.850 ;
        RECT 313.950 593.850 316.050 595.950 ;
        RECT 313.950 592.050 315.750 593.850 ;
        RECT 298.650 579.750 300.450 585.600 ;
        RECT 301.650 579.750 303.450 585.600 ;
        RECT 306.300 579.750 308.100 591.600 ;
        RECT 310.500 579.750 312.300 591.600 ;
        RECT 323.400 585.600 324.600 598.050 ;
        RECT 329.100 597.150 330.900 598.950 ;
        RECT 328.950 595.050 331.050 597.150 ;
        RECT 332.550 595.950 333.750 603.300 ;
        RECT 341.700 602.400 343.500 611.250 ;
        RECT 347.100 603.000 348.900 611.250 ;
        RECT 356.550 608.400 358.350 611.250 ;
        RECT 357.150 604.500 358.350 608.400 ;
        RECT 359.850 605.400 361.650 611.250 ;
        RECT 362.850 605.400 364.650 611.250 ;
        RECT 368.550 605.400 370.350 611.250 ;
        RECT 371.550 605.400 373.350 611.250 ;
        RECT 374.550 605.400 376.350 611.250 ;
        RECT 357.150 603.600 362.250 604.500 ;
        RECT 347.100 601.350 351.600 603.000 ;
        RECT 335.100 597.150 336.900 598.950 ;
        RECT 350.400 597.150 351.600 601.350 ;
        RECT 360.000 602.700 362.250 603.600 ;
        RECT 331.950 593.850 334.050 595.950 ;
        RECT 334.950 595.050 337.050 597.150 ;
        RECT 340.950 593.850 343.050 595.950 ;
        RECT 346.950 593.850 349.050 595.950 ;
        RECT 349.950 595.050 352.050 597.150 ;
        RECT 355.950 596.850 358.050 598.950 ;
        RECT 356.100 595.050 357.900 596.850 ;
        RECT 332.550 585.600 333.750 593.850 ;
        RECT 341.100 592.050 342.900 593.850 ;
        RECT 343.950 590.850 346.050 592.950 ;
        RECT 347.250 592.050 349.050 593.850 ;
        RECT 344.100 589.050 345.900 590.850 ;
        RECT 350.700 586.800 351.750 595.050 ;
        RECT 360.000 594.300 361.050 602.700 ;
        RECT 363.150 598.950 364.350 605.400 ;
        RECT 371.400 604.500 373.200 605.400 ;
        RECT 377.550 604.500 379.350 611.250 ;
        RECT 380.550 605.400 382.350 611.250 ;
        RECT 383.550 605.400 385.350 611.250 ;
        RECT 386.550 605.400 388.350 611.250 ;
        RECT 389.550 605.400 391.350 611.250 ;
        RECT 392.550 605.400 394.350 611.250 ;
        RECT 399.150 605.400 400.950 611.250 ;
        RECT 402.150 608.400 403.950 611.250 ;
        RECT 406.950 609.300 408.750 611.250 ;
        RECT 405.000 608.400 408.750 609.300 ;
        RECT 411.450 608.400 413.250 611.250 ;
        RECT 414.750 608.400 416.550 611.250 ;
        RECT 418.650 608.400 420.450 611.250 ;
        RECT 422.850 608.400 424.650 611.250 ;
        RECT 427.350 608.400 429.150 611.250 ;
        RECT 405.000 607.500 406.050 608.400 ;
        RECT 403.950 605.400 406.050 607.500 ;
        RECT 414.750 606.600 415.800 608.400 ;
        RECT 383.400 604.500 385.200 605.400 ;
        RECT 389.400 604.500 391.200 605.400 ;
        RECT 371.400 603.300 375.450 604.500 ;
        RECT 377.550 603.300 381.300 604.500 ;
        RECT 383.400 603.300 387.300 604.500 ;
        RECT 389.400 604.350 392.100 604.500 ;
        RECT 389.400 603.300 392.250 604.350 ;
        RECT 374.250 602.400 375.450 603.300 ;
        RECT 380.100 602.400 381.300 603.300 ;
        RECT 386.100 602.400 387.300 603.300 ;
        RECT 371.100 600.150 372.900 601.950 ;
        RECT 374.250 600.600 378.300 602.400 ;
        RECT 380.100 600.600 384.300 602.400 ;
        RECT 386.100 600.600 390.300 602.400 ;
        RECT 361.950 596.850 364.350 598.950 ;
        RECT 370.950 598.050 373.050 600.150 ;
        RECT 360.000 593.400 362.250 594.300 ;
        RECT 344.700 585.900 351.750 586.800 ;
        RECT 344.700 585.600 346.350 585.900 ;
        RECT 313.800 579.750 315.600 585.600 ;
        RECT 320.550 579.750 322.350 585.600 ;
        RECT 323.550 579.750 325.350 585.600 ;
        RECT 329.550 579.750 331.350 585.600 ;
        RECT 332.550 579.750 334.350 585.600 ;
        RECT 335.550 579.750 337.350 585.600 ;
        RECT 341.550 579.750 343.350 585.600 ;
        RECT 344.550 579.750 346.350 585.600 ;
        RECT 350.550 585.600 351.750 585.900 ;
        RECT 356.550 592.500 362.250 593.400 ;
        RECT 356.550 585.600 357.750 592.500 ;
        RECT 363.150 591.600 364.350 596.850 ;
        RECT 374.250 593.700 375.450 600.600 ;
        RECT 380.100 593.700 381.300 600.600 ;
        RECT 386.100 593.700 387.300 600.600 ;
        RECT 391.200 600.150 392.250 603.300 ;
        RECT 391.200 598.050 394.050 600.150 ;
        RECT 391.200 593.700 392.250 598.050 ;
        RECT 371.550 592.500 375.450 593.700 ;
        RECT 377.550 592.500 381.300 593.700 ;
        RECT 383.550 592.500 387.300 593.700 ;
        RECT 389.550 592.500 392.250 593.700 ;
        RECT 399.150 592.800 400.050 605.400 ;
        RECT 407.550 604.800 409.350 606.600 ;
        RECT 410.850 605.550 415.800 606.600 ;
        RECT 423.300 607.500 424.350 608.400 ;
        RECT 423.300 606.300 427.050 607.500 ;
        RECT 410.850 604.800 412.650 605.550 ;
        RECT 407.850 603.900 408.900 604.800 ;
        RECT 418.050 604.200 419.850 606.000 ;
        RECT 424.950 605.400 427.050 606.300 ;
        RECT 430.650 605.400 432.450 611.250 ;
        RECT 434.550 608.400 436.350 611.250 ;
        RECT 437.550 608.400 439.350 611.250 ;
        RECT 418.050 603.900 418.950 604.200 ;
        RECT 407.850 603.000 418.950 603.900 ;
        RECT 431.250 603.150 432.450 605.400 ;
        RECT 407.850 601.800 408.900 603.000 ;
        RECT 402.000 600.600 408.900 601.800 ;
        RECT 402.000 599.850 402.900 600.600 ;
        RECT 407.100 600.000 408.900 600.600 ;
        RECT 401.100 598.050 402.900 599.850 ;
        RECT 404.100 598.950 405.900 599.700 ;
        RECT 418.050 598.950 418.950 603.000 ;
        RECT 427.950 601.050 432.450 603.150 ;
        RECT 426.150 599.250 430.050 601.050 ;
        RECT 427.950 598.950 430.050 599.250 ;
        RECT 404.100 597.900 412.050 598.950 ;
        RECT 409.950 596.850 412.050 597.900 ;
        RECT 415.950 596.850 418.950 598.950 ;
        RECT 408.450 593.100 410.250 593.400 ;
        RECT 408.450 592.800 416.850 593.100 ;
        RECT 347.550 579.750 349.350 585.000 ;
        RECT 350.550 579.750 352.350 585.600 ;
        RECT 356.550 579.750 358.350 585.600 ;
        RECT 359.850 579.750 361.650 591.600 ;
        RECT 362.850 579.750 364.650 591.600 ;
        RECT 368.550 579.750 370.350 591.600 ;
        RECT 371.550 579.750 373.350 592.500 ;
        RECT 374.550 579.750 376.350 591.600 ;
        RECT 377.550 579.750 379.350 592.500 ;
        RECT 380.550 579.750 382.350 591.600 ;
        RECT 383.550 579.750 385.350 592.500 ;
        RECT 386.550 579.750 388.350 591.600 ;
        RECT 389.550 579.750 391.350 592.500 ;
        RECT 399.150 592.200 416.850 592.800 ;
        RECT 399.150 591.600 410.250 592.200 ;
        RECT 392.550 579.750 394.350 591.600 ;
        RECT 399.150 579.750 400.950 591.600 ;
        RECT 413.250 590.700 415.050 591.300 ;
        RECT 407.550 589.500 415.050 590.700 ;
        RECT 415.950 590.100 416.850 592.200 ;
        RECT 418.050 592.200 418.950 596.850 ;
        RECT 428.250 593.400 430.050 595.200 ;
        RECT 424.950 592.200 429.150 593.400 ;
        RECT 418.050 591.300 424.050 592.200 ;
        RECT 424.950 591.300 427.050 592.200 ;
        RECT 431.250 591.600 432.450 601.050 ;
        RECT 433.950 599.850 436.050 601.950 ;
        RECT 437.400 600.150 438.600 608.400 ;
        RECT 443.550 606.300 445.350 611.250 ;
        RECT 446.550 607.200 448.350 611.250 ;
        RECT 449.550 606.300 451.350 611.250 ;
        RECT 443.550 604.950 451.350 606.300 ;
        RECT 452.550 605.400 454.350 611.250 ;
        RECT 458.550 608.400 460.350 611.250 ;
        RECT 461.550 608.400 463.350 611.250 ;
        RECT 464.550 608.400 466.350 611.250 ;
        RECT 452.550 603.300 453.750 605.400 ;
        RECT 450.000 602.250 453.750 603.300 ;
        RECT 446.100 600.150 447.900 601.950 ;
        RECT 434.100 598.050 435.900 599.850 ;
        RECT 436.950 598.050 439.050 600.150 ;
        RECT 423.150 590.400 424.050 591.300 ;
        RECT 420.450 590.100 422.250 590.400 ;
        RECT 407.550 588.600 408.750 589.500 ;
        RECT 415.950 589.200 422.250 590.100 ;
        RECT 420.450 588.600 422.250 589.200 ;
        RECT 423.150 588.600 425.850 590.400 ;
        RECT 403.950 586.500 408.750 588.600 ;
        RECT 411.150 586.500 418.050 588.300 ;
        RECT 407.550 585.600 408.750 586.500 ;
        RECT 402.150 579.750 403.950 585.600 ;
        RECT 407.250 579.750 409.050 585.600 ;
        RECT 412.050 579.750 413.850 585.600 ;
        RECT 415.050 579.750 416.850 586.500 ;
        RECT 423.150 585.600 427.050 587.700 ;
        RECT 418.950 579.750 420.750 585.600 ;
        RECT 423.150 579.750 424.950 585.600 ;
        RECT 427.650 579.750 429.450 582.600 ;
        RECT 430.650 579.750 432.450 591.600 ;
        RECT 437.400 585.600 438.600 598.050 ;
        RECT 442.950 596.850 445.050 598.950 ;
        RECT 445.950 598.050 448.050 600.150 ;
        RECT 449.850 598.950 451.050 602.250 ;
        RECT 462.000 601.950 463.050 608.400 ;
        RECT 470.850 605.400 472.650 611.250 ;
        RECT 475.350 604.200 477.150 611.250 ;
        RECT 485.700 608.400 487.500 611.250 ;
        RECT 489.000 607.050 490.800 611.250 ;
        RECT 460.950 599.850 463.050 601.950 ;
        RECT 448.950 596.850 451.050 598.950 ;
        RECT 457.950 596.850 460.050 598.950 ;
        RECT 443.100 595.050 444.900 596.850 ;
        RECT 448.950 591.600 450.150 596.850 ;
        RECT 451.950 593.850 454.050 595.950 ;
        RECT 458.100 595.050 459.900 596.850 ;
        RECT 451.950 592.050 453.750 593.850 ;
        RECT 462.000 592.650 463.050 599.850 ;
        RECT 473.550 603.300 477.150 604.200 ;
        RECT 485.100 605.400 490.800 607.050 ;
        RECT 493.200 605.400 495.000 611.250 ;
        RECT 463.950 596.850 466.050 598.950 ;
        RECT 470.100 597.150 471.900 598.950 ;
        RECT 464.100 595.050 465.900 596.850 ;
        RECT 469.950 595.050 472.050 597.150 ;
        RECT 473.550 595.950 474.750 603.300 ;
        RECT 485.100 598.950 486.300 605.400 ;
        RECT 497.550 603.900 499.350 611.250 ;
        RECT 502.050 605.400 503.850 611.250 ;
        RECT 505.050 606.900 506.850 611.250 ;
        RECT 514.650 608.400 516.450 611.250 ;
        RECT 517.650 608.400 519.450 611.250 ;
        RECT 520.650 608.400 522.450 611.250 ;
        RECT 526.650 608.400 528.450 611.250 ;
        RECT 529.650 608.400 531.450 611.250 ;
        RECT 505.050 605.400 508.350 606.900 ;
        RECT 503.250 603.900 505.050 604.500 ;
        RECT 497.550 602.700 505.050 603.900 ;
        RECT 488.100 600.150 489.900 601.950 ;
        RECT 476.100 597.150 477.900 598.950 ;
        RECT 472.950 593.850 475.050 595.950 ;
        RECT 475.950 595.050 478.050 597.150 ;
        RECT 484.950 596.850 487.050 598.950 ;
        RECT 487.950 598.050 490.050 600.150 ;
        RECT 490.950 599.850 493.050 601.950 ;
        RECT 494.100 600.150 495.900 601.950 ;
        RECT 491.100 598.050 492.900 599.850 ;
        RECT 493.950 598.050 496.050 600.150 ;
        RECT 496.950 596.850 499.050 598.950 ;
        RECT 462.000 591.600 464.550 592.650 ;
        RECT 434.550 579.750 436.350 585.600 ;
        RECT 437.550 579.750 439.350 585.600 ;
        RECT 444.300 579.750 446.100 591.600 ;
        RECT 448.500 579.750 450.300 591.600 ;
        RECT 451.800 579.750 453.600 585.600 ;
        RECT 458.550 579.750 460.350 591.600 ;
        RECT 462.750 579.750 464.550 591.600 ;
        RECT 473.550 585.600 474.750 593.850 ;
        RECT 485.100 591.600 486.300 596.850 ;
        RECT 497.100 595.050 498.900 596.850 ;
        RECT 470.550 579.750 472.350 585.600 ;
        RECT 473.550 579.750 475.350 585.600 ;
        RECT 476.550 579.750 478.350 585.600 ;
        RECT 484.650 579.750 486.450 591.600 ;
        RECT 487.650 590.700 495.450 591.600 ;
        RECT 487.650 579.750 489.450 590.700 ;
        RECT 490.650 579.750 492.450 589.800 ;
        RECT 493.650 579.750 495.450 590.700 ;
        RECT 500.700 585.600 501.900 602.700 ;
        RECT 507.150 598.950 508.350 605.400 ;
        RECT 517.950 601.950 519.000 608.400 ;
        RECT 517.950 599.850 520.050 601.950 ;
        RECT 527.400 600.150 528.600 608.400 ;
        RECT 533.550 605.400 535.350 611.250 ;
        RECT 536.850 608.400 538.650 611.250 ;
        RECT 541.350 608.400 543.150 611.250 ;
        RECT 545.550 608.400 547.350 611.250 ;
        RECT 549.450 608.400 551.250 611.250 ;
        RECT 552.750 608.400 554.550 611.250 ;
        RECT 557.250 609.300 559.050 611.250 ;
        RECT 557.250 608.400 561.000 609.300 ;
        RECT 562.050 608.400 563.850 611.250 ;
        RECT 541.650 607.500 542.700 608.400 ;
        RECT 538.950 606.300 542.700 607.500 ;
        RECT 550.200 606.600 551.250 608.400 ;
        RECT 559.950 607.500 561.000 608.400 ;
        RECT 538.950 605.400 541.050 606.300 ;
        RECT 533.550 603.150 534.750 605.400 ;
        RECT 546.150 604.200 547.950 606.000 ;
        RECT 550.200 605.550 555.150 606.600 ;
        RECT 553.350 604.800 555.150 605.550 ;
        RECT 556.650 604.800 558.450 606.600 ;
        RECT 559.950 605.400 562.050 607.500 ;
        RECT 565.050 605.400 566.850 611.250 ;
        RECT 572.700 608.400 574.500 611.250 ;
        RECT 576.000 607.050 577.800 611.250 ;
        RECT 547.050 603.900 547.950 604.200 ;
        RECT 557.100 603.900 558.150 604.800 ;
        RECT 503.100 597.150 504.900 598.950 ;
        RECT 502.950 595.050 505.050 597.150 ;
        RECT 505.950 596.850 508.350 598.950 ;
        RECT 514.950 596.850 517.050 598.950 ;
        RECT 507.150 591.600 508.350 596.850 ;
        RECT 515.100 595.050 516.900 596.850 ;
        RECT 517.950 592.650 519.000 599.850 ;
        RECT 520.950 596.850 523.050 598.950 ;
        RECT 526.950 598.050 529.050 600.150 ;
        RECT 529.950 599.850 532.050 601.950 ;
        RECT 533.550 601.050 538.050 603.150 ;
        RECT 547.050 603.000 558.150 603.900 ;
        RECT 530.100 598.050 531.900 599.850 ;
        RECT 521.100 595.050 522.900 596.850 ;
        RECT 516.450 591.600 519.000 592.650 ;
        RECT 497.550 579.750 499.350 585.600 ;
        RECT 500.550 579.750 502.350 585.600 ;
        RECT 504.150 579.750 505.950 591.600 ;
        RECT 507.150 579.750 508.950 591.600 ;
        RECT 516.450 579.750 518.250 591.600 ;
        RECT 520.650 579.750 522.450 591.600 ;
        RECT 527.400 585.600 528.600 598.050 ;
        RECT 533.550 591.600 534.750 601.050 ;
        RECT 535.950 599.250 539.850 601.050 ;
        RECT 535.950 598.950 538.050 599.250 ;
        RECT 547.050 598.950 547.950 603.000 ;
        RECT 557.100 601.800 558.150 603.000 ;
        RECT 557.100 600.600 564.000 601.800 ;
        RECT 557.100 600.000 558.900 600.600 ;
        RECT 563.100 599.850 564.000 600.600 ;
        RECT 560.100 598.950 561.900 599.700 ;
        RECT 547.050 596.850 550.050 598.950 ;
        RECT 553.950 597.900 561.900 598.950 ;
        RECT 563.100 598.050 564.900 599.850 ;
        RECT 553.950 596.850 556.050 597.900 ;
        RECT 535.950 593.400 537.750 595.200 ;
        RECT 536.850 592.200 541.050 593.400 ;
        RECT 547.050 592.200 547.950 596.850 ;
        RECT 555.750 593.100 557.550 593.400 ;
        RECT 526.650 579.750 528.450 585.600 ;
        RECT 529.650 579.750 531.450 585.600 ;
        RECT 533.550 579.750 535.350 591.600 ;
        RECT 538.950 591.300 541.050 592.200 ;
        RECT 541.950 591.300 547.950 592.200 ;
        RECT 549.150 592.800 557.550 593.100 ;
        RECT 565.950 592.800 566.850 605.400 ;
        RECT 572.100 605.400 577.800 607.050 ;
        RECT 580.200 605.400 582.000 611.250 ;
        RECT 584.550 608.400 586.350 611.250 ;
        RECT 587.550 608.400 589.350 611.250 ;
        RECT 590.550 608.400 592.350 611.250 ;
        RECT 598.650 608.400 600.450 611.250 ;
        RECT 601.650 608.400 603.450 611.250 ;
        RECT 604.650 608.400 606.450 611.250 ;
        RECT 572.100 598.950 573.300 605.400 ;
        RECT 588.000 601.950 589.050 608.400 ;
        RECT 575.100 600.150 576.900 601.950 ;
        RECT 571.950 596.850 574.050 598.950 ;
        RECT 574.950 598.050 577.050 600.150 ;
        RECT 577.950 599.850 580.050 601.950 ;
        RECT 581.100 600.150 582.900 601.950 ;
        RECT 578.100 598.050 579.900 599.850 ;
        RECT 580.950 598.050 583.050 600.150 ;
        RECT 586.950 599.850 589.050 601.950 ;
        RECT 583.950 596.850 586.050 598.950 ;
        RECT 549.150 592.200 566.850 592.800 ;
        RECT 541.950 590.400 542.850 591.300 ;
        RECT 540.150 588.600 542.850 590.400 ;
        RECT 543.750 590.100 545.550 590.400 ;
        RECT 549.150 590.100 550.050 592.200 ;
        RECT 555.750 591.600 566.850 592.200 ;
        RECT 572.100 591.600 573.300 596.850 ;
        RECT 584.100 595.050 585.900 596.850 ;
        RECT 588.000 592.650 589.050 599.850 ;
        RECT 601.950 601.950 603.000 608.400 ;
        RECT 608.550 603.900 610.350 611.250 ;
        RECT 613.050 605.400 614.850 611.250 ;
        RECT 616.050 606.900 617.850 611.250 ;
        RECT 616.050 605.400 619.350 606.900 ;
        RECT 614.250 603.900 616.050 604.500 ;
        RECT 608.550 602.700 616.050 603.900 ;
        RECT 601.950 599.850 604.050 601.950 ;
        RECT 589.950 596.850 592.050 598.950 ;
        RECT 598.950 596.850 601.050 598.950 ;
        RECT 590.100 595.050 591.900 596.850 ;
        RECT 599.100 595.050 600.900 596.850 ;
        RECT 601.950 592.650 603.000 599.850 ;
        RECT 604.950 596.850 607.050 598.950 ;
        RECT 607.950 596.850 610.050 598.950 ;
        RECT 605.100 595.050 606.900 596.850 ;
        RECT 608.100 595.050 609.900 596.850 ;
        RECT 588.000 591.600 590.550 592.650 ;
        RECT 543.750 589.200 550.050 590.100 ;
        RECT 550.950 590.700 552.750 591.300 ;
        RECT 550.950 589.500 558.450 590.700 ;
        RECT 543.750 588.600 545.550 589.200 ;
        RECT 557.250 588.600 558.450 589.500 ;
        RECT 538.950 585.600 542.850 587.700 ;
        RECT 547.950 586.500 554.850 588.300 ;
        RECT 557.250 586.500 562.050 588.600 ;
        RECT 536.550 579.750 538.350 582.600 ;
        RECT 541.050 579.750 542.850 585.600 ;
        RECT 545.250 579.750 547.050 585.600 ;
        RECT 549.150 579.750 550.950 586.500 ;
        RECT 557.250 585.600 558.450 586.500 ;
        RECT 552.150 579.750 553.950 585.600 ;
        RECT 556.950 579.750 558.750 585.600 ;
        RECT 562.050 579.750 563.850 585.600 ;
        RECT 565.050 579.750 566.850 591.600 ;
        RECT 571.650 579.750 573.450 591.600 ;
        RECT 574.650 590.700 582.450 591.600 ;
        RECT 574.650 579.750 576.450 590.700 ;
        RECT 577.650 579.750 579.450 589.800 ;
        RECT 580.650 579.750 582.450 590.700 ;
        RECT 584.550 579.750 586.350 591.600 ;
        RECT 588.750 579.750 590.550 591.600 ;
        RECT 600.450 591.600 603.000 592.650 ;
        RECT 600.450 579.750 602.250 591.600 ;
        RECT 604.650 579.750 606.450 591.600 ;
        RECT 611.700 585.600 612.900 602.700 ;
        RECT 618.150 598.950 619.350 605.400 ;
        RECT 623.550 606.300 625.350 611.250 ;
        RECT 626.550 607.200 628.350 611.250 ;
        RECT 629.550 606.300 631.350 611.250 ;
        RECT 623.550 604.950 631.350 606.300 ;
        RECT 632.550 605.400 634.350 611.250 ;
        RECT 640.650 605.400 642.450 611.250 ;
        RECT 632.550 603.300 633.750 605.400 ;
        RECT 630.000 602.250 633.750 603.300 ;
        RECT 641.250 603.300 642.450 605.400 ;
        RECT 643.650 606.300 645.450 611.250 ;
        RECT 646.650 607.200 648.450 611.250 ;
        RECT 649.650 606.300 651.450 611.250 ;
        RECT 655.650 608.400 657.450 611.250 ;
        RECT 658.650 608.400 660.450 611.250 ;
        RECT 643.650 604.950 651.450 606.300 ;
        RECT 641.250 602.250 645.000 603.300 ;
        RECT 626.100 600.150 627.900 601.950 ;
        RECT 614.100 597.150 615.900 598.950 ;
        RECT 613.950 595.050 616.050 597.150 ;
        RECT 616.950 596.850 619.350 598.950 ;
        RECT 622.950 596.850 625.050 598.950 ;
        RECT 625.950 598.050 628.050 600.150 ;
        RECT 629.850 598.950 631.050 602.250 ;
        RECT 628.950 596.850 631.050 598.950 ;
        RECT 643.950 598.950 645.150 602.250 ;
        RECT 647.100 600.150 648.900 601.950 ;
        RECT 656.400 600.150 657.600 608.400 ;
        RECT 662.550 605.400 664.350 611.250 ;
        RECT 665.850 608.400 667.650 611.250 ;
        RECT 670.350 608.400 672.150 611.250 ;
        RECT 674.550 608.400 676.350 611.250 ;
        RECT 678.450 608.400 680.250 611.250 ;
        RECT 681.750 608.400 683.550 611.250 ;
        RECT 686.250 609.300 688.050 611.250 ;
        RECT 686.250 608.400 690.000 609.300 ;
        RECT 691.050 608.400 692.850 611.250 ;
        RECT 670.650 607.500 671.700 608.400 ;
        RECT 667.950 606.300 671.700 607.500 ;
        RECT 679.200 606.600 680.250 608.400 ;
        RECT 688.950 607.500 690.000 608.400 ;
        RECT 667.950 605.400 670.050 606.300 ;
        RECT 662.550 603.150 663.750 605.400 ;
        RECT 675.150 604.200 676.950 606.000 ;
        RECT 679.200 605.550 684.150 606.600 ;
        RECT 682.350 604.800 684.150 605.550 ;
        RECT 685.650 604.800 687.450 606.600 ;
        RECT 688.950 605.400 691.050 607.500 ;
        RECT 694.050 605.400 695.850 611.250 ;
        RECT 698.550 608.400 700.350 611.250 ;
        RECT 701.550 608.400 703.350 611.250 ;
        RECT 676.050 603.900 676.950 604.200 ;
        RECT 686.100 603.900 687.150 604.800 ;
        RECT 643.950 596.850 646.050 598.950 ;
        RECT 646.950 598.050 649.050 600.150 ;
        RECT 649.950 596.850 652.050 598.950 ;
        RECT 655.950 598.050 658.050 600.150 ;
        RECT 658.950 599.850 661.050 601.950 ;
        RECT 662.550 601.050 667.050 603.150 ;
        RECT 676.050 603.000 687.150 603.900 ;
        RECT 659.100 598.050 660.900 599.850 ;
        RECT 618.150 591.600 619.350 596.850 ;
        RECT 623.100 595.050 624.900 596.850 ;
        RECT 628.950 591.600 630.150 596.850 ;
        RECT 631.950 593.850 634.050 595.950 ;
        RECT 640.950 593.850 643.050 595.950 ;
        RECT 631.950 592.050 633.750 593.850 ;
        RECT 641.250 592.050 643.050 593.850 ;
        RECT 644.850 591.600 646.050 596.850 ;
        RECT 650.100 595.050 651.900 596.850 ;
        RECT 608.550 579.750 610.350 585.600 ;
        RECT 611.550 579.750 613.350 585.600 ;
        RECT 615.150 579.750 616.950 591.600 ;
        RECT 618.150 579.750 619.950 591.600 ;
        RECT 624.300 579.750 626.100 591.600 ;
        RECT 628.500 579.750 630.300 591.600 ;
        RECT 631.800 579.750 633.600 585.600 ;
        RECT 641.400 579.750 643.200 585.600 ;
        RECT 644.700 579.750 646.500 591.600 ;
        RECT 648.900 579.750 650.700 591.600 ;
        RECT 656.400 585.600 657.600 598.050 ;
        RECT 662.550 591.600 663.750 601.050 ;
        RECT 664.950 599.250 668.850 601.050 ;
        RECT 664.950 598.950 667.050 599.250 ;
        RECT 676.050 598.950 676.950 603.000 ;
        RECT 686.100 601.800 687.150 603.000 ;
        RECT 686.100 600.600 693.000 601.800 ;
        RECT 686.100 600.000 687.900 600.600 ;
        RECT 692.100 599.850 693.000 600.600 ;
        RECT 689.100 598.950 690.900 599.700 ;
        RECT 676.050 596.850 679.050 598.950 ;
        RECT 682.950 597.900 690.900 598.950 ;
        RECT 692.100 598.050 693.900 599.850 ;
        RECT 682.950 596.850 685.050 597.900 ;
        RECT 664.950 593.400 666.750 595.200 ;
        RECT 665.850 592.200 670.050 593.400 ;
        RECT 676.050 592.200 676.950 596.850 ;
        RECT 684.750 593.100 686.550 593.400 ;
        RECT 655.650 579.750 657.450 585.600 ;
        RECT 658.650 579.750 660.450 585.600 ;
        RECT 662.550 579.750 664.350 591.600 ;
        RECT 667.950 591.300 670.050 592.200 ;
        RECT 670.950 591.300 676.950 592.200 ;
        RECT 678.150 592.800 686.550 593.100 ;
        RECT 694.950 592.800 695.850 605.400 ;
        RECT 697.950 599.850 700.050 601.950 ;
        RECT 701.400 600.150 702.600 608.400 ;
        RECT 698.100 598.050 699.900 599.850 ;
        RECT 700.950 598.050 703.050 600.150 ;
        RECT 678.150 592.200 695.850 592.800 ;
        RECT 670.950 590.400 671.850 591.300 ;
        RECT 669.150 588.600 671.850 590.400 ;
        RECT 672.750 590.100 674.550 590.400 ;
        RECT 678.150 590.100 679.050 592.200 ;
        RECT 684.750 591.600 695.850 592.200 ;
        RECT 672.750 589.200 679.050 590.100 ;
        RECT 679.950 590.700 681.750 591.300 ;
        RECT 679.950 589.500 687.450 590.700 ;
        RECT 672.750 588.600 674.550 589.200 ;
        RECT 686.250 588.600 687.450 589.500 ;
        RECT 667.950 585.600 671.850 587.700 ;
        RECT 676.950 586.500 683.850 588.300 ;
        RECT 686.250 586.500 691.050 588.600 ;
        RECT 665.550 579.750 667.350 582.600 ;
        RECT 670.050 579.750 671.850 585.600 ;
        RECT 674.250 579.750 676.050 585.600 ;
        RECT 678.150 579.750 679.950 586.500 ;
        RECT 686.250 585.600 687.450 586.500 ;
        RECT 681.150 579.750 682.950 585.600 ;
        RECT 685.950 579.750 687.750 585.600 ;
        RECT 691.050 579.750 692.850 585.600 ;
        RECT 694.050 579.750 695.850 591.600 ;
        RECT 701.400 585.600 702.600 598.050 ;
        RECT 698.550 579.750 700.350 585.600 ;
        RECT 701.550 579.750 703.350 585.600 ;
        RECT 6.450 563.400 8.250 575.250 ;
        RECT 10.650 563.400 12.450 575.250 ;
        RECT 15.300 563.400 17.100 575.250 ;
        RECT 19.500 563.400 21.300 575.250 ;
        RECT 22.800 569.400 24.600 575.250 ;
        RECT 31.650 569.400 33.450 575.250 ;
        RECT 34.650 569.400 36.450 575.250 ;
        RECT 6.450 562.350 9.000 563.400 ;
        RECT 5.100 558.150 6.900 559.950 ;
        RECT 4.950 556.050 7.050 558.150 ;
        RECT 7.950 555.150 9.000 562.350 ;
        RECT 11.100 558.150 12.900 559.950 ;
        RECT 14.100 558.150 15.900 559.950 ;
        RECT 19.950 558.150 21.150 563.400 ;
        RECT 22.950 561.150 24.750 562.950 ;
        RECT 22.950 559.050 25.050 561.150 ;
        RECT 10.950 556.050 13.050 558.150 ;
        RECT 13.950 556.050 16.050 558.150 ;
        RECT 7.950 553.050 10.050 555.150 ;
        RECT 16.950 554.850 19.050 556.950 ;
        RECT 19.950 556.050 22.050 558.150 ;
        RECT 32.400 556.950 33.600 569.400 ;
        RECT 40.650 563.400 42.450 575.250 ;
        RECT 43.650 564.300 45.450 575.250 ;
        RECT 46.650 565.200 48.450 575.250 ;
        RECT 49.650 564.300 51.450 575.250 ;
        RECT 43.650 563.400 51.450 564.300 ;
        RECT 55.050 563.400 56.850 575.250 ;
        RECT 58.050 563.400 59.850 575.250 ;
        RECT 61.650 569.400 63.450 575.250 ;
        RECT 64.650 569.400 66.450 575.250 ;
        RECT 70.650 569.400 72.450 575.250 ;
        RECT 73.650 569.400 75.450 575.250 ;
        RECT 76.650 569.400 78.450 575.250 ;
        RECT 82.650 569.400 84.450 575.250 ;
        RECT 85.650 569.400 87.450 575.250 ;
        RECT 88.650 569.400 90.450 575.250 ;
        RECT 92.550 569.400 94.350 575.250 ;
        RECT 95.550 569.400 97.350 575.250 ;
        RECT 41.100 558.150 42.300 563.400 ;
        RECT 55.650 558.150 56.850 563.400 ;
        RECT 17.100 553.050 18.900 554.850 ;
        RECT 7.950 546.600 9.000 553.050 ;
        RECT 20.850 552.750 22.050 556.050 ;
        RECT 31.950 554.850 34.050 556.950 ;
        RECT 35.100 555.150 36.900 556.950 ;
        RECT 40.950 556.050 43.050 558.150 ;
        RECT 21.000 551.700 24.750 552.750 ;
        RECT 14.550 548.700 22.350 550.050 ;
        RECT 4.650 543.750 6.450 546.600 ;
        RECT 7.650 543.750 9.450 546.600 ;
        RECT 10.650 543.750 12.450 546.600 ;
        RECT 14.550 543.750 16.350 548.700 ;
        RECT 17.550 543.750 19.350 547.800 ;
        RECT 20.550 543.750 22.350 548.700 ;
        RECT 23.550 549.600 24.750 551.700 ;
        RECT 23.550 543.750 25.350 549.600 ;
        RECT 32.400 546.600 33.600 554.850 ;
        RECT 34.950 553.050 37.050 555.150 ;
        RECT 41.100 549.600 42.300 556.050 ;
        RECT 43.950 554.850 46.050 556.950 ;
        RECT 47.100 555.150 48.900 556.950 ;
        RECT 44.100 553.050 45.900 554.850 ;
        RECT 46.950 553.050 49.050 555.150 ;
        RECT 49.950 554.850 52.050 556.950 ;
        RECT 55.650 556.050 58.050 558.150 ;
        RECT 58.950 557.850 61.050 559.950 ;
        RECT 59.100 556.050 60.900 557.850 ;
        RECT 50.100 553.050 51.900 554.850 ;
        RECT 55.650 549.600 56.850 556.050 ;
        RECT 62.100 552.300 63.300 569.400 ;
        RECT 74.250 561.150 75.450 569.400 ;
        RECT 82.950 564.450 85.050 565.050 ;
        RECT 80.550 563.550 85.050 564.450 ;
        RECT 65.100 558.150 66.900 559.950 ;
        RECT 64.950 556.050 67.050 558.150 ;
        RECT 70.950 557.850 73.050 559.950 ;
        RECT 73.950 559.050 76.050 561.150 ;
        RECT 71.100 556.050 72.900 557.850 ;
        RECT 58.950 551.100 66.450 552.300 ;
        RECT 74.250 551.700 75.450 559.050 ;
        RECT 76.950 557.850 79.050 559.950 ;
        RECT 77.100 556.050 78.900 557.850 ;
        RECT 80.550 553.050 81.450 563.550 ;
        RECT 82.950 562.950 85.050 563.550 ;
        RECT 86.250 561.150 87.450 569.400 ;
        RECT 82.950 557.850 85.050 559.950 ;
        RECT 85.950 559.050 88.050 561.150 ;
        RECT 83.100 556.050 84.900 557.850 ;
        RECT 58.950 550.500 60.750 551.100 ;
        RECT 41.100 547.950 46.800 549.600 ;
        RECT 31.650 543.750 33.450 546.600 ;
        RECT 34.650 543.750 36.450 546.600 ;
        RECT 41.700 543.750 43.500 546.600 ;
        RECT 45.000 543.750 46.800 547.950 ;
        RECT 49.200 543.750 51.000 549.600 ;
        RECT 55.650 548.100 58.950 549.600 ;
        RECT 57.150 543.750 58.950 548.100 ;
        RECT 60.150 543.750 61.950 549.600 ;
        RECT 64.650 543.750 66.450 551.100 ;
        RECT 71.850 550.800 75.450 551.700 ;
        RECT 79.950 550.950 82.050 553.050 ;
        RECT 86.250 551.700 87.450 559.050 ;
        RECT 88.950 557.850 91.050 559.950 ;
        RECT 89.100 556.050 90.900 557.850 ;
        RECT 95.400 556.950 96.600 569.400 ;
        RECT 102.300 563.400 104.100 575.250 ;
        RECT 106.500 563.400 108.300 575.250 ;
        RECT 109.800 569.400 111.600 575.250 ;
        RECT 116.550 569.400 118.350 575.250 ;
        RECT 119.550 569.400 121.350 575.250 ;
        RECT 122.550 569.400 124.350 575.250 ;
        RECT 130.650 569.400 132.450 575.250 ;
        RECT 133.650 570.000 135.450 575.250 ;
        RECT 101.100 558.150 102.900 559.950 ;
        RECT 106.950 558.150 108.150 563.400 ;
        RECT 112.950 562.950 115.050 565.050 ;
        RECT 109.950 561.150 111.750 562.950 ;
        RECT 109.950 559.050 112.050 561.150 ;
        RECT 92.100 555.150 93.900 556.950 ;
        RECT 91.950 553.050 94.050 555.150 ;
        RECT 94.950 554.850 97.050 556.950 ;
        RECT 100.950 556.050 103.050 558.150 ;
        RECT 103.950 554.850 106.050 556.950 ;
        RECT 106.950 556.050 109.050 558.150 ;
        RECT 83.850 550.800 87.450 551.700 ;
        RECT 71.850 543.750 73.650 550.800 ;
        RECT 76.350 543.750 78.150 549.600 ;
        RECT 83.850 543.750 85.650 550.800 ;
        RECT 88.350 543.750 90.150 549.600 ;
        RECT 95.400 546.600 96.600 554.850 ;
        RECT 104.100 553.050 105.900 554.850 ;
        RECT 107.850 552.750 109.050 556.050 ;
        RECT 109.950 555.450 112.050 556.050 ;
        RECT 113.550 555.450 114.450 562.950 ;
        RECT 119.550 561.150 120.750 569.400 ;
        RECT 131.250 569.100 132.450 569.400 ;
        RECT 136.650 569.400 138.450 575.250 ;
        RECT 139.650 569.400 141.450 575.250 ;
        RECT 136.650 569.100 138.300 569.400 ;
        RECT 131.250 568.200 138.300 569.100 ;
        RECT 115.950 557.850 118.050 559.950 ;
        RECT 118.950 559.050 121.050 561.150 ;
        RECT 131.250 559.950 132.300 568.200 ;
        RECT 137.100 564.150 138.900 565.950 ;
        RECT 143.550 564.300 145.350 575.250 ;
        RECT 146.550 565.200 148.350 575.250 ;
        RECT 149.550 564.300 151.350 575.250 ;
        RECT 133.950 561.150 135.750 562.950 ;
        RECT 136.950 562.050 139.050 564.150 ;
        RECT 143.550 563.400 151.350 564.300 ;
        RECT 152.550 563.400 154.350 575.250 ;
        RECT 158.550 569.400 160.350 575.250 ;
        RECT 161.550 569.400 163.350 575.250 ;
        RECT 164.550 570.000 166.350 575.250 ;
        RECT 161.700 569.100 163.350 569.400 ;
        RECT 167.550 569.400 169.350 575.250 ;
        RECT 167.550 569.100 168.750 569.400 ;
        RECT 161.700 568.200 168.750 569.100 ;
        RECT 161.100 564.150 162.900 565.950 ;
        RECT 140.100 561.150 141.900 562.950 ;
        RECT 116.100 556.050 117.900 557.850 ;
        RECT 109.950 554.550 114.450 555.450 ;
        RECT 109.950 553.950 112.050 554.550 ;
        RECT 108.000 551.700 111.750 552.750 ;
        RECT 101.550 548.700 109.350 550.050 ;
        RECT 92.550 543.750 94.350 546.600 ;
        RECT 95.550 543.750 97.350 546.600 ;
        RECT 101.550 543.750 103.350 548.700 ;
        RECT 104.550 543.750 106.350 547.800 ;
        RECT 107.550 543.750 109.350 548.700 ;
        RECT 110.550 549.600 111.750 551.700 ;
        RECT 119.550 551.700 120.750 559.050 ;
        RECT 121.950 557.850 124.050 559.950 ;
        RECT 130.950 557.850 133.050 559.950 ;
        RECT 133.950 559.050 136.050 561.150 ;
        RECT 139.950 559.050 142.050 561.150 ;
        RECT 152.700 558.150 153.900 563.400 ;
        RECT 158.100 561.150 159.900 562.950 ;
        RECT 160.950 562.050 163.050 564.150 ;
        RECT 164.250 561.150 166.050 562.950 ;
        RECT 157.950 559.050 160.050 561.150 ;
        RECT 163.950 559.050 166.050 561.150 ;
        RECT 167.700 559.950 168.750 568.200 ;
        RECT 173.550 564.300 175.350 575.250 ;
        RECT 176.550 565.200 178.350 575.250 ;
        RECT 179.550 564.300 181.350 575.250 ;
        RECT 173.550 563.400 181.350 564.300 ;
        RECT 182.550 563.400 184.350 575.250 ;
        RECT 188.550 569.400 190.350 575.250 ;
        RECT 191.550 569.400 193.350 575.250 ;
        RECT 199.650 569.400 201.450 575.250 ;
        RECT 202.650 570.000 204.450 575.250 ;
        RECT 122.100 556.050 123.900 557.850 ;
        RECT 131.400 553.650 132.600 557.850 ;
        RECT 142.950 554.850 145.050 556.950 ;
        RECT 146.100 555.150 147.900 556.950 ;
        RECT 131.400 552.000 135.900 553.650 ;
        RECT 143.100 553.050 144.900 554.850 ;
        RECT 145.950 553.050 148.050 555.150 ;
        RECT 148.950 554.850 151.050 556.950 ;
        RECT 151.950 556.050 154.050 558.150 ;
        RECT 166.950 557.850 169.050 559.950 ;
        RECT 182.700 558.150 183.900 563.400 ;
        RECT 149.100 553.050 150.900 554.850 ;
        RECT 119.550 550.800 123.150 551.700 ;
        RECT 110.550 543.750 112.350 549.600 ;
        RECT 116.850 543.750 118.650 549.600 ;
        RECT 121.350 543.750 123.150 550.800 ;
        RECT 134.100 543.750 135.900 552.000 ;
        RECT 139.500 543.750 141.300 552.600 ;
        RECT 152.700 549.600 153.900 556.050 ;
        RECT 167.400 553.650 168.600 557.850 ;
        RECT 172.950 554.850 175.050 556.950 ;
        RECT 176.100 555.150 177.900 556.950 ;
        RECT 144.000 543.750 145.800 549.600 ;
        RECT 148.200 547.950 153.900 549.600 ;
        RECT 148.200 543.750 150.000 547.950 ;
        RECT 151.500 543.750 153.300 546.600 ;
        RECT 158.700 543.750 160.500 552.600 ;
        RECT 164.100 552.000 168.600 553.650 ;
        RECT 173.100 553.050 174.900 554.850 ;
        RECT 175.950 553.050 178.050 555.150 ;
        RECT 178.950 554.850 181.050 556.950 ;
        RECT 181.950 556.050 184.050 558.150 ;
        RECT 191.400 556.950 192.600 569.400 ;
        RECT 200.250 569.100 201.450 569.400 ;
        RECT 205.650 569.400 207.450 575.250 ;
        RECT 208.650 569.400 210.450 575.250 ;
        RECT 214.650 569.400 216.450 575.250 ;
        RECT 217.650 569.400 219.450 575.250 ;
        RECT 224.400 569.400 226.200 575.250 ;
        RECT 205.650 569.100 207.300 569.400 ;
        RECT 200.250 568.200 207.300 569.100 ;
        RECT 200.250 559.950 201.300 568.200 ;
        RECT 206.100 564.150 207.900 565.950 ;
        RECT 202.950 561.150 204.750 562.950 ;
        RECT 205.950 562.050 208.050 564.150 ;
        RECT 209.100 561.150 210.900 562.950 ;
        RECT 199.950 557.850 202.050 559.950 ;
        RECT 202.950 559.050 205.050 561.150 ;
        RECT 208.950 559.050 211.050 561.150 ;
        RECT 179.100 553.050 180.900 554.850 ;
        RECT 164.100 543.750 165.900 552.000 ;
        RECT 182.700 549.600 183.900 556.050 ;
        RECT 188.100 555.150 189.900 556.950 ;
        RECT 187.950 553.050 190.050 555.150 ;
        RECT 190.950 554.850 193.050 556.950 ;
        RECT 174.000 543.750 175.800 549.600 ;
        RECT 178.200 547.950 183.900 549.600 ;
        RECT 178.200 543.750 180.000 547.950 ;
        RECT 191.400 546.600 192.600 554.850 ;
        RECT 200.400 553.650 201.600 557.850 ;
        RECT 215.400 556.950 216.600 569.400 ;
        RECT 227.700 563.400 229.500 575.250 ;
        RECT 231.900 563.400 233.700 575.250 ;
        RECT 238.650 569.400 240.450 575.250 ;
        RECT 241.650 569.400 243.450 575.250 ;
        RECT 224.250 561.150 226.050 562.950 ;
        RECT 223.950 559.050 226.050 561.150 ;
        RECT 227.850 558.150 229.050 563.400 ;
        RECT 233.100 558.150 234.900 559.950 ;
        RECT 214.950 554.850 217.050 556.950 ;
        RECT 218.100 555.150 219.900 556.950 ;
        RECT 226.950 556.050 229.050 558.150 ;
        RECT 200.400 552.000 204.900 553.650 ;
        RECT 181.500 543.750 183.300 546.600 ;
        RECT 188.550 543.750 190.350 546.600 ;
        RECT 191.550 543.750 193.350 546.600 ;
        RECT 203.100 543.750 204.900 552.000 ;
        RECT 208.500 543.750 210.300 552.600 ;
        RECT 215.400 546.600 216.600 554.850 ;
        RECT 217.950 553.050 220.050 555.150 ;
        RECT 226.950 552.750 228.150 556.050 ;
        RECT 229.950 554.850 232.050 556.950 ;
        RECT 232.950 556.050 235.050 558.150 ;
        RECT 239.400 556.950 240.600 569.400 ;
        RECT 245.550 564.300 247.350 575.250 ;
        RECT 248.550 565.200 250.350 575.250 ;
        RECT 251.550 564.300 253.350 575.250 ;
        RECT 245.550 563.400 253.350 564.300 ;
        RECT 254.550 563.400 256.350 575.250 ;
        RECT 260.550 563.400 262.350 575.250 ;
        RECT 264.750 563.400 266.550 575.250 ;
        RECT 274.650 563.400 276.450 575.250 ;
        RECT 277.650 564.300 279.450 575.250 ;
        RECT 280.650 565.200 282.450 575.250 ;
        RECT 283.650 564.300 285.450 575.250 ;
        RECT 289.650 569.400 291.450 575.250 ;
        RECT 292.650 569.400 294.450 575.250 ;
        RECT 295.650 569.400 297.450 575.250 ;
        RECT 277.650 563.400 285.450 564.300 ;
        RECT 254.700 558.150 255.900 563.400 ;
        RECT 264.000 562.350 266.550 563.400 ;
        RECT 260.100 558.150 261.900 559.950 ;
        RECT 238.950 554.850 241.050 556.950 ;
        RECT 242.100 555.150 243.900 556.950 ;
        RECT 230.100 553.050 231.900 554.850 ;
        RECT 224.250 551.700 228.000 552.750 ;
        RECT 224.250 549.600 225.450 551.700 ;
        RECT 214.650 543.750 216.450 546.600 ;
        RECT 217.650 543.750 219.450 546.600 ;
        RECT 223.650 543.750 225.450 549.600 ;
        RECT 226.650 548.700 234.450 550.050 ;
        RECT 226.650 543.750 228.450 548.700 ;
        RECT 229.650 543.750 231.450 547.800 ;
        RECT 232.650 543.750 234.450 548.700 ;
        RECT 239.400 546.600 240.600 554.850 ;
        RECT 241.950 553.050 244.050 555.150 ;
        RECT 244.950 554.850 247.050 556.950 ;
        RECT 248.100 555.150 249.900 556.950 ;
        RECT 245.100 553.050 246.900 554.850 ;
        RECT 247.950 553.050 250.050 555.150 ;
        RECT 250.950 554.850 253.050 556.950 ;
        RECT 253.950 556.050 256.050 558.150 ;
        RECT 259.950 556.050 262.050 558.150 ;
        RECT 251.100 553.050 252.900 554.850 ;
        RECT 254.700 549.600 255.900 556.050 ;
        RECT 264.000 555.150 265.050 562.350 ;
        RECT 266.100 558.150 267.900 559.950 ;
        RECT 275.100 558.150 276.300 563.400 ;
        RECT 293.250 561.150 294.450 569.400 ;
        RECT 299.550 563.400 301.350 575.250 ;
        RECT 304.050 563.550 305.850 575.250 ;
        RECT 307.050 564.900 308.850 575.250 ;
        RECT 314.550 569.400 316.350 575.250 ;
        RECT 307.050 563.550 309.450 564.900 ;
        RECT 299.550 562.200 300.750 563.400 ;
        RECT 304.950 562.200 306.750 562.650 ;
        RECT 265.950 556.050 268.050 558.150 ;
        RECT 274.950 556.050 277.050 558.150 ;
        RECT 289.950 557.850 292.050 559.950 ;
        RECT 292.950 559.050 295.050 561.150 ;
        RECT 299.550 561.000 306.750 562.200 ;
        RECT 304.950 560.850 306.750 561.000 ;
        RECT 262.950 553.050 265.050 555.150 ;
        RECT 238.650 543.750 240.450 546.600 ;
        RECT 241.650 543.750 243.450 546.600 ;
        RECT 246.000 543.750 247.800 549.600 ;
        RECT 250.200 547.950 255.900 549.600 ;
        RECT 250.200 543.750 252.000 547.950 ;
        RECT 264.000 546.600 265.050 553.050 ;
        RECT 275.100 549.600 276.300 556.050 ;
        RECT 277.950 554.850 280.050 556.950 ;
        RECT 281.100 555.150 282.900 556.950 ;
        RECT 278.100 553.050 279.900 554.850 ;
        RECT 280.950 553.050 283.050 555.150 ;
        RECT 283.950 554.850 286.050 556.950 ;
        RECT 290.100 556.050 291.900 557.850 ;
        RECT 284.100 553.050 285.900 554.850 ;
        RECT 293.250 551.700 294.450 559.050 ;
        RECT 295.950 557.850 298.050 559.950 ;
        RECT 302.100 558.150 303.900 559.950 ;
        RECT 296.100 556.050 297.900 557.850 ;
        RECT 299.100 555.150 300.900 556.950 ;
        RECT 301.950 556.050 304.050 558.150 ;
        RECT 298.950 553.050 301.050 555.150 ;
        RECT 305.700 552.600 306.600 560.850 ;
        RECT 308.100 556.950 309.450 563.550 ;
        RECT 314.550 562.500 315.750 569.400 ;
        RECT 317.850 563.400 319.650 575.250 ;
        RECT 320.850 563.400 322.650 575.250 ;
        RECT 328.650 563.400 330.450 575.250 ;
        RECT 314.550 561.600 320.250 562.500 ;
        RECT 318.000 560.700 320.250 561.600 ;
        RECT 314.100 558.150 315.900 559.950 ;
        RECT 307.950 554.850 310.050 556.950 ;
        RECT 313.950 556.050 316.050 558.150 ;
        RECT 304.950 551.700 306.750 552.600 ;
        RECT 290.850 550.800 294.450 551.700 ;
        RECT 303.450 550.800 306.750 551.700 ;
        RECT 275.100 547.950 280.800 549.600 ;
        RECT 253.500 543.750 255.300 546.600 ;
        RECT 260.550 543.750 262.350 546.600 ;
        RECT 263.550 543.750 265.350 546.600 ;
        RECT 266.550 543.750 268.350 546.600 ;
        RECT 275.700 543.750 277.500 546.600 ;
        RECT 279.000 543.750 280.800 547.950 ;
        RECT 283.200 543.750 285.000 549.600 ;
        RECT 290.850 543.750 292.650 550.800 ;
        RECT 295.350 543.750 297.150 549.600 ;
        RECT 303.450 546.600 304.350 550.800 ;
        RECT 309.000 549.600 310.050 554.850 ;
        RECT 318.000 552.300 319.050 560.700 ;
        RECT 321.150 558.150 322.350 563.400 ;
        RECT 331.650 562.500 333.450 575.250 ;
        RECT 334.650 563.400 336.450 575.250 ;
        RECT 337.650 562.500 339.450 575.250 ;
        RECT 340.650 563.400 342.450 575.250 ;
        RECT 343.650 562.500 345.450 575.250 ;
        RECT 346.650 563.400 348.450 575.250 ;
        RECT 349.650 562.500 351.450 575.250 ;
        RECT 352.650 563.400 354.450 575.250 ;
        RECT 357.150 563.400 358.950 575.250 ;
        RECT 360.150 569.400 361.950 575.250 ;
        RECT 365.250 569.400 367.050 575.250 ;
        RECT 370.050 569.400 371.850 575.250 ;
        RECT 365.550 568.500 366.750 569.400 ;
        RECT 373.050 568.500 374.850 575.250 ;
        RECT 376.950 569.400 378.750 575.250 ;
        RECT 381.150 569.400 382.950 575.250 ;
        RECT 385.650 572.400 387.450 575.250 ;
        RECT 361.950 566.400 366.750 568.500 ;
        RECT 369.150 566.700 376.050 568.500 ;
        RECT 381.150 567.300 385.050 569.400 ;
        RECT 365.550 565.500 366.750 566.400 ;
        RECT 378.450 565.800 380.250 566.400 ;
        RECT 365.550 564.300 373.050 565.500 ;
        RECT 371.250 563.700 373.050 564.300 ;
        RECT 373.950 564.900 380.250 565.800 ;
        RECT 319.950 556.050 322.350 558.150 ;
        RECT 330.750 561.300 333.450 562.500 ;
        RECT 335.700 561.300 339.450 562.500 ;
        RECT 341.700 561.300 345.450 562.500 ;
        RECT 347.550 561.300 351.450 562.500 ;
        RECT 357.150 562.800 368.250 563.400 ;
        RECT 373.950 562.800 374.850 564.900 ;
        RECT 378.450 564.600 380.250 564.900 ;
        RECT 381.150 564.600 383.850 566.400 ;
        RECT 381.150 563.700 382.050 564.600 ;
        RECT 357.150 562.200 374.850 562.800 ;
        RECT 330.750 556.950 331.800 561.300 ;
        RECT 318.000 551.400 320.250 552.300 ;
        RECT 315.150 550.500 320.250 551.400 ;
        RECT 299.550 543.750 301.350 546.600 ;
        RECT 302.550 543.750 304.350 546.600 ;
        RECT 305.550 543.750 307.350 546.600 ;
        RECT 308.550 543.750 310.350 549.600 ;
        RECT 315.150 546.600 316.350 550.500 ;
        RECT 321.150 549.600 322.350 556.050 ;
        RECT 328.950 554.850 331.800 556.950 ;
        RECT 330.750 551.700 331.800 554.850 ;
        RECT 335.700 554.400 336.900 561.300 ;
        RECT 341.700 554.400 342.900 561.300 ;
        RECT 347.550 554.400 348.750 561.300 ;
        RECT 349.950 554.850 352.050 556.950 ;
        RECT 332.700 552.600 336.900 554.400 ;
        RECT 338.700 552.600 342.900 554.400 ;
        RECT 344.700 552.600 348.750 554.400 ;
        RECT 350.100 553.050 351.900 554.850 ;
        RECT 335.700 551.700 336.900 552.600 ;
        RECT 341.700 551.700 342.900 552.600 ;
        RECT 347.550 551.700 348.750 552.600 ;
        RECT 330.750 550.650 333.600 551.700 ;
        RECT 330.900 550.500 333.600 550.650 ;
        RECT 335.700 550.500 339.600 551.700 ;
        RECT 341.700 550.500 345.450 551.700 ;
        RECT 347.550 550.500 351.600 551.700 ;
        RECT 331.800 549.600 333.600 550.500 ;
        RECT 337.800 549.600 339.600 550.500 ;
        RECT 314.550 543.750 316.350 546.600 ;
        RECT 317.850 543.750 319.650 549.600 ;
        RECT 320.850 543.750 322.650 549.600 ;
        RECT 328.650 543.750 330.450 549.600 ;
        RECT 331.650 543.750 333.450 549.600 ;
        RECT 334.650 543.750 336.450 549.600 ;
        RECT 337.650 543.750 339.450 549.600 ;
        RECT 340.650 543.750 342.450 549.600 ;
        RECT 343.650 543.750 345.450 550.500 ;
        RECT 349.800 549.600 351.600 550.500 ;
        RECT 357.150 549.600 358.050 562.200 ;
        RECT 366.450 561.900 374.850 562.200 ;
        RECT 376.050 562.800 382.050 563.700 ;
        RECT 382.950 562.800 385.050 563.700 ;
        RECT 388.650 563.400 390.450 575.250 ;
        RECT 395.400 569.400 397.200 575.250 ;
        RECT 398.700 563.400 400.500 575.250 ;
        RECT 402.900 563.400 404.700 575.250 ;
        RECT 409.650 569.400 411.450 575.250 ;
        RECT 412.650 569.400 414.450 575.250 ;
        RECT 366.450 561.600 368.250 561.900 ;
        RECT 376.050 558.150 376.950 562.800 ;
        RECT 382.950 561.600 387.150 562.800 ;
        RECT 386.250 559.800 388.050 561.600 ;
        RECT 367.950 557.100 370.050 558.150 ;
        RECT 359.100 555.150 360.900 556.950 ;
        RECT 362.100 556.050 370.050 557.100 ;
        RECT 373.950 556.050 376.950 558.150 ;
        RECT 362.100 555.300 363.900 556.050 ;
        RECT 360.000 554.400 360.900 555.150 ;
        RECT 365.100 554.400 366.900 555.000 ;
        RECT 360.000 553.200 366.900 554.400 ;
        RECT 365.850 552.000 366.900 553.200 ;
        RECT 376.050 552.000 376.950 556.050 ;
        RECT 385.950 555.750 388.050 556.050 ;
        RECT 384.150 553.950 388.050 555.750 ;
        RECT 389.250 553.950 390.450 563.400 ;
        RECT 395.250 561.150 397.050 562.950 ;
        RECT 394.950 559.050 397.050 561.150 ;
        RECT 398.850 558.150 400.050 563.400 ;
        RECT 404.100 558.150 405.900 559.950 ;
        RECT 365.850 551.100 376.950 552.000 ;
        RECT 385.950 551.850 390.450 553.950 ;
        RECT 397.950 556.050 400.050 558.150 ;
        RECT 397.950 552.750 399.150 556.050 ;
        RECT 400.950 554.850 403.050 556.950 ;
        RECT 403.950 556.050 406.050 558.150 ;
        RECT 410.400 556.950 411.600 569.400 ;
        RECT 420.450 563.400 422.250 575.250 ;
        RECT 424.650 563.400 426.450 575.250 ;
        RECT 432.450 563.400 434.250 575.250 ;
        RECT 436.650 563.400 438.450 575.250 ;
        RECT 444.450 563.400 446.250 575.250 ;
        RECT 448.650 563.400 450.450 575.250 ;
        RECT 452.550 569.400 454.350 575.250 ;
        RECT 455.550 569.400 457.350 575.250 ;
        RECT 463.650 569.400 465.450 575.250 ;
        RECT 466.650 569.400 468.450 575.250 ;
        RECT 420.450 562.350 423.000 563.400 ;
        RECT 432.450 562.350 435.000 563.400 ;
        RECT 444.450 562.350 447.000 563.400 ;
        RECT 419.100 558.150 420.900 559.950 ;
        RECT 409.950 554.850 412.050 556.950 ;
        RECT 413.100 555.150 414.900 556.950 ;
        RECT 418.950 556.050 421.050 558.150 ;
        RECT 421.950 555.150 423.000 562.350 ;
        RECT 425.100 558.150 426.900 559.950 ;
        RECT 431.100 558.150 432.900 559.950 ;
        RECT 424.950 556.050 427.050 558.150 ;
        RECT 430.950 556.050 433.050 558.150 ;
        RECT 433.950 555.150 435.000 562.350 ;
        RECT 437.100 558.150 438.900 559.950 ;
        RECT 443.100 558.150 444.900 559.950 ;
        RECT 436.950 556.050 439.050 558.150 ;
        RECT 442.950 556.050 445.050 558.150 ;
        RECT 445.950 555.150 447.000 562.350 ;
        RECT 449.100 558.150 450.900 559.950 ;
        RECT 448.950 556.050 451.050 558.150 ;
        RECT 455.400 556.950 456.600 569.400 ;
        RECT 464.400 556.950 465.600 569.400 ;
        RECT 471.300 563.400 473.100 575.250 ;
        RECT 475.500 563.400 477.300 575.250 ;
        RECT 478.800 569.400 480.600 575.250 ;
        RECT 487.650 563.400 489.450 575.250 ;
        RECT 490.650 564.300 492.450 575.250 ;
        RECT 493.650 565.200 495.450 575.250 ;
        RECT 496.650 564.300 498.450 575.250 ;
        RECT 490.650 563.400 498.450 564.300 ;
        RECT 500.550 564.300 502.350 575.250 ;
        RECT 503.550 565.200 505.350 575.250 ;
        RECT 506.550 564.300 508.350 575.250 ;
        RECT 500.550 563.400 508.350 564.300 ;
        RECT 509.550 563.400 511.350 575.250 ;
        RECT 515.550 569.400 517.350 575.250 ;
        RECT 518.550 569.400 520.350 575.250 ;
        RECT 524.550 569.400 526.350 575.250 ;
        RECT 527.550 569.400 529.350 575.250 ;
        RECT 470.100 558.150 471.900 559.950 ;
        RECT 475.950 558.150 477.150 563.400 ;
        RECT 478.950 561.150 480.750 562.950 ;
        RECT 478.950 559.050 481.050 561.150 ;
        RECT 488.100 558.150 489.300 563.400 ;
        RECT 509.700 558.150 510.900 563.400 ;
        RECT 452.100 555.150 453.900 556.950 ;
        RECT 401.100 553.050 402.900 554.850 ;
        RECT 365.850 550.200 366.900 551.100 ;
        RECT 376.050 550.800 376.950 551.100 ;
        RECT 346.650 543.750 348.450 549.600 ;
        RECT 349.650 543.750 351.450 549.600 ;
        RECT 352.650 543.750 354.450 549.600 ;
        RECT 357.150 543.750 358.950 549.600 ;
        RECT 361.950 547.500 364.050 549.600 ;
        RECT 365.550 548.400 367.350 550.200 ;
        RECT 368.850 549.450 370.650 550.200 ;
        RECT 368.850 548.400 373.800 549.450 ;
        RECT 376.050 549.000 377.850 550.800 ;
        RECT 389.250 549.600 390.450 551.850 ;
        RECT 395.250 551.700 399.000 552.750 ;
        RECT 395.250 549.600 396.450 551.700 ;
        RECT 382.950 548.700 385.050 549.600 ;
        RECT 363.000 546.600 364.050 547.500 ;
        RECT 372.750 546.600 373.800 548.400 ;
        RECT 381.300 547.500 385.050 548.700 ;
        RECT 381.300 546.600 382.350 547.500 ;
        RECT 360.150 543.750 361.950 546.600 ;
        RECT 363.000 545.700 366.750 546.600 ;
        RECT 364.950 543.750 366.750 545.700 ;
        RECT 369.450 543.750 371.250 546.600 ;
        RECT 372.750 543.750 374.550 546.600 ;
        RECT 376.650 543.750 378.450 546.600 ;
        RECT 380.850 543.750 382.650 546.600 ;
        RECT 385.350 543.750 387.150 546.600 ;
        RECT 388.650 543.750 390.450 549.600 ;
        RECT 394.650 543.750 396.450 549.600 ;
        RECT 397.650 548.700 405.450 550.050 ;
        RECT 397.650 543.750 399.450 548.700 ;
        RECT 400.650 543.750 402.450 547.800 ;
        RECT 403.650 543.750 405.450 548.700 ;
        RECT 410.400 546.600 411.600 554.850 ;
        RECT 412.950 553.050 415.050 555.150 ;
        RECT 421.950 553.050 424.050 555.150 ;
        RECT 433.950 553.050 436.050 555.150 ;
        RECT 445.950 553.050 448.050 555.150 ;
        RECT 451.950 553.050 454.050 555.150 ;
        RECT 454.950 554.850 457.050 556.950 ;
        RECT 463.950 554.850 466.050 556.950 ;
        RECT 467.100 555.150 468.900 556.950 ;
        RECT 469.950 556.050 472.050 558.150 ;
        RECT 421.950 546.600 423.000 553.050 ;
        RECT 433.950 546.600 435.000 553.050 ;
        RECT 445.950 546.600 447.000 553.050 ;
        RECT 455.400 546.600 456.600 554.850 ;
        RECT 464.400 546.600 465.600 554.850 ;
        RECT 466.950 553.050 469.050 555.150 ;
        RECT 472.950 554.850 475.050 556.950 ;
        RECT 475.950 556.050 478.050 558.150 ;
        RECT 487.950 556.050 490.050 558.150 ;
        RECT 473.100 553.050 474.900 554.850 ;
        RECT 476.850 552.750 478.050 556.050 ;
        RECT 477.000 551.700 480.750 552.750 ;
        RECT 470.550 548.700 478.350 550.050 ;
        RECT 409.650 543.750 411.450 546.600 ;
        RECT 412.650 543.750 414.450 546.600 ;
        RECT 418.650 543.750 420.450 546.600 ;
        RECT 421.650 543.750 423.450 546.600 ;
        RECT 424.650 543.750 426.450 546.600 ;
        RECT 430.650 543.750 432.450 546.600 ;
        RECT 433.650 543.750 435.450 546.600 ;
        RECT 436.650 543.750 438.450 546.600 ;
        RECT 442.650 543.750 444.450 546.600 ;
        RECT 445.650 543.750 447.450 546.600 ;
        RECT 448.650 543.750 450.450 546.600 ;
        RECT 452.550 543.750 454.350 546.600 ;
        RECT 455.550 543.750 457.350 546.600 ;
        RECT 463.650 543.750 465.450 546.600 ;
        RECT 466.650 543.750 468.450 546.600 ;
        RECT 470.550 543.750 472.350 548.700 ;
        RECT 473.550 543.750 475.350 547.800 ;
        RECT 476.550 543.750 478.350 548.700 ;
        RECT 479.550 549.600 480.750 551.700 ;
        RECT 488.100 549.600 489.300 556.050 ;
        RECT 490.950 554.850 493.050 556.950 ;
        RECT 494.100 555.150 495.900 556.950 ;
        RECT 491.100 553.050 492.900 554.850 ;
        RECT 493.950 553.050 496.050 555.150 ;
        RECT 496.950 554.850 499.050 556.950 ;
        RECT 499.950 554.850 502.050 556.950 ;
        RECT 503.100 555.150 504.900 556.950 ;
        RECT 497.100 553.050 498.900 554.850 ;
        RECT 500.100 553.050 501.900 554.850 ;
        RECT 502.950 553.050 505.050 555.150 ;
        RECT 505.950 554.850 508.050 556.950 ;
        RECT 508.950 556.050 511.050 558.150 ;
        RECT 518.400 556.950 519.600 569.400 ;
        RECT 524.100 558.150 525.900 559.950 ;
        RECT 506.100 553.050 507.900 554.850 ;
        RECT 509.700 549.600 510.900 556.050 ;
        RECT 515.100 555.150 516.900 556.950 ;
        RECT 514.950 553.050 517.050 555.150 ;
        RECT 517.950 554.850 520.050 556.950 ;
        RECT 523.950 556.050 526.050 558.150 ;
        RECT 479.550 543.750 481.350 549.600 ;
        RECT 488.100 547.950 493.800 549.600 ;
        RECT 488.700 543.750 490.500 546.600 ;
        RECT 492.000 543.750 493.800 547.950 ;
        RECT 496.200 543.750 498.000 549.600 ;
        RECT 501.000 543.750 502.800 549.600 ;
        RECT 505.200 547.950 510.900 549.600 ;
        RECT 505.200 543.750 507.000 547.950 ;
        RECT 518.400 546.600 519.600 554.850 ;
        RECT 527.700 552.300 528.900 569.400 ;
        RECT 531.150 563.400 532.950 575.250 ;
        RECT 534.150 563.400 535.950 575.250 ;
        RECT 540.300 563.400 542.100 575.250 ;
        RECT 544.500 563.400 546.300 575.250 ;
        RECT 547.800 569.400 549.600 575.250 ;
        RECT 555.300 563.400 557.100 575.250 ;
        RECT 559.500 563.400 561.300 575.250 ;
        RECT 562.800 569.400 564.600 575.250 ;
        RECT 570.150 563.400 571.950 575.250 ;
        RECT 573.150 569.400 574.950 575.250 ;
        RECT 578.250 569.400 580.050 575.250 ;
        RECT 583.050 569.400 584.850 575.250 ;
        RECT 578.550 568.500 579.750 569.400 ;
        RECT 586.050 568.500 587.850 575.250 ;
        RECT 589.950 569.400 591.750 575.250 ;
        RECT 594.150 569.400 595.950 575.250 ;
        RECT 598.650 572.400 600.450 575.250 ;
        RECT 574.950 566.400 579.750 568.500 ;
        RECT 582.150 566.700 589.050 568.500 ;
        RECT 594.150 567.300 598.050 569.400 ;
        RECT 578.550 565.500 579.750 566.400 ;
        RECT 591.450 565.800 593.250 566.400 ;
        RECT 578.550 564.300 586.050 565.500 ;
        RECT 584.250 563.700 586.050 564.300 ;
        RECT 586.950 564.900 593.250 565.800 ;
        RECT 529.950 557.850 532.050 559.950 ;
        RECT 534.150 558.150 535.350 563.400 ;
        RECT 539.100 558.150 540.900 559.950 ;
        RECT 544.950 558.150 546.150 563.400 ;
        RECT 547.950 561.150 549.750 562.950 ;
        RECT 547.950 559.050 550.050 561.150 ;
        RECT 554.100 558.150 555.900 559.950 ;
        RECT 559.950 558.150 561.150 563.400 ;
        RECT 562.950 561.150 564.750 562.950 ;
        RECT 570.150 562.800 581.250 563.400 ;
        RECT 586.950 562.800 587.850 564.900 ;
        RECT 591.450 564.600 593.250 564.900 ;
        RECT 594.150 564.600 596.850 566.400 ;
        RECT 594.150 563.700 595.050 564.600 ;
        RECT 570.150 562.200 587.850 562.800 ;
        RECT 562.950 559.050 565.050 561.150 ;
        RECT 530.100 556.050 531.900 557.850 ;
        RECT 532.950 556.050 535.350 558.150 ;
        RECT 538.950 556.050 541.050 558.150 ;
        RECT 524.550 551.100 532.050 552.300 ;
        RECT 508.500 543.750 510.300 546.600 ;
        RECT 515.550 543.750 517.350 546.600 ;
        RECT 518.550 543.750 520.350 546.600 ;
        RECT 524.550 543.750 526.350 551.100 ;
        RECT 530.250 550.500 532.050 551.100 ;
        RECT 534.150 549.600 535.350 556.050 ;
        RECT 541.950 554.850 544.050 556.950 ;
        RECT 544.950 556.050 547.050 558.150 ;
        RECT 553.950 556.050 556.050 558.150 ;
        RECT 542.100 553.050 543.900 554.850 ;
        RECT 545.850 552.750 547.050 556.050 ;
        RECT 556.950 554.850 559.050 556.950 ;
        RECT 559.950 556.050 562.050 558.150 ;
        RECT 557.100 553.050 558.900 554.850 ;
        RECT 560.850 552.750 562.050 556.050 ;
        RECT 546.000 551.700 549.750 552.750 ;
        RECT 561.000 551.700 564.750 552.750 ;
        RECT 529.050 543.750 530.850 549.600 ;
        RECT 532.050 548.100 535.350 549.600 ;
        RECT 539.550 548.700 547.350 550.050 ;
        RECT 532.050 543.750 533.850 548.100 ;
        RECT 539.550 543.750 541.350 548.700 ;
        RECT 542.550 543.750 544.350 547.800 ;
        RECT 545.550 543.750 547.350 548.700 ;
        RECT 548.550 549.600 549.750 551.700 ;
        RECT 548.550 543.750 550.350 549.600 ;
        RECT 554.550 548.700 562.350 550.050 ;
        RECT 554.550 543.750 556.350 548.700 ;
        RECT 557.550 543.750 559.350 547.800 ;
        RECT 560.550 543.750 562.350 548.700 ;
        RECT 563.550 549.600 564.750 551.700 ;
        RECT 570.150 549.600 571.050 562.200 ;
        RECT 579.450 561.900 587.850 562.200 ;
        RECT 589.050 562.800 595.050 563.700 ;
        RECT 595.950 562.800 598.050 563.700 ;
        RECT 601.650 563.400 603.450 575.250 ;
        RECT 579.450 561.600 581.250 561.900 ;
        RECT 589.050 558.150 589.950 562.800 ;
        RECT 595.950 561.600 600.150 562.800 ;
        RECT 599.250 559.800 601.050 561.600 ;
        RECT 580.950 557.100 583.050 558.150 ;
        RECT 572.100 555.150 573.900 556.950 ;
        RECT 575.100 556.050 583.050 557.100 ;
        RECT 586.950 556.050 589.950 558.150 ;
        RECT 575.100 555.300 576.900 556.050 ;
        RECT 573.000 554.400 573.900 555.150 ;
        RECT 578.100 554.400 579.900 555.000 ;
        RECT 573.000 553.200 579.900 554.400 ;
        RECT 578.850 552.000 579.900 553.200 ;
        RECT 589.050 552.000 589.950 556.050 ;
        RECT 598.950 555.750 601.050 556.050 ;
        RECT 597.150 553.950 601.050 555.750 ;
        RECT 602.250 553.950 603.450 563.400 ;
        RECT 605.550 569.400 607.350 575.250 ;
        RECT 605.550 562.500 606.750 569.400 ;
        RECT 608.850 563.400 610.650 575.250 ;
        RECT 611.850 563.400 613.650 575.250 ;
        RECT 621.450 563.400 623.250 575.250 ;
        RECT 625.650 563.400 627.450 575.250 ;
        RECT 629.550 564.300 631.350 575.250 ;
        RECT 632.550 565.200 634.350 575.250 ;
        RECT 635.550 564.300 637.350 575.250 ;
        RECT 629.550 563.400 637.350 564.300 ;
        RECT 638.550 563.400 640.350 575.250 ;
        RECT 644.550 563.400 646.350 575.250 ;
        RECT 647.550 572.400 649.350 575.250 ;
        RECT 652.050 569.400 653.850 575.250 ;
        RECT 656.250 569.400 658.050 575.250 ;
        RECT 649.950 567.300 653.850 569.400 ;
        RECT 660.150 568.500 661.950 575.250 ;
        RECT 663.150 569.400 664.950 575.250 ;
        RECT 667.950 569.400 669.750 575.250 ;
        RECT 673.050 569.400 674.850 575.250 ;
        RECT 668.250 568.500 669.450 569.400 ;
        RECT 658.950 566.700 665.850 568.500 ;
        RECT 668.250 566.400 673.050 568.500 ;
        RECT 651.150 564.600 653.850 566.400 ;
        RECT 654.750 565.800 656.550 566.400 ;
        RECT 654.750 564.900 661.050 565.800 ;
        RECT 668.250 565.500 669.450 566.400 ;
        RECT 654.750 564.600 656.550 564.900 ;
        RECT 652.950 563.700 653.850 564.600 ;
        RECT 605.550 561.600 611.250 562.500 ;
        RECT 609.000 560.700 611.250 561.600 ;
        RECT 605.100 558.150 606.900 559.950 ;
        RECT 604.950 556.050 607.050 558.150 ;
        RECT 578.850 551.100 589.950 552.000 ;
        RECT 598.950 551.850 603.450 553.950 ;
        RECT 578.850 550.200 579.900 551.100 ;
        RECT 589.050 550.800 589.950 551.100 ;
        RECT 563.550 543.750 565.350 549.600 ;
        RECT 570.150 543.750 571.950 549.600 ;
        RECT 574.950 547.500 577.050 549.600 ;
        RECT 578.550 548.400 580.350 550.200 ;
        RECT 581.850 549.450 583.650 550.200 ;
        RECT 581.850 548.400 586.800 549.450 ;
        RECT 589.050 549.000 590.850 550.800 ;
        RECT 602.250 549.600 603.450 551.850 ;
        RECT 609.000 552.300 610.050 560.700 ;
        RECT 612.150 558.150 613.350 563.400 ;
        RECT 621.450 562.350 624.000 563.400 ;
        RECT 620.100 558.150 621.900 559.950 ;
        RECT 610.950 556.050 613.350 558.150 ;
        RECT 619.950 556.050 622.050 558.150 ;
        RECT 609.000 551.400 611.250 552.300 ;
        RECT 595.950 548.700 598.050 549.600 ;
        RECT 576.000 546.600 577.050 547.500 ;
        RECT 585.750 546.600 586.800 548.400 ;
        RECT 594.300 547.500 598.050 548.700 ;
        RECT 594.300 546.600 595.350 547.500 ;
        RECT 573.150 543.750 574.950 546.600 ;
        RECT 576.000 545.700 579.750 546.600 ;
        RECT 577.950 543.750 579.750 545.700 ;
        RECT 582.450 543.750 584.250 546.600 ;
        RECT 585.750 543.750 587.550 546.600 ;
        RECT 589.650 543.750 591.450 546.600 ;
        RECT 593.850 543.750 595.650 546.600 ;
        RECT 598.350 543.750 600.150 546.600 ;
        RECT 601.650 543.750 603.450 549.600 ;
        RECT 606.150 550.500 611.250 551.400 ;
        RECT 606.150 546.600 607.350 550.500 ;
        RECT 612.150 549.600 613.350 556.050 ;
        RECT 622.950 555.150 624.000 562.350 ;
        RECT 626.100 558.150 627.900 559.950 ;
        RECT 638.700 558.150 639.900 563.400 ;
        RECT 625.950 556.050 628.050 558.150 ;
        RECT 622.950 553.050 625.050 555.150 ;
        RECT 628.950 554.850 631.050 556.950 ;
        RECT 632.100 555.150 633.900 556.950 ;
        RECT 629.100 553.050 630.900 554.850 ;
        RECT 631.950 553.050 634.050 555.150 ;
        RECT 634.950 554.850 637.050 556.950 ;
        RECT 637.950 556.050 640.050 558.150 ;
        RECT 635.100 553.050 636.900 554.850 ;
        RECT 605.550 543.750 607.350 546.600 ;
        RECT 608.850 543.750 610.650 549.600 ;
        RECT 611.850 543.750 613.650 549.600 ;
        RECT 622.950 546.600 624.000 553.050 ;
        RECT 638.700 549.600 639.900 556.050 ;
        RECT 619.650 543.750 621.450 546.600 ;
        RECT 622.650 543.750 624.450 546.600 ;
        RECT 625.650 543.750 627.450 546.600 ;
        RECT 630.000 543.750 631.800 549.600 ;
        RECT 634.200 547.950 639.900 549.600 ;
        RECT 644.550 553.950 645.750 563.400 ;
        RECT 649.950 562.800 652.050 563.700 ;
        RECT 652.950 562.800 658.950 563.700 ;
        RECT 647.850 561.600 652.050 562.800 ;
        RECT 646.950 559.800 648.750 561.600 ;
        RECT 658.050 558.150 658.950 562.800 ;
        RECT 660.150 562.800 661.050 564.900 ;
        RECT 661.950 564.300 669.450 565.500 ;
        RECT 661.950 563.700 663.750 564.300 ;
        RECT 676.050 563.400 677.850 575.250 ;
        RECT 666.750 562.800 677.850 563.400 ;
        RECT 660.150 562.200 677.850 562.800 ;
        RECT 660.150 561.900 668.550 562.200 ;
        RECT 666.750 561.600 668.550 561.900 ;
        RECT 658.050 556.050 661.050 558.150 ;
        RECT 664.950 557.100 667.050 558.150 ;
        RECT 664.950 556.050 672.900 557.100 ;
        RECT 646.950 555.750 649.050 556.050 ;
        RECT 646.950 553.950 650.850 555.750 ;
        RECT 644.550 551.850 649.050 553.950 ;
        RECT 658.050 552.000 658.950 556.050 ;
        RECT 671.100 555.300 672.900 556.050 ;
        RECT 674.100 555.150 675.900 556.950 ;
        RECT 668.100 554.400 669.900 555.000 ;
        RECT 674.100 554.400 675.000 555.150 ;
        RECT 668.100 553.200 675.000 554.400 ;
        RECT 668.100 552.000 669.150 553.200 ;
        RECT 644.550 549.600 645.750 551.850 ;
        RECT 658.050 551.100 669.150 552.000 ;
        RECT 658.050 550.800 658.950 551.100 ;
        RECT 634.200 543.750 636.000 547.950 ;
        RECT 637.500 543.750 639.300 546.600 ;
        RECT 644.550 543.750 646.350 549.600 ;
        RECT 649.950 548.700 652.050 549.600 ;
        RECT 657.150 549.000 658.950 550.800 ;
        RECT 668.100 550.200 669.150 551.100 ;
        RECT 664.350 549.450 666.150 550.200 ;
        RECT 649.950 547.500 653.700 548.700 ;
        RECT 652.650 546.600 653.700 547.500 ;
        RECT 661.200 548.400 666.150 549.450 ;
        RECT 667.650 548.400 669.450 550.200 ;
        RECT 676.950 549.600 677.850 562.200 ;
        RECT 680.550 569.400 682.350 575.250 ;
        RECT 680.550 562.500 681.750 569.400 ;
        RECT 683.850 563.400 685.650 575.250 ;
        RECT 686.850 563.400 688.650 575.250 ;
        RECT 694.650 569.400 696.450 575.250 ;
        RECT 697.650 569.400 699.450 575.250 ;
        RECT 701.550 569.400 703.350 575.250 ;
        RECT 704.550 569.400 706.350 575.250 ;
        RECT 680.550 561.600 686.250 562.500 ;
        RECT 684.000 560.700 686.250 561.600 ;
        RECT 680.100 558.150 681.900 559.950 ;
        RECT 679.950 556.050 682.050 558.150 ;
        RECT 684.000 552.300 685.050 560.700 ;
        RECT 687.150 558.150 688.350 563.400 ;
        RECT 685.950 556.050 688.350 558.150 ;
        RECT 695.400 556.950 696.600 569.400 ;
        RECT 704.400 556.950 705.600 569.400 ;
        RECT 684.000 551.400 686.250 552.300 ;
        RECT 661.200 546.600 662.250 548.400 ;
        RECT 670.950 547.500 673.050 549.600 ;
        RECT 670.950 546.600 672.000 547.500 ;
        RECT 647.850 543.750 649.650 546.600 ;
        RECT 652.350 543.750 654.150 546.600 ;
        RECT 656.550 543.750 658.350 546.600 ;
        RECT 660.450 543.750 662.250 546.600 ;
        RECT 663.750 543.750 665.550 546.600 ;
        RECT 668.250 545.700 672.000 546.600 ;
        RECT 668.250 543.750 670.050 545.700 ;
        RECT 673.050 543.750 674.850 546.600 ;
        RECT 676.050 543.750 677.850 549.600 ;
        RECT 681.150 550.500 686.250 551.400 ;
        RECT 681.150 546.600 682.350 550.500 ;
        RECT 687.150 549.600 688.350 556.050 ;
        RECT 694.950 554.850 697.050 556.950 ;
        RECT 698.100 555.150 699.900 556.950 ;
        RECT 701.100 555.150 702.900 556.950 ;
        RECT 680.550 543.750 682.350 546.600 ;
        RECT 683.850 543.750 685.650 549.600 ;
        RECT 686.850 543.750 688.650 549.600 ;
        RECT 695.400 546.600 696.600 554.850 ;
        RECT 697.950 553.050 700.050 555.150 ;
        RECT 700.950 553.050 703.050 555.150 ;
        RECT 703.950 554.850 706.050 556.950 ;
        RECT 704.400 546.600 705.600 554.850 ;
        RECT 694.650 543.750 696.450 546.600 ;
        RECT 697.650 543.750 699.450 546.600 ;
        RECT 701.550 543.750 703.350 546.600 ;
        RECT 704.550 543.750 706.350 546.600 ;
        RECT 5.850 532.200 7.650 539.250 ;
        RECT 10.350 533.400 12.150 539.250 ;
        RECT 15.150 533.400 16.950 539.250 ;
        RECT 18.150 536.400 19.950 539.250 ;
        RECT 22.950 537.300 24.750 539.250 ;
        RECT 21.000 536.400 24.750 537.300 ;
        RECT 27.450 536.400 29.250 539.250 ;
        RECT 30.750 536.400 32.550 539.250 ;
        RECT 34.650 536.400 36.450 539.250 ;
        RECT 38.850 536.400 40.650 539.250 ;
        RECT 43.350 536.400 45.150 539.250 ;
        RECT 21.000 535.500 22.050 536.400 ;
        RECT 19.950 533.400 22.050 535.500 ;
        RECT 30.750 534.600 31.800 536.400 ;
        RECT 5.850 531.300 9.450 532.200 ;
        RECT 5.100 525.150 6.900 526.950 ;
        RECT 4.950 523.050 7.050 525.150 ;
        RECT 8.250 523.950 9.450 531.300 ;
        RECT 11.100 525.150 12.900 526.950 ;
        RECT 7.950 521.850 10.050 523.950 ;
        RECT 10.950 523.050 13.050 525.150 ;
        RECT 8.250 513.600 9.450 521.850 ;
        RECT 15.150 520.800 16.050 533.400 ;
        RECT 23.550 532.800 25.350 534.600 ;
        RECT 26.850 533.550 31.800 534.600 ;
        RECT 39.300 535.500 40.350 536.400 ;
        RECT 39.300 534.300 43.050 535.500 ;
        RECT 26.850 532.800 28.650 533.550 ;
        RECT 23.850 531.900 24.900 532.800 ;
        RECT 34.050 532.200 35.850 534.000 ;
        RECT 40.950 533.400 43.050 534.300 ;
        RECT 46.650 533.400 48.450 539.250 ;
        RECT 52.650 536.400 54.450 539.250 ;
        RECT 55.650 536.400 57.450 539.250 ;
        RECT 34.050 531.900 34.950 532.200 ;
        RECT 23.850 531.000 34.950 531.900 ;
        RECT 47.250 531.150 48.450 533.400 ;
        RECT 23.850 529.800 24.900 531.000 ;
        RECT 18.000 528.600 24.900 529.800 ;
        RECT 18.000 527.850 18.900 528.600 ;
        RECT 23.100 528.000 24.900 528.600 ;
        RECT 17.100 526.050 18.900 527.850 ;
        RECT 20.100 526.950 21.900 527.700 ;
        RECT 34.050 526.950 34.950 531.000 ;
        RECT 43.950 529.050 48.450 531.150 ;
        RECT 42.150 527.250 46.050 529.050 ;
        RECT 43.950 526.950 46.050 527.250 ;
        RECT 20.100 525.900 28.050 526.950 ;
        RECT 25.950 524.850 28.050 525.900 ;
        RECT 31.950 524.850 34.950 526.950 ;
        RECT 24.450 521.100 26.250 521.400 ;
        RECT 24.450 520.800 32.850 521.100 ;
        RECT 15.150 520.200 32.850 520.800 ;
        RECT 15.150 519.600 26.250 520.200 ;
        RECT 4.650 507.750 6.450 513.600 ;
        RECT 7.650 507.750 9.450 513.600 ;
        RECT 10.650 507.750 12.450 513.600 ;
        RECT 15.150 507.750 16.950 519.600 ;
        RECT 29.250 518.700 31.050 519.300 ;
        RECT 23.550 517.500 31.050 518.700 ;
        RECT 31.950 518.100 32.850 520.200 ;
        RECT 34.050 520.200 34.950 524.850 ;
        RECT 44.250 521.400 46.050 523.200 ;
        RECT 40.950 520.200 45.150 521.400 ;
        RECT 34.050 519.300 40.050 520.200 ;
        RECT 40.950 519.300 43.050 520.200 ;
        RECT 47.250 519.600 48.450 529.050 ;
        RECT 53.400 528.150 54.600 536.400 ;
        RECT 62.850 532.200 64.650 539.250 ;
        RECT 67.350 533.400 69.150 539.250 ;
        RECT 73.650 533.400 75.450 539.250 ;
        RECT 62.850 531.300 66.450 532.200 ;
        RECT 52.950 526.050 55.050 528.150 ;
        RECT 55.950 527.850 58.050 529.950 ;
        RECT 56.100 526.050 57.900 527.850 ;
        RECT 39.150 518.400 40.050 519.300 ;
        RECT 36.450 518.100 38.250 518.400 ;
        RECT 23.550 516.600 24.750 517.500 ;
        RECT 31.950 517.200 38.250 518.100 ;
        RECT 36.450 516.600 38.250 517.200 ;
        RECT 39.150 516.600 41.850 518.400 ;
        RECT 19.950 514.500 24.750 516.600 ;
        RECT 27.150 514.500 34.050 516.300 ;
        RECT 23.550 513.600 24.750 514.500 ;
        RECT 18.150 507.750 19.950 513.600 ;
        RECT 23.250 507.750 25.050 513.600 ;
        RECT 28.050 507.750 29.850 513.600 ;
        RECT 31.050 507.750 32.850 514.500 ;
        RECT 39.150 513.600 43.050 515.700 ;
        RECT 34.950 507.750 36.750 513.600 ;
        RECT 39.150 507.750 40.950 513.600 ;
        RECT 43.650 507.750 45.450 510.600 ;
        RECT 46.650 507.750 48.450 519.600 ;
        RECT 53.400 513.600 54.600 526.050 ;
        RECT 62.100 525.150 63.900 526.950 ;
        RECT 61.950 523.050 64.050 525.150 ;
        RECT 65.250 523.950 66.450 531.300 ;
        RECT 74.250 531.300 75.450 533.400 ;
        RECT 76.650 534.300 78.450 539.250 ;
        RECT 79.650 535.200 81.450 539.250 ;
        RECT 82.650 534.300 84.450 539.250 ;
        RECT 76.650 532.950 84.450 534.300 ;
        RECT 88.650 533.400 90.450 539.250 ;
        RECT 89.250 531.300 90.450 533.400 ;
        RECT 91.650 534.300 93.450 539.250 ;
        RECT 94.650 535.200 96.450 539.250 ;
        RECT 97.650 534.300 99.450 539.250 ;
        RECT 91.650 532.950 99.450 534.300 ;
        RECT 101.850 533.400 103.650 539.250 ;
        RECT 106.350 532.200 108.150 539.250 ;
        RECT 113.550 534.000 115.350 539.250 ;
        RECT 116.550 534.900 118.350 539.250 ;
        RECT 119.550 538.500 127.350 539.250 ;
        RECT 119.550 534.000 121.350 538.500 ;
        RECT 113.550 533.100 121.350 534.000 ;
        RECT 122.550 533.400 124.350 537.600 ;
        RECT 125.550 533.400 127.350 538.500 ;
        RECT 131.550 536.400 133.350 539.250 ;
        RECT 134.550 536.400 136.350 539.250 ;
        RECT 104.550 531.300 108.150 532.200 ;
        RECT 122.850 531.900 123.750 533.400 ;
        RECT 74.250 530.250 78.000 531.300 ;
        RECT 89.250 530.250 93.000 531.300 ;
        RECT 76.950 526.950 78.150 530.250 ;
        RECT 80.100 528.150 81.900 529.950 ;
        RECT 68.100 525.150 69.900 526.950 ;
        RECT 64.950 521.850 67.050 523.950 ;
        RECT 67.950 523.050 70.050 525.150 ;
        RECT 76.950 524.850 79.050 526.950 ;
        RECT 79.950 526.050 82.050 528.150 ;
        RECT 91.950 526.950 93.150 530.250 ;
        RECT 95.100 528.150 96.900 529.950 ;
        RECT 82.950 524.850 85.050 526.950 ;
        RECT 91.950 524.850 94.050 526.950 ;
        RECT 94.950 526.050 97.050 528.150 ;
        RECT 97.950 524.850 100.050 526.950 ;
        RECT 101.100 525.150 102.900 526.950 ;
        RECT 73.950 521.850 76.050 523.950 ;
        RECT 65.250 513.600 66.450 521.850 ;
        RECT 74.250 520.050 76.050 521.850 ;
        RECT 77.850 519.600 79.050 524.850 ;
        RECT 83.100 523.050 84.900 524.850 ;
        RECT 88.950 521.850 91.050 523.950 ;
        RECT 89.250 520.050 91.050 521.850 ;
        RECT 92.850 519.600 94.050 524.850 ;
        RECT 98.100 523.050 99.900 524.850 ;
        RECT 100.950 523.050 103.050 525.150 ;
        RECT 104.550 523.950 105.750 531.300 ;
        RECT 119.400 530.850 123.750 531.900 ;
        RECT 116.100 528.150 117.900 529.950 ;
        RECT 107.100 525.150 108.900 526.950 ;
        RECT 103.950 521.850 106.050 523.950 ;
        RECT 106.950 523.050 109.050 525.150 ;
        RECT 112.950 524.850 115.050 526.950 ;
        RECT 115.950 526.050 118.050 528.150 ;
        RECT 119.400 526.950 120.600 530.850 ;
        RECT 121.500 528.150 123.300 529.950 ;
        RECT 118.950 524.850 121.050 526.950 ;
        RECT 121.950 526.050 124.050 528.150 ;
        RECT 130.950 527.850 133.050 529.950 ;
        RECT 134.400 528.150 135.600 536.400 ;
        RECT 142.950 534.450 145.050 535.050 ;
        RECT 140.550 533.550 145.050 534.450 ;
        RECT 124.950 524.850 127.050 526.950 ;
        RECT 131.100 526.050 132.900 527.850 ;
        RECT 133.950 526.050 136.050 528.150 ;
        RECT 113.100 523.050 114.900 524.850 ;
        RECT 52.650 507.750 54.450 513.600 ;
        RECT 55.650 507.750 57.450 513.600 ;
        RECT 61.650 507.750 63.450 513.600 ;
        RECT 64.650 507.750 66.450 513.600 ;
        RECT 67.650 507.750 69.450 513.600 ;
        RECT 74.400 507.750 76.200 513.600 ;
        RECT 77.700 507.750 79.500 519.600 ;
        RECT 81.900 507.750 83.700 519.600 ;
        RECT 89.400 507.750 91.200 513.600 ;
        RECT 92.700 507.750 94.500 519.600 ;
        RECT 96.900 507.750 98.700 519.600 ;
        RECT 104.550 513.600 105.750 521.850 ;
        RECT 119.550 519.600 120.750 524.850 ;
        RECT 124.950 523.050 126.750 524.850 ;
        RECT 101.550 507.750 103.350 513.600 ;
        RECT 104.550 507.750 106.350 513.600 ;
        RECT 107.550 507.750 109.350 513.600 ;
        RECT 113.550 507.750 115.350 519.600 ;
        RECT 118.050 507.750 121.350 519.600 ;
        RECT 124.050 507.750 125.850 519.600 ;
        RECT 134.400 513.600 135.600 526.050 ;
        RECT 140.550 520.050 141.450 533.550 ;
        RECT 142.950 532.950 145.050 533.550 ;
        RECT 146.100 531.000 147.900 539.250 ;
        RECT 143.400 529.350 147.900 531.000 ;
        RECT 151.500 530.400 153.300 539.250 ;
        RECT 156.000 533.400 157.800 539.250 ;
        RECT 160.200 535.050 162.000 539.250 ;
        RECT 163.500 536.400 165.300 539.250 ;
        RECT 170.550 536.400 172.350 539.250 ;
        RECT 173.550 536.400 175.350 539.250 ;
        RECT 176.550 536.400 178.350 539.250 ;
        RECT 160.200 533.400 165.900 535.050 ;
        RECT 143.400 525.150 144.600 529.350 ;
        RECT 155.100 528.150 156.900 529.950 ;
        RECT 154.950 526.050 157.050 528.150 ;
        RECT 157.950 527.850 160.050 529.950 ;
        RECT 161.100 528.150 162.900 529.950 ;
        RECT 158.100 526.050 159.900 527.850 ;
        RECT 160.950 526.050 163.050 528.150 ;
        RECT 164.700 526.950 165.900 533.400 ;
        RECT 174.000 529.950 175.050 536.400 ;
        RECT 182.850 533.400 184.650 539.250 ;
        RECT 187.350 532.200 189.150 539.250 ;
        RECT 194.850 533.400 196.650 539.250 ;
        RECT 199.350 532.200 201.150 539.250 ;
        RECT 206.550 534.300 208.350 539.250 ;
        RECT 209.550 535.200 211.350 539.250 ;
        RECT 212.550 534.300 214.350 539.250 ;
        RECT 206.550 532.950 214.350 534.300 ;
        RECT 215.550 533.400 217.350 539.250 ;
        RECT 222.150 533.400 223.950 539.250 ;
        RECT 225.150 536.400 226.950 539.250 ;
        RECT 229.950 537.300 231.750 539.250 ;
        RECT 228.000 536.400 231.750 537.300 ;
        RECT 234.450 536.400 236.250 539.250 ;
        RECT 237.750 536.400 239.550 539.250 ;
        RECT 241.650 536.400 243.450 539.250 ;
        RECT 245.850 536.400 247.650 539.250 ;
        RECT 250.350 536.400 252.150 539.250 ;
        RECT 228.000 535.500 229.050 536.400 ;
        RECT 226.950 533.400 229.050 535.500 ;
        RECT 237.750 534.600 238.800 536.400 ;
        RECT 172.950 527.850 175.050 529.950 ;
        RECT 142.950 523.050 145.050 525.150 ;
        RECT 163.950 524.850 166.050 526.950 ;
        RECT 169.950 524.850 172.050 526.950 ;
        RECT 139.950 517.950 142.050 520.050 ;
        RECT 143.250 514.800 144.300 523.050 ;
        RECT 145.950 521.850 148.050 523.950 ;
        RECT 151.950 521.850 154.050 523.950 ;
        RECT 145.950 520.050 147.750 521.850 ;
        RECT 148.950 518.850 151.050 520.950 ;
        RECT 152.100 520.050 153.900 521.850 ;
        RECT 164.700 519.600 165.900 524.850 ;
        RECT 170.100 523.050 171.900 524.850 ;
        RECT 174.000 520.650 175.050 527.850 ;
        RECT 185.550 531.300 189.150 532.200 ;
        RECT 197.550 531.300 201.150 532.200 ;
        RECT 215.550 531.300 216.750 533.400 ;
        RECT 175.950 524.850 178.050 526.950 ;
        RECT 182.100 525.150 183.900 526.950 ;
        RECT 176.100 523.050 177.900 524.850 ;
        RECT 181.950 523.050 184.050 525.150 ;
        RECT 185.550 523.950 186.750 531.300 ;
        RECT 188.100 525.150 189.900 526.950 ;
        RECT 194.100 525.150 195.900 526.950 ;
        RECT 184.950 521.850 187.050 523.950 ;
        RECT 187.950 523.050 190.050 525.150 ;
        RECT 193.950 523.050 196.050 525.150 ;
        RECT 197.550 523.950 198.750 531.300 ;
        RECT 213.000 530.250 216.750 531.300 ;
        RECT 209.100 528.150 210.900 529.950 ;
        RECT 200.100 525.150 201.900 526.950 ;
        RECT 196.950 521.850 199.050 523.950 ;
        RECT 199.950 523.050 202.050 525.150 ;
        RECT 205.950 524.850 208.050 526.950 ;
        RECT 208.950 526.050 211.050 528.150 ;
        RECT 212.850 526.950 214.050 530.250 ;
        RECT 211.950 524.850 214.050 526.950 ;
        RECT 206.100 523.050 207.900 524.850 ;
        RECT 174.000 519.600 176.550 520.650 ;
        RECT 149.100 517.050 150.900 518.850 ;
        RECT 155.550 518.700 163.350 519.600 ;
        RECT 143.250 513.900 150.300 514.800 ;
        RECT 143.250 513.600 144.450 513.900 ;
        RECT 131.550 507.750 133.350 513.600 ;
        RECT 134.550 507.750 136.350 513.600 ;
        RECT 142.650 507.750 144.450 513.600 ;
        RECT 148.650 513.600 150.300 513.900 ;
        RECT 145.650 507.750 147.450 513.000 ;
        RECT 148.650 507.750 150.450 513.600 ;
        RECT 151.650 507.750 153.450 513.600 ;
        RECT 155.550 507.750 157.350 518.700 ;
        RECT 158.550 507.750 160.350 517.800 ;
        RECT 161.550 507.750 163.350 518.700 ;
        RECT 164.550 507.750 166.350 519.600 ;
        RECT 170.550 507.750 172.350 519.600 ;
        RECT 174.750 507.750 176.550 519.600 ;
        RECT 185.550 513.600 186.750 521.850 ;
        RECT 197.550 513.600 198.750 521.850 ;
        RECT 211.950 519.600 213.150 524.850 ;
        RECT 214.950 521.850 217.050 523.950 ;
        RECT 214.950 520.050 216.750 521.850 ;
        RECT 222.150 520.800 223.050 533.400 ;
        RECT 230.550 532.800 232.350 534.600 ;
        RECT 233.850 533.550 238.800 534.600 ;
        RECT 246.300 535.500 247.350 536.400 ;
        RECT 246.300 534.300 250.050 535.500 ;
        RECT 233.850 532.800 235.650 533.550 ;
        RECT 230.850 531.900 231.900 532.800 ;
        RECT 241.050 532.200 242.850 534.000 ;
        RECT 247.950 533.400 250.050 534.300 ;
        RECT 253.650 533.400 255.450 539.250 ;
        RECT 241.050 531.900 241.950 532.200 ;
        RECT 230.850 531.000 241.950 531.900 ;
        RECT 254.250 531.150 255.450 533.400 ;
        RECT 260.850 532.200 262.650 539.250 ;
        RECT 265.350 533.400 267.150 539.250 ;
        RECT 269.550 534.300 271.350 539.250 ;
        RECT 272.550 535.200 274.350 539.250 ;
        RECT 275.550 534.300 277.350 539.250 ;
        RECT 269.550 532.950 277.350 534.300 ;
        RECT 278.550 533.400 280.350 539.250 ;
        RECT 284.550 533.400 286.350 539.250 ;
        RECT 287.550 533.400 289.350 539.250 ;
        RECT 260.850 531.300 264.450 532.200 ;
        RECT 278.550 531.300 279.750 533.400 ;
        RECT 230.850 529.800 231.900 531.000 ;
        RECT 225.000 528.600 231.900 529.800 ;
        RECT 225.000 527.850 225.900 528.600 ;
        RECT 230.100 528.000 231.900 528.600 ;
        RECT 224.100 526.050 225.900 527.850 ;
        RECT 227.100 526.950 228.900 527.700 ;
        RECT 241.050 526.950 241.950 531.000 ;
        RECT 250.950 529.050 255.450 531.150 ;
        RECT 249.150 527.250 253.050 529.050 ;
        RECT 250.950 526.950 253.050 527.250 ;
        RECT 227.100 525.900 235.050 526.950 ;
        RECT 232.950 524.850 235.050 525.900 ;
        RECT 238.950 524.850 241.950 526.950 ;
        RECT 231.450 521.100 233.250 521.400 ;
        RECT 231.450 520.800 239.850 521.100 ;
        RECT 222.150 520.200 239.850 520.800 ;
        RECT 222.150 519.600 233.250 520.200 ;
        RECT 182.550 507.750 184.350 513.600 ;
        RECT 185.550 507.750 187.350 513.600 ;
        RECT 188.550 507.750 190.350 513.600 ;
        RECT 194.550 507.750 196.350 513.600 ;
        RECT 197.550 507.750 199.350 513.600 ;
        RECT 200.550 507.750 202.350 513.600 ;
        RECT 207.300 507.750 209.100 519.600 ;
        RECT 211.500 507.750 213.300 519.600 ;
        RECT 214.800 507.750 216.600 513.600 ;
        RECT 222.150 507.750 223.950 519.600 ;
        RECT 236.250 518.700 238.050 519.300 ;
        RECT 230.550 517.500 238.050 518.700 ;
        RECT 238.950 518.100 239.850 520.200 ;
        RECT 241.050 520.200 241.950 524.850 ;
        RECT 251.250 521.400 253.050 523.200 ;
        RECT 247.950 520.200 252.150 521.400 ;
        RECT 241.050 519.300 247.050 520.200 ;
        RECT 247.950 519.300 250.050 520.200 ;
        RECT 254.250 519.600 255.450 529.050 ;
        RECT 260.100 525.150 261.900 526.950 ;
        RECT 259.950 523.050 262.050 525.150 ;
        RECT 263.250 523.950 264.450 531.300 ;
        RECT 276.000 530.250 279.750 531.300 ;
        RECT 272.100 528.150 273.900 529.950 ;
        RECT 266.100 525.150 267.900 526.950 ;
        RECT 262.950 521.850 265.050 523.950 ;
        RECT 265.950 523.050 268.050 525.150 ;
        RECT 268.950 524.850 271.050 526.950 ;
        RECT 271.950 526.050 274.050 528.150 ;
        RECT 275.850 526.950 277.050 530.250 ;
        RECT 284.100 528.150 285.900 529.950 ;
        RECT 274.950 524.850 277.050 526.950 ;
        RECT 283.950 526.050 286.050 528.150 ;
        RECT 287.400 526.950 288.600 533.400 ;
        RECT 296.850 532.200 298.650 539.250 ;
        RECT 301.350 533.400 303.150 539.250 ;
        RECT 309.150 534.900 310.950 539.250 ;
        RECT 307.650 533.400 310.950 534.900 ;
        RECT 312.150 533.400 313.950 539.250 ;
        RECT 296.850 531.300 300.450 532.200 ;
        RECT 286.950 524.850 289.050 526.950 ;
        RECT 296.100 525.150 297.900 526.950 ;
        RECT 269.100 523.050 270.900 524.850 ;
        RECT 246.150 518.400 247.050 519.300 ;
        RECT 243.450 518.100 245.250 518.400 ;
        RECT 230.550 516.600 231.750 517.500 ;
        RECT 238.950 517.200 245.250 518.100 ;
        RECT 243.450 516.600 245.250 517.200 ;
        RECT 246.150 516.600 248.850 518.400 ;
        RECT 226.950 514.500 231.750 516.600 ;
        RECT 234.150 514.500 241.050 516.300 ;
        RECT 230.550 513.600 231.750 514.500 ;
        RECT 225.150 507.750 226.950 513.600 ;
        RECT 230.250 507.750 232.050 513.600 ;
        RECT 235.050 507.750 236.850 513.600 ;
        RECT 238.050 507.750 239.850 514.500 ;
        RECT 246.150 513.600 250.050 515.700 ;
        RECT 241.950 507.750 243.750 513.600 ;
        RECT 246.150 507.750 247.950 513.600 ;
        RECT 250.650 507.750 252.450 510.600 ;
        RECT 253.650 507.750 255.450 519.600 ;
        RECT 263.250 513.600 264.450 521.850 ;
        RECT 274.950 519.600 276.150 524.850 ;
        RECT 277.950 521.850 280.050 523.950 ;
        RECT 277.950 520.050 279.750 521.850 ;
        RECT 287.400 519.600 288.600 524.850 ;
        RECT 295.950 523.050 298.050 525.150 ;
        RECT 299.250 523.950 300.450 531.300 ;
        RECT 307.650 526.950 308.850 533.400 ;
        RECT 310.950 531.900 312.750 532.500 ;
        RECT 316.650 531.900 318.450 539.250 ;
        RECT 320.850 533.400 322.650 539.250 ;
        RECT 325.350 532.200 327.150 539.250 ;
        RECT 310.950 530.700 318.450 531.900 ;
        RECT 323.550 531.300 327.150 532.200 ;
        RECT 302.100 525.150 303.900 526.950 ;
        RECT 298.950 521.850 301.050 523.950 ;
        RECT 301.950 523.050 304.050 525.150 ;
        RECT 307.650 524.850 310.050 526.950 ;
        RECT 311.100 525.150 312.900 526.950 ;
        RECT 259.650 507.750 261.450 513.600 ;
        RECT 262.650 507.750 264.450 513.600 ;
        RECT 265.650 507.750 267.450 513.600 ;
        RECT 270.300 507.750 272.100 519.600 ;
        RECT 274.500 507.750 276.300 519.600 ;
        RECT 277.800 507.750 279.600 513.600 ;
        RECT 284.550 507.750 286.350 519.600 ;
        RECT 287.550 507.750 289.350 519.600 ;
        RECT 299.250 513.600 300.450 521.850 ;
        RECT 307.650 519.600 308.850 524.850 ;
        RECT 310.950 523.050 313.050 525.150 ;
        RECT 295.650 507.750 297.450 513.600 ;
        RECT 298.650 507.750 300.450 513.600 ;
        RECT 301.650 507.750 303.450 513.600 ;
        RECT 307.050 507.750 308.850 519.600 ;
        RECT 310.050 507.750 311.850 519.600 ;
        RECT 314.100 513.600 315.300 530.700 ;
        RECT 316.950 524.850 319.050 526.950 ;
        RECT 320.100 525.150 321.900 526.950 ;
        RECT 317.100 523.050 318.900 524.850 ;
        RECT 319.950 523.050 322.050 525.150 ;
        RECT 323.550 523.950 324.750 531.300 ;
        RECT 332.700 530.400 334.500 539.250 ;
        RECT 338.100 531.000 339.900 539.250 ;
        RECT 347.550 536.400 349.350 539.250 ;
        RECT 350.550 536.400 352.350 539.250 ;
        RECT 356.550 536.400 358.350 539.250 ;
        RECT 359.550 536.400 361.350 539.250 ;
        RECT 338.100 529.350 342.600 531.000 ;
        RECT 326.100 525.150 327.900 526.950 ;
        RECT 341.400 525.150 342.600 529.350 ;
        RECT 346.950 527.850 349.050 529.950 ;
        RECT 350.400 528.150 351.600 536.400 ;
        RECT 347.100 526.050 348.900 527.850 ;
        RECT 349.950 526.050 352.050 528.150 ;
        RECT 355.950 527.850 358.050 529.950 ;
        RECT 359.400 528.150 360.600 536.400 ;
        RECT 365.550 533.400 367.350 539.250 ;
        RECT 368.850 536.400 370.650 539.250 ;
        RECT 373.350 536.400 375.150 539.250 ;
        RECT 377.550 536.400 379.350 539.250 ;
        RECT 381.450 536.400 383.250 539.250 ;
        RECT 384.750 536.400 386.550 539.250 ;
        RECT 389.250 537.300 391.050 539.250 ;
        RECT 389.250 536.400 393.000 537.300 ;
        RECT 394.050 536.400 395.850 539.250 ;
        RECT 373.650 535.500 374.700 536.400 ;
        RECT 370.950 534.300 374.700 535.500 ;
        RECT 382.200 534.600 383.250 536.400 ;
        RECT 391.950 535.500 393.000 536.400 ;
        RECT 370.950 533.400 373.050 534.300 ;
        RECT 365.550 531.150 366.750 533.400 ;
        RECT 378.150 532.200 379.950 534.000 ;
        RECT 382.200 533.550 387.150 534.600 ;
        RECT 385.350 532.800 387.150 533.550 ;
        RECT 388.650 532.800 390.450 534.600 ;
        RECT 391.950 533.400 394.050 535.500 ;
        RECT 397.050 533.400 398.850 539.250 ;
        RECT 379.050 531.900 379.950 532.200 ;
        RECT 389.100 531.900 390.150 532.800 ;
        RECT 365.550 529.050 370.050 531.150 ;
        RECT 379.050 531.000 390.150 531.900 ;
        RECT 356.100 526.050 357.900 527.850 ;
        RECT 358.950 526.050 361.050 528.150 ;
        RECT 322.950 521.850 325.050 523.950 ;
        RECT 325.950 523.050 328.050 525.150 ;
        RECT 331.950 521.850 334.050 523.950 ;
        RECT 337.950 521.850 340.050 523.950 ;
        RECT 340.950 523.050 343.050 525.150 ;
        RECT 323.550 513.600 324.750 521.850 ;
        RECT 332.100 520.050 333.900 521.850 ;
        RECT 334.950 518.850 337.050 520.950 ;
        RECT 338.250 520.050 340.050 521.850 ;
        RECT 335.100 517.050 336.900 518.850 ;
        RECT 341.700 514.800 342.750 523.050 ;
        RECT 335.700 513.900 342.750 514.800 ;
        RECT 335.700 513.600 337.350 513.900 ;
        RECT 313.650 507.750 315.450 513.600 ;
        RECT 316.650 507.750 318.450 513.600 ;
        RECT 320.550 507.750 322.350 513.600 ;
        RECT 323.550 507.750 325.350 513.600 ;
        RECT 326.550 507.750 328.350 513.600 ;
        RECT 332.550 507.750 334.350 513.600 ;
        RECT 335.550 507.750 337.350 513.600 ;
        RECT 341.550 513.600 342.750 513.900 ;
        RECT 350.400 513.600 351.600 526.050 ;
        RECT 359.400 513.600 360.600 526.050 ;
        RECT 365.550 519.600 366.750 529.050 ;
        RECT 367.950 527.250 371.850 529.050 ;
        RECT 367.950 526.950 370.050 527.250 ;
        RECT 379.050 526.950 379.950 531.000 ;
        RECT 389.100 529.800 390.150 531.000 ;
        RECT 389.100 528.600 396.000 529.800 ;
        RECT 389.100 528.000 390.900 528.600 ;
        RECT 395.100 527.850 396.000 528.600 ;
        RECT 392.100 526.950 393.900 527.700 ;
        RECT 379.050 524.850 382.050 526.950 ;
        RECT 385.950 525.900 393.900 526.950 ;
        RECT 395.100 526.050 396.900 527.850 ;
        RECT 385.950 524.850 388.050 525.900 ;
        RECT 367.950 521.400 369.750 523.200 ;
        RECT 368.850 520.200 373.050 521.400 ;
        RECT 379.050 520.200 379.950 524.850 ;
        RECT 387.750 521.100 389.550 521.400 ;
        RECT 338.550 507.750 340.350 513.000 ;
        RECT 341.550 507.750 343.350 513.600 ;
        RECT 347.550 507.750 349.350 513.600 ;
        RECT 350.550 507.750 352.350 513.600 ;
        RECT 356.550 507.750 358.350 513.600 ;
        RECT 359.550 507.750 361.350 513.600 ;
        RECT 365.550 507.750 367.350 519.600 ;
        RECT 370.950 519.300 373.050 520.200 ;
        RECT 373.950 519.300 379.950 520.200 ;
        RECT 381.150 520.800 389.550 521.100 ;
        RECT 397.950 520.800 398.850 533.400 ;
        RECT 401.550 534.300 403.350 539.250 ;
        RECT 404.550 535.200 406.350 539.250 ;
        RECT 407.550 534.300 409.350 539.250 ;
        RECT 401.550 532.950 409.350 534.300 ;
        RECT 410.550 533.400 412.350 539.250 ;
        RECT 416.550 536.400 418.350 539.250 ;
        RECT 410.550 531.300 411.750 533.400 ;
        RECT 417.150 532.500 418.350 536.400 ;
        RECT 419.850 533.400 421.650 539.250 ;
        RECT 422.850 533.400 424.650 539.250 ;
        RECT 428.850 533.400 430.650 539.250 ;
        RECT 417.150 531.600 422.250 532.500 ;
        RECT 408.000 530.250 411.750 531.300 ;
        RECT 420.000 530.700 422.250 531.600 ;
        RECT 404.100 528.150 405.900 529.950 ;
        RECT 400.950 524.850 403.050 526.950 ;
        RECT 403.950 526.050 406.050 528.150 ;
        RECT 407.850 526.950 409.050 530.250 ;
        RECT 406.950 524.850 409.050 526.950 ;
        RECT 415.950 524.850 418.050 526.950 ;
        RECT 401.100 523.050 402.900 524.850 ;
        RECT 381.150 520.200 398.850 520.800 ;
        RECT 373.950 518.400 374.850 519.300 ;
        RECT 372.150 516.600 374.850 518.400 ;
        RECT 375.750 518.100 377.550 518.400 ;
        RECT 381.150 518.100 382.050 520.200 ;
        RECT 387.750 519.600 398.850 520.200 ;
        RECT 406.950 519.600 408.150 524.850 ;
        RECT 409.950 521.850 412.050 523.950 ;
        RECT 416.100 523.050 417.900 524.850 ;
        RECT 420.000 522.300 421.050 530.700 ;
        RECT 423.150 526.950 424.350 533.400 ;
        RECT 433.350 532.200 435.150 539.250 ;
        RECT 431.550 531.300 435.150 532.200 ;
        RECT 440.550 533.400 442.350 539.250 ;
        RECT 443.850 536.400 445.650 539.250 ;
        RECT 448.350 536.400 450.150 539.250 ;
        RECT 452.550 536.400 454.350 539.250 ;
        RECT 456.450 536.400 458.250 539.250 ;
        RECT 459.750 536.400 461.550 539.250 ;
        RECT 464.250 537.300 466.050 539.250 ;
        RECT 464.250 536.400 468.000 537.300 ;
        RECT 469.050 536.400 470.850 539.250 ;
        RECT 448.650 535.500 449.700 536.400 ;
        RECT 445.950 534.300 449.700 535.500 ;
        RECT 457.200 534.600 458.250 536.400 ;
        RECT 466.950 535.500 468.000 536.400 ;
        RECT 445.950 533.400 448.050 534.300 ;
        RECT 421.950 524.850 424.350 526.950 ;
        RECT 428.100 525.150 429.900 526.950 ;
        RECT 409.950 520.050 411.750 521.850 ;
        RECT 420.000 521.400 422.250 522.300 ;
        RECT 416.550 520.500 422.250 521.400 ;
        RECT 375.750 517.200 382.050 518.100 ;
        RECT 382.950 518.700 384.750 519.300 ;
        RECT 382.950 517.500 390.450 518.700 ;
        RECT 375.750 516.600 377.550 517.200 ;
        RECT 389.250 516.600 390.450 517.500 ;
        RECT 370.950 513.600 374.850 515.700 ;
        RECT 379.950 514.500 386.850 516.300 ;
        RECT 389.250 514.500 394.050 516.600 ;
        RECT 368.550 507.750 370.350 510.600 ;
        RECT 373.050 507.750 374.850 513.600 ;
        RECT 377.250 507.750 379.050 513.600 ;
        RECT 381.150 507.750 382.950 514.500 ;
        RECT 389.250 513.600 390.450 514.500 ;
        RECT 384.150 507.750 385.950 513.600 ;
        RECT 388.950 507.750 390.750 513.600 ;
        RECT 394.050 507.750 395.850 513.600 ;
        RECT 397.050 507.750 398.850 519.600 ;
        RECT 402.300 507.750 404.100 519.600 ;
        RECT 406.500 507.750 408.300 519.600 ;
        RECT 416.550 513.600 417.750 520.500 ;
        RECT 423.150 519.600 424.350 524.850 ;
        RECT 427.950 523.050 430.050 525.150 ;
        RECT 431.550 523.950 432.750 531.300 ;
        RECT 440.550 531.150 441.750 533.400 ;
        RECT 453.150 532.200 454.950 534.000 ;
        RECT 457.200 533.550 462.150 534.600 ;
        RECT 460.350 532.800 462.150 533.550 ;
        RECT 463.650 532.800 465.450 534.600 ;
        RECT 466.950 533.400 469.050 535.500 ;
        RECT 472.050 533.400 473.850 539.250 ;
        RECT 478.650 533.400 480.450 539.250 ;
        RECT 454.050 531.900 454.950 532.200 ;
        RECT 464.100 531.900 465.150 532.800 ;
        RECT 440.550 529.050 445.050 531.150 ;
        RECT 454.050 531.000 465.150 531.900 ;
        RECT 434.100 525.150 435.900 526.950 ;
        RECT 430.950 521.850 433.050 523.950 ;
        RECT 433.950 523.050 436.050 525.150 ;
        RECT 409.800 507.750 411.600 513.600 ;
        RECT 416.550 507.750 418.350 513.600 ;
        RECT 419.850 507.750 421.650 519.600 ;
        RECT 422.850 507.750 424.650 519.600 ;
        RECT 431.550 513.600 432.750 521.850 ;
        RECT 440.550 519.600 441.750 529.050 ;
        RECT 442.950 527.250 446.850 529.050 ;
        RECT 442.950 526.950 445.050 527.250 ;
        RECT 454.050 526.950 454.950 531.000 ;
        RECT 464.100 529.800 465.150 531.000 ;
        RECT 464.100 528.600 471.000 529.800 ;
        RECT 464.100 528.000 465.900 528.600 ;
        RECT 470.100 527.850 471.000 528.600 ;
        RECT 467.100 526.950 468.900 527.700 ;
        RECT 454.050 524.850 457.050 526.950 ;
        RECT 460.950 525.900 468.900 526.950 ;
        RECT 470.100 526.050 471.900 527.850 ;
        RECT 460.950 524.850 463.050 525.900 ;
        RECT 442.950 521.400 444.750 523.200 ;
        RECT 443.850 520.200 448.050 521.400 ;
        RECT 454.050 520.200 454.950 524.850 ;
        RECT 462.750 521.100 464.550 521.400 ;
        RECT 428.550 507.750 430.350 513.600 ;
        RECT 431.550 507.750 433.350 513.600 ;
        RECT 434.550 507.750 436.350 513.600 ;
        RECT 440.550 507.750 442.350 519.600 ;
        RECT 445.950 519.300 448.050 520.200 ;
        RECT 448.950 519.300 454.950 520.200 ;
        RECT 456.150 520.800 464.550 521.100 ;
        RECT 472.950 520.800 473.850 533.400 ;
        RECT 479.250 531.300 480.450 533.400 ;
        RECT 481.650 534.300 483.450 539.250 ;
        RECT 484.650 535.200 486.450 539.250 ;
        RECT 487.650 534.300 489.450 539.250 ;
        RECT 493.650 536.400 495.450 539.250 ;
        RECT 496.650 536.400 498.450 539.250 ;
        RECT 500.550 536.400 502.350 539.250 ;
        RECT 503.550 536.400 505.350 539.250 ;
        RECT 506.550 536.400 508.350 539.250 ;
        RECT 512.550 536.400 514.350 539.250 ;
        RECT 515.550 536.400 517.350 539.250 ;
        RECT 523.650 536.400 525.450 539.250 ;
        RECT 526.650 536.400 528.450 539.250 ;
        RECT 529.650 536.400 531.450 539.250 ;
        RECT 481.650 532.950 489.450 534.300 ;
        RECT 479.250 530.250 483.000 531.300 ;
        RECT 481.950 526.950 483.150 530.250 ;
        RECT 485.100 528.150 486.900 529.950 ;
        RECT 494.400 528.150 495.600 536.400 ;
        RECT 504.000 529.950 505.050 536.400 ;
        RECT 508.950 529.950 511.050 532.050 ;
        RECT 481.950 524.850 484.050 526.950 ;
        RECT 484.950 526.050 487.050 528.150 ;
        RECT 487.950 524.850 490.050 526.950 ;
        RECT 493.950 526.050 496.050 528.150 ;
        RECT 496.950 527.850 499.050 529.950 ;
        RECT 502.950 527.850 505.050 529.950 ;
        RECT 497.100 526.050 498.900 527.850 ;
        RECT 478.950 521.850 481.050 523.950 ;
        RECT 456.150 520.200 473.850 520.800 ;
        RECT 448.950 518.400 449.850 519.300 ;
        RECT 447.150 516.600 449.850 518.400 ;
        RECT 450.750 518.100 452.550 518.400 ;
        RECT 456.150 518.100 457.050 520.200 ;
        RECT 462.750 519.600 473.850 520.200 ;
        RECT 479.250 520.050 481.050 521.850 ;
        RECT 482.850 519.600 484.050 524.850 ;
        RECT 488.100 523.050 489.900 524.850 ;
        RECT 450.750 517.200 457.050 518.100 ;
        RECT 457.950 518.700 459.750 519.300 ;
        RECT 457.950 517.500 465.450 518.700 ;
        RECT 450.750 516.600 452.550 517.200 ;
        RECT 464.250 516.600 465.450 517.500 ;
        RECT 445.950 513.600 449.850 515.700 ;
        RECT 454.950 514.500 461.850 516.300 ;
        RECT 464.250 514.500 469.050 516.600 ;
        RECT 443.550 507.750 445.350 510.600 ;
        RECT 448.050 507.750 449.850 513.600 ;
        RECT 452.250 507.750 454.050 513.600 ;
        RECT 456.150 507.750 457.950 514.500 ;
        RECT 464.250 513.600 465.450 514.500 ;
        RECT 459.150 507.750 460.950 513.600 ;
        RECT 463.950 507.750 465.750 513.600 ;
        RECT 469.050 507.750 470.850 513.600 ;
        RECT 472.050 507.750 473.850 519.600 ;
        RECT 479.400 507.750 481.200 513.600 ;
        RECT 482.700 507.750 484.500 519.600 ;
        RECT 486.900 507.750 488.700 519.600 ;
        RECT 494.400 513.600 495.600 526.050 ;
        RECT 499.950 524.850 502.050 526.950 ;
        RECT 500.100 523.050 501.900 524.850 ;
        RECT 504.000 520.650 505.050 527.850 ;
        RECT 505.950 524.850 508.050 526.950 ;
        RECT 506.100 523.050 507.900 524.850 ;
        RECT 509.550 522.450 510.450 529.950 ;
        RECT 511.950 527.850 514.050 529.950 ;
        RECT 515.400 528.150 516.600 536.400 ;
        RECT 526.950 529.950 528.000 536.400 ;
        RECT 534.000 533.400 535.800 539.250 ;
        RECT 538.200 535.050 540.000 539.250 ;
        RECT 541.500 536.400 543.300 539.250 ;
        RECT 548.550 536.400 550.350 539.250 ;
        RECT 551.550 536.400 553.350 539.250 ;
        RECT 554.550 536.400 556.350 539.250 ;
        RECT 538.200 533.400 543.900 535.050 ;
        RECT 512.100 526.050 513.900 527.850 ;
        RECT 514.950 526.050 517.050 528.150 ;
        RECT 526.950 527.850 529.050 529.950 ;
        RECT 533.100 528.150 534.900 529.950 ;
        RECT 511.950 522.450 514.050 523.050 ;
        RECT 509.550 521.550 514.050 522.450 ;
        RECT 511.950 520.950 514.050 521.550 ;
        RECT 504.000 519.600 506.550 520.650 ;
        RECT 493.650 507.750 495.450 513.600 ;
        RECT 496.650 507.750 498.450 513.600 ;
        RECT 500.550 507.750 502.350 519.600 ;
        RECT 504.750 507.750 506.550 519.600 ;
        RECT 515.400 513.600 516.600 526.050 ;
        RECT 523.950 524.850 526.050 526.950 ;
        RECT 524.100 523.050 525.900 524.850 ;
        RECT 526.950 520.650 528.000 527.850 ;
        RECT 529.950 524.850 532.050 526.950 ;
        RECT 532.950 526.050 535.050 528.150 ;
        RECT 535.950 527.850 538.050 529.950 ;
        RECT 539.100 528.150 540.900 529.950 ;
        RECT 536.100 526.050 537.900 527.850 ;
        RECT 538.950 526.050 541.050 528.150 ;
        RECT 542.700 526.950 543.900 533.400 ;
        RECT 552.450 532.200 553.350 536.400 ;
        RECT 557.550 533.400 559.350 539.250 ;
        RECT 568.800 533.400 570.600 539.250 ;
        RECT 573.000 533.400 574.800 539.250 ;
        RECT 577.200 533.400 579.000 539.250 ;
        RECT 552.450 531.300 555.750 532.200 ;
        RECT 553.950 530.400 555.750 531.300 ;
        RECT 547.950 527.850 550.050 529.950 ;
        RECT 541.950 524.850 544.050 526.950 ;
        RECT 548.100 526.050 549.900 527.850 ;
        RECT 550.950 524.850 553.050 526.950 ;
        RECT 530.100 523.050 531.900 524.850 ;
        RECT 525.450 519.600 528.000 520.650 ;
        RECT 542.700 519.600 543.900 524.850 ;
        RECT 551.100 523.050 552.900 524.850 ;
        RECT 554.700 522.150 555.600 530.400 ;
        RECT 558.000 528.150 559.050 533.400 ;
        RECT 569.250 528.150 571.050 529.950 ;
        RECT 556.950 526.050 559.050 528.150 ;
        RECT 553.950 522.000 555.750 522.150 ;
        RECT 548.550 520.800 555.750 522.000 ;
        RECT 548.550 519.600 549.750 520.800 ;
        RECT 553.950 520.350 555.750 520.800 ;
        RECT 512.550 507.750 514.350 513.600 ;
        RECT 515.550 507.750 517.350 513.600 ;
        RECT 525.450 507.750 527.250 519.600 ;
        RECT 529.650 507.750 531.450 519.600 ;
        RECT 533.550 518.700 541.350 519.600 ;
        RECT 533.550 507.750 535.350 518.700 ;
        RECT 536.550 507.750 538.350 517.800 ;
        RECT 539.550 507.750 541.350 518.700 ;
        RECT 542.550 507.750 544.350 519.600 ;
        RECT 548.550 507.750 550.350 519.600 ;
        RECT 557.100 519.450 558.450 526.050 ;
        RECT 565.950 524.850 568.050 526.950 ;
        RECT 568.950 526.050 571.050 528.150 ;
        RECT 573.000 526.950 574.050 533.400 ;
        RECT 584.850 532.200 586.650 539.250 ;
        RECT 589.350 533.400 591.150 539.250 ;
        RECT 593.550 533.400 595.350 539.250 ;
        RECT 596.850 536.400 598.650 539.250 ;
        RECT 601.350 536.400 603.150 539.250 ;
        RECT 605.550 536.400 607.350 539.250 ;
        RECT 609.450 536.400 611.250 539.250 ;
        RECT 612.750 536.400 614.550 539.250 ;
        RECT 617.250 537.300 619.050 539.250 ;
        RECT 617.250 536.400 621.000 537.300 ;
        RECT 622.050 536.400 623.850 539.250 ;
        RECT 601.650 535.500 602.700 536.400 ;
        RECT 598.950 534.300 602.700 535.500 ;
        RECT 610.200 534.600 611.250 536.400 ;
        RECT 619.950 535.500 621.000 536.400 ;
        RECT 598.950 533.400 601.050 534.300 ;
        RECT 584.850 531.300 588.450 532.200 ;
        RECT 571.950 524.850 574.050 526.950 ;
        RECT 574.950 528.150 576.750 529.950 ;
        RECT 574.950 526.050 577.050 528.150 ;
        RECT 577.950 524.850 580.050 526.950 ;
        RECT 584.100 525.150 585.900 526.950 ;
        RECT 566.100 523.050 567.900 524.850 ;
        RECT 571.950 521.400 572.850 524.850 ;
        RECT 577.950 523.050 579.750 524.850 ;
        RECT 583.950 523.050 586.050 525.150 ;
        RECT 587.250 523.950 588.450 531.300 ;
        RECT 593.550 531.150 594.750 533.400 ;
        RECT 606.150 532.200 607.950 534.000 ;
        RECT 610.200 533.550 615.150 534.600 ;
        RECT 613.350 532.800 615.150 533.550 ;
        RECT 616.650 532.800 618.450 534.600 ;
        RECT 619.950 533.400 622.050 535.500 ;
        RECT 625.050 533.400 626.850 539.250 ;
        RECT 607.050 531.900 607.950 532.200 ;
        RECT 617.100 531.900 618.150 532.800 ;
        RECT 593.550 529.050 598.050 531.150 ;
        RECT 607.050 531.000 618.150 531.900 ;
        RECT 590.100 525.150 591.900 526.950 ;
        RECT 586.950 521.850 589.050 523.950 ;
        RECT 589.950 523.050 592.050 525.150 ;
        RECT 568.800 520.500 572.850 521.400 ;
        RECT 568.800 519.600 570.600 520.500 ;
        RECT 553.050 507.750 554.850 519.450 ;
        RECT 556.050 518.100 558.450 519.450 ;
        RECT 556.050 507.750 557.850 518.100 ;
        RECT 565.650 508.500 567.450 519.600 ;
        RECT 568.650 509.400 570.450 519.600 ;
        RECT 571.650 518.400 579.450 519.300 ;
        RECT 571.650 508.500 573.450 518.400 ;
        RECT 565.650 507.750 573.450 508.500 ;
        RECT 574.650 507.750 576.450 517.500 ;
        RECT 577.650 507.750 579.450 518.400 ;
        RECT 587.250 513.600 588.450 521.850 ;
        RECT 593.550 519.600 594.750 529.050 ;
        RECT 595.950 527.250 599.850 529.050 ;
        RECT 595.950 526.950 598.050 527.250 ;
        RECT 607.050 526.950 607.950 531.000 ;
        RECT 617.100 529.800 618.150 531.000 ;
        RECT 617.100 528.600 624.000 529.800 ;
        RECT 617.100 528.000 618.900 528.600 ;
        RECT 623.100 527.850 624.000 528.600 ;
        RECT 620.100 526.950 621.900 527.700 ;
        RECT 607.050 524.850 610.050 526.950 ;
        RECT 613.950 525.900 621.900 526.950 ;
        RECT 623.100 526.050 624.900 527.850 ;
        RECT 613.950 524.850 616.050 525.900 ;
        RECT 595.950 521.400 597.750 523.200 ;
        RECT 596.850 520.200 601.050 521.400 ;
        RECT 607.050 520.200 607.950 524.850 ;
        RECT 615.750 521.100 617.550 521.400 ;
        RECT 583.650 507.750 585.450 513.600 ;
        RECT 586.650 507.750 588.450 513.600 ;
        RECT 589.650 507.750 591.450 513.600 ;
        RECT 593.550 507.750 595.350 519.600 ;
        RECT 598.950 519.300 601.050 520.200 ;
        RECT 601.950 519.300 607.950 520.200 ;
        RECT 609.150 520.800 617.550 521.100 ;
        RECT 625.950 520.800 626.850 533.400 ;
        RECT 609.150 520.200 626.850 520.800 ;
        RECT 601.950 518.400 602.850 519.300 ;
        RECT 600.150 516.600 602.850 518.400 ;
        RECT 603.750 518.100 605.550 518.400 ;
        RECT 609.150 518.100 610.050 520.200 ;
        RECT 615.750 519.600 626.850 520.200 ;
        RECT 603.750 517.200 610.050 518.100 ;
        RECT 610.950 518.700 612.750 519.300 ;
        RECT 610.950 517.500 618.450 518.700 ;
        RECT 603.750 516.600 605.550 517.200 ;
        RECT 617.250 516.600 618.450 517.500 ;
        RECT 598.950 513.600 602.850 515.700 ;
        RECT 607.950 514.500 614.850 516.300 ;
        RECT 617.250 514.500 622.050 516.600 ;
        RECT 596.550 507.750 598.350 510.600 ;
        RECT 601.050 507.750 602.850 513.600 ;
        RECT 605.250 507.750 607.050 513.600 ;
        RECT 609.150 507.750 610.950 514.500 ;
        RECT 617.250 513.600 618.450 514.500 ;
        RECT 612.150 507.750 613.950 513.600 ;
        RECT 616.950 507.750 618.750 513.600 ;
        RECT 622.050 507.750 623.850 513.600 ;
        RECT 625.050 507.750 626.850 519.600 ;
        RECT 629.550 533.400 631.350 539.250 ;
        RECT 632.850 536.400 634.650 539.250 ;
        RECT 637.350 536.400 639.150 539.250 ;
        RECT 641.550 536.400 643.350 539.250 ;
        RECT 645.450 536.400 647.250 539.250 ;
        RECT 648.750 536.400 650.550 539.250 ;
        RECT 653.250 537.300 655.050 539.250 ;
        RECT 653.250 536.400 657.000 537.300 ;
        RECT 658.050 536.400 659.850 539.250 ;
        RECT 637.650 535.500 638.700 536.400 ;
        RECT 634.950 534.300 638.700 535.500 ;
        RECT 646.200 534.600 647.250 536.400 ;
        RECT 655.950 535.500 657.000 536.400 ;
        RECT 634.950 533.400 637.050 534.300 ;
        RECT 629.550 531.150 630.750 533.400 ;
        RECT 642.150 532.200 643.950 534.000 ;
        RECT 646.200 533.550 651.150 534.600 ;
        RECT 649.350 532.800 651.150 533.550 ;
        RECT 652.650 532.800 654.450 534.600 ;
        RECT 655.950 533.400 658.050 535.500 ;
        RECT 661.050 533.400 662.850 539.250 ;
        RECT 667.650 533.400 669.450 539.250 ;
        RECT 670.650 533.400 672.450 539.250 ;
        RECT 673.650 533.400 675.450 539.250 ;
        RECT 676.650 533.400 678.450 539.250 ;
        RECT 679.650 533.400 681.450 539.250 ;
        RECT 643.050 531.900 643.950 532.200 ;
        RECT 653.100 531.900 654.150 532.800 ;
        RECT 629.550 529.050 634.050 531.150 ;
        RECT 643.050 531.000 654.150 531.900 ;
        RECT 629.550 519.600 630.750 529.050 ;
        RECT 631.950 527.250 635.850 529.050 ;
        RECT 631.950 526.950 634.050 527.250 ;
        RECT 643.050 526.950 643.950 531.000 ;
        RECT 653.100 529.800 654.150 531.000 ;
        RECT 653.100 528.600 660.000 529.800 ;
        RECT 653.100 528.000 654.900 528.600 ;
        RECT 659.100 527.850 660.000 528.600 ;
        RECT 656.100 526.950 657.900 527.700 ;
        RECT 643.050 524.850 646.050 526.950 ;
        RECT 649.950 525.900 657.900 526.950 ;
        RECT 659.100 526.050 660.900 527.850 ;
        RECT 649.950 524.850 652.050 525.900 ;
        RECT 631.950 521.400 633.750 523.200 ;
        RECT 632.850 520.200 637.050 521.400 ;
        RECT 643.050 520.200 643.950 524.850 ;
        RECT 651.750 521.100 653.550 521.400 ;
        RECT 629.550 507.750 631.350 519.600 ;
        RECT 634.950 519.300 637.050 520.200 ;
        RECT 637.950 519.300 643.950 520.200 ;
        RECT 645.150 520.800 653.550 521.100 ;
        RECT 661.950 520.800 662.850 533.400 ;
        RECT 670.800 532.500 672.600 533.400 ;
        RECT 676.800 532.500 678.600 533.400 ;
        RECT 682.650 532.500 684.450 539.250 ;
        RECT 685.650 533.400 687.450 539.250 ;
        RECT 688.650 533.400 690.450 539.250 ;
        RECT 691.650 533.400 693.450 539.250 ;
        RECT 695.550 534.300 697.350 539.250 ;
        RECT 698.550 535.200 700.350 539.250 ;
        RECT 701.550 534.300 703.350 539.250 ;
        RECT 688.800 532.500 690.600 533.400 ;
        RECT 695.550 532.950 703.350 534.300 ;
        RECT 704.550 533.400 706.350 539.250 ;
        RECT 669.900 532.350 672.600 532.500 ;
        RECT 669.750 531.300 672.600 532.350 ;
        RECT 674.700 531.300 678.600 532.500 ;
        RECT 680.700 531.300 684.450 532.500 ;
        RECT 686.550 531.300 690.600 532.500 ;
        RECT 704.550 531.300 705.750 533.400 ;
        RECT 669.750 528.150 670.800 531.300 ;
        RECT 674.700 530.400 675.900 531.300 ;
        RECT 680.700 530.400 681.900 531.300 ;
        RECT 686.550 530.400 687.750 531.300 ;
        RECT 671.700 528.600 675.900 530.400 ;
        RECT 677.700 528.600 681.900 530.400 ;
        RECT 683.700 528.600 687.750 530.400 ;
        RECT 702.000 530.250 705.750 531.300 ;
        RECT 667.950 526.050 670.800 528.150 ;
        RECT 645.150 520.200 662.850 520.800 ;
        RECT 669.750 521.700 670.800 526.050 ;
        RECT 674.700 521.700 675.900 528.600 ;
        RECT 680.700 521.700 681.900 528.600 ;
        RECT 686.550 521.700 687.750 528.600 ;
        RECT 689.100 528.150 690.900 529.950 ;
        RECT 698.100 528.150 699.900 529.950 ;
        RECT 688.950 526.050 691.050 528.150 ;
        RECT 694.950 524.850 697.050 526.950 ;
        RECT 697.950 526.050 700.050 528.150 ;
        RECT 701.850 526.950 703.050 530.250 ;
        RECT 700.950 524.850 703.050 526.950 ;
        RECT 695.100 523.050 696.900 524.850 ;
        RECT 669.750 520.500 672.450 521.700 ;
        RECT 674.700 520.500 678.450 521.700 ;
        RECT 680.700 520.500 684.450 521.700 ;
        RECT 686.550 520.500 690.450 521.700 ;
        RECT 637.950 518.400 638.850 519.300 ;
        RECT 636.150 516.600 638.850 518.400 ;
        RECT 639.750 518.100 641.550 518.400 ;
        RECT 645.150 518.100 646.050 520.200 ;
        RECT 651.750 519.600 662.850 520.200 ;
        RECT 639.750 517.200 646.050 518.100 ;
        RECT 646.950 518.700 648.750 519.300 ;
        RECT 646.950 517.500 654.450 518.700 ;
        RECT 639.750 516.600 641.550 517.200 ;
        RECT 653.250 516.600 654.450 517.500 ;
        RECT 634.950 513.600 638.850 515.700 ;
        RECT 643.950 514.500 650.850 516.300 ;
        RECT 653.250 514.500 658.050 516.600 ;
        RECT 632.550 507.750 634.350 510.600 ;
        RECT 637.050 507.750 638.850 513.600 ;
        RECT 641.250 507.750 643.050 513.600 ;
        RECT 645.150 507.750 646.950 514.500 ;
        RECT 653.250 513.600 654.450 514.500 ;
        RECT 648.150 507.750 649.950 513.600 ;
        RECT 652.950 507.750 654.750 513.600 ;
        RECT 658.050 507.750 659.850 513.600 ;
        RECT 661.050 507.750 662.850 519.600 ;
        RECT 667.650 507.750 669.450 519.600 ;
        RECT 670.650 507.750 672.450 520.500 ;
        RECT 673.650 507.750 675.450 519.600 ;
        RECT 676.650 507.750 678.450 520.500 ;
        RECT 679.650 507.750 681.450 519.600 ;
        RECT 682.650 507.750 684.450 520.500 ;
        RECT 685.650 507.750 687.450 519.600 ;
        RECT 688.650 507.750 690.450 520.500 ;
        RECT 700.950 519.600 702.150 524.850 ;
        RECT 703.950 521.850 706.050 523.950 ;
        RECT 703.950 520.050 705.750 521.850 ;
        RECT 691.650 507.750 693.450 519.600 ;
        RECT 696.300 507.750 698.100 519.600 ;
        RECT 700.500 507.750 702.300 519.600 ;
        RECT 703.800 507.750 705.600 513.600 ;
        RECT 3.150 491.400 4.950 503.250 ;
        RECT 6.150 497.400 7.950 503.250 ;
        RECT 11.250 497.400 13.050 503.250 ;
        RECT 16.050 497.400 17.850 503.250 ;
        RECT 11.550 496.500 12.750 497.400 ;
        RECT 19.050 496.500 20.850 503.250 ;
        RECT 22.950 497.400 24.750 503.250 ;
        RECT 27.150 497.400 28.950 503.250 ;
        RECT 31.650 500.400 33.450 503.250 ;
        RECT 7.950 494.400 12.750 496.500 ;
        RECT 15.150 494.700 22.050 496.500 ;
        RECT 27.150 495.300 31.050 497.400 ;
        RECT 11.550 493.500 12.750 494.400 ;
        RECT 24.450 493.800 26.250 494.400 ;
        RECT 11.550 492.300 19.050 493.500 ;
        RECT 17.250 491.700 19.050 492.300 ;
        RECT 19.950 492.900 26.250 493.800 ;
        RECT 3.150 490.800 14.250 491.400 ;
        RECT 19.950 490.800 20.850 492.900 ;
        RECT 24.450 492.600 26.250 492.900 ;
        RECT 27.150 492.600 29.850 494.400 ;
        RECT 27.150 491.700 28.050 492.600 ;
        RECT 3.150 490.200 20.850 490.800 ;
        RECT 3.150 477.600 4.050 490.200 ;
        RECT 12.450 489.900 20.850 490.200 ;
        RECT 22.050 490.800 28.050 491.700 ;
        RECT 28.950 490.800 31.050 491.700 ;
        RECT 34.650 491.400 36.450 503.250 ;
        RECT 40.650 502.500 48.450 503.250 ;
        RECT 40.650 491.400 42.450 502.500 ;
        RECT 43.650 491.400 45.450 501.600 ;
        RECT 46.650 492.600 48.450 502.500 ;
        RECT 49.650 493.500 51.450 503.250 ;
        RECT 52.650 492.600 54.450 503.250 ;
        RECT 58.650 497.400 60.450 503.250 ;
        RECT 61.650 497.400 63.450 503.250 ;
        RECT 64.650 497.400 66.450 503.250 ;
        RECT 58.950 493.950 61.050 496.050 ;
        RECT 46.650 491.700 54.450 492.600 ;
        RECT 59.550 492.450 60.450 493.950 ;
        RECT 56.550 491.550 60.450 492.450 ;
        RECT 12.450 489.600 14.250 489.900 ;
        RECT 22.050 486.150 22.950 490.800 ;
        RECT 28.950 489.600 33.150 490.800 ;
        RECT 32.250 487.800 34.050 489.600 ;
        RECT 13.950 485.100 16.050 486.150 ;
        RECT 5.100 483.150 6.900 484.950 ;
        RECT 8.100 484.050 16.050 485.100 ;
        RECT 19.950 484.050 22.950 486.150 ;
        RECT 8.100 483.300 9.900 484.050 ;
        RECT 6.000 482.400 6.900 483.150 ;
        RECT 11.100 482.400 12.900 483.000 ;
        RECT 6.000 481.200 12.900 482.400 ;
        RECT 11.850 480.000 12.900 481.200 ;
        RECT 22.050 480.000 22.950 484.050 ;
        RECT 31.950 483.750 34.050 484.050 ;
        RECT 30.150 481.950 34.050 483.750 ;
        RECT 35.250 481.950 36.450 491.400 ;
        RECT 43.800 490.500 45.600 491.400 ;
        RECT 43.800 489.600 47.850 490.500 ;
        RECT 41.100 486.150 42.900 487.950 ;
        RECT 46.950 486.150 47.850 489.600 ;
        RECT 52.950 486.150 54.750 487.950 ;
        RECT 40.950 484.050 43.050 486.150 ;
        RECT 43.950 482.850 46.050 484.950 ;
        RECT 46.950 484.050 49.050 486.150 ;
        RECT 11.850 479.100 22.950 480.000 ;
        RECT 31.950 479.850 36.450 481.950 ;
        RECT 44.250 481.050 46.050 482.850 ;
        RECT 11.850 478.200 12.900 479.100 ;
        RECT 22.050 478.800 22.950 479.100 ;
        RECT 3.150 471.750 4.950 477.600 ;
        RECT 7.950 475.500 10.050 477.600 ;
        RECT 11.550 476.400 13.350 478.200 ;
        RECT 14.850 477.450 16.650 478.200 ;
        RECT 14.850 476.400 19.800 477.450 ;
        RECT 22.050 477.000 23.850 478.800 ;
        RECT 35.250 477.600 36.450 479.850 ;
        RECT 48.000 477.600 49.050 484.050 ;
        RECT 49.950 482.850 52.050 484.950 ;
        RECT 52.950 484.050 55.050 486.150 ;
        RECT 56.550 484.050 57.450 491.550 ;
        RECT 62.250 489.150 63.450 497.400 ;
        RECT 68.550 491.400 70.350 503.250 ;
        RECT 71.550 500.400 73.350 503.250 ;
        RECT 76.050 497.400 77.850 503.250 ;
        RECT 80.250 497.400 82.050 503.250 ;
        RECT 73.950 495.300 77.850 497.400 ;
        RECT 84.150 496.500 85.950 503.250 ;
        RECT 87.150 497.400 88.950 503.250 ;
        RECT 91.950 497.400 93.750 503.250 ;
        RECT 97.050 497.400 98.850 503.250 ;
        RECT 92.250 496.500 93.450 497.400 ;
        RECT 82.950 494.700 89.850 496.500 ;
        RECT 92.250 494.400 97.050 496.500 ;
        RECT 75.150 492.600 77.850 494.400 ;
        RECT 78.750 493.800 80.550 494.400 ;
        RECT 78.750 492.900 85.050 493.800 ;
        RECT 92.250 493.500 93.450 494.400 ;
        RECT 78.750 492.600 80.550 492.900 ;
        RECT 76.950 491.700 77.850 492.600 ;
        RECT 58.950 485.850 61.050 487.950 ;
        RECT 61.950 487.050 64.050 489.150 ;
        RECT 59.100 484.050 60.900 485.850 ;
        RECT 49.950 481.050 51.750 482.850 ;
        RECT 55.950 481.950 58.050 484.050 ;
        RECT 62.250 479.700 63.450 487.050 ;
        RECT 64.950 485.850 67.050 487.950 ;
        RECT 65.100 484.050 66.900 485.850 ;
        RECT 59.850 478.800 63.450 479.700 ;
        RECT 68.550 481.950 69.750 491.400 ;
        RECT 73.950 490.800 76.050 491.700 ;
        RECT 76.950 490.800 82.950 491.700 ;
        RECT 71.850 489.600 76.050 490.800 ;
        RECT 70.950 487.800 72.750 489.600 ;
        RECT 82.050 486.150 82.950 490.800 ;
        RECT 84.150 490.800 85.050 492.900 ;
        RECT 85.950 492.300 93.450 493.500 ;
        RECT 85.950 491.700 87.750 492.300 ;
        RECT 100.050 491.400 101.850 503.250 ;
        RECT 107.400 497.400 109.200 503.250 ;
        RECT 110.700 491.400 112.500 503.250 ;
        RECT 114.900 491.400 116.700 503.250 ;
        RECT 121.650 502.500 129.450 503.250 ;
        RECT 121.650 491.400 123.450 502.500 ;
        RECT 124.650 491.400 126.450 501.600 ;
        RECT 127.650 492.600 129.450 502.500 ;
        RECT 130.650 493.500 132.450 503.250 ;
        RECT 133.650 492.600 135.450 503.250 ;
        RECT 137.550 497.400 139.350 503.250 ;
        RECT 140.550 497.400 142.350 503.250 ;
        RECT 143.550 497.400 145.350 503.250 ;
        RECT 151.650 497.400 153.450 503.250 ;
        RECT 154.650 498.000 156.450 503.250 ;
        RECT 127.650 491.700 135.450 492.600 ;
        RECT 90.750 490.800 101.850 491.400 ;
        RECT 84.150 490.200 101.850 490.800 ;
        RECT 84.150 489.900 92.550 490.200 ;
        RECT 90.750 489.600 92.550 489.900 ;
        RECT 82.050 484.050 85.050 486.150 ;
        RECT 88.950 485.100 91.050 486.150 ;
        RECT 88.950 484.050 96.900 485.100 ;
        RECT 70.950 483.750 73.050 484.050 ;
        RECT 70.950 481.950 74.850 483.750 ;
        RECT 68.550 479.850 73.050 481.950 ;
        RECT 82.050 480.000 82.950 484.050 ;
        RECT 95.100 483.300 96.900 484.050 ;
        RECT 98.100 483.150 99.900 484.950 ;
        RECT 92.100 482.400 93.900 483.000 ;
        RECT 98.100 482.400 99.000 483.150 ;
        RECT 92.100 481.200 99.000 482.400 ;
        RECT 92.100 480.000 93.150 481.200 ;
        RECT 28.950 476.700 31.050 477.600 ;
        RECT 9.000 474.600 10.050 475.500 ;
        RECT 18.750 474.600 19.800 476.400 ;
        RECT 27.300 475.500 31.050 476.700 ;
        RECT 27.300 474.600 28.350 475.500 ;
        RECT 6.150 471.750 7.950 474.600 ;
        RECT 9.000 473.700 12.750 474.600 ;
        RECT 10.950 471.750 12.750 473.700 ;
        RECT 15.450 471.750 17.250 474.600 ;
        RECT 18.750 471.750 20.550 474.600 ;
        RECT 22.650 471.750 24.450 474.600 ;
        RECT 26.850 471.750 28.650 474.600 ;
        RECT 31.350 471.750 33.150 474.600 ;
        RECT 34.650 471.750 36.450 477.600 ;
        RECT 43.800 471.750 45.600 477.600 ;
        RECT 48.000 471.750 49.800 477.600 ;
        RECT 52.200 471.750 54.000 477.600 ;
        RECT 59.850 471.750 61.650 478.800 ;
        RECT 68.550 477.600 69.750 479.850 ;
        RECT 82.050 479.100 93.150 480.000 ;
        RECT 82.050 478.800 82.950 479.100 ;
        RECT 64.350 471.750 66.150 477.600 ;
        RECT 68.550 471.750 70.350 477.600 ;
        RECT 73.950 476.700 76.050 477.600 ;
        RECT 81.150 477.000 82.950 478.800 ;
        RECT 92.100 478.200 93.150 479.100 ;
        RECT 88.350 477.450 90.150 478.200 ;
        RECT 73.950 475.500 77.700 476.700 ;
        RECT 76.650 474.600 77.700 475.500 ;
        RECT 85.200 476.400 90.150 477.450 ;
        RECT 91.650 476.400 93.450 478.200 ;
        RECT 100.950 477.600 101.850 490.200 ;
        RECT 107.250 489.150 109.050 490.950 ;
        RECT 106.950 487.050 109.050 489.150 ;
        RECT 110.850 486.150 112.050 491.400 ;
        RECT 124.800 490.500 126.600 491.400 ;
        RECT 124.800 489.600 128.850 490.500 ;
        RECT 116.100 486.150 117.900 487.950 ;
        RECT 122.100 486.150 123.900 487.950 ;
        RECT 127.950 486.150 128.850 489.600 ;
        RECT 140.550 489.150 141.750 497.400 ;
        RECT 152.250 497.100 153.450 497.400 ;
        RECT 157.650 497.400 159.450 503.250 ;
        RECT 160.650 497.400 162.450 503.250 ;
        RECT 157.650 497.100 159.300 497.400 ;
        RECT 152.250 496.200 159.300 497.100 ;
        RECT 133.950 486.150 135.750 487.950 ;
        RECT 109.950 484.050 112.050 486.150 ;
        RECT 109.950 480.750 111.150 484.050 ;
        RECT 112.950 482.850 115.050 484.950 ;
        RECT 115.950 484.050 118.050 486.150 ;
        RECT 121.950 484.050 124.050 486.150 ;
        RECT 124.950 482.850 127.050 484.950 ;
        RECT 127.950 484.050 130.050 486.150 ;
        RECT 113.100 481.050 114.900 482.850 ;
        RECT 125.250 481.050 127.050 482.850 ;
        RECT 107.250 479.700 111.000 480.750 ;
        RECT 107.250 477.600 108.450 479.700 ;
        RECT 85.200 474.600 86.250 476.400 ;
        RECT 94.950 475.500 97.050 477.600 ;
        RECT 94.950 474.600 96.000 475.500 ;
        RECT 71.850 471.750 73.650 474.600 ;
        RECT 76.350 471.750 78.150 474.600 ;
        RECT 80.550 471.750 82.350 474.600 ;
        RECT 84.450 471.750 86.250 474.600 ;
        RECT 87.750 471.750 89.550 474.600 ;
        RECT 92.250 473.700 96.000 474.600 ;
        RECT 92.250 471.750 94.050 473.700 ;
        RECT 97.050 471.750 98.850 474.600 ;
        RECT 100.050 471.750 101.850 477.600 ;
        RECT 106.650 471.750 108.450 477.600 ;
        RECT 109.650 476.700 117.450 478.050 ;
        RECT 129.000 477.600 130.050 484.050 ;
        RECT 130.950 482.850 133.050 484.950 ;
        RECT 133.950 484.050 136.050 486.150 ;
        RECT 136.950 485.850 139.050 487.950 ;
        RECT 139.950 487.050 142.050 489.150 ;
        RECT 152.250 487.950 153.300 496.200 ;
        RECT 158.100 492.150 159.900 493.950 ;
        RECT 154.950 489.150 156.750 490.950 ;
        RECT 157.950 490.050 160.050 492.150 ;
        RECT 166.050 491.400 167.850 503.250 ;
        RECT 169.050 491.400 170.850 503.250 ;
        RECT 172.650 497.400 174.450 503.250 ;
        RECT 175.650 497.400 177.450 503.250 ;
        RECT 179.550 497.400 181.350 503.250 ;
        RECT 182.550 497.400 184.350 503.250 ;
        RECT 185.550 498.000 187.350 503.250 ;
        RECT 161.100 489.150 162.900 490.950 ;
        RECT 137.100 484.050 138.900 485.850 ;
        RECT 130.950 481.050 132.750 482.850 ;
        RECT 140.550 479.700 141.750 487.050 ;
        RECT 142.950 485.850 145.050 487.950 ;
        RECT 151.950 485.850 154.050 487.950 ;
        RECT 154.950 487.050 157.050 489.150 ;
        RECT 160.950 487.050 163.050 489.150 ;
        RECT 166.650 486.150 167.850 491.400 ;
        RECT 143.100 484.050 144.900 485.850 ;
        RECT 152.400 481.650 153.600 485.850 ;
        RECT 166.650 484.050 169.050 486.150 ;
        RECT 169.950 485.850 172.050 487.950 ;
        RECT 170.100 484.050 171.900 485.850 ;
        RECT 152.400 480.000 156.900 481.650 ;
        RECT 140.550 478.800 144.150 479.700 ;
        RECT 109.650 471.750 111.450 476.700 ;
        RECT 112.650 471.750 114.450 475.800 ;
        RECT 115.650 471.750 117.450 476.700 ;
        RECT 124.800 471.750 126.600 477.600 ;
        RECT 129.000 471.750 130.800 477.600 ;
        RECT 133.200 471.750 135.000 477.600 ;
        RECT 137.850 471.750 139.650 477.600 ;
        RECT 142.350 471.750 144.150 478.800 ;
        RECT 155.100 471.750 156.900 480.000 ;
        RECT 160.500 471.750 162.300 480.600 ;
        RECT 166.650 477.600 167.850 484.050 ;
        RECT 173.100 480.300 174.300 497.400 ;
        RECT 182.700 497.100 184.350 497.400 ;
        RECT 188.550 497.400 190.350 503.250 ;
        RECT 188.550 497.100 189.750 497.400 ;
        RECT 182.700 496.200 189.750 497.100 ;
        RECT 182.100 492.150 183.900 493.950 ;
        RECT 179.100 489.150 180.900 490.950 ;
        RECT 181.950 490.050 184.050 492.150 ;
        RECT 185.250 489.150 187.050 490.950 ;
        RECT 176.100 486.150 177.900 487.950 ;
        RECT 178.950 487.050 181.050 489.150 ;
        RECT 184.950 487.050 187.050 489.150 ;
        RECT 188.700 487.950 189.750 496.200 ;
        RECT 195.300 491.400 197.100 503.250 ;
        RECT 199.500 491.400 201.300 503.250 ;
        RECT 202.800 497.400 204.600 503.250 ;
        RECT 209.550 497.400 211.350 503.250 ;
        RECT 212.550 497.400 214.350 503.250 ;
        RECT 215.550 497.400 217.350 503.250 ;
        RECT 175.950 484.050 178.050 486.150 ;
        RECT 187.950 485.850 190.050 487.950 ;
        RECT 194.100 486.150 195.900 487.950 ;
        RECT 199.950 486.150 201.150 491.400 ;
        RECT 202.950 489.150 204.750 490.950 ;
        RECT 212.550 489.150 213.750 497.400 ;
        RECT 225.150 492.900 226.950 503.250 ;
        RECT 224.550 491.550 226.950 492.900 ;
        RECT 228.150 491.550 229.950 503.250 ;
        RECT 202.950 487.050 205.050 489.150 ;
        RECT 188.400 481.650 189.600 485.850 ;
        RECT 193.950 484.050 196.050 486.150 ;
        RECT 196.950 482.850 199.050 484.950 ;
        RECT 199.950 484.050 202.050 486.150 ;
        RECT 208.950 485.850 211.050 487.950 ;
        RECT 211.950 487.050 214.050 489.150 ;
        RECT 209.100 484.050 210.900 485.850 ;
        RECT 169.950 479.100 177.450 480.300 ;
        RECT 169.950 478.500 171.750 479.100 ;
        RECT 166.650 476.100 169.950 477.600 ;
        RECT 168.150 471.750 169.950 476.100 ;
        RECT 171.150 471.750 172.950 477.600 ;
        RECT 175.650 471.750 177.450 479.100 ;
        RECT 179.700 471.750 181.500 480.600 ;
        RECT 185.100 480.000 189.600 481.650 ;
        RECT 197.100 481.050 198.900 482.850 ;
        RECT 200.850 480.750 202.050 484.050 ;
        RECT 185.100 471.750 186.900 480.000 ;
        RECT 201.000 479.700 204.750 480.750 ;
        RECT 194.550 476.700 202.350 478.050 ;
        RECT 194.550 471.750 196.350 476.700 ;
        RECT 197.550 471.750 199.350 475.800 ;
        RECT 200.550 471.750 202.350 476.700 ;
        RECT 203.550 477.600 204.750 479.700 ;
        RECT 212.550 479.700 213.750 487.050 ;
        RECT 214.950 485.850 217.050 487.950 ;
        RECT 215.100 484.050 216.900 485.850 ;
        RECT 224.550 484.950 225.900 491.550 ;
        RECT 232.650 491.400 234.450 503.250 ;
        RECT 238.650 497.400 240.450 503.250 ;
        RECT 241.650 497.400 243.450 503.250 ;
        RECT 244.650 497.400 246.450 503.250 ;
        RECT 238.950 492.450 241.050 493.050 ;
        RECT 227.250 490.200 229.050 490.650 ;
        RECT 233.250 490.200 234.450 491.400 ;
        RECT 227.250 489.000 234.450 490.200 ;
        RECT 236.550 491.550 241.050 492.450 ;
        RECT 227.250 488.850 229.050 489.000 ;
        RECT 223.950 482.850 226.050 484.950 ;
        RECT 212.550 478.800 216.150 479.700 ;
        RECT 203.550 471.750 205.350 477.600 ;
        RECT 209.850 471.750 211.650 477.600 ;
        RECT 214.350 471.750 216.150 478.800 ;
        RECT 223.950 477.600 225.000 482.850 ;
        RECT 227.400 480.600 228.300 488.850 ;
        RECT 230.100 486.150 231.900 487.950 ;
        RECT 229.950 484.050 232.050 486.150 ;
        RECT 233.100 483.150 234.900 484.950 ;
        RECT 232.950 481.050 235.050 483.150 ;
        RECT 227.250 479.700 229.050 480.600 ;
        RECT 227.250 478.800 230.550 479.700 ;
        RECT 223.650 471.750 225.450 477.600 ;
        RECT 229.650 474.600 230.550 478.800 ;
        RECT 232.950 477.450 235.050 478.050 ;
        RECT 236.550 477.450 237.450 491.550 ;
        RECT 238.950 490.950 241.050 491.550 ;
        RECT 242.250 489.150 243.450 497.400 ;
        RECT 249.300 491.400 251.100 503.250 ;
        RECT 253.500 491.400 255.300 503.250 ;
        RECT 256.800 497.400 258.600 503.250 ;
        RECT 266.400 497.400 268.200 503.250 ;
        RECT 269.700 491.400 271.500 503.250 ;
        RECT 273.900 491.400 275.700 503.250 ;
        RECT 278.550 497.400 280.350 503.250 ;
        RECT 281.550 497.400 283.350 503.250 ;
        RECT 284.550 497.400 286.350 503.250 ;
        RECT 238.950 485.850 241.050 487.950 ;
        RECT 241.950 487.050 244.050 489.150 ;
        RECT 239.100 484.050 240.900 485.850 ;
        RECT 242.250 479.700 243.450 487.050 ;
        RECT 244.950 485.850 247.050 487.950 ;
        RECT 248.100 486.150 249.900 487.950 ;
        RECT 253.950 486.150 255.150 491.400 ;
        RECT 256.950 489.150 258.750 490.950 ;
        RECT 266.250 489.150 268.050 490.950 ;
        RECT 256.950 487.050 259.050 489.150 ;
        RECT 265.950 487.050 268.050 489.150 ;
        RECT 269.850 486.150 271.050 491.400 ;
        RECT 281.550 489.150 282.750 497.400 ;
        RECT 283.950 492.450 286.050 493.050 ;
        RECT 283.950 491.550 288.450 492.450 ;
        RECT 283.950 490.950 286.050 491.550 ;
        RECT 275.100 486.150 276.900 487.950 ;
        RECT 245.100 484.050 246.900 485.850 ;
        RECT 247.950 484.050 250.050 486.150 ;
        RECT 250.950 482.850 253.050 484.950 ;
        RECT 253.950 484.050 256.050 486.150 ;
        RECT 251.100 481.050 252.900 482.850 ;
        RECT 254.850 480.750 256.050 484.050 ;
        RECT 268.950 484.050 271.050 486.150 ;
        RECT 268.950 480.750 270.150 484.050 ;
        RECT 271.950 482.850 274.050 484.950 ;
        RECT 274.950 484.050 277.050 486.150 ;
        RECT 277.950 485.850 280.050 487.950 ;
        RECT 280.950 487.050 283.050 489.150 ;
        RECT 278.100 484.050 279.900 485.850 ;
        RECT 272.100 481.050 273.900 482.850 ;
        RECT 255.000 479.700 258.750 480.750 ;
        RECT 232.950 476.550 237.450 477.450 ;
        RECT 239.850 478.800 243.450 479.700 ;
        RECT 232.950 475.950 235.050 476.550 ;
        RECT 226.650 471.750 228.450 474.600 ;
        RECT 229.650 471.750 231.450 474.600 ;
        RECT 232.650 471.750 234.450 474.600 ;
        RECT 239.850 471.750 241.650 478.800 ;
        RECT 244.350 471.750 246.150 477.600 ;
        RECT 248.550 476.700 256.350 478.050 ;
        RECT 248.550 471.750 250.350 476.700 ;
        RECT 251.550 471.750 253.350 475.800 ;
        RECT 254.550 471.750 256.350 476.700 ;
        RECT 257.550 477.600 258.750 479.700 ;
        RECT 266.250 479.700 270.000 480.750 ;
        RECT 281.550 479.700 282.750 487.050 ;
        RECT 283.950 485.850 286.050 487.950 ;
        RECT 284.100 484.050 285.900 485.850 ;
        RECT 287.550 480.450 288.450 491.550 ;
        RECT 291.300 491.400 293.100 503.250 ;
        RECT 295.500 491.400 297.300 503.250 ;
        RECT 298.800 497.400 300.600 503.250 ;
        RECT 308.400 497.400 310.200 503.250 ;
        RECT 311.700 491.400 313.500 503.250 ;
        RECT 315.900 491.400 317.700 503.250 ;
        RECT 320.550 497.400 322.350 503.250 ;
        RECT 323.550 497.400 325.350 503.250 ;
        RECT 290.100 486.150 291.900 487.950 ;
        RECT 295.950 486.150 297.150 491.400 ;
        RECT 298.950 489.150 300.750 490.950 ;
        RECT 308.250 489.150 310.050 490.950 ;
        RECT 298.950 487.050 301.050 489.150 ;
        RECT 307.950 487.050 310.050 489.150 ;
        RECT 311.850 486.150 313.050 491.400 ;
        RECT 317.100 486.150 318.900 487.950 ;
        RECT 289.950 484.050 292.050 486.150 ;
        RECT 292.950 482.850 295.050 484.950 ;
        RECT 295.950 484.050 298.050 486.150 ;
        RECT 293.100 481.050 294.900 482.850 ;
        RECT 289.950 480.450 292.050 481.050 ;
        RECT 296.850 480.750 298.050 484.050 ;
        RECT 310.950 484.050 313.050 486.150 ;
        RECT 310.950 480.750 312.150 484.050 ;
        RECT 313.950 482.850 316.050 484.950 ;
        RECT 316.950 484.050 319.050 486.150 ;
        RECT 323.400 484.950 324.600 497.400 ;
        RECT 330.300 491.400 332.100 503.250 ;
        RECT 334.500 491.400 336.300 503.250 ;
        RECT 337.800 497.400 339.600 503.250 ;
        RECT 346.650 497.400 348.450 503.250 ;
        RECT 349.650 497.400 351.450 503.250 ;
        RECT 353.550 497.400 355.350 503.250 ;
        RECT 356.550 497.400 358.350 503.250 ;
        RECT 359.550 497.400 361.350 503.250 ;
        RECT 329.100 486.150 330.900 487.950 ;
        RECT 334.950 486.150 336.150 491.400 ;
        RECT 337.950 489.150 339.750 490.950 ;
        RECT 337.950 487.050 340.050 489.150 ;
        RECT 320.100 483.150 321.900 484.950 ;
        RECT 314.100 481.050 315.900 482.850 ;
        RECT 319.950 481.050 322.050 483.150 ;
        RECT 322.950 482.850 325.050 484.950 ;
        RECT 328.950 484.050 331.050 486.150 ;
        RECT 331.950 482.850 334.050 484.950 ;
        RECT 334.950 484.050 337.050 486.150 ;
        RECT 347.400 484.950 348.600 497.400 ;
        RECT 356.550 489.150 357.750 497.400 ;
        RECT 365.550 491.400 367.350 503.250 ;
        RECT 368.550 500.400 370.350 503.250 ;
        RECT 373.050 497.400 374.850 503.250 ;
        RECT 377.250 497.400 379.050 503.250 ;
        RECT 370.950 495.300 374.850 497.400 ;
        RECT 381.150 496.500 382.950 503.250 ;
        RECT 384.150 497.400 385.950 503.250 ;
        RECT 388.950 497.400 390.750 503.250 ;
        RECT 394.050 497.400 395.850 503.250 ;
        RECT 389.250 496.500 390.450 497.400 ;
        RECT 379.950 494.700 386.850 496.500 ;
        RECT 389.250 494.400 394.050 496.500 ;
        RECT 372.150 492.600 374.850 494.400 ;
        RECT 375.750 493.800 377.550 494.400 ;
        RECT 375.750 492.900 382.050 493.800 ;
        RECT 389.250 493.500 390.450 494.400 ;
        RECT 375.750 492.600 377.550 492.900 ;
        RECT 373.950 491.700 374.850 492.600 ;
        RECT 352.950 485.850 355.050 487.950 ;
        RECT 355.950 487.050 358.050 489.150 ;
        RECT 266.250 477.600 267.450 479.700 ;
        RECT 281.550 478.800 285.150 479.700 ;
        RECT 287.550 479.550 292.050 480.450 ;
        RECT 297.000 479.700 300.750 480.750 ;
        RECT 289.950 478.950 292.050 479.550 ;
        RECT 257.550 471.750 259.350 477.600 ;
        RECT 265.650 471.750 267.450 477.600 ;
        RECT 268.650 476.700 276.450 478.050 ;
        RECT 268.650 471.750 270.450 476.700 ;
        RECT 271.650 471.750 273.450 475.800 ;
        RECT 274.650 471.750 276.450 476.700 ;
        RECT 278.850 471.750 280.650 477.600 ;
        RECT 283.350 471.750 285.150 478.800 ;
        RECT 290.550 476.700 298.350 478.050 ;
        RECT 290.550 471.750 292.350 476.700 ;
        RECT 293.550 471.750 295.350 475.800 ;
        RECT 296.550 471.750 298.350 476.700 ;
        RECT 299.550 477.600 300.750 479.700 ;
        RECT 308.250 479.700 312.000 480.750 ;
        RECT 308.250 477.600 309.450 479.700 ;
        RECT 299.550 471.750 301.350 477.600 ;
        RECT 307.650 471.750 309.450 477.600 ;
        RECT 310.650 476.700 318.450 478.050 ;
        RECT 310.650 471.750 312.450 476.700 ;
        RECT 313.650 471.750 315.450 475.800 ;
        RECT 316.650 471.750 318.450 476.700 ;
        RECT 323.400 474.600 324.600 482.850 ;
        RECT 332.100 481.050 333.900 482.850 ;
        RECT 335.850 480.750 337.050 484.050 ;
        RECT 346.950 482.850 349.050 484.950 ;
        RECT 350.100 483.150 351.900 484.950 ;
        RECT 353.100 484.050 354.900 485.850 ;
        RECT 336.000 479.700 339.750 480.750 ;
        RECT 329.550 476.700 337.350 478.050 ;
        RECT 320.550 471.750 322.350 474.600 ;
        RECT 323.550 471.750 325.350 474.600 ;
        RECT 329.550 471.750 331.350 476.700 ;
        RECT 332.550 471.750 334.350 475.800 ;
        RECT 335.550 471.750 337.350 476.700 ;
        RECT 338.550 477.600 339.750 479.700 ;
        RECT 338.550 471.750 340.350 477.600 ;
        RECT 347.400 474.600 348.600 482.850 ;
        RECT 349.950 481.050 352.050 483.150 ;
        RECT 356.550 479.700 357.750 487.050 ;
        RECT 358.950 485.850 361.050 487.950 ;
        RECT 359.100 484.050 360.900 485.850 ;
        RECT 365.550 481.950 366.750 491.400 ;
        RECT 370.950 490.800 373.050 491.700 ;
        RECT 373.950 490.800 379.950 491.700 ;
        RECT 368.850 489.600 373.050 490.800 ;
        RECT 367.950 487.800 369.750 489.600 ;
        RECT 379.050 486.150 379.950 490.800 ;
        RECT 381.150 490.800 382.050 492.900 ;
        RECT 382.950 492.300 390.450 493.500 ;
        RECT 382.950 491.700 384.750 492.300 ;
        RECT 397.050 491.400 398.850 503.250 ;
        RECT 387.750 490.800 398.850 491.400 ;
        RECT 381.150 490.200 398.850 490.800 ;
        RECT 381.150 489.900 389.550 490.200 ;
        RECT 387.750 489.600 389.550 489.900 ;
        RECT 379.050 484.050 382.050 486.150 ;
        RECT 385.950 485.100 388.050 486.150 ;
        RECT 385.950 484.050 393.900 485.100 ;
        RECT 367.950 483.750 370.050 484.050 ;
        RECT 367.950 481.950 371.850 483.750 ;
        RECT 365.550 479.850 370.050 481.950 ;
        RECT 379.050 480.000 379.950 484.050 ;
        RECT 392.100 483.300 393.900 484.050 ;
        RECT 395.100 483.150 396.900 484.950 ;
        RECT 389.100 482.400 390.900 483.000 ;
        RECT 395.100 482.400 396.000 483.150 ;
        RECT 389.100 481.200 396.000 482.400 ;
        RECT 389.100 480.000 390.150 481.200 ;
        RECT 356.550 478.800 360.150 479.700 ;
        RECT 346.650 471.750 348.450 474.600 ;
        RECT 349.650 471.750 351.450 474.600 ;
        RECT 353.850 471.750 355.650 477.600 ;
        RECT 358.350 471.750 360.150 478.800 ;
        RECT 365.550 477.600 366.750 479.850 ;
        RECT 379.050 479.100 390.150 480.000 ;
        RECT 379.050 478.800 379.950 479.100 ;
        RECT 365.550 471.750 367.350 477.600 ;
        RECT 370.950 476.700 373.050 477.600 ;
        RECT 378.150 477.000 379.950 478.800 ;
        RECT 389.100 478.200 390.150 479.100 ;
        RECT 385.350 477.450 387.150 478.200 ;
        RECT 370.950 475.500 374.700 476.700 ;
        RECT 373.650 474.600 374.700 475.500 ;
        RECT 382.200 476.400 387.150 477.450 ;
        RECT 388.650 476.400 390.450 478.200 ;
        RECT 397.950 477.600 398.850 490.200 ;
        RECT 401.550 497.400 403.350 503.250 ;
        RECT 401.550 490.500 402.750 497.400 ;
        RECT 404.850 491.400 406.650 503.250 ;
        RECT 407.850 491.400 409.650 503.250 ;
        RECT 413.550 491.400 415.350 503.250 ;
        RECT 416.550 500.400 418.350 503.250 ;
        RECT 421.050 497.400 422.850 503.250 ;
        RECT 425.250 497.400 427.050 503.250 ;
        RECT 418.950 495.300 422.850 497.400 ;
        RECT 429.150 496.500 430.950 503.250 ;
        RECT 432.150 497.400 433.950 503.250 ;
        RECT 436.950 497.400 438.750 503.250 ;
        RECT 442.050 497.400 443.850 503.250 ;
        RECT 437.250 496.500 438.450 497.400 ;
        RECT 427.950 494.700 434.850 496.500 ;
        RECT 437.250 494.400 442.050 496.500 ;
        RECT 420.150 492.600 422.850 494.400 ;
        RECT 423.750 493.800 425.550 494.400 ;
        RECT 423.750 492.900 430.050 493.800 ;
        RECT 437.250 493.500 438.450 494.400 ;
        RECT 423.750 492.600 425.550 492.900 ;
        RECT 421.950 491.700 422.850 492.600 ;
        RECT 401.550 489.600 407.250 490.500 ;
        RECT 405.000 488.700 407.250 489.600 ;
        RECT 401.100 486.150 402.900 487.950 ;
        RECT 400.950 484.050 403.050 486.150 ;
        RECT 405.000 480.300 406.050 488.700 ;
        RECT 408.150 486.150 409.350 491.400 ;
        RECT 406.950 484.050 409.350 486.150 ;
        RECT 405.000 479.400 407.250 480.300 ;
        RECT 382.200 474.600 383.250 476.400 ;
        RECT 391.950 475.500 394.050 477.600 ;
        RECT 391.950 474.600 393.000 475.500 ;
        RECT 368.850 471.750 370.650 474.600 ;
        RECT 373.350 471.750 375.150 474.600 ;
        RECT 377.550 471.750 379.350 474.600 ;
        RECT 381.450 471.750 383.250 474.600 ;
        RECT 384.750 471.750 386.550 474.600 ;
        RECT 389.250 473.700 393.000 474.600 ;
        RECT 389.250 471.750 391.050 473.700 ;
        RECT 394.050 471.750 395.850 474.600 ;
        RECT 397.050 471.750 398.850 477.600 ;
        RECT 402.150 478.500 407.250 479.400 ;
        RECT 402.150 474.600 403.350 478.500 ;
        RECT 408.150 477.600 409.350 484.050 ;
        RECT 413.550 481.950 414.750 491.400 ;
        RECT 418.950 490.800 421.050 491.700 ;
        RECT 421.950 490.800 427.950 491.700 ;
        RECT 416.850 489.600 421.050 490.800 ;
        RECT 415.950 487.800 417.750 489.600 ;
        RECT 427.050 486.150 427.950 490.800 ;
        RECT 429.150 490.800 430.050 492.900 ;
        RECT 430.950 492.300 438.450 493.500 ;
        RECT 430.950 491.700 432.750 492.300 ;
        RECT 445.050 491.400 446.850 503.250 ;
        RECT 452.400 497.400 454.200 503.250 ;
        RECT 455.700 491.400 457.500 503.250 ;
        RECT 459.900 491.400 461.700 503.250 ;
        RECT 467.400 497.400 469.200 503.250 ;
        RECT 470.700 491.400 472.500 503.250 ;
        RECT 474.900 491.400 476.700 503.250 ;
        RECT 480.300 491.400 482.100 503.250 ;
        RECT 484.500 491.400 486.300 503.250 ;
        RECT 487.800 497.400 489.600 503.250 ;
        RECT 497.400 497.400 499.200 503.250 ;
        RECT 500.700 491.400 502.500 503.250 ;
        RECT 504.900 491.400 506.700 503.250 ;
        RECT 510.300 491.400 512.100 503.250 ;
        RECT 514.500 491.400 516.300 503.250 ;
        RECT 517.800 497.400 519.600 503.250 ;
        RECT 524.550 497.400 526.350 503.250 ;
        RECT 527.550 497.400 529.350 503.250 ;
        RECT 530.550 497.400 532.350 503.250 ;
        RECT 536.550 497.400 538.350 503.250 ;
        RECT 539.550 497.400 541.350 503.250 ;
        RECT 542.550 497.400 544.350 503.250 ;
        RECT 548.550 497.400 550.350 503.250 ;
        RECT 551.550 497.400 553.350 503.250 ;
        RECT 554.550 497.400 556.350 503.250 ;
        RECT 560.550 497.400 562.350 503.250 ;
        RECT 563.550 497.400 565.350 503.250 ;
        RECT 566.550 497.400 568.350 503.250 ;
        RECT 572.550 497.400 574.350 503.250 ;
        RECT 435.750 490.800 446.850 491.400 ;
        RECT 429.150 490.200 446.850 490.800 ;
        RECT 429.150 489.900 437.550 490.200 ;
        RECT 435.750 489.600 437.550 489.900 ;
        RECT 427.050 484.050 430.050 486.150 ;
        RECT 433.950 485.100 436.050 486.150 ;
        RECT 433.950 484.050 441.900 485.100 ;
        RECT 415.950 483.750 418.050 484.050 ;
        RECT 415.950 481.950 419.850 483.750 ;
        RECT 413.550 479.850 418.050 481.950 ;
        RECT 427.050 480.000 427.950 484.050 ;
        RECT 440.100 483.300 441.900 484.050 ;
        RECT 443.100 483.150 444.900 484.950 ;
        RECT 437.100 482.400 438.900 483.000 ;
        RECT 443.100 482.400 444.000 483.150 ;
        RECT 437.100 481.200 444.000 482.400 ;
        RECT 437.100 480.000 438.150 481.200 ;
        RECT 413.550 477.600 414.750 479.850 ;
        RECT 427.050 479.100 438.150 480.000 ;
        RECT 427.050 478.800 427.950 479.100 ;
        RECT 401.550 471.750 403.350 474.600 ;
        RECT 404.850 471.750 406.650 477.600 ;
        RECT 407.850 471.750 409.650 477.600 ;
        RECT 413.550 471.750 415.350 477.600 ;
        RECT 418.950 476.700 421.050 477.600 ;
        RECT 426.150 477.000 427.950 478.800 ;
        RECT 437.100 478.200 438.150 479.100 ;
        RECT 433.350 477.450 435.150 478.200 ;
        RECT 418.950 475.500 422.700 476.700 ;
        RECT 421.650 474.600 422.700 475.500 ;
        RECT 430.200 476.400 435.150 477.450 ;
        RECT 436.650 476.400 438.450 478.200 ;
        RECT 445.950 477.600 446.850 490.200 ;
        RECT 452.250 489.150 454.050 490.950 ;
        RECT 451.950 487.050 454.050 489.150 ;
        RECT 455.850 486.150 457.050 491.400 ;
        RECT 467.250 489.150 469.050 490.950 ;
        RECT 461.100 486.150 462.900 487.950 ;
        RECT 466.950 487.050 469.050 489.150 ;
        RECT 470.850 486.150 472.050 491.400 ;
        RECT 476.100 486.150 477.900 487.950 ;
        RECT 479.100 486.150 480.900 487.950 ;
        RECT 484.950 486.150 486.150 491.400 ;
        RECT 487.950 489.150 489.750 490.950 ;
        RECT 497.250 489.150 499.050 490.950 ;
        RECT 487.950 487.050 490.050 489.150 ;
        RECT 496.950 487.050 499.050 489.150 ;
        RECT 500.850 486.150 502.050 491.400 ;
        RECT 506.100 486.150 507.900 487.950 ;
        RECT 509.100 486.150 510.900 487.950 ;
        RECT 514.950 486.150 516.150 491.400 ;
        RECT 517.950 489.150 519.750 490.950 ;
        RECT 527.550 489.150 528.750 497.400 ;
        RECT 539.550 489.150 540.750 497.400 ;
        RECT 551.550 489.150 552.750 497.400 ;
        RECT 563.550 489.150 564.750 497.400 ;
        RECT 572.550 490.500 573.750 497.400 ;
        RECT 575.850 491.400 577.650 503.250 ;
        RECT 578.850 491.400 580.650 503.250 ;
        RECT 586.650 497.400 588.450 503.250 ;
        RECT 589.650 497.400 591.450 503.250 ;
        RECT 592.650 497.400 594.450 503.250 ;
        RECT 572.550 489.600 578.250 490.500 ;
        RECT 517.950 487.050 520.050 489.150 ;
        RECT 454.950 484.050 457.050 486.150 ;
        RECT 454.950 480.750 456.150 484.050 ;
        RECT 457.950 482.850 460.050 484.950 ;
        RECT 460.950 484.050 463.050 486.150 ;
        RECT 469.950 484.050 472.050 486.150 ;
        RECT 458.100 481.050 459.900 482.850 ;
        RECT 469.950 480.750 471.150 484.050 ;
        RECT 472.950 482.850 475.050 484.950 ;
        RECT 475.950 484.050 478.050 486.150 ;
        RECT 478.950 484.050 481.050 486.150 ;
        RECT 481.950 482.850 484.050 484.950 ;
        RECT 484.950 484.050 487.050 486.150 ;
        RECT 473.100 481.050 474.900 482.850 ;
        RECT 482.100 481.050 483.900 482.850 ;
        RECT 485.850 480.750 487.050 484.050 ;
        RECT 499.950 484.050 502.050 486.150 ;
        RECT 499.950 480.750 501.150 484.050 ;
        RECT 502.950 482.850 505.050 484.950 ;
        RECT 505.950 484.050 508.050 486.150 ;
        RECT 508.950 484.050 511.050 486.150 ;
        RECT 511.950 482.850 514.050 484.950 ;
        RECT 514.950 484.050 517.050 486.150 ;
        RECT 523.950 485.850 526.050 487.950 ;
        RECT 526.950 487.050 529.050 489.150 ;
        RECT 524.100 484.050 525.900 485.850 ;
        RECT 503.100 481.050 504.900 482.850 ;
        RECT 512.100 481.050 513.900 482.850 ;
        RECT 515.850 480.750 517.050 484.050 ;
        RECT 452.250 479.700 456.000 480.750 ;
        RECT 467.250 479.700 471.000 480.750 ;
        RECT 486.000 479.700 489.750 480.750 ;
        RECT 452.250 477.600 453.450 479.700 ;
        RECT 430.200 474.600 431.250 476.400 ;
        RECT 439.950 475.500 442.050 477.600 ;
        RECT 439.950 474.600 441.000 475.500 ;
        RECT 416.850 471.750 418.650 474.600 ;
        RECT 421.350 471.750 423.150 474.600 ;
        RECT 425.550 471.750 427.350 474.600 ;
        RECT 429.450 471.750 431.250 474.600 ;
        RECT 432.750 471.750 434.550 474.600 ;
        RECT 437.250 473.700 441.000 474.600 ;
        RECT 437.250 471.750 439.050 473.700 ;
        RECT 442.050 471.750 443.850 474.600 ;
        RECT 445.050 471.750 446.850 477.600 ;
        RECT 451.650 471.750 453.450 477.600 ;
        RECT 454.650 476.700 462.450 478.050 ;
        RECT 467.250 477.600 468.450 479.700 ;
        RECT 454.650 471.750 456.450 476.700 ;
        RECT 457.650 471.750 459.450 475.800 ;
        RECT 460.650 471.750 462.450 476.700 ;
        RECT 466.650 471.750 468.450 477.600 ;
        RECT 469.650 476.700 477.450 478.050 ;
        RECT 469.650 471.750 471.450 476.700 ;
        RECT 472.650 471.750 474.450 475.800 ;
        RECT 475.650 471.750 477.450 476.700 ;
        RECT 479.550 476.700 487.350 478.050 ;
        RECT 479.550 471.750 481.350 476.700 ;
        RECT 482.550 471.750 484.350 475.800 ;
        RECT 485.550 471.750 487.350 476.700 ;
        RECT 488.550 477.600 489.750 479.700 ;
        RECT 497.250 479.700 501.000 480.750 ;
        RECT 516.000 479.700 519.750 480.750 ;
        RECT 497.250 477.600 498.450 479.700 ;
        RECT 488.550 471.750 490.350 477.600 ;
        RECT 496.650 471.750 498.450 477.600 ;
        RECT 499.650 476.700 507.450 478.050 ;
        RECT 499.650 471.750 501.450 476.700 ;
        RECT 502.650 471.750 504.450 475.800 ;
        RECT 505.650 471.750 507.450 476.700 ;
        RECT 509.550 476.700 517.350 478.050 ;
        RECT 509.550 471.750 511.350 476.700 ;
        RECT 512.550 471.750 514.350 475.800 ;
        RECT 515.550 471.750 517.350 476.700 ;
        RECT 518.550 477.600 519.750 479.700 ;
        RECT 527.550 479.700 528.750 487.050 ;
        RECT 529.950 485.850 532.050 487.950 ;
        RECT 535.950 485.850 538.050 487.950 ;
        RECT 538.950 487.050 541.050 489.150 ;
        RECT 530.100 484.050 531.900 485.850 ;
        RECT 536.100 484.050 537.900 485.850 ;
        RECT 539.550 479.700 540.750 487.050 ;
        RECT 541.950 485.850 544.050 487.950 ;
        RECT 547.950 485.850 550.050 487.950 ;
        RECT 550.950 487.050 553.050 489.150 ;
        RECT 542.100 484.050 543.900 485.850 ;
        RECT 548.100 484.050 549.900 485.850 ;
        RECT 551.550 479.700 552.750 487.050 ;
        RECT 553.950 485.850 556.050 487.950 ;
        RECT 559.950 485.850 562.050 487.950 ;
        RECT 562.950 487.050 565.050 489.150 ;
        RECT 576.000 488.700 578.250 489.600 ;
        RECT 554.100 484.050 555.900 485.850 ;
        RECT 560.100 484.050 561.900 485.850 ;
        RECT 563.550 479.700 564.750 487.050 ;
        RECT 565.950 485.850 568.050 487.950 ;
        RECT 572.100 486.150 573.900 487.950 ;
        RECT 566.100 484.050 567.900 485.850 ;
        RECT 571.950 484.050 574.050 486.150 ;
        RECT 576.000 480.300 577.050 488.700 ;
        RECT 579.150 486.150 580.350 491.400 ;
        RECT 590.250 489.150 591.450 497.400 ;
        RECT 600.450 491.400 602.250 503.250 ;
        RECT 604.650 491.400 606.450 503.250 ;
        RECT 608.550 497.400 610.350 503.250 ;
        RECT 600.450 490.350 603.000 491.400 ;
        RECT 577.950 484.050 580.350 486.150 ;
        RECT 586.950 485.850 589.050 487.950 ;
        RECT 589.950 487.050 592.050 489.150 ;
        RECT 587.100 484.050 588.900 485.850 ;
        RECT 527.550 478.800 531.150 479.700 ;
        RECT 539.550 478.800 543.150 479.700 ;
        RECT 551.550 478.800 555.150 479.700 ;
        RECT 563.550 478.800 567.150 479.700 ;
        RECT 576.000 479.400 578.250 480.300 ;
        RECT 518.550 471.750 520.350 477.600 ;
        RECT 524.850 471.750 526.650 477.600 ;
        RECT 529.350 471.750 531.150 478.800 ;
        RECT 536.850 471.750 538.650 477.600 ;
        RECT 541.350 471.750 543.150 478.800 ;
        RECT 548.850 471.750 550.650 477.600 ;
        RECT 553.350 471.750 555.150 478.800 ;
        RECT 560.850 471.750 562.650 477.600 ;
        RECT 565.350 471.750 567.150 478.800 ;
        RECT 573.150 478.500 578.250 479.400 ;
        RECT 573.150 474.600 574.350 478.500 ;
        RECT 579.150 477.600 580.350 484.050 ;
        RECT 590.250 479.700 591.450 487.050 ;
        RECT 592.950 485.850 595.050 487.950 ;
        RECT 599.100 486.150 600.900 487.950 ;
        RECT 593.100 484.050 594.900 485.850 ;
        RECT 598.950 484.050 601.050 486.150 ;
        RECT 587.850 478.800 591.450 479.700 ;
        RECT 601.950 483.150 603.000 490.350 ;
        RECT 608.550 490.500 609.750 497.400 ;
        RECT 611.850 491.400 613.650 503.250 ;
        RECT 614.850 491.400 616.650 503.250 ;
        RECT 622.650 497.400 624.450 503.250 ;
        RECT 625.650 497.400 627.450 503.250 ;
        RECT 632.400 497.400 634.200 503.250 ;
        RECT 608.550 489.600 614.250 490.500 ;
        RECT 612.000 488.700 614.250 489.600 ;
        RECT 605.100 486.150 606.900 487.950 ;
        RECT 608.100 486.150 609.900 487.950 ;
        RECT 604.950 484.050 607.050 486.150 ;
        RECT 607.950 484.050 610.050 486.150 ;
        RECT 601.950 481.050 604.050 483.150 ;
        RECT 572.550 471.750 574.350 474.600 ;
        RECT 575.850 471.750 577.650 477.600 ;
        RECT 578.850 471.750 580.650 477.600 ;
        RECT 587.850 471.750 589.650 478.800 ;
        RECT 592.350 471.750 594.150 477.600 ;
        RECT 601.950 474.600 603.000 481.050 ;
        RECT 612.000 480.300 613.050 488.700 ;
        RECT 615.150 486.150 616.350 491.400 ;
        RECT 613.950 484.050 616.350 486.150 ;
        RECT 623.400 484.950 624.600 497.400 ;
        RECT 635.700 491.400 637.500 503.250 ;
        RECT 639.900 491.400 641.700 503.250 ;
        RECT 646.650 497.400 648.450 503.250 ;
        RECT 649.650 497.400 651.450 503.250 ;
        RECT 632.250 489.150 634.050 490.950 ;
        RECT 631.950 487.050 634.050 489.150 ;
        RECT 635.850 486.150 637.050 491.400 ;
        RECT 641.100 486.150 642.900 487.950 ;
        RECT 612.000 479.400 614.250 480.300 ;
        RECT 609.150 478.500 614.250 479.400 ;
        RECT 609.150 474.600 610.350 478.500 ;
        RECT 615.150 477.600 616.350 484.050 ;
        RECT 622.950 482.850 625.050 484.950 ;
        RECT 626.100 483.150 627.900 484.950 ;
        RECT 634.950 484.050 637.050 486.150 ;
        RECT 598.650 471.750 600.450 474.600 ;
        RECT 601.650 471.750 603.450 474.600 ;
        RECT 604.650 471.750 606.450 474.600 ;
        RECT 608.550 471.750 610.350 474.600 ;
        RECT 611.850 471.750 613.650 477.600 ;
        RECT 614.850 471.750 616.650 477.600 ;
        RECT 623.400 474.600 624.600 482.850 ;
        RECT 625.950 481.050 628.050 483.150 ;
        RECT 634.950 480.750 636.150 484.050 ;
        RECT 637.950 482.850 640.050 484.950 ;
        RECT 640.950 484.050 643.050 486.150 ;
        RECT 647.400 484.950 648.600 497.400 ;
        RECT 654.300 491.400 656.100 503.250 ;
        RECT 658.500 491.400 660.300 503.250 ;
        RECT 661.800 497.400 663.600 503.250 ;
        RECT 670.650 497.400 672.450 503.250 ;
        RECT 673.650 497.400 675.450 503.250 ;
        RECT 676.650 497.400 678.450 503.250 ;
        RECT 653.100 486.150 654.900 487.950 ;
        RECT 658.950 486.150 660.150 491.400 ;
        RECT 661.950 489.150 663.750 490.950 ;
        RECT 674.250 489.150 675.450 497.400 ;
        RECT 681.150 491.400 682.950 503.250 ;
        RECT 684.150 497.400 685.950 503.250 ;
        RECT 689.250 497.400 691.050 503.250 ;
        RECT 694.050 497.400 695.850 503.250 ;
        RECT 689.550 496.500 690.750 497.400 ;
        RECT 697.050 496.500 698.850 503.250 ;
        RECT 700.950 497.400 702.750 503.250 ;
        RECT 705.150 497.400 706.950 503.250 ;
        RECT 709.650 500.400 711.450 503.250 ;
        RECT 685.950 494.400 690.750 496.500 ;
        RECT 693.150 494.700 700.050 496.500 ;
        RECT 705.150 495.300 709.050 497.400 ;
        RECT 689.550 493.500 690.750 494.400 ;
        RECT 702.450 493.800 704.250 494.400 ;
        RECT 689.550 492.300 697.050 493.500 ;
        RECT 695.250 491.700 697.050 492.300 ;
        RECT 697.950 492.900 704.250 493.800 ;
        RECT 681.150 490.800 692.250 491.400 ;
        RECT 697.950 490.800 698.850 492.900 ;
        RECT 702.450 492.600 704.250 492.900 ;
        RECT 705.150 492.600 707.850 494.400 ;
        RECT 705.150 491.700 706.050 492.600 ;
        RECT 681.150 490.200 698.850 490.800 ;
        RECT 661.950 487.050 664.050 489.150 ;
        RECT 646.950 482.850 649.050 484.950 ;
        RECT 650.100 483.150 651.900 484.950 ;
        RECT 652.950 484.050 655.050 486.150 ;
        RECT 638.100 481.050 639.900 482.850 ;
        RECT 632.250 479.700 636.000 480.750 ;
        RECT 632.250 477.600 633.450 479.700 ;
        RECT 622.650 471.750 624.450 474.600 ;
        RECT 625.650 471.750 627.450 474.600 ;
        RECT 631.650 471.750 633.450 477.600 ;
        RECT 634.650 476.700 642.450 478.050 ;
        RECT 634.650 471.750 636.450 476.700 ;
        RECT 637.650 471.750 639.450 475.800 ;
        RECT 640.650 471.750 642.450 476.700 ;
        RECT 647.400 474.600 648.600 482.850 ;
        RECT 649.950 481.050 652.050 483.150 ;
        RECT 655.950 482.850 658.050 484.950 ;
        RECT 658.950 484.050 661.050 486.150 ;
        RECT 670.950 485.850 673.050 487.950 ;
        RECT 673.950 487.050 676.050 489.150 ;
        RECT 671.100 484.050 672.900 485.850 ;
        RECT 656.100 481.050 657.900 482.850 ;
        RECT 659.850 480.750 661.050 484.050 ;
        RECT 660.000 479.700 663.750 480.750 ;
        RECT 674.250 479.700 675.450 487.050 ;
        RECT 676.950 485.850 679.050 487.950 ;
        RECT 677.100 484.050 678.900 485.850 ;
        RECT 653.550 476.700 661.350 478.050 ;
        RECT 646.650 471.750 648.450 474.600 ;
        RECT 649.650 471.750 651.450 474.600 ;
        RECT 653.550 471.750 655.350 476.700 ;
        RECT 656.550 471.750 658.350 475.800 ;
        RECT 659.550 471.750 661.350 476.700 ;
        RECT 662.550 477.600 663.750 479.700 ;
        RECT 671.850 478.800 675.450 479.700 ;
        RECT 662.550 471.750 664.350 477.600 ;
        RECT 671.850 471.750 673.650 478.800 ;
        RECT 681.150 477.600 682.050 490.200 ;
        RECT 690.450 489.900 698.850 490.200 ;
        RECT 700.050 490.800 706.050 491.700 ;
        RECT 706.950 490.800 709.050 491.700 ;
        RECT 712.650 491.400 714.450 503.250 ;
        RECT 690.450 489.600 692.250 489.900 ;
        RECT 700.050 486.150 700.950 490.800 ;
        RECT 706.950 489.600 711.150 490.800 ;
        RECT 710.250 487.800 712.050 489.600 ;
        RECT 691.950 485.100 694.050 486.150 ;
        RECT 683.100 483.150 684.900 484.950 ;
        RECT 686.100 484.050 694.050 485.100 ;
        RECT 697.950 484.050 700.950 486.150 ;
        RECT 686.100 483.300 687.900 484.050 ;
        RECT 684.000 482.400 684.900 483.150 ;
        RECT 689.100 482.400 690.900 483.000 ;
        RECT 684.000 481.200 690.900 482.400 ;
        RECT 689.850 480.000 690.900 481.200 ;
        RECT 700.050 480.000 700.950 484.050 ;
        RECT 709.950 483.750 712.050 484.050 ;
        RECT 708.150 481.950 712.050 483.750 ;
        RECT 713.250 481.950 714.450 491.400 ;
        RECT 689.850 479.100 700.950 480.000 ;
        RECT 709.950 479.850 714.450 481.950 ;
        RECT 689.850 478.200 690.900 479.100 ;
        RECT 700.050 478.800 700.950 479.100 ;
        RECT 676.350 471.750 678.150 477.600 ;
        RECT 681.150 471.750 682.950 477.600 ;
        RECT 685.950 475.500 688.050 477.600 ;
        RECT 689.550 476.400 691.350 478.200 ;
        RECT 692.850 477.450 694.650 478.200 ;
        RECT 692.850 476.400 697.800 477.450 ;
        RECT 700.050 477.000 701.850 478.800 ;
        RECT 713.250 477.600 714.450 479.850 ;
        RECT 706.950 476.700 709.050 477.600 ;
        RECT 687.000 474.600 688.050 475.500 ;
        RECT 696.750 474.600 697.800 476.400 ;
        RECT 705.300 475.500 709.050 476.700 ;
        RECT 705.300 474.600 706.350 475.500 ;
        RECT 684.150 471.750 685.950 474.600 ;
        RECT 687.000 473.700 690.750 474.600 ;
        RECT 688.950 471.750 690.750 473.700 ;
        RECT 693.450 471.750 695.250 474.600 ;
        RECT 696.750 471.750 698.550 474.600 ;
        RECT 700.650 471.750 702.450 474.600 ;
        RECT 704.850 471.750 706.650 474.600 ;
        RECT 709.350 471.750 711.150 474.600 ;
        RECT 712.650 471.750 714.450 477.600 ;
        RECT 7.800 461.400 9.600 467.250 ;
        RECT 12.000 461.400 13.800 467.250 ;
        RECT 16.200 461.400 18.000 467.250 ;
        RECT 24.150 462.900 25.950 467.250 ;
        RECT 22.650 461.400 25.950 462.900 ;
        RECT 27.150 461.400 28.950 467.250 ;
        RECT 8.250 456.150 10.050 457.950 ;
        RECT 4.950 452.850 7.050 454.950 ;
        RECT 7.950 454.050 10.050 456.150 ;
        RECT 12.000 454.950 13.050 461.400 ;
        RECT 10.950 452.850 13.050 454.950 ;
        RECT 13.950 456.150 15.750 457.950 ;
        RECT 13.950 454.050 16.050 456.150 ;
        RECT 22.650 454.950 23.850 461.400 ;
        RECT 25.950 459.900 27.750 460.500 ;
        RECT 31.650 459.900 33.450 467.250 ;
        RECT 25.950 458.700 33.450 459.900 ;
        RECT 35.550 461.400 37.350 467.250 ;
        RECT 38.850 464.400 40.650 467.250 ;
        RECT 43.350 464.400 45.150 467.250 ;
        RECT 47.550 464.400 49.350 467.250 ;
        RECT 51.450 464.400 53.250 467.250 ;
        RECT 54.750 464.400 56.550 467.250 ;
        RECT 59.250 465.300 61.050 467.250 ;
        RECT 59.250 464.400 63.000 465.300 ;
        RECT 64.050 464.400 65.850 467.250 ;
        RECT 43.650 463.500 44.700 464.400 ;
        RECT 40.950 462.300 44.700 463.500 ;
        RECT 52.200 462.600 53.250 464.400 ;
        RECT 61.950 463.500 63.000 464.400 ;
        RECT 40.950 461.400 43.050 462.300 ;
        RECT 35.550 459.150 36.750 461.400 ;
        RECT 48.150 460.200 49.950 462.000 ;
        RECT 52.200 461.550 57.150 462.600 ;
        RECT 55.350 460.800 57.150 461.550 ;
        RECT 58.650 460.800 60.450 462.600 ;
        RECT 61.950 461.400 64.050 463.500 ;
        RECT 67.050 461.400 68.850 467.250 ;
        RECT 49.050 459.900 49.950 460.200 ;
        RECT 59.100 459.900 60.150 460.800 ;
        RECT 16.950 452.850 19.050 454.950 ;
        RECT 22.650 452.850 25.050 454.950 ;
        RECT 26.100 453.150 27.900 454.950 ;
        RECT 5.100 451.050 6.900 452.850 ;
        RECT 10.950 449.400 11.850 452.850 ;
        RECT 16.950 451.050 18.750 452.850 ;
        RECT 7.800 448.500 11.850 449.400 ;
        RECT 7.800 447.600 9.600 448.500 ;
        RECT 22.650 447.600 23.850 452.850 ;
        RECT 25.950 451.050 28.050 453.150 ;
        RECT 4.650 436.500 6.450 447.600 ;
        RECT 7.650 437.400 9.450 447.600 ;
        RECT 10.650 446.400 18.450 447.300 ;
        RECT 10.650 436.500 12.450 446.400 ;
        RECT 4.650 435.750 12.450 436.500 ;
        RECT 13.650 435.750 15.450 445.500 ;
        RECT 16.650 435.750 18.450 446.400 ;
        RECT 22.050 435.750 23.850 447.600 ;
        RECT 25.050 435.750 26.850 447.600 ;
        RECT 29.100 441.600 30.300 458.700 ;
        RECT 35.550 457.050 40.050 459.150 ;
        RECT 49.050 459.000 60.150 459.900 ;
        RECT 31.950 452.850 34.050 454.950 ;
        RECT 32.100 451.050 33.900 452.850 ;
        RECT 35.550 447.600 36.750 457.050 ;
        RECT 37.950 455.250 41.850 457.050 ;
        RECT 37.950 454.950 40.050 455.250 ;
        RECT 49.050 454.950 49.950 459.000 ;
        RECT 59.100 457.800 60.150 459.000 ;
        RECT 59.100 456.600 66.000 457.800 ;
        RECT 59.100 456.000 60.900 456.600 ;
        RECT 65.100 455.850 66.000 456.600 ;
        RECT 62.100 454.950 63.900 455.700 ;
        RECT 49.050 452.850 52.050 454.950 ;
        RECT 55.950 453.900 63.900 454.950 ;
        RECT 65.100 454.050 66.900 455.850 ;
        RECT 55.950 452.850 58.050 453.900 ;
        RECT 37.950 449.400 39.750 451.200 ;
        RECT 38.850 448.200 43.050 449.400 ;
        RECT 49.050 448.200 49.950 452.850 ;
        RECT 57.750 449.100 59.550 449.400 ;
        RECT 28.650 435.750 30.450 441.600 ;
        RECT 31.650 435.750 33.450 441.600 ;
        RECT 35.550 435.750 37.350 447.600 ;
        RECT 40.950 447.300 43.050 448.200 ;
        RECT 43.950 447.300 49.950 448.200 ;
        RECT 51.150 448.800 59.550 449.100 ;
        RECT 67.950 448.800 68.850 461.400 ;
        RECT 71.550 462.300 73.350 467.250 ;
        RECT 74.550 463.200 76.350 467.250 ;
        RECT 77.550 462.300 79.350 467.250 ;
        RECT 71.550 460.950 79.350 462.300 ;
        RECT 80.550 461.400 82.350 467.250 ;
        RECT 86.850 461.400 88.650 467.250 ;
        RECT 80.550 459.300 81.750 461.400 ;
        RECT 91.350 460.200 93.150 467.250 ;
        RECT 85.950 459.450 88.050 460.050 ;
        RECT 78.000 458.250 81.750 459.300 ;
        RECT 83.550 458.550 88.050 459.450 ;
        RECT 74.100 456.150 75.900 457.950 ;
        RECT 70.950 452.850 73.050 454.950 ;
        RECT 73.950 454.050 76.050 456.150 ;
        RECT 77.850 454.950 79.050 458.250 ;
        RECT 76.950 452.850 79.050 454.950 ;
        RECT 71.100 451.050 72.900 452.850 ;
        RECT 51.150 448.200 68.850 448.800 ;
        RECT 43.950 446.400 44.850 447.300 ;
        RECT 42.150 444.600 44.850 446.400 ;
        RECT 45.750 446.100 47.550 446.400 ;
        RECT 51.150 446.100 52.050 448.200 ;
        RECT 57.750 447.600 68.850 448.200 ;
        RECT 76.950 447.600 78.150 452.850 ;
        RECT 79.950 449.850 82.050 451.950 ;
        RECT 79.950 448.050 81.750 449.850 ;
        RECT 45.750 445.200 52.050 446.100 ;
        RECT 52.950 446.700 54.750 447.300 ;
        RECT 52.950 445.500 60.450 446.700 ;
        RECT 45.750 444.600 47.550 445.200 ;
        RECT 59.250 444.600 60.450 445.500 ;
        RECT 40.950 441.600 44.850 443.700 ;
        RECT 49.950 442.500 56.850 444.300 ;
        RECT 59.250 442.500 64.050 444.600 ;
        RECT 38.550 435.750 40.350 438.600 ;
        RECT 43.050 435.750 44.850 441.600 ;
        RECT 47.250 435.750 49.050 441.600 ;
        RECT 51.150 435.750 52.950 442.500 ;
        RECT 59.250 441.600 60.450 442.500 ;
        RECT 54.150 435.750 55.950 441.600 ;
        RECT 58.950 435.750 60.750 441.600 ;
        RECT 64.050 435.750 65.850 441.600 ;
        RECT 67.050 435.750 68.850 447.600 ;
        RECT 72.300 435.750 74.100 447.600 ;
        RECT 76.500 435.750 78.300 447.600 ;
        RECT 79.950 444.450 82.050 445.050 ;
        RECT 83.550 444.450 84.450 458.550 ;
        RECT 85.950 457.950 88.050 458.550 ;
        RECT 89.550 459.300 93.150 460.200 ;
        RECT 101.850 460.200 103.650 467.250 ;
        RECT 106.350 461.400 108.150 467.250 ;
        RECT 112.650 464.400 114.450 467.250 ;
        RECT 115.650 464.400 117.450 467.250 ;
        RECT 118.650 464.400 120.450 467.250 ;
        RECT 101.850 459.300 105.450 460.200 ;
        RECT 86.100 453.150 87.900 454.950 ;
        RECT 85.950 451.050 88.050 453.150 ;
        RECT 89.550 451.950 90.750 459.300 ;
        RECT 92.100 453.150 93.900 454.950 ;
        RECT 101.100 453.150 102.900 454.950 ;
        RECT 88.950 449.850 91.050 451.950 ;
        RECT 91.950 451.050 94.050 453.150 ;
        RECT 100.950 451.050 103.050 453.150 ;
        RECT 104.250 451.950 105.450 459.300 ;
        RECT 115.950 457.950 117.000 464.400 ;
        RECT 122.850 461.400 124.650 467.250 ;
        RECT 127.350 460.200 129.150 467.250 ;
        RECT 136.650 461.400 138.450 467.250 ;
        RECT 125.550 459.300 129.150 460.200 ;
        RECT 137.250 459.300 138.450 461.400 ;
        RECT 139.650 462.300 141.450 467.250 ;
        RECT 142.650 463.200 144.450 467.250 ;
        RECT 145.650 462.300 147.450 467.250 ;
        RECT 139.650 460.950 147.450 462.300 ;
        RECT 151.650 461.400 153.450 467.250 ;
        RECT 152.250 459.300 153.450 461.400 ;
        RECT 154.650 462.300 156.450 467.250 ;
        RECT 157.650 463.200 159.450 467.250 ;
        RECT 160.650 462.300 162.450 467.250 ;
        RECT 166.650 464.400 168.450 467.250 ;
        RECT 169.650 464.400 171.450 467.250 ;
        RECT 172.650 464.400 174.450 467.250 ;
        RECT 154.650 460.950 162.450 462.300 ;
        RECT 115.950 455.850 118.050 457.950 ;
        RECT 107.100 453.150 108.900 454.950 ;
        RECT 103.950 449.850 106.050 451.950 ;
        RECT 106.950 451.050 109.050 453.150 ;
        RECT 112.950 452.850 115.050 454.950 ;
        RECT 113.100 451.050 114.900 452.850 ;
        RECT 79.950 443.550 84.450 444.450 ;
        RECT 79.950 442.950 82.050 443.550 ;
        RECT 89.550 441.600 90.750 449.850 ;
        RECT 104.250 441.600 105.450 449.850 ;
        RECT 115.950 448.650 117.000 455.850 ;
        RECT 118.950 452.850 121.050 454.950 ;
        RECT 122.100 453.150 123.900 454.950 ;
        RECT 119.100 451.050 120.900 452.850 ;
        RECT 121.950 451.050 124.050 453.150 ;
        RECT 125.550 451.950 126.750 459.300 ;
        RECT 137.250 458.250 141.000 459.300 ;
        RECT 152.250 458.250 156.000 459.300 ;
        RECT 139.950 454.950 141.150 458.250 ;
        RECT 143.100 456.150 144.900 457.950 ;
        RECT 128.100 453.150 129.900 454.950 ;
        RECT 124.950 449.850 127.050 451.950 ;
        RECT 127.950 451.050 130.050 453.150 ;
        RECT 139.950 452.850 142.050 454.950 ;
        RECT 142.950 454.050 145.050 456.150 ;
        RECT 154.950 454.950 156.150 458.250 ;
        RECT 169.950 457.950 171.000 464.400 ;
        RECT 178.650 461.400 180.450 467.250 ;
        RECT 179.250 459.300 180.450 461.400 ;
        RECT 181.650 462.300 183.450 467.250 ;
        RECT 184.650 463.200 186.450 467.250 ;
        RECT 187.650 462.300 189.450 467.250 ;
        RECT 181.650 460.950 189.450 462.300 ;
        RECT 191.850 461.400 193.650 467.250 ;
        RECT 196.350 460.200 198.150 467.250 ;
        RECT 205.650 461.400 207.450 467.250 ;
        RECT 208.650 461.400 210.450 467.250 ;
        RECT 212.850 461.400 214.650 467.250 ;
        RECT 194.550 459.300 198.150 460.200 ;
        RECT 179.250 458.250 183.000 459.300 ;
        RECT 158.100 456.150 159.900 457.950 ;
        RECT 145.950 452.850 148.050 454.950 ;
        RECT 154.950 452.850 157.050 454.950 ;
        RECT 157.950 454.050 160.050 456.150 ;
        RECT 169.950 455.850 172.050 457.950 ;
        RECT 160.950 452.850 163.050 454.950 ;
        RECT 166.950 452.850 169.050 454.950 ;
        RECT 136.950 449.850 139.050 451.950 ;
        RECT 114.450 447.600 117.000 448.650 ;
        RECT 79.800 435.750 81.600 441.600 ;
        RECT 86.550 435.750 88.350 441.600 ;
        RECT 89.550 435.750 91.350 441.600 ;
        RECT 92.550 435.750 94.350 441.600 ;
        RECT 100.650 435.750 102.450 441.600 ;
        RECT 103.650 435.750 105.450 441.600 ;
        RECT 106.650 435.750 108.450 441.600 ;
        RECT 114.450 435.750 116.250 447.600 ;
        RECT 118.650 435.750 120.450 447.600 ;
        RECT 125.550 441.600 126.750 449.850 ;
        RECT 137.250 448.050 139.050 449.850 ;
        RECT 140.850 447.600 142.050 452.850 ;
        RECT 146.100 451.050 147.900 452.850 ;
        RECT 151.950 449.850 154.050 451.950 ;
        RECT 152.250 448.050 154.050 449.850 ;
        RECT 155.850 447.600 157.050 452.850 ;
        RECT 161.100 451.050 162.900 452.850 ;
        RECT 167.100 451.050 168.900 452.850 ;
        RECT 169.950 448.650 171.000 455.850 ;
        RECT 181.950 454.950 183.150 458.250 ;
        RECT 185.100 456.150 186.900 457.950 ;
        RECT 172.950 452.850 175.050 454.950 ;
        RECT 181.950 452.850 184.050 454.950 ;
        RECT 184.950 454.050 187.050 456.150 ;
        RECT 187.950 452.850 190.050 454.950 ;
        RECT 191.100 453.150 192.900 454.950 ;
        RECT 173.100 451.050 174.900 452.850 ;
        RECT 178.950 449.850 181.050 451.950 ;
        RECT 168.450 447.600 171.000 448.650 ;
        RECT 179.250 448.050 181.050 449.850 ;
        RECT 182.850 447.600 184.050 452.850 ;
        RECT 188.100 451.050 189.900 452.850 ;
        RECT 190.950 451.050 193.050 453.150 ;
        RECT 194.550 451.950 195.750 459.300 ;
        RECT 206.400 454.950 207.600 461.400 ;
        RECT 217.350 460.200 219.150 467.250 ;
        RECT 224.850 461.400 226.650 467.250 ;
        RECT 229.350 460.200 231.150 467.250 ;
        RECT 236.550 464.400 238.350 467.250 ;
        RECT 215.550 459.300 219.150 460.200 ;
        RECT 227.550 459.300 231.150 460.200 ;
        RECT 237.150 460.500 238.350 464.400 ;
        RECT 239.850 461.400 241.650 467.250 ;
        RECT 242.850 461.400 244.650 467.250 ;
        RECT 248.550 462.300 250.350 467.250 ;
        RECT 251.550 463.200 253.350 467.250 ;
        RECT 254.550 462.300 256.350 467.250 ;
        RECT 237.150 459.600 242.250 460.500 ;
        RECT 209.100 456.150 210.900 457.950 ;
        RECT 197.100 453.150 198.900 454.950 ;
        RECT 193.950 449.850 196.050 451.950 ;
        RECT 196.950 451.050 199.050 453.150 ;
        RECT 205.950 452.850 208.050 454.950 ;
        RECT 208.950 454.050 211.050 456.150 ;
        RECT 212.100 453.150 213.900 454.950 ;
        RECT 122.550 435.750 124.350 441.600 ;
        RECT 125.550 435.750 127.350 441.600 ;
        RECT 128.550 435.750 130.350 441.600 ;
        RECT 137.400 435.750 139.200 441.600 ;
        RECT 140.700 435.750 142.500 447.600 ;
        RECT 144.900 435.750 146.700 447.600 ;
        RECT 152.400 435.750 154.200 441.600 ;
        RECT 155.700 435.750 157.500 447.600 ;
        RECT 159.900 435.750 161.700 447.600 ;
        RECT 168.450 435.750 170.250 447.600 ;
        RECT 172.650 435.750 174.450 447.600 ;
        RECT 179.400 435.750 181.200 441.600 ;
        RECT 182.700 435.750 184.500 447.600 ;
        RECT 186.900 435.750 188.700 447.600 ;
        RECT 194.550 441.600 195.750 449.850 ;
        RECT 206.400 447.600 207.600 452.850 ;
        RECT 211.950 451.050 214.050 453.150 ;
        RECT 215.550 451.950 216.750 459.300 ;
        RECT 218.100 453.150 219.900 454.950 ;
        RECT 224.100 453.150 225.900 454.950 ;
        RECT 214.950 449.850 217.050 451.950 ;
        RECT 217.950 451.050 220.050 453.150 ;
        RECT 223.950 451.050 226.050 453.150 ;
        RECT 227.550 451.950 228.750 459.300 ;
        RECT 240.000 458.700 242.250 459.600 ;
        RECT 230.100 453.150 231.900 454.950 ;
        RECT 226.950 449.850 229.050 451.950 ;
        RECT 229.950 451.050 232.050 453.150 ;
        RECT 235.950 452.850 238.050 454.950 ;
        RECT 236.100 451.050 237.900 452.850 ;
        RECT 240.000 450.300 241.050 458.700 ;
        RECT 243.150 454.950 244.350 461.400 ;
        RECT 248.550 460.950 256.350 462.300 ;
        RECT 257.550 461.400 259.350 467.250 ;
        RECT 263.550 462.300 265.350 467.250 ;
        RECT 266.550 463.200 268.350 467.250 ;
        RECT 269.550 462.300 271.350 467.250 ;
        RECT 257.550 459.300 258.750 461.400 ;
        RECT 263.550 460.950 271.350 462.300 ;
        RECT 272.550 461.400 274.350 467.250 ;
        RECT 278.550 464.400 280.350 467.250 ;
        RECT 281.550 464.400 283.350 467.250 ;
        RECT 284.550 464.400 286.350 467.250 ;
        RECT 272.550 459.300 273.750 461.400 ;
        RECT 255.000 458.250 258.750 459.300 ;
        RECT 270.000 458.250 273.750 459.300 ;
        RECT 251.100 456.150 252.900 457.950 ;
        RECT 241.950 452.850 244.350 454.950 ;
        RECT 247.950 452.850 250.050 454.950 ;
        RECT 250.950 454.050 253.050 456.150 ;
        RECT 254.850 454.950 256.050 458.250 ;
        RECT 266.100 456.150 267.900 457.950 ;
        RECT 253.950 452.850 256.050 454.950 ;
        RECT 262.950 452.850 265.050 454.950 ;
        RECT 265.950 454.050 268.050 456.150 ;
        RECT 269.850 454.950 271.050 458.250 ;
        RECT 282.000 457.950 283.050 464.400 ;
        RECT 291.000 461.400 292.800 467.250 ;
        RECT 295.200 463.050 297.000 467.250 ;
        RECT 298.500 464.400 300.300 467.250 ;
        RECT 305.550 464.400 307.350 467.250 ;
        RECT 308.550 464.400 310.350 467.250 ;
        RECT 295.200 461.400 300.900 463.050 ;
        RECT 271.950 456.450 274.050 457.050 ;
        RECT 271.950 455.550 276.450 456.450 ;
        RECT 280.950 455.850 283.050 457.950 ;
        RECT 290.100 456.150 291.900 457.950 ;
        RECT 271.950 454.950 274.050 455.550 ;
        RECT 268.950 452.850 271.050 454.950 ;
        RECT 191.550 435.750 193.350 441.600 ;
        RECT 194.550 435.750 196.350 441.600 ;
        RECT 197.550 435.750 199.350 441.600 ;
        RECT 205.650 435.750 207.450 447.600 ;
        RECT 208.650 435.750 210.450 447.600 ;
        RECT 215.550 441.600 216.750 449.850 ;
        RECT 227.550 441.600 228.750 449.850 ;
        RECT 240.000 449.400 242.250 450.300 ;
        RECT 236.550 448.500 242.250 449.400 ;
        RECT 236.550 441.600 237.750 448.500 ;
        RECT 243.150 447.600 244.350 452.850 ;
        RECT 248.100 451.050 249.900 452.850 ;
        RECT 253.950 447.600 255.150 452.850 ;
        RECT 256.950 449.850 259.050 451.950 ;
        RECT 263.100 451.050 264.900 452.850 ;
        RECT 256.950 448.050 258.750 449.850 ;
        RECT 268.950 447.600 270.150 452.850 ;
        RECT 271.950 449.850 274.050 451.950 ;
        RECT 271.950 448.050 273.750 449.850 ;
        RECT 275.550 448.050 276.450 455.550 ;
        RECT 277.950 452.850 280.050 454.950 ;
        RECT 278.100 451.050 279.900 452.850 ;
        RECT 282.000 448.650 283.050 455.850 ;
        RECT 283.950 452.850 286.050 454.950 ;
        RECT 289.950 454.050 292.050 456.150 ;
        RECT 292.950 455.850 295.050 457.950 ;
        RECT 296.100 456.150 297.900 457.950 ;
        RECT 293.100 454.050 294.900 455.850 ;
        RECT 295.950 454.050 298.050 456.150 ;
        RECT 299.700 454.950 300.900 461.400 ;
        RECT 304.950 455.850 307.050 457.950 ;
        RECT 308.400 456.150 309.600 464.400 ;
        RECT 314.550 462.300 316.350 467.250 ;
        RECT 317.550 463.200 319.350 467.250 ;
        RECT 320.550 462.300 322.350 467.250 ;
        RECT 314.550 460.950 322.350 462.300 ;
        RECT 323.550 461.400 325.350 467.250 ;
        RECT 329.550 464.400 331.350 467.250 ;
        RECT 332.550 464.400 334.350 467.250 ;
        RECT 335.550 464.400 337.350 467.250 ;
        RECT 323.550 459.300 324.750 461.400 ;
        RECT 321.000 458.250 324.750 459.300 ;
        RECT 317.100 456.150 318.900 457.950 ;
        RECT 298.950 452.850 301.050 454.950 ;
        RECT 305.100 454.050 306.900 455.850 ;
        RECT 307.950 454.050 310.050 456.150 ;
        RECT 284.100 451.050 285.900 452.850 ;
        RECT 212.550 435.750 214.350 441.600 ;
        RECT 215.550 435.750 217.350 441.600 ;
        RECT 218.550 435.750 220.350 441.600 ;
        RECT 224.550 435.750 226.350 441.600 ;
        RECT 227.550 435.750 229.350 441.600 ;
        RECT 230.550 435.750 232.350 441.600 ;
        RECT 236.550 435.750 238.350 441.600 ;
        RECT 239.850 435.750 241.650 447.600 ;
        RECT 242.850 435.750 244.650 447.600 ;
        RECT 249.300 435.750 251.100 447.600 ;
        RECT 253.500 435.750 255.300 447.600 ;
        RECT 256.800 435.750 258.600 441.600 ;
        RECT 264.300 435.750 266.100 447.600 ;
        RECT 268.500 435.750 270.300 447.600 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 282.000 447.600 284.550 448.650 ;
        RECT 299.700 447.600 300.900 452.850 ;
        RECT 271.800 435.750 273.600 441.600 ;
        RECT 278.550 435.750 280.350 447.600 ;
        RECT 282.750 435.750 284.550 447.600 ;
        RECT 290.550 446.700 298.350 447.600 ;
        RECT 290.550 435.750 292.350 446.700 ;
        RECT 293.550 435.750 295.350 445.800 ;
        RECT 296.550 435.750 298.350 446.700 ;
        RECT 299.550 435.750 301.350 447.600 ;
        RECT 308.400 441.600 309.600 454.050 ;
        RECT 313.950 452.850 316.050 454.950 ;
        RECT 316.950 454.050 319.050 456.150 ;
        RECT 320.850 454.950 322.050 458.250 ;
        RECT 333.000 457.950 334.050 464.400 ;
        RECT 344.850 460.200 346.650 467.250 ;
        RECT 349.350 461.400 351.150 467.250 ;
        RECT 353.550 462.300 355.350 467.250 ;
        RECT 356.550 463.200 358.350 467.250 ;
        RECT 359.550 462.300 361.350 467.250 ;
        RECT 353.550 460.950 361.350 462.300 ;
        RECT 362.550 461.400 364.350 467.250 ;
        RECT 368.550 464.400 370.350 467.250 ;
        RECT 371.550 464.400 373.350 467.250 ;
        RECT 344.850 459.300 348.450 460.200 ;
        RECT 362.550 459.300 363.750 461.400 ;
        RECT 331.950 455.850 334.050 457.950 ;
        RECT 319.950 452.850 322.050 454.950 ;
        RECT 328.950 452.850 331.050 454.950 ;
        RECT 314.100 451.050 315.900 452.850 ;
        RECT 319.950 447.600 321.150 452.850 ;
        RECT 322.950 449.850 325.050 451.950 ;
        RECT 329.100 451.050 330.900 452.850 ;
        RECT 322.950 448.050 324.750 449.850 ;
        RECT 333.000 448.650 334.050 455.850 ;
        RECT 334.950 452.850 337.050 454.950 ;
        RECT 344.100 453.150 345.900 454.950 ;
        RECT 335.100 451.050 336.900 452.850 ;
        RECT 343.950 451.050 346.050 453.150 ;
        RECT 347.250 451.950 348.450 459.300 ;
        RECT 360.000 458.250 363.750 459.300 ;
        RECT 356.100 456.150 357.900 457.950 ;
        RECT 350.100 453.150 351.900 454.950 ;
        RECT 346.950 449.850 349.050 451.950 ;
        RECT 349.950 451.050 352.050 453.150 ;
        RECT 352.950 452.850 355.050 454.950 ;
        RECT 355.950 454.050 358.050 456.150 ;
        RECT 359.850 454.950 361.050 458.250 ;
        RECT 367.950 455.850 370.050 457.950 ;
        RECT 371.400 456.150 372.600 464.400 ;
        RECT 377.550 462.300 379.350 467.250 ;
        RECT 380.550 463.200 382.350 467.250 ;
        RECT 383.550 462.300 385.350 467.250 ;
        RECT 377.550 460.950 385.350 462.300 ;
        RECT 386.550 461.400 388.350 467.250 ;
        RECT 392.550 464.400 394.350 467.250 ;
        RECT 386.550 459.300 387.750 461.400 ;
        RECT 393.150 460.500 394.350 464.400 ;
        RECT 395.850 461.400 397.650 467.250 ;
        RECT 398.850 461.400 400.650 467.250 ;
        RECT 404.850 461.400 406.650 467.250 ;
        RECT 393.150 459.600 398.250 460.500 ;
        RECT 384.000 458.250 387.750 459.300 ;
        RECT 396.000 458.700 398.250 459.600 ;
        RECT 380.100 456.150 381.900 457.950 ;
        RECT 358.950 452.850 361.050 454.950 ;
        RECT 368.100 454.050 369.900 455.850 ;
        RECT 370.950 454.050 373.050 456.150 ;
        RECT 353.100 451.050 354.900 452.850 ;
        RECT 333.000 447.600 335.550 448.650 ;
        RECT 305.550 435.750 307.350 441.600 ;
        RECT 308.550 435.750 310.350 441.600 ;
        RECT 315.300 435.750 317.100 447.600 ;
        RECT 319.500 435.750 321.300 447.600 ;
        RECT 322.800 435.750 324.600 441.600 ;
        RECT 329.550 435.750 331.350 447.600 ;
        RECT 333.750 435.750 335.550 447.600 ;
        RECT 347.250 441.600 348.450 449.850 ;
        RECT 358.950 447.600 360.150 452.850 ;
        RECT 361.950 449.850 364.050 451.950 ;
        RECT 361.950 448.050 363.750 449.850 ;
        RECT 343.650 435.750 345.450 441.600 ;
        RECT 346.650 435.750 348.450 441.600 ;
        RECT 349.650 435.750 351.450 441.600 ;
        RECT 354.300 435.750 356.100 447.600 ;
        RECT 358.500 435.750 360.300 447.600 ;
        RECT 371.400 441.600 372.600 454.050 ;
        RECT 376.950 452.850 379.050 454.950 ;
        RECT 379.950 454.050 382.050 456.150 ;
        RECT 383.850 454.950 385.050 458.250 ;
        RECT 382.950 452.850 385.050 454.950 ;
        RECT 391.950 452.850 394.050 454.950 ;
        RECT 377.100 451.050 378.900 452.850 ;
        RECT 382.950 447.600 384.150 452.850 ;
        RECT 385.950 449.850 388.050 451.950 ;
        RECT 392.100 451.050 393.900 452.850 ;
        RECT 396.000 450.300 397.050 458.700 ;
        RECT 399.150 454.950 400.350 461.400 ;
        RECT 409.350 460.200 411.150 467.250 ;
        RECT 407.550 459.300 411.150 460.200 ;
        RECT 417.150 461.400 418.950 467.250 ;
        RECT 420.150 464.400 421.950 467.250 ;
        RECT 424.950 465.300 426.750 467.250 ;
        RECT 423.000 464.400 426.750 465.300 ;
        RECT 429.450 464.400 431.250 467.250 ;
        RECT 432.750 464.400 434.550 467.250 ;
        RECT 436.650 464.400 438.450 467.250 ;
        RECT 440.850 464.400 442.650 467.250 ;
        RECT 445.350 464.400 447.150 467.250 ;
        RECT 423.000 463.500 424.050 464.400 ;
        RECT 421.950 461.400 424.050 463.500 ;
        RECT 432.750 462.600 433.800 464.400 ;
        RECT 397.950 452.850 400.350 454.950 ;
        RECT 404.100 453.150 405.900 454.950 ;
        RECT 385.950 448.050 387.750 449.850 ;
        RECT 396.000 449.400 398.250 450.300 ;
        RECT 392.550 448.500 398.250 449.400 ;
        RECT 361.800 435.750 363.600 441.600 ;
        RECT 368.550 435.750 370.350 441.600 ;
        RECT 371.550 435.750 373.350 441.600 ;
        RECT 378.300 435.750 380.100 447.600 ;
        RECT 382.500 435.750 384.300 447.600 ;
        RECT 392.550 441.600 393.750 448.500 ;
        RECT 399.150 447.600 400.350 452.850 ;
        RECT 403.950 451.050 406.050 453.150 ;
        RECT 407.550 451.950 408.750 459.300 ;
        RECT 410.100 453.150 411.900 454.950 ;
        RECT 406.950 449.850 409.050 451.950 ;
        RECT 409.950 451.050 412.050 453.150 ;
        RECT 385.800 435.750 387.600 441.600 ;
        RECT 392.550 435.750 394.350 441.600 ;
        RECT 395.850 435.750 397.650 447.600 ;
        RECT 398.850 435.750 400.650 447.600 ;
        RECT 407.550 441.600 408.750 449.850 ;
        RECT 417.150 448.800 418.050 461.400 ;
        RECT 425.550 460.800 427.350 462.600 ;
        RECT 428.850 461.550 433.800 462.600 ;
        RECT 441.300 463.500 442.350 464.400 ;
        RECT 441.300 462.300 445.050 463.500 ;
        RECT 428.850 460.800 430.650 461.550 ;
        RECT 425.850 459.900 426.900 460.800 ;
        RECT 436.050 460.200 437.850 462.000 ;
        RECT 442.950 461.400 445.050 462.300 ;
        RECT 448.650 461.400 450.450 467.250 ;
        RECT 454.650 464.400 456.450 467.250 ;
        RECT 457.650 464.400 459.450 467.250 ;
        RECT 460.650 464.400 462.450 467.250 ;
        RECT 467.700 464.400 469.500 467.250 ;
        RECT 436.050 459.900 436.950 460.200 ;
        RECT 425.850 459.000 436.950 459.900 ;
        RECT 449.250 459.150 450.450 461.400 ;
        RECT 425.850 457.800 426.900 459.000 ;
        RECT 420.000 456.600 426.900 457.800 ;
        RECT 420.000 455.850 420.900 456.600 ;
        RECT 425.100 456.000 426.900 456.600 ;
        RECT 419.100 454.050 420.900 455.850 ;
        RECT 422.100 454.950 423.900 455.700 ;
        RECT 436.050 454.950 436.950 459.000 ;
        RECT 445.950 457.050 450.450 459.150 ;
        RECT 444.150 455.250 448.050 457.050 ;
        RECT 445.950 454.950 448.050 455.250 ;
        RECT 422.100 453.900 430.050 454.950 ;
        RECT 427.950 452.850 430.050 453.900 ;
        RECT 433.950 452.850 436.950 454.950 ;
        RECT 426.450 449.100 428.250 449.400 ;
        RECT 426.450 448.800 434.850 449.100 ;
        RECT 417.150 448.200 434.850 448.800 ;
        RECT 417.150 447.600 428.250 448.200 ;
        RECT 404.550 435.750 406.350 441.600 ;
        RECT 407.550 435.750 409.350 441.600 ;
        RECT 410.550 435.750 412.350 441.600 ;
        RECT 417.150 435.750 418.950 447.600 ;
        RECT 431.250 446.700 433.050 447.300 ;
        RECT 425.550 445.500 433.050 446.700 ;
        RECT 433.950 446.100 434.850 448.200 ;
        RECT 436.050 448.200 436.950 452.850 ;
        RECT 446.250 449.400 448.050 451.200 ;
        RECT 442.950 448.200 447.150 449.400 ;
        RECT 436.050 447.300 442.050 448.200 ;
        RECT 442.950 447.300 445.050 448.200 ;
        RECT 449.250 447.600 450.450 457.050 ;
        RECT 457.950 457.950 459.000 464.400 ;
        RECT 471.000 463.050 472.800 467.250 ;
        RECT 467.100 461.400 472.800 463.050 ;
        RECT 475.200 461.400 477.000 467.250 ;
        RECT 479.550 464.400 481.350 467.250 ;
        RECT 482.550 464.400 484.350 467.250 ;
        RECT 485.550 464.400 487.350 467.250 ;
        RECT 457.950 455.850 460.050 457.950 ;
        RECT 454.950 452.850 457.050 454.950 ;
        RECT 455.100 451.050 456.900 452.850 ;
        RECT 457.950 448.650 459.000 455.850 ;
        RECT 467.100 454.950 468.300 461.400 ;
        RECT 483.000 457.950 484.050 464.400 ;
        RECT 470.100 456.150 471.900 457.950 ;
        RECT 460.950 452.850 463.050 454.950 ;
        RECT 466.950 452.850 469.050 454.950 ;
        RECT 469.950 454.050 472.050 456.150 ;
        RECT 472.950 455.850 475.050 457.950 ;
        RECT 476.100 456.150 477.900 457.950 ;
        RECT 473.100 454.050 474.900 455.850 ;
        RECT 475.950 454.050 478.050 456.150 ;
        RECT 481.950 455.850 484.050 457.950 ;
        RECT 478.950 452.850 481.050 454.950 ;
        RECT 461.100 451.050 462.900 452.850 ;
        RECT 441.150 446.400 442.050 447.300 ;
        RECT 438.450 446.100 440.250 446.400 ;
        RECT 425.550 444.600 426.750 445.500 ;
        RECT 433.950 445.200 440.250 446.100 ;
        RECT 438.450 444.600 440.250 445.200 ;
        RECT 441.150 444.600 443.850 446.400 ;
        RECT 421.950 442.500 426.750 444.600 ;
        RECT 429.150 442.500 436.050 444.300 ;
        RECT 425.550 441.600 426.750 442.500 ;
        RECT 420.150 435.750 421.950 441.600 ;
        RECT 425.250 435.750 427.050 441.600 ;
        RECT 430.050 435.750 431.850 441.600 ;
        RECT 433.050 435.750 434.850 442.500 ;
        RECT 441.150 441.600 445.050 443.700 ;
        RECT 436.950 435.750 438.750 441.600 ;
        RECT 441.150 435.750 442.950 441.600 ;
        RECT 445.650 435.750 447.450 438.600 ;
        RECT 448.650 435.750 450.450 447.600 ;
        RECT 456.450 447.600 459.000 448.650 ;
        RECT 467.100 447.600 468.300 452.850 ;
        RECT 479.100 451.050 480.900 452.850 ;
        RECT 483.000 448.650 484.050 455.850 ;
        RECT 492.150 461.400 493.950 467.250 ;
        RECT 495.150 464.400 496.950 467.250 ;
        RECT 499.950 465.300 501.750 467.250 ;
        RECT 498.000 464.400 501.750 465.300 ;
        RECT 504.450 464.400 506.250 467.250 ;
        RECT 507.750 464.400 509.550 467.250 ;
        RECT 511.650 464.400 513.450 467.250 ;
        RECT 515.850 464.400 517.650 467.250 ;
        RECT 520.350 464.400 522.150 467.250 ;
        RECT 498.000 463.500 499.050 464.400 ;
        RECT 496.950 461.400 499.050 463.500 ;
        RECT 507.750 462.600 508.800 464.400 ;
        RECT 484.950 452.850 487.050 454.950 ;
        RECT 485.100 451.050 486.900 452.850 ;
        RECT 492.150 448.800 493.050 461.400 ;
        RECT 500.550 460.800 502.350 462.600 ;
        RECT 503.850 461.550 508.800 462.600 ;
        RECT 516.300 463.500 517.350 464.400 ;
        RECT 516.300 462.300 520.050 463.500 ;
        RECT 503.850 460.800 505.650 461.550 ;
        RECT 500.850 459.900 501.900 460.800 ;
        RECT 511.050 460.200 512.850 462.000 ;
        RECT 517.950 461.400 520.050 462.300 ;
        RECT 523.650 461.400 525.450 467.250 ;
        RECT 511.050 459.900 511.950 460.200 ;
        RECT 500.850 459.000 511.950 459.900 ;
        RECT 524.250 459.150 525.450 461.400 ;
        RECT 500.850 457.800 501.900 459.000 ;
        RECT 495.000 456.600 501.900 457.800 ;
        RECT 495.000 455.850 495.900 456.600 ;
        RECT 500.100 456.000 501.900 456.600 ;
        RECT 494.100 454.050 495.900 455.850 ;
        RECT 497.100 454.950 498.900 455.700 ;
        RECT 511.050 454.950 511.950 459.000 ;
        RECT 520.950 457.050 525.450 459.150 ;
        RECT 519.150 455.250 523.050 457.050 ;
        RECT 520.950 454.950 523.050 455.250 ;
        RECT 497.100 453.900 505.050 454.950 ;
        RECT 502.950 452.850 505.050 453.900 ;
        RECT 508.950 452.850 511.950 454.950 ;
        RECT 501.450 449.100 503.250 449.400 ;
        RECT 501.450 448.800 509.850 449.100 ;
        RECT 483.000 447.600 485.550 448.650 ;
        RECT 456.450 435.750 458.250 447.600 ;
        RECT 460.650 435.750 462.450 447.600 ;
        RECT 466.650 435.750 468.450 447.600 ;
        RECT 469.650 446.700 477.450 447.600 ;
        RECT 469.650 435.750 471.450 446.700 ;
        RECT 472.650 435.750 474.450 445.800 ;
        RECT 475.650 435.750 477.450 446.700 ;
        RECT 479.550 435.750 481.350 447.600 ;
        RECT 483.750 435.750 485.550 447.600 ;
        RECT 492.150 448.200 509.850 448.800 ;
        RECT 492.150 447.600 503.250 448.200 ;
        RECT 492.150 435.750 493.950 447.600 ;
        RECT 506.250 446.700 508.050 447.300 ;
        RECT 500.550 445.500 508.050 446.700 ;
        RECT 508.950 446.100 509.850 448.200 ;
        RECT 511.050 448.200 511.950 452.850 ;
        RECT 521.250 449.400 523.050 451.200 ;
        RECT 517.950 448.200 522.150 449.400 ;
        RECT 511.050 447.300 517.050 448.200 ;
        RECT 517.950 447.300 520.050 448.200 ;
        RECT 524.250 447.600 525.450 457.050 ;
        RECT 516.150 446.400 517.050 447.300 ;
        RECT 513.450 446.100 515.250 446.400 ;
        RECT 500.550 444.600 501.750 445.500 ;
        RECT 508.950 445.200 515.250 446.100 ;
        RECT 513.450 444.600 515.250 445.200 ;
        RECT 516.150 444.600 518.850 446.400 ;
        RECT 496.950 442.500 501.750 444.600 ;
        RECT 504.150 442.500 511.050 444.300 ;
        RECT 500.550 441.600 501.750 442.500 ;
        RECT 495.150 435.750 496.950 441.600 ;
        RECT 500.250 435.750 502.050 441.600 ;
        RECT 505.050 435.750 506.850 441.600 ;
        RECT 508.050 435.750 509.850 442.500 ;
        RECT 516.150 441.600 520.050 443.700 ;
        RECT 511.950 435.750 513.750 441.600 ;
        RECT 516.150 435.750 517.950 441.600 ;
        RECT 520.650 435.750 522.450 438.600 ;
        RECT 523.650 435.750 525.450 447.600 ;
        RECT 528.150 461.400 529.950 467.250 ;
        RECT 531.150 464.400 532.950 467.250 ;
        RECT 535.950 465.300 537.750 467.250 ;
        RECT 534.000 464.400 537.750 465.300 ;
        RECT 540.450 464.400 542.250 467.250 ;
        RECT 543.750 464.400 545.550 467.250 ;
        RECT 547.650 464.400 549.450 467.250 ;
        RECT 551.850 464.400 553.650 467.250 ;
        RECT 556.350 464.400 558.150 467.250 ;
        RECT 534.000 463.500 535.050 464.400 ;
        RECT 532.950 461.400 535.050 463.500 ;
        RECT 543.750 462.600 544.800 464.400 ;
        RECT 528.150 448.800 529.050 461.400 ;
        RECT 536.550 460.800 538.350 462.600 ;
        RECT 539.850 461.550 544.800 462.600 ;
        RECT 552.300 463.500 553.350 464.400 ;
        RECT 552.300 462.300 556.050 463.500 ;
        RECT 539.850 460.800 541.650 461.550 ;
        RECT 536.850 459.900 537.900 460.800 ;
        RECT 547.050 460.200 548.850 462.000 ;
        RECT 553.950 461.400 556.050 462.300 ;
        RECT 559.650 461.400 561.450 467.250 ;
        RECT 563.550 464.400 565.350 467.250 ;
        RECT 566.550 464.400 568.350 467.250 ;
        RECT 569.550 464.400 571.350 467.250 ;
        RECT 547.050 459.900 547.950 460.200 ;
        RECT 536.850 459.000 547.950 459.900 ;
        RECT 560.250 459.150 561.450 461.400 ;
        RECT 536.850 457.800 537.900 459.000 ;
        RECT 531.000 456.600 537.900 457.800 ;
        RECT 531.000 455.850 531.900 456.600 ;
        RECT 536.100 456.000 537.900 456.600 ;
        RECT 530.100 454.050 531.900 455.850 ;
        RECT 533.100 454.950 534.900 455.700 ;
        RECT 547.050 454.950 547.950 459.000 ;
        RECT 556.950 457.050 561.450 459.150 ;
        RECT 567.000 457.950 568.050 464.400 ;
        RECT 577.650 461.400 579.450 467.250 ;
        RECT 578.250 459.300 579.450 461.400 ;
        RECT 580.650 462.300 582.450 467.250 ;
        RECT 583.650 463.200 585.450 467.250 ;
        RECT 586.650 462.300 588.450 467.250 ;
        RECT 580.650 460.950 588.450 462.300 ;
        RECT 592.650 461.400 594.450 467.250 ;
        RECT 593.250 459.300 594.450 461.400 ;
        RECT 595.650 462.300 597.450 467.250 ;
        RECT 598.650 463.200 600.450 467.250 ;
        RECT 601.650 462.300 603.450 467.250 ;
        RECT 595.650 460.950 603.450 462.300 ;
        RECT 605.550 462.300 607.350 467.250 ;
        RECT 608.550 463.200 610.350 467.250 ;
        RECT 611.550 462.300 613.350 467.250 ;
        RECT 605.550 460.950 613.350 462.300 ;
        RECT 614.550 461.400 616.350 467.250 ;
        RECT 620.550 462.300 622.350 467.250 ;
        RECT 623.550 463.200 625.350 467.250 ;
        RECT 626.550 462.300 628.350 467.250 ;
        RECT 614.550 459.300 615.750 461.400 ;
        RECT 620.550 460.950 628.350 462.300 ;
        RECT 629.550 461.400 631.350 467.250 ;
        RECT 635.550 464.400 637.350 467.250 ;
        RECT 638.550 464.400 640.350 467.250 ;
        RECT 629.550 459.300 630.750 461.400 ;
        RECT 578.250 458.250 582.000 459.300 ;
        RECT 593.250 458.250 597.000 459.300 ;
        RECT 612.000 458.250 615.750 459.300 ;
        RECT 627.000 458.250 630.750 459.300 ;
        RECT 555.150 455.250 559.050 457.050 ;
        RECT 556.950 454.950 559.050 455.250 ;
        RECT 533.100 453.900 541.050 454.950 ;
        RECT 538.950 452.850 541.050 453.900 ;
        RECT 544.950 452.850 547.950 454.950 ;
        RECT 537.450 449.100 539.250 449.400 ;
        RECT 537.450 448.800 545.850 449.100 ;
        RECT 528.150 448.200 545.850 448.800 ;
        RECT 528.150 447.600 539.250 448.200 ;
        RECT 528.150 435.750 529.950 447.600 ;
        RECT 542.250 446.700 544.050 447.300 ;
        RECT 536.550 445.500 544.050 446.700 ;
        RECT 544.950 446.100 545.850 448.200 ;
        RECT 547.050 448.200 547.950 452.850 ;
        RECT 557.250 449.400 559.050 451.200 ;
        RECT 553.950 448.200 558.150 449.400 ;
        RECT 547.050 447.300 553.050 448.200 ;
        RECT 553.950 447.300 556.050 448.200 ;
        RECT 560.250 447.600 561.450 457.050 ;
        RECT 565.950 455.850 568.050 457.950 ;
        RECT 562.950 452.850 565.050 454.950 ;
        RECT 563.100 451.050 564.900 452.850 ;
        RECT 567.000 448.650 568.050 455.850 ;
        RECT 580.950 454.950 582.150 458.250 ;
        RECT 584.100 456.150 585.900 457.950 ;
        RECT 568.950 452.850 571.050 454.950 ;
        RECT 580.950 452.850 583.050 454.950 ;
        RECT 583.950 454.050 586.050 456.150 ;
        RECT 595.950 454.950 597.150 458.250 ;
        RECT 599.100 456.150 600.900 457.950 ;
        RECT 608.100 456.150 609.900 457.950 ;
        RECT 586.950 452.850 589.050 454.950 ;
        RECT 595.950 452.850 598.050 454.950 ;
        RECT 598.950 454.050 601.050 456.150 ;
        RECT 601.950 452.850 604.050 454.950 ;
        RECT 604.950 452.850 607.050 454.950 ;
        RECT 607.950 454.050 610.050 456.150 ;
        RECT 611.850 454.950 613.050 458.250 ;
        RECT 623.100 456.150 624.900 457.950 ;
        RECT 610.950 452.850 613.050 454.950 ;
        RECT 619.950 452.850 622.050 454.950 ;
        RECT 622.950 454.050 625.050 456.150 ;
        RECT 626.850 454.950 628.050 458.250 ;
        RECT 634.950 455.850 637.050 457.950 ;
        RECT 638.400 456.150 639.600 464.400 ;
        RECT 640.950 460.950 643.050 463.050 ;
        RECT 625.950 452.850 628.050 454.950 ;
        RECT 635.100 454.050 636.900 455.850 ;
        RECT 637.950 454.050 640.050 456.150 ;
        RECT 569.100 451.050 570.900 452.850 ;
        RECT 577.950 449.850 580.050 451.950 ;
        RECT 567.000 447.600 569.550 448.650 ;
        RECT 578.250 448.050 580.050 449.850 ;
        RECT 581.850 447.600 583.050 452.850 ;
        RECT 587.100 451.050 588.900 452.850 ;
        RECT 592.950 449.850 595.050 451.950 ;
        RECT 593.250 448.050 595.050 449.850 ;
        RECT 596.850 447.600 598.050 452.850 ;
        RECT 602.100 451.050 603.900 452.850 ;
        RECT 605.100 451.050 606.900 452.850 ;
        RECT 610.950 447.600 612.150 452.850 ;
        RECT 613.950 449.850 616.050 451.950 ;
        RECT 620.100 451.050 621.900 452.850 ;
        RECT 613.950 448.050 615.750 449.850 ;
        RECT 625.950 447.600 627.150 452.850 ;
        RECT 628.950 449.850 631.050 451.950 ;
        RECT 628.950 448.050 630.750 449.850 ;
        RECT 552.150 446.400 553.050 447.300 ;
        RECT 549.450 446.100 551.250 446.400 ;
        RECT 536.550 444.600 537.750 445.500 ;
        RECT 544.950 445.200 551.250 446.100 ;
        RECT 549.450 444.600 551.250 445.200 ;
        RECT 552.150 444.600 554.850 446.400 ;
        RECT 532.950 442.500 537.750 444.600 ;
        RECT 540.150 442.500 547.050 444.300 ;
        RECT 536.550 441.600 537.750 442.500 ;
        RECT 531.150 435.750 532.950 441.600 ;
        RECT 536.250 435.750 538.050 441.600 ;
        RECT 541.050 435.750 542.850 441.600 ;
        RECT 544.050 435.750 545.850 442.500 ;
        RECT 552.150 441.600 556.050 443.700 ;
        RECT 547.950 435.750 549.750 441.600 ;
        RECT 552.150 435.750 553.950 441.600 ;
        RECT 556.650 435.750 558.450 438.600 ;
        RECT 559.650 435.750 561.450 447.600 ;
        RECT 563.550 435.750 565.350 447.600 ;
        RECT 567.750 435.750 569.550 447.600 ;
        RECT 578.400 435.750 580.200 441.600 ;
        RECT 581.700 435.750 583.500 447.600 ;
        RECT 585.900 435.750 587.700 447.600 ;
        RECT 593.400 435.750 595.200 441.600 ;
        RECT 596.700 435.750 598.500 447.600 ;
        RECT 600.900 435.750 602.700 447.600 ;
        RECT 606.300 435.750 608.100 447.600 ;
        RECT 610.500 435.750 612.300 447.600 ;
        RECT 613.800 435.750 615.600 441.600 ;
        RECT 621.300 435.750 623.100 447.600 ;
        RECT 625.500 435.750 627.300 447.600 ;
        RECT 638.400 441.600 639.600 454.050 ;
        RECT 641.550 451.050 642.450 460.950 ;
        RECT 644.700 458.400 646.500 467.250 ;
        RECT 650.100 459.000 651.900 467.250 ;
        RECT 659.550 461.400 661.350 467.250 ;
        RECT 662.850 464.400 664.650 467.250 ;
        RECT 667.350 464.400 669.150 467.250 ;
        RECT 671.550 464.400 673.350 467.250 ;
        RECT 675.450 464.400 677.250 467.250 ;
        RECT 678.750 464.400 680.550 467.250 ;
        RECT 683.250 465.300 685.050 467.250 ;
        RECT 683.250 464.400 687.000 465.300 ;
        RECT 688.050 464.400 689.850 467.250 ;
        RECT 667.650 463.500 668.700 464.400 ;
        RECT 664.950 462.300 668.700 463.500 ;
        RECT 676.200 462.600 677.250 464.400 ;
        RECT 685.950 463.500 687.000 464.400 ;
        RECT 664.950 461.400 667.050 462.300 ;
        RECT 659.550 459.150 660.750 461.400 ;
        RECT 672.150 460.200 673.950 462.000 ;
        RECT 676.200 461.550 681.150 462.600 ;
        RECT 679.350 460.800 681.150 461.550 ;
        RECT 682.650 460.800 684.450 462.600 ;
        RECT 685.950 461.400 688.050 463.500 ;
        RECT 691.050 461.400 692.850 467.250 ;
        RECT 673.050 459.900 673.950 460.200 ;
        RECT 683.100 459.900 684.150 460.800 ;
        RECT 650.100 457.350 654.600 459.000 ;
        RECT 653.400 453.150 654.600 457.350 ;
        RECT 659.550 457.050 664.050 459.150 ;
        RECT 673.050 459.000 684.150 459.900 ;
        RECT 640.950 448.950 643.050 451.050 ;
        RECT 643.950 449.850 646.050 451.950 ;
        RECT 649.950 449.850 652.050 451.950 ;
        RECT 652.950 451.050 655.050 453.150 ;
        RECT 644.100 448.050 645.900 449.850 ;
        RECT 646.950 446.850 649.050 448.950 ;
        RECT 650.250 448.050 652.050 449.850 ;
        RECT 647.100 445.050 648.900 446.850 ;
        RECT 653.700 442.800 654.750 451.050 ;
        RECT 647.700 441.900 654.750 442.800 ;
        RECT 647.700 441.600 649.350 441.900 ;
        RECT 628.800 435.750 630.600 441.600 ;
        RECT 635.550 435.750 637.350 441.600 ;
        RECT 638.550 435.750 640.350 441.600 ;
        RECT 644.550 435.750 646.350 441.600 ;
        RECT 647.550 435.750 649.350 441.600 ;
        RECT 653.550 441.600 654.750 441.900 ;
        RECT 659.550 447.600 660.750 457.050 ;
        RECT 661.950 455.250 665.850 457.050 ;
        RECT 661.950 454.950 664.050 455.250 ;
        RECT 673.050 454.950 673.950 459.000 ;
        RECT 683.100 457.800 684.150 459.000 ;
        RECT 683.100 456.600 690.000 457.800 ;
        RECT 683.100 456.000 684.900 456.600 ;
        RECT 689.100 455.850 690.000 456.600 ;
        RECT 686.100 454.950 687.900 455.700 ;
        RECT 673.050 452.850 676.050 454.950 ;
        RECT 679.950 453.900 687.900 454.950 ;
        RECT 689.100 454.050 690.900 455.850 ;
        RECT 679.950 452.850 682.050 453.900 ;
        RECT 661.950 449.400 663.750 451.200 ;
        RECT 662.850 448.200 667.050 449.400 ;
        RECT 673.050 448.200 673.950 452.850 ;
        RECT 681.750 449.100 683.550 449.400 ;
        RECT 650.550 435.750 652.350 441.000 ;
        RECT 653.550 435.750 655.350 441.600 ;
        RECT 659.550 435.750 661.350 447.600 ;
        RECT 664.950 447.300 667.050 448.200 ;
        RECT 667.950 447.300 673.950 448.200 ;
        RECT 675.150 448.800 683.550 449.100 ;
        RECT 691.950 448.800 692.850 461.400 ;
        RECT 695.550 462.300 697.350 467.250 ;
        RECT 698.550 463.200 700.350 467.250 ;
        RECT 701.550 462.300 703.350 467.250 ;
        RECT 695.550 460.950 703.350 462.300 ;
        RECT 704.550 461.400 706.350 467.250 ;
        RECT 704.550 459.300 705.750 461.400 ;
        RECT 709.950 460.950 712.050 463.050 ;
        RECT 702.000 458.250 705.750 459.300 ;
        RECT 698.100 456.150 699.900 457.950 ;
        RECT 694.950 452.850 697.050 454.950 ;
        RECT 697.950 454.050 700.050 456.150 ;
        RECT 701.850 454.950 703.050 458.250 ;
        RECT 700.950 452.850 703.050 454.950 ;
        RECT 695.100 451.050 696.900 452.850 ;
        RECT 675.150 448.200 692.850 448.800 ;
        RECT 667.950 446.400 668.850 447.300 ;
        RECT 666.150 444.600 668.850 446.400 ;
        RECT 669.750 446.100 671.550 446.400 ;
        RECT 675.150 446.100 676.050 448.200 ;
        RECT 681.750 447.600 692.850 448.200 ;
        RECT 700.950 447.600 702.150 452.850 ;
        RECT 703.950 449.850 706.050 451.950 ;
        RECT 710.550 451.050 711.450 460.950 ;
        RECT 703.950 448.050 705.750 449.850 ;
        RECT 709.950 448.950 712.050 451.050 ;
        RECT 669.750 445.200 676.050 446.100 ;
        RECT 676.950 446.700 678.750 447.300 ;
        RECT 676.950 445.500 684.450 446.700 ;
        RECT 669.750 444.600 671.550 445.200 ;
        RECT 683.250 444.600 684.450 445.500 ;
        RECT 664.950 441.600 668.850 443.700 ;
        RECT 673.950 442.500 680.850 444.300 ;
        RECT 683.250 442.500 688.050 444.600 ;
        RECT 662.550 435.750 664.350 438.600 ;
        RECT 667.050 435.750 668.850 441.600 ;
        RECT 671.250 435.750 673.050 441.600 ;
        RECT 675.150 435.750 676.950 442.500 ;
        RECT 683.250 441.600 684.450 442.500 ;
        RECT 678.150 435.750 679.950 441.600 ;
        RECT 682.950 435.750 684.750 441.600 ;
        RECT 688.050 435.750 689.850 441.600 ;
        RECT 691.050 435.750 692.850 447.600 ;
        RECT 696.300 435.750 698.100 447.600 ;
        RECT 700.500 435.750 702.300 447.600 ;
        RECT 703.800 435.750 705.600 441.600 ;
        RECT 4.650 425.400 6.450 431.250 ;
        RECT 7.650 425.400 9.450 431.250 ;
        RECT 14.400 425.400 16.200 431.250 ;
        RECT 5.400 412.950 6.600 425.400 ;
        RECT 17.700 419.400 19.500 431.250 ;
        RECT 21.900 419.400 23.700 431.250 ;
        RECT 26.550 420.600 28.350 431.250 ;
        RECT 29.550 421.500 31.350 431.250 ;
        RECT 32.550 430.500 40.350 431.250 ;
        RECT 32.550 420.600 34.350 430.500 ;
        RECT 26.550 419.700 34.350 420.600 ;
        RECT 35.550 419.400 37.350 429.600 ;
        RECT 38.550 419.400 40.350 430.500 ;
        RECT 44.550 425.400 46.350 431.250 ;
        RECT 47.550 425.400 49.350 431.250 ;
        RECT 50.550 425.400 52.350 431.250 ;
        RECT 56.550 425.400 58.350 431.250 ;
        RECT 59.550 425.400 61.350 431.250 ;
        RECT 14.250 417.150 16.050 418.950 ;
        RECT 13.950 415.050 16.050 417.150 ;
        RECT 17.850 414.150 19.050 419.400 ;
        RECT 35.400 418.500 37.200 419.400 ;
        RECT 33.150 417.600 37.200 418.500 ;
        RECT 23.100 414.150 24.900 415.950 ;
        RECT 26.250 414.150 28.050 415.950 ;
        RECT 33.150 414.150 34.050 417.600 ;
        RECT 47.550 417.150 48.750 425.400 ;
        RECT 38.100 414.150 39.900 415.950 ;
        RECT 4.950 410.850 7.050 412.950 ;
        RECT 8.100 411.150 9.900 412.950 ;
        RECT 16.950 412.050 19.050 414.150 ;
        RECT 5.400 402.600 6.600 410.850 ;
        RECT 7.950 409.050 10.050 411.150 ;
        RECT 16.950 408.750 18.150 412.050 ;
        RECT 19.950 410.850 22.050 412.950 ;
        RECT 22.950 412.050 25.050 414.150 ;
        RECT 25.950 412.050 28.050 414.150 ;
        RECT 28.950 410.850 31.050 412.950 ;
        RECT 20.100 409.050 21.900 410.850 ;
        RECT 29.250 409.050 31.050 410.850 ;
        RECT 31.950 412.050 34.050 414.150 ;
        RECT 14.250 407.700 18.000 408.750 ;
        RECT 14.250 405.600 15.450 407.700 ;
        RECT 4.650 399.750 6.450 402.600 ;
        RECT 7.650 399.750 9.450 402.600 ;
        RECT 13.650 399.750 15.450 405.600 ;
        RECT 16.650 404.700 24.450 406.050 ;
        RECT 31.950 405.600 33.000 412.050 ;
        RECT 34.950 410.850 37.050 412.950 ;
        RECT 37.950 412.050 40.050 414.150 ;
        RECT 43.950 413.850 46.050 415.950 ;
        RECT 46.950 415.050 49.050 417.150 ;
        RECT 44.100 412.050 45.900 413.850 ;
        RECT 34.950 409.050 36.750 410.850 ;
        RECT 47.550 407.700 48.750 415.050 ;
        RECT 49.950 413.850 52.050 415.950 ;
        RECT 56.100 414.150 57.900 415.950 ;
        RECT 50.100 412.050 51.900 413.850 ;
        RECT 55.950 412.050 58.050 414.150 ;
        RECT 59.700 408.300 60.900 425.400 ;
        RECT 63.150 419.400 64.950 431.250 ;
        RECT 66.150 419.400 67.950 431.250 ;
        RECT 74.400 425.400 76.200 431.250 ;
        RECT 77.700 419.400 79.500 431.250 ;
        RECT 81.900 419.400 83.700 431.250 ;
        RECT 86.550 425.400 88.350 431.250 ;
        RECT 89.550 425.400 91.350 431.250 ;
        RECT 92.550 425.400 94.350 431.250 ;
        RECT 61.950 413.850 64.050 415.950 ;
        RECT 66.150 414.150 67.350 419.400 ;
        RECT 74.250 417.150 76.050 418.950 ;
        RECT 73.950 415.050 76.050 417.150 ;
        RECT 77.850 414.150 79.050 419.400 ;
        RECT 89.550 417.150 90.750 425.400 ;
        RECT 100.650 419.400 102.450 431.250 ;
        RECT 103.650 419.400 105.450 431.250 ;
        RECT 109.650 419.400 111.450 431.250 ;
        RECT 112.650 419.400 114.450 431.250 ;
        RECT 116.550 425.400 118.350 431.250 ;
        RECT 119.550 425.400 121.350 431.250 ;
        RECT 122.550 425.400 124.350 431.250 ;
        RECT 128.550 425.400 130.350 431.250 ;
        RECT 131.550 425.400 133.350 431.250 ;
        RECT 83.100 414.150 84.900 415.950 ;
        RECT 62.100 412.050 63.900 413.850 ;
        RECT 64.950 412.050 67.350 414.150 ;
        RECT 47.550 406.800 51.150 407.700 ;
        RECT 16.650 399.750 18.450 404.700 ;
        RECT 19.650 399.750 21.450 403.800 ;
        RECT 22.650 399.750 24.450 404.700 ;
        RECT 27.000 399.750 28.800 405.600 ;
        RECT 31.200 399.750 33.000 405.600 ;
        RECT 35.400 399.750 37.200 405.600 ;
        RECT 44.850 399.750 46.650 405.600 ;
        RECT 49.350 399.750 51.150 406.800 ;
        RECT 56.550 407.100 64.050 408.300 ;
        RECT 56.550 399.750 58.350 407.100 ;
        RECT 62.250 406.500 64.050 407.100 ;
        RECT 66.150 405.600 67.350 412.050 ;
        RECT 76.950 412.050 79.050 414.150 ;
        RECT 76.950 408.750 78.150 412.050 ;
        RECT 79.950 410.850 82.050 412.950 ;
        RECT 82.950 412.050 85.050 414.150 ;
        RECT 85.950 413.850 88.050 415.950 ;
        RECT 88.950 415.050 91.050 417.150 ;
        RECT 86.100 412.050 87.900 413.850 ;
        RECT 80.100 409.050 81.900 410.850 ;
        RECT 74.250 407.700 78.000 408.750 ;
        RECT 89.550 407.700 90.750 415.050 ;
        RECT 91.950 413.850 94.050 415.950 ;
        RECT 101.400 414.150 102.600 419.400 ;
        RECT 110.400 414.150 111.600 419.400 ;
        RECT 119.550 417.150 120.750 425.400 ;
        RECT 92.100 412.050 93.900 413.850 ;
        RECT 100.950 412.050 103.050 414.150 ;
        RECT 74.250 405.600 75.450 407.700 ;
        RECT 89.550 406.800 93.150 407.700 ;
        RECT 61.050 399.750 62.850 405.600 ;
        RECT 64.050 404.100 67.350 405.600 ;
        RECT 64.050 399.750 65.850 404.100 ;
        RECT 73.650 399.750 75.450 405.600 ;
        RECT 76.650 404.700 84.450 406.050 ;
        RECT 76.650 399.750 78.450 404.700 ;
        RECT 79.650 399.750 81.450 403.800 ;
        RECT 82.650 399.750 84.450 404.700 ;
        RECT 86.850 399.750 88.650 405.600 ;
        RECT 91.350 399.750 93.150 406.800 ;
        RECT 101.400 405.600 102.600 412.050 ;
        RECT 103.950 410.850 106.050 412.950 ;
        RECT 109.950 412.050 112.050 414.150 ;
        RECT 115.950 413.850 118.050 415.950 ;
        RECT 118.950 415.050 121.050 417.150 ;
        RECT 104.100 409.050 105.900 410.850 ;
        RECT 110.400 405.600 111.600 412.050 ;
        RECT 112.950 410.850 115.050 412.950 ;
        RECT 116.100 412.050 117.900 413.850 ;
        RECT 113.100 409.050 114.900 410.850 ;
        RECT 119.550 407.700 120.750 415.050 ;
        RECT 121.950 413.850 124.050 415.950 ;
        RECT 128.100 414.150 129.900 415.950 ;
        RECT 122.100 412.050 123.900 413.850 ;
        RECT 127.950 412.050 130.050 414.150 ;
        RECT 131.700 408.300 132.900 425.400 ;
        RECT 135.150 419.400 136.950 431.250 ;
        RECT 138.150 419.400 139.950 431.250 ;
        RECT 146.400 425.400 148.200 431.250 ;
        RECT 149.700 419.400 151.500 431.250 ;
        RECT 153.900 419.400 155.700 431.250 ;
        RECT 158.550 425.400 160.350 431.250 ;
        RECT 161.550 425.400 163.350 431.250 ;
        RECT 164.550 425.400 166.350 431.250 ;
        RECT 173.400 425.400 175.200 431.250 ;
        RECT 133.950 413.850 136.050 415.950 ;
        RECT 138.150 414.150 139.350 419.400 ;
        RECT 146.250 417.150 148.050 418.950 ;
        RECT 145.950 415.050 148.050 417.150 ;
        RECT 149.850 414.150 151.050 419.400 ;
        RECT 161.550 417.150 162.750 425.400 ;
        RECT 176.700 419.400 178.500 431.250 ;
        RECT 180.900 419.400 182.700 431.250 ;
        RECT 185.550 419.400 187.350 431.250 ;
        RECT 188.550 428.400 190.350 431.250 ;
        RECT 193.050 425.400 194.850 431.250 ;
        RECT 197.250 425.400 199.050 431.250 ;
        RECT 190.950 423.300 194.850 425.400 ;
        RECT 201.150 424.500 202.950 431.250 ;
        RECT 204.150 425.400 205.950 431.250 ;
        RECT 208.950 425.400 210.750 431.250 ;
        RECT 214.050 425.400 215.850 431.250 ;
        RECT 209.250 424.500 210.450 425.400 ;
        RECT 199.950 422.700 206.850 424.500 ;
        RECT 209.250 422.400 214.050 424.500 ;
        RECT 192.150 420.600 194.850 422.400 ;
        RECT 195.750 421.800 197.550 422.400 ;
        RECT 195.750 420.900 202.050 421.800 ;
        RECT 209.250 421.500 210.450 422.400 ;
        RECT 195.750 420.600 197.550 420.900 ;
        RECT 193.950 419.700 194.850 420.600 ;
        RECT 173.250 417.150 175.050 418.950 ;
        RECT 155.100 414.150 156.900 415.950 ;
        RECT 134.100 412.050 135.900 413.850 ;
        RECT 136.950 412.050 139.350 414.150 ;
        RECT 119.550 406.800 123.150 407.700 ;
        RECT 100.650 399.750 102.450 405.600 ;
        RECT 103.650 399.750 105.450 405.600 ;
        RECT 109.650 399.750 111.450 405.600 ;
        RECT 112.650 399.750 114.450 405.600 ;
        RECT 116.850 399.750 118.650 405.600 ;
        RECT 121.350 399.750 123.150 406.800 ;
        RECT 128.550 407.100 136.050 408.300 ;
        RECT 128.550 399.750 130.350 407.100 ;
        RECT 134.250 406.500 136.050 407.100 ;
        RECT 138.150 405.600 139.350 412.050 ;
        RECT 148.950 412.050 151.050 414.150 ;
        RECT 148.950 408.750 150.150 412.050 ;
        RECT 151.950 410.850 154.050 412.950 ;
        RECT 154.950 412.050 157.050 414.150 ;
        RECT 157.950 413.850 160.050 415.950 ;
        RECT 160.950 415.050 163.050 417.150 ;
        RECT 158.100 412.050 159.900 413.850 ;
        RECT 152.100 409.050 153.900 410.850 ;
        RECT 146.250 407.700 150.000 408.750 ;
        RECT 161.550 407.700 162.750 415.050 ;
        RECT 163.950 413.850 166.050 415.950 ;
        RECT 172.950 415.050 175.050 417.150 ;
        RECT 176.850 414.150 178.050 419.400 ;
        RECT 182.100 414.150 183.900 415.950 ;
        RECT 164.100 412.050 165.900 413.850 ;
        RECT 175.950 412.050 178.050 414.150 ;
        RECT 175.950 408.750 177.150 412.050 ;
        RECT 178.950 410.850 181.050 412.950 ;
        RECT 181.950 412.050 184.050 414.150 ;
        RECT 179.100 409.050 180.900 410.850 ;
        RECT 185.550 409.950 186.750 419.400 ;
        RECT 190.950 418.800 193.050 419.700 ;
        RECT 193.950 418.800 199.950 419.700 ;
        RECT 188.850 417.600 193.050 418.800 ;
        RECT 187.950 415.800 189.750 417.600 ;
        RECT 199.050 414.150 199.950 418.800 ;
        RECT 201.150 418.800 202.050 420.900 ;
        RECT 202.950 420.300 210.450 421.500 ;
        RECT 202.950 419.700 204.750 420.300 ;
        RECT 217.050 419.400 218.850 431.250 ;
        RECT 223.350 419.400 225.150 431.250 ;
        RECT 226.350 419.400 228.150 431.250 ;
        RECT 229.650 425.400 231.450 431.250 ;
        RECT 207.750 418.800 218.850 419.400 ;
        RECT 201.150 418.200 218.850 418.800 ;
        RECT 201.150 417.900 209.550 418.200 ;
        RECT 207.750 417.600 209.550 417.900 ;
        RECT 199.050 412.050 202.050 414.150 ;
        RECT 205.950 413.100 208.050 414.150 ;
        RECT 205.950 412.050 213.900 413.100 ;
        RECT 187.950 411.750 190.050 412.050 ;
        RECT 187.950 409.950 191.850 411.750 ;
        RECT 173.250 407.700 177.000 408.750 ;
        RECT 185.550 407.850 190.050 409.950 ;
        RECT 199.050 408.000 199.950 412.050 ;
        RECT 212.100 411.300 213.900 412.050 ;
        RECT 215.100 411.150 216.900 412.950 ;
        RECT 209.100 410.400 210.900 411.000 ;
        RECT 215.100 410.400 216.000 411.150 ;
        RECT 209.100 409.200 216.000 410.400 ;
        RECT 209.100 408.000 210.150 409.200 ;
        RECT 146.250 405.600 147.450 407.700 ;
        RECT 161.550 406.800 165.150 407.700 ;
        RECT 133.050 399.750 134.850 405.600 ;
        RECT 136.050 404.100 139.350 405.600 ;
        RECT 136.050 399.750 137.850 404.100 ;
        RECT 145.650 399.750 147.450 405.600 ;
        RECT 148.650 404.700 156.450 406.050 ;
        RECT 148.650 399.750 150.450 404.700 ;
        RECT 151.650 399.750 153.450 403.800 ;
        RECT 154.650 399.750 156.450 404.700 ;
        RECT 158.850 399.750 160.650 405.600 ;
        RECT 163.350 399.750 165.150 406.800 ;
        RECT 173.250 405.600 174.450 407.700 ;
        RECT 172.650 399.750 174.450 405.600 ;
        RECT 175.650 404.700 183.450 406.050 ;
        RECT 175.650 399.750 177.450 404.700 ;
        RECT 178.650 399.750 180.450 403.800 ;
        RECT 181.650 399.750 183.450 404.700 ;
        RECT 185.550 405.600 186.750 407.850 ;
        RECT 199.050 407.100 210.150 408.000 ;
        RECT 199.050 406.800 199.950 407.100 ;
        RECT 185.550 399.750 187.350 405.600 ;
        RECT 190.950 404.700 193.050 405.600 ;
        RECT 198.150 405.000 199.950 406.800 ;
        RECT 209.100 406.200 210.150 407.100 ;
        RECT 205.350 405.450 207.150 406.200 ;
        RECT 190.950 403.500 194.700 404.700 ;
        RECT 193.650 402.600 194.700 403.500 ;
        RECT 202.200 404.400 207.150 405.450 ;
        RECT 208.650 404.400 210.450 406.200 ;
        RECT 217.950 405.600 218.850 418.200 ;
        RECT 223.650 414.150 224.850 419.400 ;
        RECT 230.250 418.500 231.450 425.400 ;
        RECT 225.750 417.600 231.450 418.500 ;
        RECT 234.150 419.400 235.950 431.250 ;
        RECT 237.150 425.400 238.950 431.250 ;
        RECT 242.250 425.400 244.050 431.250 ;
        RECT 247.050 425.400 248.850 431.250 ;
        RECT 242.550 424.500 243.750 425.400 ;
        RECT 250.050 424.500 251.850 431.250 ;
        RECT 253.950 425.400 255.750 431.250 ;
        RECT 258.150 425.400 259.950 431.250 ;
        RECT 262.650 428.400 264.450 431.250 ;
        RECT 238.950 422.400 243.750 424.500 ;
        RECT 246.150 422.700 253.050 424.500 ;
        RECT 258.150 423.300 262.050 425.400 ;
        RECT 242.550 421.500 243.750 422.400 ;
        RECT 255.450 421.800 257.250 422.400 ;
        RECT 242.550 420.300 250.050 421.500 ;
        RECT 248.250 419.700 250.050 420.300 ;
        RECT 250.950 420.900 257.250 421.800 ;
        RECT 234.150 418.800 245.250 419.400 ;
        RECT 250.950 418.800 251.850 420.900 ;
        RECT 255.450 420.600 257.250 420.900 ;
        RECT 258.150 420.600 260.850 422.400 ;
        RECT 258.150 419.700 259.050 420.600 ;
        RECT 234.150 418.200 251.850 418.800 ;
        RECT 225.750 416.700 228.000 417.600 ;
        RECT 223.650 412.050 226.050 414.150 ;
        RECT 223.650 405.600 224.850 412.050 ;
        RECT 226.950 408.300 228.000 416.700 ;
        RECT 230.100 414.150 231.900 415.950 ;
        RECT 229.950 412.050 232.050 414.150 ;
        RECT 225.750 407.400 228.000 408.300 ;
        RECT 225.750 406.500 230.850 407.400 ;
        RECT 202.200 402.600 203.250 404.400 ;
        RECT 211.950 403.500 214.050 405.600 ;
        RECT 211.950 402.600 213.000 403.500 ;
        RECT 188.850 399.750 190.650 402.600 ;
        RECT 193.350 399.750 195.150 402.600 ;
        RECT 197.550 399.750 199.350 402.600 ;
        RECT 201.450 399.750 203.250 402.600 ;
        RECT 204.750 399.750 206.550 402.600 ;
        RECT 209.250 401.700 213.000 402.600 ;
        RECT 209.250 399.750 211.050 401.700 ;
        RECT 214.050 399.750 215.850 402.600 ;
        RECT 217.050 399.750 218.850 405.600 ;
        RECT 223.350 399.750 225.150 405.600 ;
        RECT 226.350 399.750 228.150 405.600 ;
        RECT 229.650 402.600 230.850 406.500 ;
        RECT 234.150 405.600 235.050 418.200 ;
        RECT 243.450 417.900 251.850 418.200 ;
        RECT 253.050 418.800 259.050 419.700 ;
        RECT 259.950 418.800 262.050 419.700 ;
        RECT 265.650 419.400 267.450 431.250 ;
        RECT 270.300 419.400 272.100 431.250 ;
        RECT 274.500 419.400 276.300 431.250 ;
        RECT 277.800 425.400 279.600 431.250 ;
        RECT 284.550 425.400 286.350 431.250 ;
        RECT 287.550 425.400 289.350 431.250 ;
        RECT 243.450 417.600 245.250 417.900 ;
        RECT 253.050 414.150 253.950 418.800 ;
        RECT 259.950 417.600 264.150 418.800 ;
        RECT 263.250 415.800 265.050 417.600 ;
        RECT 244.950 413.100 247.050 414.150 ;
        RECT 236.100 411.150 237.900 412.950 ;
        RECT 239.100 412.050 247.050 413.100 ;
        RECT 250.950 412.050 253.950 414.150 ;
        RECT 239.100 411.300 240.900 412.050 ;
        RECT 237.000 410.400 237.900 411.150 ;
        RECT 242.100 410.400 243.900 411.000 ;
        RECT 237.000 409.200 243.900 410.400 ;
        RECT 242.850 408.000 243.900 409.200 ;
        RECT 253.050 408.000 253.950 412.050 ;
        RECT 262.950 411.750 265.050 412.050 ;
        RECT 261.150 409.950 265.050 411.750 ;
        RECT 266.250 409.950 267.450 419.400 ;
        RECT 269.100 414.150 270.900 415.950 ;
        RECT 274.950 414.150 276.150 419.400 ;
        RECT 277.950 417.150 279.750 418.950 ;
        RECT 277.950 415.050 280.050 417.150 ;
        RECT 268.950 412.050 271.050 414.150 ;
        RECT 271.950 410.850 274.050 412.950 ;
        RECT 274.950 412.050 277.050 414.150 ;
        RECT 287.400 412.950 288.600 425.400 ;
        RECT 293.550 419.400 295.350 431.250 ;
        RECT 298.050 419.400 301.350 431.250 ;
        RECT 304.050 419.400 305.850 431.250 ;
        RECT 315.450 419.400 317.250 431.250 ;
        RECT 319.650 419.400 321.450 431.250 ;
        RECT 327.450 419.400 329.250 431.250 ;
        RECT 331.650 419.400 333.450 431.250 ;
        RECT 339.450 419.400 341.250 431.250 ;
        RECT 343.650 419.400 345.450 431.250 ;
        RECT 347.550 425.400 349.350 431.250 ;
        RECT 350.550 425.400 352.350 431.250 ;
        RECT 289.950 415.950 292.050 418.050 ;
        RECT 242.850 407.100 253.950 408.000 ;
        RECT 262.950 407.850 267.450 409.950 ;
        RECT 272.100 409.050 273.900 410.850 ;
        RECT 275.850 408.750 277.050 412.050 ;
        RECT 284.100 411.150 285.900 412.950 ;
        RECT 283.950 409.050 286.050 411.150 ;
        RECT 286.950 410.850 289.050 412.950 ;
        RECT 242.850 406.200 243.900 407.100 ;
        RECT 253.050 406.800 253.950 407.100 ;
        RECT 229.650 399.750 231.450 402.600 ;
        RECT 234.150 399.750 235.950 405.600 ;
        RECT 238.950 403.500 241.050 405.600 ;
        RECT 242.550 404.400 244.350 406.200 ;
        RECT 245.850 405.450 247.650 406.200 ;
        RECT 245.850 404.400 250.800 405.450 ;
        RECT 253.050 405.000 254.850 406.800 ;
        RECT 266.250 405.600 267.450 407.850 ;
        RECT 276.000 407.700 279.750 408.750 ;
        RECT 259.950 404.700 262.050 405.600 ;
        RECT 240.000 402.600 241.050 403.500 ;
        RECT 249.750 402.600 250.800 404.400 ;
        RECT 258.300 403.500 262.050 404.700 ;
        RECT 258.300 402.600 259.350 403.500 ;
        RECT 237.150 399.750 238.950 402.600 ;
        RECT 240.000 401.700 243.750 402.600 ;
        RECT 241.950 399.750 243.750 401.700 ;
        RECT 246.450 399.750 248.250 402.600 ;
        RECT 249.750 399.750 251.550 402.600 ;
        RECT 253.650 399.750 255.450 402.600 ;
        RECT 257.850 399.750 259.650 402.600 ;
        RECT 262.350 399.750 264.150 402.600 ;
        RECT 265.650 399.750 267.450 405.600 ;
        RECT 269.550 404.700 277.350 406.050 ;
        RECT 269.550 399.750 271.350 404.700 ;
        RECT 272.550 399.750 274.350 403.800 ;
        RECT 275.550 399.750 277.350 404.700 ;
        RECT 278.550 405.600 279.750 407.700 ;
        RECT 278.550 399.750 280.350 405.600 ;
        RECT 287.400 402.600 288.600 410.850 ;
        RECT 290.550 409.050 291.450 415.950 ;
        RECT 293.100 414.150 294.900 415.950 ;
        RECT 299.550 414.150 300.750 419.400 ;
        RECT 315.450 418.350 318.000 419.400 ;
        RECT 327.450 418.350 330.000 419.400 ;
        RECT 339.450 418.350 342.000 419.400 ;
        RECT 304.950 414.150 306.750 415.950 ;
        RECT 314.100 414.150 315.900 415.950 ;
        RECT 292.950 412.050 295.050 414.150 ;
        RECT 295.950 410.850 298.050 412.950 ;
        RECT 298.950 412.050 301.050 414.150 ;
        RECT 296.100 409.050 297.900 410.850 ;
        RECT 289.950 406.950 292.050 409.050 ;
        RECT 299.400 408.150 300.600 412.050 ;
        RECT 301.950 410.850 304.050 412.950 ;
        RECT 304.950 412.050 307.050 414.150 ;
        RECT 313.950 412.050 316.050 414.150 ;
        RECT 316.950 411.150 318.000 418.350 ;
        RECT 320.100 414.150 321.900 415.950 ;
        RECT 326.100 414.150 327.900 415.950 ;
        RECT 319.950 412.050 322.050 414.150 ;
        RECT 325.950 412.050 328.050 414.150 ;
        RECT 328.950 411.150 330.000 418.350 ;
        RECT 332.100 414.150 333.900 415.950 ;
        RECT 338.100 414.150 339.900 415.950 ;
        RECT 331.950 412.050 334.050 414.150 ;
        RECT 337.950 412.050 340.050 414.150 ;
        RECT 340.950 411.150 342.000 418.350 ;
        RECT 344.100 414.150 345.900 415.950 ;
        RECT 343.950 412.050 346.050 414.150 ;
        RECT 350.400 412.950 351.600 425.400 ;
        RECT 360.450 419.400 362.250 431.250 ;
        RECT 364.650 419.400 366.450 431.250 ;
        RECT 368.550 425.400 370.350 431.250 ;
        RECT 371.550 425.400 373.350 431.250 ;
        RECT 377.550 425.400 379.350 431.250 ;
        RECT 380.550 425.400 382.350 431.250 ;
        RECT 360.450 418.350 363.000 419.400 ;
        RECT 359.100 414.150 360.900 415.950 ;
        RECT 347.100 411.150 348.900 412.950 ;
        RECT 301.500 409.050 303.300 410.850 ;
        RECT 316.950 409.050 319.050 411.150 ;
        RECT 328.950 409.050 331.050 411.150 ;
        RECT 340.950 409.050 343.050 411.150 ;
        RECT 346.950 409.050 349.050 411.150 ;
        RECT 349.950 410.850 352.050 412.950 ;
        RECT 358.950 412.050 361.050 414.150 ;
        RECT 361.950 411.150 363.000 418.350 ;
        RECT 365.100 414.150 366.900 415.950 ;
        RECT 364.950 412.050 367.050 414.150 ;
        RECT 371.400 412.950 372.600 425.400 ;
        RECT 377.100 414.150 378.900 415.950 ;
        RECT 368.100 411.150 369.900 412.950 ;
        RECT 299.400 407.100 303.750 408.150 ;
        RECT 293.550 405.000 301.350 405.900 ;
        RECT 302.850 405.600 303.750 407.100 ;
        RECT 284.550 399.750 286.350 402.600 ;
        RECT 287.550 399.750 289.350 402.600 ;
        RECT 293.550 399.750 295.350 405.000 ;
        RECT 296.550 399.750 298.350 404.100 ;
        RECT 299.550 400.500 301.350 405.000 ;
        RECT 302.550 401.400 304.350 405.600 ;
        RECT 305.550 400.500 307.350 405.600 ;
        RECT 316.950 402.600 318.000 409.050 ;
        RECT 328.950 402.600 330.000 409.050 ;
        RECT 340.950 402.600 342.000 409.050 ;
        RECT 350.400 402.600 351.600 410.850 ;
        RECT 361.950 409.050 364.050 411.150 ;
        RECT 367.950 409.050 370.050 411.150 ;
        RECT 370.950 410.850 373.050 412.950 ;
        RECT 376.950 412.050 379.050 414.150 ;
        RECT 361.950 402.600 363.000 409.050 ;
        RECT 371.400 402.600 372.600 410.850 ;
        RECT 380.700 408.300 381.900 425.400 ;
        RECT 384.150 419.400 385.950 431.250 ;
        RECT 387.150 419.400 388.950 431.250 ;
        RECT 393.300 419.400 395.100 431.250 ;
        RECT 397.500 419.400 399.300 431.250 ;
        RECT 400.800 425.400 402.600 431.250 ;
        RECT 408.300 419.400 410.100 431.250 ;
        RECT 412.500 419.400 414.300 431.250 ;
        RECT 415.800 425.400 417.600 431.250 ;
        RECT 422.550 425.400 424.350 431.250 ;
        RECT 425.550 425.400 427.350 431.250 ;
        RECT 428.550 425.400 430.350 431.250 ;
        RECT 382.950 413.850 385.050 415.950 ;
        RECT 387.150 414.150 388.350 419.400 ;
        RECT 392.100 414.150 393.900 415.950 ;
        RECT 397.950 414.150 399.150 419.400 ;
        RECT 400.950 417.150 402.750 418.950 ;
        RECT 400.950 415.050 403.050 417.150 ;
        RECT 407.100 414.150 408.900 415.950 ;
        RECT 412.950 414.150 414.150 419.400 ;
        RECT 415.950 417.150 417.750 418.950 ;
        RECT 425.550 417.150 426.750 425.400 ;
        RECT 435.150 419.400 436.950 431.250 ;
        RECT 438.150 425.400 439.950 431.250 ;
        RECT 443.250 425.400 445.050 431.250 ;
        RECT 448.050 425.400 449.850 431.250 ;
        RECT 443.550 424.500 444.750 425.400 ;
        RECT 451.050 424.500 452.850 431.250 ;
        RECT 454.950 425.400 456.750 431.250 ;
        RECT 459.150 425.400 460.950 431.250 ;
        RECT 463.650 428.400 465.450 431.250 ;
        RECT 439.950 422.400 444.750 424.500 ;
        RECT 447.150 422.700 454.050 424.500 ;
        RECT 459.150 423.300 463.050 425.400 ;
        RECT 443.550 421.500 444.750 422.400 ;
        RECT 456.450 421.800 458.250 422.400 ;
        RECT 443.550 420.300 451.050 421.500 ;
        RECT 449.250 419.700 451.050 420.300 ;
        RECT 451.950 420.900 458.250 421.800 ;
        RECT 435.150 418.800 446.250 419.400 ;
        RECT 451.950 418.800 452.850 420.900 ;
        RECT 456.450 420.600 458.250 420.900 ;
        RECT 459.150 420.600 461.850 422.400 ;
        RECT 459.150 419.700 460.050 420.600 ;
        RECT 435.150 418.200 452.850 418.800 ;
        RECT 415.950 415.050 418.050 417.150 ;
        RECT 383.100 412.050 384.900 413.850 ;
        RECT 385.950 412.050 388.350 414.150 ;
        RECT 391.950 412.050 394.050 414.150 ;
        RECT 377.550 407.100 385.050 408.300 ;
        RECT 299.550 399.750 307.350 400.500 ;
        RECT 313.650 399.750 315.450 402.600 ;
        RECT 316.650 399.750 318.450 402.600 ;
        RECT 319.650 399.750 321.450 402.600 ;
        RECT 325.650 399.750 327.450 402.600 ;
        RECT 328.650 399.750 330.450 402.600 ;
        RECT 331.650 399.750 333.450 402.600 ;
        RECT 337.650 399.750 339.450 402.600 ;
        RECT 340.650 399.750 342.450 402.600 ;
        RECT 343.650 399.750 345.450 402.600 ;
        RECT 347.550 399.750 349.350 402.600 ;
        RECT 350.550 399.750 352.350 402.600 ;
        RECT 358.650 399.750 360.450 402.600 ;
        RECT 361.650 399.750 363.450 402.600 ;
        RECT 364.650 399.750 366.450 402.600 ;
        RECT 368.550 399.750 370.350 402.600 ;
        RECT 371.550 399.750 373.350 402.600 ;
        RECT 377.550 399.750 379.350 407.100 ;
        RECT 383.250 406.500 385.050 407.100 ;
        RECT 387.150 405.600 388.350 412.050 ;
        RECT 394.950 410.850 397.050 412.950 ;
        RECT 397.950 412.050 400.050 414.150 ;
        RECT 406.950 412.050 409.050 414.150 ;
        RECT 395.100 409.050 396.900 410.850 ;
        RECT 398.850 408.750 400.050 412.050 ;
        RECT 409.950 410.850 412.050 412.950 ;
        RECT 412.950 412.050 415.050 414.150 ;
        RECT 421.950 413.850 424.050 415.950 ;
        RECT 424.950 415.050 427.050 417.150 ;
        RECT 422.100 412.050 423.900 413.850 ;
        RECT 410.100 409.050 411.900 410.850 ;
        RECT 413.850 408.750 415.050 412.050 ;
        RECT 399.000 407.700 402.750 408.750 ;
        RECT 414.000 407.700 417.750 408.750 ;
        RECT 382.050 399.750 383.850 405.600 ;
        RECT 385.050 404.100 388.350 405.600 ;
        RECT 392.550 404.700 400.350 406.050 ;
        RECT 385.050 399.750 386.850 404.100 ;
        RECT 392.550 399.750 394.350 404.700 ;
        RECT 395.550 399.750 397.350 403.800 ;
        RECT 398.550 399.750 400.350 404.700 ;
        RECT 401.550 405.600 402.750 407.700 ;
        RECT 401.550 399.750 403.350 405.600 ;
        RECT 407.550 404.700 415.350 406.050 ;
        RECT 407.550 399.750 409.350 404.700 ;
        RECT 410.550 399.750 412.350 403.800 ;
        RECT 413.550 399.750 415.350 404.700 ;
        RECT 416.550 405.600 417.750 407.700 ;
        RECT 425.550 407.700 426.750 415.050 ;
        RECT 427.950 413.850 430.050 415.950 ;
        RECT 428.100 412.050 429.900 413.850 ;
        RECT 425.550 406.800 429.150 407.700 ;
        RECT 416.550 399.750 418.350 405.600 ;
        RECT 422.850 399.750 424.650 405.600 ;
        RECT 427.350 399.750 429.150 406.800 ;
        RECT 435.150 405.600 436.050 418.200 ;
        RECT 444.450 417.900 452.850 418.200 ;
        RECT 454.050 418.800 460.050 419.700 ;
        RECT 460.950 418.800 463.050 419.700 ;
        RECT 466.650 419.400 468.450 431.250 ;
        RECT 444.450 417.600 446.250 417.900 ;
        RECT 454.050 414.150 454.950 418.800 ;
        RECT 460.950 417.600 465.150 418.800 ;
        RECT 464.250 415.800 466.050 417.600 ;
        RECT 445.950 413.100 448.050 414.150 ;
        RECT 437.100 411.150 438.900 412.950 ;
        RECT 440.100 412.050 448.050 413.100 ;
        RECT 451.950 412.050 454.950 414.150 ;
        RECT 440.100 411.300 441.900 412.050 ;
        RECT 438.000 410.400 438.900 411.150 ;
        RECT 443.100 410.400 444.900 411.000 ;
        RECT 438.000 409.200 444.900 410.400 ;
        RECT 443.850 408.000 444.900 409.200 ;
        RECT 454.050 408.000 454.950 412.050 ;
        RECT 463.950 411.750 466.050 412.050 ;
        RECT 462.150 409.950 466.050 411.750 ;
        RECT 467.250 409.950 468.450 419.400 ;
        RECT 443.850 407.100 454.950 408.000 ;
        RECT 463.950 407.850 468.450 409.950 ;
        RECT 443.850 406.200 444.900 407.100 ;
        RECT 454.050 406.800 454.950 407.100 ;
        RECT 435.150 399.750 436.950 405.600 ;
        RECT 439.950 403.500 442.050 405.600 ;
        RECT 443.550 404.400 445.350 406.200 ;
        RECT 446.850 405.450 448.650 406.200 ;
        RECT 446.850 404.400 451.800 405.450 ;
        RECT 454.050 405.000 455.850 406.800 ;
        RECT 467.250 405.600 468.450 407.850 ;
        RECT 460.950 404.700 463.050 405.600 ;
        RECT 441.000 402.600 442.050 403.500 ;
        RECT 450.750 402.600 451.800 404.400 ;
        RECT 459.300 403.500 463.050 404.700 ;
        RECT 459.300 402.600 460.350 403.500 ;
        RECT 438.150 399.750 439.950 402.600 ;
        RECT 441.000 401.700 444.750 402.600 ;
        RECT 442.950 399.750 444.750 401.700 ;
        RECT 447.450 399.750 449.250 402.600 ;
        RECT 450.750 399.750 452.550 402.600 ;
        RECT 454.650 399.750 456.450 402.600 ;
        RECT 458.850 399.750 460.650 402.600 ;
        RECT 463.350 399.750 465.150 402.600 ;
        RECT 466.650 399.750 468.450 405.600 ;
        RECT 471.150 419.400 472.950 431.250 ;
        RECT 474.150 425.400 475.950 431.250 ;
        RECT 479.250 425.400 481.050 431.250 ;
        RECT 484.050 425.400 485.850 431.250 ;
        RECT 479.550 424.500 480.750 425.400 ;
        RECT 487.050 424.500 488.850 431.250 ;
        RECT 490.950 425.400 492.750 431.250 ;
        RECT 495.150 425.400 496.950 431.250 ;
        RECT 499.650 428.400 501.450 431.250 ;
        RECT 475.950 422.400 480.750 424.500 ;
        RECT 483.150 422.700 490.050 424.500 ;
        RECT 495.150 423.300 499.050 425.400 ;
        RECT 479.550 421.500 480.750 422.400 ;
        RECT 492.450 421.800 494.250 422.400 ;
        RECT 479.550 420.300 487.050 421.500 ;
        RECT 485.250 419.700 487.050 420.300 ;
        RECT 487.950 420.900 494.250 421.800 ;
        RECT 471.150 418.800 482.250 419.400 ;
        RECT 487.950 418.800 488.850 420.900 ;
        RECT 492.450 420.600 494.250 420.900 ;
        RECT 495.150 420.600 497.850 422.400 ;
        RECT 495.150 419.700 496.050 420.600 ;
        RECT 471.150 418.200 488.850 418.800 ;
        RECT 471.150 405.600 472.050 418.200 ;
        RECT 480.450 417.900 488.850 418.200 ;
        RECT 490.050 418.800 496.050 419.700 ;
        RECT 496.950 418.800 499.050 419.700 ;
        RECT 502.650 419.400 504.450 431.250 ;
        RECT 508.650 425.400 510.450 431.250 ;
        RECT 511.650 425.400 513.450 431.250 ;
        RECT 480.450 417.600 482.250 417.900 ;
        RECT 490.050 414.150 490.950 418.800 ;
        RECT 496.950 417.600 501.150 418.800 ;
        RECT 500.250 415.800 502.050 417.600 ;
        RECT 481.950 413.100 484.050 414.150 ;
        RECT 473.100 411.150 474.900 412.950 ;
        RECT 476.100 412.050 484.050 413.100 ;
        RECT 487.950 412.050 490.950 414.150 ;
        RECT 476.100 411.300 477.900 412.050 ;
        RECT 474.000 410.400 474.900 411.150 ;
        RECT 479.100 410.400 480.900 411.000 ;
        RECT 474.000 409.200 480.900 410.400 ;
        RECT 479.850 408.000 480.900 409.200 ;
        RECT 490.050 408.000 490.950 412.050 ;
        RECT 499.950 411.750 502.050 412.050 ;
        RECT 498.150 409.950 502.050 411.750 ;
        RECT 503.250 409.950 504.450 419.400 ;
        RECT 509.400 412.950 510.600 425.400 ;
        RECT 519.450 419.400 521.250 431.250 ;
        RECT 523.650 419.400 525.450 431.250 ;
        RECT 529.650 419.400 531.450 431.250 ;
        RECT 532.650 419.400 534.450 431.250 ;
        RECT 537.150 419.400 538.950 431.250 ;
        RECT 540.150 425.400 541.950 431.250 ;
        RECT 545.250 425.400 547.050 431.250 ;
        RECT 550.050 425.400 551.850 431.250 ;
        RECT 545.550 424.500 546.750 425.400 ;
        RECT 553.050 424.500 554.850 431.250 ;
        RECT 556.950 425.400 558.750 431.250 ;
        RECT 561.150 425.400 562.950 431.250 ;
        RECT 565.650 428.400 567.450 431.250 ;
        RECT 541.950 422.400 546.750 424.500 ;
        RECT 549.150 422.700 556.050 424.500 ;
        RECT 561.150 423.300 565.050 425.400 ;
        RECT 545.550 421.500 546.750 422.400 ;
        RECT 558.450 421.800 560.250 422.400 ;
        RECT 545.550 420.300 553.050 421.500 ;
        RECT 551.250 419.700 553.050 420.300 ;
        RECT 553.950 420.900 560.250 421.800 ;
        RECT 519.450 418.350 522.000 419.400 ;
        RECT 518.100 414.150 519.900 415.950 ;
        RECT 508.950 410.850 511.050 412.950 ;
        RECT 512.100 411.150 513.900 412.950 ;
        RECT 517.950 412.050 520.050 414.150 ;
        RECT 520.950 411.150 522.000 418.350 ;
        RECT 524.100 414.150 525.900 415.950 ;
        RECT 530.400 414.150 531.600 419.400 ;
        RECT 537.150 418.800 548.250 419.400 ;
        RECT 553.950 418.800 554.850 420.900 ;
        RECT 558.450 420.600 560.250 420.900 ;
        RECT 561.150 420.600 563.850 422.400 ;
        RECT 561.150 419.700 562.050 420.600 ;
        RECT 537.150 418.200 554.850 418.800 ;
        RECT 523.950 412.050 526.050 414.150 ;
        RECT 529.950 412.050 532.050 414.150 ;
        RECT 479.850 407.100 490.950 408.000 ;
        RECT 499.950 407.850 504.450 409.950 ;
        RECT 479.850 406.200 480.900 407.100 ;
        RECT 490.050 406.800 490.950 407.100 ;
        RECT 471.150 399.750 472.950 405.600 ;
        RECT 475.950 403.500 478.050 405.600 ;
        RECT 479.550 404.400 481.350 406.200 ;
        RECT 482.850 405.450 484.650 406.200 ;
        RECT 482.850 404.400 487.800 405.450 ;
        RECT 490.050 405.000 491.850 406.800 ;
        RECT 503.250 405.600 504.450 407.850 ;
        RECT 496.950 404.700 499.050 405.600 ;
        RECT 477.000 402.600 478.050 403.500 ;
        RECT 486.750 402.600 487.800 404.400 ;
        RECT 495.300 403.500 499.050 404.700 ;
        RECT 495.300 402.600 496.350 403.500 ;
        RECT 474.150 399.750 475.950 402.600 ;
        RECT 477.000 401.700 480.750 402.600 ;
        RECT 478.950 399.750 480.750 401.700 ;
        RECT 483.450 399.750 485.250 402.600 ;
        RECT 486.750 399.750 488.550 402.600 ;
        RECT 490.650 399.750 492.450 402.600 ;
        RECT 494.850 399.750 496.650 402.600 ;
        RECT 499.350 399.750 501.150 402.600 ;
        RECT 502.650 399.750 504.450 405.600 ;
        RECT 509.400 402.600 510.600 410.850 ;
        RECT 511.950 409.050 514.050 411.150 ;
        RECT 520.950 409.050 523.050 411.150 ;
        RECT 520.950 402.600 522.000 409.050 ;
        RECT 530.400 405.600 531.600 412.050 ;
        RECT 532.950 410.850 535.050 412.950 ;
        RECT 533.100 409.050 534.900 410.850 ;
        RECT 537.150 405.600 538.050 418.200 ;
        RECT 546.450 417.900 554.850 418.200 ;
        RECT 556.050 418.800 562.050 419.700 ;
        RECT 562.950 418.800 565.050 419.700 ;
        RECT 568.650 419.400 570.450 431.250 ;
        RECT 574.650 430.500 582.450 431.250 ;
        RECT 574.650 419.400 576.450 430.500 ;
        RECT 577.650 419.400 579.450 429.600 ;
        RECT 580.650 420.600 582.450 430.500 ;
        RECT 583.650 421.500 585.450 431.250 ;
        RECT 586.650 420.600 588.450 431.250 ;
        RECT 580.650 419.700 588.450 420.600 ;
        RECT 594.450 419.400 596.250 431.250 ;
        RECT 598.650 419.400 600.450 431.250 ;
        RECT 603.300 419.400 605.100 431.250 ;
        RECT 607.500 419.400 609.300 431.250 ;
        RECT 610.800 425.400 612.600 431.250 ;
        RECT 620.400 425.400 622.200 431.250 ;
        RECT 623.700 419.400 625.500 431.250 ;
        RECT 627.900 419.400 629.700 431.250 ;
        RECT 632.550 419.400 634.350 431.250 ;
        RECT 636.750 419.400 638.550 431.250 ;
        RECT 546.450 417.600 548.250 417.900 ;
        RECT 556.050 414.150 556.950 418.800 ;
        RECT 562.950 417.600 567.150 418.800 ;
        RECT 566.250 415.800 568.050 417.600 ;
        RECT 547.950 413.100 550.050 414.150 ;
        RECT 539.100 411.150 540.900 412.950 ;
        RECT 542.100 412.050 550.050 413.100 ;
        RECT 553.950 412.050 556.950 414.150 ;
        RECT 542.100 411.300 543.900 412.050 ;
        RECT 540.000 410.400 540.900 411.150 ;
        RECT 545.100 410.400 546.900 411.000 ;
        RECT 540.000 409.200 546.900 410.400 ;
        RECT 545.850 408.000 546.900 409.200 ;
        RECT 556.050 408.000 556.950 412.050 ;
        RECT 565.950 411.750 568.050 412.050 ;
        RECT 564.150 409.950 568.050 411.750 ;
        RECT 569.250 409.950 570.450 419.400 ;
        RECT 577.800 418.500 579.600 419.400 ;
        RECT 577.800 417.600 581.850 418.500 ;
        RECT 594.450 418.350 597.000 419.400 ;
        RECT 575.100 414.150 576.900 415.950 ;
        RECT 580.950 414.150 581.850 417.600 ;
        RECT 586.950 414.150 588.750 415.950 ;
        RECT 593.100 414.150 594.900 415.950 ;
        RECT 574.950 412.050 577.050 414.150 ;
        RECT 577.950 410.850 580.050 412.950 ;
        RECT 580.950 412.050 583.050 414.150 ;
        RECT 545.850 407.100 556.950 408.000 ;
        RECT 565.950 407.850 570.450 409.950 ;
        RECT 578.250 409.050 580.050 410.850 ;
        RECT 545.850 406.200 546.900 407.100 ;
        RECT 556.050 406.800 556.950 407.100 ;
        RECT 508.650 399.750 510.450 402.600 ;
        RECT 511.650 399.750 513.450 402.600 ;
        RECT 517.650 399.750 519.450 402.600 ;
        RECT 520.650 399.750 522.450 402.600 ;
        RECT 523.650 399.750 525.450 402.600 ;
        RECT 529.650 399.750 531.450 405.600 ;
        RECT 532.650 399.750 534.450 405.600 ;
        RECT 537.150 399.750 538.950 405.600 ;
        RECT 541.950 403.500 544.050 405.600 ;
        RECT 545.550 404.400 547.350 406.200 ;
        RECT 548.850 405.450 550.650 406.200 ;
        RECT 548.850 404.400 553.800 405.450 ;
        RECT 556.050 405.000 557.850 406.800 ;
        RECT 569.250 405.600 570.450 407.850 ;
        RECT 582.000 405.600 583.050 412.050 ;
        RECT 583.950 410.850 586.050 412.950 ;
        RECT 586.950 412.050 589.050 414.150 ;
        RECT 592.950 412.050 595.050 414.150 ;
        RECT 595.950 411.150 597.000 418.350 ;
        RECT 599.100 414.150 600.900 415.950 ;
        RECT 602.100 414.150 603.900 415.950 ;
        RECT 607.950 414.150 609.150 419.400 ;
        RECT 610.950 417.150 612.750 418.950 ;
        RECT 620.250 417.150 622.050 418.950 ;
        RECT 610.950 415.050 613.050 417.150 ;
        RECT 619.950 415.050 622.050 417.150 ;
        RECT 623.850 414.150 625.050 419.400 ;
        RECT 636.000 418.350 638.550 419.400 ;
        RECT 645.150 419.400 646.950 431.250 ;
        RECT 648.150 425.400 649.950 431.250 ;
        RECT 653.250 425.400 655.050 431.250 ;
        RECT 658.050 425.400 659.850 431.250 ;
        RECT 653.550 424.500 654.750 425.400 ;
        RECT 661.050 424.500 662.850 431.250 ;
        RECT 664.950 425.400 666.750 431.250 ;
        RECT 669.150 425.400 670.950 431.250 ;
        RECT 673.650 428.400 675.450 431.250 ;
        RECT 649.950 422.400 654.750 424.500 ;
        RECT 657.150 422.700 664.050 424.500 ;
        RECT 669.150 423.300 673.050 425.400 ;
        RECT 653.550 421.500 654.750 422.400 ;
        RECT 666.450 421.800 668.250 422.400 ;
        RECT 653.550 420.300 661.050 421.500 ;
        RECT 659.250 419.700 661.050 420.300 ;
        RECT 661.950 420.900 668.250 421.800 ;
        RECT 645.150 418.800 656.250 419.400 ;
        RECT 661.950 418.800 662.850 420.900 ;
        RECT 666.450 420.600 668.250 420.900 ;
        RECT 669.150 420.600 671.850 422.400 ;
        RECT 669.150 419.700 670.050 420.600 ;
        RECT 629.100 414.150 630.900 415.950 ;
        RECT 632.100 414.150 633.900 415.950 ;
        RECT 598.950 412.050 601.050 414.150 ;
        RECT 601.950 412.050 604.050 414.150 ;
        RECT 583.950 409.050 585.750 410.850 ;
        RECT 595.950 409.050 598.050 411.150 ;
        RECT 604.950 410.850 607.050 412.950 ;
        RECT 607.950 412.050 610.050 414.150 ;
        RECT 605.100 409.050 606.900 410.850 ;
        RECT 562.950 404.700 565.050 405.600 ;
        RECT 543.000 402.600 544.050 403.500 ;
        RECT 552.750 402.600 553.800 404.400 ;
        RECT 561.300 403.500 565.050 404.700 ;
        RECT 561.300 402.600 562.350 403.500 ;
        RECT 540.150 399.750 541.950 402.600 ;
        RECT 543.000 401.700 546.750 402.600 ;
        RECT 544.950 399.750 546.750 401.700 ;
        RECT 549.450 399.750 551.250 402.600 ;
        RECT 552.750 399.750 554.550 402.600 ;
        RECT 556.650 399.750 558.450 402.600 ;
        RECT 560.850 399.750 562.650 402.600 ;
        RECT 565.350 399.750 567.150 402.600 ;
        RECT 568.650 399.750 570.450 405.600 ;
        RECT 577.800 399.750 579.600 405.600 ;
        RECT 582.000 399.750 583.800 405.600 ;
        RECT 586.200 399.750 588.000 405.600 ;
        RECT 595.950 402.600 597.000 409.050 ;
        RECT 608.850 408.750 610.050 412.050 ;
        RECT 622.950 412.050 625.050 414.150 ;
        RECT 622.950 408.750 624.150 412.050 ;
        RECT 625.950 410.850 628.050 412.950 ;
        RECT 628.950 412.050 631.050 414.150 ;
        RECT 631.950 412.050 634.050 414.150 ;
        RECT 636.000 411.150 637.050 418.350 ;
        RECT 645.150 418.200 662.850 418.800 ;
        RECT 638.100 414.150 639.900 415.950 ;
        RECT 637.950 412.050 640.050 414.150 ;
        RECT 626.100 409.050 627.900 410.850 ;
        RECT 634.950 409.050 637.050 411.150 ;
        RECT 609.000 407.700 612.750 408.750 ;
        RECT 602.550 404.700 610.350 406.050 ;
        RECT 592.650 399.750 594.450 402.600 ;
        RECT 595.650 399.750 597.450 402.600 ;
        RECT 598.650 399.750 600.450 402.600 ;
        RECT 602.550 399.750 604.350 404.700 ;
        RECT 605.550 399.750 607.350 403.800 ;
        RECT 608.550 399.750 610.350 404.700 ;
        RECT 611.550 405.600 612.750 407.700 ;
        RECT 620.250 407.700 624.000 408.750 ;
        RECT 620.250 405.600 621.450 407.700 ;
        RECT 611.550 399.750 613.350 405.600 ;
        RECT 619.650 399.750 621.450 405.600 ;
        RECT 622.650 404.700 630.450 406.050 ;
        RECT 622.650 399.750 624.450 404.700 ;
        RECT 625.650 399.750 627.450 403.800 ;
        RECT 628.650 399.750 630.450 404.700 ;
        RECT 636.000 402.600 637.050 409.050 ;
        RECT 645.150 405.600 646.050 418.200 ;
        RECT 654.450 417.900 662.850 418.200 ;
        RECT 664.050 418.800 670.050 419.700 ;
        RECT 670.950 418.800 673.050 419.700 ;
        RECT 676.650 419.400 678.450 431.250 ;
        RECT 681.300 419.400 683.100 431.250 ;
        RECT 685.500 419.400 687.300 431.250 ;
        RECT 688.800 425.400 690.600 431.250 ;
        RECT 695.550 425.400 697.350 431.250 ;
        RECT 698.550 425.400 700.350 431.250 ;
        RECT 701.550 425.400 703.350 431.250 ;
        RECT 654.450 417.600 656.250 417.900 ;
        RECT 664.050 414.150 664.950 418.800 ;
        RECT 670.950 417.600 675.150 418.800 ;
        RECT 674.250 415.800 676.050 417.600 ;
        RECT 655.950 413.100 658.050 414.150 ;
        RECT 647.100 411.150 648.900 412.950 ;
        RECT 650.100 412.050 658.050 413.100 ;
        RECT 661.950 412.050 664.950 414.150 ;
        RECT 650.100 411.300 651.900 412.050 ;
        RECT 648.000 410.400 648.900 411.150 ;
        RECT 653.100 410.400 654.900 411.000 ;
        RECT 648.000 409.200 654.900 410.400 ;
        RECT 653.850 408.000 654.900 409.200 ;
        RECT 664.050 408.000 664.950 412.050 ;
        RECT 673.950 411.750 676.050 412.050 ;
        RECT 672.150 409.950 676.050 411.750 ;
        RECT 677.250 409.950 678.450 419.400 ;
        RECT 680.100 414.150 681.900 415.950 ;
        RECT 685.950 414.150 687.150 419.400 ;
        RECT 688.950 417.150 690.750 418.950 ;
        RECT 698.550 417.150 699.750 425.400 ;
        RECT 688.950 415.050 691.050 417.150 ;
        RECT 679.950 412.050 682.050 414.150 ;
        RECT 682.950 410.850 685.050 412.950 ;
        RECT 685.950 412.050 688.050 414.150 ;
        RECT 694.950 413.850 697.050 415.950 ;
        RECT 697.950 415.050 700.050 417.150 ;
        RECT 695.100 412.050 696.900 413.850 ;
        RECT 653.850 407.100 664.950 408.000 ;
        RECT 673.950 407.850 678.450 409.950 ;
        RECT 683.100 409.050 684.900 410.850 ;
        RECT 686.850 408.750 688.050 412.050 ;
        RECT 653.850 406.200 654.900 407.100 ;
        RECT 664.050 406.800 664.950 407.100 ;
        RECT 632.550 399.750 634.350 402.600 ;
        RECT 635.550 399.750 637.350 402.600 ;
        RECT 638.550 399.750 640.350 402.600 ;
        RECT 645.150 399.750 646.950 405.600 ;
        RECT 649.950 403.500 652.050 405.600 ;
        RECT 653.550 404.400 655.350 406.200 ;
        RECT 656.850 405.450 658.650 406.200 ;
        RECT 656.850 404.400 661.800 405.450 ;
        RECT 664.050 405.000 665.850 406.800 ;
        RECT 677.250 405.600 678.450 407.850 ;
        RECT 687.000 407.700 690.750 408.750 ;
        RECT 670.950 404.700 673.050 405.600 ;
        RECT 651.000 402.600 652.050 403.500 ;
        RECT 660.750 402.600 661.800 404.400 ;
        RECT 669.300 403.500 673.050 404.700 ;
        RECT 669.300 402.600 670.350 403.500 ;
        RECT 648.150 399.750 649.950 402.600 ;
        RECT 651.000 401.700 654.750 402.600 ;
        RECT 652.950 399.750 654.750 401.700 ;
        RECT 657.450 399.750 659.250 402.600 ;
        RECT 660.750 399.750 662.550 402.600 ;
        RECT 664.650 399.750 666.450 402.600 ;
        RECT 668.850 399.750 670.650 402.600 ;
        RECT 673.350 399.750 675.150 402.600 ;
        RECT 676.650 399.750 678.450 405.600 ;
        RECT 680.550 404.700 688.350 406.050 ;
        RECT 680.550 399.750 682.350 404.700 ;
        RECT 683.550 399.750 685.350 403.800 ;
        RECT 686.550 399.750 688.350 404.700 ;
        RECT 689.550 405.600 690.750 407.700 ;
        RECT 698.550 407.700 699.750 415.050 ;
        RECT 700.950 413.850 703.050 415.950 ;
        RECT 701.100 412.050 702.900 413.850 ;
        RECT 698.550 406.800 702.150 407.700 ;
        RECT 689.550 399.750 691.350 405.600 ;
        RECT 695.850 399.750 697.650 405.600 ;
        RECT 700.350 399.750 702.150 406.800 ;
        RECT 2.700 386.400 4.500 395.250 ;
        RECT 8.100 387.000 9.900 395.250 ;
        RECT 18.000 389.400 19.800 395.250 ;
        RECT 22.200 391.050 24.000 395.250 ;
        RECT 25.500 392.400 27.300 395.250 ;
        RECT 34.650 392.400 36.450 395.250 ;
        RECT 37.650 392.400 39.450 395.250 ;
        RECT 22.200 389.400 27.900 391.050 ;
        RECT 8.100 385.350 12.600 387.000 ;
        RECT 11.400 381.150 12.600 385.350 ;
        RECT 17.100 384.150 18.900 385.950 ;
        RECT 16.950 382.050 19.050 384.150 ;
        RECT 19.950 383.850 22.050 385.950 ;
        RECT 23.100 384.150 24.900 385.950 ;
        RECT 20.100 382.050 21.900 383.850 ;
        RECT 22.950 382.050 25.050 384.150 ;
        RECT 26.700 382.950 27.900 389.400 ;
        RECT 35.400 384.150 36.600 392.400 ;
        RECT 45.150 390.900 46.950 395.250 ;
        RECT 43.650 389.400 46.950 390.900 ;
        RECT 48.150 389.400 49.950 395.250 ;
        RECT 1.950 377.850 4.050 379.950 ;
        RECT 7.950 377.850 10.050 379.950 ;
        RECT 10.950 379.050 13.050 381.150 ;
        RECT 25.950 380.850 28.050 382.950 ;
        RECT 34.950 382.050 37.050 384.150 ;
        RECT 37.950 383.850 40.050 385.950 ;
        RECT 38.100 382.050 39.900 383.850 ;
        RECT 43.650 382.950 44.850 389.400 ;
        RECT 46.950 387.900 48.750 388.500 ;
        RECT 52.650 387.900 54.450 395.250 ;
        RECT 59.700 392.400 61.500 395.250 ;
        RECT 63.000 391.050 64.800 395.250 ;
        RECT 46.950 386.700 54.450 387.900 ;
        RECT 59.100 389.400 64.800 391.050 ;
        RECT 67.200 389.400 69.000 395.250 ;
        RECT 73.950 390.450 76.050 391.050 ;
        RECT 71.550 389.550 76.050 390.450 ;
        RECT 2.100 376.050 3.900 377.850 ;
        RECT 4.950 374.850 7.050 376.950 ;
        RECT 8.250 376.050 10.050 377.850 ;
        RECT 5.100 373.050 6.900 374.850 ;
        RECT 11.700 370.800 12.750 379.050 ;
        RECT 26.700 375.600 27.900 380.850 ;
        RECT 5.700 369.900 12.750 370.800 ;
        RECT 5.700 369.600 7.350 369.900 ;
        RECT 2.550 363.750 4.350 369.600 ;
        RECT 5.550 363.750 7.350 369.600 ;
        RECT 11.550 369.600 12.750 369.900 ;
        RECT 17.550 374.700 25.350 375.600 ;
        RECT 8.550 363.750 10.350 369.000 ;
        RECT 11.550 363.750 13.350 369.600 ;
        RECT 17.550 363.750 19.350 374.700 ;
        RECT 20.550 363.750 22.350 373.800 ;
        RECT 23.550 363.750 25.350 374.700 ;
        RECT 26.550 363.750 28.350 375.600 ;
        RECT 35.400 369.600 36.600 382.050 ;
        RECT 43.650 380.850 46.050 382.950 ;
        RECT 47.100 381.150 48.900 382.950 ;
        RECT 43.650 375.600 44.850 380.850 ;
        RECT 46.950 379.050 49.050 381.150 ;
        RECT 34.650 363.750 36.450 369.600 ;
        RECT 37.650 363.750 39.450 369.600 ;
        RECT 43.050 363.750 44.850 375.600 ;
        RECT 46.050 363.750 47.850 375.600 ;
        RECT 50.100 369.600 51.300 386.700 ;
        RECT 59.100 382.950 60.300 389.400 ;
        RECT 62.100 384.150 63.900 385.950 ;
        RECT 52.950 380.850 55.050 382.950 ;
        RECT 58.950 380.850 61.050 382.950 ;
        RECT 61.950 382.050 64.050 384.150 ;
        RECT 64.950 383.850 67.050 385.950 ;
        RECT 68.100 384.150 69.900 385.950 ;
        RECT 65.100 382.050 66.900 383.850 ;
        RECT 67.950 382.050 70.050 384.150 ;
        RECT 53.100 379.050 54.900 380.850 ;
        RECT 59.100 375.600 60.300 380.850 ;
        RECT 67.950 378.450 70.050 379.050 ;
        RECT 71.550 378.450 72.450 389.550 ;
        RECT 73.950 388.950 76.050 389.550 ;
        RECT 77.100 387.000 78.900 395.250 ;
        RECT 74.400 385.350 78.900 387.000 ;
        RECT 82.500 386.400 84.300 395.250 ;
        RECT 88.650 389.400 90.450 395.250 ;
        RECT 89.250 387.300 90.450 389.400 ;
        RECT 91.650 390.300 93.450 395.250 ;
        RECT 94.650 391.200 96.450 395.250 ;
        RECT 97.650 390.300 99.450 395.250 ;
        RECT 91.650 388.950 99.450 390.300 ;
        RECT 103.650 389.400 105.450 395.250 ;
        RECT 106.650 389.400 108.450 395.250 ;
        RECT 89.250 386.250 93.000 387.300 ;
        RECT 74.400 381.150 75.600 385.350 ;
        RECT 79.950 384.450 82.050 385.050 ;
        RECT 88.950 384.450 91.050 385.050 ;
        RECT 79.950 383.550 91.050 384.450 ;
        RECT 79.950 382.950 82.050 383.550 ;
        RECT 88.950 382.950 91.050 383.550 ;
        RECT 91.950 382.950 93.150 386.250 ;
        RECT 95.100 384.150 96.900 385.950 ;
        RECT 73.950 379.050 76.050 381.150 ;
        RECT 91.950 380.850 94.050 382.950 ;
        RECT 94.950 382.050 97.050 384.150 ;
        RECT 104.400 382.950 105.600 389.400 ;
        RECT 113.850 388.200 115.650 395.250 ;
        RECT 118.350 389.400 120.150 395.250 ;
        RECT 113.850 387.300 117.450 388.200 ;
        RECT 107.100 384.150 108.900 385.950 ;
        RECT 97.950 380.850 100.050 382.950 ;
        RECT 103.950 380.850 106.050 382.950 ;
        RECT 106.950 382.050 109.050 384.150 ;
        RECT 113.100 381.150 114.900 382.950 ;
        RECT 67.950 377.550 72.450 378.450 ;
        RECT 67.950 376.950 70.050 377.550 ;
        RECT 49.650 363.750 51.450 369.600 ;
        RECT 52.650 363.750 54.450 369.600 ;
        RECT 58.650 363.750 60.450 375.600 ;
        RECT 61.650 374.700 69.450 375.600 ;
        RECT 61.650 363.750 63.450 374.700 ;
        RECT 64.650 363.750 66.450 373.800 ;
        RECT 67.650 363.750 69.450 374.700 ;
        RECT 74.250 370.800 75.300 379.050 ;
        RECT 76.950 377.850 79.050 379.950 ;
        RECT 82.950 377.850 85.050 379.950 ;
        RECT 88.950 377.850 91.050 379.950 ;
        RECT 76.950 376.050 78.750 377.850 ;
        RECT 79.950 374.850 82.050 376.950 ;
        RECT 83.100 376.050 84.900 377.850 ;
        RECT 89.250 376.050 91.050 377.850 ;
        RECT 92.850 375.600 94.050 380.850 ;
        RECT 98.100 379.050 99.900 380.850 ;
        RECT 104.400 375.600 105.600 380.850 ;
        RECT 112.950 379.050 115.050 381.150 ;
        RECT 116.250 379.950 117.450 387.300 ;
        RECT 118.950 387.450 121.050 388.050 ;
        RECT 118.950 386.550 123.450 387.450 ;
        RECT 128.100 387.000 129.900 395.250 ;
        RECT 118.950 385.950 121.050 386.550 ;
        RECT 119.100 381.150 120.900 382.950 ;
        RECT 115.950 377.850 118.050 379.950 ;
        RECT 118.950 379.050 121.050 381.150 ;
        RECT 80.100 373.050 81.900 374.850 ;
        RECT 74.250 369.900 81.300 370.800 ;
        RECT 74.250 369.600 75.450 369.900 ;
        RECT 73.650 363.750 75.450 369.600 ;
        RECT 79.650 369.600 81.300 369.900 ;
        RECT 76.650 363.750 78.450 369.000 ;
        RECT 79.650 363.750 81.450 369.600 ;
        RECT 82.650 363.750 84.450 369.600 ;
        RECT 89.400 363.750 91.200 369.600 ;
        RECT 92.700 363.750 94.500 375.600 ;
        RECT 96.900 363.750 98.700 375.600 ;
        RECT 103.650 363.750 105.450 375.600 ;
        RECT 106.650 363.750 108.450 375.600 ;
        RECT 116.250 369.600 117.450 377.850 ;
        RECT 118.950 375.450 121.050 376.050 ;
        RECT 122.550 375.450 123.450 386.550 ;
        RECT 125.400 385.350 129.900 387.000 ;
        RECT 133.500 386.400 135.300 395.250 ;
        RECT 139.650 389.400 141.450 395.250 ;
        RECT 140.250 387.300 141.450 389.400 ;
        RECT 142.650 390.300 144.450 395.250 ;
        RECT 145.650 391.200 147.450 395.250 ;
        RECT 148.650 390.300 150.450 395.250 ;
        RECT 142.650 388.950 150.450 390.300 ;
        RECT 152.850 389.400 154.650 395.250 ;
        RECT 157.350 388.200 159.150 395.250 ;
        RECT 155.550 387.300 159.150 388.200 ;
        RECT 140.250 386.250 144.000 387.300 ;
        RECT 125.400 381.150 126.600 385.350 ;
        RECT 142.950 382.950 144.150 386.250 ;
        RECT 146.100 384.150 147.900 385.950 ;
        RECT 124.950 379.050 127.050 381.150 ;
        RECT 142.950 380.850 145.050 382.950 ;
        RECT 145.950 382.050 148.050 384.150 ;
        RECT 148.950 380.850 151.050 382.950 ;
        RECT 152.100 381.150 153.900 382.950 ;
        RECT 118.950 374.550 123.450 375.450 ;
        RECT 118.950 373.950 121.050 374.550 ;
        RECT 125.250 370.800 126.300 379.050 ;
        RECT 127.950 377.850 130.050 379.950 ;
        RECT 133.950 377.850 136.050 379.950 ;
        RECT 139.950 377.850 142.050 379.950 ;
        RECT 127.950 376.050 129.750 377.850 ;
        RECT 130.950 374.850 133.050 376.950 ;
        RECT 134.100 376.050 135.900 377.850 ;
        RECT 140.250 376.050 142.050 377.850 ;
        RECT 143.850 375.600 145.050 380.850 ;
        RECT 149.100 379.050 150.900 380.850 ;
        RECT 151.950 379.050 154.050 381.150 ;
        RECT 155.550 379.950 156.750 387.300 ;
        RECT 170.100 387.000 171.900 395.250 ;
        RECT 167.400 385.350 171.900 387.000 ;
        RECT 175.500 386.400 177.300 395.250 ;
        RECT 181.650 392.400 183.450 395.250 ;
        RECT 184.650 392.400 186.450 395.250 ;
        RECT 158.100 381.150 159.900 382.950 ;
        RECT 167.400 381.150 168.600 385.350 ;
        RECT 182.400 384.150 183.600 392.400 ;
        RECT 190.650 389.400 192.450 395.250 ;
        RECT 191.250 387.300 192.450 389.400 ;
        RECT 193.650 390.300 195.450 395.250 ;
        RECT 196.650 391.200 198.450 395.250 ;
        RECT 199.650 390.300 201.450 395.250 ;
        RECT 193.650 388.950 201.450 390.300 ;
        RECT 203.850 389.400 205.650 395.250 ;
        RECT 208.350 388.200 210.150 395.250 ;
        RECT 215.550 389.400 217.350 395.250 ;
        RECT 218.550 389.400 220.350 395.250 ;
        RECT 206.550 387.300 210.150 388.200 ;
        RECT 191.250 386.250 195.000 387.300 ;
        RECT 181.950 382.050 184.050 384.150 ;
        RECT 184.950 383.850 187.050 385.950 ;
        RECT 185.100 382.050 186.900 383.850 ;
        RECT 193.950 382.950 195.150 386.250 ;
        RECT 197.100 384.150 198.900 385.950 ;
        RECT 154.950 377.850 157.050 379.950 ;
        RECT 157.950 379.050 160.050 381.150 ;
        RECT 166.950 379.050 169.050 381.150 ;
        RECT 131.100 373.050 132.900 374.850 ;
        RECT 125.250 369.900 132.300 370.800 ;
        RECT 125.250 369.600 126.450 369.900 ;
        RECT 112.650 363.750 114.450 369.600 ;
        RECT 115.650 363.750 117.450 369.600 ;
        RECT 118.650 363.750 120.450 369.600 ;
        RECT 124.650 363.750 126.450 369.600 ;
        RECT 130.650 369.600 132.300 369.900 ;
        RECT 127.650 363.750 129.450 369.000 ;
        RECT 130.650 363.750 132.450 369.600 ;
        RECT 133.650 363.750 135.450 369.600 ;
        RECT 140.400 363.750 142.200 369.600 ;
        RECT 143.700 363.750 145.500 375.600 ;
        RECT 147.900 363.750 149.700 375.600 ;
        RECT 155.550 369.600 156.750 377.850 ;
        RECT 167.250 370.800 168.300 379.050 ;
        RECT 169.950 377.850 172.050 379.950 ;
        RECT 175.950 377.850 178.050 379.950 ;
        RECT 169.950 376.050 171.750 377.850 ;
        RECT 172.950 374.850 175.050 376.950 ;
        RECT 176.100 376.050 177.900 377.850 ;
        RECT 173.100 373.050 174.900 374.850 ;
        RECT 167.250 369.900 174.300 370.800 ;
        RECT 167.250 369.600 168.450 369.900 ;
        RECT 152.550 363.750 154.350 369.600 ;
        RECT 155.550 363.750 157.350 369.600 ;
        RECT 158.550 363.750 160.350 369.600 ;
        RECT 166.650 363.750 168.450 369.600 ;
        RECT 172.650 369.600 174.300 369.900 ;
        RECT 182.400 369.600 183.600 382.050 ;
        RECT 193.950 380.850 196.050 382.950 ;
        RECT 196.950 382.050 199.050 384.150 ;
        RECT 199.950 380.850 202.050 382.950 ;
        RECT 203.100 381.150 204.900 382.950 ;
        RECT 190.950 377.850 193.050 379.950 ;
        RECT 191.250 376.050 193.050 377.850 ;
        RECT 194.850 375.600 196.050 380.850 ;
        RECT 200.100 379.050 201.900 380.850 ;
        RECT 202.950 379.050 205.050 381.150 ;
        RECT 206.550 379.950 207.750 387.300 ;
        RECT 215.100 384.150 216.900 385.950 ;
        RECT 209.100 381.150 210.900 382.950 ;
        RECT 214.950 382.050 217.050 384.150 ;
        RECT 218.400 382.950 219.600 389.400 ;
        RECT 227.850 388.200 229.650 395.250 ;
        RECT 232.350 389.400 234.150 395.250 ;
        RECT 237.150 389.400 238.950 395.250 ;
        RECT 240.150 392.400 241.950 395.250 ;
        RECT 244.950 393.300 246.750 395.250 ;
        RECT 243.000 392.400 246.750 393.300 ;
        RECT 249.450 392.400 251.250 395.250 ;
        RECT 252.750 392.400 254.550 395.250 ;
        RECT 256.650 392.400 258.450 395.250 ;
        RECT 260.850 392.400 262.650 395.250 ;
        RECT 265.350 392.400 267.150 395.250 ;
        RECT 243.000 391.500 244.050 392.400 ;
        RECT 241.950 389.400 244.050 391.500 ;
        RECT 252.750 390.600 253.800 392.400 ;
        RECT 227.850 387.300 231.450 388.200 ;
        RECT 205.950 377.850 208.050 379.950 ;
        RECT 208.950 379.050 211.050 381.150 ;
        RECT 217.950 380.850 220.050 382.950 ;
        RECT 227.100 381.150 228.900 382.950 ;
        RECT 169.650 363.750 171.450 369.000 ;
        RECT 172.650 363.750 174.450 369.600 ;
        RECT 175.650 363.750 177.450 369.600 ;
        RECT 181.650 363.750 183.450 369.600 ;
        RECT 184.650 363.750 186.450 369.600 ;
        RECT 191.400 363.750 193.200 369.600 ;
        RECT 194.700 363.750 196.500 375.600 ;
        RECT 198.900 363.750 200.700 375.600 ;
        RECT 206.550 369.600 207.750 377.850 ;
        RECT 218.400 375.600 219.600 380.850 ;
        RECT 226.950 379.050 229.050 381.150 ;
        RECT 230.250 379.950 231.450 387.300 ;
        RECT 233.100 381.150 234.900 382.950 ;
        RECT 229.950 377.850 232.050 379.950 ;
        RECT 232.950 379.050 235.050 381.150 ;
        RECT 203.550 363.750 205.350 369.600 ;
        RECT 206.550 363.750 208.350 369.600 ;
        RECT 209.550 363.750 211.350 369.600 ;
        RECT 215.550 363.750 217.350 375.600 ;
        RECT 218.550 363.750 220.350 375.600 ;
        RECT 230.250 369.600 231.450 377.850 ;
        RECT 237.150 376.800 238.050 389.400 ;
        RECT 245.550 388.800 247.350 390.600 ;
        RECT 248.850 389.550 253.800 390.600 ;
        RECT 261.300 391.500 262.350 392.400 ;
        RECT 261.300 390.300 265.050 391.500 ;
        RECT 248.850 388.800 250.650 389.550 ;
        RECT 245.850 387.900 246.900 388.800 ;
        RECT 256.050 388.200 257.850 390.000 ;
        RECT 262.950 389.400 265.050 390.300 ;
        RECT 268.650 389.400 270.450 395.250 ;
        RECT 272.850 389.400 274.650 395.250 ;
        RECT 256.050 387.900 256.950 388.200 ;
        RECT 245.850 387.000 256.950 387.900 ;
        RECT 269.250 387.150 270.450 389.400 ;
        RECT 277.350 388.200 279.150 395.250 ;
        RECT 284.850 389.400 286.650 395.250 ;
        RECT 289.350 388.200 291.150 395.250 ;
        RECT 245.850 385.800 246.900 387.000 ;
        RECT 240.000 384.600 246.900 385.800 ;
        RECT 240.000 383.850 240.900 384.600 ;
        RECT 245.100 384.000 246.900 384.600 ;
        RECT 239.100 382.050 240.900 383.850 ;
        RECT 242.100 382.950 243.900 383.700 ;
        RECT 256.050 382.950 256.950 387.000 ;
        RECT 265.950 385.050 270.450 387.150 ;
        RECT 264.150 383.250 268.050 385.050 ;
        RECT 265.950 382.950 268.050 383.250 ;
        RECT 242.100 381.900 250.050 382.950 ;
        RECT 247.950 380.850 250.050 381.900 ;
        RECT 253.950 380.850 256.950 382.950 ;
        RECT 246.450 377.100 248.250 377.400 ;
        RECT 246.450 376.800 254.850 377.100 ;
        RECT 237.150 376.200 254.850 376.800 ;
        RECT 237.150 375.600 248.250 376.200 ;
        RECT 226.650 363.750 228.450 369.600 ;
        RECT 229.650 363.750 231.450 369.600 ;
        RECT 232.650 363.750 234.450 369.600 ;
        RECT 237.150 363.750 238.950 375.600 ;
        RECT 251.250 374.700 253.050 375.300 ;
        RECT 245.550 373.500 253.050 374.700 ;
        RECT 253.950 374.100 254.850 376.200 ;
        RECT 256.050 376.200 256.950 380.850 ;
        RECT 266.250 377.400 268.050 379.200 ;
        RECT 262.950 376.200 267.150 377.400 ;
        RECT 256.050 375.300 262.050 376.200 ;
        RECT 262.950 375.300 265.050 376.200 ;
        RECT 269.250 375.600 270.450 385.050 ;
        RECT 275.550 387.300 279.150 388.200 ;
        RECT 287.550 387.300 291.150 388.200 ;
        RECT 272.100 381.150 273.900 382.950 ;
        RECT 271.950 379.050 274.050 381.150 ;
        RECT 275.550 379.950 276.750 387.300 ;
        RECT 278.100 381.150 279.900 382.950 ;
        RECT 284.100 381.150 285.900 382.950 ;
        RECT 274.950 377.850 277.050 379.950 ;
        RECT 277.950 379.050 280.050 381.150 ;
        RECT 283.950 379.050 286.050 381.150 ;
        RECT 287.550 379.950 288.750 387.300 ;
        RECT 296.700 386.400 298.500 395.250 ;
        RECT 302.100 387.000 303.900 395.250 ;
        RECT 311.550 392.400 313.350 395.250 ;
        RECT 314.550 392.400 316.350 395.250 ;
        RECT 317.550 392.400 319.350 395.250 ;
        RECT 325.650 392.400 327.450 395.250 ;
        RECT 328.650 392.400 330.450 395.250 ;
        RECT 334.650 392.400 336.450 395.250 ;
        RECT 337.650 392.400 339.450 395.250 ;
        RECT 340.650 392.400 342.450 395.250 ;
        RECT 346.650 392.400 348.450 395.250 ;
        RECT 349.650 392.400 351.450 395.250 ;
        RECT 302.100 385.350 306.600 387.000 ;
        RECT 315.000 385.950 316.050 392.400 ;
        RECT 290.100 381.150 291.900 382.950 ;
        RECT 305.400 381.150 306.600 385.350 ;
        RECT 313.950 383.850 316.050 385.950 ;
        RECT 326.400 384.150 327.600 392.400 ;
        RECT 337.950 385.950 339.000 392.400 ;
        RECT 286.950 377.850 289.050 379.950 ;
        RECT 289.950 379.050 292.050 381.150 ;
        RECT 295.950 377.850 298.050 379.950 ;
        RECT 301.950 377.850 304.050 379.950 ;
        RECT 304.950 379.050 307.050 381.150 ;
        RECT 310.950 380.850 313.050 382.950 ;
        RECT 311.100 379.050 312.900 380.850 ;
        RECT 261.150 374.400 262.050 375.300 ;
        RECT 258.450 374.100 260.250 374.400 ;
        RECT 245.550 372.600 246.750 373.500 ;
        RECT 253.950 373.200 260.250 374.100 ;
        RECT 258.450 372.600 260.250 373.200 ;
        RECT 261.150 372.600 263.850 374.400 ;
        RECT 241.950 370.500 246.750 372.600 ;
        RECT 249.150 370.500 256.050 372.300 ;
        RECT 245.550 369.600 246.750 370.500 ;
        RECT 240.150 363.750 241.950 369.600 ;
        RECT 245.250 363.750 247.050 369.600 ;
        RECT 250.050 363.750 251.850 369.600 ;
        RECT 253.050 363.750 254.850 370.500 ;
        RECT 261.150 369.600 265.050 371.700 ;
        RECT 256.950 363.750 258.750 369.600 ;
        RECT 261.150 363.750 262.950 369.600 ;
        RECT 265.650 363.750 267.450 366.600 ;
        RECT 268.650 363.750 270.450 375.600 ;
        RECT 275.550 369.600 276.750 377.850 ;
        RECT 287.550 369.600 288.750 377.850 ;
        RECT 296.100 376.050 297.900 377.850 ;
        RECT 298.950 374.850 301.050 376.950 ;
        RECT 302.250 376.050 304.050 377.850 ;
        RECT 299.100 373.050 300.900 374.850 ;
        RECT 305.700 370.800 306.750 379.050 ;
        RECT 315.000 376.650 316.050 383.850 ;
        RECT 316.950 380.850 319.050 382.950 ;
        RECT 325.950 382.050 328.050 384.150 ;
        RECT 328.950 383.850 331.050 385.950 ;
        RECT 337.950 383.850 340.050 385.950 ;
        RECT 347.400 384.150 348.600 392.400 ;
        RECT 355.650 389.400 357.450 395.250 ;
        RECT 356.250 387.300 357.450 389.400 ;
        RECT 358.650 390.300 360.450 395.250 ;
        RECT 361.650 391.200 363.450 395.250 ;
        RECT 364.650 390.300 366.450 395.250 ;
        RECT 368.550 392.400 370.350 395.250 ;
        RECT 371.550 392.400 373.350 395.250 ;
        RECT 374.550 392.400 376.350 395.250 ;
        RECT 358.650 388.950 366.450 390.300 ;
        RECT 356.250 386.250 360.000 387.300 ;
        RECT 329.100 382.050 330.900 383.850 ;
        RECT 317.100 379.050 318.900 380.850 ;
        RECT 315.000 375.600 317.550 376.650 ;
        RECT 299.700 369.900 306.750 370.800 ;
        RECT 299.700 369.600 301.350 369.900 ;
        RECT 272.550 363.750 274.350 369.600 ;
        RECT 275.550 363.750 277.350 369.600 ;
        RECT 278.550 363.750 280.350 369.600 ;
        RECT 284.550 363.750 286.350 369.600 ;
        RECT 287.550 363.750 289.350 369.600 ;
        RECT 290.550 363.750 292.350 369.600 ;
        RECT 296.550 363.750 298.350 369.600 ;
        RECT 299.550 363.750 301.350 369.600 ;
        RECT 305.550 369.600 306.750 369.900 ;
        RECT 302.550 363.750 304.350 369.000 ;
        RECT 305.550 363.750 307.350 369.600 ;
        RECT 311.550 363.750 313.350 375.600 ;
        RECT 315.750 363.750 317.550 375.600 ;
        RECT 326.400 369.600 327.600 382.050 ;
        RECT 334.950 380.850 337.050 382.950 ;
        RECT 335.100 379.050 336.900 380.850 ;
        RECT 337.950 376.650 339.000 383.850 ;
        RECT 340.950 380.850 343.050 382.950 ;
        RECT 346.950 382.050 349.050 384.150 ;
        RECT 349.950 383.850 352.050 385.950 ;
        RECT 350.100 382.050 351.900 383.850 ;
        RECT 358.950 382.950 360.150 386.250 ;
        RECT 372.000 385.950 373.050 392.400 ;
        RECT 380.550 387.900 382.350 395.250 ;
        RECT 385.050 389.400 386.850 395.250 ;
        RECT 388.050 390.900 389.850 395.250 ;
        RECT 388.050 389.400 391.350 390.900 ;
        RECT 386.250 387.900 388.050 388.500 ;
        RECT 380.550 386.700 388.050 387.900 ;
        RECT 362.100 384.150 363.900 385.950 ;
        RECT 341.100 379.050 342.900 380.850 ;
        RECT 336.450 375.600 339.000 376.650 ;
        RECT 325.650 363.750 327.450 369.600 ;
        RECT 328.650 363.750 330.450 369.600 ;
        RECT 336.450 363.750 338.250 375.600 ;
        RECT 340.650 363.750 342.450 375.600 ;
        RECT 347.400 369.600 348.600 382.050 ;
        RECT 358.950 380.850 361.050 382.950 ;
        RECT 361.950 382.050 364.050 384.150 ;
        RECT 370.950 383.850 373.050 385.950 ;
        RECT 364.950 380.850 367.050 382.950 ;
        RECT 367.950 380.850 370.050 382.950 ;
        RECT 355.950 377.850 358.050 379.950 ;
        RECT 356.250 376.050 358.050 377.850 ;
        RECT 359.850 375.600 361.050 380.850 ;
        RECT 365.100 379.050 366.900 380.850 ;
        RECT 368.100 379.050 369.900 380.850 ;
        RECT 372.000 376.650 373.050 383.850 ;
        RECT 373.950 380.850 376.050 382.950 ;
        RECT 379.950 380.850 382.050 382.950 ;
        RECT 374.100 379.050 375.900 380.850 ;
        RECT 380.100 379.050 381.900 380.850 ;
        RECT 372.000 375.600 374.550 376.650 ;
        RECT 346.650 363.750 348.450 369.600 ;
        RECT 349.650 363.750 351.450 369.600 ;
        RECT 356.400 363.750 358.200 369.600 ;
        RECT 359.700 363.750 361.500 375.600 ;
        RECT 363.900 363.750 365.700 375.600 ;
        RECT 368.550 363.750 370.350 375.600 ;
        RECT 372.750 363.750 374.550 375.600 ;
        RECT 383.700 369.600 384.900 386.700 ;
        RECT 390.150 382.950 391.350 389.400 ;
        RECT 395.550 390.300 397.350 395.250 ;
        RECT 398.550 391.200 400.350 395.250 ;
        RECT 401.550 390.300 403.350 395.250 ;
        RECT 395.550 388.950 403.350 390.300 ;
        RECT 404.550 389.400 406.350 395.250 ;
        RECT 404.550 387.300 405.750 389.400 ;
        RECT 413.850 388.200 415.650 395.250 ;
        RECT 418.350 389.400 420.150 395.250 ;
        RECT 422.550 392.400 424.350 395.250 ;
        RECT 425.550 392.400 427.350 395.250 ;
        RECT 428.550 392.400 430.350 395.250 ;
        RECT 426.450 388.200 427.350 392.400 ;
        RECT 431.550 389.400 433.350 395.250 ;
        RECT 437.850 389.400 439.650 395.250 ;
        RECT 413.850 387.300 417.450 388.200 ;
        RECT 426.450 387.300 429.750 388.200 ;
        RECT 402.000 386.250 405.750 387.300 ;
        RECT 398.100 384.150 399.900 385.950 ;
        RECT 386.100 381.150 387.900 382.950 ;
        RECT 385.950 379.050 388.050 381.150 ;
        RECT 388.950 380.850 391.350 382.950 ;
        RECT 394.950 380.850 397.050 382.950 ;
        RECT 397.950 382.050 400.050 384.150 ;
        RECT 401.850 382.950 403.050 386.250 ;
        RECT 400.950 380.850 403.050 382.950 ;
        RECT 413.100 381.150 414.900 382.950 ;
        RECT 390.150 375.600 391.350 380.850 ;
        RECT 395.100 379.050 396.900 380.850 ;
        RECT 400.950 375.600 402.150 380.850 ;
        RECT 403.950 377.850 406.050 379.950 ;
        RECT 412.950 379.050 415.050 381.150 ;
        RECT 416.250 379.950 417.450 387.300 ;
        RECT 427.950 386.400 429.750 387.300 ;
        RECT 421.950 383.850 424.050 385.950 ;
        RECT 419.100 381.150 420.900 382.950 ;
        RECT 422.100 382.050 423.900 383.850 ;
        RECT 415.950 377.850 418.050 379.950 ;
        RECT 418.950 379.050 421.050 381.150 ;
        RECT 424.950 380.850 427.050 382.950 ;
        RECT 425.100 379.050 426.900 380.850 ;
        RECT 428.700 378.150 429.600 386.400 ;
        RECT 432.000 384.150 433.050 389.400 ;
        RECT 442.350 388.200 444.150 395.250 ;
        RECT 449.550 392.400 451.350 395.250 ;
        RECT 430.950 382.050 433.050 384.150 ;
        RECT 440.550 387.300 444.150 388.200 ;
        RECT 450.150 388.500 451.350 392.400 ;
        RECT 452.850 389.400 454.650 395.250 ;
        RECT 455.850 389.400 457.650 395.250 ;
        RECT 461.550 390.300 463.350 395.250 ;
        RECT 464.550 391.200 466.350 395.250 ;
        RECT 467.550 390.300 469.350 395.250 ;
        RECT 450.150 387.600 455.250 388.500 ;
        RECT 427.950 378.000 429.750 378.150 ;
        RECT 403.950 376.050 405.750 377.850 ;
        RECT 380.550 363.750 382.350 369.600 ;
        RECT 383.550 363.750 385.350 369.600 ;
        RECT 387.150 363.750 388.950 375.600 ;
        RECT 390.150 363.750 391.950 375.600 ;
        RECT 396.300 363.750 398.100 375.600 ;
        RECT 400.500 363.750 402.300 375.600 ;
        RECT 416.250 369.600 417.450 377.850 ;
        RECT 422.550 376.800 429.750 378.000 ;
        RECT 422.550 375.600 423.750 376.800 ;
        RECT 427.950 376.350 429.750 376.800 ;
        RECT 403.800 363.750 405.600 369.600 ;
        RECT 412.650 363.750 414.450 369.600 ;
        RECT 415.650 363.750 417.450 369.600 ;
        RECT 418.650 363.750 420.450 369.600 ;
        RECT 422.550 363.750 424.350 375.600 ;
        RECT 431.100 375.450 432.450 382.050 ;
        RECT 437.100 381.150 438.900 382.950 ;
        RECT 436.950 379.050 439.050 381.150 ;
        RECT 440.550 379.950 441.750 387.300 ;
        RECT 453.000 386.700 455.250 387.600 ;
        RECT 443.100 381.150 444.900 382.950 ;
        RECT 439.950 377.850 442.050 379.950 ;
        RECT 442.950 379.050 445.050 381.150 ;
        RECT 448.950 380.850 451.050 382.950 ;
        RECT 449.100 379.050 450.900 380.850 ;
        RECT 453.000 378.300 454.050 386.700 ;
        RECT 456.150 382.950 457.350 389.400 ;
        RECT 461.550 388.950 469.350 390.300 ;
        RECT 470.550 389.400 472.350 395.250 ;
        RECT 478.350 389.400 480.150 395.250 ;
        RECT 481.350 389.400 483.150 395.250 ;
        RECT 484.650 392.400 486.450 395.250 ;
        RECT 470.550 387.300 471.750 389.400 ;
        RECT 468.000 386.250 471.750 387.300 ;
        RECT 464.100 384.150 465.900 385.950 ;
        RECT 454.950 380.850 457.350 382.950 ;
        RECT 460.950 380.850 463.050 382.950 ;
        RECT 463.950 382.050 466.050 384.150 ;
        RECT 467.850 382.950 469.050 386.250 ;
        RECT 466.950 380.850 469.050 382.950 ;
        RECT 478.650 382.950 479.850 389.400 ;
        RECT 484.650 388.500 485.850 392.400 ;
        RECT 480.750 387.600 485.850 388.500 ;
        RECT 491.850 388.200 493.650 395.250 ;
        RECT 496.350 389.400 498.150 395.250 ;
        RECT 501.000 389.400 502.800 395.250 ;
        RECT 505.200 389.400 507.000 395.250 ;
        RECT 509.400 389.400 511.200 395.250 ;
        RECT 518.550 392.400 520.350 395.250 ;
        RECT 480.750 386.700 483.000 387.600 ;
        RECT 491.850 387.300 495.450 388.200 ;
        RECT 478.650 380.850 481.050 382.950 ;
        RECT 427.050 363.750 428.850 375.450 ;
        RECT 430.050 374.100 432.450 375.450 ;
        RECT 430.050 363.750 431.850 374.100 ;
        RECT 440.550 369.600 441.750 377.850 ;
        RECT 453.000 377.400 455.250 378.300 ;
        RECT 449.550 376.500 455.250 377.400 ;
        RECT 449.550 369.600 450.750 376.500 ;
        RECT 456.150 375.600 457.350 380.850 ;
        RECT 461.100 379.050 462.900 380.850 ;
        RECT 466.950 375.600 468.150 380.850 ;
        RECT 469.950 377.850 472.050 379.950 ;
        RECT 469.950 376.050 471.750 377.850 ;
        RECT 478.650 375.600 479.850 380.850 ;
        RECT 481.950 378.300 483.000 386.700 ;
        RECT 484.950 380.850 487.050 382.950 ;
        RECT 491.100 381.150 492.900 382.950 ;
        RECT 485.100 379.050 486.900 380.850 ;
        RECT 490.950 379.050 493.050 381.150 ;
        RECT 494.250 379.950 495.450 387.300 ;
        RECT 503.250 384.150 505.050 385.950 ;
        RECT 497.100 381.150 498.900 382.950 ;
        RECT 480.750 377.400 483.000 378.300 ;
        RECT 493.950 377.850 496.050 379.950 ;
        RECT 496.950 379.050 499.050 381.150 ;
        RECT 499.950 380.850 502.050 382.950 ;
        RECT 502.950 382.050 505.050 384.150 ;
        RECT 505.950 382.950 507.000 389.400 ;
        RECT 519.150 388.500 520.350 392.400 ;
        RECT 521.850 389.400 523.650 395.250 ;
        RECT 524.850 389.400 526.650 395.250 ;
        RECT 532.350 389.400 534.150 395.250 ;
        RECT 535.350 389.400 537.150 395.250 ;
        RECT 538.650 392.400 540.450 395.250 ;
        RECT 519.150 387.600 524.250 388.500 ;
        RECT 522.000 386.700 524.250 387.600 ;
        RECT 508.950 384.150 510.750 385.950 ;
        RECT 505.950 380.850 508.050 382.950 ;
        RECT 508.950 382.050 511.050 384.150 ;
        RECT 511.950 380.850 514.050 382.950 ;
        RECT 517.950 380.850 520.050 382.950 ;
        RECT 500.250 379.050 502.050 380.850 ;
        RECT 480.750 376.500 486.450 377.400 ;
        RECT 437.550 363.750 439.350 369.600 ;
        RECT 440.550 363.750 442.350 369.600 ;
        RECT 443.550 363.750 445.350 369.600 ;
        RECT 449.550 363.750 451.350 369.600 ;
        RECT 452.850 363.750 454.650 375.600 ;
        RECT 455.850 363.750 457.650 375.600 ;
        RECT 462.300 363.750 464.100 375.600 ;
        RECT 466.500 363.750 468.300 375.600 ;
        RECT 469.800 363.750 471.600 369.600 ;
        RECT 478.350 363.750 480.150 375.600 ;
        RECT 481.350 363.750 483.150 375.600 ;
        RECT 485.250 369.600 486.450 376.500 ;
        RECT 494.250 369.600 495.450 377.850 ;
        RECT 507.150 377.400 508.050 380.850 ;
        RECT 512.100 379.050 513.900 380.850 ;
        RECT 518.100 379.050 519.900 380.850 ;
        RECT 522.000 378.300 523.050 386.700 ;
        RECT 525.150 382.950 526.350 389.400 ;
        RECT 523.950 380.850 526.350 382.950 ;
        RECT 522.000 377.400 524.250 378.300 ;
        RECT 507.150 376.500 511.200 377.400 ;
        RECT 509.400 375.600 511.200 376.500 ;
        RECT 518.550 376.500 524.250 377.400 ;
        RECT 500.550 374.400 508.350 375.300 ;
        RECT 484.650 363.750 486.450 369.600 ;
        RECT 490.650 363.750 492.450 369.600 ;
        RECT 493.650 363.750 495.450 369.600 ;
        RECT 496.650 363.750 498.450 369.600 ;
        RECT 500.550 363.750 502.350 374.400 ;
        RECT 503.550 363.750 505.350 373.500 ;
        RECT 506.550 364.500 508.350 374.400 ;
        RECT 509.550 365.400 511.350 375.600 ;
        RECT 512.550 364.500 514.350 375.600 ;
        RECT 506.550 363.750 514.350 364.500 ;
        RECT 518.550 369.600 519.750 376.500 ;
        RECT 525.150 375.600 526.350 380.850 ;
        RECT 532.650 382.950 533.850 389.400 ;
        RECT 538.650 388.500 539.850 392.400 ;
        RECT 534.750 387.600 539.850 388.500 ;
        RECT 543.150 389.400 544.950 395.250 ;
        RECT 546.150 392.400 547.950 395.250 ;
        RECT 550.950 393.300 552.750 395.250 ;
        RECT 549.000 392.400 552.750 393.300 ;
        RECT 555.450 392.400 557.250 395.250 ;
        RECT 558.750 392.400 560.550 395.250 ;
        RECT 562.650 392.400 564.450 395.250 ;
        RECT 566.850 392.400 568.650 395.250 ;
        RECT 571.350 392.400 573.150 395.250 ;
        RECT 549.000 391.500 550.050 392.400 ;
        RECT 547.950 389.400 550.050 391.500 ;
        RECT 558.750 390.600 559.800 392.400 ;
        RECT 534.750 386.700 537.000 387.600 ;
        RECT 532.650 380.850 535.050 382.950 ;
        RECT 532.650 375.600 533.850 380.850 ;
        RECT 535.950 378.300 537.000 386.700 ;
        RECT 538.950 380.850 541.050 382.950 ;
        RECT 539.100 379.050 540.900 380.850 ;
        RECT 534.750 377.400 537.000 378.300 ;
        RECT 534.750 376.500 540.450 377.400 ;
        RECT 518.550 363.750 520.350 369.600 ;
        RECT 521.850 363.750 523.650 375.600 ;
        RECT 524.850 363.750 526.650 375.600 ;
        RECT 532.350 363.750 534.150 375.600 ;
        RECT 535.350 363.750 537.150 375.600 ;
        RECT 539.250 369.600 540.450 376.500 ;
        RECT 538.650 363.750 540.450 369.600 ;
        RECT 543.150 376.800 544.050 389.400 ;
        RECT 551.550 388.800 553.350 390.600 ;
        RECT 554.850 389.550 559.800 390.600 ;
        RECT 567.300 391.500 568.350 392.400 ;
        RECT 567.300 390.300 571.050 391.500 ;
        RECT 554.850 388.800 556.650 389.550 ;
        RECT 551.850 387.900 552.900 388.800 ;
        RECT 562.050 388.200 563.850 390.000 ;
        RECT 568.950 389.400 571.050 390.300 ;
        RECT 574.650 389.400 576.450 395.250 ;
        RECT 581.700 392.400 583.500 395.250 ;
        RECT 585.000 391.050 586.800 395.250 ;
        RECT 562.050 387.900 562.950 388.200 ;
        RECT 551.850 387.000 562.950 387.900 ;
        RECT 575.250 387.150 576.450 389.400 ;
        RECT 551.850 385.800 552.900 387.000 ;
        RECT 546.000 384.600 552.900 385.800 ;
        RECT 546.000 383.850 546.900 384.600 ;
        RECT 551.100 384.000 552.900 384.600 ;
        RECT 545.100 382.050 546.900 383.850 ;
        RECT 548.100 382.950 549.900 383.700 ;
        RECT 562.050 382.950 562.950 387.000 ;
        RECT 571.950 385.050 576.450 387.150 ;
        RECT 570.150 383.250 574.050 385.050 ;
        RECT 571.950 382.950 574.050 383.250 ;
        RECT 548.100 381.900 556.050 382.950 ;
        RECT 553.950 380.850 556.050 381.900 ;
        RECT 559.950 380.850 562.950 382.950 ;
        RECT 552.450 377.100 554.250 377.400 ;
        RECT 552.450 376.800 560.850 377.100 ;
        RECT 543.150 376.200 560.850 376.800 ;
        RECT 543.150 375.600 554.250 376.200 ;
        RECT 543.150 363.750 544.950 375.600 ;
        RECT 557.250 374.700 559.050 375.300 ;
        RECT 551.550 373.500 559.050 374.700 ;
        RECT 559.950 374.100 560.850 376.200 ;
        RECT 562.050 376.200 562.950 380.850 ;
        RECT 572.250 377.400 574.050 379.200 ;
        RECT 568.950 376.200 573.150 377.400 ;
        RECT 562.050 375.300 568.050 376.200 ;
        RECT 568.950 375.300 571.050 376.200 ;
        RECT 575.250 375.600 576.450 385.050 ;
        RECT 581.100 389.400 586.800 391.050 ;
        RECT 589.200 389.400 591.000 395.250 ;
        RECT 593.550 392.400 595.350 395.250 ;
        RECT 596.550 392.400 598.350 395.250 ;
        RECT 599.550 392.400 601.350 395.250 ;
        RECT 581.100 382.950 582.300 389.400 ;
        RECT 597.000 385.950 598.050 392.400 ;
        RECT 605.550 389.400 607.350 395.250 ;
        RECT 608.550 389.400 610.350 395.250 ;
        RECT 611.550 389.400 613.350 395.250 ;
        RECT 608.400 388.500 610.200 389.400 ;
        RECT 614.550 388.500 616.350 395.250 ;
        RECT 617.550 389.400 619.350 395.250 ;
        RECT 620.550 389.400 622.350 395.250 ;
        RECT 623.550 389.400 625.350 395.250 ;
        RECT 626.550 389.400 628.350 395.250 ;
        RECT 629.550 389.400 631.350 395.250 ;
        RECT 636.150 389.400 637.950 395.250 ;
        RECT 639.150 392.400 640.950 395.250 ;
        RECT 643.950 393.300 645.750 395.250 ;
        RECT 642.000 392.400 645.750 393.300 ;
        RECT 648.450 392.400 650.250 395.250 ;
        RECT 651.750 392.400 653.550 395.250 ;
        RECT 655.650 392.400 657.450 395.250 ;
        RECT 659.850 392.400 661.650 395.250 ;
        RECT 664.350 392.400 666.150 395.250 ;
        RECT 642.000 391.500 643.050 392.400 ;
        RECT 640.950 389.400 643.050 391.500 ;
        RECT 651.750 390.600 652.800 392.400 ;
        RECT 620.400 388.500 622.200 389.400 ;
        RECT 626.400 388.500 628.200 389.400 ;
        RECT 608.400 387.300 612.450 388.500 ;
        RECT 614.550 387.300 618.300 388.500 ;
        RECT 620.400 387.300 624.300 388.500 ;
        RECT 626.400 388.350 629.100 388.500 ;
        RECT 626.400 387.300 629.250 388.350 ;
        RECT 611.250 386.400 612.450 387.300 ;
        RECT 617.100 386.400 618.300 387.300 ;
        RECT 623.100 386.400 624.300 387.300 ;
        RECT 584.100 384.150 585.900 385.950 ;
        RECT 580.950 380.850 583.050 382.950 ;
        RECT 583.950 382.050 586.050 384.150 ;
        RECT 586.950 383.850 589.050 385.950 ;
        RECT 590.100 384.150 591.900 385.950 ;
        RECT 587.100 382.050 588.900 383.850 ;
        RECT 589.950 382.050 592.050 384.150 ;
        RECT 595.950 383.850 598.050 385.950 ;
        RECT 608.100 384.150 609.900 385.950 ;
        RECT 611.250 384.600 615.300 386.400 ;
        RECT 617.100 384.600 621.300 386.400 ;
        RECT 623.100 384.600 627.300 386.400 ;
        RECT 592.950 380.850 595.050 382.950 ;
        RECT 581.100 375.600 582.300 380.850 ;
        RECT 593.100 379.050 594.900 380.850 ;
        RECT 597.000 376.650 598.050 383.850 ;
        RECT 598.950 380.850 601.050 382.950 ;
        RECT 607.950 382.050 610.050 384.150 ;
        RECT 599.100 379.050 600.900 380.850 ;
        RECT 611.250 377.700 612.450 384.600 ;
        RECT 617.100 377.700 618.300 384.600 ;
        RECT 623.100 377.700 624.300 384.600 ;
        RECT 628.200 384.150 629.250 387.300 ;
        RECT 628.200 382.050 631.050 384.150 ;
        RECT 628.200 377.700 629.250 382.050 ;
        RECT 597.000 375.600 599.550 376.650 ;
        RECT 608.550 376.500 612.450 377.700 ;
        RECT 614.550 376.500 618.300 377.700 ;
        RECT 620.550 376.500 624.300 377.700 ;
        RECT 626.550 376.500 629.250 377.700 ;
        RECT 636.150 376.800 637.050 389.400 ;
        RECT 644.550 388.800 646.350 390.600 ;
        RECT 647.850 389.550 652.800 390.600 ;
        RECT 660.300 391.500 661.350 392.400 ;
        RECT 660.300 390.300 664.050 391.500 ;
        RECT 647.850 388.800 649.650 389.550 ;
        RECT 644.850 387.900 645.900 388.800 ;
        RECT 655.050 388.200 656.850 390.000 ;
        RECT 661.950 389.400 664.050 390.300 ;
        RECT 667.650 389.400 669.450 395.250 ;
        RECT 655.050 387.900 655.950 388.200 ;
        RECT 644.850 387.000 655.950 387.900 ;
        RECT 668.250 387.150 669.450 389.400 ;
        RECT 671.550 390.300 673.350 395.250 ;
        RECT 674.550 391.200 676.350 395.250 ;
        RECT 677.550 390.300 679.350 395.250 ;
        RECT 671.550 388.950 679.350 390.300 ;
        RECT 680.550 389.400 682.350 395.250 ;
        RECT 686.850 389.400 688.650 395.250 ;
        RECT 680.550 387.300 681.750 389.400 ;
        RECT 691.350 388.200 693.150 395.250 ;
        RECT 698.850 389.400 700.650 395.250 ;
        RECT 703.350 388.200 705.150 395.250 ;
        RECT 644.850 385.800 645.900 387.000 ;
        RECT 639.000 384.600 645.900 385.800 ;
        RECT 639.000 383.850 639.900 384.600 ;
        RECT 644.100 384.000 645.900 384.600 ;
        RECT 638.100 382.050 639.900 383.850 ;
        RECT 641.100 382.950 642.900 383.700 ;
        RECT 655.050 382.950 655.950 387.000 ;
        RECT 664.950 385.050 669.450 387.150 ;
        RECT 678.000 386.250 681.750 387.300 ;
        RECT 689.550 387.300 693.150 388.200 ;
        RECT 701.550 387.300 705.150 388.200 ;
        RECT 663.150 383.250 667.050 385.050 ;
        RECT 664.950 382.950 667.050 383.250 ;
        RECT 641.100 381.900 649.050 382.950 ;
        RECT 646.950 380.850 649.050 381.900 ;
        RECT 652.950 380.850 655.950 382.950 ;
        RECT 645.450 377.100 647.250 377.400 ;
        RECT 645.450 376.800 653.850 377.100 ;
        RECT 567.150 374.400 568.050 375.300 ;
        RECT 564.450 374.100 566.250 374.400 ;
        RECT 551.550 372.600 552.750 373.500 ;
        RECT 559.950 373.200 566.250 374.100 ;
        RECT 564.450 372.600 566.250 373.200 ;
        RECT 567.150 372.600 569.850 374.400 ;
        RECT 547.950 370.500 552.750 372.600 ;
        RECT 555.150 370.500 562.050 372.300 ;
        RECT 551.550 369.600 552.750 370.500 ;
        RECT 546.150 363.750 547.950 369.600 ;
        RECT 551.250 363.750 553.050 369.600 ;
        RECT 556.050 363.750 557.850 369.600 ;
        RECT 559.050 363.750 560.850 370.500 ;
        RECT 567.150 369.600 571.050 371.700 ;
        RECT 562.950 363.750 564.750 369.600 ;
        RECT 567.150 363.750 568.950 369.600 ;
        RECT 571.650 363.750 573.450 366.600 ;
        RECT 574.650 363.750 576.450 375.600 ;
        RECT 580.650 363.750 582.450 375.600 ;
        RECT 583.650 374.700 591.450 375.600 ;
        RECT 583.650 363.750 585.450 374.700 ;
        RECT 586.650 363.750 588.450 373.800 ;
        RECT 589.650 363.750 591.450 374.700 ;
        RECT 593.550 363.750 595.350 375.600 ;
        RECT 597.750 363.750 599.550 375.600 ;
        RECT 605.550 363.750 607.350 375.600 ;
        RECT 608.550 363.750 610.350 376.500 ;
        RECT 611.550 363.750 613.350 375.600 ;
        RECT 614.550 363.750 616.350 376.500 ;
        RECT 617.550 363.750 619.350 375.600 ;
        RECT 620.550 363.750 622.350 376.500 ;
        RECT 623.550 363.750 625.350 375.600 ;
        RECT 626.550 363.750 628.350 376.500 ;
        RECT 636.150 376.200 653.850 376.800 ;
        RECT 636.150 375.600 647.250 376.200 ;
        RECT 629.550 363.750 631.350 375.600 ;
        RECT 636.150 363.750 637.950 375.600 ;
        RECT 650.250 374.700 652.050 375.300 ;
        RECT 644.550 373.500 652.050 374.700 ;
        RECT 652.950 374.100 653.850 376.200 ;
        RECT 655.050 376.200 655.950 380.850 ;
        RECT 665.250 377.400 667.050 379.200 ;
        RECT 661.950 376.200 666.150 377.400 ;
        RECT 655.050 375.300 661.050 376.200 ;
        RECT 661.950 375.300 664.050 376.200 ;
        RECT 668.250 375.600 669.450 385.050 ;
        RECT 674.100 384.150 675.900 385.950 ;
        RECT 670.950 380.850 673.050 382.950 ;
        RECT 673.950 382.050 676.050 384.150 ;
        RECT 677.850 382.950 679.050 386.250 ;
        RECT 676.950 380.850 679.050 382.950 ;
        RECT 686.100 381.150 687.900 382.950 ;
        RECT 671.100 379.050 672.900 380.850 ;
        RECT 676.950 375.600 678.150 380.850 ;
        RECT 679.950 377.850 682.050 379.950 ;
        RECT 685.950 379.050 688.050 381.150 ;
        RECT 689.550 379.950 690.750 387.300 ;
        RECT 692.100 381.150 693.900 382.950 ;
        RECT 698.100 381.150 699.900 382.950 ;
        RECT 688.950 377.850 691.050 379.950 ;
        RECT 691.950 379.050 694.050 381.150 ;
        RECT 697.950 379.050 700.050 381.150 ;
        RECT 701.550 379.950 702.750 387.300 ;
        RECT 704.100 381.150 705.900 382.950 ;
        RECT 700.950 377.850 703.050 379.950 ;
        RECT 703.950 379.050 706.050 381.150 ;
        RECT 679.950 376.050 681.750 377.850 ;
        RECT 660.150 374.400 661.050 375.300 ;
        RECT 657.450 374.100 659.250 374.400 ;
        RECT 644.550 372.600 645.750 373.500 ;
        RECT 652.950 373.200 659.250 374.100 ;
        RECT 657.450 372.600 659.250 373.200 ;
        RECT 660.150 372.600 662.850 374.400 ;
        RECT 640.950 370.500 645.750 372.600 ;
        RECT 648.150 370.500 655.050 372.300 ;
        RECT 644.550 369.600 645.750 370.500 ;
        RECT 639.150 363.750 640.950 369.600 ;
        RECT 644.250 363.750 646.050 369.600 ;
        RECT 649.050 363.750 650.850 369.600 ;
        RECT 652.050 363.750 653.850 370.500 ;
        RECT 660.150 369.600 664.050 371.700 ;
        RECT 655.950 363.750 657.750 369.600 ;
        RECT 660.150 363.750 661.950 369.600 ;
        RECT 664.650 363.750 666.450 366.600 ;
        RECT 667.650 363.750 669.450 375.600 ;
        RECT 672.300 363.750 674.100 375.600 ;
        RECT 676.500 363.750 678.300 375.600 ;
        RECT 689.550 369.600 690.750 377.850 ;
        RECT 701.550 369.600 702.750 377.850 ;
        RECT 679.800 363.750 681.600 369.600 ;
        RECT 686.550 363.750 688.350 369.600 ;
        RECT 689.550 363.750 691.350 369.600 ;
        RECT 692.550 363.750 694.350 369.600 ;
        RECT 698.550 363.750 700.350 369.600 ;
        RECT 701.550 363.750 703.350 369.600 ;
        RECT 704.550 363.750 706.350 369.600 ;
        RECT 4.650 353.400 6.450 359.250 ;
        RECT 7.650 354.000 9.450 359.250 ;
        RECT 5.250 353.100 6.450 353.400 ;
        RECT 10.650 353.400 12.450 359.250 ;
        RECT 13.650 353.400 15.450 359.250 ;
        RECT 20.400 353.400 22.200 359.250 ;
        RECT 10.650 353.100 12.300 353.400 ;
        RECT 5.250 352.200 12.300 353.100 ;
        RECT 5.250 343.950 6.300 352.200 ;
        RECT 19.950 351.450 22.050 352.050 ;
        RECT 17.550 350.550 22.050 351.450 ;
        RECT 11.100 348.150 12.900 349.950 ;
        RECT 7.950 345.150 9.750 346.950 ;
        RECT 10.950 346.050 13.050 348.150 ;
        RECT 14.100 345.150 15.900 346.950 ;
        RECT 4.950 341.850 7.050 343.950 ;
        RECT 7.950 343.050 10.050 345.150 ;
        RECT 13.950 343.050 16.050 345.150 ;
        RECT 5.400 337.650 6.600 341.850 ;
        RECT 13.950 339.450 16.050 340.050 ;
        RECT 17.550 339.450 18.450 350.550 ;
        RECT 19.950 349.950 22.050 350.550 ;
        RECT 23.700 347.400 25.500 359.250 ;
        RECT 27.900 347.400 29.700 359.250 ;
        RECT 33.300 347.400 35.100 359.250 ;
        RECT 37.500 347.400 39.300 359.250 ;
        RECT 40.800 353.400 42.600 359.250 ;
        RECT 47.550 353.400 49.350 359.250 ;
        RECT 50.550 353.400 52.350 359.250 ;
        RECT 53.550 354.000 55.350 359.250 ;
        RECT 50.700 353.100 52.350 353.400 ;
        RECT 56.550 353.400 58.350 359.250 ;
        RECT 56.550 353.100 57.750 353.400 ;
        RECT 50.700 352.200 57.750 353.100 ;
        RECT 50.100 348.150 51.900 349.950 ;
        RECT 20.250 345.150 22.050 346.950 ;
        RECT 19.950 343.050 22.050 345.150 ;
        RECT 23.850 342.150 25.050 347.400 ;
        RECT 29.100 342.150 30.900 343.950 ;
        RECT 32.100 342.150 33.900 343.950 ;
        RECT 37.950 342.150 39.150 347.400 ;
        RECT 40.950 345.150 42.750 346.950 ;
        RECT 47.100 345.150 48.900 346.950 ;
        RECT 49.950 346.050 52.050 348.150 ;
        RECT 53.250 345.150 55.050 346.950 ;
        RECT 40.950 343.050 43.050 345.150 ;
        RECT 46.950 343.050 49.050 345.150 ;
        RECT 52.950 343.050 55.050 345.150 ;
        RECT 56.700 343.950 57.750 352.200 ;
        RECT 62.550 348.300 64.350 359.250 ;
        RECT 65.550 349.200 67.350 359.250 ;
        RECT 68.550 348.300 70.350 359.250 ;
        RECT 62.550 347.400 70.350 348.300 ;
        RECT 71.550 347.400 73.350 359.250 ;
        RECT 78.300 347.400 80.100 359.250 ;
        RECT 82.500 347.400 84.300 359.250 ;
        RECT 85.800 353.400 87.600 359.250 ;
        RECT 94.650 347.400 96.450 359.250 ;
        RECT 97.650 348.300 99.450 359.250 ;
        RECT 100.650 349.200 102.450 359.250 ;
        RECT 103.650 348.300 105.450 359.250 ;
        RECT 107.550 353.400 109.350 359.250 ;
        RECT 110.550 353.400 112.350 359.250 ;
        RECT 97.650 347.400 105.450 348.300 ;
        RECT 13.950 338.550 18.450 339.450 ;
        RECT 22.950 340.050 25.050 342.150 ;
        RECT 13.950 337.950 16.050 338.550 ;
        RECT 5.400 336.000 9.900 337.650 ;
        RECT 22.950 336.750 24.150 340.050 ;
        RECT 25.950 338.850 28.050 340.950 ;
        RECT 28.950 340.050 31.050 342.150 ;
        RECT 31.950 340.050 34.050 342.150 ;
        RECT 34.950 338.850 37.050 340.950 ;
        RECT 37.950 340.050 40.050 342.150 ;
        RECT 55.950 341.850 58.050 343.950 ;
        RECT 71.700 342.150 72.900 347.400 ;
        RECT 77.100 342.150 78.900 343.950 ;
        RECT 82.950 342.150 84.150 347.400 ;
        RECT 85.950 345.150 87.750 346.950 ;
        RECT 85.950 343.050 88.050 345.150 ;
        RECT 95.100 342.150 96.300 347.400 ;
        RECT 26.100 337.050 27.900 338.850 ;
        RECT 35.100 337.050 36.900 338.850 ;
        RECT 38.850 336.750 40.050 340.050 ;
        RECT 56.400 337.650 57.600 341.850 ;
        RECT 61.950 338.850 64.050 340.950 ;
        RECT 65.100 339.150 66.900 340.950 ;
        RECT 8.100 327.750 9.900 336.000 ;
        RECT 13.500 327.750 15.300 336.600 ;
        RECT 20.250 335.700 24.000 336.750 ;
        RECT 39.000 335.700 42.750 336.750 ;
        RECT 20.250 333.600 21.450 335.700 ;
        RECT 19.650 327.750 21.450 333.600 ;
        RECT 22.650 332.700 30.450 334.050 ;
        RECT 22.650 327.750 24.450 332.700 ;
        RECT 25.650 327.750 27.450 331.800 ;
        RECT 28.650 327.750 30.450 332.700 ;
        RECT 32.550 332.700 40.350 334.050 ;
        RECT 32.550 327.750 34.350 332.700 ;
        RECT 35.550 327.750 37.350 331.800 ;
        RECT 38.550 327.750 40.350 332.700 ;
        RECT 41.550 333.600 42.750 335.700 ;
        RECT 41.550 327.750 43.350 333.600 ;
        RECT 47.700 327.750 49.500 336.600 ;
        RECT 53.100 336.000 57.600 337.650 ;
        RECT 62.100 337.050 63.900 338.850 ;
        RECT 64.950 337.050 67.050 339.150 ;
        RECT 67.950 338.850 70.050 340.950 ;
        RECT 70.950 340.050 73.050 342.150 ;
        RECT 76.950 340.050 79.050 342.150 ;
        RECT 68.100 337.050 69.900 338.850 ;
        RECT 53.100 327.750 54.900 336.000 ;
        RECT 71.700 333.600 72.900 340.050 ;
        RECT 79.950 338.850 82.050 340.950 ;
        RECT 82.950 340.050 85.050 342.150 ;
        RECT 94.950 340.050 97.050 342.150 ;
        RECT 110.400 340.950 111.600 353.400 ;
        RECT 118.050 347.400 119.850 359.250 ;
        RECT 121.050 347.400 122.850 359.250 ;
        RECT 124.650 353.400 126.450 359.250 ;
        RECT 127.650 353.400 129.450 359.250 ;
        RECT 131.550 353.400 133.350 359.250 ;
        RECT 134.550 353.400 136.350 359.250 ;
        RECT 137.550 353.400 139.350 359.250 ;
        RECT 143.550 353.400 145.350 359.250 ;
        RECT 146.550 353.400 148.350 359.250 ;
        RECT 118.650 342.150 119.850 347.400 ;
        RECT 80.100 337.050 81.900 338.850 ;
        RECT 83.850 336.750 85.050 340.050 ;
        RECT 84.000 335.700 87.750 336.750 ;
        RECT 63.000 327.750 64.800 333.600 ;
        RECT 67.200 331.950 72.900 333.600 ;
        RECT 77.550 332.700 85.350 334.050 ;
        RECT 67.200 327.750 69.000 331.950 ;
        RECT 70.500 327.750 72.300 330.600 ;
        RECT 77.550 327.750 79.350 332.700 ;
        RECT 80.550 327.750 82.350 331.800 ;
        RECT 83.550 327.750 85.350 332.700 ;
        RECT 86.550 333.600 87.750 335.700 ;
        RECT 95.100 333.600 96.300 340.050 ;
        RECT 97.950 338.850 100.050 340.950 ;
        RECT 101.100 339.150 102.900 340.950 ;
        RECT 98.100 337.050 99.900 338.850 ;
        RECT 100.950 337.050 103.050 339.150 ;
        RECT 103.950 338.850 106.050 340.950 ;
        RECT 107.100 339.150 108.900 340.950 ;
        RECT 104.100 337.050 105.900 338.850 ;
        RECT 106.950 337.050 109.050 339.150 ;
        RECT 109.950 338.850 112.050 340.950 ;
        RECT 118.650 340.050 121.050 342.150 ;
        RECT 121.950 341.850 124.050 343.950 ;
        RECT 122.100 340.050 123.900 341.850 ;
        RECT 86.550 327.750 88.350 333.600 ;
        RECT 95.100 331.950 100.800 333.600 ;
        RECT 95.700 327.750 97.500 330.600 ;
        RECT 99.000 327.750 100.800 331.950 ;
        RECT 103.200 327.750 105.000 333.600 ;
        RECT 110.400 330.600 111.600 338.850 ;
        RECT 118.650 333.600 119.850 340.050 ;
        RECT 125.100 336.300 126.300 353.400 ;
        RECT 134.550 345.150 135.750 353.400 ;
        RECT 128.100 342.150 129.900 343.950 ;
        RECT 127.950 340.050 130.050 342.150 ;
        RECT 130.950 341.850 133.050 343.950 ;
        RECT 133.950 343.050 136.050 345.150 ;
        RECT 131.100 340.050 132.900 341.850 ;
        RECT 121.950 335.100 129.450 336.300 ;
        RECT 121.950 334.500 123.750 335.100 ;
        RECT 118.650 332.100 121.950 333.600 ;
        RECT 107.550 327.750 109.350 330.600 ;
        RECT 110.550 327.750 112.350 330.600 ;
        RECT 120.150 327.750 121.950 332.100 ;
        RECT 123.150 327.750 124.950 333.600 ;
        RECT 127.650 327.750 129.450 335.100 ;
        RECT 134.550 335.700 135.750 343.050 ;
        RECT 136.950 341.850 139.050 343.950 ;
        RECT 143.100 342.150 144.900 343.950 ;
        RECT 137.100 340.050 138.900 341.850 ;
        RECT 142.950 340.050 145.050 342.150 ;
        RECT 146.700 336.300 147.900 353.400 ;
        RECT 150.150 347.400 151.950 359.250 ;
        RECT 153.150 347.400 154.950 359.250 ;
        RECT 161.400 353.400 163.200 359.250 ;
        RECT 164.700 347.400 166.500 359.250 ;
        RECT 168.900 347.400 170.700 359.250 ;
        RECT 176.400 353.400 178.200 359.250 ;
        RECT 179.700 347.400 181.500 359.250 ;
        RECT 183.900 347.400 185.700 359.250 ;
        RECT 189.150 347.400 190.950 359.250 ;
        RECT 192.150 353.400 193.950 359.250 ;
        RECT 197.250 353.400 199.050 359.250 ;
        RECT 202.050 353.400 203.850 359.250 ;
        RECT 197.550 352.500 198.750 353.400 ;
        RECT 205.050 352.500 206.850 359.250 ;
        RECT 208.950 353.400 210.750 359.250 ;
        RECT 213.150 353.400 214.950 359.250 ;
        RECT 217.650 356.400 219.450 359.250 ;
        RECT 193.950 350.400 198.750 352.500 ;
        RECT 201.150 350.700 208.050 352.500 ;
        RECT 213.150 351.300 217.050 353.400 ;
        RECT 197.550 349.500 198.750 350.400 ;
        RECT 210.450 349.800 212.250 350.400 ;
        RECT 197.550 348.300 205.050 349.500 ;
        RECT 203.250 347.700 205.050 348.300 ;
        RECT 205.950 348.900 212.250 349.800 ;
        RECT 148.950 341.850 151.050 343.950 ;
        RECT 153.150 342.150 154.350 347.400 ;
        RECT 161.250 345.150 163.050 346.950 ;
        RECT 160.950 343.050 163.050 345.150 ;
        RECT 164.850 342.150 166.050 347.400 ;
        RECT 176.250 345.150 178.050 346.950 ;
        RECT 170.100 342.150 171.900 343.950 ;
        RECT 175.950 343.050 178.050 345.150 ;
        RECT 179.850 342.150 181.050 347.400 ;
        RECT 189.150 346.800 200.250 347.400 ;
        RECT 205.950 346.800 206.850 348.900 ;
        RECT 210.450 348.600 212.250 348.900 ;
        RECT 213.150 348.600 215.850 350.400 ;
        RECT 213.150 347.700 214.050 348.600 ;
        RECT 189.150 346.200 206.850 346.800 ;
        RECT 185.100 342.150 186.900 343.950 ;
        RECT 149.100 340.050 150.900 341.850 ;
        RECT 151.950 340.050 154.350 342.150 ;
        RECT 134.550 334.800 138.150 335.700 ;
        RECT 131.850 327.750 133.650 333.600 ;
        RECT 136.350 327.750 138.150 334.800 ;
        RECT 143.550 335.100 151.050 336.300 ;
        RECT 143.550 327.750 145.350 335.100 ;
        RECT 149.250 334.500 151.050 335.100 ;
        RECT 153.150 333.600 154.350 340.050 ;
        RECT 163.950 340.050 166.050 342.150 ;
        RECT 163.950 336.750 165.150 340.050 ;
        RECT 166.950 338.850 169.050 340.950 ;
        RECT 169.950 340.050 172.050 342.150 ;
        RECT 178.950 340.050 181.050 342.150 ;
        RECT 167.100 337.050 168.900 338.850 ;
        RECT 178.950 336.750 180.150 340.050 ;
        RECT 181.950 338.850 184.050 340.950 ;
        RECT 184.950 340.050 187.050 342.150 ;
        RECT 182.100 337.050 183.900 338.850 ;
        RECT 161.250 335.700 165.000 336.750 ;
        RECT 176.250 335.700 180.000 336.750 ;
        RECT 161.250 333.600 162.450 335.700 ;
        RECT 148.050 327.750 149.850 333.600 ;
        RECT 151.050 332.100 154.350 333.600 ;
        RECT 151.050 327.750 152.850 332.100 ;
        RECT 160.650 327.750 162.450 333.600 ;
        RECT 163.650 332.700 171.450 334.050 ;
        RECT 176.250 333.600 177.450 335.700 ;
        RECT 163.650 327.750 165.450 332.700 ;
        RECT 166.650 327.750 168.450 331.800 ;
        RECT 169.650 327.750 171.450 332.700 ;
        RECT 175.650 327.750 177.450 333.600 ;
        RECT 178.650 332.700 186.450 334.050 ;
        RECT 178.650 327.750 180.450 332.700 ;
        RECT 181.650 327.750 183.450 331.800 ;
        RECT 184.650 327.750 186.450 332.700 ;
        RECT 189.150 333.600 190.050 346.200 ;
        RECT 198.450 345.900 206.850 346.200 ;
        RECT 208.050 346.800 214.050 347.700 ;
        RECT 214.950 346.800 217.050 347.700 ;
        RECT 220.650 347.400 222.450 359.250 ;
        RECT 227.400 353.400 229.200 359.250 ;
        RECT 230.700 347.400 232.500 359.250 ;
        RECT 234.900 347.400 236.700 359.250 ;
        RECT 240.150 347.400 241.950 359.250 ;
        RECT 243.150 353.400 244.950 359.250 ;
        RECT 248.250 353.400 250.050 359.250 ;
        RECT 253.050 353.400 254.850 359.250 ;
        RECT 248.550 352.500 249.750 353.400 ;
        RECT 256.050 352.500 257.850 359.250 ;
        RECT 259.950 353.400 261.750 359.250 ;
        RECT 264.150 353.400 265.950 359.250 ;
        RECT 268.650 356.400 270.450 359.250 ;
        RECT 244.950 350.400 249.750 352.500 ;
        RECT 252.150 350.700 259.050 352.500 ;
        RECT 264.150 351.300 268.050 353.400 ;
        RECT 248.550 349.500 249.750 350.400 ;
        RECT 261.450 349.800 263.250 350.400 ;
        RECT 248.550 348.300 256.050 349.500 ;
        RECT 254.250 347.700 256.050 348.300 ;
        RECT 256.950 348.900 263.250 349.800 ;
        RECT 198.450 345.600 200.250 345.900 ;
        RECT 208.050 342.150 208.950 346.800 ;
        RECT 214.950 345.600 219.150 346.800 ;
        RECT 218.250 343.800 220.050 345.600 ;
        RECT 199.950 341.100 202.050 342.150 ;
        RECT 191.100 339.150 192.900 340.950 ;
        RECT 194.100 340.050 202.050 341.100 ;
        RECT 205.950 340.050 208.950 342.150 ;
        RECT 194.100 339.300 195.900 340.050 ;
        RECT 192.000 338.400 192.900 339.150 ;
        RECT 197.100 338.400 198.900 339.000 ;
        RECT 192.000 337.200 198.900 338.400 ;
        RECT 197.850 336.000 198.900 337.200 ;
        RECT 208.050 336.000 208.950 340.050 ;
        RECT 217.950 339.750 220.050 340.050 ;
        RECT 216.150 337.950 220.050 339.750 ;
        RECT 221.250 337.950 222.450 347.400 ;
        RECT 227.250 345.150 229.050 346.950 ;
        RECT 226.950 343.050 229.050 345.150 ;
        RECT 230.850 342.150 232.050 347.400 ;
        RECT 240.150 346.800 251.250 347.400 ;
        RECT 256.950 346.800 257.850 348.900 ;
        RECT 261.450 348.600 263.250 348.900 ;
        RECT 264.150 348.600 266.850 350.400 ;
        RECT 264.150 347.700 265.050 348.600 ;
        RECT 240.150 346.200 257.850 346.800 ;
        RECT 236.100 342.150 237.900 343.950 ;
        RECT 197.850 335.100 208.950 336.000 ;
        RECT 217.950 335.850 222.450 337.950 ;
        RECT 229.950 340.050 232.050 342.150 ;
        RECT 229.950 336.750 231.150 340.050 ;
        RECT 232.950 338.850 235.050 340.950 ;
        RECT 235.950 340.050 238.050 342.150 ;
        RECT 233.100 337.050 234.900 338.850 ;
        RECT 197.850 334.200 198.900 335.100 ;
        RECT 208.050 334.800 208.950 335.100 ;
        RECT 189.150 327.750 190.950 333.600 ;
        RECT 193.950 331.500 196.050 333.600 ;
        RECT 197.550 332.400 199.350 334.200 ;
        RECT 200.850 333.450 202.650 334.200 ;
        RECT 200.850 332.400 205.800 333.450 ;
        RECT 208.050 333.000 209.850 334.800 ;
        RECT 221.250 333.600 222.450 335.850 ;
        RECT 227.250 335.700 231.000 336.750 ;
        RECT 227.250 333.600 228.450 335.700 ;
        RECT 214.950 332.700 217.050 333.600 ;
        RECT 195.000 330.600 196.050 331.500 ;
        RECT 204.750 330.600 205.800 332.400 ;
        RECT 213.300 331.500 217.050 332.700 ;
        RECT 213.300 330.600 214.350 331.500 ;
        RECT 192.150 327.750 193.950 330.600 ;
        RECT 195.000 329.700 198.750 330.600 ;
        RECT 196.950 327.750 198.750 329.700 ;
        RECT 201.450 327.750 203.250 330.600 ;
        RECT 204.750 327.750 206.550 330.600 ;
        RECT 208.650 327.750 210.450 330.600 ;
        RECT 212.850 327.750 214.650 330.600 ;
        RECT 217.350 327.750 219.150 330.600 ;
        RECT 220.650 327.750 222.450 333.600 ;
        RECT 226.650 327.750 228.450 333.600 ;
        RECT 229.650 332.700 237.450 334.050 ;
        RECT 229.650 327.750 231.450 332.700 ;
        RECT 232.650 327.750 234.450 331.800 ;
        RECT 235.650 327.750 237.450 332.700 ;
        RECT 240.150 333.600 241.050 346.200 ;
        RECT 249.450 345.900 257.850 346.200 ;
        RECT 259.050 346.800 265.050 347.700 ;
        RECT 265.950 346.800 268.050 347.700 ;
        RECT 271.650 347.400 273.450 359.250 ;
        RECT 277.650 353.400 279.450 359.250 ;
        RECT 280.650 353.400 282.450 359.250 ;
        RECT 286.650 353.400 288.450 359.250 ;
        RECT 289.650 353.400 291.450 359.250 ;
        RECT 249.450 345.600 251.250 345.900 ;
        RECT 259.050 342.150 259.950 346.800 ;
        RECT 265.950 345.600 270.150 346.800 ;
        RECT 269.250 343.800 271.050 345.600 ;
        RECT 250.950 341.100 253.050 342.150 ;
        RECT 242.100 339.150 243.900 340.950 ;
        RECT 245.100 340.050 253.050 341.100 ;
        RECT 256.950 340.050 259.950 342.150 ;
        RECT 245.100 339.300 246.900 340.050 ;
        RECT 243.000 338.400 243.900 339.150 ;
        RECT 248.100 338.400 249.900 339.000 ;
        RECT 243.000 337.200 249.900 338.400 ;
        RECT 248.850 336.000 249.900 337.200 ;
        RECT 259.050 336.000 259.950 340.050 ;
        RECT 268.950 339.750 271.050 340.050 ;
        RECT 267.150 337.950 271.050 339.750 ;
        RECT 272.250 337.950 273.450 347.400 ;
        RECT 278.400 340.950 279.600 353.400 ;
        RECT 287.400 340.950 288.600 353.400 ;
        RECT 294.300 347.400 296.100 359.250 ;
        RECT 298.500 347.400 300.300 359.250 ;
        RECT 301.800 353.400 303.600 359.250 ;
        RECT 309.150 347.400 310.950 359.250 ;
        RECT 312.150 353.400 313.950 359.250 ;
        RECT 317.250 353.400 319.050 359.250 ;
        RECT 322.050 353.400 323.850 359.250 ;
        RECT 317.550 352.500 318.750 353.400 ;
        RECT 325.050 352.500 326.850 359.250 ;
        RECT 328.950 353.400 330.750 359.250 ;
        RECT 333.150 353.400 334.950 359.250 ;
        RECT 337.650 356.400 339.450 359.250 ;
        RECT 313.950 350.400 318.750 352.500 ;
        RECT 321.150 350.700 328.050 352.500 ;
        RECT 333.150 351.300 337.050 353.400 ;
        RECT 317.550 349.500 318.750 350.400 ;
        RECT 330.450 349.800 332.250 350.400 ;
        RECT 317.550 348.300 325.050 349.500 ;
        RECT 323.250 347.700 325.050 348.300 ;
        RECT 325.950 348.900 332.250 349.800 ;
        RECT 293.100 342.150 294.900 343.950 ;
        RECT 298.950 342.150 300.150 347.400 ;
        RECT 301.950 345.150 303.750 346.950 ;
        RECT 309.150 346.800 320.250 347.400 ;
        RECT 325.950 346.800 326.850 348.900 ;
        RECT 330.450 348.600 332.250 348.900 ;
        RECT 333.150 348.600 335.850 350.400 ;
        RECT 333.150 347.700 334.050 348.600 ;
        RECT 309.150 346.200 326.850 346.800 ;
        RECT 301.950 343.050 304.050 345.150 ;
        RECT 277.950 338.850 280.050 340.950 ;
        RECT 281.100 339.150 282.900 340.950 ;
        RECT 248.850 335.100 259.950 336.000 ;
        RECT 268.950 335.850 273.450 337.950 ;
        RECT 248.850 334.200 249.900 335.100 ;
        RECT 259.050 334.800 259.950 335.100 ;
        RECT 240.150 327.750 241.950 333.600 ;
        RECT 244.950 331.500 247.050 333.600 ;
        RECT 248.550 332.400 250.350 334.200 ;
        RECT 251.850 333.450 253.650 334.200 ;
        RECT 251.850 332.400 256.800 333.450 ;
        RECT 259.050 333.000 260.850 334.800 ;
        RECT 272.250 333.600 273.450 335.850 ;
        RECT 265.950 332.700 268.050 333.600 ;
        RECT 246.000 330.600 247.050 331.500 ;
        RECT 255.750 330.600 256.800 332.400 ;
        RECT 264.300 331.500 268.050 332.700 ;
        RECT 264.300 330.600 265.350 331.500 ;
        RECT 243.150 327.750 244.950 330.600 ;
        RECT 246.000 329.700 249.750 330.600 ;
        RECT 247.950 327.750 249.750 329.700 ;
        RECT 252.450 327.750 254.250 330.600 ;
        RECT 255.750 327.750 257.550 330.600 ;
        RECT 259.650 327.750 261.450 330.600 ;
        RECT 263.850 327.750 265.650 330.600 ;
        RECT 268.350 327.750 270.150 330.600 ;
        RECT 271.650 327.750 273.450 333.600 ;
        RECT 278.400 330.600 279.600 338.850 ;
        RECT 280.950 337.050 283.050 339.150 ;
        RECT 286.950 338.850 289.050 340.950 ;
        RECT 290.100 339.150 291.900 340.950 ;
        RECT 292.950 340.050 295.050 342.150 ;
        RECT 287.400 330.600 288.600 338.850 ;
        RECT 289.950 337.050 292.050 339.150 ;
        RECT 295.950 338.850 298.050 340.950 ;
        RECT 298.950 340.050 301.050 342.150 ;
        RECT 296.100 337.050 297.900 338.850 ;
        RECT 299.850 336.750 301.050 340.050 ;
        RECT 300.000 335.700 303.750 336.750 ;
        RECT 293.550 332.700 301.350 334.050 ;
        RECT 277.650 327.750 279.450 330.600 ;
        RECT 280.650 327.750 282.450 330.600 ;
        RECT 286.650 327.750 288.450 330.600 ;
        RECT 289.650 327.750 291.450 330.600 ;
        RECT 293.550 327.750 295.350 332.700 ;
        RECT 296.550 327.750 298.350 331.800 ;
        RECT 299.550 327.750 301.350 332.700 ;
        RECT 302.550 333.600 303.750 335.700 ;
        RECT 309.150 333.600 310.050 346.200 ;
        RECT 318.450 345.900 326.850 346.200 ;
        RECT 328.050 346.800 334.050 347.700 ;
        RECT 334.950 346.800 337.050 347.700 ;
        RECT 340.650 347.400 342.450 359.250 ;
        RECT 346.650 347.400 348.450 359.250 ;
        RECT 349.650 348.300 351.450 359.250 ;
        RECT 352.650 349.200 354.450 359.250 ;
        RECT 355.650 348.300 357.450 359.250 ;
        RECT 349.650 347.400 357.450 348.300 ;
        RECT 361.650 347.400 363.450 359.250 ;
        RECT 364.650 348.300 366.450 359.250 ;
        RECT 367.650 349.200 369.450 359.250 ;
        RECT 370.650 348.300 372.450 359.250 ;
        RECT 374.550 353.400 376.350 359.250 ;
        RECT 377.550 353.400 379.350 359.250 ;
        RECT 380.550 354.000 382.350 359.250 ;
        RECT 377.700 353.100 379.350 353.400 ;
        RECT 383.550 353.400 385.350 359.250 ;
        RECT 389.550 353.400 391.350 359.250 ;
        RECT 392.550 353.400 394.350 359.250 ;
        RECT 383.550 353.100 384.750 353.400 ;
        RECT 377.700 352.200 384.750 353.100 ;
        RECT 364.650 347.400 372.450 348.300 ;
        RECT 377.100 348.150 378.900 349.950 ;
        RECT 318.450 345.600 320.250 345.900 ;
        RECT 328.050 342.150 328.950 346.800 ;
        RECT 334.950 345.600 339.150 346.800 ;
        RECT 338.250 343.800 340.050 345.600 ;
        RECT 319.950 341.100 322.050 342.150 ;
        RECT 311.100 339.150 312.900 340.950 ;
        RECT 314.100 340.050 322.050 341.100 ;
        RECT 325.950 340.050 328.950 342.150 ;
        RECT 314.100 339.300 315.900 340.050 ;
        RECT 312.000 338.400 312.900 339.150 ;
        RECT 317.100 338.400 318.900 339.000 ;
        RECT 312.000 337.200 318.900 338.400 ;
        RECT 317.850 336.000 318.900 337.200 ;
        RECT 328.050 336.000 328.950 340.050 ;
        RECT 337.950 339.750 340.050 340.050 ;
        RECT 336.150 337.950 340.050 339.750 ;
        RECT 341.250 337.950 342.450 347.400 ;
        RECT 347.100 342.150 348.300 347.400 ;
        RECT 362.100 342.150 363.300 347.400 ;
        RECT 374.100 345.150 375.900 346.950 ;
        RECT 376.950 346.050 379.050 348.150 ;
        RECT 380.250 345.150 382.050 346.950 ;
        RECT 373.950 343.050 376.050 345.150 ;
        RECT 379.950 343.050 382.050 345.150 ;
        RECT 383.700 343.950 384.750 352.200 ;
        RECT 346.950 340.050 349.050 342.150 ;
        RECT 317.850 335.100 328.950 336.000 ;
        RECT 337.950 335.850 342.450 337.950 ;
        RECT 317.850 334.200 318.900 335.100 ;
        RECT 328.050 334.800 328.950 335.100 ;
        RECT 302.550 327.750 304.350 333.600 ;
        RECT 309.150 327.750 310.950 333.600 ;
        RECT 313.950 331.500 316.050 333.600 ;
        RECT 317.550 332.400 319.350 334.200 ;
        RECT 320.850 333.450 322.650 334.200 ;
        RECT 320.850 332.400 325.800 333.450 ;
        RECT 328.050 333.000 329.850 334.800 ;
        RECT 341.250 333.600 342.450 335.850 ;
        RECT 334.950 332.700 337.050 333.600 ;
        RECT 315.000 330.600 316.050 331.500 ;
        RECT 324.750 330.600 325.800 332.400 ;
        RECT 333.300 331.500 337.050 332.700 ;
        RECT 333.300 330.600 334.350 331.500 ;
        RECT 312.150 327.750 313.950 330.600 ;
        RECT 315.000 329.700 318.750 330.600 ;
        RECT 316.950 327.750 318.750 329.700 ;
        RECT 321.450 327.750 323.250 330.600 ;
        RECT 324.750 327.750 326.550 330.600 ;
        RECT 328.650 327.750 330.450 330.600 ;
        RECT 332.850 327.750 334.650 330.600 ;
        RECT 337.350 327.750 339.150 330.600 ;
        RECT 340.650 327.750 342.450 333.600 ;
        RECT 347.100 333.600 348.300 340.050 ;
        RECT 349.950 338.850 352.050 340.950 ;
        RECT 353.100 339.150 354.900 340.950 ;
        RECT 350.100 337.050 351.900 338.850 ;
        RECT 352.950 337.050 355.050 339.150 ;
        RECT 355.950 338.850 358.050 340.950 ;
        RECT 361.950 340.050 364.050 342.150 ;
        RECT 382.950 341.850 385.050 343.950 ;
        RECT 389.100 342.150 390.900 343.950 ;
        RECT 356.100 337.050 357.900 338.850 ;
        RECT 362.100 333.600 363.300 340.050 ;
        RECT 364.950 338.850 367.050 340.950 ;
        RECT 368.100 339.150 369.900 340.950 ;
        RECT 365.100 337.050 366.900 338.850 ;
        RECT 367.950 337.050 370.050 339.150 ;
        RECT 370.950 338.850 373.050 340.950 ;
        RECT 371.100 337.050 372.900 338.850 ;
        RECT 383.400 337.650 384.600 341.850 ;
        RECT 388.950 340.050 391.050 342.150 ;
        RECT 347.100 331.950 352.800 333.600 ;
        RECT 347.700 327.750 349.500 330.600 ;
        RECT 351.000 327.750 352.800 331.950 ;
        RECT 355.200 327.750 357.000 333.600 ;
        RECT 362.100 331.950 367.800 333.600 ;
        RECT 362.700 327.750 364.500 330.600 ;
        RECT 366.000 327.750 367.800 331.950 ;
        RECT 370.200 327.750 372.000 333.600 ;
        RECT 374.700 327.750 376.500 336.600 ;
        RECT 380.100 336.000 384.600 337.650 ;
        RECT 392.700 336.300 393.900 353.400 ;
        RECT 396.150 347.400 397.950 359.250 ;
        RECT 399.150 347.400 400.950 359.250 ;
        RECT 404.550 347.400 406.350 359.250 ;
        RECT 407.550 356.400 409.350 359.250 ;
        RECT 412.050 353.400 413.850 359.250 ;
        RECT 416.250 353.400 418.050 359.250 ;
        RECT 409.950 351.300 413.850 353.400 ;
        RECT 420.150 352.500 421.950 359.250 ;
        RECT 423.150 353.400 424.950 359.250 ;
        RECT 427.950 353.400 429.750 359.250 ;
        RECT 433.050 353.400 434.850 359.250 ;
        RECT 428.250 352.500 429.450 353.400 ;
        RECT 418.950 350.700 425.850 352.500 ;
        RECT 428.250 350.400 433.050 352.500 ;
        RECT 411.150 348.600 413.850 350.400 ;
        RECT 414.750 349.800 416.550 350.400 ;
        RECT 414.750 348.900 421.050 349.800 ;
        RECT 428.250 349.500 429.450 350.400 ;
        RECT 414.750 348.600 416.550 348.900 ;
        RECT 412.950 347.700 413.850 348.600 ;
        RECT 394.950 341.850 397.050 343.950 ;
        RECT 399.150 342.150 400.350 347.400 ;
        RECT 395.100 340.050 396.900 341.850 ;
        RECT 397.950 340.050 400.350 342.150 ;
        RECT 380.100 327.750 381.900 336.000 ;
        RECT 389.550 335.100 397.050 336.300 ;
        RECT 389.550 327.750 391.350 335.100 ;
        RECT 395.250 334.500 397.050 335.100 ;
        RECT 399.150 333.600 400.350 340.050 ;
        RECT 394.050 327.750 395.850 333.600 ;
        RECT 397.050 332.100 400.350 333.600 ;
        RECT 404.550 337.950 405.750 347.400 ;
        RECT 409.950 346.800 412.050 347.700 ;
        RECT 412.950 346.800 418.950 347.700 ;
        RECT 407.850 345.600 412.050 346.800 ;
        RECT 406.950 343.800 408.750 345.600 ;
        RECT 418.050 342.150 418.950 346.800 ;
        RECT 420.150 346.800 421.050 348.900 ;
        RECT 421.950 348.300 429.450 349.500 ;
        RECT 421.950 347.700 423.750 348.300 ;
        RECT 436.050 347.400 437.850 359.250 ;
        RECT 443.400 353.400 445.200 359.250 ;
        RECT 446.700 347.400 448.500 359.250 ;
        RECT 450.900 347.400 452.700 359.250 ;
        RECT 458.400 353.400 460.200 359.250 ;
        RECT 461.700 347.400 463.500 359.250 ;
        RECT 465.900 347.400 467.700 359.250 ;
        RECT 471.300 347.400 473.100 359.250 ;
        RECT 475.500 347.400 477.300 359.250 ;
        RECT 478.800 353.400 480.600 359.250 ;
        RECT 485.550 347.400 487.350 359.250 ;
        RECT 488.550 356.400 490.350 359.250 ;
        RECT 493.050 353.400 494.850 359.250 ;
        RECT 497.250 353.400 499.050 359.250 ;
        RECT 490.950 351.300 494.850 353.400 ;
        RECT 501.150 352.500 502.950 359.250 ;
        RECT 504.150 353.400 505.950 359.250 ;
        RECT 508.950 353.400 510.750 359.250 ;
        RECT 514.050 353.400 515.850 359.250 ;
        RECT 509.250 352.500 510.450 353.400 ;
        RECT 499.950 350.700 506.850 352.500 ;
        RECT 509.250 350.400 514.050 352.500 ;
        RECT 492.150 348.600 494.850 350.400 ;
        RECT 495.750 349.800 497.550 350.400 ;
        RECT 495.750 348.900 502.050 349.800 ;
        RECT 509.250 349.500 510.450 350.400 ;
        RECT 495.750 348.600 497.550 348.900 ;
        RECT 493.950 347.700 494.850 348.600 ;
        RECT 426.750 346.800 437.850 347.400 ;
        RECT 420.150 346.200 437.850 346.800 ;
        RECT 420.150 345.900 428.550 346.200 ;
        RECT 426.750 345.600 428.550 345.900 ;
        RECT 418.050 340.050 421.050 342.150 ;
        RECT 424.950 341.100 427.050 342.150 ;
        RECT 424.950 340.050 432.900 341.100 ;
        RECT 406.950 339.750 409.050 340.050 ;
        RECT 406.950 337.950 410.850 339.750 ;
        RECT 404.550 335.850 409.050 337.950 ;
        RECT 418.050 336.000 418.950 340.050 ;
        RECT 431.100 339.300 432.900 340.050 ;
        RECT 434.100 339.150 435.900 340.950 ;
        RECT 428.100 338.400 429.900 339.000 ;
        RECT 434.100 338.400 435.000 339.150 ;
        RECT 428.100 337.200 435.000 338.400 ;
        RECT 428.100 336.000 429.150 337.200 ;
        RECT 404.550 333.600 405.750 335.850 ;
        RECT 418.050 335.100 429.150 336.000 ;
        RECT 418.050 334.800 418.950 335.100 ;
        RECT 397.050 327.750 398.850 332.100 ;
        RECT 404.550 327.750 406.350 333.600 ;
        RECT 409.950 332.700 412.050 333.600 ;
        RECT 417.150 333.000 418.950 334.800 ;
        RECT 428.100 334.200 429.150 335.100 ;
        RECT 424.350 333.450 426.150 334.200 ;
        RECT 409.950 331.500 413.700 332.700 ;
        RECT 412.650 330.600 413.700 331.500 ;
        RECT 421.200 332.400 426.150 333.450 ;
        RECT 427.650 332.400 429.450 334.200 ;
        RECT 436.950 333.600 437.850 346.200 ;
        RECT 443.250 345.150 445.050 346.950 ;
        RECT 442.950 343.050 445.050 345.150 ;
        RECT 446.850 342.150 448.050 347.400 ;
        RECT 458.250 345.150 460.050 346.950 ;
        RECT 452.100 342.150 453.900 343.950 ;
        RECT 457.950 343.050 460.050 345.150 ;
        RECT 461.850 342.150 463.050 347.400 ;
        RECT 467.100 342.150 468.900 343.950 ;
        RECT 470.100 342.150 471.900 343.950 ;
        RECT 475.950 342.150 477.150 347.400 ;
        RECT 478.950 345.150 480.750 346.950 ;
        RECT 478.950 343.050 481.050 345.150 ;
        RECT 445.950 340.050 448.050 342.150 ;
        RECT 445.950 336.750 447.150 340.050 ;
        RECT 448.950 338.850 451.050 340.950 ;
        RECT 451.950 340.050 454.050 342.150 ;
        RECT 460.950 340.050 463.050 342.150 ;
        RECT 449.100 337.050 450.900 338.850 ;
        RECT 460.950 336.750 462.150 340.050 ;
        RECT 463.950 338.850 466.050 340.950 ;
        RECT 466.950 340.050 469.050 342.150 ;
        RECT 469.950 340.050 472.050 342.150 ;
        RECT 472.950 338.850 475.050 340.950 ;
        RECT 475.950 340.050 478.050 342.150 ;
        RECT 464.100 337.050 465.900 338.850 ;
        RECT 473.100 337.050 474.900 338.850 ;
        RECT 476.850 336.750 478.050 340.050 ;
        RECT 485.550 337.950 486.750 347.400 ;
        RECT 490.950 346.800 493.050 347.700 ;
        RECT 493.950 346.800 499.950 347.700 ;
        RECT 488.850 345.600 493.050 346.800 ;
        RECT 487.950 343.800 489.750 345.600 ;
        RECT 499.050 342.150 499.950 346.800 ;
        RECT 501.150 346.800 502.050 348.900 ;
        RECT 502.950 348.300 510.450 349.500 ;
        RECT 502.950 347.700 504.750 348.300 ;
        RECT 517.050 347.400 518.850 359.250 ;
        RECT 524.400 353.400 526.200 359.250 ;
        RECT 527.700 347.400 529.500 359.250 ;
        RECT 531.900 347.400 533.700 359.250 ;
        RECT 540.450 347.400 542.250 359.250 ;
        RECT 544.650 347.400 546.450 359.250 ;
        RECT 548.550 347.400 550.350 359.250 ;
        RECT 553.050 347.550 554.850 359.250 ;
        RECT 556.050 348.900 557.850 359.250 ;
        RECT 565.650 353.400 567.450 359.250 ;
        RECT 568.650 353.400 570.450 359.250 ;
        RECT 571.650 353.400 573.450 359.250 ;
        RECT 577.650 358.500 585.450 359.250 ;
        RECT 556.050 347.550 558.450 348.900 ;
        RECT 565.950 348.450 568.050 349.050 ;
        RECT 507.750 346.800 518.850 347.400 ;
        RECT 501.150 346.200 518.850 346.800 ;
        RECT 501.150 345.900 509.550 346.200 ;
        RECT 507.750 345.600 509.550 345.900 ;
        RECT 499.050 340.050 502.050 342.150 ;
        RECT 505.950 341.100 508.050 342.150 ;
        RECT 505.950 340.050 513.900 341.100 ;
        RECT 487.950 339.750 490.050 340.050 ;
        RECT 487.950 337.950 491.850 339.750 ;
        RECT 443.250 335.700 447.000 336.750 ;
        RECT 458.250 335.700 462.000 336.750 ;
        RECT 477.000 335.700 480.750 336.750 ;
        RECT 443.250 333.600 444.450 335.700 ;
        RECT 421.200 330.600 422.250 332.400 ;
        RECT 430.950 331.500 433.050 333.600 ;
        RECT 430.950 330.600 432.000 331.500 ;
        RECT 407.850 327.750 409.650 330.600 ;
        RECT 412.350 327.750 414.150 330.600 ;
        RECT 416.550 327.750 418.350 330.600 ;
        RECT 420.450 327.750 422.250 330.600 ;
        RECT 423.750 327.750 425.550 330.600 ;
        RECT 428.250 329.700 432.000 330.600 ;
        RECT 428.250 327.750 430.050 329.700 ;
        RECT 433.050 327.750 434.850 330.600 ;
        RECT 436.050 327.750 437.850 333.600 ;
        RECT 442.650 327.750 444.450 333.600 ;
        RECT 445.650 332.700 453.450 334.050 ;
        RECT 458.250 333.600 459.450 335.700 ;
        RECT 445.650 327.750 447.450 332.700 ;
        RECT 448.650 327.750 450.450 331.800 ;
        RECT 451.650 327.750 453.450 332.700 ;
        RECT 457.650 327.750 459.450 333.600 ;
        RECT 460.650 332.700 468.450 334.050 ;
        RECT 460.650 327.750 462.450 332.700 ;
        RECT 463.650 327.750 465.450 331.800 ;
        RECT 466.650 327.750 468.450 332.700 ;
        RECT 470.550 332.700 478.350 334.050 ;
        RECT 470.550 327.750 472.350 332.700 ;
        RECT 473.550 327.750 475.350 331.800 ;
        RECT 476.550 327.750 478.350 332.700 ;
        RECT 479.550 333.600 480.750 335.700 ;
        RECT 485.550 335.850 490.050 337.950 ;
        RECT 499.050 336.000 499.950 340.050 ;
        RECT 512.100 339.300 513.900 340.050 ;
        RECT 515.100 339.150 516.900 340.950 ;
        RECT 509.100 338.400 510.900 339.000 ;
        RECT 515.100 338.400 516.000 339.150 ;
        RECT 509.100 337.200 516.000 338.400 ;
        RECT 509.100 336.000 510.150 337.200 ;
        RECT 485.550 333.600 486.750 335.850 ;
        RECT 499.050 335.100 510.150 336.000 ;
        RECT 499.050 334.800 499.950 335.100 ;
        RECT 479.550 327.750 481.350 333.600 ;
        RECT 485.550 327.750 487.350 333.600 ;
        RECT 490.950 332.700 493.050 333.600 ;
        RECT 498.150 333.000 499.950 334.800 ;
        RECT 509.100 334.200 510.150 335.100 ;
        RECT 505.350 333.450 507.150 334.200 ;
        RECT 490.950 331.500 494.700 332.700 ;
        RECT 493.650 330.600 494.700 331.500 ;
        RECT 502.200 332.400 507.150 333.450 ;
        RECT 508.650 332.400 510.450 334.200 ;
        RECT 517.950 333.600 518.850 346.200 ;
        RECT 524.250 345.150 526.050 346.950 ;
        RECT 523.950 343.050 526.050 345.150 ;
        RECT 527.850 342.150 529.050 347.400 ;
        RECT 540.450 346.350 543.000 347.400 ;
        RECT 533.100 342.150 534.900 343.950 ;
        RECT 539.100 342.150 540.900 343.950 ;
        RECT 526.950 340.050 529.050 342.150 ;
        RECT 526.950 336.750 528.150 340.050 ;
        RECT 529.950 338.850 532.050 340.950 ;
        RECT 532.950 340.050 535.050 342.150 ;
        RECT 538.950 340.050 541.050 342.150 ;
        RECT 541.950 339.150 543.000 346.350 ;
        RECT 548.550 346.200 549.750 347.400 ;
        RECT 553.950 346.200 555.750 346.650 ;
        RECT 548.550 345.000 555.750 346.200 ;
        RECT 553.950 344.850 555.750 345.000 ;
        RECT 545.100 342.150 546.900 343.950 ;
        RECT 551.100 342.150 552.900 343.950 ;
        RECT 544.950 340.050 547.050 342.150 ;
        RECT 548.100 339.150 549.900 340.950 ;
        RECT 550.950 340.050 553.050 342.150 ;
        RECT 530.100 337.050 531.900 338.850 ;
        RECT 541.950 337.050 544.050 339.150 ;
        RECT 547.950 337.050 550.050 339.150 ;
        RECT 524.250 335.700 528.000 336.750 ;
        RECT 524.250 333.600 525.450 335.700 ;
        RECT 502.200 330.600 503.250 332.400 ;
        RECT 511.950 331.500 514.050 333.600 ;
        RECT 511.950 330.600 513.000 331.500 ;
        RECT 488.850 327.750 490.650 330.600 ;
        RECT 493.350 327.750 495.150 330.600 ;
        RECT 497.550 327.750 499.350 330.600 ;
        RECT 501.450 327.750 503.250 330.600 ;
        RECT 504.750 327.750 506.550 330.600 ;
        RECT 509.250 329.700 513.000 330.600 ;
        RECT 509.250 327.750 511.050 329.700 ;
        RECT 514.050 327.750 515.850 330.600 ;
        RECT 517.050 327.750 518.850 333.600 ;
        RECT 523.650 327.750 525.450 333.600 ;
        RECT 526.650 332.700 534.450 334.050 ;
        RECT 526.650 327.750 528.450 332.700 ;
        RECT 529.650 327.750 531.450 331.800 ;
        RECT 532.650 327.750 534.450 332.700 ;
        RECT 541.950 330.600 543.000 337.050 ;
        RECT 554.700 336.600 555.600 344.850 ;
        RECT 557.100 340.950 558.450 347.550 ;
        RECT 560.550 347.550 568.050 348.450 ;
        RECT 560.550 343.050 561.450 347.550 ;
        RECT 565.950 346.950 568.050 347.550 ;
        RECT 569.250 345.150 570.450 353.400 ;
        RECT 577.650 347.400 579.450 358.500 ;
        RECT 580.650 347.400 582.450 357.600 ;
        RECT 583.650 348.600 585.450 358.500 ;
        RECT 586.650 349.500 588.450 359.250 ;
        RECT 589.650 348.600 591.450 359.250 ;
        RECT 583.650 347.700 591.450 348.600 ;
        RECT 595.650 358.500 603.450 359.250 ;
        RECT 595.650 347.400 597.450 358.500 ;
        RECT 598.650 347.400 600.450 357.600 ;
        RECT 601.650 348.600 603.450 358.500 ;
        RECT 604.650 349.500 606.450 359.250 ;
        RECT 607.650 348.600 609.450 359.250 ;
        RECT 601.650 347.700 609.450 348.600 ;
        RECT 612.150 347.400 613.950 359.250 ;
        RECT 615.150 353.400 616.950 359.250 ;
        RECT 620.250 353.400 622.050 359.250 ;
        RECT 625.050 353.400 626.850 359.250 ;
        RECT 620.550 352.500 621.750 353.400 ;
        RECT 628.050 352.500 629.850 359.250 ;
        RECT 631.950 353.400 633.750 359.250 ;
        RECT 636.150 353.400 637.950 359.250 ;
        RECT 640.650 356.400 642.450 359.250 ;
        RECT 616.950 350.400 621.750 352.500 ;
        RECT 624.150 350.700 631.050 352.500 ;
        RECT 636.150 351.300 640.050 353.400 ;
        RECT 620.550 349.500 621.750 350.400 ;
        RECT 633.450 349.800 635.250 350.400 ;
        RECT 620.550 348.300 628.050 349.500 ;
        RECT 626.250 347.700 628.050 348.300 ;
        RECT 628.950 348.900 635.250 349.800 ;
        RECT 580.800 346.500 582.600 347.400 ;
        RECT 598.800 346.500 600.600 347.400 ;
        RECT 612.150 346.800 623.250 347.400 ;
        RECT 628.950 346.800 629.850 348.900 ;
        RECT 633.450 348.600 635.250 348.900 ;
        RECT 636.150 348.600 638.850 350.400 ;
        RECT 636.150 347.700 637.050 348.600 ;
        RECT 580.800 345.600 584.850 346.500 ;
        RECT 559.950 340.950 562.050 343.050 ;
        RECT 565.950 341.850 568.050 343.950 ;
        RECT 568.950 343.050 571.050 345.150 ;
        RECT 556.950 338.850 559.050 340.950 ;
        RECT 566.100 340.050 567.900 341.850 ;
        RECT 553.950 335.700 555.750 336.600 ;
        RECT 552.450 334.800 555.750 335.700 ;
        RECT 552.450 330.600 553.350 334.800 ;
        RECT 558.000 333.600 559.050 338.850 ;
        RECT 569.250 335.700 570.450 343.050 ;
        RECT 571.950 341.850 574.050 343.950 ;
        RECT 578.100 342.150 579.900 343.950 ;
        RECT 583.950 342.150 584.850 345.600 ;
        RECT 592.950 343.950 595.050 346.050 ;
        RECT 598.800 345.600 602.850 346.500 ;
        RECT 589.950 342.150 591.750 343.950 ;
        RECT 572.100 340.050 573.900 341.850 ;
        RECT 577.950 340.050 580.050 342.150 ;
        RECT 580.950 338.850 583.050 340.950 ;
        RECT 583.950 340.050 586.050 342.150 ;
        RECT 581.250 337.050 583.050 338.850 ;
        RECT 566.850 334.800 570.450 335.700 ;
        RECT 538.650 327.750 540.450 330.600 ;
        RECT 541.650 327.750 543.450 330.600 ;
        RECT 544.650 327.750 546.450 330.600 ;
        RECT 548.550 327.750 550.350 330.600 ;
        RECT 551.550 327.750 553.350 330.600 ;
        RECT 554.550 327.750 556.350 330.600 ;
        RECT 557.550 327.750 559.350 333.600 ;
        RECT 566.850 327.750 568.650 334.800 ;
        RECT 585.000 333.600 586.050 340.050 ;
        RECT 586.950 338.850 589.050 340.950 ;
        RECT 589.950 340.050 592.050 342.150 ;
        RECT 586.950 337.050 588.750 338.850 ;
        RECT 589.950 336.450 592.050 337.050 ;
        RECT 593.550 336.450 594.450 343.950 ;
        RECT 596.100 342.150 597.900 343.950 ;
        RECT 601.950 342.150 602.850 345.600 ;
        RECT 612.150 346.200 629.850 346.800 ;
        RECT 607.950 342.150 609.750 343.950 ;
        RECT 595.950 340.050 598.050 342.150 ;
        RECT 598.950 338.850 601.050 340.950 ;
        RECT 601.950 340.050 604.050 342.150 ;
        RECT 599.250 337.050 601.050 338.850 ;
        RECT 589.950 335.550 594.450 336.450 ;
        RECT 589.950 334.950 592.050 335.550 ;
        RECT 603.000 333.600 604.050 340.050 ;
        RECT 604.950 338.850 607.050 340.950 ;
        RECT 607.950 340.050 610.050 342.150 ;
        RECT 604.950 337.050 606.750 338.850 ;
        RECT 612.150 333.600 613.050 346.200 ;
        RECT 621.450 345.900 629.850 346.200 ;
        RECT 631.050 346.800 637.050 347.700 ;
        RECT 637.950 346.800 640.050 347.700 ;
        RECT 643.650 347.400 645.450 359.250 ;
        RECT 621.450 345.600 623.250 345.900 ;
        RECT 631.050 342.150 631.950 346.800 ;
        RECT 637.950 345.600 642.150 346.800 ;
        RECT 641.250 343.800 643.050 345.600 ;
        RECT 622.950 341.100 625.050 342.150 ;
        RECT 614.100 339.150 615.900 340.950 ;
        RECT 617.100 340.050 625.050 341.100 ;
        RECT 628.950 340.050 631.950 342.150 ;
        RECT 617.100 339.300 618.900 340.050 ;
        RECT 615.000 338.400 615.900 339.150 ;
        RECT 620.100 338.400 621.900 339.000 ;
        RECT 615.000 337.200 621.900 338.400 ;
        RECT 620.850 336.000 621.900 337.200 ;
        RECT 631.050 336.000 631.950 340.050 ;
        RECT 640.950 339.750 643.050 340.050 ;
        RECT 639.150 337.950 643.050 339.750 ;
        RECT 644.250 337.950 645.450 347.400 ;
        RECT 620.850 335.100 631.950 336.000 ;
        RECT 640.950 335.850 645.450 337.950 ;
        RECT 620.850 334.200 621.900 335.100 ;
        RECT 631.050 334.800 631.950 335.100 ;
        RECT 571.350 327.750 573.150 333.600 ;
        RECT 580.800 327.750 582.600 333.600 ;
        RECT 585.000 327.750 586.800 333.600 ;
        RECT 589.200 327.750 591.000 333.600 ;
        RECT 598.800 327.750 600.600 333.600 ;
        RECT 603.000 327.750 604.800 333.600 ;
        RECT 607.200 327.750 609.000 333.600 ;
        RECT 612.150 327.750 613.950 333.600 ;
        RECT 616.950 331.500 619.050 333.600 ;
        RECT 620.550 332.400 622.350 334.200 ;
        RECT 623.850 333.450 625.650 334.200 ;
        RECT 623.850 332.400 628.800 333.450 ;
        RECT 631.050 333.000 632.850 334.800 ;
        RECT 644.250 333.600 645.450 335.850 ;
        RECT 637.950 332.700 640.050 333.600 ;
        RECT 618.000 330.600 619.050 331.500 ;
        RECT 627.750 330.600 628.800 332.400 ;
        RECT 636.300 331.500 640.050 332.700 ;
        RECT 636.300 330.600 637.350 331.500 ;
        RECT 615.150 327.750 616.950 330.600 ;
        RECT 618.000 329.700 621.750 330.600 ;
        RECT 619.950 327.750 621.750 329.700 ;
        RECT 624.450 327.750 626.250 330.600 ;
        RECT 627.750 327.750 629.550 330.600 ;
        RECT 631.650 327.750 633.450 330.600 ;
        RECT 635.850 327.750 637.650 330.600 ;
        RECT 640.350 327.750 642.150 330.600 ;
        RECT 643.650 327.750 645.450 333.600 ;
        RECT 647.550 347.400 649.350 359.250 ;
        RECT 650.550 356.400 652.350 359.250 ;
        RECT 655.050 353.400 656.850 359.250 ;
        RECT 659.250 353.400 661.050 359.250 ;
        RECT 652.950 351.300 656.850 353.400 ;
        RECT 663.150 352.500 664.950 359.250 ;
        RECT 666.150 353.400 667.950 359.250 ;
        RECT 670.950 353.400 672.750 359.250 ;
        RECT 676.050 353.400 677.850 359.250 ;
        RECT 671.250 352.500 672.450 353.400 ;
        RECT 661.950 350.700 668.850 352.500 ;
        RECT 671.250 350.400 676.050 352.500 ;
        RECT 654.150 348.600 656.850 350.400 ;
        RECT 657.750 349.800 659.550 350.400 ;
        RECT 657.750 348.900 664.050 349.800 ;
        RECT 671.250 349.500 672.450 350.400 ;
        RECT 657.750 348.600 659.550 348.900 ;
        RECT 655.950 347.700 656.850 348.600 ;
        RECT 647.550 337.950 648.750 347.400 ;
        RECT 652.950 346.800 655.050 347.700 ;
        RECT 655.950 346.800 661.950 347.700 ;
        RECT 650.850 345.600 655.050 346.800 ;
        RECT 649.950 343.800 651.750 345.600 ;
        RECT 661.050 342.150 661.950 346.800 ;
        RECT 663.150 346.800 664.050 348.900 ;
        RECT 664.950 348.300 672.450 349.500 ;
        RECT 664.950 347.700 666.750 348.300 ;
        RECT 679.050 347.400 680.850 359.250 ;
        RECT 684.300 347.400 686.100 359.250 ;
        RECT 688.500 347.400 690.300 359.250 ;
        RECT 691.800 353.400 693.600 359.250 ;
        RECT 698.550 353.400 700.350 359.250 ;
        RECT 701.550 353.400 703.350 359.250 ;
        RECT 704.550 353.400 706.350 359.250 ;
        RECT 669.750 346.800 680.850 347.400 ;
        RECT 663.150 346.200 680.850 346.800 ;
        RECT 663.150 345.900 671.550 346.200 ;
        RECT 669.750 345.600 671.550 345.900 ;
        RECT 661.050 340.050 664.050 342.150 ;
        RECT 667.950 341.100 670.050 342.150 ;
        RECT 667.950 340.050 675.900 341.100 ;
        RECT 649.950 339.750 652.050 340.050 ;
        RECT 649.950 337.950 653.850 339.750 ;
        RECT 647.550 335.850 652.050 337.950 ;
        RECT 661.050 336.000 661.950 340.050 ;
        RECT 674.100 339.300 675.900 340.050 ;
        RECT 677.100 339.150 678.900 340.950 ;
        RECT 671.100 338.400 672.900 339.000 ;
        RECT 677.100 338.400 678.000 339.150 ;
        RECT 671.100 337.200 678.000 338.400 ;
        RECT 671.100 336.000 672.150 337.200 ;
        RECT 647.550 333.600 648.750 335.850 ;
        RECT 661.050 335.100 672.150 336.000 ;
        RECT 661.050 334.800 661.950 335.100 ;
        RECT 647.550 327.750 649.350 333.600 ;
        RECT 652.950 332.700 655.050 333.600 ;
        RECT 660.150 333.000 661.950 334.800 ;
        RECT 671.100 334.200 672.150 335.100 ;
        RECT 667.350 333.450 669.150 334.200 ;
        RECT 652.950 331.500 656.700 332.700 ;
        RECT 655.650 330.600 656.700 331.500 ;
        RECT 664.200 332.400 669.150 333.450 ;
        RECT 670.650 332.400 672.450 334.200 ;
        RECT 679.950 333.600 680.850 346.200 ;
        RECT 683.100 342.150 684.900 343.950 ;
        RECT 688.950 342.150 690.150 347.400 ;
        RECT 691.950 345.150 693.750 346.950 ;
        RECT 701.550 345.150 702.750 353.400 ;
        RECT 691.950 343.050 694.050 345.150 ;
        RECT 682.950 340.050 685.050 342.150 ;
        RECT 685.950 338.850 688.050 340.950 ;
        RECT 688.950 340.050 691.050 342.150 ;
        RECT 697.950 341.850 700.050 343.950 ;
        RECT 700.950 343.050 703.050 345.150 ;
        RECT 698.100 340.050 699.900 341.850 ;
        RECT 686.100 337.050 687.900 338.850 ;
        RECT 689.850 336.750 691.050 340.050 ;
        RECT 690.000 335.700 693.750 336.750 ;
        RECT 664.200 330.600 665.250 332.400 ;
        RECT 673.950 331.500 676.050 333.600 ;
        RECT 673.950 330.600 675.000 331.500 ;
        RECT 650.850 327.750 652.650 330.600 ;
        RECT 655.350 327.750 657.150 330.600 ;
        RECT 659.550 327.750 661.350 330.600 ;
        RECT 663.450 327.750 665.250 330.600 ;
        RECT 666.750 327.750 668.550 330.600 ;
        RECT 671.250 329.700 675.000 330.600 ;
        RECT 671.250 327.750 673.050 329.700 ;
        RECT 676.050 327.750 677.850 330.600 ;
        RECT 679.050 327.750 680.850 333.600 ;
        RECT 683.550 332.700 691.350 334.050 ;
        RECT 683.550 327.750 685.350 332.700 ;
        RECT 686.550 327.750 688.350 331.800 ;
        RECT 689.550 327.750 691.350 332.700 ;
        RECT 692.550 333.600 693.750 335.700 ;
        RECT 701.550 335.700 702.750 343.050 ;
        RECT 703.950 341.850 706.050 343.950 ;
        RECT 704.100 340.050 705.900 341.850 ;
        RECT 701.550 334.800 705.150 335.700 ;
        RECT 692.550 327.750 694.350 333.600 ;
        RECT 698.850 327.750 700.650 333.600 ;
        RECT 703.350 327.750 705.150 334.800 ;
        RECT 4.350 317.400 6.150 323.250 ;
        RECT 7.350 317.400 9.150 323.250 ;
        RECT 10.650 320.400 12.450 323.250 ;
        RECT 4.650 310.950 5.850 317.400 ;
        RECT 10.650 316.500 11.850 320.400 ;
        RECT 16.650 317.400 18.450 323.250 ;
        RECT 6.750 315.600 11.850 316.500 ;
        RECT 6.750 314.700 9.000 315.600 ;
        RECT 4.650 308.850 7.050 310.950 ;
        RECT 4.650 303.600 5.850 308.850 ;
        RECT 7.950 306.300 9.000 314.700 ;
        RECT 17.250 315.300 18.450 317.400 ;
        RECT 19.650 318.300 21.450 323.250 ;
        RECT 22.650 319.200 24.450 323.250 ;
        RECT 25.650 318.300 27.450 323.250 ;
        RECT 19.650 316.950 27.450 318.300 ;
        RECT 17.250 314.250 21.000 315.300 ;
        RECT 35.100 315.000 36.900 323.250 ;
        RECT 16.950 312.450 19.050 313.050 ;
        RECT 14.550 311.550 19.050 312.450 ;
        RECT 10.950 308.850 13.050 310.950 ;
        RECT 11.100 307.050 12.900 308.850 ;
        RECT 6.750 305.400 9.000 306.300 ;
        RECT 6.750 304.500 12.450 305.400 ;
        RECT 4.350 291.750 6.150 303.600 ;
        RECT 7.350 291.750 9.150 303.600 ;
        RECT 11.250 297.600 12.450 304.500 ;
        RECT 14.550 300.450 15.450 311.550 ;
        RECT 16.950 310.950 19.050 311.550 ;
        RECT 19.950 310.950 21.150 314.250 ;
        RECT 23.100 312.150 24.900 313.950 ;
        RECT 32.400 313.350 36.900 315.000 ;
        RECT 40.500 314.400 42.300 323.250 ;
        RECT 45.000 317.400 46.800 323.250 ;
        RECT 49.200 319.050 51.000 323.250 ;
        RECT 52.500 320.400 54.300 323.250 ;
        RECT 49.200 317.400 54.900 319.050 ;
        RECT 60.000 317.400 61.800 323.250 ;
        RECT 64.200 319.050 66.000 323.250 ;
        RECT 67.500 320.400 69.300 323.250 ;
        RECT 64.200 317.400 69.900 319.050 ;
        RECT 19.950 308.850 22.050 310.950 ;
        RECT 22.950 310.050 25.050 312.150 ;
        RECT 25.950 308.850 28.050 310.950 ;
        RECT 32.400 309.150 33.600 313.350 ;
        RECT 44.100 312.150 45.900 313.950 ;
        RECT 43.950 310.050 46.050 312.150 ;
        RECT 46.950 311.850 49.050 313.950 ;
        RECT 50.100 312.150 51.900 313.950 ;
        RECT 47.100 310.050 48.900 311.850 ;
        RECT 49.950 310.050 52.050 312.150 ;
        RECT 53.700 310.950 54.900 317.400 ;
        RECT 59.100 312.150 60.900 313.950 ;
        RECT 16.950 305.850 19.050 307.950 ;
        RECT 17.250 304.050 19.050 305.850 ;
        RECT 20.850 303.600 22.050 308.850 ;
        RECT 26.100 307.050 27.900 308.850 ;
        RECT 31.950 307.050 34.050 309.150 ;
        RECT 52.950 308.850 55.050 310.950 ;
        RECT 58.950 310.050 61.050 312.150 ;
        RECT 61.950 311.850 64.050 313.950 ;
        RECT 65.100 312.150 66.900 313.950 ;
        RECT 62.100 310.050 63.900 311.850 ;
        RECT 64.950 310.050 67.050 312.150 ;
        RECT 68.700 310.950 69.900 317.400 ;
        RECT 74.700 314.400 76.500 323.250 ;
        RECT 80.100 315.000 81.900 323.250 ;
        RECT 80.100 313.350 84.600 315.000 ;
        RECT 89.700 314.400 91.500 323.250 ;
        RECT 95.100 315.000 96.900 323.250 ;
        RECT 105.000 317.400 106.800 323.250 ;
        RECT 109.200 319.050 111.000 323.250 ;
        RECT 112.500 320.400 114.300 323.250 ;
        RECT 109.200 317.400 114.900 319.050 ;
        RECT 121.650 317.400 123.450 323.250 ;
        RECT 95.100 313.350 99.600 315.000 ;
        RECT 67.950 308.850 70.050 310.950 ;
        RECT 83.400 309.150 84.600 313.350 ;
        RECT 98.400 309.150 99.600 313.350 ;
        RECT 104.100 312.150 105.900 313.950 ;
        RECT 103.950 310.050 106.050 312.150 ;
        RECT 106.950 311.850 109.050 313.950 ;
        RECT 110.100 312.150 111.900 313.950 ;
        RECT 107.100 310.050 108.900 311.850 ;
        RECT 109.950 310.050 112.050 312.150 ;
        RECT 113.700 310.950 114.900 317.400 ;
        RECT 122.250 315.300 123.450 317.400 ;
        RECT 124.650 318.300 126.450 323.250 ;
        RECT 127.650 319.200 129.450 323.250 ;
        RECT 130.650 318.300 132.450 323.250 ;
        RECT 124.650 316.950 132.450 318.300 ;
        RECT 122.250 314.250 126.000 315.300 ;
        RECT 134.700 314.400 136.500 323.250 ;
        RECT 140.100 315.000 141.900 323.250 ;
        RECT 124.950 310.950 126.150 314.250 ;
        RECT 128.100 312.150 129.900 313.950 ;
        RECT 140.100 313.350 144.600 315.000 ;
        RECT 149.700 314.400 151.500 323.250 ;
        RECT 155.100 315.000 156.900 323.250 ;
        RECT 155.100 313.350 159.600 315.000 ;
        RECT 164.700 314.400 166.500 323.250 ;
        RECT 170.100 315.000 171.900 323.250 ;
        RECT 180.000 317.400 181.800 323.250 ;
        RECT 184.200 319.050 186.000 323.250 ;
        RECT 187.500 320.400 189.300 323.250 ;
        RECT 194.550 320.400 196.350 323.250 ;
        RECT 197.550 320.400 199.350 323.250 ;
        RECT 200.550 320.400 202.350 323.250 ;
        RECT 184.200 317.400 189.900 319.050 ;
        RECT 170.100 313.350 174.600 315.000 ;
        RECT 16.950 300.450 19.050 301.050 ;
        RECT 14.550 299.550 19.050 300.450 ;
        RECT 16.950 298.950 19.050 299.550 ;
        RECT 10.650 291.750 12.450 297.600 ;
        RECT 17.400 291.750 19.200 297.600 ;
        RECT 20.700 291.750 22.500 303.600 ;
        RECT 24.900 291.750 26.700 303.600 ;
        RECT 32.250 298.800 33.300 307.050 ;
        RECT 34.950 305.850 37.050 307.950 ;
        RECT 40.950 305.850 43.050 307.950 ;
        RECT 34.950 304.050 36.750 305.850 ;
        RECT 37.950 302.850 40.050 304.950 ;
        RECT 41.100 304.050 42.900 305.850 ;
        RECT 53.700 303.600 54.900 308.850 ;
        RECT 68.700 303.600 69.900 308.850 ;
        RECT 73.950 305.850 76.050 307.950 ;
        RECT 79.950 305.850 82.050 307.950 ;
        RECT 82.950 307.050 85.050 309.150 ;
        RECT 74.100 304.050 75.900 305.850 ;
        RECT 38.100 301.050 39.900 302.850 ;
        RECT 44.550 302.700 52.350 303.600 ;
        RECT 32.250 297.900 39.300 298.800 ;
        RECT 32.250 297.600 33.450 297.900 ;
        RECT 31.650 291.750 33.450 297.600 ;
        RECT 37.650 297.600 39.300 297.900 ;
        RECT 34.650 291.750 36.450 297.000 ;
        RECT 37.650 291.750 39.450 297.600 ;
        RECT 40.650 291.750 42.450 297.600 ;
        RECT 44.550 291.750 46.350 302.700 ;
        RECT 47.550 291.750 49.350 301.800 ;
        RECT 50.550 291.750 52.350 302.700 ;
        RECT 53.550 291.750 55.350 303.600 ;
        RECT 59.550 302.700 67.350 303.600 ;
        RECT 59.550 291.750 61.350 302.700 ;
        RECT 62.550 291.750 64.350 301.800 ;
        RECT 65.550 291.750 67.350 302.700 ;
        RECT 68.550 291.750 70.350 303.600 ;
        RECT 76.950 302.850 79.050 304.950 ;
        RECT 80.250 304.050 82.050 305.850 ;
        RECT 77.100 301.050 78.900 302.850 ;
        RECT 83.700 298.800 84.750 307.050 ;
        RECT 88.950 305.850 91.050 307.950 ;
        RECT 94.950 305.850 97.050 307.950 ;
        RECT 97.950 307.050 100.050 309.150 ;
        RECT 112.950 308.850 115.050 310.950 ;
        RECT 124.950 308.850 127.050 310.950 ;
        RECT 127.950 310.050 130.050 312.150 ;
        RECT 130.950 308.850 133.050 310.950 ;
        RECT 143.400 309.150 144.600 313.350 ;
        RECT 158.400 309.150 159.600 313.350 ;
        RECT 160.950 312.450 163.050 313.050 ;
        RECT 166.950 312.450 169.050 313.050 ;
        RECT 160.950 311.550 169.050 312.450 ;
        RECT 160.950 310.950 163.050 311.550 ;
        RECT 166.950 310.950 169.050 311.550 ;
        RECT 173.400 309.150 174.600 313.350 ;
        RECT 179.100 312.150 180.900 313.950 ;
        RECT 178.950 310.050 181.050 312.150 ;
        RECT 181.950 311.850 184.050 313.950 ;
        RECT 185.100 312.150 186.900 313.950 ;
        RECT 182.100 310.050 183.900 311.850 ;
        RECT 184.950 310.050 187.050 312.150 ;
        RECT 188.700 310.950 189.900 317.400 ;
        RECT 193.950 315.450 196.050 316.050 ;
        RECT 191.550 314.550 196.050 315.450 ;
        RECT 89.100 304.050 90.900 305.850 ;
        RECT 91.950 302.850 94.050 304.950 ;
        RECT 95.250 304.050 97.050 305.850 ;
        RECT 92.100 301.050 93.900 302.850 ;
        RECT 98.700 298.800 99.750 307.050 ;
        RECT 113.700 303.600 114.900 308.850 ;
        RECT 121.950 305.850 124.050 307.950 ;
        RECT 122.250 304.050 124.050 305.850 ;
        RECT 125.850 303.600 127.050 308.850 ;
        RECT 131.100 307.050 132.900 308.850 ;
        RECT 133.950 305.850 136.050 307.950 ;
        RECT 139.950 305.850 142.050 307.950 ;
        RECT 142.950 307.050 145.050 309.150 ;
        RECT 134.100 304.050 135.900 305.850 ;
        RECT 77.700 297.900 84.750 298.800 ;
        RECT 77.700 297.600 79.350 297.900 ;
        RECT 74.550 291.750 76.350 297.600 ;
        RECT 77.550 291.750 79.350 297.600 ;
        RECT 83.550 297.600 84.750 297.900 ;
        RECT 92.700 297.900 99.750 298.800 ;
        RECT 92.700 297.600 94.350 297.900 ;
        RECT 80.550 291.750 82.350 297.000 ;
        RECT 83.550 291.750 85.350 297.600 ;
        RECT 89.550 291.750 91.350 297.600 ;
        RECT 92.550 291.750 94.350 297.600 ;
        RECT 98.550 297.600 99.750 297.900 ;
        RECT 104.550 302.700 112.350 303.600 ;
        RECT 95.550 291.750 97.350 297.000 ;
        RECT 98.550 291.750 100.350 297.600 ;
        RECT 104.550 291.750 106.350 302.700 ;
        RECT 107.550 291.750 109.350 301.800 ;
        RECT 110.550 291.750 112.350 302.700 ;
        RECT 113.550 291.750 115.350 303.600 ;
        RECT 122.400 291.750 124.200 297.600 ;
        RECT 125.700 291.750 127.500 303.600 ;
        RECT 129.900 291.750 131.700 303.600 ;
        RECT 136.950 302.850 139.050 304.950 ;
        RECT 140.250 304.050 142.050 305.850 ;
        RECT 137.100 301.050 138.900 302.850 ;
        RECT 143.700 298.800 144.750 307.050 ;
        RECT 148.950 305.850 151.050 307.950 ;
        RECT 154.950 305.850 157.050 307.950 ;
        RECT 157.950 307.050 160.050 309.150 ;
        RECT 149.100 304.050 150.900 305.850 ;
        RECT 151.950 302.850 154.050 304.950 ;
        RECT 155.250 304.050 157.050 305.850 ;
        RECT 152.100 301.050 153.900 302.850 ;
        RECT 158.700 298.800 159.750 307.050 ;
        RECT 163.950 305.850 166.050 307.950 ;
        RECT 169.950 305.850 172.050 307.950 ;
        RECT 172.950 307.050 175.050 309.150 ;
        RECT 187.950 308.850 190.050 310.950 ;
        RECT 164.100 304.050 165.900 305.850 ;
        RECT 166.950 302.850 169.050 304.950 ;
        RECT 170.250 304.050 172.050 305.850 ;
        RECT 167.100 301.050 168.900 302.850 ;
        RECT 173.700 298.800 174.750 307.050 ;
        RECT 188.700 303.600 189.900 308.850 ;
        RECT 191.550 307.050 192.450 314.550 ;
        RECT 193.950 313.950 196.050 314.550 ;
        RECT 198.000 313.950 199.050 320.400 ;
        RECT 209.850 316.200 211.650 323.250 ;
        RECT 214.350 317.400 216.150 323.250 ;
        RECT 221.850 316.200 223.650 323.250 ;
        RECT 226.350 317.400 228.150 323.250 ;
        RECT 230.850 317.400 232.650 323.250 ;
        RECT 235.350 316.200 237.150 323.250 ;
        RECT 244.650 317.400 246.450 323.250 ;
        RECT 209.850 315.300 213.450 316.200 ;
        RECT 196.950 311.850 199.050 313.950 ;
        RECT 193.950 308.850 196.050 310.950 ;
        RECT 194.100 307.050 195.900 308.850 ;
        RECT 190.950 304.950 193.050 307.050 ;
        RECT 198.000 304.650 199.050 311.850 ;
        RECT 199.950 308.850 202.050 310.950 ;
        RECT 200.100 307.050 201.900 308.850 ;
        RECT 205.950 307.950 208.050 310.050 ;
        RECT 209.100 309.150 210.900 310.950 ;
        RECT 198.000 303.600 200.550 304.650 ;
        RECT 137.700 297.900 144.750 298.800 ;
        RECT 137.700 297.600 139.350 297.900 ;
        RECT 134.550 291.750 136.350 297.600 ;
        RECT 137.550 291.750 139.350 297.600 ;
        RECT 143.550 297.600 144.750 297.900 ;
        RECT 152.700 297.900 159.750 298.800 ;
        RECT 152.700 297.600 154.350 297.900 ;
        RECT 140.550 291.750 142.350 297.000 ;
        RECT 143.550 291.750 145.350 297.600 ;
        RECT 149.550 291.750 151.350 297.600 ;
        RECT 152.550 291.750 154.350 297.600 ;
        RECT 158.550 297.600 159.750 297.900 ;
        RECT 167.700 297.900 174.750 298.800 ;
        RECT 167.700 297.600 169.350 297.900 ;
        RECT 155.550 291.750 157.350 297.000 ;
        RECT 158.550 291.750 160.350 297.600 ;
        RECT 164.550 291.750 166.350 297.600 ;
        RECT 167.550 291.750 169.350 297.600 ;
        RECT 173.550 297.600 174.750 297.900 ;
        RECT 179.550 302.700 187.350 303.600 ;
        RECT 170.550 291.750 172.350 297.000 ;
        RECT 173.550 291.750 175.350 297.600 ;
        RECT 179.550 291.750 181.350 302.700 ;
        RECT 182.550 291.750 184.350 301.800 ;
        RECT 185.550 291.750 187.350 302.700 ;
        RECT 188.550 291.750 190.350 303.600 ;
        RECT 194.550 291.750 196.350 303.600 ;
        RECT 198.750 291.750 200.550 303.600 ;
        RECT 202.950 303.450 205.050 304.050 ;
        RECT 206.550 303.450 207.450 307.950 ;
        RECT 208.950 307.050 211.050 309.150 ;
        RECT 212.250 307.950 213.450 315.300 ;
        RECT 214.950 315.450 217.050 316.050 ;
        RECT 214.950 314.550 219.450 315.450 ;
        RECT 221.850 315.300 225.450 316.200 ;
        RECT 214.950 313.950 217.050 314.550 ;
        RECT 215.100 309.150 216.900 310.950 ;
        RECT 211.950 305.850 214.050 307.950 ;
        RECT 214.950 307.050 217.050 309.150 ;
        RECT 202.950 302.550 207.450 303.450 ;
        RECT 202.950 301.950 205.050 302.550 ;
        RECT 212.250 297.600 213.450 305.850 ;
        RECT 218.550 303.450 219.450 314.550 ;
        RECT 221.100 309.150 222.900 310.950 ;
        RECT 220.950 307.050 223.050 309.150 ;
        RECT 224.250 307.950 225.450 315.300 ;
        RECT 233.550 315.300 237.150 316.200 ;
        RECT 245.250 315.300 246.450 317.400 ;
        RECT 247.650 318.300 249.450 323.250 ;
        RECT 250.650 319.200 252.450 323.250 ;
        RECT 253.650 318.300 255.450 323.250 ;
        RECT 247.650 316.950 255.450 318.300 ;
        RECT 258.000 317.400 259.800 323.250 ;
        RECT 262.200 319.050 264.000 323.250 ;
        RECT 265.500 320.400 267.300 323.250 ;
        RECT 272.550 320.400 274.350 323.250 ;
        RECT 275.550 320.400 277.350 323.250 ;
        RECT 278.550 320.400 280.350 323.250 ;
        RECT 262.200 317.400 267.900 319.050 ;
        RECT 227.100 309.150 228.900 310.950 ;
        RECT 230.100 309.150 231.900 310.950 ;
        RECT 223.950 305.850 226.050 307.950 ;
        RECT 226.950 307.050 229.050 309.150 ;
        RECT 229.950 307.050 232.050 309.150 ;
        RECT 233.550 307.950 234.750 315.300 ;
        RECT 245.250 314.250 249.000 315.300 ;
        RECT 247.950 310.950 249.150 314.250 ;
        RECT 251.100 312.150 252.900 313.950 ;
        RECT 257.100 312.150 258.900 313.950 ;
        RECT 236.100 309.150 237.900 310.950 ;
        RECT 232.950 305.850 235.050 307.950 ;
        RECT 235.950 307.050 238.050 309.150 ;
        RECT 247.950 308.850 250.050 310.950 ;
        RECT 250.950 310.050 253.050 312.150 ;
        RECT 253.950 308.850 256.050 310.950 ;
        RECT 256.950 310.050 259.050 312.150 ;
        RECT 259.950 311.850 262.050 313.950 ;
        RECT 263.100 312.150 264.900 313.950 ;
        RECT 260.100 310.050 261.900 311.850 ;
        RECT 262.950 310.050 265.050 312.150 ;
        RECT 266.700 310.950 267.900 317.400 ;
        RECT 276.000 313.950 277.050 320.400 ;
        RECT 286.650 317.400 288.450 323.250 ;
        RECT 287.250 315.300 288.450 317.400 ;
        RECT 289.650 318.300 291.450 323.250 ;
        RECT 292.650 319.200 294.450 323.250 ;
        RECT 295.650 318.300 297.450 323.250 ;
        RECT 289.650 316.950 297.450 318.300 ;
        RECT 299.550 318.300 301.350 323.250 ;
        RECT 302.550 319.200 304.350 323.250 ;
        RECT 305.550 318.300 307.350 323.250 ;
        RECT 299.550 316.950 307.350 318.300 ;
        RECT 308.550 317.400 310.350 323.250 ;
        RECT 316.650 317.400 318.450 323.250 ;
        RECT 308.550 315.300 309.750 317.400 ;
        RECT 287.250 314.250 291.000 315.300 ;
        RECT 306.000 314.250 309.750 315.300 ;
        RECT 317.250 315.300 318.450 317.400 ;
        RECT 319.650 318.300 321.450 323.250 ;
        RECT 322.650 319.200 324.450 323.250 ;
        RECT 325.650 318.300 327.450 323.250 ;
        RECT 319.650 316.950 327.450 318.300 ;
        RECT 331.650 317.400 333.450 323.250 ;
        RECT 334.650 317.400 336.450 323.250 ;
        RECT 337.650 317.400 339.450 323.250 ;
        RECT 340.650 317.400 342.450 323.250 ;
        RECT 343.650 317.400 345.450 323.250 ;
        RECT 334.800 316.500 336.600 317.400 ;
        RECT 340.800 316.500 342.600 317.400 ;
        RECT 346.650 316.500 348.450 323.250 ;
        RECT 349.650 317.400 351.450 323.250 ;
        RECT 352.650 317.400 354.450 323.250 ;
        RECT 355.650 317.400 357.450 323.250 ;
        RECT 359.850 317.400 361.650 323.250 ;
        RECT 352.800 316.500 354.600 317.400 ;
        RECT 333.900 316.350 336.600 316.500 ;
        RECT 333.750 315.300 336.600 316.350 ;
        RECT 338.700 315.300 342.600 316.500 ;
        RECT 344.700 315.300 348.450 316.500 ;
        RECT 350.550 315.300 354.600 316.500 ;
        RECT 364.350 316.200 366.150 323.250 ;
        RECT 375.150 318.900 376.950 323.250 ;
        RECT 362.550 315.300 366.150 316.200 ;
        RECT 373.650 317.400 376.950 318.900 ;
        RECT 378.150 317.400 379.950 323.250 ;
        RECT 317.250 314.250 321.000 315.300 ;
        RECT 274.950 311.850 277.050 313.950 ;
        RECT 265.950 308.850 268.050 310.950 ;
        RECT 271.950 308.850 274.050 310.950 ;
        RECT 244.950 305.850 247.050 307.950 ;
        RECT 220.950 303.450 223.050 304.050 ;
        RECT 218.550 302.550 223.050 303.450 ;
        RECT 220.950 301.950 223.050 302.550 ;
        RECT 224.250 297.600 225.450 305.850 ;
        RECT 233.550 297.600 234.750 305.850 ;
        RECT 245.250 304.050 247.050 305.850 ;
        RECT 248.850 303.600 250.050 308.850 ;
        RECT 254.100 307.050 255.900 308.850 ;
        RECT 266.700 303.600 267.900 308.850 ;
        RECT 272.100 307.050 273.900 308.850 ;
        RECT 276.000 304.650 277.050 311.850 ;
        RECT 289.950 310.950 291.150 314.250 ;
        RECT 293.100 312.150 294.900 313.950 ;
        RECT 302.100 312.150 303.900 313.950 ;
        RECT 277.950 308.850 280.050 310.950 ;
        RECT 289.950 308.850 292.050 310.950 ;
        RECT 292.950 310.050 295.050 312.150 ;
        RECT 295.950 308.850 298.050 310.950 ;
        RECT 298.950 308.850 301.050 310.950 ;
        RECT 301.950 310.050 304.050 312.150 ;
        RECT 305.850 310.950 307.050 314.250 ;
        RECT 304.950 308.850 307.050 310.950 ;
        RECT 319.950 310.950 321.150 314.250 ;
        RECT 323.100 312.150 324.900 313.950 ;
        RECT 333.750 312.150 334.800 315.300 ;
        RECT 338.700 314.400 339.900 315.300 ;
        RECT 344.700 314.400 345.900 315.300 ;
        RECT 350.550 314.400 351.750 315.300 ;
        RECT 335.700 312.600 339.900 314.400 ;
        RECT 341.700 312.600 345.900 314.400 ;
        RECT 347.700 312.600 351.750 314.400 ;
        RECT 319.950 308.850 322.050 310.950 ;
        RECT 322.950 310.050 325.050 312.150 ;
        RECT 325.950 308.850 328.050 310.950 ;
        RECT 331.950 310.050 334.800 312.150 ;
        RECT 278.100 307.050 279.900 308.850 ;
        RECT 286.950 305.850 289.050 307.950 ;
        RECT 276.000 303.600 278.550 304.650 ;
        RECT 287.250 304.050 289.050 305.850 ;
        RECT 290.850 303.600 292.050 308.850 ;
        RECT 296.100 307.050 297.900 308.850 ;
        RECT 299.100 307.050 300.900 308.850 ;
        RECT 304.950 303.600 306.150 308.850 ;
        RECT 307.950 305.850 310.050 307.950 ;
        RECT 316.950 305.850 319.050 307.950 ;
        RECT 307.950 304.050 309.750 305.850 ;
        RECT 317.250 304.050 319.050 305.850 ;
        RECT 320.850 303.600 322.050 308.850 ;
        RECT 326.100 307.050 327.900 308.850 ;
        RECT 333.750 305.700 334.800 310.050 ;
        RECT 338.700 305.700 339.900 312.600 ;
        RECT 344.700 305.700 345.900 312.600 ;
        RECT 350.550 305.700 351.750 312.600 ;
        RECT 353.100 312.150 354.900 313.950 ;
        RECT 352.950 310.050 355.050 312.150 ;
        RECT 359.100 309.150 360.900 310.950 ;
        RECT 358.950 307.050 361.050 309.150 ;
        RECT 362.550 307.950 363.750 315.300 ;
        RECT 373.650 310.950 374.850 317.400 ;
        RECT 376.950 315.900 378.750 316.500 ;
        RECT 382.650 315.900 384.450 323.250 ;
        RECT 386.550 320.400 388.350 323.250 ;
        RECT 389.550 320.400 391.350 323.250 ;
        RECT 392.550 320.400 394.350 323.250 ;
        RECT 376.950 314.700 384.450 315.900 ;
        RECT 390.450 316.200 391.350 320.400 ;
        RECT 395.550 317.400 397.350 323.250 ;
        RECT 390.450 315.300 393.750 316.200 ;
        RECT 365.100 309.150 366.900 310.950 ;
        RECT 361.950 305.850 364.050 307.950 ;
        RECT 364.950 307.050 367.050 309.150 ;
        RECT 373.650 308.850 376.050 310.950 ;
        RECT 377.100 309.150 378.900 310.950 ;
        RECT 333.750 304.500 336.450 305.700 ;
        RECT 338.700 304.500 342.450 305.700 ;
        RECT 344.700 304.500 348.450 305.700 ;
        RECT 350.550 304.500 354.450 305.700 ;
        RECT 208.650 291.750 210.450 297.600 ;
        RECT 211.650 291.750 213.450 297.600 ;
        RECT 214.650 291.750 216.450 297.600 ;
        RECT 220.650 291.750 222.450 297.600 ;
        RECT 223.650 291.750 225.450 297.600 ;
        RECT 226.650 291.750 228.450 297.600 ;
        RECT 230.550 291.750 232.350 297.600 ;
        RECT 233.550 291.750 235.350 297.600 ;
        RECT 236.550 291.750 238.350 297.600 ;
        RECT 245.400 291.750 247.200 297.600 ;
        RECT 248.700 291.750 250.500 303.600 ;
        RECT 252.900 291.750 254.700 303.600 ;
        RECT 257.550 302.700 265.350 303.600 ;
        RECT 257.550 291.750 259.350 302.700 ;
        RECT 260.550 291.750 262.350 301.800 ;
        RECT 263.550 291.750 265.350 302.700 ;
        RECT 266.550 291.750 268.350 303.600 ;
        RECT 272.550 291.750 274.350 303.600 ;
        RECT 276.750 291.750 278.550 303.600 ;
        RECT 287.400 291.750 289.200 297.600 ;
        RECT 290.700 291.750 292.500 303.600 ;
        RECT 294.900 291.750 296.700 303.600 ;
        RECT 300.300 291.750 302.100 303.600 ;
        RECT 304.500 291.750 306.300 303.600 ;
        RECT 307.800 291.750 309.600 297.600 ;
        RECT 317.400 291.750 319.200 297.600 ;
        RECT 320.700 291.750 322.500 303.600 ;
        RECT 324.900 291.750 326.700 303.600 ;
        RECT 331.650 291.750 333.450 303.600 ;
        RECT 334.650 291.750 336.450 304.500 ;
        RECT 337.650 291.750 339.450 303.600 ;
        RECT 340.650 291.750 342.450 304.500 ;
        RECT 343.650 291.750 345.450 303.600 ;
        RECT 346.650 291.750 348.450 304.500 ;
        RECT 349.650 291.750 351.450 303.600 ;
        RECT 352.650 291.750 354.450 304.500 ;
        RECT 355.650 291.750 357.450 303.600 ;
        RECT 362.550 297.600 363.750 305.850 ;
        RECT 373.650 303.600 374.850 308.850 ;
        RECT 376.950 307.050 379.050 309.150 ;
        RECT 359.550 291.750 361.350 297.600 ;
        RECT 362.550 291.750 364.350 297.600 ;
        RECT 365.550 291.750 367.350 297.600 ;
        RECT 373.050 291.750 374.850 303.600 ;
        RECT 376.050 291.750 377.850 303.600 ;
        RECT 380.100 297.600 381.300 314.700 ;
        RECT 391.950 314.400 393.750 315.300 ;
        RECT 385.950 311.850 388.050 313.950 ;
        RECT 382.950 308.850 385.050 310.950 ;
        RECT 386.100 310.050 387.900 311.850 ;
        RECT 388.950 308.850 391.050 310.950 ;
        RECT 383.100 307.050 384.900 308.850 ;
        RECT 389.100 307.050 390.900 308.850 ;
        RECT 392.700 306.150 393.600 314.400 ;
        RECT 396.000 312.150 397.050 317.400 ;
        RECT 404.850 316.200 406.650 323.250 ;
        RECT 409.350 317.400 411.150 323.250 ;
        RECT 413.850 317.400 415.650 323.250 ;
        RECT 418.350 316.200 420.150 323.250 ;
        RECT 404.850 315.300 408.450 316.200 ;
        RECT 394.950 310.050 397.050 312.150 ;
        RECT 391.950 306.000 393.750 306.150 ;
        RECT 386.550 304.800 393.750 306.000 ;
        RECT 386.550 303.600 387.750 304.800 ;
        RECT 391.950 304.350 393.750 304.800 ;
        RECT 379.650 291.750 381.450 297.600 ;
        RECT 382.650 291.750 384.450 297.600 ;
        RECT 386.550 291.750 388.350 303.600 ;
        RECT 395.100 303.450 396.450 310.050 ;
        RECT 404.100 309.150 405.900 310.950 ;
        RECT 403.950 307.050 406.050 309.150 ;
        RECT 407.250 307.950 408.450 315.300 ;
        RECT 416.550 315.300 420.150 316.200 ;
        RECT 426.150 317.400 427.950 323.250 ;
        RECT 429.150 320.400 430.950 323.250 ;
        RECT 433.950 321.300 435.750 323.250 ;
        RECT 432.000 320.400 435.750 321.300 ;
        RECT 438.450 320.400 440.250 323.250 ;
        RECT 441.750 320.400 443.550 323.250 ;
        RECT 445.650 320.400 447.450 323.250 ;
        RECT 449.850 320.400 451.650 323.250 ;
        RECT 454.350 320.400 456.150 323.250 ;
        RECT 432.000 319.500 433.050 320.400 ;
        RECT 430.950 317.400 433.050 319.500 ;
        RECT 441.750 318.600 442.800 320.400 ;
        RECT 410.100 309.150 411.900 310.950 ;
        RECT 413.100 309.150 414.900 310.950 ;
        RECT 406.950 305.850 409.050 307.950 ;
        RECT 409.950 307.050 412.050 309.150 ;
        RECT 412.950 307.050 415.050 309.150 ;
        RECT 416.550 307.950 417.750 315.300 ;
        RECT 419.100 309.150 420.900 310.950 ;
        RECT 415.950 305.850 418.050 307.950 ;
        RECT 418.950 307.050 421.050 309.150 ;
        RECT 391.050 291.750 392.850 303.450 ;
        RECT 394.050 302.100 396.450 303.450 ;
        RECT 394.050 291.750 395.850 302.100 ;
        RECT 407.250 297.600 408.450 305.850 ;
        RECT 416.550 297.600 417.750 305.850 ;
        RECT 426.150 304.800 427.050 317.400 ;
        RECT 434.550 316.800 436.350 318.600 ;
        RECT 437.850 317.550 442.800 318.600 ;
        RECT 450.300 319.500 451.350 320.400 ;
        RECT 450.300 318.300 454.050 319.500 ;
        RECT 437.850 316.800 439.650 317.550 ;
        RECT 434.850 315.900 435.900 316.800 ;
        RECT 445.050 316.200 446.850 318.000 ;
        RECT 451.950 317.400 454.050 318.300 ;
        RECT 457.650 317.400 459.450 323.250 ;
        RECT 464.700 320.400 466.500 323.250 ;
        RECT 468.000 319.050 469.800 323.250 ;
        RECT 445.050 315.900 445.950 316.200 ;
        RECT 434.850 315.000 445.950 315.900 ;
        RECT 458.250 315.150 459.450 317.400 ;
        RECT 434.850 313.800 435.900 315.000 ;
        RECT 429.000 312.600 435.900 313.800 ;
        RECT 429.000 311.850 429.900 312.600 ;
        RECT 434.100 312.000 435.900 312.600 ;
        RECT 428.100 310.050 429.900 311.850 ;
        RECT 431.100 310.950 432.900 311.700 ;
        RECT 445.050 310.950 445.950 315.000 ;
        RECT 454.950 313.050 459.450 315.150 ;
        RECT 453.150 311.250 457.050 313.050 ;
        RECT 454.950 310.950 457.050 311.250 ;
        RECT 431.100 309.900 439.050 310.950 ;
        RECT 436.950 308.850 439.050 309.900 ;
        RECT 442.950 308.850 445.950 310.950 ;
        RECT 435.450 305.100 437.250 305.400 ;
        RECT 435.450 304.800 443.850 305.100 ;
        RECT 426.150 304.200 443.850 304.800 ;
        RECT 426.150 303.600 437.250 304.200 ;
        RECT 403.650 291.750 405.450 297.600 ;
        RECT 406.650 291.750 408.450 297.600 ;
        RECT 409.650 291.750 411.450 297.600 ;
        RECT 413.550 291.750 415.350 297.600 ;
        RECT 416.550 291.750 418.350 297.600 ;
        RECT 419.550 291.750 421.350 297.600 ;
        RECT 426.150 291.750 427.950 303.600 ;
        RECT 440.250 302.700 442.050 303.300 ;
        RECT 434.550 301.500 442.050 302.700 ;
        RECT 442.950 302.100 443.850 304.200 ;
        RECT 445.050 304.200 445.950 308.850 ;
        RECT 455.250 305.400 457.050 307.200 ;
        RECT 451.950 304.200 456.150 305.400 ;
        RECT 445.050 303.300 451.050 304.200 ;
        RECT 451.950 303.300 454.050 304.200 ;
        RECT 458.250 303.600 459.450 313.050 ;
        RECT 464.100 317.400 469.800 319.050 ;
        RECT 472.200 317.400 474.000 323.250 ;
        RECT 476.550 320.400 478.350 323.250 ;
        RECT 479.550 320.400 481.350 323.250 ;
        RECT 482.550 320.400 484.350 323.250 ;
        RECT 464.100 310.950 465.300 317.400 ;
        RECT 480.000 313.950 481.050 320.400 ;
        RECT 493.800 317.400 495.600 323.250 ;
        RECT 498.000 317.400 499.800 323.250 ;
        RECT 502.200 317.400 504.000 323.250 ;
        RECT 507.150 317.400 508.950 323.250 ;
        RECT 510.150 320.400 511.950 323.250 ;
        RECT 514.950 321.300 516.750 323.250 ;
        RECT 513.000 320.400 516.750 321.300 ;
        RECT 519.450 320.400 521.250 323.250 ;
        RECT 522.750 320.400 524.550 323.250 ;
        RECT 526.650 320.400 528.450 323.250 ;
        RECT 530.850 320.400 532.650 323.250 ;
        RECT 535.350 320.400 537.150 323.250 ;
        RECT 513.000 319.500 514.050 320.400 ;
        RECT 511.950 317.400 514.050 319.500 ;
        RECT 522.750 318.600 523.800 320.400 ;
        RECT 467.100 312.150 468.900 313.950 ;
        RECT 463.950 308.850 466.050 310.950 ;
        RECT 466.950 310.050 469.050 312.150 ;
        RECT 469.950 311.850 472.050 313.950 ;
        RECT 473.100 312.150 474.900 313.950 ;
        RECT 470.100 310.050 471.900 311.850 ;
        RECT 472.950 310.050 475.050 312.150 ;
        RECT 478.950 311.850 481.050 313.950 ;
        RECT 494.250 312.150 496.050 313.950 ;
        RECT 475.950 308.850 478.050 310.950 ;
        RECT 464.100 303.600 465.300 308.850 ;
        RECT 476.100 307.050 477.900 308.850 ;
        RECT 480.000 304.650 481.050 311.850 ;
        RECT 481.950 308.850 484.050 310.950 ;
        RECT 490.950 308.850 493.050 310.950 ;
        RECT 493.950 310.050 496.050 312.150 ;
        RECT 498.000 310.950 499.050 317.400 ;
        RECT 496.950 308.850 499.050 310.950 ;
        RECT 499.950 312.150 501.750 313.950 ;
        RECT 499.950 310.050 502.050 312.150 ;
        RECT 502.950 308.850 505.050 310.950 ;
        RECT 482.100 307.050 483.900 308.850 ;
        RECT 491.100 307.050 492.900 308.850 ;
        RECT 496.950 305.400 497.850 308.850 ;
        RECT 502.950 307.050 504.750 308.850 ;
        RECT 480.000 303.600 482.550 304.650 ;
        RECT 493.800 304.500 497.850 305.400 ;
        RECT 507.150 304.800 508.050 317.400 ;
        RECT 515.550 316.800 517.350 318.600 ;
        RECT 518.850 317.550 523.800 318.600 ;
        RECT 531.300 319.500 532.350 320.400 ;
        RECT 531.300 318.300 535.050 319.500 ;
        RECT 518.850 316.800 520.650 317.550 ;
        RECT 515.850 315.900 516.900 316.800 ;
        RECT 526.050 316.200 527.850 318.000 ;
        RECT 532.950 317.400 535.050 318.300 ;
        RECT 538.650 317.400 540.450 323.250 ;
        RECT 526.050 315.900 526.950 316.200 ;
        RECT 515.850 315.000 526.950 315.900 ;
        RECT 539.250 315.150 540.450 317.400 ;
        RECT 542.550 318.300 544.350 323.250 ;
        RECT 545.550 319.200 547.350 323.250 ;
        RECT 548.550 318.300 550.350 323.250 ;
        RECT 542.550 316.950 550.350 318.300 ;
        RECT 551.550 317.400 553.350 323.250 ;
        RECT 558.150 317.400 559.950 323.250 ;
        RECT 561.150 320.400 562.950 323.250 ;
        RECT 565.950 321.300 567.750 323.250 ;
        RECT 564.000 320.400 567.750 321.300 ;
        RECT 570.450 320.400 572.250 323.250 ;
        RECT 573.750 320.400 575.550 323.250 ;
        RECT 577.650 320.400 579.450 323.250 ;
        RECT 581.850 320.400 583.650 323.250 ;
        RECT 586.350 320.400 588.150 323.250 ;
        RECT 564.000 319.500 565.050 320.400 ;
        RECT 562.950 317.400 565.050 319.500 ;
        RECT 573.750 318.600 574.800 320.400 ;
        RECT 551.550 315.300 552.750 317.400 ;
        RECT 515.850 313.800 516.900 315.000 ;
        RECT 510.000 312.600 516.900 313.800 ;
        RECT 510.000 311.850 510.900 312.600 ;
        RECT 515.100 312.000 516.900 312.600 ;
        RECT 509.100 310.050 510.900 311.850 ;
        RECT 512.100 310.950 513.900 311.700 ;
        RECT 526.050 310.950 526.950 315.000 ;
        RECT 535.950 313.050 540.450 315.150 ;
        RECT 549.000 314.250 552.750 315.300 ;
        RECT 534.150 311.250 538.050 313.050 ;
        RECT 535.950 310.950 538.050 311.250 ;
        RECT 512.100 309.900 520.050 310.950 ;
        RECT 517.950 308.850 520.050 309.900 ;
        RECT 523.950 308.850 526.950 310.950 ;
        RECT 516.450 305.100 518.250 305.400 ;
        RECT 516.450 304.800 524.850 305.100 ;
        RECT 493.800 303.600 495.600 304.500 ;
        RECT 507.150 304.200 524.850 304.800 ;
        RECT 507.150 303.600 518.250 304.200 ;
        RECT 450.150 302.400 451.050 303.300 ;
        RECT 447.450 302.100 449.250 302.400 ;
        RECT 434.550 300.600 435.750 301.500 ;
        RECT 442.950 301.200 449.250 302.100 ;
        RECT 447.450 300.600 449.250 301.200 ;
        RECT 450.150 300.600 452.850 302.400 ;
        RECT 430.950 298.500 435.750 300.600 ;
        RECT 438.150 298.500 445.050 300.300 ;
        RECT 434.550 297.600 435.750 298.500 ;
        RECT 429.150 291.750 430.950 297.600 ;
        RECT 434.250 291.750 436.050 297.600 ;
        RECT 439.050 291.750 440.850 297.600 ;
        RECT 442.050 291.750 443.850 298.500 ;
        RECT 450.150 297.600 454.050 299.700 ;
        RECT 445.950 291.750 447.750 297.600 ;
        RECT 450.150 291.750 451.950 297.600 ;
        RECT 454.650 291.750 456.450 294.600 ;
        RECT 457.650 291.750 459.450 303.600 ;
        RECT 463.650 291.750 465.450 303.600 ;
        RECT 466.650 302.700 474.450 303.600 ;
        RECT 466.650 291.750 468.450 302.700 ;
        RECT 469.650 291.750 471.450 301.800 ;
        RECT 472.650 291.750 474.450 302.700 ;
        RECT 476.550 291.750 478.350 303.600 ;
        RECT 480.750 291.750 482.550 303.600 ;
        RECT 490.650 292.500 492.450 303.600 ;
        RECT 493.650 293.400 495.450 303.600 ;
        RECT 496.650 302.400 504.450 303.300 ;
        RECT 496.650 292.500 498.450 302.400 ;
        RECT 490.650 291.750 498.450 292.500 ;
        RECT 499.650 291.750 501.450 301.500 ;
        RECT 502.650 291.750 504.450 302.400 ;
        RECT 507.150 291.750 508.950 303.600 ;
        RECT 521.250 302.700 523.050 303.300 ;
        RECT 515.550 301.500 523.050 302.700 ;
        RECT 523.950 302.100 524.850 304.200 ;
        RECT 526.050 304.200 526.950 308.850 ;
        RECT 536.250 305.400 538.050 307.200 ;
        RECT 532.950 304.200 537.150 305.400 ;
        RECT 526.050 303.300 532.050 304.200 ;
        RECT 532.950 303.300 535.050 304.200 ;
        RECT 539.250 303.600 540.450 313.050 ;
        RECT 545.100 312.150 546.900 313.950 ;
        RECT 541.950 308.850 544.050 310.950 ;
        RECT 544.950 310.050 547.050 312.150 ;
        RECT 548.850 310.950 550.050 314.250 ;
        RECT 547.950 308.850 550.050 310.950 ;
        RECT 542.100 307.050 543.900 308.850 ;
        RECT 547.950 303.600 549.150 308.850 ;
        RECT 550.950 305.850 553.050 307.950 ;
        RECT 550.950 304.050 552.750 305.850 ;
        RECT 558.150 304.800 559.050 317.400 ;
        RECT 566.550 316.800 568.350 318.600 ;
        RECT 569.850 317.550 574.800 318.600 ;
        RECT 582.300 319.500 583.350 320.400 ;
        RECT 582.300 318.300 586.050 319.500 ;
        RECT 569.850 316.800 571.650 317.550 ;
        RECT 566.850 315.900 567.900 316.800 ;
        RECT 577.050 316.200 578.850 318.000 ;
        RECT 583.950 317.400 586.050 318.300 ;
        RECT 589.650 317.400 591.450 323.250 ;
        RECT 577.050 315.900 577.950 316.200 ;
        RECT 566.850 315.000 577.950 315.900 ;
        RECT 590.250 315.150 591.450 317.400 ;
        RECT 566.850 313.800 567.900 315.000 ;
        RECT 561.000 312.600 567.900 313.800 ;
        RECT 561.000 311.850 561.900 312.600 ;
        RECT 566.100 312.000 567.900 312.600 ;
        RECT 560.100 310.050 561.900 311.850 ;
        RECT 563.100 310.950 564.900 311.700 ;
        RECT 577.050 310.950 577.950 315.000 ;
        RECT 586.950 313.050 591.450 315.150 ;
        RECT 585.150 311.250 589.050 313.050 ;
        RECT 586.950 310.950 589.050 311.250 ;
        RECT 563.100 309.900 571.050 310.950 ;
        RECT 568.950 308.850 571.050 309.900 ;
        RECT 574.950 308.850 577.950 310.950 ;
        RECT 567.450 305.100 569.250 305.400 ;
        RECT 567.450 304.800 575.850 305.100 ;
        RECT 558.150 304.200 575.850 304.800 ;
        RECT 558.150 303.600 569.250 304.200 ;
        RECT 531.150 302.400 532.050 303.300 ;
        RECT 528.450 302.100 530.250 302.400 ;
        RECT 515.550 300.600 516.750 301.500 ;
        RECT 523.950 301.200 530.250 302.100 ;
        RECT 528.450 300.600 530.250 301.200 ;
        RECT 531.150 300.600 533.850 302.400 ;
        RECT 511.950 298.500 516.750 300.600 ;
        RECT 519.150 298.500 526.050 300.300 ;
        RECT 515.550 297.600 516.750 298.500 ;
        RECT 510.150 291.750 511.950 297.600 ;
        RECT 515.250 291.750 517.050 297.600 ;
        RECT 520.050 291.750 521.850 297.600 ;
        RECT 523.050 291.750 524.850 298.500 ;
        RECT 531.150 297.600 535.050 299.700 ;
        RECT 526.950 291.750 528.750 297.600 ;
        RECT 531.150 291.750 532.950 297.600 ;
        RECT 535.650 291.750 537.450 294.600 ;
        RECT 538.650 291.750 540.450 303.600 ;
        RECT 543.300 291.750 545.100 303.600 ;
        RECT 547.500 291.750 549.300 303.600 ;
        RECT 550.800 291.750 552.600 297.600 ;
        RECT 558.150 291.750 559.950 303.600 ;
        RECT 572.250 302.700 574.050 303.300 ;
        RECT 566.550 301.500 574.050 302.700 ;
        RECT 574.950 302.100 575.850 304.200 ;
        RECT 577.050 304.200 577.950 308.850 ;
        RECT 587.250 305.400 589.050 307.200 ;
        RECT 583.950 304.200 588.150 305.400 ;
        RECT 577.050 303.300 583.050 304.200 ;
        RECT 583.950 303.300 586.050 304.200 ;
        RECT 590.250 303.600 591.450 313.050 ;
        RECT 582.150 302.400 583.050 303.300 ;
        RECT 579.450 302.100 581.250 302.400 ;
        RECT 566.550 300.600 567.750 301.500 ;
        RECT 574.950 301.200 581.250 302.100 ;
        RECT 579.450 300.600 581.250 301.200 ;
        RECT 582.150 300.600 584.850 302.400 ;
        RECT 562.950 298.500 567.750 300.600 ;
        RECT 570.150 298.500 577.050 300.300 ;
        RECT 566.550 297.600 567.750 298.500 ;
        RECT 561.150 291.750 562.950 297.600 ;
        RECT 566.250 291.750 568.050 297.600 ;
        RECT 571.050 291.750 572.850 297.600 ;
        RECT 574.050 291.750 575.850 298.500 ;
        RECT 582.150 297.600 586.050 299.700 ;
        RECT 577.950 291.750 579.750 297.600 ;
        RECT 582.150 291.750 583.950 297.600 ;
        RECT 586.650 291.750 588.450 294.600 ;
        RECT 589.650 291.750 591.450 303.600 ;
        RECT 593.550 317.400 595.350 323.250 ;
        RECT 596.850 320.400 598.650 323.250 ;
        RECT 601.350 320.400 603.150 323.250 ;
        RECT 605.550 320.400 607.350 323.250 ;
        RECT 609.450 320.400 611.250 323.250 ;
        RECT 612.750 320.400 614.550 323.250 ;
        RECT 617.250 321.300 619.050 323.250 ;
        RECT 617.250 320.400 621.000 321.300 ;
        RECT 622.050 320.400 623.850 323.250 ;
        RECT 601.650 319.500 602.700 320.400 ;
        RECT 598.950 318.300 602.700 319.500 ;
        RECT 610.200 318.600 611.250 320.400 ;
        RECT 619.950 319.500 621.000 320.400 ;
        RECT 598.950 317.400 601.050 318.300 ;
        RECT 593.550 315.150 594.750 317.400 ;
        RECT 606.150 316.200 607.950 318.000 ;
        RECT 610.200 317.550 615.150 318.600 ;
        RECT 613.350 316.800 615.150 317.550 ;
        RECT 616.650 316.800 618.450 318.600 ;
        RECT 619.950 317.400 622.050 319.500 ;
        RECT 625.050 317.400 626.850 323.250 ;
        RECT 634.800 317.400 636.600 323.250 ;
        RECT 639.000 317.400 640.800 323.250 ;
        RECT 643.200 317.400 645.000 323.250 ;
        RECT 647.550 320.400 649.350 323.250 ;
        RECT 650.550 320.400 652.350 323.250 ;
        RECT 658.650 320.400 660.450 323.250 ;
        RECT 661.650 320.400 663.450 323.250 ;
        RECT 664.650 320.400 666.450 323.250 ;
        RECT 670.650 320.400 672.450 323.250 ;
        RECT 673.650 320.400 675.450 323.250 ;
        RECT 676.650 320.400 678.450 323.250 ;
        RECT 607.050 315.900 607.950 316.200 ;
        RECT 617.100 315.900 618.150 316.800 ;
        RECT 593.550 313.050 598.050 315.150 ;
        RECT 607.050 315.000 618.150 315.900 ;
        RECT 593.550 303.600 594.750 313.050 ;
        RECT 595.950 311.250 599.850 313.050 ;
        RECT 595.950 310.950 598.050 311.250 ;
        RECT 607.050 310.950 607.950 315.000 ;
        RECT 617.100 313.800 618.150 315.000 ;
        RECT 617.100 312.600 624.000 313.800 ;
        RECT 617.100 312.000 618.900 312.600 ;
        RECT 623.100 311.850 624.000 312.600 ;
        RECT 620.100 310.950 621.900 311.700 ;
        RECT 607.050 308.850 610.050 310.950 ;
        RECT 613.950 309.900 621.900 310.950 ;
        RECT 623.100 310.050 624.900 311.850 ;
        RECT 613.950 308.850 616.050 309.900 ;
        RECT 595.950 305.400 597.750 307.200 ;
        RECT 596.850 304.200 601.050 305.400 ;
        RECT 607.050 304.200 607.950 308.850 ;
        RECT 615.750 305.100 617.550 305.400 ;
        RECT 593.550 291.750 595.350 303.600 ;
        RECT 598.950 303.300 601.050 304.200 ;
        RECT 601.950 303.300 607.950 304.200 ;
        RECT 609.150 304.800 617.550 305.100 ;
        RECT 625.950 304.800 626.850 317.400 ;
        RECT 635.250 312.150 637.050 313.950 ;
        RECT 631.950 308.850 634.050 310.950 ;
        RECT 634.950 310.050 637.050 312.150 ;
        RECT 639.000 310.950 640.050 317.400 ;
        RECT 637.950 308.850 640.050 310.950 ;
        RECT 640.950 312.150 642.750 313.950 ;
        RECT 640.950 310.050 643.050 312.150 ;
        RECT 646.950 311.850 649.050 313.950 ;
        RECT 650.400 312.150 651.600 320.400 ;
        RECT 661.950 313.950 663.000 320.400 ;
        RECT 673.950 313.950 675.000 320.400 ;
        RECT 680.550 317.400 682.350 323.250 ;
        RECT 683.850 320.400 685.650 323.250 ;
        RECT 688.350 320.400 690.150 323.250 ;
        RECT 692.550 320.400 694.350 323.250 ;
        RECT 696.450 320.400 698.250 323.250 ;
        RECT 699.750 320.400 701.550 323.250 ;
        RECT 704.250 321.300 706.050 323.250 ;
        RECT 704.250 320.400 708.000 321.300 ;
        RECT 709.050 320.400 710.850 323.250 ;
        RECT 688.650 319.500 689.700 320.400 ;
        RECT 685.950 318.300 689.700 319.500 ;
        RECT 697.200 318.600 698.250 320.400 ;
        RECT 706.950 319.500 708.000 320.400 ;
        RECT 685.950 317.400 688.050 318.300 ;
        RECT 680.550 315.150 681.750 317.400 ;
        RECT 693.150 316.200 694.950 318.000 ;
        RECT 697.200 317.550 702.150 318.600 ;
        RECT 700.350 316.800 702.150 317.550 ;
        RECT 703.650 316.800 705.450 318.600 ;
        RECT 706.950 317.400 709.050 319.500 ;
        RECT 712.050 317.400 713.850 323.250 ;
        RECT 694.050 315.900 694.950 316.200 ;
        RECT 704.100 315.900 705.150 316.800 ;
        RECT 643.950 308.850 646.050 310.950 ;
        RECT 647.100 310.050 648.900 311.850 ;
        RECT 649.950 310.050 652.050 312.150 ;
        RECT 661.950 311.850 664.050 313.950 ;
        RECT 673.950 311.850 676.050 313.950 ;
        RECT 680.550 313.050 685.050 315.150 ;
        RECT 694.050 315.000 705.150 315.900 ;
        RECT 632.100 307.050 633.900 308.850 ;
        RECT 637.950 305.400 638.850 308.850 ;
        RECT 643.950 307.050 645.750 308.850 ;
        RECT 609.150 304.200 626.850 304.800 ;
        RECT 601.950 302.400 602.850 303.300 ;
        RECT 600.150 300.600 602.850 302.400 ;
        RECT 603.750 302.100 605.550 302.400 ;
        RECT 609.150 302.100 610.050 304.200 ;
        RECT 615.750 303.600 626.850 304.200 ;
        RECT 634.800 304.500 638.850 305.400 ;
        RECT 634.800 303.600 636.600 304.500 ;
        RECT 603.750 301.200 610.050 302.100 ;
        RECT 610.950 302.700 612.750 303.300 ;
        RECT 610.950 301.500 618.450 302.700 ;
        RECT 603.750 300.600 605.550 301.200 ;
        RECT 617.250 300.600 618.450 301.500 ;
        RECT 598.950 297.600 602.850 299.700 ;
        RECT 607.950 298.500 614.850 300.300 ;
        RECT 617.250 298.500 622.050 300.600 ;
        RECT 596.550 291.750 598.350 294.600 ;
        RECT 601.050 291.750 602.850 297.600 ;
        RECT 605.250 291.750 607.050 297.600 ;
        RECT 609.150 291.750 610.950 298.500 ;
        RECT 617.250 297.600 618.450 298.500 ;
        RECT 612.150 291.750 613.950 297.600 ;
        RECT 616.950 291.750 618.750 297.600 ;
        RECT 622.050 291.750 623.850 297.600 ;
        RECT 625.050 291.750 626.850 303.600 ;
        RECT 631.650 292.500 633.450 303.600 ;
        RECT 634.650 293.400 636.450 303.600 ;
        RECT 637.650 302.400 645.450 303.300 ;
        RECT 637.650 292.500 639.450 302.400 ;
        RECT 631.650 291.750 639.450 292.500 ;
        RECT 640.650 291.750 642.450 301.500 ;
        RECT 643.650 291.750 645.450 302.400 ;
        RECT 650.400 297.600 651.600 310.050 ;
        RECT 658.950 308.850 661.050 310.950 ;
        RECT 659.100 307.050 660.900 308.850 ;
        RECT 661.950 304.650 663.000 311.850 ;
        RECT 664.950 308.850 667.050 310.950 ;
        RECT 670.950 308.850 673.050 310.950 ;
        RECT 665.100 307.050 666.900 308.850 ;
        RECT 671.100 307.050 672.900 308.850 ;
        RECT 673.950 304.650 675.000 311.850 ;
        RECT 676.950 308.850 679.050 310.950 ;
        RECT 677.100 307.050 678.900 308.850 ;
        RECT 660.450 303.600 663.000 304.650 ;
        RECT 672.450 303.600 675.000 304.650 ;
        RECT 680.550 303.600 681.750 313.050 ;
        RECT 682.950 311.250 686.850 313.050 ;
        RECT 682.950 310.950 685.050 311.250 ;
        RECT 694.050 310.950 694.950 315.000 ;
        RECT 704.100 313.800 705.150 315.000 ;
        RECT 704.100 312.600 711.000 313.800 ;
        RECT 704.100 312.000 705.900 312.600 ;
        RECT 710.100 311.850 711.000 312.600 ;
        RECT 707.100 310.950 708.900 311.700 ;
        RECT 694.050 308.850 697.050 310.950 ;
        RECT 700.950 309.900 708.900 310.950 ;
        RECT 710.100 310.050 711.900 311.850 ;
        RECT 700.950 308.850 703.050 309.900 ;
        RECT 682.950 305.400 684.750 307.200 ;
        RECT 683.850 304.200 688.050 305.400 ;
        RECT 694.050 304.200 694.950 308.850 ;
        RECT 702.750 305.100 704.550 305.400 ;
        RECT 647.550 291.750 649.350 297.600 ;
        RECT 650.550 291.750 652.350 297.600 ;
        RECT 660.450 291.750 662.250 303.600 ;
        RECT 664.650 291.750 666.450 303.600 ;
        RECT 672.450 291.750 674.250 303.600 ;
        RECT 676.650 291.750 678.450 303.600 ;
        RECT 680.550 291.750 682.350 303.600 ;
        RECT 685.950 303.300 688.050 304.200 ;
        RECT 688.950 303.300 694.950 304.200 ;
        RECT 696.150 304.800 704.550 305.100 ;
        RECT 712.950 304.800 713.850 317.400 ;
        RECT 696.150 304.200 713.850 304.800 ;
        RECT 688.950 302.400 689.850 303.300 ;
        RECT 687.150 300.600 689.850 302.400 ;
        RECT 690.750 302.100 692.550 302.400 ;
        RECT 696.150 302.100 697.050 304.200 ;
        RECT 702.750 303.600 713.850 304.200 ;
        RECT 690.750 301.200 697.050 302.100 ;
        RECT 697.950 302.700 699.750 303.300 ;
        RECT 697.950 301.500 705.450 302.700 ;
        RECT 690.750 300.600 692.550 301.200 ;
        RECT 704.250 300.600 705.450 301.500 ;
        RECT 685.950 297.600 689.850 299.700 ;
        RECT 694.950 298.500 701.850 300.300 ;
        RECT 704.250 298.500 709.050 300.600 ;
        RECT 683.550 291.750 685.350 294.600 ;
        RECT 688.050 291.750 689.850 297.600 ;
        RECT 692.250 291.750 694.050 297.600 ;
        RECT 696.150 291.750 697.950 298.500 ;
        RECT 704.250 297.600 705.450 298.500 ;
        RECT 699.150 291.750 700.950 297.600 ;
        RECT 703.950 291.750 705.750 297.600 ;
        RECT 709.050 291.750 710.850 297.600 ;
        RECT 712.050 291.750 713.850 303.600 ;
        RECT 4.650 286.500 12.450 287.250 ;
        RECT 4.650 275.400 6.450 286.500 ;
        RECT 7.650 275.400 9.450 285.600 ;
        RECT 10.650 276.600 12.450 286.500 ;
        RECT 13.650 277.500 15.450 287.250 ;
        RECT 16.650 276.600 18.450 287.250 ;
        RECT 10.650 275.700 18.450 276.600 ;
        RECT 21.300 275.400 23.100 287.250 ;
        RECT 25.500 275.400 27.300 287.250 ;
        RECT 28.800 281.400 30.600 287.250 ;
        RECT 35.550 281.400 37.350 287.250 ;
        RECT 38.550 281.400 40.350 287.250 ;
        RECT 41.550 281.400 43.350 287.250 ;
        RECT 49.650 281.400 51.450 287.250 ;
        RECT 52.650 282.000 54.450 287.250 ;
        RECT 7.800 274.500 9.600 275.400 ;
        RECT 7.800 273.600 11.850 274.500 ;
        RECT 5.100 270.150 6.900 271.950 ;
        RECT 10.950 270.150 11.850 273.600 ;
        RECT 16.950 270.150 18.750 271.950 ;
        RECT 20.100 270.150 21.900 271.950 ;
        RECT 25.950 270.150 27.150 275.400 ;
        RECT 31.950 274.950 34.050 277.050 ;
        RECT 28.950 273.150 30.750 274.950 ;
        RECT 28.950 271.050 31.050 273.150 ;
        RECT 4.950 268.050 7.050 270.150 ;
        RECT 7.950 266.850 10.050 268.950 ;
        RECT 10.950 268.050 13.050 270.150 ;
        RECT 8.250 265.050 10.050 266.850 ;
        RECT 12.000 261.600 13.050 268.050 ;
        RECT 13.950 266.850 16.050 268.950 ;
        RECT 16.950 268.050 19.050 270.150 ;
        RECT 19.950 268.050 22.050 270.150 ;
        RECT 22.950 266.850 25.050 268.950 ;
        RECT 25.950 268.050 28.050 270.150 ;
        RECT 13.950 265.050 15.750 266.850 ;
        RECT 23.100 265.050 24.900 266.850 ;
        RECT 26.850 264.750 28.050 268.050 ;
        RECT 28.950 267.450 31.050 268.050 ;
        RECT 32.550 267.450 33.450 274.950 ;
        RECT 38.550 273.150 39.750 281.400 ;
        RECT 50.250 281.100 51.450 281.400 ;
        RECT 55.650 281.400 57.450 287.250 ;
        RECT 58.650 281.400 60.450 287.250 ;
        RECT 55.650 281.100 57.300 281.400 ;
        RECT 50.250 280.200 57.300 281.100 ;
        RECT 34.950 269.850 37.050 271.950 ;
        RECT 37.950 271.050 40.050 273.150 ;
        RECT 50.250 271.950 51.300 280.200 ;
        RECT 56.100 276.150 57.900 277.950 ;
        RECT 62.550 276.600 64.350 287.250 ;
        RECT 65.550 277.500 67.350 287.250 ;
        RECT 68.550 286.500 76.350 287.250 ;
        RECT 68.550 276.600 70.350 286.500 ;
        RECT 52.950 273.150 54.750 274.950 ;
        RECT 55.950 274.050 58.050 276.150 ;
        RECT 62.550 275.700 70.350 276.600 ;
        RECT 71.550 275.400 73.350 285.600 ;
        RECT 74.550 275.400 76.350 286.500 ;
        RECT 80.550 281.400 82.350 287.250 ;
        RECT 83.550 281.400 85.350 287.250 ;
        RECT 59.100 273.150 60.900 274.950 ;
        RECT 71.400 274.500 73.200 275.400 ;
        RECT 69.150 273.600 73.200 274.500 ;
        RECT 35.100 268.050 36.900 269.850 ;
        RECT 28.950 266.550 33.450 267.450 ;
        RECT 28.950 265.950 31.050 266.550 ;
        RECT 27.000 263.700 30.750 264.750 ;
        RECT 7.800 255.750 9.600 261.600 ;
        RECT 12.000 255.750 13.800 261.600 ;
        RECT 16.200 255.750 18.000 261.600 ;
        RECT 20.550 260.700 28.350 262.050 ;
        RECT 20.550 255.750 22.350 260.700 ;
        RECT 23.550 255.750 25.350 259.800 ;
        RECT 26.550 255.750 28.350 260.700 ;
        RECT 29.550 261.600 30.750 263.700 ;
        RECT 38.550 263.700 39.750 271.050 ;
        RECT 40.950 269.850 43.050 271.950 ;
        RECT 49.950 269.850 52.050 271.950 ;
        RECT 52.950 271.050 55.050 273.150 ;
        RECT 58.950 271.050 61.050 273.150 ;
        RECT 62.250 270.150 64.050 271.950 ;
        RECT 69.150 270.150 70.050 273.600 ;
        RECT 74.100 270.150 75.900 271.950 ;
        RECT 80.100 270.150 81.900 271.950 ;
        RECT 41.100 268.050 42.900 269.850 ;
        RECT 50.400 265.650 51.600 269.850 ;
        RECT 61.950 268.050 64.050 270.150 ;
        RECT 64.950 266.850 67.050 268.950 ;
        RECT 50.400 264.000 54.900 265.650 ;
        RECT 65.250 265.050 67.050 266.850 ;
        RECT 67.950 268.050 70.050 270.150 ;
        RECT 38.550 262.800 42.150 263.700 ;
        RECT 29.550 255.750 31.350 261.600 ;
        RECT 35.850 255.750 37.650 261.600 ;
        RECT 40.350 255.750 42.150 262.800 ;
        RECT 53.100 255.750 54.900 264.000 ;
        RECT 58.500 255.750 60.300 264.600 ;
        RECT 67.950 261.600 69.000 268.050 ;
        RECT 70.950 266.850 73.050 268.950 ;
        RECT 73.950 268.050 76.050 270.150 ;
        RECT 79.950 268.050 82.050 270.150 ;
        RECT 70.950 265.050 72.750 266.850 ;
        RECT 83.700 264.300 84.900 281.400 ;
        RECT 87.150 275.400 88.950 287.250 ;
        RECT 90.150 275.400 91.950 287.250 ;
        RECT 97.650 275.400 99.450 287.250 ;
        RECT 100.650 275.400 102.450 287.250 ;
        RECT 104.550 281.400 106.350 287.250 ;
        RECT 85.950 269.850 88.050 271.950 ;
        RECT 90.150 270.150 91.350 275.400 ;
        RECT 98.400 270.150 99.600 275.400 ;
        RECT 104.550 274.500 105.750 281.400 ;
        RECT 107.850 275.400 109.650 287.250 ;
        RECT 110.850 275.400 112.650 287.250 ;
        RECT 119.400 281.400 121.200 287.250 ;
        RECT 122.700 275.400 124.500 287.250 ;
        RECT 126.900 275.400 128.700 287.250 ;
        RECT 132.300 275.400 134.100 287.250 ;
        RECT 136.500 275.400 138.300 287.250 ;
        RECT 139.800 281.400 141.600 287.250 ;
        RECT 146.550 281.400 148.350 287.250 ;
        RECT 149.550 281.400 151.350 287.250 ;
        RECT 152.550 282.000 154.350 287.250 ;
        RECT 149.700 281.100 151.350 281.400 ;
        RECT 155.550 281.400 157.350 287.250 ;
        RECT 161.550 281.400 163.350 287.250 ;
        RECT 164.550 281.400 166.350 287.250 ;
        RECT 170.550 281.400 172.350 287.250 ;
        RECT 173.550 281.400 175.350 287.250 ;
        RECT 176.550 282.000 178.350 287.250 ;
        RECT 155.550 281.100 156.750 281.400 ;
        RECT 149.700 280.200 156.750 281.100 ;
        RECT 149.100 276.150 150.900 277.950 ;
        RECT 104.550 273.600 110.250 274.500 ;
        RECT 108.000 272.700 110.250 273.600 ;
        RECT 104.100 270.150 105.900 271.950 ;
        RECT 86.100 268.050 87.900 269.850 ;
        RECT 88.950 268.050 91.350 270.150 ;
        RECT 97.950 268.050 100.050 270.150 ;
        RECT 80.550 263.100 88.050 264.300 ;
        RECT 63.000 255.750 64.800 261.600 ;
        RECT 67.200 255.750 69.000 261.600 ;
        RECT 71.400 255.750 73.200 261.600 ;
        RECT 80.550 255.750 82.350 263.100 ;
        RECT 86.250 262.500 88.050 263.100 ;
        RECT 90.150 261.600 91.350 268.050 ;
        RECT 98.400 261.600 99.600 268.050 ;
        RECT 100.950 266.850 103.050 268.950 ;
        RECT 103.950 268.050 106.050 270.150 ;
        RECT 101.100 265.050 102.900 266.850 ;
        RECT 108.000 264.300 109.050 272.700 ;
        RECT 111.150 270.150 112.350 275.400 ;
        RECT 119.250 273.150 121.050 274.950 ;
        RECT 118.950 271.050 121.050 273.150 ;
        RECT 122.850 270.150 124.050 275.400 ;
        RECT 128.100 270.150 129.900 271.950 ;
        RECT 131.100 270.150 132.900 271.950 ;
        RECT 136.950 270.150 138.150 275.400 ;
        RECT 139.950 273.150 141.750 274.950 ;
        RECT 146.100 273.150 147.900 274.950 ;
        RECT 148.950 274.050 151.050 276.150 ;
        RECT 152.250 273.150 154.050 274.950 ;
        RECT 139.950 271.050 142.050 273.150 ;
        RECT 145.950 271.050 148.050 273.150 ;
        RECT 151.950 271.050 154.050 273.150 ;
        RECT 155.700 271.950 156.750 280.200 ;
        RECT 109.950 268.050 112.350 270.150 ;
        RECT 108.000 263.400 110.250 264.300 ;
        RECT 105.150 262.500 110.250 263.400 ;
        RECT 85.050 255.750 86.850 261.600 ;
        RECT 88.050 260.100 91.350 261.600 ;
        RECT 88.050 255.750 89.850 260.100 ;
        RECT 97.650 255.750 99.450 261.600 ;
        RECT 100.650 255.750 102.450 261.600 ;
        RECT 105.150 258.600 106.350 262.500 ;
        RECT 111.150 261.600 112.350 268.050 ;
        RECT 121.950 268.050 124.050 270.150 ;
        RECT 121.950 264.750 123.150 268.050 ;
        RECT 124.950 266.850 127.050 268.950 ;
        RECT 127.950 268.050 130.050 270.150 ;
        RECT 130.950 268.050 133.050 270.150 ;
        RECT 133.950 266.850 136.050 268.950 ;
        RECT 136.950 268.050 139.050 270.150 ;
        RECT 154.950 269.850 157.050 271.950 ;
        RECT 125.100 265.050 126.900 266.850 ;
        RECT 134.100 265.050 135.900 266.850 ;
        RECT 137.850 264.750 139.050 268.050 ;
        RECT 155.400 265.650 156.600 269.850 ;
        RECT 164.400 268.950 165.600 281.400 ;
        RECT 173.700 281.100 175.350 281.400 ;
        RECT 179.550 281.400 181.350 287.250 ;
        RECT 185.550 281.400 187.350 287.250 ;
        RECT 188.550 281.400 190.350 287.250 ;
        RECT 191.550 282.000 193.350 287.250 ;
        RECT 179.550 281.100 180.750 281.400 ;
        RECT 173.700 280.200 180.750 281.100 ;
        RECT 188.700 281.100 190.350 281.400 ;
        RECT 194.550 281.400 196.350 287.250 ;
        RECT 202.650 281.400 204.450 287.250 ;
        RECT 205.650 281.400 207.450 287.250 ;
        RECT 211.650 286.500 219.450 287.250 ;
        RECT 194.550 281.100 195.750 281.400 ;
        RECT 188.700 280.200 195.750 281.100 ;
        RECT 169.950 279.450 172.050 280.050 ;
        RECT 167.550 278.550 172.050 279.450 ;
        RECT 161.100 267.150 162.900 268.950 ;
        RECT 119.250 263.700 123.000 264.750 ;
        RECT 138.000 263.700 141.750 264.750 ;
        RECT 119.250 261.600 120.450 263.700 ;
        RECT 104.550 255.750 106.350 258.600 ;
        RECT 107.850 255.750 109.650 261.600 ;
        RECT 110.850 255.750 112.650 261.600 ;
        RECT 118.650 255.750 120.450 261.600 ;
        RECT 121.650 260.700 129.450 262.050 ;
        RECT 121.650 255.750 123.450 260.700 ;
        RECT 124.650 255.750 126.450 259.800 ;
        RECT 127.650 255.750 129.450 260.700 ;
        RECT 131.550 260.700 139.350 262.050 ;
        RECT 131.550 255.750 133.350 260.700 ;
        RECT 134.550 255.750 136.350 259.800 ;
        RECT 137.550 255.750 139.350 260.700 ;
        RECT 140.550 261.600 141.750 263.700 ;
        RECT 140.550 255.750 142.350 261.600 ;
        RECT 146.700 255.750 148.500 264.600 ;
        RECT 152.100 264.000 156.600 265.650 ;
        RECT 160.950 265.050 163.050 267.150 ;
        RECT 163.950 266.850 166.050 268.950 ;
        RECT 167.550 267.450 168.450 278.550 ;
        RECT 169.950 277.950 172.050 278.550 ;
        RECT 173.100 276.150 174.900 277.950 ;
        RECT 170.100 273.150 171.900 274.950 ;
        RECT 172.950 274.050 175.050 276.150 ;
        RECT 176.250 273.150 178.050 274.950 ;
        RECT 169.950 271.050 172.050 273.150 ;
        RECT 175.950 271.050 178.050 273.150 ;
        RECT 179.700 271.950 180.750 280.200 ;
        RECT 188.100 276.150 189.900 277.950 ;
        RECT 185.100 273.150 186.900 274.950 ;
        RECT 187.950 274.050 190.050 276.150 ;
        RECT 191.250 273.150 193.050 274.950 ;
        RECT 178.950 269.850 181.050 271.950 ;
        RECT 184.950 271.050 187.050 273.150 ;
        RECT 190.950 271.050 193.050 273.150 ;
        RECT 194.700 271.950 195.750 280.200 ;
        RECT 193.950 269.850 196.050 271.950 ;
        RECT 172.950 267.450 175.050 268.050 ;
        RECT 152.100 255.750 153.900 264.000 ;
        RECT 164.400 258.600 165.600 266.850 ;
        RECT 167.550 266.550 175.050 267.450 ;
        RECT 172.950 265.950 175.050 266.550 ;
        RECT 179.400 265.650 180.600 269.850 ;
        RECT 194.400 265.650 195.600 269.850 ;
        RECT 203.400 268.950 204.600 281.400 ;
        RECT 211.650 275.400 213.450 286.500 ;
        RECT 214.650 275.400 216.450 285.600 ;
        RECT 217.650 276.600 219.450 286.500 ;
        RECT 220.650 277.500 222.450 287.250 ;
        RECT 223.650 276.600 225.450 287.250 ;
        RECT 227.550 281.400 229.350 287.250 ;
        RECT 230.550 281.400 232.350 287.250 ;
        RECT 233.550 282.000 235.350 287.250 ;
        RECT 230.700 281.100 232.350 281.400 ;
        RECT 236.550 281.400 238.350 287.250 ;
        RECT 242.550 281.400 244.350 287.250 ;
        RECT 245.550 281.400 247.350 287.250 ;
        RECT 236.550 281.100 237.750 281.400 ;
        RECT 230.700 280.200 237.750 281.100 ;
        RECT 217.650 275.700 225.450 276.600 ;
        RECT 230.100 276.150 231.900 277.950 ;
        RECT 214.800 274.500 216.600 275.400 ;
        RECT 214.800 273.600 218.850 274.500 ;
        RECT 212.100 270.150 213.900 271.950 ;
        RECT 217.950 270.150 218.850 273.600 ;
        RECT 227.100 273.150 228.900 274.950 ;
        RECT 229.950 274.050 232.050 276.150 ;
        RECT 233.250 273.150 235.050 274.950 ;
        RECT 223.950 270.150 225.750 271.950 ;
        RECT 226.950 271.050 229.050 273.150 ;
        RECT 232.950 271.050 235.050 273.150 ;
        RECT 236.700 271.950 237.750 280.200 ;
        RECT 202.950 266.850 205.050 268.950 ;
        RECT 206.100 267.150 207.900 268.950 ;
        RECT 211.950 268.050 214.050 270.150 ;
        RECT 161.550 255.750 163.350 258.600 ;
        RECT 164.550 255.750 166.350 258.600 ;
        RECT 170.700 255.750 172.500 264.600 ;
        RECT 176.100 264.000 180.600 265.650 ;
        RECT 176.100 255.750 177.900 264.000 ;
        RECT 185.700 255.750 187.500 264.600 ;
        RECT 191.100 264.000 195.600 265.650 ;
        RECT 191.100 255.750 192.900 264.000 ;
        RECT 203.400 258.600 204.600 266.850 ;
        RECT 205.950 265.050 208.050 267.150 ;
        RECT 214.950 266.850 217.050 268.950 ;
        RECT 217.950 268.050 220.050 270.150 ;
        RECT 215.250 265.050 217.050 266.850 ;
        RECT 219.000 261.600 220.050 268.050 ;
        RECT 220.950 266.850 223.050 268.950 ;
        RECT 223.950 268.050 226.050 270.150 ;
        RECT 235.950 269.850 238.050 271.950 ;
        RECT 220.950 265.050 222.750 266.850 ;
        RECT 236.400 265.650 237.600 269.850 ;
        RECT 245.400 268.950 246.600 281.400 ;
        RECT 253.650 275.400 255.450 287.250 ;
        RECT 256.650 275.400 258.450 287.250 ;
        RECT 262.650 281.400 264.450 287.250 ;
        RECT 265.650 282.000 267.450 287.250 ;
        RECT 263.250 281.100 264.450 281.400 ;
        RECT 268.650 281.400 270.450 287.250 ;
        RECT 271.650 281.400 273.450 287.250 ;
        RECT 275.550 281.400 277.350 287.250 ;
        RECT 278.550 281.400 280.350 287.250 ;
        RECT 268.650 281.100 270.300 281.400 ;
        RECT 263.250 280.200 270.300 281.100 ;
        RECT 254.400 270.150 255.600 275.400 ;
        RECT 263.250 271.950 264.300 280.200 ;
        RECT 269.100 276.150 270.900 277.950 ;
        RECT 265.950 273.150 267.750 274.950 ;
        RECT 268.950 274.050 271.050 276.150 ;
        RECT 272.100 273.150 273.900 274.950 ;
        RECT 242.100 267.150 243.900 268.950 ;
        RECT 202.650 255.750 204.450 258.600 ;
        RECT 205.650 255.750 207.450 258.600 ;
        RECT 214.800 255.750 216.600 261.600 ;
        RECT 219.000 255.750 220.800 261.600 ;
        RECT 223.200 255.750 225.000 261.600 ;
        RECT 227.700 255.750 229.500 264.600 ;
        RECT 233.100 264.000 237.600 265.650 ;
        RECT 241.950 265.050 244.050 267.150 ;
        RECT 244.950 266.850 247.050 268.950 ;
        RECT 253.950 268.050 256.050 270.150 ;
        RECT 262.950 269.850 265.050 271.950 ;
        RECT 265.950 271.050 268.050 273.150 ;
        RECT 271.950 271.050 274.050 273.150 ;
        RECT 275.100 270.150 276.900 271.950 ;
        RECT 233.100 255.750 234.900 264.000 ;
        RECT 245.400 258.600 246.600 266.850 ;
        RECT 254.400 261.600 255.600 268.050 ;
        RECT 256.950 266.850 259.050 268.950 ;
        RECT 257.100 265.050 258.900 266.850 ;
        RECT 263.400 265.650 264.600 269.850 ;
        RECT 274.950 268.050 277.050 270.150 ;
        RECT 263.400 264.000 267.900 265.650 ;
        RECT 242.550 255.750 244.350 258.600 ;
        RECT 245.550 255.750 247.350 258.600 ;
        RECT 253.650 255.750 255.450 261.600 ;
        RECT 256.650 255.750 258.450 261.600 ;
        RECT 266.100 255.750 267.900 264.000 ;
        RECT 271.500 255.750 273.300 264.600 ;
        RECT 278.700 264.300 279.900 281.400 ;
        RECT 282.150 275.400 283.950 287.250 ;
        RECT 285.150 275.400 286.950 287.250 ;
        RECT 291.150 275.400 292.950 287.250 ;
        RECT 294.150 281.400 295.950 287.250 ;
        RECT 299.250 281.400 301.050 287.250 ;
        RECT 304.050 281.400 305.850 287.250 ;
        RECT 299.550 280.500 300.750 281.400 ;
        RECT 307.050 280.500 308.850 287.250 ;
        RECT 310.950 281.400 312.750 287.250 ;
        RECT 315.150 281.400 316.950 287.250 ;
        RECT 319.650 284.400 321.450 287.250 ;
        RECT 295.950 278.400 300.750 280.500 ;
        RECT 303.150 278.700 310.050 280.500 ;
        RECT 315.150 279.300 319.050 281.400 ;
        RECT 299.550 277.500 300.750 278.400 ;
        RECT 312.450 277.800 314.250 278.400 ;
        RECT 299.550 276.300 307.050 277.500 ;
        RECT 305.250 275.700 307.050 276.300 ;
        RECT 307.950 276.900 314.250 277.800 ;
        RECT 280.950 269.850 283.050 271.950 ;
        RECT 285.150 270.150 286.350 275.400 ;
        RECT 281.100 268.050 282.900 269.850 ;
        RECT 283.950 268.050 286.350 270.150 ;
        RECT 275.550 263.100 283.050 264.300 ;
        RECT 275.550 255.750 277.350 263.100 ;
        RECT 281.250 262.500 283.050 263.100 ;
        RECT 285.150 261.600 286.350 268.050 ;
        RECT 280.050 255.750 281.850 261.600 ;
        RECT 283.050 260.100 286.350 261.600 ;
        RECT 291.150 274.800 302.250 275.400 ;
        RECT 307.950 274.800 308.850 276.900 ;
        RECT 312.450 276.600 314.250 276.900 ;
        RECT 315.150 276.600 317.850 278.400 ;
        RECT 315.150 275.700 316.050 276.600 ;
        RECT 291.150 274.200 308.850 274.800 ;
        RECT 291.150 261.600 292.050 274.200 ;
        RECT 300.450 273.900 308.850 274.200 ;
        RECT 310.050 274.800 316.050 275.700 ;
        RECT 316.950 274.800 319.050 275.700 ;
        RECT 322.650 275.400 324.450 287.250 ;
        RECT 300.450 273.600 302.250 273.900 ;
        RECT 310.050 270.150 310.950 274.800 ;
        RECT 316.950 273.600 321.150 274.800 ;
        RECT 320.250 271.800 322.050 273.600 ;
        RECT 301.950 269.100 304.050 270.150 ;
        RECT 293.100 267.150 294.900 268.950 ;
        RECT 296.100 268.050 304.050 269.100 ;
        RECT 307.950 268.050 310.950 270.150 ;
        RECT 296.100 267.300 297.900 268.050 ;
        RECT 294.000 266.400 294.900 267.150 ;
        RECT 299.100 266.400 300.900 267.000 ;
        RECT 294.000 265.200 300.900 266.400 ;
        RECT 299.850 264.000 300.900 265.200 ;
        RECT 310.050 264.000 310.950 268.050 ;
        RECT 319.950 267.750 322.050 268.050 ;
        RECT 318.150 265.950 322.050 267.750 ;
        RECT 323.250 265.950 324.450 275.400 ;
        RECT 330.450 275.400 332.250 287.250 ;
        RECT 334.650 275.400 336.450 287.250 ;
        RECT 338.550 281.400 340.350 287.250 ;
        RECT 341.550 281.400 343.350 287.250 ;
        RECT 330.450 274.350 333.000 275.400 ;
        RECT 329.100 270.150 330.900 271.950 ;
        RECT 328.950 268.050 331.050 270.150 ;
        RECT 299.850 263.100 310.950 264.000 ;
        RECT 319.950 263.850 324.450 265.950 ;
        RECT 299.850 262.200 300.900 263.100 ;
        RECT 310.050 262.800 310.950 263.100 ;
        RECT 283.050 255.750 284.850 260.100 ;
        RECT 291.150 255.750 292.950 261.600 ;
        RECT 295.950 259.500 298.050 261.600 ;
        RECT 299.550 260.400 301.350 262.200 ;
        RECT 302.850 261.450 304.650 262.200 ;
        RECT 302.850 260.400 307.800 261.450 ;
        RECT 310.050 261.000 311.850 262.800 ;
        RECT 323.250 261.600 324.450 263.850 ;
        RECT 316.950 260.700 319.050 261.600 ;
        RECT 297.000 258.600 298.050 259.500 ;
        RECT 306.750 258.600 307.800 260.400 ;
        RECT 315.300 259.500 319.050 260.700 ;
        RECT 315.300 258.600 316.350 259.500 ;
        RECT 294.150 255.750 295.950 258.600 ;
        RECT 297.000 257.700 300.750 258.600 ;
        RECT 298.950 255.750 300.750 257.700 ;
        RECT 303.450 255.750 305.250 258.600 ;
        RECT 306.750 255.750 308.550 258.600 ;
        RECT 310.650 255.750 312.450 258.600 ;
        RECT 314.850 255.750 316.650 258.600 ;
        RECT 319.350 255.750 321.150 258.600 ;
        RECT 322.650 255.750 324.450 261.600 ;
        RECT 331.950 267.150 333.000 274.350 ;
        RECT 335.100 270.150 336.900 271.950 ;
        RECT 334.950 268.050 337.050 270.150 ;
        RECT 341.400 268.950 342.600 281.400 ;
        RECT 348.300 275.400 350.100 287.250 ;
        RECT 352.500 275.400 354.300 287.250 ;
        RECT 355.800 281.400 357.600 287.250 ;
        RECT 362.550 275.400 364.350 287.250 ;
        RECT 366.750 275.400 368.550 287.250 ;
        RECT 374.550 275.400 376.350 287.250 ;
        RECT 378.750 275.400 380.550 287.250 ;
        RECT 387.300 275.400 389.100 287.250 ;
        RECT 391.500 275.400 393.300 287.250 ;
        RECT 394.800 281.400 396.600 287.250 ;
        RECT 403.650 281.400 405.450 287.250 ;
        RECT 406.650 281.400 408.450 287.250 ;
        RECT 409.650 281.400 411.450 287.250 ;
        RECT 347.100 270.150 348.900 271.950 ;
        RECT 352.950 270.150 354.150 275.400 ;
        RECT 355.950 273.150 357.750 274.950 ;
        RECT 366.000 274.350 368.550 275.400 ;
        RECT 378.000 274.350 380.550 275.400 ;
        RECT 355.950 271.050 358.050 273.150 ;
        RECT 362.100 270.150 363.900 271.950 ;
        RECT 338.100 267.150 339.900 268.950 ;
        RECT 331.950 265.050 334.050 267.150 ;
        RECT 337.950 265.050 340.050 267.150 ;
        RECT 340.950 266.850 343.050 268.950 ;
        RECT 346.950 268.050 349.050 270.150 ;
        RECT 349.950 266.850 352.050 268.950 ;
        RECT 352.950 268.050 355.050 270.150 ;
        RECT 361.950 268.050 364.050 270.150 ;
        RECT 331.950 258.600 333.000 265.050 ;
        RECT 341.400 258.600 342.600 266.850 ;
        RECT 350.100 265.050 351.900 266.850 ;
        RECT 353.850 264.750 355.050 268.050 ;
        RECT 366.000 267.150 367.050 274.350 ;
        RECT 368.100 270.150 369.900 271.950 ;
        RECT 374.100 270.150 375.900 271.950 ;
        RECT 367.950 268.050 370.050 270.150 ;
        RECT 373.950 268.050 376.050 270.150 ;
        RECT 378.000 267.150 379.050 274.350 ;
        RECT 380.100 270.150 381.900 271.950 ;
        RECT 386.100 270.150 387.900 271.950 ;
        RECT 391.950 270.150 393.150 275.400 ;
        RECT 394.950 273.150 396.750 274.950 ;
        RECT 407.250 273.150 408.450 281.400 ;
        RECT 417.450 275.400 419.250 287.250 ;
        RECT 421.650 275.400 423.450 287.250 ;
        RECT 426.300 275.400 428.100 287.250 ;
        RECT 430.500 275.400 432.300 287.250 ;
        RECT 433.800 281.400 435.600 287.250 ;
        RECT 440.550 281.400 442.350 287.250 ;
        RECT 443.550 281.400 445.350 287.250 ;
        RECT 417.450 274.350 420.000 275.400 ;
        RECT 394.950 271.050 397.050 273.150 ;
        RECT 379.950 268.050 382.050 270.150 ;
        RECT 385.950 268.050 388.050 270.150 ;
        RECT 364.950 265.050 367.050 267.150 ;
        RECT 376.950 265.050 379.050 267.150 ;
        RECT 388.950 266.850 391.050 268.950 ;
        RECT 391.950 268.050 394.050 270.150 ;
        RECT 403.950 269.850 406.050 271.950 ;
        RECT 406.950 271.050 409.050 273.150 ;
        RECT 404.100 268.050 405.900 269.850 ;
        RECT 389.100 265.050 390.900 266.850 ;
        RECT 354.000 263.700 357.750 264.750 ;
        RECT 347.550 260.700 355.350 262.050 ;
        RECT 328.650 255.750 330.450 258.600 ;
        RECT 331.650 255.750 333.450 258.600 ;
        RECT 334.650 255.750 336.450 258.600 ;
        RECT 338.550 255.750 340.350 258.600 ;
        RECT 341.550 255.750 343.350 258.600 ;
        RECT 347.550 255.750 349.350 260.700 ;
        RECT 350.550 255.750 352.350 259.800 ;
        RECT 353.550 255.750 355.350 260.700 ;
        RECT 356.550 261.600 357.750 263.700 ;
        RECT 356.550 255.750 358.350 261.600 ;
        RECT 366.000 258.600 367.050 265.050 ;
        RECT 378.000 258.600 379.050 265.050 ;
        RECT 392.850 264.750 394.050 268.050 ;
        RECT 393.000 263.700 396.750 264.750 ;
        RECT 407.250 263.700 408.450 271.050 ;
        RECT 409.950 269.850 412.050 271.950 ;
        RECT 416.100 270.150 417.900 271.950 ;
        RECT 410.100 268.050 411.900 269.850 ;
        RECT 415.950 268.050 418.050 270.150 ;
        RECT 386.550 260.700 394.350 262.050 ;
        RECT 362.550 255.750 364.350 258.600 ;
        RECT 365.550 255.750 367.350 258.600 ;
        RECT 368.550 255.750 370.350 258.600 ;
        RECT 374.550 255.750 376.350 258.600 ;
        RECT 377.550 255.750 379.350 258.600 ;
        RECT 380.550 255.750 382.350 258.600 ;
        RECT 386.550 255.750 388.350 260.700 ;
        RECT 389.550 255.750 391.350 259.800 ;
        RECT 392.550 255.750 394.350 260.700 ;
        RECT 395.550 261.600 396.750 263.700 ;
        RECT 404.850 262.800 408.450 263.700 ;
        RECT 418.950 267.150 420.000 274.350 ;
        RECT 422.100 270.150 423.900 271.950 ;
        RECT 425.100 270.150 426.900 271.950 ;
        RECT 430.950 270.150 432.150 275.400 ;
        RECT 433.950 273.150 435.750 274.950 ;
        RECT 433.950 271.050 436.050 273.150 ;
        RECT 421.950 268.050 424.050 270.150 ;
        RECT 424.950 268.050 427.050 270.150 ;
        RECT 418.950 265.050 421.050 267.150 ;
        RECT 427.950 266.850 430.050 268.950 ;
        RECT 430.950 268.050 433.050 270.150 ;
        RECT 443.400 268.950 444.600 281.400 ;
        RECT 453.450 275.400 455.250 287.250 ;
        RECT 457.650 275.400 459.450 287.250 ;
        RECT 461.550 275.400 463.350 287.250 ;
        RECT 464.550 284.400 466.350 287.250 ;
        RECT 469.050 281.400 470.850 287.250 ;
        RECT 473.250 281.400 475.050 287.250 ;
        RECT 466.950 279.300 470.850 281.400 ;
        RECT 477.150 280.500 478.950 287.250 ;
        RECT 480.150 281.400 481.950 287.250 ;
        RECT 484.950 281.400 486.750 287.250 ;
        RECT 490.050 281.400 491.850 287.250 ;
        RECT 485.250 280.500 486.450 281.400 ;
        RECT 475.950 278.700 482.850 280.500 ;
        RECT 485.250 278.400 490.050 280.500 ;
        RECT 468.150 276.600 470.850 278.400 ;
        RECT 471.750 277.800 473.550 278.400 ;
        RECT 471.750 276.900 478.050 277.800 ;
        RECT 485.250 277.500 486.450 278.400 ;
        RECT 471.750 276.600 473.550 276.900 ;
        RECT 469.950 275.700 470.850 276.600 ;
        RECT 453.450 274.350 456.000 275.400 ;
        RECT 452.100 270.150 453.900 271.950 ;
        RECT 428.100 265.050 429.900 266.850 ;
        RECT 395.550 255.750 397.350 261.600 ;
        RECT 404.850 255.750 406.650 262.800 ;
        RECT 409.350 255.750 411.150 261.600 ;
        RECT 418.950 258.600 420.000 265.050 ;
        RECT 431.850 264.750 433.050 268.050 ;
        RECT 440.100 267.150 441.900 268.950 ;
        RECT 439.950 265.050 442.050 267.150 ;
        RECT 442.950 266.850 445.050 268.950 ;
        RECT 451.950 268.050 454.050 270.150 ;
        RECT 454.950 267.150 456.000 274.350 ;
        RECT 458.100 270.150 459.900 271.950 ;
        RECT 457.950 268.050 460.050 270.150 ;
        RECT 432.000 263.700 435.750 264.750 ;
        RECT 425.550 260.700 433.350 262.050 ;
        RECT 415.650 255.750 417.450 258.600 ;
        RECT 418.650 255.750 420.450 258.600 ;
        RECT 421.650 255.750 423.450 258.600 ;
        RECT 425.550 255.750 427.350 260.700 ;
        RECT 428.550 255.750 430.350 259.800 ;
        RECT 431.550 255.750 433.350 260.700 ;
        RECT 434.550 261.600 435.750 263.700 ;
        RECT 434.550 255.750 436.350 261.600 ;
        RECT 443.400 258.600 444.600 266.850 ;
        RECT 454.950 265.050 457.050 267.150 ;
        RECT 461.550 265.950 462.750 275.400 ;
        RECT 466.950 274.800 469.050 275.700 ;
        RECT 469.950 274.800 475.950 275.700 ;
        RECT 464.850 273.600 469.050 274.800 ;
        RECT 463.950 271.800 465.750 273.600 ;
        RECT 475.050 270.150 475.950 274.800 ;
        RECT 477.150 274.800 478.050 276.900 ;
        RECT 478.950 276.300 486.450 277.500 ;
        RECT 478.950 275.700 480.750 276.300 ;
        RECT 493.050 275.400 494.850 287.250 ;
        RECT 498.300 275.400 500.100 287.250 ;
        RECT 502.500 275.400 504.300 287.250 ;
        RECT 505.800 281.400 507.600 287.250 ;
        RECT 512.550 281.400 514.350 287.250 ;
        RECT 515.550 281.400 517.350 287.250 ;
        RECT 518.550 281.400 520.350 287.250 ;
        RECT 483.750 274.800 494.850 275.400 ;
        RECT 477.150 274.200 494.850 274.800 ;
        RECT 477.150 273.900 485.550 274.200 ;
        RECT 483.750 273.600 485.550 273.900 ;
        RECT 475.050 268.050 478.050 270.150 ;
        RECT 481.950 269.100 484.050 270.150 ;
        RECT 481.950 268.050 489.900 269.100 ;
        RECT 463.950 267.750 466.050 268.050 ;
        RECT 463.950 265.950 467.850 267.750 ;
        RECT 454.950 258.600 456.000 265.050 ;
        RECT 461.550 263.850 466.050 265.950 ;
        RECT 475.050 264.000 475.950 268.050 ;
        RECT 488.100 267.300 489.900 268.050 ;
        RECT 491.100 267.150 492.900 268.950 ;
        RECT 485.100 266.400 486.900 267.000 ;
        RECT 491.100 266.400 492.000 267.150 ;
        RECT 485.100 265.200 492.000 266.400 ;
        RECT 485.100 264.000 486.150 265.200 ;
        RECT 461.550 261.600 462.750 263.850 ;
        RECT 475.050 263.100 486.150 264.000 ;
        RECT 475.050 262.800 475.950 263.100 ;
        RECT 440.550 255.750 442.350 258.600 ;
        RECT 443.550 255.750 445.350 258.600 ;
        RECT 451.650 255.750 453.450 258.600 ;
        RECT 454.650 255.750 456.450 258.600 ;
        RECT 457.650 255.750 459.450 258.600 ;
        RECT 461.550 255.750 463.350 261.600 ;
        RECT 466.950 260.700 469.050 261.600 ;
        RECT 474.150 261.000 475.950 262.800 ;
        RECT 485.100 262.200 486.150 263.100 ;
        RECT 481.350 261.450 483.150 262.200 ;
        RECT 466.950 259.500 470.700 260.700 ;
        RECT 469.650 258.600 470.700 259.500 ;
        RECT 478.200 260.400 483.150 261.450 ;
        RECT 484.650 260.400 486.450 262.200 ;
        RECT 493.950 261.600 494.850 274.200 ;
        RECT 497.100 270.150 498.900 271.950 ;
        RECT 502.950 270.150 504.150 275.400 ;
        RECT 505.950 273.150 507.750 274.950 ;
        RECT 515.550 273.150 516.750 281.400 ;
        RECT 524.550 275.400 526.350 287.250 ;
        RECT 527.550 284.400 529.350 287.250 ;
        RECT 532.050 281.400 533.850 287.250 ;
        RECT 536.250 281.400 538.050 287.250 ;
        RECT 529.950 279.300 533.850 281.400 ;
        RECT 540.150 280.500 541.950 287.250 ;
        RECT 543.150 281.400 544.950 287.250 ;
        RECT 547.950 281.400 549.750 287.250 ;
        RECT 553.050 281.400 554.850 287.250 ;
        RECT 548.250 280.500 549.450 281.400 ;
        RECT 538.950 278.700 545.850 280.500 ;
        RECT 548.250 278.400 553.050 280.500 ;
        RECT 531.150 276.600 533.850 278.400 ;
        RECT 534.750 277.800 536.550 278.400 ;
        RECT 534.750 276.900 541.050 277.800 ;
        RECT 548.250 277.500 549.450 278.400 ;
        RECT 534.750 276.600 536.550 276.900 ;
        RECT 532.950 275.700 533.850 276.600 ;
        RECT 505.950 271.050 508.050 273.150 ;
        RECT 496.950 268.050 499.050 270.150 ;
        RECT 499.950 266.850 502.050 268.950 ;
        RECT 502.950 268.050 505.050 270.150 ;
        RECT 511.950 269.850 514.050 271.950 ;
        RECT 514.950 271.050 517.050 273.150 ;
        RECT 512.100 268.050 513.900 269.850 ;
        RECT 500.100 265.050 501.900 266.850 ;
        RECT 503.850 264.750 505.050 268.050 ;
        RECT 504.000 263.700 507.750 264.750 ;
        RECT 478.200 258.600 479.250 260.400 ;
        RECT 487.950 259.500 490.050 261.600 ;
        RECT 487.950 258.600 489.000 259.500 ;
        RECT 464.850 255.750 466.650 258.600 ;
        RECT 469.350 255.750 471.150 258.600 ;
        RECT 473.550 255.750 475.350 258.600 ;
        RECT 477.450 255.750 479.250 258.600 ;
        RECT 480.750 255.750 482.550 258.600 ;
        RECT 485.250 257.700 489.000 258.600 ;
        RECT 485.250 255.750 487.050 257.700 ;
        RECT 490.050 255.750 491.850 258.600 ;
        RECT 493.050 255.750 494.850 261.600 ;
        RECT 497.550 260.700 505.350 262.050 ;
        RECT 497.550 255.750 499.350 260.700 ;
        RECT 500.550 255.750 502.350 259.800 ;
        RECT 503.550 255.750 505.350 260.700 ;
        RECT 506.550 261.600 507.750 263.700 ;
        RECT 515.550 263.700 516.750 271.050 ;
        RECT 517.950 269.850 520.050 271.950 ;
        RECT 518.100 268.050 519.900 269.850 ;
        RECT 524.550 265.950 525.750 275.400 ;
        RECT 529.950 274.800 532.050 275.700 ;
        RECT 532.950 274.800 538.950 275.700 ;
        RECT 527.850 273.600 532.050 274.800 ;
        RECT 526.950 271.800 528.750 273.600 ;
        RECT 538.050 270.150 538.950 274.800 ;
        RECT 540.150 274.800 541.050 276.900 ;
        RECT 541.950 276.300 549.450 277.500 ;
        RECT 541.950 275.700 543.750 276.300 ;
        RECT 556.050 275.400 557.850 287.250 ;
        RECT 546.750 274.800 557.850 275.400 ;
        RECT 540.150 274.200 557.850 274.800 ;
        RECT 540.150 273.900 548.550 274.200 ;
        RECT 546.750 273.600 548.550 273.900 ;
        RECT 538.050 268.050 541.050 270.150 ;
        RECT 544.950 269.100 547.050 270.150 ;
        RECT 544.950 268.050 552.900 269.100 ;
        RECT 526.950 267.750 529.050 268.050 ;
        RECT 526.950 265.950 530.850 267.750 ;
        RECT 524.550 263.850 529.050 265.950 ;
        RECT 538.050 264.000 538.950 268.050 ;
        RECT 551.100 267.300 552.900 268.050 ;
        RECT 554.100 267.150 555.900 268.950 ;
        RECT 548.100 266.400 549.900 267.000 ;
        RECT 554.100 266.400 555.000 267.150 ;
        RECT 548.100 265.200 555.000 266.400 ;
        RECT 548.100 264.000 549.150 265.200 ;
        RECT 515.550 262.800 519.150 263.700 ;
        RECT 506.550 255.750 508.350 261.600 ;
        RECT 512.850 255.750 514.650 261.600 ;
        RECT 517.350 255.750 519.150 262.800 ;
        RECT 524.550 261.600 525.750 263.850 ;
        RECT 538.050 263.100 549.150 264.000 ;
        RECT 538.050 262.800 538.950 263.100 ;
        RECT 524.550 255.750 526.350 261.600 ;
        RECT 529.950 260.700 532.050 261.600 ;
        RECT 537.150 261.000 538.950 262.800 ;
        RECT 548.100 262.200 549.150 263.100 ;
        RECT 544.350 261.450 546.150 262.200 ;
        RECT 529.950 259.500 533.700 260.700 ;
        RECT 532.650 258.600 533.700 259.500 ;
        RECT 541.200 260.400 546.150 261.450 ;
        RECT 547.650 260.400 549.450 262.200 ;
        RECT 556.950 261.600 557.850 274.200 ;
        RECT 560.550 281.400 562.350 287.250 ;
        RECT 560.550 274.500 561.750 281.400 ;
        RECT 563.850 275.400 565.650 287.250 ;
        RECT 566.850 275.400 568.650 287.250 ;
        RECT 574.650 281.400 576.450 287.250 ;
        RECT 577.650 281.400 579.450 287.250 ;
        RECT 580.650 281.400 582.450 287.250 ;
        RECT 587.400 281.400 589.200 287.250 ;
        RECT 560.550 273.600 566.250 274.500 ;
        RECT 564.000 272.700 566.250 273.600 ;
        RECT 560.100 270.150 561.900 271.950 ;
        RECT 559.950 268.050 562.050 270.150 ;
        RECT 564.000 264.300 565.050 272.700 ;
        RECT 567.150 270.150 568.350 275.400 ;
        RECT 578.250 273.150 579.450 281.400 ;
        RECT 586.950 279.450 589.050 280.050 ;
        RECT 584.550 278.550 589.050 279.450 ;
        RECT 565.950 268.050 568.350 270.150 ;
        RECT 574.950 269.850 577.050 271.950 ;
        RECT 577.950 271.050 580.050 273.150 ;
        RECT 575.100 268.050 576.900 269.850 ;
        RECT 564.000 263.400 566.250 264.300 ;
        RECT 541.200 258.600 542.250 260.400 ;
        RECT 550.950 259.500 553.050 261.600 ;
        RECT 550.950 258.600 552.000 259.500 ;
        RECT 527.850 255.750 529.650 258.600 ;
        RECT 532.350 255.750 534.150 258.600 ;
        RECT 536.550 255.750 538.350 258.600 ;
        RECT 540.450 255.750 542.250 258.600 ;
        RECT 543.750 255.750 545.550 258.600 ;
        RECT 548.250 257.700 552.000 258.600 ;
        RECT 548.250 255.750 550.050 257.700 ;
        RECT 553.050 255.750 554.850 258.600 ;
        RECT 556.050 255.750 557.850 261.600 ;
        RECT 561.150 262.500 566.250 263.400 ;
        RECT 561.150 258.600 562.350 262.500 ;
        RECT 567.150 261.600 568.350 268.050 ;
        RECT 578.250 263.700 579.450 271.050 ;
        RECT 580.950 269.850 583.050 271.950 ;
        RECT 581.100 268.050 582.900 269.850 ;
        RECT 584.550 267.450 585.450 278.550 ;
        RECT 586.950 277.950 589.050 278.550 ;
        RECT 590.700 275.400 592.500 287.250 ;
        RECT 594.900 275.400 596.700 287.250 ;
        RECT 602.400 281.400 604.200 287.250 ;
        RECT 605.700 275.400 607.500 287.250 ;
        RECT 609.900 275.400 611.700 287.250 ;
        RECT 614.550 275.400 616.350 287.250 ;
        RECT 619.050 275.550 620.850 287.250 ;
        RECT 622.050 276.900 623.850 287.250 ;
        RECT 631.650 281.400 633.450 287.250 ;
        RECT 634.650 281.400 636.450 287.250 ;
        RECT 622.050 275.550 624.450 276.900 ;
        RECT 587.250 273.150 589.050 274.950 ;
        RECT 586.950 271.050 589.050 273.150 ;
        RECT 590.850 270.150 592.050 275.400 ;
        RECT 602.250 273.150 604.050 274.950 ;
        RECT 596.100 270.150 597.900 271.950 ;
        RECT 601.950 271.050 604.050 273.150 ;
        RECT 605.850 270.150 607.050 275.400 ;
        RECT 614.550 274.200 615.750 275.400 ;
        RECT 619.950 274.200 621.750 274.650 ;
        RECT 614.550 273.000 621.750 274.200 ;
        RECT 619.950 272.850 621.750 273.000 ;
        RECT 611.100 270.150 612.900 271.950 ;
        RECT 617.100 270.150 618.900 271.950 ;
        RECT 589.950 268.050 592.050 270.150 ;
        RECT 586.950 267.450 589.050 268.050 ;
        RECT 584.550 266.550 589.050 267.450 ;
        RECT 586.950 265.950 589.050 266.550 ;
        RECT 589.950 264.750 591.150 268.050 ;
        RECT 592.950 266.850 595.050 268.950 ;
        RECT 595.950 268.050 598.050 270.150 ;
        RECT 604.950 268.050 607.050 270.150 ;
        RECT 593.100 265.050 594.900 266.850 ;
        RECT 604.950 264.750 606.150 268.050 ;
        RECT 607.950 266.850 610.050 268.950 ;
        RECT 610.950 268.050 613.050 270.150 ;
        RECT 614.100 267.150 615.900 268.950 ;
        RECT 616.950 268.050 619.050 270.150 ;
        RECT 608.100 265.050 609.900 266.850 ;
        RECT 613.950 265.050 616.050 267.150 ;
        RECT 575.850 262.800 579.450 263.700 ;
        RECT 587.250 263.700 591.000 264.750 ;
        RECT 602.250 263.700 606.000 264.750 ;
        RECT 620.700 264.600 621.600 272.850 ;
        RECT 623.100 268.950 624.450 275.550 ;
        RECT 632.400 268.950 633.600 281.400 ;
        RECT 638.550 276.300 640.350 287.250 ;
        RECT 641.550 277.200 643.350 287.250 ;
        RECT 644.550 276.300 646.350 287.250 ;
        RECT 638.550 275.400 646.350 276.300 ;
        RECT 647.550 275.400 649.350 287.250 ;
        RECT 657.450 275.400 659.250 287.250 ;
        RECT 661.650 275.400 663.450 287.250 ;
        RECT 665.550 275.400 667.350 287.250 ;
        RECT 668.550 284.400 670.350 287.250 ;
        RECT 673.050 281.400 674.850 287.250 ;
        RECT 677.250 281.400 679.050 287.250 ;
        RECT 670.950 279.300 674.850 281.400 ;
        RECT 681.150 280.500 682.950 287.250 ;
        RECT 684.150 281.400 685.950 287.250 ;
        RECT 688.950 281.400 690.750 287.250 ;
        RECT 694.050 281.400 695.850 287.250 ;
        RECT 689.250 280.500 690.450 281.400 ;
        RECT 679.950 278.700 686.850 280.500 ;
        RECT 689.250 278.400 694.050 280.500 ;
        RECT 672.150 276.600 674.850 278.400 ;
        RECT 675.750 277.800 677.550 278.400 ;
        RECT 675.750 276.900 682.050 277.800 ;
        RECT 689.250 277.500 690.450 278.400 ;
        RECT 675.750 276.600 677.550 276.900 ;
        RECT 673.950 275.700 674.850 276.600 ;
        RECT 647.700 270.150 648.900 275.400 ;
        RECT 657.450 274.350 660.000 275.400 ;
        RECT 656.100 270.150 657.900 271.950 ;
        RECT 622.950 266.850 625.050 268.950 ;
        RECT 631.950 266.850 634.050 268.950 ;
        RECT 635.100 267.150 636.900 268.950 ;
        RECT 619.950 263.700 621.750 264.600 ;
        RECT 560.550 255.750 562.350 258.600 ;
        RECT 563.850 255.750 565.650 261.600 ;
        RECT 566.850 255.750 568.650 261.600 ;
        RECT 575.850 255.750 577.650 262.800 ;
        RECT 587.250 261.600 588.450 263.700 ;
        RECT 580.350 255.750 582.150 261.600 ;
        RECT 586.650 255.750 588.450 261.600 ;
        RECT 589.650 260.700 597.450 262.050 ;
        RECT 602.250 261.600 603.450 263.700 ;
        RECT 618.450 262.800 621.750 263.700 ;
        RECT 589.650 255.750 591.450 260.700 ;
        RECT 592.650 255.750 594.450 259.800 ;
        RECT 595.650 255.750 597.450 260.700 ;
        RECT 601.650 255.750 603.450 261.600 ;
        RECT 604.650 260.700 612.450 262.050 ;
        RECT 604.650 255.750 606.450 260.700 ;
        RECT 607.650 255.750 609.450 259.800 ;
        RECT 610.650 255.750 612.450 260.700 ;
        RECT 618.450 258.600 619.350 262.800 ;
        RECT 624.000 261.600 625.050 266.850 ;
        RECT 614.550 255.750 616.350 258.600 ;
        RECT 617.550 255.750 619.350 258.600 ;
        RECT 620.550 255.750 622.350 258.600 ;
        RECT 623.550 255.750 625.350 261.600 ;
        RECT 632.400 258.600 633.600 266.850 ;
        RECT 634.950 265.050 637.050 267.150 ;
        RECT 637.950 266.850 640.050 268.950 ;
        RECT 641.100 267.150 642.900 268.950 ;
        RECT 638.100 265.050 639.900 266.850 ;
        RECT 640.950 265.050 643.050 267.150 ;
        RECT 643.950 266.850 646.050 268.950 ;
        RECT 646.950 268.050 649.050 270.150 ;
        RECT 655.950 268.050 658.050 270.150 ;
        RECT 644.100 265.050 645.900 266.850 ;
        RECT 647.700 261.600 648.900 268.050 ;
        RECT 631.650 255.750 633.450 258.600 ;
        RECT 634.650 255.750 636.450 258.600 ;
        RECT 639.000 255.750 640.800 261.600 ;
        RECT 643.200 259.950 648.900 261.600 ;
        RECT 658.950 267.150 660.000 274.350 ;
        RECT 662.100 270.150 663.900 271.950 ;
        RECT 661.950 268.050 664.050 270.150 ;
        RECT 658.950 265.050 661.050 267.150 ;
        RECT 665.550 265.950 666.750 275.400 ;
        RECT 670.950 274.800 673.050 275.700 ;
        RECT 673.950 274.800 679.950 275.700 ;
        RECT 668.850 273.600 673.050 274.800 ;
        RECT 667.950 271.800 669.750 273.600 ;
        RECT 679.050 270.150 679.950 274.800 ;
        RECT 681.150 274.800 682.050 276.900 ;
        RECT 682.950 276.300 690.450 277.500 ;
        RECT 682.950 275.700 684.750 276.300 ;
        RECT 697.050 275.400 698.850 287.250 ;
        RECT 703.650 281.400 705.450 287.250 ;
        RECT 706.650 281.400 708.450 287.250 ;
        RECT 709.650 281.400 711.450 287.250 ;
        RECT 687.750 274.800 698.850 275.400 ;
        RECT 681.150 274.200 698.850 274.800 ;
        RECT 681.150 273.900 689.550 274.200 ;
        RECT 687.750 273.600 689.550 273.900 ;
        RECT 679.050 268.050 682.050 270.150 ;
        RECT 685.950 269.100 688.050 270.150 ;
        RECT 685.950 268.050 693.900 269.100 ;
        RECT 667.950 267.750 670.050 268.050 ;
        RECT 667.950 265.950 671.850 267.750 ;
        RECT 643.200 255.750 645.000 259.950 ;
        RECT 658.950 258.600 660.000 265.050 ;
        RECT 665.550 263.850 670.050 265.950 ;
        RECT 679.050 264.000 679.950 268.050 ;
        RECT 692.100 267.300 693.900 268.050 ;
        RECT 695.100 267.150 696.900 268.950 ;
        RECT 689.100 266.400 690.900 267.000 ;
        RECT 695.100 266.400 696.000 267.150 ;
        RECT 689.100 265.200 696.000 266.400 ;
        RECT 689.100 264.000 690.150 265.200 ;
        RECT 665.550 261.600 666.750 263.850 ;
        RECT 679.050 263.100 690.150 264.000 ;
        RECT 679.050 262.800 679.950 263.100 ;
        RECT 646.500 255.750 648.300 258.600 ;
        RECT 655.650 255.750 657.450 258.600 ;
        RECT 658.650 255.750 660.450 258.600 ;
        RECT 661.650 255.750 663.450 258.600 ;
        RECT 665.550 255.750 667.350 261.600 ;
        RECT 670.950 260.700 673.050 261.600 ;
        RECT 678.150 261.000 679.950 262.800 ;
        RECT 689.100 262.200 690.150 263.100 ;
        RECT 685.350 261.450 687.150 262.200 ;
        RECT 670.950 259.500 674.700 260.700 ;
        RECT 673.650 258.600 674.700 259.500 ;
        RECT 682.200 260.400 687.150 261.450 ;
        RECT 688.650 260.400 690.450 262.200 ;
        RECT 697.950 261.600 698.850 274.200 ;
        RECT 707.250 273.150 708.450 281.400 ;
        RECT 703.950 269.850 706.050 271.950 ;
        RECT 706.950 271.050 709.050 273.150 ;
        RECT 704.100 268.050 705.900 269.850 ;
        RECT 707.250 263.700 708.450 271.050 ;
        RECT 709.950 269.850 712.050 271.950 ;
        RECT 710.100 268.050 711.900 269.850 ;
        RECT 682.200 258.600 683.250 260.400 ;
        RECT 691.950 259.500 694.050 261.600 ;
        RECT 691.950 258.600 693.000 259.500 ;
        RECT 668.850 255.750 670.650 258.600 ;
        RECT 673.350 255.750 675.150 258.600 ;
        RECT 677.550 255.750 679.350 258.600 ;
        RECT 681.450 255.750 683.250 258.600 ;
        RECT 684.750 255.750 686.550 258.600 ;
        RECT 689.250 257.700 693.000 258.600 ;
        RECT 689.250 255.750 691.050 257.700 ;
        RECT 694.050 255.750 695.850 258.600 ;
        RECT 697.050 255.750 698.850 261.600 ;
        RECT 704.850 262.800 708.450 263.700 ;
        RECT 704.850 255.750 706.650 262.800 ;
        RECT 709.350 255.750 711.150 261.600 ;
        RECT 4.650 248.400 6.450 251.250 ;
        RECT 7.650 248.400 9.450 251.250 ;
        RECT 14.700 248.400 16.500 251.250 ;
        RECT 5.400 240.150 6.600 248.400 ;
        RECT 18.000 247.050 19.800 251.250 ;
        RECT 14.100 245.400 19.800 247.050 ;
        RECT 22.200 245.400 24.000 251.250 ;
        RECT 4.950 238.050 7.050 240.150 ;
        RECT 7.950 239.850 10.050 241.950 ;
        RECT 8.100 238.050 9.900 239.850 ;
        RECT 14.100 238.950 15.300 245.400 ;
        RECT 26.700 242.400 28.500 251.250 ;
        RECT 32.100 243.000 33.900 251.250 ;
        RECT 41.850 245.400 43.650 251.250 ;
        RECT 46.350 244.200 48.150 251.250 ;
        RECT 55.650 245.400 57.450 251.250 ;
        RECT 40.950 243.450 43.050 244.050 ;
        RECT 17.100 240.150 18.900 241.950 ;
        RECT 5.400 225.600 6.600 238.050 ;
        RECT 13.950 236.850 16.050 238.950 ;
        RECT 16.950 238.050 19.050 240.150 ;
        RECT 19.950 239.850 22.050 241.950 ;
        RECT 23.100 240.150 24.900 241.950 ;
        RECT 32.100 241.350 36.600 243.000 ;
        RECT 20.100 238.050 21.900 239.850 ;
        RECT 22.950 238.050 25.050 240.150 ;
        RECT 35.400 237.150 36.600 241.350 ;
        RECT 38.550 242.550 43.050 243.450 ;
        RECT 14.100 231.600 15.300 236.850 ;
        RECT 25.950 233.850 28.050 235.950 ;
        RECT 31.950 233.850 34.050 235.950 ;
        RECT 34.950 235.050 37.050 237.150 ;
        RECT 26.100 232.050 27.900 233.850 ;
        RECT 4.650 219.750 6.450 225.600 ;
        RECT 7.650 219.750 9.450 225.600 ;
        RECT 13.650 219.750 15.450 231.600 ;
        RECT 16.650 230.700 24.450 231.600 ;
        RECT 28.950 230.850 31.050 232.950 ;
        RECT 32.250 232.050 34.050 233.850 ;
        RECT 16.650 219.750 18.450 230.700 ;
        RECT 19.650 219.750 21.450 229.800 ;
        RECT 22.650 219.750 24.450 230.700 ;
        RECT 29.100 229.050 30.900 230.850 ;
        RECT 35.700 226.800 36.750 235.050 ;
        RECT 38.550 231.450 39.450 242.550 ;
        RECT 40.950 241.950 43.050 242.550 ;
        RECT 44.550 243.300 48.150 244.200 ;
        RECT 56.250 243.300 57.450 245.400 ;
        RECT 58.650 246.300 60.450 251.250 ;
        RECT 61.650 247.200 63.450 251.250 ;
        RECT 64.650 246.300 66.450 251.250 ;
        RECT 58.650 244.950 66.450 246.300 ;
        RECT 70.350 245.400 72.150 251.250 ;
        RECT 73.350 245.400 75.150 251.250 ;
        RECT 76.650 248.400 78.450 251.250 ;
        RECT 82.650 248.400 84.450 251.250 ;
        RECT 85.650 248.400 87.450 251.250 ;
        RECT 41.100 237.150 42.900 238.950 ;
        RECT 40.950 235.050 43.050 237.150 ;
        RECT 44.550 235.950 45.750 243.300 ;
        RECT 56.250 242.250 60.000 243.300 ;
        RECT 58.950 238.950 60.150 242.250 ;
        RECT 62.100 240.150 63.900 241.950 ;
        RECT 47.100 237.150 48.900 238.950 ;
        RECT 43.950 233.850 46.050 235.950 ;
        RECT 46.950 235.050 49.050 237.150 ;
        RECT 58.950 236.850 61.050 238.950 ;
        RECT 61.950 238.050 64.050 240.150 ;
        RECT 70.650 238.950 71.850 245.400 ;
        RECT 76.650 244.500 77.850 248.400 ;
        RECT 72.750 243.600 77.850 244.500 ;
        RECT 72.750 242.700 75.000 243.600 ;
        RECT 64.950 236.850 67.050 238.950 ;
        RECT 70.650 236.850 73.050 238.950 ;
        RECT 55.950 233.850 58.050 235.950 ;
        RECT 40.950 231.450 43.050 232.050 ;
        RECT 38.550 230.550 43.050 231.450 ;
        RECT 40.950 229.950 43.050 230.550 ;
        RECT 29.700 225.900 36.750 226.800 ;
        RECT 29.700 225.600 31.350 225.900 ;
        RECT 26.550 219.750 28.350 225.600 ;
        RECT 29.550 219.750 31.350 225.600 ;
        RECT 35.550 225.600 36.750 225.900 ;
        RECT 44.550 225.600 45.750 233.850 ;
        RECT 56.250 232.050 58.050 233.850 ;
        RECT 59.850 231.600 61.050 236.850 ;
        RECT 65.100 235.050 66.900 236.850 ;
        RECT 70.650 231.600 71.850 236.850 ;
        RECT 73.950 234.300 75.000 242.700 ;
        RECT 83.400 240.150 84.600 248.400 ;
        RECT 89.700 242.400 91.500 251.250 ;
        RECT 95.100 243.000 96.900 251.250 ;
        RECT 105.000 245.400 106.800 251.250 ;
        RECT 109.200 247.050 111.000 251.250 ;
        RECT 112.500 248.400 114.300 251.250 ;
        RECT 109.200 245.400 114.900 247.050 ;
        RECT 76.950 236.850 79.050 238.950 ;
        RECT 82.950 238.050 85.050 240.150 ;
        RECT 85.950 239.850 88.050 241.950 ;
        RECT 95.100 241.350 99.600 243.000 ;
        RECT 86.100 238.050 87.900 239.850 ;
        RECT 77.100 235.050 78.900 236.850 ;
        RECT 72.750 233.400 75.000 234.300 ;
        RECT 72.750 232.500 78.450 233.400 ;
        RECT 32.550 219.750 34.350 225.000 ;
        RECT 35.550 219.750 37.350 225.600 ;
        RECT 41.550 219.750 43.350 225.600 ;
        RECT 44.550 219.750 46.350 225.600 ;
        RECT 47.550 219.750 49.350 225.600 ;
        RECT 56.400 219.750 58.200 225.600 ;
        RECT 59.700 219.750 61.500 231.600 ;
        RECT 63.900 219.750 65.700 231.600 ;
        RECT 70.350 219.750 72.150 231.600 ;
        RECT 73.350 219.750 75.150 231.600 ;
        RECT 77.250 225.600 78.450 232.500 ;
        RECT 83.400 225.600 84.600 238.050 ;
        RECT 98.400 237.150 99.600 241.350 ;
        RECT 104.100 240.150 105.900 241.950 ;
        RECT 103.950 238.050 106.050 240.150 ;
        RECT 106.950 239.850 109.050 241.950 ;
        RECT 110.100 240.150 111.900 241.950 ;
        RECT 107.100 238.050 108.900 239.850 ;
        RECT 109.950 238.050 112.050 240.150 ;
        RECT 113.700 238.950 114.900 245.400 ;
        RECT 119.700 242.400 121.500 251.250 ;
        RECT 125.100 243.000 126.900 251.250 ;
        RECT 135.000 245.400 136.800 251.250 ;
        RECT 139.200 247.050 141.000 251.250 ;
        RECT 142.500 248.400 144.300 251.250 ;
        RECT 139.200 245.400 144.900 247.050 ;
        RECT 125.100 241.350 129.600 243.000 ;
        RECT 88.950 233.850 91.050 235.950 ;
        RECT 94.950 233.850 97.050 235.950 ;
        RECT 97.950 235.050 100.050 237.150 ;
        RECT 112.950 236.850 115.050 238.950 ;
        RECT 128.400 237.150 129.600 241.350 ;
        RECT 134.100 240.150 135.900 241.950 ;
        RECT 133.950 238.050 136.050 240.150 ;
        RECT 136.950 239.850 139.050 241.950 ;
        RECT 140.100 240.150 141.900 241.950 ;
        RECT 137.100 238.050 138.900 239.850 ;
        RECT 139.950 238.050 142.050 240.150 ;
        RECT 143.700 238.950 144.900 245.400 ;
        RECT 149.700 242.400 151.500 251.250 ;
        RECT 155.100 243.000 156.900 251.250 ;
        RECT 166.650 245.400 168.450 251.250 ;
        RECT 155.100 241.350 159.600 243.000 ;
        RECT 160.950 241.950 163.050 244.050 ;
        RECT 167.250 243.300 168.450 245.400 ;
        RECT 169.650 246.300 171.450 251.250 ;
        RECT 172.650 247.200 174.450 251.250 ;
        RECT 175.650 246.300 177.450 251.250 ;
        RECT 169.650 244.950 177.450 246.300 ;
        RECT 167.250 242.250 171.000 243.300 ;
        RECT 179.700 242.400 181.500 251.250 ;
        RECT 185.100 243.000 186.900 251.250 ;
        RECT 187.950 246.450 190.050 247.050 ;
        RECT 187.950 245.550 192.450 246.450 ;
        RECT 187.950 244.950 190.050 245.550 ;
        RECT 89.100 232.050 90.900 233.850 ;
        RECT 91.950 230.850 94.050 232.950 ;
        RECT 95.250 232.050 97.050 233.850 ;
        RECT 92.100 229.050 93.900 230.850 ;
        RECT 98.700 226.800 99.750 235.050 ;
        RECT 113.700 231.600 114.900 236.850 ;
        RECT 118.950 233.850 121.050 235.950 ;
        RECT 124.950 233.850 127.050 235.950 ;
        RECT 127.950 235.050 130.050 237.150 ;
        RECT 142.950 236.850 145.050 238.950 ;
        RECT 158.400 237.150 159.600 241.350 ;
        RECT 119.100 232.050 120.900 233.850 ;
        RECT 92.700 225.900 99.750 226.800 ;
        RECT 92.700 225.600 94.350 225.900 ;
        RECT 76.650 219.750 78.450 225.600 ;
        RECT 82.650 219.750 84.450 225.600 ;
        RECT 85.650 219.750 87.450 225.600 ;
        RECT 89.550 219.750 91.350 225.600 ;
        RECT 92.550 219.750 94.350 225.600 ;
        RECT 98.550 225.600 99.750 225.900 ;
        RECT 104.550 230.700 112.350 231.600 ;
        RECT 95.550 219.750 97.350 225.000 ;
        RECT 98.550 219.750 100.350 225.600 ;
        RECT 104.550 219.750 106.350 230.700 ;
        RECT 107.550 219.750 109.350 229.800 ;
        RECT 110.550 219.750 112.350 230.700 ;
        RECT 113.550 219.750 115.350 231.600 ;
        RECT 121.950 230.850 124.050 232.950 ;
        RECT 125.250 232.050 127.050 233.850 ;
        RECT 122.100 229.050 123.900 230.850 ;
        RECT 128.700 226.800 129.750 235.050 ;
        RECT 143.700 231.600 144.900 236.850 ;
        RECT 148.950 233.850 151.050 235.950 ;
        RECT 154.950 233.850 157.050 235.950 ;
        RECT 157.950 235.050 160.050 237.150 ;
        RECT 149.100 232.050 150.900 233.850 ;
        RECT 122.700 225.900 129.750 226.800 ;
        RECT 122.700 225.600 124.350 225.900 ;
        RECT 119.550 219.750 121.350 225.600 ;
        RECT 122.550 219.750 124.350 225.600 ;
        RECT 128.550 225.600 129.750 225.900 ;
        RECT 134.550 230.700 142.350 231.600 ;
        RECT 125.550 219.750 127.350 225.000 ;
        RECT 128.550 219.750 130.350 225.600 ;
        RECT 134.550 219.750 136.350 230.700 ;
        RECT 137.550 219.750 139.350 229.800 ;
        RECT 140.550 219.750 142.350 230.700 ;
        RECT 143.550 219.750 145.350 231.600 ;
        RECT 151.950 230.850 154.050 232.950 ;
        RECT 155.250 232.050 157.050 233.850 ;
        RECT 152.100 229.050 153.900 230.850 ;
        RECT 158.700 226.800 159.750 235.050 ;
        RECT 161.550 231.450 162.450 241.950 ;
        RECT 169.950 238.950 171.150 242.250 ;
        RECT 173.100 240.150 174.900 241.950 ;
        RECT 185.100 241.350 189.600 243.000 ;
        RECT 169.950 236.850 172.050 238.950 ;
        RECT 172.950 238.050 175.050 240.150 ;
        RECT 175.950 236.850 178.050 238.950 ;
        RECT 188.400 237.150 189.600 241.350 ;
        RECT 166.950 233.850 169.050 235.950 ;
        RECT 167.250 232.050 169.050 233.850 ;
        RECT 163.950 231.450 166.050 232.050 ;
        RECT 170.850 231.600 172.050 236.850 ;
        RECT 176.100 235.050 177.900 236.850 ;
        RECT 178.950 233.850 181.050 235.950 ;
        RECT 184.950 233.850 187.050 235.950 ;
        RECT 187.950 235.050 190.050 237.150 ;
        RECT 179.100 232.050 180.900 233.850 ;
        RECT 161.550 230.550 166.050 231.450 ;
        RECT 163.950 229.950 166.050 230.550 ;
        RECT 152.700 225.900 159.750 226.800 ;
        RECT 152.700 225.600 154.350 225.900 ;
        RECT 149.550 219.750 151.350 225.600 ;
        RECT 152.550 219.750 154.350 225.600 ;
        RECT 158.550 225.600 159.750 225.900 ;
        RECT 155.550 219.750 157.350 225.000 ;
        RECT 158.550 219.750 160.350 225.600 ;
        RECT 167.400 219.750 169.200 225.600 ;
        RECT 170.700 219.750 172.500 231.600 ;
        RECT 174.900 219.750 176.700 231.600 ;
        RECT 181.950 230.850 184.050 232.950 ;
        RECT 185.250 232.050 187.050 233.850 ;
        RECT 182.100 229.050 183.900 230.850 ;
        RECT 188.700 226.800 189.750 235.050 ;
        RECT 191.550 234.450 192.450 245.550 ;
        RECT 195.000 245.400 196.800 251.250 ;
        RECT 199.200 247.050 201.000 251.250 ;
        RECT 202.500 248.400 204.300 251.250 ;
        RECT 211.650 248.400 213.450 251.250 ;
        RECT 214.650 248.400 216.450 251.250 ;
        RECT 199.200 245.400 204.900 247.050 ;
        RECT 194.100 240.150 195.900 241.950 ;
        RECT 193.950 238.050 196.050 240.150 ;
        RECT 196.950 239.850 199.050 241.950 ;
        RECT 200.100 240.150 201.900 241.950 ;
        RECT 197.100 238.050 198.900 239.850 ;
        RECT 199.950 238.050 202.050 240.150 ;
        RECT 203.700 238.950 204.900 245.400 ;
        RECT 212.400 240.150 213.600 248.400 ;
        RECT 218.700 242.400 220.500 251.250 ;
        RECT 224.100 243.000 225.900 251.250 ;
        RECT 234.000 245.400 235.800 251.250 ;
        RECT 238.200 247.050 240.000 251.250 ;
        RECT 241.500 248.400 243.300 251.250 ;
        RECT 238.200 245.400 243.900 247.050 ;
        RECT 202.950 236.850 205.050 238.950 ;
        RECT 211.950 238.050 214.050 240.150 ;
        RECT 214.950 239.850 217.050 241.950 ;
        RECT 224.100 241.350 228.600 243.000 ;
        RECT 215.100 238.050 216.900 239.850 ;
        RECT 193.950 234.450 196.050 235.050 ;
        RECT 191.550 233.550 196.050 234.450 ;
        RECT 193.950 232.950 196.050 233.550 ;
        RECT 203.700 231.600 204.900 236.850 ;
        RECT 182.700 225.900 189.750 226.800 ;
        RECT 182.700 225.600 184.350 225.900 ;
        RECT 179.550 219.750 181.350 225.600 ;
        RECT 182.550 219.750 184.350 225.600 ;
        RECT 188.550 225.600 189.750 225.900 ;
        RECT 194.550 230.700 202.350 231.600 ;
        RECT 185.550 219.750 187.350 225.000 ;
        RECT 188.550 219.750 190.350 225.600 ;
        RECT 194.550 219.750 196.350 230.700 ;
        RECT 197.550 219.750 199.350 229.800 ;
        RECT 200.550 219.750 202.350 230.700 ;
        RECT 203.550 219.750 205.350 231.600 ;
        RECT 212.400 225.600 213.600 238.050 ;
        RECT 227.400 237.150 228.600 241.350 ;
        RECT 233.100 240.150 234.900 241.950 ;
        RECT 232.950 238.050 235.050 240.150 ;
        RECT 235.950 239.850 238.050 241.950 ;
        RECT 239.100 240.150 240.900 241.950 ;
        RECT 236.100 238.050 237.900 239.850 ;
        RECT 238.950 238.050 241.050 240.150 ;
        RECT 242.700 238.950 243.900 245.400 ;
        RECT 248.700 242.400 250.500 251.250 ;
        RECT 254.100 243.000 255.900 251.250 ;
        RECT 263.550 246.300 265.350 251.250 ;
        RECT 266.550 247.200 268.350 251.250 ;
        RECT 269.550 246.300 271.350 251.250 ;
        RECT 263.550 244.950 271.350 246.300 ;
        RECT 272.550 245.400 274.350 251.250 ;
        RECT 281.700 248.400 283.500 251.250 ;
        RECT 285.000 247.050 286.800 251.250 ;
        RECT 281.100 245.400 286.800 247.050 ;
        RECT 289.200 245.400 291.000 251.250 ;
        RECT 293.550 248.400 295.350 251.250 ;
        RECT 296.550 248.400 298.350 251.250 ;
        RECT 272.550 243.300 273.750 245.400 ;
        RECT 254.100 241.350 258.600 243.000 ;
        RECT 270.000 242.250 273.750 243.300 ;
        RECT 217.950 233.850 220.050 235.950 ;
        RECT 223.950 233.850 226.050 235.950 ;
        RECT 226.950 235.050 229.050 237.150 ;
        RECT 241.950 236.850 244.050 238.950 ;
        RECT 257.400 237.150 258.600 241.350 ;
        RECT 266.100 240.150 267.900 241.950 ;
        RECT 218.100 232.050 219.900 233.850 ;
        RECT 220.950 230.850 223.050 232.950 ;
        RECT 224.250 232.050 226.050 233.850 ;
        RECT 221.100 229.050 222.900 230.850 ;
        RECT 227.700 226.800 228.750 235.050 ;
        RECT 242.700 231.600 243.900 236.850 ;
        RECT 247.950 233.850 250.050 235.950 ;
        RECT 253.950 233.850 256.050 235.950 ;
        RECT 256.950 235.050 259.050 237.150 ;
        RECT 262.950 236.850 265.050 238.950 ;
        RECT 265.950 238.050 268.050 240.150 ;
        RECT 269.850 238.950 271.050 242.250 ;
        RECT 281.100 238.950 282.300 245.400 ;
        RECT 284.100 240.150 285.900 241.950 ;
        RECT 268.950 236.850 271.050 238.950 ;
        RECT 280.950 236.850 283.050 238.950 ;
        RECT 283.950 238.050 286.050 240.150 ;
        RECT 286.950 239.850 289.050 241.950 ;
        RECT 290.100 240.150 291.900 241.950 ;
        RECT 287.100 238.050 288.900 239.850 ;
        RECT 289.950 238.050 292.050 240.150 ;
        RECT 292.950 239.850 295.050 241.950 ;
        RECT 296.400 240.150 297.600 248.400 ;
        RECT 302.700 242.400 304.500 251.250 ;
        RECT 308.100 243.000 309.900 251.250 ;
        RECT 319.650 245.400 321.450 251.250 ;
        RECT 320.250 243.300 321.450 245.400 ;
        RECT 322.650 246.300 324.450 251.250 ;
        RECT 325.650 247.200 327.450 251.250 ;
        RECT 328.650 246.300 330.450 251.250 ;
        RECT 332.550 248.400 334.350 251.250 ;
        RECT 335.550 248.400 337.350 251.250 ;
        RECT 322.650 244.950 330.450 246.300 ;
        RECT 308.100 241.350 312.600 243.000 ;
        RECT 320.250 242.250 324.000 243.300 ;
        RECT 304.950 240.450 307.050 241.050 ;
        RECT 293.100 238.050 294.900 239.850 ;
        RECT 295.950 238.050 298.050 240.150 ;
        RECT 299.550 239.550 307.050 240.450 ;
        RECT 263.100 235.050 264.900 236.850 ;
        RECT 248.100 232.050 249.900 233.850 ;
        RECT 221.700 225.900 228.750 226.800 ;
        RECT 221.700 225.600 223.350 225.900 ;
        RECT 211.650 219.750 213.450 225.600 ;
        RECT 214.650 219.750 216.450 225.600 ;
        RECT 218.550 219.750 220.350 225.600 ;
        RECT 221.550 219.750 223.350 225.600 ;
        RECT 227.550 225.600 228.750 225.900 ;
        RECT 233.550 230.700 241.350 231.600 ;
        RECT 224.550 219.750 226.350 225.000 ;
        RECT 227.550 219.750 229.350 225.600 ;
        RECT 233.550 219.750 235.350 230.700 ;
        RECT 236.550 219.750 238.350 229.800 ;
        RECT 239.550 219.750 241.350 230.700 ;
        RECT 242.550 219.750 244.350 231.600 ;
        RECT 250.950 230.850 253.050 232.950 ;
        RECT 254.250 232.050 256.050 233.850 ;
        RECT 251.100 229.050 252.900 230.850 ;
        RECT 257.700 226.800 258.750 235.050 ;
        RECT 268.950 231.600 270.150 236.850 ;
        RECT 271.950 233.850 274.050 235.950 ;
        RECT 271.950 232.050 273.750 233.850 ;
        RECT 281.100 231.600 282.300 236.850 ;
        RECT 251.700 225.900 258.750 226.800 ;
        RECT 251.700 225.600 253.350 225.900 ;
        RECT 248.550 219.750 250.350 225.600 ;
        RECT 251.550 219.750 253.350 225.600 ;
        RECT 257.550 225.600 258.750 225.900 ;
        RECT 254.550 219.750 256.350 225.000 ;
        RECT 257.550 219.750 259.350 225.600 ;
        RECT 264.300 219.750 266.100 231.600 ;
        RECT 268.500 219.750 270.300 231.600 ;
        RECT 271.800 219.750 273.600 225.600 ;
        RECT 280.650 219.750 282.450 231.600 ;
        RECT 283.650 230.700 291.450 231.600 ;
        RECT 283.650 219.750 285.450 230.700 ;
        RECT 286.650 219.750 288.450 229.800 ;
        RECT 289.650 219.750 291.450 230.700 ;
        RECT 296.400 225.600 297.600 238.050 ;
        RECT 299.550 232.050 300.450 239.550 ;
        RECT 304.950 238.950 307.050 239.550 ;
        RECT 311.400 237.150 312.600 241.350 ;
        RECT 319.950 240.450 322.050 241.050 ;
        RECT 317.550 239.550 322.050 240.450 ;
        RECT 301.950 233.850 304.050 235.950 ;
        RECT 307.950 233.850 310.050 235.950 ;
        RECT 310.950 235.050 313.050 237.150 ;
        RECT 302.100 232.050 303.900 233.850 ;
        RECT 298.950 229.950 301.050 232.050 ;
        RECT 304.950 230.850 307.050 232.950 ;
        RECT 308.250 232.050 310.050 233.850 ;
        RECT 305.100 229.050 306.900 230.850 ;
        RECT 311.700 226.800 312.750 235.050 ;
        RECT 313.950 231.450 316.050 232.050 ;
        RECT 317.550 231.450 318.450 239.550 ;
        RECT 319.950 238.950 322.050 239.550 ;
        RECT 322.950 238.950 324.150 242.250 ;
        RECT 326.100 240.150 327.900 241.950 ;
        RECT 322.950 236.850 325.050 238.950 ;
        RECT 325.950 238.050 328.050 240.150 ;
        RECT 331.950 239.850 334.050 241.950 ;
        RECT 335.400 240.150 336.600 248.400 ;
        RECT 341.550 245.400 343.350 251.250 ;
        RECT 344.850 248.400 346.650 251.250 ;
        RECT 349.350 248.400 351.150 251.250 ;
        RECT 353.550 248.400 355.350 251.250 ;
        RECT 357.450 248.400 359.250 251.250 ;
        RECT 360.750 248.400 362.550 251.250 ;
        RECT 365.250 249.300 367.050 251.250 ;
        RECT 365.250 248.400 369.000 249.300 ;
        RECT 370.050 248.400 371.850 251.250 ;
        RECT 349.650 247.500 350.700 248.400 ;
        RECT 346.950 246.300 350.700 247.500 ;
        RECT 358.200 246.600 359.250 248.400 ;
        RECT 367.950 247.500 369.000 248.400 ;
        RECT 346.950 245.400 349.050 246.300 ;
        RECT 341.550 243.150 342.750 245.400 ;
        RECT 354.150 244.200 355.950 246.000 ;
        RECT 358.200 245.550 363.150 246.600 ;
        RECT 361.350 244.800 363.150 245.550 ;
        RECT 364.650 244.800 366.450 246.600 ;
        RECT 367.950 245.400 370.050 247.500 ;
        RECT 373.050 245.400 374.850 251.250 ;
        RECT 379.650 245.400 381.450 251.250 ;
        RECT 355.050 243.900 355.950 244.200 ;
        RECT 365.100 243.900 366.150 244.800 ;
        RECT 341.550 241.050 346.050 243.150 ;
        RECT 355.050 243.000 366.150 243.900 ;
        RECT 328.950 236.850 331.050 238.950 ;
        RECT 332.100 238.050 333.900 239.850 ;
        RECT 334.950 238.050 337.050 240.150 ;
        RECT 319.950 233.850 322.050 235.950 ;
        RECT 320.250 232.050 322.050 233.850 ;
        RECT 323.850 231.600 325.050 236.850 ;
        RECT 329.100 235.050 330.900 236.850 ;
        RECT 313.950 230.550 318.450 231.450 ;
        RECT 313.950 229.950 316.050 230.550 ;
        RECT 305.700 225.900 312.750 226.800 ;
        RECT 305.700 225.600 307.350 225.900 ;
        RECT 293.550 219.750 295.350 225.600 ;
        RECT 296.550 219.750 298.350 225.600 ;
        RECT 302.550 219.750 304.350 225.600 ;
        RECT 305.550 219.750 307.350 225.600 ;
        RECT 311.550 225.600 312.750 225.900 ;
        RECT 308.550 219.750 310.350 225.000 ;
        RECT 311.550 219.750 313.350 225.600 ;
        RECT 320.400 219.750 322.200 225.600 ;
        RECT 323.700 219.750 325.500 231.600 ;
        RECT 327.900 219.750 329.700 231.600 ;
        RECT 335.400 225.600 336.600 238.050 ;
        RECT 341.550 231.600 342.750 241.050 ;
        RECT 343.950 239.250 347.850 241.050 ;
        RECT 343.950 238.950 346.050 239.250 ;
        RECT 355.050 238.950 355.950 243.000 ;
        RECT 365.100 241.800 366.150 243.000 ;
        RECT 365.100 240.600 372.000 241.800 ;
        RECT 365.100 240.000 366.900 240.600 ;
        RECT 371.100 239.850 372.000 240.600 ;
        RECT 368.100 238.950 369.900 239.700 ;
        RECT 355.050 236.850 358.050 238.950 ;
        RECT 361.950 237.900 369.900 238.950 ;
        RECT 371.100 238.050 372.900 239.850 ;
        RECT 361.950 236.850 364.050 237.900 ;
        RECT 343.950 233.400 345.750 235.200 ;
        RECT 344.850 232.200 349.050 233.400 ;
        RECT 355.050 232.200 355.950 236.850 ;
        RECT 363.750 233.100 365.550 233.400 ;
        RECT 332.550 219.750 334.350 225.600 ;
        RECT 335.550 219.750 337.350 225.600 ;
        RECT 341.550 219.750 343.350 231.600 ;
        RECT 346.950 231.300 349.050 232.200 ;
        RECT 349.950 231.300 355.950 232.200 ;
        RECT 357.150 232.800 365.550 233.100 ;
        RECT 373.950 232.800 374.850 245.400 ;
        RECT 380.250 243.300 381.450 245.400 ;
        RECT 382.650 246.300 384.450 251.250 ;
        RECT 385.650 247.200 387.450 251.250 ;
        RECT 388.650 246.300 390.450 251.250 ;
        RECT 396.150 246.900 397.950 251.250 ;
        RECT 382.650 244.950 390.450 246.300 ;
        RECT 394.650 245.400 397.950 246.900 ;
        RECT 399.150 245.400 400.950 251.250 ;
        RECT 380.250 242.250 384.000 243.300 ;
        RECT 382.950 238.950 384.150 242.250 ;
        RECT 386.100 240.150 387.900 241.950 ;
        RECT 382.950 236.850 385.050 238.950 ;
        RECT 385.950 238.050 388.050 240.150 ;
        RECT 394.650 238.950 395.850 245.400 ;
        RECT 397.950 243.900 399.750 244.500 ;
        RECT 403.650 243.900 405.450 251.250 ;
        RECT 407.550 248.400 409.350 251.250 ;
        RECT 410.550 248.400 412.350 251.250 ;
        RECT 413.550 248.400 415.350 251.250 ;
        RECT 397.950 242.700 405.450 243.900 ;
        RECT 388.950 236.850 391.050 238.950 ;
        RECT 394.650 236.850 397.050 238.950 ;
        RECT 398.100 237.150 399.900 238.950 ;
        RECT 379.950 233.850 382.050 235.950 ;
        RECT 357.150 232.200 374.850 232.800 ;
        RECT 349.950 230.400 350.850 231.300 ;
        RECT 348.150 228.600 350.850 230.400 ;
        RECT 351.750 230.100 353.550 230.400 ;
        RECT 357.150 230.100 358.050 232.200 ;
        RECT 363.750 231.600 374.850 232.200 ;
        RECT 380.250 232.050 382.050 233.850 ;
        RECT 383.850 231.600 385.050 236.850 ;
        RECT 389.100 235.050 390.900 236.850 ;
        RECT 394.650 231.600 395.850 236.850 ;
        RECT 397.950 235.050 400.050 237.150 ;
        RECT 351.750 229.200 358.050 230.100 ;
        RECT 358.950 230.700 360.750 231.300 ;
        RECT 358.950 229.500 366.450 230.700 ;
        RECT 351.750 228.600 353.550 229.200 ;
        RECT 365.250 228.600 366.450 229.500 ;
        RECT 346.950 225.600 350.850 227.700 ;
        RECT 355.950 226.500 362.850 228.300 ;
        RECT 365.250 226.500 370.050 228.600 ;
        RECT 344.550 219.750 346.350 222.600 ;
        RECT 349.050 219.750 350.850 225.600 ;
        RECT 353.250 219.750 355.050 225.600 ;
        RECT 357.150 219.750 358.950 226.500 ;
        RECT 365.250 225.600 366.450 226.500 ;
        RECT 360.150 219.750 361.950 225.600 ;
        RECT 364.950 219.750 366.750 225.600 ;
        RECT 370.050 219.750 371.850 225.600 ;
        RECT 373.050 219.750 374.850 231.600 ;
        RECT 380.400 219.750 382.200 225.600 ;
        RECT 383.700 219.750 385.500 231.600 ;
        RECT 387.900 219.750 389.700 231.600 ;
        RECT 394.050 219.750 395.850 231.600 ;
        RECT 397.050 219.750 398.850 231.600 ;
        RECT 401.100 225.600 402.300 242.700 ;
        RECT 411.000 241.950 412.050 248.400 ;
        RECT 420.000 245.400 421.800 251.250 ;
        RECT 424.200 247.050 426.000 251.250 ;
        RECT 427.500 248.400 429.300 251.250 ;
        RECT 436.650 248.400 438.450 251.250 ;
        RECT 439.650 248.400 441.450 251.250 ;
        RECT 442.650 248.400 444.450 251.250 ;
        RECT 448.650 248.400 450.450 251.250 ;
        RECT 451.650 248.400 453.450 251.250 ;
        RECT 457.650 248.400 459.450 251.250 ;
        RECT 460.650 248.400 462.450 251.250 ;
        RECT 424.200 245.400 429.900 247.050 ;
        RECT 409.950 239.850 412.050 241.950 ;
        RECT 419.100 240.150 420.900 241.950 ;
        RECT 403.950 236.850 406.050 238.950 ;
        RECT 406.950 236.850 409.050 238.950 ;
        RECT 404.100 235.050 405.900 236.850 ;
        RECT 407.100 235.050 408.900 236.850 ;
        RECT 411.000 232.650 412.050 239.850 ;
        RECT 412.950 236.850 415.050 238.950 ;
        RECT 418.950 238.050 421.050 240.150 ;
        RECT 421.950 239.850 424.050 241.950 ;
        RECT 425.100 240.150 426.900 241.950 ;
        RECT 422.100 238.050 423.900 239.850 ;
        RECT 424.950 238.050 427.050 240.150 ;
        RECT 428.700 238.950 429.900 245.400 ;
        RECT 439.950 241.950 441.000 248.400 ;
        RECT 439.950 239.850 442.050 241.950 ;
        RECT 449.400 240.150 450.600 248.400 ;
        RECT 427.950 236.850 430.050 238.950 ;
        RECT 436.950 236.850 439.050 238.950 ;
        RECT 413.100 235.050 414.900 236.850 ;
        RECT 411.000 231.600 413.550 232.650 ;
        RECT 428.700 231.600 429.900 236.850 ;
        RECT 437.100 235.050 438.900 236.850 ;
        RECT 439.950 232.650 441.000 239.850 ;
        RECT 442.950 236.850 445.050 238.950 ;
        RECT 448.950 238.050 451.050 240.150 ;
        RECT 451.950 239.850 454.050 241.950 ;
        RECT 458.400 240.150 459.600 248.400 ;
        RECT 464.550 246.300 466.350 251.250 ;
        RECT 467.550 247.200 469.350 251.250 ;
        RECT 470.550 246.300 472.350 251.250 ;
        RECT 464.550 244.950 472.350 246.300 ;
        RECT 473.550 245.400 475.350 251.250 ;
        RECT 479.850 245.400 481.650 251.250 ;
        RECT 473.550 243.300 474.750 245.400 ;
        RECT 484.350 244.200 486.150 251.250 ;
        RECT 471.000 242.250 474.750 243.300 ;
        RECT 482.550 243.300 486.150 244.200 ;
        RECT 494.850 244.200 496.650 251.250 ;
        RECT 499.350 245.400 501.150 251.250 ;
        RECT 505.650 245.400 507.450 251.250 ;
        RECT 494.850 243.300 498.450 244.200 ;
        RECT 452.100 238.050 453.900 239.850 ;
        RECT 457.950 238.050 460.050 240.150 ;
        RECT 460.950 239.850 463.050 241.950 ;
        RECT 467.100 240.150 468.900 241.950 ;
        RECT 461.100 238.050 462.900 239.850 ;
        RECT 443.100 235.050 444.900 236.850 ;
        RECT 438.450 231.600 441.000 232.650 ;
        RECT 400.650 219.750 402.450 225.600 ;
        RECT 403.650 219.750 405.450 225.600 ;
        RECT 407.550 219.750 409.350 231.600 ;
        RECT 411.750 219.750 413.550 231.600 ;
        RECT 419.550 230.700 427.350 231.600 ;
        RECT 419.550 219.750 421.350 230.700 ;
        RECT 422.550 219.750 424.350 229.800 ;
        RECT 425.550 219.750 427.350 230.700 ;
        RECT 428.550 219.750 430.350 231.600 ;
        RECT 438.450 219.750 440.250 231.600 ;
        RECT 442.650 219.750 444.450 231.600 ;
        RECT 449.400 225.600 450.600 238.050 ;
        RECT 458.400 225.600 459.600 238.050 ;
        RECT 463.950 236.850 466.050 238.950 ;
        RECT 466.950 238.050 469.050 240.150 ;
        RECT 470.850 238.950 472.050 242.250 ;
        RECT 469.950 236.850 472.050 238.950 ;
        RECT 479.100 237.150 480.900 238.950 ;
        RECT 464.100 235.050 465.900 236.850 ;
        RECT 469.950 231.600 471.150 236.850 ;
        RECT 472.950 233.850 475.050 235.950 ;
        RECT 478.950 235.050 481.050 237.150 ;
        RECT 482.550 235.950 483.750 243.300 ;
        RECT 485.100 237.150 486.900 238.950 ;
        RECT 494.100 237.150 495.900 238.950 ;
        RECT 481.950 233.850 484.050 235.950 ;
        RECT 484.950 235.050 487.050 237.150 ;
        RECT 493.950 235.050 496.050 237.150 ;
        RECT 497.250 235.950 498.450 243.300 ;
        RECT 506.250 243.300 507.450 245.400 ;
        RECT 508.650 246.300 510.450 251.250 ;
        RECT 511.650 247.200 513.450 251.250 ;
        RECT 514.650 246.300 516.450 251.250 ;
        RECT 508.650 244.950 516.450 246.300 ;
        RECT 519.150 245.400 520.950 251.250 ;
        RECT 522.150 248.400 523.950 251.250 ;
        RECT 526.950 249.300 528.750 251.250 ;
        RECT 525.000 248.400 528.750 249.300 ;
        RECT 531.450 248.400 533.250 251.250 ;
        RECT 534.750 248.400 536.550 251.250 ;
        RECT 538.650 248.400 540.450 251.250 ;
        RECT 542.850 248.400 544.650 251.250 ;
        RECT 547.350 248.400 549.150 251.250 ;
        RECT 525.000 247.500 526.050 248.400 ;
        RECT 523.950 245.400 526.050 247.500 ;
        RECT 534.750 246.600 535.800 248.400 ;
        RECT 506.250 242.250 510.000 243.300 ;
        RECT 505.950 240.450 508.050 241.050 ;
        RECT 503.550 239.550 508.050 240.450 ;
        RECT 500.100 237.150 501.900 238.950 ;
        RECT 496.950 233.850 499.050 235.950 ;
        RECT 499.950 235.050 502.050 237.150 ;
        RECT 472.950 232.050 474.750 233.850 ;
        RECT 448.650 219.750 450.450 225.600 ;
        RECT 451.650 219.750 453.450 225.600 ;
        RECT 457.650 219.750 459.450 225.600 ;
        RECT 460.650 219.750 462.450 225.600 ;
        RECT 465.300 219.750 467.100 231.600 ;
        RECT 469.500 219.750 471.300 231.600 ;
        RECT 482.550 225.600 483.750 233.850 ;
        RECT 497.250 225.600 498.450 233.850 ;
        RECT 503.550 228.450 504.450 239.550 ;
        RECT 505.950 238.950 508.050 239.550 ;
        RECT 508.950 238.950 510.150 242.250 ;
        RECT 512.100 240.150 513.900 241.950 ;
        RECT 508.950 236.850 511.050 238.950 ;
        RECT 511.950 238.050 514.050 240.150 ;
        RECT 514.950 236.850 517.050 238.950 ;
        RECT 505.950 233.850 508.050 235.950 ;
        RECT 506.250 232.050 508.050 233.850 ;
        RECT 509.850 231.600 511.050 236.850 ;
        RECT 515.100 235.050 516.900 236.850 ;
        RECT 519.150 232.800 520.050 245.400 ;
        RECT 527.550 244.800 529.350 246.600 ;
        RECT 530.850 245.550 535.800 246.600 ;
        RECT 543.300 247.500 544.350 248.400 ;
        RECT 543.300 246.300 547.050 247.500 ;
        RECT 530.850 244.800 532.650 245.550 ;
        RECT 527.850 243.900 528.900 244.800 ;
        RECT 538.050 244.200 539.850 246.000 ;
        RECT 544.950 245.400 547.050 246.300 ;
        RECT 550.650 245.400 552.450 251.250 ;
        RECT 554.550 248.400 556.350 251.250 ;
        RECT 557.550 248.400 559.350 251.250 ;
        RECT 565.650 248.400 567.450 251.250 ;
        RECT 568.650 248.400 570.450 251.250 ;
        RECT 538.050 243.900 538.950 244.200 ;
        RECT 527.850 243.000 538.950 243.900 ;
        RECT 551.250 243.150 552.450 245.400 ;
        RECT 527.850 241.800 528.900 243.000 ;
        RECT 522.000 240.600 528.900 241.800 ;
        RECT 522.000 239.850 522.900 240.600 ;
        RECT 527.100 240.000 528.900 240.600 ;
        RECT 521.100 238.050 522.900 239.850 ;
        RECT 524.100 238.950 525.900 239.700 ;
        RECT 538.050 238.950 538.950 243.000 ;
        RECT 547.950 241.050 552.450 243.150 ;
        RECT 546.150 239.250 550.050 241.050 ;
        RECT 547.950 238.950 550.050 239.250 ;
        RECT 524.100 237.900 532.050 238.950 ;
        RECT 529.950 236.850 532.050 237.900 ;
        RECT 535.950 236.850 538.950 238.950 ;
        RECT 528.450 233.100 530.250 233.400 ;
        RECT 528.450 232.800 536.850 233.100 ;
        RECT 519.150 232.200 536.850 232.800 ;
        RECT 519.150 231.600 530.250 232.200 ;
        RECT 505.950 228.450 508.050 229.050 ;
        RECT 503.550 227.550 508.050 228.450 ;
        RECT 505.950 226.950 508.050 227.550 ;
        RECT 472.800 219.750 474.600 225.600 ;
        RECT 479.550 219.750 481.350 225.600 ;
        RECT 482.550 219.750 484.350 225.600 ;
        RECT 485.550 219.750 487.350 225.600 ;
        RECT 493.650 219.750 495.450 225.600 ;
        RECT 496.650 219.750 498.450 225.600 ;
        RECT 499.650 219.750 501.450 225.600 ;
        RECT 506.400 219.750 508.200 225.600 ;
        RECT 509.700 219.750 511.500 231.600 ;
        RECT 513.900 219.750 515.700 231.600 ;
        RECT 519.150 219.750 520.950 231.600 ;
        RECT 533.250 230.700 535.050 231.300 ;
        RECT 527.550 229.500 535.050 230.700 ;
        RECT 535.950 230.100 536.850 232.200 ;
        RECT 538.050 232.200 538.950 236.850 ;
        RECT 548.250 233.400 550.050 235.200 ;
        RECT 544.950 232.200 549.150 233.400 ;
        RECT 538.050 231.300 544.050 232.200 ;
        RECT 544.950 231.300 547.050 232.200 ;
        RECT 551.250 231.600 552.450 241.050 ;
        RECT 553.950 239.850 556.050 241.950 ;
        RECT 557.400 240.150 558.600 248.400 ;
        RECT 566.400 240.150 567.600 248.400 ;
        RECT 574.650 245.400 576.450 251.250 ;
        RECT 575.250 243.300 576.450 245.400 ;
        RECT 577.650 246.300 579.450 251.250 ;
        RECT 580.650 247.200 582.450 251.250 ;
        RECT 583.650 246.300 585.450 251.250 ;
        RECT 587.550 248.400 589.350 251.250 ;
        RECT 590.550 248.400 592.350 251.250 ;
        RECT 593.550 248.400 595.350 251.250 ;
        RECT 599.550 248.400 601.350 251.250 ;
        RECT 602.550 248.400 604.350 251.250 ;
        RECT 605.550 248.400 607.350 251.250 ;
        RECT 611.550 248.400 613.350 251.250 ;
        RECT 614.550 248.400 616.350 251.250 ;
        RECT 577.650 244.950 585.450 246.300 ;
        RECT 575.250 242.250 579.000 243.300 ;
        RECT 554.100 238.050 555.900 239.850 ;
        RECT 556.950 238.050 559.050 240.150 ;
        RECT 565.950 238.050 568.050 240.150 ;
        RECT 568.950 239.850 571.050 241.950 ;
        RECT 569.100 238.050 570.900 239.850 ;
        RECT 577.950 238.950 579.150 242.250 ;
        RECT 591.000 241.950 592.050 248.400 ;
        RECT 603.000 241.950 604.050 248.400 ;
        RECT 581.100 240.150 582.900 241.950 ;
        RECT 543.150 230.400 544.050 231.300 ;
        RECT 540.450 230.100 542.250 230.400 ;
        RECT 527.550 228.600 528.750 229.500 ;
        RECT 535.950 229.200 542.250 230.100 ;
        RECT 540.450 228.600 542.250 229.200 ;
        RECT 543.150 228.600 545.850 230.400 ;
        RECT 523.950 226.500 528.750 228.600 ;
        RECT 531.150 226.500 538.050 228.300 ;
        RECT 527.550 225.600 528.750 226.500 ;
        RECT 522.150 219.750 523.950 225.600 ;
        RECT 527.250 219.750 529.050 225.600 ;
        RECT 532.050 219.750 533.850 225.600 ;
        RECT 535.050 219.750 536.850 226.500 ;
        RECT 543.150 225.600 547.050 227.700 ;
        RECT 538.950 219.750 540.750 225.600 ;
        RECT 543.150 219.750 544.950 225.600 ;
        RECT 547.650 219.750 549.450 222.600 ;
        RECT 550.650 219.750 552.450 231.600 ;
        RECT 557.400 225.600 558.600 238.050 ;
        RECT 566.400 225.600 567.600 238.050 ;
        RECT 577.950 236.850 580.050 238.950 ;
        RECT 580.950 238.050 583.050 240.150 ;
        RECT 589.950 239.850 592.050 241.950 ;
        RECT 601.950 239.850 604.050 241.950 ;
        RECT 610.950 239.850 613.050 241.950 ;
        RECT 614.400 240.150 615.600 248.400 ;
        RECT 621.000 245.400 622.800 251.250 ;
        RECT 625.200 247.050 627.000 251.250 ;
        RECT 628.500 248.400 630.300 251.250 ;
        RECT 635.550 248.400 637.350 251.250 ;
        RECT 638.550 248.400 640.350 251.250 ;
        RECT 641.550 248.400 643.350 251.250 ;
        RECT 625.200 245.400 630.900 247.050 ;
        RECT 620.100 240.150 621.900 241.950 ;
        RECT 583.950 236.850 586.050 238.950 ;
        RECT 586.950 236.850 589.050 238.950 ;
        RECT 574.950 233.850 577.050 235.950 ;
        RECT 575.250 232.050 577.050 233.850 ;
        RECT 578.850 231.600 580.050 236.850 ;
        RECT 584.100 235.050 585.900 236.850 ;
        RECT 587.100 235.050 588.900 236.850 ;
        RECT 591.000 232.650 592.050 239.850 ;
        RECT 592.950 236.850 595.050 238.950 ;
        RECT 598.950 236.850 601.050 238.950 ;
        RECT 593.100 235.050 594.900 236.850 ;
        RECT 599.100 235.050 600.900 236.850 ;
        RECT 603.000 232.650 604.050 239.850 ;
        RECT 604.950 236.850 607.050 238.950 ;
        RECT 611.100 238.050 612.900 239.850 ;
        RECT 613.950 238.050 616.050 240.150 ;
        RECT 619.950 238.050 622.050 240.150 ;
        RECT 622.950 239.850 625.050 241.950 ;
        RECT 626.100 240.150 627.900 241.950 ;
        RECT 623.100 238.050 624.900 239.850 ;
        RECT 625.950 238.050 628.050 240.150 ;
        RECT 629.700 238.950 630.900 245.400 ;
        RECT 631.950 241.950 634.050 244.050 ;
        RECT 639.000 241.950 640.050 248.400 ;
        RECT 648.000 245.400 649.800 251.250 ;
        RECT 652.200 247.050 654.000 251.250 ;
        RECT 655.500 248.400 657.300 251.250 ;
        RECT 662.550 248.400 664.350 251.250 ;
        RECT 665.550 248.400 667.350 251.250 ;
        RECT 671.550 248.400 673.350 251.250 ;
        RECT 674.550 248.400 676.350 251.250 ;
        RECT 682.650 248.400 684.450 251.250 ;
        RECT 685.650 248.400 687.450 251.250 ;
        RECT 652.200 245.400 657.900 247.050 ;
        RECT 605.100 235.050 606.900 236.850 ;
        RECT 591.000 231.600 593.550 232.650 ;
        RECT 603.000 231.600 605.550 232.650 ;
        RECT 554.550 219.750 556.350 225.600 ;
        RECT 557.550 219.750 559.350 225.600 ;
        RECT 565.650 219.750 567.450 225.600 ;
        RECT 568.650 219.750 570.450 225.600 ;
        RECT 575.400 219.750 577.200 225.600 ;
        RECT 578.700 219.750 580.500 231.600 ;
        RECT 582.900 219.750 584.700 231.600 ;
        RECT 587.550 219.750 589.350 231.600 ;
        RECT 591.750 219.750 593.550 231.600 ;
        RECT 599.550 219.750 601.350 231.600 ;
        RECT 603.750 219.750 605.550 231.600 ;
        RECT 614.400 225.600 615.600 238.050 ;
        RECT 628.950 236.850 631.050 238.950 ;
        RECT 629.700 231.600 630.900 236.850 ;
        RECT 632.550 235.050 633.450 241.950 ;
        RECT 637.950 239.850 640.050 241.950 ;
        RECT 647.100 240.150 648.900 241.950 ;
        RECT 634.950 236.850 637.050 238.950 ;
        RECT 635.100 235.050 636.900 236.850 ;
        RECT 631.950 232.950 634.050 235.050 ;
        RECT 639.000 232.650 640.050 239.850 ;
        RECT 640.950 236.850 643.050 238.950 ;
        RECT 646.950 238.050 649.050 240.150 ;
        RECT 649.950 239.850 652.050 241.950 ;
        RECT 653.100 240.150 654.900 241.950 ;
        RECT 650.100 238.050 651.900 239.850 ;
        RECT 652.950 238.050 655.050 240.150 ;
        RECT 656.700 238.950 657.900 245.400 ;
        RECT 661.950 239.850 664.050 241.950 ;
        RECT 665.400 240.150 666.600 248.400 ;
        RECT 655.950 236.850 658.050 238.950 ;
        RECT 662.100 238.050 663.900 239.850 ;
        RECT 664.950 238.050 667.050 240.150 ;
        RECT 670.950 239.850 673.050 241.950 ;
        RECT 674.400 240.150 675.600 248.400 ;
        RECT 683.400 240.150 684.600 248.400 ;
        RECT 689.550 246.300 691.350 251.250 ;
        RECT 692.550 247.200 694.350 251.250 ;
        RECT 695.550 246.300 697.350 251.250 ;
        RECT 689.550 244.950 697.350 246.300 ;
        RECT 698.550 245.400 700.350 251.250 ;
        RECT 704.850 245.400 706.650 251.250 ;
        RECT 698.550 243.300 699.750 245.400 ;
        RECT 709.350 244.200 711.150 251.250 ;
        RECT 696.000 242.250 699.750 243.300 ;
        RECT 671.100 238.050 672.900 239.850 ;
        RECT 673.950 238.050 676.050 240.150 ;
        RECT 682.950 238.050 685.050 240.150 ;
        RECT 685.950 239.850 688.050 241.950 ;
        RECT 692.100 240.150 693.900 241.950 ;
        RECT 686.100 238.050 687.900 239.850 ;
        RECT 641.100 235.050 642.900 236.850 ;
        RECT 639.000 231.600 641.550 232.650 ;
        RECT 656.700 231.600 657.900 236.850 ;
        RECT 620.550 230.700 628.350 231.600 ;
        RECT 611.550 219.750 613.350 225.600 ;
        RECT 614.550 219.750 616.350 225.600 ;
        RECT 620.550 219.750 622.350 230.700 ;
        RECT 623.550 219.750 625.350 229.800 ;
        RECT 626.550 219.750 628.350 230.700 ;
        RECT 629.550 219.750 631.350 231.600 ;
        RECT 635.550 219.750 637.350 231.600 ;
        RECT 639.750 219.750 641.550 231.600 ;
        RECT 647.550 230.700 655.350 231.600 ;
        RECT 647.550 219.750 649.350 230.700 ;
        RECT 650.550 219.750 652.350 229.800 ;
        RECT 653.550 219.750 655.350 230.700 ;
        RECT 656.550 219.750 658.350 231.600 ;
        RECT 665.400 225.600 666.600 238.050 ;
        RECT 674.400 225.600 675.600 238.050 ;
        RECT 683.400 225.600 684.600 238.050 ;
        RECT 688.950 236.850 691.050 238.950 ;
        RECT 691.950 238.050 694.050 240.150 ;
        RECT 695.850 238.950 697.050 242.250 ;
        RECT 700.950 241.950 703.050 244.050 ;
        RECT 707.550 243.300 711.150 244.200 ;
        RECT 694.950 236.850 697.050 238.950 ;
        RECT 689.100 235.050 690.900 236.850 ;
        RECT 694.950 231.600 696.150 236.850 ;
        RECT 697.950 233.850 700.050 235.950 ;
        RECT 697.950 232.050 699.750 233.850 ;
        RECT 662.550 219.750 664.350 225.600 ;
        RECT 665.550 219.750 667.350 225.600 ;
        RECT 671.550 219.750 673.350 225.600 ;
        RECT 674.550 219.750 676.350 225.600 ;
        RECT 682.650 219.750 684.450 225.600 ;
        RECT 685.650 219.750 687.450 225.600 ;
        RECT 690.300 219.750 692.100 231.600 ;
        RECT 694.500 219.750 696.300 231.600 ;
        RECT 697.950 228.450 700.050 229.050 ;
        RECT 701.550 228.450 702.450 241.950 ;
        RECT 704.100 237.150 705.900 238.950 ;
        RECT 703.950 235.050 706.050 237.150 ;
        RECT 707.550 235.950 708.750 243.300 ;
        RECT 710.100 237.150 711.900 238.950 ;
        RECT 706.950 233.850 709.050 235.950 ;
        RECT 709.950 235.050 712.050 237.150 ;
        RECT 697.950 227.550 702.450 228.450 ;
        RECT 697.950 226.950 700.050 227.550 ;
        RECT 707.550 225.600 708.750 233.850 ;
        RECT 697.800 219.750 699.600 225.600 ;
        RECT 704.550 219.750 706.350 225.600 ;
        RECT 707.550 219.750 709.350 225.600 ;
        RECT 710.550 219.750 712.350 225.600 ;
        RECT 4.650 203.400 6.450 215.250 ;
        RECT 7.650 204.300 9.450 215.250 ;
        RECT 10.650 205.200 12.450 215.250 ;
        RECT 13.650 204.300 15.450 215.250 ;
        RECT 17.550 209.400 19.350 215.250 ;
        RECT 20.550 209.400 22.350 215.250 ;
        RECT 23.550 210.000 25.350 215.250 ;
        RECT 20.700 209.100 22.350 209.400 ;
        RECT 26.550 209.400 28.350 215.250 ;
        RECT 32.550 209.400 34.350 215.250 ;
        RECT 35.550 209.400 37.350 215.250 ;
        RECT 38.550 210.000 40.350 215.250 ;
        RECT 26.550 209.100 27.750 209.400 ;
        RECT 20.700 208.200 27.750 209.100 ;
        RECT 35.700 209.100 37.350 209.400 ;
        RECT 41.550 209.400 43.350 215.250 ;
        RECT 49.650 209.400 51.450 215.250 ;
        RECT 52.650 209.400 54.450 215.250 ;
        RECT 55.650 209.400 57.450 215.250 ;
        RECT 41.550 209.100 42.750 209.400 ;
        RECT 35.700 208.200 42.750 209.100 ;
        RECT 7.650 203.400 15.450 204.300 ;
        RECT 20.100 204.150 21.900 205.950 ;
        RECT 5.100 198.150 6.300 203.400 ;
        RECT 17.100 201.150 18.900 202.950 ;
        RECT 19.950 202.050 22.050 204.150 ;
        RECT 23.250 201.150 25.050 202.950 ;
        RECT 16.950 199.050 19.050 201.150 ;
        RECT 22.950 199.050 25.050 201.150 ;
        RECT 26.700 199.950 27.750 208.200 ;
        RECT 28.950 202.950 31.050 205.050 ;
        RECT 35.100 204.150 36.900 205.950 ;
        RECT 4.950 196.050 7.050 198.150 ;
        RECT 25.950 197.850 28.050 199.950 ;
        RECT 5.100 189.600 6.300 196.050 ;
        RECT 7.950 194.850 10.050 196.950 ;
        RECT 11.100 195.150 12.900 196.950 ;
        RECT 8.100 193.050 9.900 194.850 ;
        RECT 10.950 193.050 13.050 195.150 ;
        RECT 13.950 194.850 16.050 196.950 ;
        RECT 14.100 193.050 15.900 194.850 ;
        RECT 26.400 193.650 27.600 197.850 ;
        RECT 29.550 195.450 30.450 202.950 ;
        RECT 32.100 201.150 33.900 202.950 ;
        RECT 34.950 202.050 37.050 204.150 ;
        RECT 38.250 201.150 40.050 202.950 ;
        RECT 31.950 199.050 34.050 201.150 ;
        RECT 37.950 199.050 40.050 201.150 ;
        RECT 41.700 199.950 42.750 208.200 ;
        RECT 43.950 202.950 46.050 205.050 ;
        RECT 40.950 197.850 43.050 199.950 ;
        RECT 31.950 195.450 34.050 196.050 ;
        RECT 29.550 194.550 34.050 195.450 ;
        RECT 31.950 193.950 34.050 194.550 ;
        RECT 41.400 193.650 42.600 197.850 ;
        RECT 5.100 187.950 10.800 189.600 ;
        RECT 5.700 183.750 7.500 186.600 ;
        RECT 9.000 183.750 10.800 187.950 ;
        RECT 13.200 183.750 15.000 189.600 ;
        RECT 17.700 183.750 19.500 192.600 ;
        RECT 23.100 192.000 27.600 193.650 ;
        RECT 23.100 183.750 24.900 192.000 ;
        RECT 32.700 183.750 34.500 192.600 ;
        RECT 38.100 192.000 42.600 193.650 ;
        RECT 44.550 193.050 45.450 202.950 ;
        RECT 53.250 201.150 54.450 209.400 ;
        RECT 60.300 203.400 62.100 215.250 ;
        RECT 64.500 203.400 66.300 215.250 ;
        RECT 67.800 209.400 69.600 215.250 ;
        RECT 49.950 197.850 52.050 199.950 ;
        RECT 52.950 199.050 55.050 201.150 ;
        RECT 50.100 196.050 51.900 197.850 ;
        RECT 38.100 183.750 39.900 192.000 ;
        RECT 43.950 190.950 46.050 193.050 ;
        RECT 53.250 191.700 54.450 199.050 ;
        RECT 55.950 197.850 58.050 199.950 ;
        RECT 59.100 198.150 60.900 199.950 ;
        RECT 64.950 198.150 66.150 203.400 ;
        RECT 70.950 202.950 73.050 205.050 ;
        RECT 74.550 204.300 76.350 215.250 ;
        RECT 77.550 205.200 79.350 215.250 ;
        RECT 80.550 204.300 82.350 215.250 ;
        RECT 74.550 203.400 82.350 204.300 ;
        RECT 83.550 203.400 85.350 215.250 ;
        RECT 90.300 203.400 92.100 215.250 ;
        RECT 94.500 203.400 96.300 215.250 ;
        RECT 97.800 209.400 99.600 215.250 ;
        RECT 105.300 203.400 107.100 215.250 ;
        RECT 109.500 203.400 111.300 215.250 ;
        RECT 112.800 209.400 114.600 215.250 ;
        RECT 119.550 209.400 121.350 215.250 ;
        RECT 122.550 209.400 124.350 215.250 ;
        RECT 67.950 201.150 69.750 202.950 ;
        RECT 67.950 199.050 70.050 201.150 ;
        RECT 56.100 196.050 57.900 197.850 ;
        RECT 58.950 196.050 61.050 198.150 ;
        RECT 61.950 194.850 64.050 196.950 ;
        RECT 64.950 196.050 67.050 198.150 ;
        RECT 71.550 196.050 72.450 202.950 ;
        RECT 83.700 198.150 84.900 203.400 ;
        RECT 89.100 198.150 90.900 199.950 ;
        RECT 94.950 198.150 96.150 203.400 ;
        RECT 97.950 201.150 99.750 202.950 ;
        RECT 97.950 199.050 100.050 201.150 ;
        RECT 104.100 198.150 105.900 199.950 ;
        RECT 109.950 198.150 111.150 203.400 ;
        RECT 112.950 201.150 114.750 202.950 ;
        RECT 112.950 199.050 115.050 201.150 ;
        RECT 119.100 198.150 120.900 199.950 ;
        RECT 62.100 193.050 63.900 194.850 ;
        RECT 65.850 192.750 67.050 196.050 ;
        RECT 70.950 193.950 73.050 196.050 ;
        RECT 73.950 194.850 76.050 196.950 ;
        RECT 77.100 195.150 78.900 196.950 ;
        RECT 74.100 193.050 75.900 194.850 ;
        RECT 76.950 193.050 79.050 195.150 ;
        RECT 79.950 194.850 82.050 196.950 ;
        RECT 82.950 196.050 85.050 198.150 ;
        RECT 88.950 196.050 91.050 198.150 ;
        RECT 80.100 193.050 81.900 194.850 ;
        RECT 66.000 191.700 69.750 192.750 ;
        RECT 50.850 190.800 54.450 191.700 ;
        RECT 50.850 183.750 52.650 190.800 ;
        RECT 55.350 183.750 57.150 189.600 ;
        RECT 59.550 188.700 67.350 190.050 ;
        RECT 59.550 183.750 61.350 188.700 ;
        RECT 62.550 183.750 64.350 187.800 ;
        RECT 65.550 183.750 67.350 188.700 ;
        RECT 68.550 189.600 69.750 191.700 ;
        RECT 83.700 189.600 84.900 196.050 ;
        RECT 91.950 194.850 94.050 196.950 ;
        RECT 94.950 196.050 97.050 198.150 ;
        RECT 103.950 196.050 106.050 198.150 ;
        RECT 92.100 193.050 93.900 194.850 ;
        RECT 95.850 192.750 97.050 196.050 ;
        RECT 106.950 194.850 109.050 196.950 ;
        RECT 109.950 196.050 112.050 198.150 ;
        RECT 118.950 196.050 121.050 198.150 ;
        RECT 107.100 193.050 108.900 194.850 ;
        RECT 110.850 192.750 112.050 196.050 ;
        RECT 96.000 191.700 99.750 192.750 ;
        RECT 111.000 191.700 114.750 192.750 ;
        RECT 122.700 192.300 123.900 209.400 ;
        RECT 126.150 203.400 127.950 215.250 ;
        RECT 129.150 203.400 130.950 215.250 ;
        RECT 136.650 209.400 138.450 215.250 ;
        RECT 139.650 209.400 141.450 215.250 ;
        RECT 142.650 209.400 144.450 215.250 ;
        RECT 146.550 209.400 148.350 215.250 ;
        RECT 149.550 209.400 151.350 215.250 ;
        RECT 152.550 209.400 154.350 215.250 ;
        RECT 160.650 209.400 162.450 215.250 ;
        RECT 163.650 210.000 165.450 215.250 ;
        RECT 124.950 197.850 127.050 199.950 ;
        RECT 129.150 198.150 130.350 203.400 ;
        RECT 140.250 201.150 141.450 209.400 ;
        RECT 149.550 201.150 150.750 209.400 ;
        RECT 161.250 209.100 162.450 209.400 ;
        RECT 166.650 209.400 168.450 215.250 ;
        RECT 169.650 209.400 171.450 215.250 ;
        RECT 175.650 209.400 177.450 215.250 ;
        RECT 178.650 209.400 180.450 215.250 ;
        RECT 166.650 209.100 168.300 209.400 ;
        RECT 161.250 208.200 168.300 209.100 ;
        RECT 125.100 196.050 126.900 197.850 ;
        RECT 127.950 196.050 130.350 198.150 ;
        RECT 136.950 197.850 139.050 199.950 ;
        RECT 139.950 199.050 142.050 201.150 ;
        RECT 137.100 196.050 138.900 197.850 ;
        RECT 68.550 183.750 70.350 189.600 ;
        RECT 75.000 183.750 76.800 189.600 ;
        RECT 79.200 187.950 84.900 189.600 ;
        RECT 89.550 188.700 97.350 190.050 ;
        RECT 79.200 183.750 81.000 187.950 ;
        RECT 82.500 183.750 84.300 186.600 ;
        RECT 89.550 183.750 91.350 188.700 ;
        RECT 92.550 183.750 94.350 187.800 ;
        RECT 95.550 183.750 97.350 188.700 ;
        RECT 98.550 189.600 99.750 191.700 ;
        RECT 98.550 183.750 100.350 189.600 ;
        RECT 104.550 188.700 112.350 190.050 ;
        RECT 104.550 183.750 106.350 188.700 ;
        RECT 107.550 183.750 109.350 187.800 ;
        RECT 110.550 183.750 112.350 188.700 ;
        RECT 113.550 189.600 114.750 191.700 ;
        RECT 119.550 191.100 127.050 192.300 ;
        RECT 113.550 183.750 115.350 189.600 ;
        RECT 119.550 183.750 121.350 191.100 ;
        RECT 125.250 190.500 127.050 191.100 ;
        RECT 129.150 189.600 130.350 196.050 ;
        RECT 140.250 191.700 141.450 199.050 ;
        RECT 142.950 197.850 145.050 199.950 ;
        RECT 145.950 197.850 148.050 199.950 ;
        RECT 148.950 199.050 151.050 201.150 ;
        RECT 161.250 199.950 162.300 208.200 ;
        RECT 167.100 204.150 168.900 205.950 ;
        RECT 163.950 201.150 165.750 202.950 ;
        RECT 166.950 202.050 169.050 204.150 ;
        RECT 170.100 201.150 171.900 202.950 ;
        RECT 143.100 196.050 144.900 197.850 ;
        RECT 146.100 196.050 147.900 197.850 ;
        RECT 124.050 183.750 125.850 189.600 ;
        RECT 127.050 188.100 130.350 189.600 ;
        RECT 137.850 190.800 141.450 191.700 ;
        RECT 149.550 191.700 150.750 199.050 ;
        RECT 151.950 197.850 154.050 199.950 ;
        RECT 160.950 197.850 163.050 199.950 ;
        RECT 163.950 199.050 166.050 201.150 ;
        RECT 169.950 199.050 172.050 201.150 ;
        RECT 152.100 196.050 153.900 197.850 ;
        RECT 161.400 193.650 162.600 197.850 ;
        RECT 176.400 196.950 177.600 209.400 ;
        RECT 184.050 203.400 185.850 215.250 ;
        RECT 187.050 203.400 188.850 215.250 ;
        RECT 190.650 209.400 192.450 215.250 ;
        RECT 193.650 209.400 195.450 215.250 ;
        RECT 184.650 198.150 185.850 203.400 ;
        RECT 175.950 194.850 178.050 196.950 ;
        RECT 179.100 195.150 180.900 196.950 ;
        RECT 184.650 196.050 187.050 198.150 ;
        RECT 187.950 197.850 190.050 199.950 ;
        RECT 188.100 196.050 189.900 197.850 ;
        RECT 161.400 192.000 165.900 193.650 ;
        RECT 149.550 190.800 153.150 191.700 ;
        RECT 127.050 183.750 128.850 188.100 ;
        RECT 137.850 183.750 139.650 190.800 ;
        RECT 142.350 183.750 144.150 189.600 ;
        RECT 146.850 183.750 148.650 189.600 ;
        RECT 151.350 183.750 153.150 190.800 ;
        RECT 164.100 183.750 165.900 192.000 ;
        RECT 169.500 183.750 171.300 192.600 ;
        RECT 176.400 186.600 177.600 194.850 ;
        RECT 178.950 193.050 181.050 195.150 ;
        RECT 184.650 189.600 185.850 196.050 ;
        RECT 191.100 192.300 192.300 209.400 ;
        RECT 198.300 203.400 200.100 215.250 ;
        RECT 202.500 203.400 204.300 215.250 ;
        RECT 205.800 209.400 207.600 215.250 ;
        RECT 215.400 209.400 217.200 215.250 ;
        RECT 218.700 203.400 220.500 215.250 ;
        RECT 222.900 203.400 224.700 215.250 ;
        RECT 227.550 209.400 229.350 215.250 ;
        RECT 230.550 209.400 232.350 215.250 ;
        RECT 233.550 209.400 235.350 215.250 ;
        RECT 194.100 198.150 195.900 199.950 ;
        RECT 197.100 198.150 198.900 199.950 ;
        RECT 202.950 198.150 204.150 203.400 ;
        RECT 205.950 201.150 207.750 202.950 ;
        RECT 215.250 201.150 217.050 202.950 ;
        RECT 205.950 199.050 208.050 201.150 ;
        RECT 214.950 199.050 217.050 201.150 ;
        RECT 218.850 198.150 220.050 203.400 ;
        RECT 230.550 201.150 231.750 209.400 ;
        RECT 240.300 203.400 242.100 215.250 ;
        RECT 244.500 203.400 246.300 215.250 ;
        RECT 247.800 209.400 249.600 215.250 ;
        RECT 254.550 209.400 256.350 215.250 ;
        RECT 257.550 209.400 259.350 215.250 ;
        RECT 260.550 209.400 262.350 215.250 ;
        RECT 224.100 198.150 225.900 199.950 ;
        RECT 193.950 196.050 196.050 198.150 ;
        RECT 196.950 196.050 199.050 198.150 ;
        RECT 199.950 194.850 202.050 196.950 ;
        RECT 202.950 196.050 205.050 198.150 ;
        RECT 200.100 193.050 201.900 194.850 ;
        RECT 203.850 192.750 205.050 196.050 ;
        RECT 217.950 196.050 220.050 198.150 ;
        RECT 217.950 192.750 219.150 196.050 ;
        RECT 220.950 194.850 223.050 196.950 ;
        RECT 223.950 196.050 226.050 198.150 ;
        RECT 226.950 197.850 229.050 199.950 ;
        RECT 229.950 199.050 232.050 201.150 ;
        RECT 227.100 196.050 228.900 197.850 ;
        RECT 221.100 193.050 222.900 194.850 ;
        RECT 187.950 191.100 195.450 192.300 ;
        RECT 204.000 191.700 207.750 192.750 ;
        RECT 187.950 190.500 189.750 191.100 ;
        RECT 184.650 188.100 187.950 189.600 ;
        RECT 175.650 183.750 177.450 186.600 ;
        RECT 178.650 183.750 180.450 186.600 ;
        RECT 186.150 183.750 187.950 188.100 ;
        RECT 189.150 183.750 190.950 189.600 ;
        RECT 193.650 183.750 195.450 191.100 ;
        RECT 197.550 188.700 205.350 190.050 ;
        RECT 197.550 183.750 199.350 188.700 ;
        RECT 200.550 183.750 202.350 187.800 ;
        RECT 203.550 183.750 205.350 188.700 ;
        RECT 206.550 189.600 207.750 191.700 ;
        RECT 215.250 191.700 219.000 192.750 ;
        RECT 230.550 191.700 231.750 199.050 ;
        RECT 232.950 197.850 235.050 199.950 ;
        RECT 239.100 198.150 240.900 199.950 ;
        RECT 244.950 198.150 246.150 203.400 ;
        RECT 247.950 201.150 249.750 202.950 ;
        RECT 257.550 201.150 258.750 209.400 ;
        RECT 266.550 204.300 268.350 215.250 ;
        RECT 269.550 205.200 271.350 215.250 ;
        RECT 272.550 204.300 274.350 215.250 ;
        RECT 266.550 203.400 274.350 204.300 ;
        RECT 275.550 203.400 277.350 215.250 ;
        RECT 281.550 209.400 283.350 215.250 ;
        RECT 284.550 209.400 286.350 215.250 ;
        RECT 287.550 210.000 289.350 215.250 ;
        RECT 284.700 209.100 286.350 209.400 ;
        RECT 290.550 209.400 292.350 215.250 ;
        RECT 290.550 209.100 291.750 209.400 ;
        RECT 284.700 208.200 291.750 209.100 ;
        RECT 284.100 204.150 285.900 205.950 ;
        RECT 247.950 199.050 250.050 201.150 ;
        RECT 233.100 196.050 234.900 197.850 ;
        RECT 238.950 196.050 241.050 198.150 ;
        RECT 241.950 194.850 244.050 196.950 ;
        RECT 244.950 196.050 247.050 198.150 ;
        RECT 253.950 197.850 256.050 199.950 ;
        RECT 256.950 199.050 259.050 201.150 ;
        RECT 254.100 196.050 255.900 197.850 ;
        RECT 242.100 193.050 243.900 194.850 ;
        RECT 245.850 192.750 247.050 196.050 ;
        RECT 246.000 191.700 249.750 192.750 ;
        RECT 215.250 189.600 216.450 191.700 ;
        RECT 230.550 190.800 234.150 191.700 ;
        RECT 206.550 183.750 208.350 189.600 ;
        RECT 214.650 183.750 216.450 189.600 ;
        RECT 217.650 188.700 225.450 190.050 ;
        RECT 217.650 183.750 219.450 188.700 ;
        RECT 220.650 183.750 222.450 187.800 ;
        RECT 223.650 183.750 225.450 188.700 ;
        RECT 227.850 183.750 229.650 189.600 ;
        RECT 232.350 183.750 234.150 190.800 ;
        RECT 239.550 188.700 247.350 190.050 ;
        RECT 239.550 183.750 241.350 188.700 ;
        RECT 242.550 183.750 244.350 187.800 ;
        RECT 245.550 183.750 247.350 188.700 ;
        RECT 248.550 189.600 249.750 191.700 ;
        RECT 257.550 191.700 258.750 199.050 ;
        RECT 259.950 197.850 262.050 199.950 ;
        RECT 275.700 198.150 276.900 203.400 ;
        RECT 281.100 201.150 282.900 202.950 ;
        RECT 283.950 202.050 286.050 204.150 ;
        RECT 287.250 201.150 289.050 202.950 ;
        RECT 280.950 199.050 283.050 201.150 ;
        RECT 286.950 199.050 289.050 201.150 ;
        RECT 290.700 199.950 291.750 208.200 ;
        RECT 297.300 203.400 299.100 215.250 ;
        RECT 301.500 203.400 303.300 215.250 ;
        RECT 304.800 209.400 306.600 215.250 ;
        RECT 311.550 209.400 313.350 215.250 ;
        RECT 314.550 209.400 316.350 215.250 ;
        RECT 320.550 209.400 322.350 215.250 ;
        RECT 323.550 209.400 325.350 215.250 ;
        RECT 326.550 210.000 328.350 215.250 ;
        RECT 260.100 196.050 261.900 197.850 ;
        RECT 265.950 194.850 268.050 196.950 ;
        RECT 269.100 195.150 270.900 196.950 ;
        RECT 266.100 193.050 267.900 194.850 ;
        RECT 268.950 193.050 271.050 195.150 ;
        RECT 271.950 194.850 274.050 196.950 ;
        RECT 274.950 196.050 277.050 198.150 ;
        RECT 289.950 197.850 292.050 199.950 ;
        RECT 296.100 198.150 297.900 199.950 ;
        RECT 301.950 198.150 303.150 203.400 ;
        RECT 304.950 201.150 306.750 202.950 ;
        RECT 304.950 199.050 307.050 201.150 ;
        RECT 272.100 193.050 273.900 194.850 ;
        RECT 257.550 190.800 261.150 191.700 ;
        RECT 248.550 183.750 250.350 189.600 ;
        RECT 254.850 183.750 256.650 189.600 ;
        RECT 259.350 183.750 261.150 190.800 ;
        RECT 275.700 189.600 276.900 196.050 ;
        RECT 290.400 193.650 291.600 197.850 ;
        RECT 295.950 196.050 298.050 198.150 ;
        RECT 298.950 194.850 301.050 196.950 ;
        RECT 301.950 196.050 304.050 198.150 ;
        RECT 314.400 196.950 315.600 209.400 ;
        RECT 323.700 209.100 325.350 209.400 ;
        RECT 329.550 209.400 331.350 215.250 ;
        RECT 335.550 209.400 337.350 215.250 ;
        RECT 338.550 209.400 340.350 215.250 ;
        RECT 341.550 209.400 343.350 215.250 ;
        RECT 329.550 209.100 330.750 209.400 ;
        RECT 323.700 208.200 330.750 209.100 ;
        RECT 323.100 204.150 324.900 205.950 ;
        RECT 320.100 201.150 321.900 202.950 ;
        RECT 322.950 202.050 325.050 204.150 ;
        RECT 326.250 201.150 328.050 202.950 ;
        RECT 319.950 199.050 322.050 201.150 ;
        RECT 325.950 199.050 328.050 201.150 ;
        RECT 329.700 199.950 330.750 208.200 ;
        RECT 338.550 201.150 339.750 209.400 ;
        RECT 347.550 203.400 349.350 215.250 ;
        RECT 352.050 203.550 353.850 215.250 ;
        RECT 355.050 204.900 356.850 215.250 ;
        RECT 364.650 209.400 366.450 215.250 ;
        RECT 367.650 209.400 369.450 215.250 ;
        RECT 370.650 209.400 372.450 215.250 ;
        RECT 374.550 209.400 376.350 215.250 ;
        RECT 377.550 209.400 379.350 215.250 ;
        RECT 355.050 203.550 357.450 204.900 ;
        RECT 347.550 202.200 348.750 203.400 ;
        RECT 352.950 202.200 354.750 202.650 ;
        RECT 328.950 197.850 331.050 199.950 ;
        RECT 334.950 197.850 337.050 199.950 ;
        RECT 337.950 199.050 340.050 201.150 ;
        RECT 347.550 201.000 354.750 202.200 ;
        RECT 352.950 200.850 354.750 201.000 ;
        RECT 267.000 183.750 268.800 189.600 ;
        RECT 271.200 187.950 276.900 189.600 ;
        RECT 271.200 183.750 273.000 187.950 ;
        RECT 274.500 183.750 276.300 186.600 ;
        RECT 281.700 183.750 283.500 192.600 ;
        RECT 287.100 192.000 291.600 193.650 ;
        RECT 299.100 193.050 300.900 194.850 ;
        RECT 302.850 192.750 304.050 196.050 ;
        RECT 311.100 195.150 312.900 196.950 ;
        RECT 310.950 193.050 313.050 195.150 ;
        RECT 313.950 194.850 316.050 196.950 ;
        RECT 287.100 183.750 288.900 192.000 ;
        RECT 303.000 191.700 306.750 192.750 ;
        RECT 296.550 188.700 304.350 190.050 ;
        RECT 296.550 183.750 298.350 188.700 ;
        RECT 299.550 183.750 301.350 187.800 ;
        RECT 302.550 183.750 304.350 188.700 ;
        RECT 305.550 189.600 306.750 191.700 ;
        RECT 305.550 183.750 307.350 189.600 ;
        RECT 314.400 186.600 315.600 194.850 ;
        RECT 329.400 193.650 330.600 197.850 ;
        RECT 335.100 196.050 336.900 197.850 ;
        RECT 311.550 183.750 313.350 186.600 ;
        RECT 314.550 183.750 316.350 186.600 ;
        RECT 320.700 183.750 322.500 192.600 ;
        RECT 326.100 192.000 330.600 193.650 ;
        RECT 326.100 183.750 327.900 192.000 ;
        RECT 338.550 191.700 339.750 199.050 ;
        RECT 340.950 197.850 343.050 199.950 ;
        RECT 350.100 198.150 351.900 199.950 ;
        RECT 341.100 196.050 342.900 197.850 ;
        RECT 347.100 195.150 348.900 196.950 ;
        RECT 349.950 196.050 352.050 198.150 ;
        RECT 346.950 193.050 349.050 195.150 ;
        RECT 353.700 192.600 354.600 200.850 ;
        RECT 356.100 196.950 357.450 203.550 ;
        RECT 368.250 201.150 369.450 209.400 ;
        RECT 364.950 197.850 367.050 199.950 ;
        RECT 367.950 199.050 370.050 201.150 ;
        RECT 355.950 194.850 358.050 196.950 ;
        RECT 365.100 196.050 366.900 197.850 ;
        RECT 352.950 191.700 354.750 192.600 ;
        RECT 338.550 190.800 342.150 191.700 ;
        RECT 335.850 183.750 337.650 189.600 ;
        RECT 340.350 183.750 342.150 190.800 ;
        RECT 351.450 190.800 354.750 191.700 ;
        RECT 351.450 186.600 352.350 190.800 ;
        RECT 357.000 189.600 358.050 194.850 ;
        RECT 368.250 191.700 369.450 199.050 ;
        RECT 370.950 197.850 373.050 199.950 ;
        RECT 371.100 196.050 372.900 197.850 ;
        RECT 377.400 196.950 378.600 209.400 ;
        RECT 385.350 203.400 387.150 215.250 ;
        RECT 388.350 203.400 390.150 215.250 ;
        RECT 391.650 209.400 393.450 215.250 ;
        RECT 385.650 198.150 386.850 203.400 ;
        RECT 392.250 202.500 393.450 209.400 ;
        RECT 396.300 203.400 398.100 215.250 ;
        RECT 400.500 203.400 402.300 215.250 ;
        RECT 403.800 209.400 405.600 215.250 ;
        RECT 414.150 203.400 415.950 215.250 ;
        RECT 418.650 203.400 421.950 215.250 ;
        RECT 424.650 203.400 426.450 215.250 ;
        RECT 429.150 203.400 430.950 215.250 ;
        RECT 432.150 209.400 433.950 215.250 ;
        RECT 437.250 209.400 439.050 215.250 ;
        RECT 442.050 209.400 443.850 215.250 ;
        RECT 437.550 208.500 438.750 209.400 ;
        RECT 445.050 208.500 446.850 215.250 ;
        RECT 448.950 209.400 450.750 215.250 ;
        RECT 453.150 209.400 454.950 215.250 ;
        RECT 457.650 212.400 459.450 215.250 ;
        RECT 433.950 206.400 438.750 208.500 ;
        RECT 441.150 206.700 448.050 208.500 ;
        RECT 453.150 207.300 457.050 209.400 ;
        RECT 437.550 205.500 438.750 206.400 ;
        RECT 450.450 205.800 452.250 206.400 ;
        RECT 437.550 204.300 445.050 205.500 ;
        RECT 443.250 203.700 445.050 204.300 ;
        RECT 445.950 204.900 452.250 205.800 ;
        RECT 387.750 201.600 393.450 202.500 ;
        RECT 387.750 200.700 390.000 201.600 ;
        RECT 374.100 195.150 375.900 196.950 ;
        RECT 373.950 193.050 376.050 195.150 ;
        RECT 376.950 194.850 379.050 196.950 ;
        RECT 385.650 196.050 388.050 198.150 ;
        RECT 365.850 190.800 369.450 191.700 ;
        RECT 347.550 183.750 349.350 186.600 ;
        RECT 350.550 183.750 352.350 186.600 ;
        RECT 353.550 183.750 355.350 186.600 ;
        RECT 356.550 183.750 358.350 189.600 ;
        RECT 365.850 183.750 367.650 190.800 ;
        RECT 370.350 183.750 372.150 189.600 ;
        RECT 377.400 186.600 378.600 194.850 ;
        RECT 385.650 189.600 386.850 196.050 ;
        RECT 388.950 192.300 390.000 200.700 ;
        RECT 392.100 198.150 393.900 199.950 ;
        RECT 395.100 198.150 396.900 199.950 ;
        RECT 400.950 198.150 402.150 203.400 ;
        RECT 403.950 201.150 405.750 202.950 ;
        RECT 403.950 199.050 406.050 201.150 ;
        RECT 413.250 198.150 415.050 199.950 ;
        RECT 419.250 198.150 420.450 203.400 ;
        RECT 429.150 202.800 440.250 203.400 ;
        RECT 445.950 202.800 446.850 204.900 ;
        RECT 450.450 204.600 452.250 204.900 ;
        RECT 453.150 204.600 455.850 206.400 ;
        RECT 453.150 203.700 454.050 204.600 ;
        RECT 429.150 202.200 446.850 202.800 ;
        RECT 425.100 198.150 426.900 199.950 ;
        RECT 391.950 196.050 394.050 198.150 ;
        RECT 394.950 196.050 397.050 198.150 ;
        RECT 397.950 194.850 400.050 196.950 ;
        RECT 400.950 196.050 403.050 198.150 ;
        RECT 412.950 196.050 415.050 198.150 ;
        RECT 398.100 193.050 399.900 194.850 ;
        RECT 401.850 192.750 403.050 196.050 ;
        RECT 415.950 194.850 418.050 196.950 ;
        RECT 418.950 196.050 421.050 198.150 ;
        RECT 416.700 193.050 418.500 194.850 ;
        RECT 387.750 191.400 390.000 192.300 ;
        RECT 402.000 191.700 405.750 192.750 ;
        RECT 419.400 192.150 420.600 196.050 ;
        RECT 421.950 194.850 424.050 196.950 ;
        RECT 424.950 196.050 427.050 198.150 ;
        RECT 422.100 193.050 423.900 194.850 ;
        RECT 387.750 190.500 392.850 191.400 ;
        RECT 374.550 183.750 376.350 186.600 ;
        RECT 377.550 183.750 379.350 186.600 ;
        RECT 385.350 183.750 387.150 189.600 ;
        RECT 388.350 183.750 390.150 189.600 ;
        RECT 391.650 186.600 392.850 190.500 ;
        RECT 395.550 188.700 403.350 190.050 ;
        RECT 391.650 183.750 393.450 186.600 ;
        RECT 395.550 183.750 397.350 188.700 ;
        RECT 398.550 183.750 400.350 187.800 ;
        RECT 401.550 183.750 403.350 188.700 ;
        RECT 404.550 189.600 405.750 191.700 ;
        RECT 416.250 191.100 420.600 192.150 ;
        RECT 416.250 189.600 417.150 191.100 ;
        RECT 404.550 183.750 406.350 189.600 ;
        RECT 412.650 184.500 414.450 189.600 ;
        RECT 415.650 185.400 417.450 189.600 ;
        RECT 418.650 189.000 426.450 189.900 ;
        RECT 418.650 184.500 420.450 189.000 ;
        RECT 412.650 183.750 420.450 184.500 ;
        RECT 421.650 183.750 423.450 188.100 ;
        RECT 424.650 183.750 426.450 189.000 ;
        RECT 429.150 189.600 430.050 202.200 ;
        RECT 438.450 201.900 446.850 202.200 ;
        RECT 448.050 202.800 454.050 203.700 ;
        RECT 454.950 202.800 457.050 203.700 ;
        RECT 460.650 203.400 462.450 215.250 ;
        RECT 438.450 201.600 440.250 201.900 ;
        RECT 448.050 198.150 448.950 202.800 ;
        RECT 454.950 201.600 459.150 202.800 ;
        RECT 458.250 199.800 460.050 201.600 ;
        RECT 439.950 197.100 442.050 198.150 ;
        RECT 431.100 195.150 432.900 196.950 ;
        RECT 434.100 196.050 442.050 197.100 ;
        RECT 445.950 196.050 448.950 198.150 ;
        RECT 434.100 195.300 435.900 196.050 ;
        RECT 432.000 194.400 432.900 195.150 ;
        RECT 437.100 194.400 438.900 195.000 ;
        RECT 432.000 193.200 438.900 194.400 ;
        RECT 437.850 192.000 438.900 193.200 ;
        RECT 448.050 192.000 448.950 196.050 ;
        RECT 457.950 195.750 460.050 196.050 ;
        RECT 456.150 193.950 460.050 195.750 ;
        RECT 461.250 193.950 462.450 203.400 ;
        RECT 468.450 203.400 470.250 215.250 ;
        RECT 472.650 203.400 474.450 215.250 ;
        RECT 478.650 203.400 480.450 215.250 ;
        RECT 481.650 204.300 483.450 215.250 ;
        RECT 484.650 205.200 486.450 215.250 ;
        RECT 487.650 204.300 489.450 215.250 ;
        RECT 481.650 203.400 489.450 204.300 ;
        RECT 492.150 203.400 493.950 215.250 ;
        RECT 495.150 209.400 496.950 215.250 ;
        RECT 500.250 209.400 502.050 215.250 ;
        RECT 505.050 209.400 506.850 215.250 ;
        RECT 500.550 208.500 501.750 209.400 ;
        RECT 508.050 208.500 509.850 215.250 ;
        RECT 511.950 209.400 513.750 215.250 ;
        RECT 516.150 209.400 517.950 215.250 ;
        RECT 520.650 212.400 522.450 215.250 ;
        RECT 496.950 206.400 501.750 208.500 ;
        RECT 504.150 206.700 511.050 208.500 ;
        RECT 516.150 207.300 520.050 209.400 ;
        RECT 500.550 205.500 501.750 206.400 ;
        RECT 513.450 205.800 515.250 206.400 ;
        RECT 500.550 204.300 508.050 205.500 ;
        RECT 506.250 203.700 508.050 204.300 ;
        RECT 508.950 204.900 515.250 205.800 ;
        RECT 468.450 202.350 471.000 203.400 ;
        RECT 467.100 198.150 468.900 199.950 ;
        RECT 466.950 196.050 469.050 198.150 ;
        RECT 437.850 191.100 448.950 192.000 ;
        RECT 457.950 191.850 462.450 193.950 ;
        RECT 437.850 190.200 438.900 191.100 ;
        RECT 448.050 190.800 448.950 191.100 ;
        RECT 429.150 183.750 430.950 189.600 ;
        RECT 433.950 187.500 436.050 189.600 ;
        RECT 437.550 188.400 439.350 190.200 ;
        RECT 440.850 189.450 442.650 190.200 ;
        RECT 440.850 188.400 445.800 189.450 ;
        RECT 448.050 189.000 449.850 190.800 ;
        RECT 461.250 189.600 462.450 191.850 ;
        RECT 454.950 188.700 457.050 189.600 ;
        RECT 435.000 186.600 436.050 187.500 ;
        RECT 444.750 186.600 445.800 188.400 ;
        RECT 453.300 187.500 457.050 188.700 ;
        RECT 453.300 186.600 454.350 187.500 ;
        RECT 432.150 183.750 433.950 186.600 ;
        RECT 435.000 185.700 438.750 186.600 ;
        RECT 436.950 183.750 438.750 185.700 ;
        RECT 441.450 183.750 443.250 186.600 ;
        RECT 444.750 183.750 446.550 186.600 ;
        RECT 448.650 183.750 450.450 186.600 ;
        RECT 452.850 183.750 454.650 186.600 ;
        RECT 457.350 183.750 459.150 186.600 ;
        RECT 460.650 183.750 462.450 189.600 ;
        RECT 469.950 195.150 471.000 202.350 ;
        RECT 473.100 198.150 474.900 199.950 ;
        RECT 479.100 198.150 480.300 203.400 ;
        RECT 492.150 202.800 503.250 203.400 ;
        RECT 508.950 202.800 509.850 204.900 ;
        RECT 513.450 204.600 515.250 204.900 ;
        RECT 516.150 204.600 518.850 206.400 ;
        RECT 516.150 203.700 517.050 204.600 ;
        RECT 492.150 202.200 509.850 202.800 ;
        RECT 472.950 196.050 475.050 198.150 ;
        RECT 478.950 196.050 481.050 198.150 ;
        RECT 469.950 193.050 472.050 195.150 ;
        RECT 469.950 186.600 471.000 193.050 ;
        RECT 479.100 189.600 480.300 196.050 ;
        RECT 481.950 194.850 484.050 196.950 ;
        RECT 485.100 195.150 486.900 196.950 ;
        RECT 482.100 193.050 483.900 194.850 ;
        RECT 484.950 193.050 487.050 195.150 ;
        RECT 487.950 194.850 490.050 196.950 ;
        RECT 488.100 193.050 489.900 194.850 ;
        RECT 492.150 189.600 493.050 202.200 ;
        RECT 501.450 201.900 509.850 202.200 ;
        RECT 511.050 202.800 517.050 203.700 ;
        RECT 517.950 202.800 520.050 203.700 ;
        RECT 523.650 203.400 525.450 215.250 ;
        RECT 529.650 209.400 531.450 215.250 ;
        RECT 532.650 209.400 534.450 215.250 ;
        RECT 501.450 201.600 503.250 201.900 ;
        RECT 511.050 198.150 511.950 202.800 ;
        RECT 517.950 201.600 522.150 202.800 ;
        RECT 521.250 199.800 523.050 201.600 ;
        RECT 502.950 197.100 505.050 198.150 ;
        RECT 494.100 195.150 495.900 196.950 ;
        RECT 497.100 196.050 505.050 197.100 ;
        RECT 508.950 196.050 511.950 198.150 ;
        RECT 497.100 195.300 498.900 196.050 ;
        RECT 495.000 194.400 495.900 195.150 ;
        RECT 500.100 194.400 501.900 195.000 ;
        RECT 495.000 193.200 501.900 194.400 ;
        RECT 500.850 192.000 501.900 193.200 ;
        RECT 511.050 192.000 511.950 196.050 ;
        RECT 520.950 195.750 523.050 196.050 ;
        RECT 519.150 193.950 523.050 195.750 ;
        RECT 524.250 193.950 525.450 203.400 ;
        RECT 530.400 196.950 531.600 209.400 ;
        RECT 540.450 203.400 542.250 215.250 ;
        RECT 544.650 203.400 546.450 215.250 ;
        RECT 552.450 203.400 554.250 215.250 ;
        RECT 556.650 203.400 558.450 215.250 ;
        RECT 560.550 209.400 562.350 215.250 ;
        RECT 563.550 209.400 565.350 215.250 ;
        RECT 540.450 202.350 543.000 203.400 ;
        RECT 552.450 202.350 555.000 203.400 ;
        RECT 539.100 198.150 540.900 199.950 ;
        RECT 529.950 194.850 532.050 196.950 ;
        RECT 533.100 195.150 534.900 196.950 ;
        RECT 538.950 196.050 541.050 198.150 ;
        RECT 541.950 195.150 543.000 202.350 ;
        RECT 545.100 198.150 546.900 199.950 ;
        RECT 551.100 198.150 552.900 199.950 ;
        RECT 544.950 196.050 547.050 198.150 ;
        RECT 550.950 196.050 553.050 198.150 ;
        RECT 553.950 195.150 555.000 202.350 ;
        RECT 557.100 198.150 558.900 199.950 ;
        RECT 556.950 196.050 559.050 198.150 ;
        RECT 563.400 196.950 564.600 209.400 ;
        RECT 569.550 203.400 571.350 215.250 ;
        RECT 572.550 212.400 574.350 215.250 ;
        RECT 577.050 209.400 578.850 215.250 ;
        RECT 581.250 209.400 583.050 215.250 ;
        RECT 574.950 207.300 578.850 209.400 ;
        RECT 585.150 208.500 586.950 215.250 ;
        RECT 588.150 209.400 589.950 215.250 ;
        RECT 592.950 209.400 594.750 215.250 ;
        RECT 598.050 209.400 599.850 215.250 ;
        RECT 593.250 208.500 594.450 209.400 ;
        RECT 583.950 206.700 590.850 208.500 ;
        RECT 593.250 206.400 598.050 208.500 ;
        RECT 576.150 204.600 578.850 206.400 ;
        RECT 579.750 205.800 581.550 206.400 ;
        RECT 579.750 204.900 586.050 205.800 ;
        RECT 593.250 205.500 594.450 206.400 ;
        RECT 579.750 204.600 581.550 204.900 ;
        RECT 577.950 203.700 578.850 204.600 ;
        RECT 560.100 195.150 561.900 196.950 ;
        RECT 500.850 191.100 511.950 192.000 ;
        RECT 520.950 191.850 525.450 193.950 ;
        RECT 500.850 190.200 501.900 191.100 ;
        RECT 511.050 190.800 511.950 191.100 ;
        RECT 479.100 187.950 484.800 189.600 ;
        RECT 466.650 183.750 468.450 186.600 ;
        RECT 469.650 183.750 471.450 186.600 ;
        RECT 472.650 183.750 474.450 186.600 ;
        RECT 479.700 183.750 481.500 186.600 ;
        RECT 483.000 183.750 484.800 187.950 ;
        RECT 487.200 183.750 489.000 189.600 ;
        RECT 492.150 183.750 493.950 189.600 ;
        RECT 496.950 187.500 499.050 189.600 ;
        RECT 500.550 188.400 502.350 190.200 ;
        RECT 503.850 189.450 505.650 190.200 ;
        RECT 503.850 188.400 508.800 189.450 ;
        RECT 511.050 189.000 512.850 190.800 ;
        RECT 524.250 189.600 525.450 191.850 ;
        RECT 517.950 188.700 520.050 189.600 ;
        RECT 498.000 186.600 499.050 187.500 ;
        RECT 507.750 186.600 508.800 188.400 ;
        RECT 516.300 187.500 520.050 188.700 ;
        RECT 516.300 186.600 517.350 187.500 ;
        RECT 495.150 183.750 496.950 186.600 ;
        RECT 498.000 185.700 501.750 186.600 ;
        RECT 499.950 183.750 501.750 185.700 ;
        RECT 504.450 183.750 506.250 186.600 ;
        RECT 507.750 183.750 509.550 186.600 ;
        RECT 511.650 183.750 513.450 186.600 ;
        RECT 515.850 183.750 517.650 186.600 ;
        RECT 520.350 183.750 522.150 186.600 ;
        RECT 523.650 183.750 525.450 189.600 ;
        RECT 530.400 186.600 531.600 194.850 ;
        RECT 532.950 193.050 535.050 195.150 ;
        RECT 541.950 193.050 544.050 195.150 ;
        RECT 553.950 193.050 556.050 195.150 ;
        RECT 559.950 193.050 562.050 195.150 ;
        RECT 562.950 194.850 565.050 196.950 ;
        RECT 541.950 186.600 543.000 193.050 ;
        RECT 553.950 186.600 555.000 193.050 ;
        RECT 563.400 186.600 564.600 194.850 ;
        RECT 569.550 193.950 570.750 203.400 ;
        RECT 574.950 202.800 577.050 203.700 ;
        RECT 577.950 202.800 583.950 203.700 ;
        RECT 572.850 201.600 577.050 202.800 ;
        RECT 571.950 199.800 573.750 201.600 ;
        RECT 583.050 198.150 583.950 202.800 ;
        RECT 585.150 202.800 586.050 204.900 ;
        RECT 586.950 204.300 594.450 205.500 ;
        RECT 586.950 203.700 588.750 204.300 ;
        RECT 601.050 203.400 602.850 215.250 ;
        RECT 606.300 203.400 608.100 215.250 ;
        RECT 610.500 203.400 612.300 215.250 ;
        RECT 613.800 209.400 615.600 215.250 ;
        RECT 620.550 209.400 622.350 215.250 ;
        RECT 623.550 209.400 625.350 215.250 ;
        RECT 626.550 209.400 628.350 215.250 ;
        RECT 591.750 202.800 602.850 203.400 ;
        RECT 585.150 202.200 602.850 202.800 ;
        RECT 585.150 201.900 593.550 202.200 ;
        RECT 591.750 201.600 593.550 201.900 ;
        RECT 583.050 196.050 586.050 198.150 ;
        RECT 589.950 197.100 592.050 198.150 ;
        RECT 589.950 196.050 597.900 197.100 ;
        RECT 571.950 195.750 574.050 196.050 ;
        RECT 571.950 193.950 575.850 195.750 ;
        RECT 569.550 191.850 574.050 193.950 ;
        RECT 583.050 192.000 583.950 196.050 ;
        RECT 596.100 195.300 597.900 196.050 ;
        RECT 599.100 195.150 600.900 196.950 ;
        RECT 593.100 194.400 594.900 195.000 ;
        RECT 599.100 194.400 600.000 195.150 ;
        RECT 593.100 193.200 600.000 194.400 ;
        RECT 593.100 192.000 594.150 193.200 ;
        RECT 569.550 189.600 570.750 191.850 ;
        RECT 583.050 191.100 594.150 192.000 ;
        RECT 583.050 190.800 583.950 191.100 ;
        RECT 529.650 183.750 531.450 186.600 ;
        RECT 532.650 183.750 534.450 186.600 ;
        RECT 538.650 183.750 540.450 186.600 ;
        RECT 541.650 183.750 543.450 186.600 ;
        RECT 544.650 183.750 546.450 186.600 ;
        RECT 550.650 183.750 552.450 186.600 ;
        RECT 553.650 183.750 555.450 186.600 ;
        RECT 556.650 183.750 558.450 186.600 ;
        RECT 560.550 183.750 562.350 186.600 ;
        RECT 563.550 183.750 565.350 186.600 ;
        RECT 569.550 183.750 571.350 189.600 ;
        RECT 574.950 188.700 577.050 189.600 ;
        RECT 582.150 189.000 583.950 190.800 ;
        RECT 593.100 190.200 594.150 191.100 ;
        RECT 589.350 189.450 591.150 190.200 ;
        RECT 574.950 187.500 578.700 188.700 ;
        RECT 577.650 186.600 578.700 187.500 ;
        RECT 586.200 188.400 591.150 189.450 ;
        RECT 592.650 188.400 594.450 190.200 ;
        RECT 601.950 189.600 602.850 202.200 ;
        RECT 605.100 198.150 606.900 199.950 ;
        RECT 610.950 198.150 612.150 203.400 ;
        RECT 613.950 201.150 615.750 202.950 ;
        RECT 623.550 201.150 624.750 209.400 ;
        RECT 634.350 203.400 636.150 215.250 ;
        RECT 637.350 203.400 639.150 215.250 ;
        RECT 640.650 209.400 642.450 215.250 ;
        RECT 646.650 209.400 648.450 215.250 ;
        RECT 649.650 209.400 651.450 215.250 ;
        RECT 652.650 209.400 654.450 215.250 ;
        RECT 659.400 209.400 661.200 215.250 ;
        RECT 613.950 199.050 616.050 201.150 ;
        RECT 604.950 196.050 607.050 198.150 ;
        RECT 607.950 194.850 610.050 196.950 ;
        RECT 610.950 196.050 613.050 198.150 ;
        RECT 619.950 197.850 622.050 199.950 ;
        RECT 622.950 199.050 625.050 201.150 ;
        RECT 620.100 196.050 621.900 197.850 ;
        RECT 608.100 193.050 609.900 194.850 ;
        RECT 611.850 192.750 613.050 196.050 ;
        RECT 612.000 191.700 615.750 192.750 ;
        RECT 586.200 186.600 587.250 188.400 ;
        RECT 595.950 187.500 598.050 189.600 ;
        RECT 595.950 186.600 597.000 187.500 ;
        RECT 572.850 183.750 574.650 186.600 ;
        RECT 577.350 183.750 579.150 186.600 ;
        RECT 581.550 183.750 583.350 186.600 ;
        RECT 585.450 183.750 587.250 186.600 ;
        RECT 588.750 183.750 590.550 186.600 ;
        RECT 593.250 185.700 597.000 186.600 ;
        RECT 593.250 183.750 595.050 185.700 ;
        RECT 598.050 183.750 599.850 186.600 ;
        RECT 601.050 183.750 602.850 189.600 ;
        RECT 605.550 188.700 613.350 190.050 ;
        RECT 605.550 183.750 607.350 188.700 ;
        RECT 608.550 183.750 610.350 187.800 ;
        RECT 611.550 183.750 613.350 188.700 ;
        RECT 614.550 189.600 615.750 191.700 ;
        RECT 623.550 191.700 624.750 199.050 ;
        RECT 625.950 197.850 628.050 199.950 ;
        RECT 634.650 198.150 635.850 203.400 ;
        RECT 641.250 202.500 642.450 209.400 ;
        RECT 636.750 201.600 642.450 202.500 ;
        RECT 636.750 200.700 639.000 201.600 ;
        RECT 650.250 201.150 651.450 209.400 ;
        RECT 662.700 203.400 664.500 215.250 ;
        RECT 666.900 203.400 668.700 215.250 ;
        RECT 674.400 209.400 676.200 215.250 ;
        RECT 677.700 203.400 679.500 215.250 ;
        RECT 681.900 203.400 683.700 215.250 ;
        RECT 686.550 203.400 688.350 215.250 ;
        RECT 690.750 203.400 692.550 215.250 ;
        RECT 698.550 209.400 700.350 215.250 ;
        RECT 701.550 209.400 703.350 215.250 ;
        RECT 709.650 209.400 711.450 215.250 ;
        RECT 712.650 209.400 714.450 215.250 ;
        RECT 659.250 201.150 661.050 202.950 ;
        RECT 626.100 196.050 627.900 197.850 ;
        RECT 634.650 196.050 637.050 198.150 ;
        RECT 623.550 190.800 627.150 191.700 ;
        RECT 614.550 183.750 616.350 189.600 ;
        RECT 620.850 183.750 622.650 189.600 ;
        RECT 625.350 183.750 627.150 190.800 ;
        RECT 634.650 189.600 635.850 196.050 ;
        RECT 637.950 192.300 639.000 200.700 ;
        RECT 641.100 198.150 642.900 199.950 ;
        RECT 640.950 196.050 643.050 198.150 ;
        RECT 646.950 197.850 649.050 199.950 ;
        RECT 649.950 199.050 652.050 201.150 ;
        RECT 647.100 196.050 648.900 197.850 ;
        RECT 636.750 191.400 639.000 192.300 ;
        RECT 650.250 191.700 651.450 199.050 ;
        RECT 652.950 197.850 655.050 199.950 ;
        RECT 658.950 199.050 661.050 201.150 ;
        RECT 662.850 198.150 664.050 203.400 ;
        RECT 674.250 201.150 676.050 202.950 ;
        RECT 668.100 198.150 669.900 199.950 ;
        RECT 673.950 199.050 676.050 201.150 ;
        RECT 677.850 198.150 679.050 203.400 ;
        RECT 690.000 202.350 692.550 203.400 ;
        RECT 683.100 198.150 684.900 199.950 ;
        RECT 686.100 198.150 687.900 199.950 ;
        RECT 653.100 196.050 654.900 197.850 ;
        RECT 661.950 196.050 664.050 198.150 ;
        RECT 661.950 192.750 663.150 196.050 ;
        RECT 664.950 194.850 667.050 196.950 ;
        RECT 667.950 196.050 670.050 198.150 ;
        RECT 676.950 196.050 679.050 198.150 ;
        RECT 665.100 193.050 666.900 194.850 ;
        RECT 676.950 192.750 678.150 196.050 ;
        RECT 679.950 194.850 682.050 196.950 ;
        RECT 682.950 196.050 685.050 198.150 ;
        RECT 685.950 196.050 688.050 198.150 ;
        RECT 690.000 195.150 691.050 202.350 ;
        RECT 692.100 198.150 693.900 199.950 ;
        RECT 691.950 196.050 694.050 198.150 ;
        RECT 701.400 196.950 702.600 209.400 ;
        RECT 710.400 196.950 711.600 209.400 ;
        RECT 698.100 195.150 699.900 196.950 ;
        RECT 680.100 193.050 681.900 194.850 ;
        RECT 688.950 193.050 691.050 195.150 ;
        RECT 697.950 193.050 700.050 195.150 ;
        RECT 700.950 194.850 703.050 196.950 ;
        RECT 709.950 194.850 712.050 196.950 ;
        RECT 713.100 195.150 714.900 196.950 ;
        RECT 636.750 190.500 641.850 191.400 ;
        RECT 634.350 183.750 636.150 189.600 ;
        RECT 637.350 183.750 639.150 189.600 ;
        RECT 640.650 186.600 641.850 190.500 ;
        RECT 647.850 190.800 651.450 191.700 ;
        RECT 659.250 191.700 663.000 192.750 ;
        RECT 674.250 191.700 678.000 192.750 ;
        RECT 640.650 183.750 642.450 186.600 ;
        RECT 647.850 183.750 649.650 190.800 ;
        RECT 659.250 189.600 660.450 191.700 ;
        RECT 652.350 183.750 654.150 189.600 ;
        RECT 658.650 183.750 660.450 189.600 ;
        RECT 661.650 188.700 669.450 190.050 ;
        RECT 674.250 189.600 675.450 191.700 ;
        RECT 661.650 183.750 663.450 188.700 ;
        RECT 664.650 183.750 666.450 187.800 ;
        RECT 667.650 183.750 669.450 188.700 ;
        RECT 673.650 183.750 675.450 189.600 ;
        RECT 676.650 188.700 684.450 190.050 ;
        RECT 676.650 183.750 678.450 188.700 ;
        RECT 679.650 183.750 681.450 187.800 ;
        RECT 682.650 183.750 684.450 188.700 ;
        RECT 690.000 186.600 691.050 193.050 ;
        RECT 701.400 186.600 702.600 194.850 ;
        RECT 710.400 186.600 711.600 194.850 ;
        RECT 712.950 193.050 715.050 195.150 ;
        RECT 686.550 183.750 688.350 186.600 ;
        RECT 689.550 183.750 691.350 186.600 ;
        RECT 692.550 183.750 694.350 186.600 ;
        RECT 698.550 183.750 700.350 186.600 ;
        RECT 701.550 183.750 703.350 186.600 ;
        RECT 709.650 183.750 711.450 186.600 ;
        RECT 712.650 183.750 714.450 186.600 ;
        RECT 4.650 173.400 6.450 179.250 ;
        RECT 5.250 171.300 6.450 173.400 ;
        RECT 7.650 174.300 9.450 179.250 ;
        RECT 10.650 175.200 12.450 179.250 ;
        RECT 13.650 174.300 15.450 179.250 ;
        RECT 7.650 172.950 15.450 174.300 ;
        RECT 17.550 174.300 19.350 179.250 ;
        RECT 20.550 175.200 22.350 179.250 ;
        RECT 23.550 174.300 25.350 179.250 ;
        RECT 17.550 172.950 25.350 174.300 ;
        RECT 26.550 173.400 28.350 179.250 ;
        RECT 26.550 171.300 27.750 173.400 ;
        RECT 5.250 170.250 9.000 171.300 ;
        RECT 24.000 170.250 27.750 171.300 ;
        RECT 32.700 170.400 34.500 179.250 ;
        RECT 38.100 171.000 39.900 179.250 ;
        RECT 48.000 173.400 49.800 179.250 ;
        RECT 52.200 175.050 54.000 179.250 ;
        RECT 55.500 176.400 57.300 179.250 ;
        RECT 52.200 173.400 57.900 175.050 ;
        RECT 7.950 166.950 9.150 170.250 ;
        RECT 11.100 168.150 12.900 169.950 ;
        RECT 20.100 168.150 21.900 169.950 ;
        RECT 7.950 164.850 10.050 166.950 ;
        RECT 10.950 166.050 13.050 168.150 ;
        RECT 13.950 164.850 16.050 166.950 ;
        RECT 16.950 164.850 19.050 166.950 ;
        RECT 19.950 166.050 22.050 168.150 ;
        RECT 23.850 166.950 25.050 170.250 ;
        RECT 38.100 169.350 42.600 171.000 ;
        RECT 43.950 169.950 46.050 172.050 ;
        RECT 22.950 164.850 25.050 166.950 ;
        RECT 41.400 165.150 42.600 169.350 ;
        RECT 4.950 161.850 7.050 163.950 ;
        RECT 5.250 160.050 7.050 161.850 ;
        RECT 8.850 159.600 10.050 164.850 ;
        RECT 14.100 163.050 15.900 164.850 ;
        RECT 17.100 163.050 18.900 164.850 ;
        RECT 22.950 159.600 24.150 164.850 ;
        RECT 25.950 161.850 28.050 163.950 ;
        RECT 31.950 161.850 34.050 163.950 ;
        RECT 37.950 161.850 40.050 163.950 ;
        RECT 40.950 163.050 43.050 165.150 ;
        RECT 44.550 163.050 45.450 169.950 ;
        RECT 47.100 168.150 48.900 169.950 ;
        RECT 46.950 166.050 49.050 168.150 ;
        RECT 49.950 167.850 52.050 169.950 ;
        RECT 53.100 168.150 54.900 169.950 ;
        RECT 50.100 166.050 51.900 167.850 ;
        RECT 52.950 166.050 55.050 168.150 ;
        RECT 56.700 166.950 57.900 173.400 ;
        RECT 62.700 170.400 64.500 179.250 ;
        RECT 68.100 171.000 69.900 179.250 ;
        RECT 70.950 174.450 73.050 175.050 ;
        RECT 70.950 173.550 75.450 174.450 ;
        RECT 70.950 172.950 73.050 173.550 ;
        RECT 68.100 169.350 72.600 171.000 ;
        RECT 55.950 164.850 58.050 166.950 ;
        RECT 71.400 165.150 72.600 169.350 ;
        RECT 25.950 160.050 27.750 161.850 ;
        RECT 32.100 160.050 33.900 161.850 ;
        RECT 5.400 147.750 7.200 153.600 ;
        RECT 8.700 147.750 10.500 159.600 ;
        RECT 12.900 147.750 14.700 159.600 ;
        RECT 18.300 147.750 20.100 159.600 ;
        RECT 22.500 147.750 24.300 159.600 ;
        RECT 34.950 158.850 37.050 160.950 ;
        RECT 38.250 160.050 40.050 161.850 ;
        RECT 35.100 157.050 36.900 158.850 ;
        RECT 41.700 154.800 42.750 163.050 ;
        RECT 43.950 160.950 46.050 163.050 ;
        RECT 56.700 159.600 57.900 164.850 ;
        RECT 61.950 161.850 64.050 163.950 ;
        RECT 67.950 161.850 70.050 163.950 ;
        RECT 70.950 163.050 73.050 165.150 ;
        RECT 62.100 160.050 63.900 161.850 ;
        RECT 35.700 153.900 42.750 154.800 ;
        RECT 35.700 153.600 37.350 153.900 ;
        RECT 25.800 147.750 27.600 153.600 ;
        RECT 32.550 147.750 34.350 153.600 ;
        RECT 35.550 147.750 37.350 153.600 ;
        RECT 41.550 153.600 42.750 153.900 ;
        RECT 47.550 158.700 55.350 159.600 ;
        RECT 38.550 147.750 40.350 153.000 ;
        RECT 41.550 147.750 43.350 153.600 ;
        RECT 47.550 147.750 49.350 158.700 ;
        RECT 50.550 147.750 52.350 157.800 ;
        RECT 53.550 147.750 55.350 158.700 ;
        RECT 56.550 147.750 58.350 159.600 ;
        RECT 64.950 158.850 67.050 160.950 ;
        RECT 68.250 160.050 70.050 161.850 ;
        RECT 65.100 157.050 66.900 158.850 ;
        RECT 71.700 154.800 72.750 163.050 ;
        RECT 74.550 162.450 75.450 173.550 ;
        RECT 78.000 173.400 79.800 179.250 ;
        RECT 82.200 175.050 84.000 179.250 ;
        RECT 85.500 176.400 87.300 179.250 ;
        RECT 82.200 173.400 87.900 175.050 ;
        RECT 77.100 168.150 78.900 169.950 ;
        RECT 76.950 166.050 79.050 168.150 ;
        RECT 79.950 167.850 82.050 169.950 ;
        RECT 83.100 168.150 84.900 169.950 ;
        RECT 80.100 166.050 81.900 167.850 ;
        RECT 82.950 166.050 85.050 168.150 ;
        RECT 86.700 166.950 87.900 173.400 ;
        RECT 95.850 172.200 97.650 179.250 ;
        RECT 100.350 173.400 102.150 179.250 ;
        RECT 108.150 174.900 109.950 179.250 ;
        RECT 106.650 173.400 109.950 174.900 ;
        RECT 111.150 173.400 112.950 179.250 ;
        RECT 95.850 171.300 99.450 172.200 ;
        RECT 85.950 164.850 88.050 166.950 ;
        RECT 95.100 165.150 96.900 166.950 ;
        RECT 76.950 162.450 79.050 163.050 ;
        RECT 74.550 161.550 79.050 162.450 ;
        RECT 76.950 160.950 79.050 161.550 ;
        RECT 86.700 159.600 87.900 164.850 ;
        RECT 94.950 163.050 97.050 165.150 ;
        RECT 98.250 163.950 99.450 171.300 ;
        RECT 106.650 166.950 107.850 173.400 ;
        RECT 109.950 171.900 111.750 172.500 ;
        RECT 115.650 171.900 117.450 179.250 ;
        RECT 109.950 170.700 117.450 171.900 ;
        RECT 125.100 171.000 126.900 179.250 ;
        RECT 101.100 165.150 102.900 166.950 ;
        RECT 97.950 161.850 100.050 163.950 ;
        RECT 100.950 163.050 103.050 165.150 ;
        RECT 106.650 164.850 109.050 166.950 ;
        RECT 110.100 165.150 111.900 166.950 ;
        RECT 65.700 153.900 72.750 154.800 ;
        RECT 65.700 153.600 67.350 153.900 ;
        RECT 62.550 147.750 64.350 153.600 ;
        RECT 65.550 147.750 67.350 153.600 ;
        RECT 71.550 153.600 72.750 153.900 ;
        RECT 77.550 158.700 85.350 159.600 ;
        RECT 68.550 147.750 70.350 153.000 ;
        RECT 71.550 147.750 73.350 153.600 ;
        RECT 77.550 147.750 79.350 158.700 ;
        RECT 80.550 147.750 82.350 157.800 ;
        RECT 83.550 147.750 85.350 158.700 ;
        RECT 86.550 147.750 88.350 159.600 ;
        RECT 98.250 153.600 99.450 161.850 ;
        RECT 106.650 159.600 107.850 164.850 ;
        RECT 109.950 163.050 112.050 165.150 ;
        RECT 94.650 147.750 96.450 153.600 ;
        RECT 97.650 147.750 99.450 153.600 ;
        RECT 100.650 147.750 102.450 153.600 ;
        RECT 106.050 147.750 107.850 159.600 ;
        RECT 109.050 147.750 110.850 159.600 ;
        RECT 113.100 153.600 114.300 170.700 ;
        RECT 122.400 169.350 126.900 171.000 ;
        RECT 130.500 170.400 132.300 179.250 ;
        RECT 136.650 173.400 138.450 179.250 ;
        RECT 137.250 171.300 138.450 173.400 ;
        RECT 139.650 174.300 141.450 179.250 ;
        RECT 142.650 175.200 144.450 179.250 ;
        RECT 145.650 174.300 147.450 179.250 ;
        RECT 139.650 172.950 147.450 174.300 ;
        RECT 149.550 174.300 151.350 179.250 ;
        RECT 152.550 175.200 154.350 179.250 ;
        RECT 155.550 174.300 157.350 179.250 ;
        RECT 149.550 172.950 157.350 174.300 ;
        RECT 158.550 173.400 160.350 179.250 ;
        RECT 166.650 173.400 168.450 179.250 ;
        RECT 158.550 171.300 159.750 173.400 ;
        RECT 137.250 170.250 141.000 171.300 ;
        RECT 156.000 170.250 159.750 171.300 ;
        RECT 167.250 171.300 168.450 173.400 ;
        RECT 169.650 174.300 171.450 179.250 ;
        RECT 172.650 175.200 174.450 179.250 ;
        RECT 175.650 174.300 177.450 179.250 ;
        RECT 169.650 172.950 177.450 174.300 ;
        RECT 182.850 172.200 184.650 179.250 ;
        RECT 187.350 173.400 189.150 179.250 ;
        RECT 195.150 174.900 196.950 179.250 ;
        RECT 193.650 173.400 196.950 174.900 ;
        RECT 198.150 173.400 199.950 179.250 ;
        RECT 182.850 171.300 186.450 172.200 ;
        RECT 167.250 170.250 171.000 171.300 ;
        RECT 115.950 164.850 118.050 166.950 ;
        RECT 122.400 165.150 123.600 169.350 ;
        RECT 127.950 168.450 130.050 169.050 ;
        RECT 127.950 167.550 135.450 168.450 ;
        RECT 127.950 166.950 130.050 167.550 ;
        RECT 116.100 163.050 117.900 164.850 ;
        RECT 121.950 163.050 124.050 165.150 ;
        RECT 122.250 154.800 123.300 163.050 ;
        RECT 124.950 161.850 127.050 163.950 ;
        RECT 130.950 161.850 133.050 163.950 ;
        RECT 124.950 160.050 126.750 161.850 ;
        RECT 127.950 158.850 130.050 160.950 ;
        RECT 131.100 160.050 132.900 161.850 ;
        RECT 128.100 157.050 129.900 158.850 ;
        RECT 134.550 157.050 135.450 167.550 ;
        RECT 139.950 166.950 141.150 170.250 ;
        RECT 143.100 168.150 144.900 169.950 ;
        RECT 152.100 168.150 153.900 169.950 ;
        RECT 139.950 164.850 142.050 166.950 ;
        RECT 142.950 166.050 145.050 168.150 ;
        RECT 145.950 164.850 148.050 166.950 ;
        RECT 148.950 164.850 151.050 166.950 ;
        RECT 151.950 166.050 154.050 168.150 ;
        RECT 155.850 166.950 157.050 170.250 ;
        RECT 154.950 164.850 157.050 166.950 ;
        RECT 169.950 166.950 171.150 170.250 ;
        RECT 173.100 168.150 174.900 169.950 ;
        RECT 169.950 164.850 172.050 166.950 ;
        RECT 172.950 166.050 175.050 168.150 ;
        RECT 175.950 164.850 178.050 166.950 ;
        RECT 182.100 165.150 183.900 166.950 ;
        RECT 136.950 161.850 139.050 163.950 ;
        RECT 137.250 160.050 139.050 161.850 ;
        RECT 140.850 159.600 142.050 164.850 ;
        RECT 146.100 163.050 147.900 164.850 ;
        RECT 149.100 163.050 150.900 164.850 ;
        RECT 154.950 159.600 156.150 164.850 ;
        RECT 157.950 161.850 160.050 163.950 ;
        RECT 166.950 161.850 169.050 163.950 ;
        RECT 157.950 160.050 159.750 161.850 ;
        RECT 167.250 160.050 169.050 161.850 ;
        RECT 170.850 159.600 172.050 164.850 ;
        RECT 176.100 163.050 177.900 164.850 ;
        RECT 181.950 163.050 184.050 165.150 ;
        RECT 185.250 163.950 186.450 171.300 ;
        RECT 193.650 166.950 194.850 173.400 ;
        RECT 196.950 171.900 198.750 172.500 ;
        RECT 202.650 171.900 204.450 179.250 ;
        RECT 206.850 173.400 208.650 179.250 ;
        RECT 211.350 172.200 213.150 179.250 ;
        RECT 220.650 173.400 222.450 179.250 ;
        RECT 223.650 173.400 225.450 179.250 ;
        RECT 196.950 170.700 204.450 171.900 ;
        RECT 209.550 171.300 213.150 172.200 ;
        RECT 188.100 165.150 189.900 166.950 ;
        RECT 184.950 161.850 187.050 163.950 ;
        RECT 187.950 163.050 190.050 165.150 ;
        RECT 193.650 164.850 196.050 166.950 ;
        RECT 197.100 165.150 198.900 166.950 ;
        RECT 133.950 154.950 136.050 157.050 ;
        RECT 122.250 153.900 129.300 154.800 ;
        RECT 122.250 153.600 123.450 153.900 ;
        RECT 112.650 147.750 114.450 153.600 ;
        RECT 115.650 147.750 117.450 153.600 ;
        RECT 121.650 147.750 123.450 153.600 ;
        RECT 127.650 153.600 129.300 153.900 ;
        RECT 124.650 147.750 126.450 153.000 ;
        RECT 127.650 147.750 129.450 153.600 ;
        RECT 130.650 147.750 132.450 153.600 ;
        RECT 137.400 147.750 139.200 153.600 ;
        RECT 140.700 147.750 142.500 159.600 ;
        RECT 144.900 147.750 146.700 159.600 ;
        RECT 150.300 147.750 152.100 159.600 ;
        RECT 154.500 147.750 156.300 159.600 ;
        RECT 157.800 147.750 159.600 153.600 ;
        RECT 167.400 147.750 169.200 153.600 ;
        RECT 170.700 147.750 172.500 159.600 ;
        RECT 174.900 147.750 176.700 159.600 ;
        RECT 185.250 153.600 186.450 161.850 ;
        RECT 193.650 159.600 194.850 164.850 ;
        RECT 196.950 163.050 199.050 165.150 ;
        RECT 181.650 147.750 183.450 153.600 ;
        RECT 184.650 147.750 186.450 153.600 ;
        RECT 187.650 147.750 189.450 153.600 ;
        RECT 193.050 147.750 194.850 159.600 ;
        RECT 196.050 147.750 197.850 159.600 ;
        RECT 200.100 153.600 201.300 170.700 ;
        RECT 202.950 164.850 205.050 166.950 ;
        RECT 206.100 165.150 207.900 166.950 ;
        RECT 203.100 163.050 204.900 164.850 ;
        RECT 205.950 163.050 208.050 165.150 ;
        RECT 209.550 163.950 210.750 171.300 ;
        RECT 221.400 166.950 222.600 173.400 ;
        RECT 230.850 172.200 232.650 179.250 ;
        RECT 235.350 173.400 237.150 179.250 ;
        RECT 242.850 172.200 244.650 179.250 ;
        RECT 247.350 173.400 249.150 179.250 ;
        RECT 230.850 171.300 234.450 172.200 ;
        RECT 224.100 168.150 225.900 169.950 ;
        RECT 212.100 165.150 213.900 166.950 ;
        RECT 208.950 161.850 211.050 163.950 ;
        RECT 211.950 163.050 214.050 165.150 ;
        RECT 220.950 164.850 223.050 166.950 ;
        RECT 223.950 166.050 226.050 168.150 ;
        RECT 230.100 165.150 231.900 166.950 ;
        RECT 209.550 153.600 210.750 161.850 ;
        RECT 221.400 159.600 222.600 164.850 ;
        RECT 229.950 163.050 232.050 165.150 ;
        RECT 233.250 163.950 234.450 171.300 ;
        RECT 235.950 171.450 238.050 172.050 ;
        RECT 235.950 170.550 240.450 171.450 ;
        RECT 242.850 171.300 246.450 172.200 ;
        RECT 235.950 169.950 238.050 170.550 ;
        RECT 236.100 165.150 237.900 166.950 ;
        RECT 232.950 161.850 235.050 163.950 ;
        RECT 235.950 163.050 238.050 165.150 ;
        RECT 199.650 147.750 201.450 153.600 ;
        RECT 202.650 147.750 204.450 153.600 ;
        RECT 206.550 147.750 208.350 153.600 ;
        RECT 209.550 147.750 211.350 153.600 ;
        RECT 212.550 147.750 214.350 153.600 ;
        RECT 220.650 147.750 222.450 159.600 ;
        RECT 223.650 147.750 225.450 159.600 ;
        RECT 233.250 153.600 234.450 161.850 ;
        RECT 239.550 159.450 240.450 170.550 ;
        RECT 242.100 165.150 243.900 166.950 ;
        RECT 241.950 163.050 244.050 165.150 ;
        RECT 245.250 163.950 246.450 171.300 ;
        RECT 251.700 170.400 253.500 179.250 ;
        RECT 257.100 171.000 258.900 179.250 ;
        RECT 269.850 172.200 271.650 179.250 ;
        RECT 274.350 173.400 276.150 179.250 ;
        RECT 269.850 171.300 273.450 172.200 ;
        RECT 257.100 169.350 261.600 171.000 ;
        RECT 248.100 165.150 249.900 166.950 ;
        RECT 260.400 165.150 261.600 169.350 ;
        RECT 269.100 165.150 270.900 166.950 ;
        RECT 244.950 161.850 247.050 163.950 ;
        RECT 247.950 163.050 250.050 165.150 ;
        RECT 250.950 161.850 253.050 163.950 ;
        RECT 256.950 161.850 259.050 163.950 ;
        RECT 259.950 163.050 262.050 165.150 ;
        RECT 268.950 163.050 271.050 165.150 ;
        RECT 272.250 163.950 273.450 171.300 ;
        RECT 278.700 170.400 280.500 179.250 ;
        RECT 284.100 171.000 285.900 179.250 ;
        RECT 293.850 173.400 295.650 179.250 ;
        RECT 298.350 172.200 300.150 179.250 ;
        RECT 310.800 173.400 312.600 179.250 ;
        RECT 315.000 173.400 316.800 179.250 ;
        RECT 319.200 173.400 321.000 179.250 ;
        RECT 296.550 171.300 300.150 172.200 ;
        RECT 284.100 169.350 288.600 171.000 ;
        RECT 275.100 165.150 276.900 166.950 ;
        RECT 287.400 165.150 288.600 169.350 ;
        RECT 293.100 165.150 294.900 166.950 ;
        RECT 239.550 158.550 243.450 159.450 ;
        RECT 242.550 157.050 243.450 158.550 ;
        RECT 241.950 154.950 244.050 157.050 ;
        RECT 245.250 153.600 246.450 161.850 ;
        RECT 251.100 160.050 252.900 161.850 ;
        RECT 253.950 158.850 256.050 160.950 ;
        RECT 257.250 160.050 259.050 161.850 ;
        RECT 254.100 157.050 255.900 158.850 ;
        RECT 260.700 154.800 261.750 163.050 ;
        RECT 271.950 161.850 274.050 163.950 ;
        RECT 274.950 163.050 277.050 165.150 ;
        RECT 277.950 161.850 280.050 163.950 ;
        RECT 283.950 161.850 286.050 163.950 ;
        RECT 286.950 163.050 289.050 165.150 ;
        RECT 292.950 163.050 295.050 165.150 ;
        RECT 296.550 163.950 297.750 171.300 ;
        RECT 311.250 168.150 313.050 169.950 ;
        RECT 299.100 165.150 300.900 166.950 ;
        RECT 254.700 153.900 261.750 154.800 ;
        RECT 254.700 153.600 256.350 153.900 ;
        RECT 229.650 147.750 231.450 153.600 ;
        RECT 232.650 147.750 234.450 153.600 ;
        RECT 235.650 147.750 237.450 153.600 ;
        RECT 241.650 147.750 243.450 153.600 ;
        RECT 244.650 147.750 246.450 153.600 ;
        RECT 247.650 147.750 249.450 153.600 ;
        RECT 251.550 147.750 253.350 153.600 ;
        RECT 254.550 147.750 256.350 153.600 ;
        RECT 260.550 153.600 261.750 153.900 ;
        RECT 272.250 153.600 273.450 161.850 ;
        RECT 278.100 160.050 279.900 161.850 ;
        RECT 280.950 158.850 283.050 160.950 ;
        RECT 284.250 160.050 286.050 161.850 ;
        RECT 281.100 157.050 282.900 158.850 ;
        RECT 287.700 154.800 288.750 163.050 ;
        RECT 295.950 161.850 298.050 163.950 ;
        RECT 298.950 163.050 301.050 165.150 ;
        RECT 307.950 164.850 310.050 166.950 ;
        RECT 310.950 166.050 313.050 168.150 ;
        RECT 315.000 166.950 316.050 173.400 ;
        RECT 329.100 171.000 330.900 179.250 ;
        RECT 313.950 164.850 316.050 166.950 ;
        RECT 316.950 168.150 318.750 169.950 ;
        RECT 326.400 169.350 330.900 171.000 ;
        RECT 334.500 170.400 336.300 179.250 ;
        RECT 341.850 172.200 343.650 179.250 ;
        RECT 346.350 173.400 348.150 179.250 ;
        RECT 351.000 173.400 352.800 179.250 ;
        RECT 355.200 175.050 357.000 179.250 ;
        RECT 358.500 176.400 360.300 179.250 ;
        RECT 367.650 176.400 369.450 179.250 ;
        RECT 370.650 176.400 372.450 179.250 ;
        RECT 355.200 173.400 360.900 175.050 ;
        RECT 341.850 171.300 345.450 172.200 ;
        RECT 316.950 166.050 319.050 168.150 ;
        RECT 319.950 164.850 322.050 166.950 ;
        RECT 326.400 165.150 327.600 169.350 ;
        RECT 331.950 168.450 334.050 169.050 ;
        RECT 331.950 167.550 339.450 168.450 ;
        RECT 331.950 166.950 334.050 167.550 ;
        RECT 308.100 163.050 309.900 164.850 ;
        RECT 281.700 153.900 288.750 154.800 ;
        RECT 281.700 153.600 283.350 153.900 ;
        RECT 257.550 147.750 259.350 153.000 ;
        RECT 260.550 147.750 262.350 153.600 ;
        RECT 268.650 147.750 270.450 153.600 ;
        RECT 271.650 147.750 273.450 153.600 ;
        RECT 274.650 147.750 276.450 153.600 ;
        RECT 278.550 147.750 280.350 153.600 ;
        RECT 281.550 147.750 283.350 153.600 ;
        RECT 287.550 153.600 288.750 153.900 ;
        RECT 296.550 153.600 297.750 161.850 ;
        RECT 313.950 161.400 314.850 164.850 ;
        RECT 319.950 163.050 321.750 164.850 ;
        RECT 325.950 163.050 328.050 165.150 ;
        RECT 310.800 160.500 314.850 161.400 ;
        RECT 310.800 159.600 312.600 160.500 ;
        RECT 284.550 147.750 286.350 153.000 ;
        RECT 287.550 147.750 289.350 153.600 ;
        RECT 293.550 147.750 295.350 153.600 ;
        RECT 296.550 147.750 298.350 153.600 ;
        RECT 299.550 147.750 301.350 153.600 ;
        RECT 307.650 148.500 309.450 159.600 ;
        RECT 310.650 149.400 312.450 159.600 ;
        RECT 313.650 158.400 321.450 159.300 ;
        RECT 313.650 148.500 315.450 158.400 ;
        RECT 307.650 147.750 315.450 148.500 ;
        RECT 316.650 147.750 318.450 157.500 ;
        RECT 319.650 147.750 321.450 158.400 ;
        RECT 326.250 154.800 327.300 163.050 ;
        RECT 328.950 161.850 331.050 163.950 ;
        RECT 334.950 161.850 337.050 163.950 ;
        RECT 328.950 160.050 330.750 161.850 ;
        RECT 331.950 158.850 334.050 160.950 ;
        RECT 335.100 160.050 336.900 161.850 ;
        RECT 338.550 159.450 339.450 167.550 ;
        RECT 341.100 165.150 342.900 166.950 ;
        RECT 340.950 163.050 343.050 165.150 ;
        RECT 344.250 163.950 345.450 171.300 ;
        RECT 350.100 168.150 351.900 169.950 ;
        RECT 347.100 165.150 348.900 166.950 ;
        RECT 349.950 166.050 352.050 168.150 ;
        RECT 352.950 167.850 355.050 169.950 ;
        RECT 356.100 168.150 357.900 169.950 ;
        RECT 353.100 166.050 354.900 167.850 ;
        RECT 355.950 166.050 358.050 168.150 ;
        RECT 359.700 166.950 360.900 173.400 ;
        RECT 368.400 168.150 369.600 176.400 ;
        RECT 377.850 172.200 379.650 179.250 ;
        RECT 382.350 173.400 384.150 179.250 ;
        RECT 388.650 178.500 396.450 179.250 ;
        RECT 388.650 173.400 390.450 178.500 ;
        RECT 391.650 173.400 393.450 177.600 ;
        RECT 394.650 174.000 396.450 178.500 ;
        RECT 397.650 174.900 399.450 179.250 ;
        RECT 400.650 174.000 402.450 179.250 ;
        RECT 404.550 176.400 406.350 179.250 ;
        RECT 377.850 171.300 381.450 172.200 ;
        RECT 343.950 161.850 346.050 163.950 ;
        RECT 346.950 163.050 349.050 165.150 ;
        RECT 358.950 164.850 361.050 166.950 ;
        RECT 367.950 166.050 370.050 168.150 ;
        RECT 370.950 167.850 373.050 169.950 ;
        RECT 371.100 166.050 372.900 167.850 ;
        RECT 340.950 159.450 343.050 160.050 ;
        RECT 332.100 157.050 333.900 158.850 ;
        RECT 338.550 158.550 343.050 159.450 ;
        RECT 340.950 157.950 343.050 158.550 ;
        RECT 326.250 153.900 333.300 154.800 ;
        RECT 326.250 153.600 327.450 153.900 ;
        RECT 325.650 147.750 327.450 153.600 ;
        RECT 331.650 153.600 333.300 153.900 ;
        RECT 344.250 153.600 345.450 161.850 ;
        RECT 359.700 159.600 360.900 164.850 ;
        RECT 350.550 158.700 358.350 159.600 ;
        RECT 328.650 147.750 330.450 153.000 ;
        RECT 331.650 147.750 333.450 153.600 ;
        RECT 334.650 147.750 336.450 153.600 ;
        RECT 340.650 147.750 342.450 153.600 ;
        RECT 343.650 147.750 345.450 153.600 ;
        RECT 346.650 147.750 348.450 153.600 ;
        RECT 350.550 147.750 352.350 158.700 ;
        RECT 353.550 147.750 355.350 157.800 ;
        RECT 356.550 147.750 358.350 158.700 ;
        RECT 359.550 147.750 361.350 159.600 ;
        RECT 368.400 153.600 369.600 166.050 ;
        RECT 377.100 165.150 378.900 166.950 ;
        RECT 376.950 163.050 379.050 165.150 ;
        RECT 380.250 163.950 381.450 171.300 ;
        RECT 392.250 171.900 393.150 173.400 ;
        RECT 394.650 173.100 402.450 174.000 ;
        RECT 405.150 172.500 406.350 176.400 ;
        RECT 407.850 173.400 409.650 179.250 ;
        RECT 410.850 173.400 412.650 179.250 ;
        RECT 417.150 173.400 418.950 179.250 ;
        RECT 420.150 176.400 421.950 179.250 ;
        RECT 424.950 177.300 426.750 179.250 ;
        RECT 423.000 176.400 426.750 177.300 ;
        RECT 429.450 176.400 431.250 179.250 ;
        RECT 432.750 176.400 434.550 179.250 ;
        RECT 436.650 176.400 438.450 179.250 ;
        RECT 440.850 176.400 442.650 179.250 ;
        RECT 445.350 176.400 447.150 179.250 ;
        RECT 423.000 175.500 424.050 176.400 ;
        RECT 421.950 173.400 424.050 175.500 ;
        RECT 432.750 174.600 433.800 176.400 ;
        RECT 392.250 170.850 396.600 171.900 ;
        RECT 405.150 171.600 410.250 172.500 ;
        RECT 392.700 168.150 394.500 169.950 ;
        RECT 383.100 165.150 384.900 166.950 ;
        RECT 379.950 161.850 382.050 163.950 ;
        RECT 382.950 163.050 385.050 165.150 ;
        RECT 388.950 164.850 391.050 166.950 ;
        RECT 391.950 166.050 394.050 168.150 ;
        RECT 395.400 166.950 396.600 170.850 ;
        RECT 408.000 170.700 410.250 171.600 ;
        RECT 398.100 168.150 399.900 169.950 ;
        RECT 394.950 164.850 397.050 166.950 ;
        RECT 397.950 166.050 400.050 168.150 ;
        RECT 400.950 164.850 403.050 166.950 ;
        RECT 403.950 164.850 406.050 166.950 ;
        RECT 389.250 163.050 391.050 164.850 ;
        RECT 380.250 153.600 381.450 161.850 ;
        RECT 395.250 159.600 396.450 164.850 ;
        RECT 401.100 163.050 402.900 164.850 ;
        RECT 404.100 163.050 405.900 164.850 ;
        RECT 408.000 162.300 409.050 170.700 ;
        RECT 411.150 166.950 412.350 173.400 ;
        RECT 409.950 164.850 412.350 166.950 ;
        RECT 408.000 161.400 410.250 162.300 ;
        RECT 404.550 160.500 410.250 161.400 ;
        RECT 367.650 147.750 369.450 153.600 ;
        RECT 370.650 147.750 372.450 153.600 ;
        RECT 376.650 147.750 378.450 153.600 ;
        RECT 379.650 147.750 381.450 153.600 ;
        RECT 382.650 147.750 384.450 153.600 ;
        RECT 390.150 147.750 391.950 159.600 ;
        RECT 394.650 147.750 397.950 159.600 ;
        RECT 400.650 147.750 402.450 159.600 ;
        RECT 404.550 153.600 405.750 160.500 ;
        RECT 411.150 159.600 412.350 164.850 ;
        RECT 417.150 160.800 418.050 173.400 ;
        RECT 425.550 172.800 427.350 174.600 ;
        RECT 428.850 173.550 433.800 174.600 ;
        RECT 441.300 175.500 442.350 176.400 ;
        RECT 441.300 174.300 445.050 175.500 ;
        RECT 428.850 172.800 430.650 173.550 ;
        RECT 425.850 171.900 426.900 172.800 ;
        RECT 436.050 172.200 437.850 174.000 ;
        RECT 442.950 173.400 445.050 174.300 ;
        RECT 448.650 173.400 450.450 179.250 ;
        RECT 452.850 173.400 454.650 179.250 ;
        RECT 436.050 171.900 436.950 172.200 ;
        RECT 425.850 171.000 436.950 171.900 ;
        RECT 449.250 171.150 450.450 173.400 ;
        RECT 457.350 172.200 459.150 179.250 ;
        RECT 466.650 173.400 468.450 179.250 ;
        RECT 425.850 169.800 426.900 171.000 ;
        RECT 420.000 168.600 426.900 169.800 ;
        RECT 420.000 167.850 420.900 168.600 ;
        RECT 425.100 168.000 426.900 168.600 ;
        RECT 419.100 166.050 420.900 167.850 ;
        RECT 422.100 166.950 423.900 167.700 ;
        RECT 436.050 166.950 436.950 171.000 ;
        RECT 445.950 169.050 450.450 171.150 ;
        RECT 444.150 167.250 448.050 169.050 ;
        RECT 445.950 166.950 448.050 167.250 ;
        RECT 422.100 165.900 430.050 166.950 ;
        RECT 427.950 164.850 430.050 165.900 ;
        RECT 433.950 164.850 436.950 166.950 ;
        RECT 426.450 161.100 428.250 161.400 ;
        RECT 426.450 160.800 434.850 161.100 ;
        RECT 417.150 160.200 434.850 160.800 ;
        RECT 417.150 159.600 428.250 160.200 ;
        RECT 404.550 147.750 406.350 153.600 ;
        RECT 407.850 147.750 409.650 159.600 ;
        RECT 410.850 147.750 412.650 159.600 ;
        RECT 417.150 147.750 418.950 159.600 ;
        RECT 431.250 158.700 433.050 159.300 ;
        RECT 425.550 157.500 433.050 158.700 ;
        RECT 433.950 158.100 434.850 160.200 ;
        RECT 436.050 160.200 436.950 164.850 ;
        RECT 446.250 161.400 448.050 163.200 ;
        RECT 442.950 160.200 447.150 161.400 ;
        RECT 436.050 159.300 442.050 160.200 ;
        RECT 442.950 159.300 445.050 160.200 ;
        RECT 449.250 159.600 450.450 169.050 ;
        RECT 455.550 171.300 459.150 172.200 ;
        RECT 467.250 171.300 468.450 173.400 ;
        RECT 469.650 174.300 471.450 179.250 ;
        RECT 472.650 175.200 474.450 179.250 ;
        RECT 475.650 174.300 477.450 179.250 ;
        RECT 469.650 172.950 477.450 174.300 ;
        RECT 479.550 173.400 481.350 179.250 ;
        RECT 482.550 173.400 484.350 179.250 ;
        RECT 485.550 173.400 487.350 179.250 ;
        RECT 488.550 173.400 490.350 179.250 ;
        RECT 491.550 173.400 493.350 179.250 ;
        RECT 499.350 173.400 501.150 179.250 ;
        RECT 502.350 173.400 504.150 179.250 ;
        RECT 505.650 176.400 507.450 179.250 ;
        RECT 509.550 176.400 511.350 179.250 ;
        RECT 482.550 172.500 483.750 173.400 ;
        RECT 488.550 172.500 489.750 173.400 ;
        RECT 482.550 171.300 489.750 172.500 ;
        RECT 452.100 165.150 453.900 166.950 ;
        RECT 451.950 163.050 454.050 165.150 ;
        RECT 455.550 163.950 456.750 171.300 ;
        RECT 467.250 170.250 471.000 171.300 ;
        RECT 469.950 166.950 471.150 170.250 ;
        RECT 473.100 168.150 474.900 169.950 ;
        RECT 458.100 165.150 459.900 166.950 ;
        RECT 454.950 161.850 457.050 163.950 ;
        RECT 457.950 163.050 460.050 165.150 ;
        RECT 469.950 164.850 472.050 166.950 ;
        RECT 472.950 166.050 475.050 168.150 ;
        RECT 488.550 166.950 489.750 171.300 ;
        RECT 499.650 166.950 500.850 173.400 ;
        RECT 505.650 172.500 506.850 176.400 ;
        RECT 501.750 171.600 506.850 172.500 ;
        RECT 510.150 172.500 511.350 176.400 ;
        RECT 512.850 173.400 514.650 179.250 ;
        RECT 515.850 173.400 517.650 179.250 ;
        RECT 521.550 173.400 523.350 179.250 ;
        RECT 524.550 173.400 526.350 179.250 ;
        RECT 527.550 173.400 529.350 179.250 ;
        RECT 510.150 171.600 515.250 172.500 ;
        RECT 501.750 170.700 504.000 171.600 ;
        RECT 475.950 164.850 478.050 166.950 ;
        RECT 481.950 164.850 484.050 166.950 ;
        RECT 487.950 164.850 490.050 166.950 ;
        RECT 499.650 164.850 502.050 166.950 ;
        RECT 466.950 161.850 469.050 163.950 ;
        RECT 441.150 158.400 442.050 159.300 ;
        RECT 438.450 158.100 440.250 158.400 ;
        RECT 425.550 156.600 426.750 157.500 ;
        RECT 433.950 157.200 440.250 158.100 ;
        RECT 438.450 156.600 440.250 157.200 ;
        RECT 441.150 156.600 443.850 158.400 ;
        RECT 421.950 154.500 426.750 156.600 ;
        RECT 429.150 154.500 436.050 156.300 ;
        RECT 425.550 153.600 426.750 154.500 ;
        RECT 420.150 147.750 421.950 153.600 ;
        RECT 425.250 147.750 427.050 153.600 ;
        RECT 430.050 147.750 431.850 153.600 ;
        RECT 433.050 147.750 434.850 154.500 ;
        RECT 441.150 153.600 445.050 155.700 ;
        RECT 436.950 147.750 438.750 153.600 ;
        RECT 441.150 147.750 442.950 153.600 ;
        RECT 445.650 147.750 447.450 150.600 ;
        RECT 448.650 147.750 450.450 159.600 ;
        RECT 455.550 153.600 456.750 161.850 ;
        RECT 467.250 160.050 469.050 161.850 ;
        RECT 470.850 159.600 472.050 164.850 ;
        RECT 476.100 163.050 477.900 164.850 ;
        RECT 482.100 163.050 483.900 164.850 ;
        RECT 488.550 161.400 489.750 164.850 ;
        RECT 482.550 160.500 489.750 161.400 ;
        RECT 452.550 147.750 454.350 153.600 ;
        RECT 455.550 147.750 457.350 153.600 ;
        RECT 458.550 147.750 460.350 153.600 ;
        RECT 467.400 147.750 469.200 153.600 ;
        RECT 470.700 147.750 472.500 159.600 ;
        RECT 474.900 147.750 476.700 159.600 ;
        RECT 479.550 147.750 481.350 159.600 ;
        RECT 482.550 147.750 484.350 160.500 ;
        RECT 488.550 159.600 489.750 160.500 ;
        RECT 499.650 159.600 500.850 164.850 ;
        RECT 502.950 162.300 504.000 170.700 ;
        RECT 513.000 170.700 515.250 171.600 ;
        RECT 505.950 164.850 508.050 166.950 ;
        RECT 508.950 164.850 511.050 166.950 ;
        RECT 506.100 163.050 507.900 164.850 ;
        RECT 509.100 163.050 510.900 164.850 ;
        RECT 501.750 161.400 504.000 162.300 ;
        RECT 513.000 162.300 514.050 170.700 ;
        RECT 516.150 166.950 517.350 173.400 ;
        RECT 524.400 172.500 526.200 173.400 ;
        RECT 530.550 172.500 532.350 179.250 ;
        RECT 533.550 173.400 535.350 179.250 ;
        RECT 536.550 173.400 538.350 179.250 ;
        RECT 539.550 173.400 541.350 179.250 ;
        RECT 542.550 173.400 544.350 179.250 ;
        RECT 545.550 173.400 547.350 179.250 ;
        RECT 551.550 173.400 553.350 179.250 ;
        RECT 554.550 173.400 556.350 179.250 ;
        RECT 557.550 173.400 559.350 179.250 ;
        RECT 536.400 172.500 538.200 173.400 ;
        RECT 542.400 172.500 544.200 173.400 ;
        RECT 554.400 172.500 556.200 173.400 ;
        RECT 560.550 172.500 562.350 179.250 ;
        RECT 563.550 173.400 565.350 179.250 ;
        RECT 566.550 173.400 568.350 179.250 ;
        RECT 569.550 173.400 571.350 179.250 ;
        RECT 572.550 173.400 574.350 179.250 ;
        RECT 575.550 173.400 577.350 179.250 ;
        RECT 581.550 176.400 583.350 179.250 ;
        RECT 566.400 172.500 568.200 173.400 ;
        RECT 572.400 172.500 574.200 173.400 ;
        RECT 582.150 172.500 583.350 176.400 ;
        RECT 584.850 173.400 586.650 179.250 ;
        RECT 587.850 173.400 589.650 179.250 ;
        RECT 593.850 173.400 595.650 179.250 ;
        RECT 524.400 171.300 528.450 172.500 ;
        RECT 530.550 171.300 534.300 172.500 ;
        RECT 536.400 171.300 540.300 172.500 ;
        RECT 542.400 172.350 545.100 172.500 ;
        RECT 542.400 171.300 545.250 172.350 ;
        RECT 554.400 171.300 558.450 172.500 ;
        RECT 560.550 171.300 564.300 172.500 ;
        RECT 566.400 171.300 570.300 172.500 ;
        RECT 572.400 172.350 575.100 172.500 ;
        RECT 572.400 171.300 575.250 172.350 ;
        RECT 582.150 171.600 587.250 172.500 ;
        RECT 527.250 170.400 528.450 171.300 ;
        RECT 533.100 170.400 534.300 171.300 ;
        RECT 539.100 170.400 540.300 171.300 ;
        RECT 524.100 168.150 525.900 169.950 ;
        RECT 527.250 168.600 531.300 170.400 ;
        RECT 533.100 168.600 537.300 170.400 ;
        RECT 539.100 168.600 543.300 170.400 ;
        RECT 514.950 164.850 517.350 166.950 ;
        RECT 523.950 166.050 526.050 168.150 ;
        RECT 513.000 161.400 515.250 162.300 ;
        RECT 501.750 160.500 507.450 161.400 ;
        RECT 485.550 147.750 487.350 159.600 ;
        RECT 488.550 147.750 490.350 159.600 ;
        RECT 491.550 147.750 493.350 159.600 ;
        RECT 499.350 147.750 501.150 159.600 ;
        RECT 502.350 147.750 504.150 159.600 ;
        RECT 506.250 153.600 507.450 160.500 ;
        RECT 505.650 147.750 507.450 153.600 ;
        RECT 509.550 160.500 515.250 161.400 ;
        RECT 509.550 153.600 510.750 160.500 ;
        RECT 516.150 159.600 517.350 164.850 ;
        RECT 527.250 161.700 528.450 168.600 ;
        RECT 533.100 161.700 534.300 168.600 ;
        RECT 539.100 161.700 540.300 168.600 ;
        RECT 544.200 168.150 545.250 171.300 ;
        RECT 557.250 170.400 558.450 171.300 ;
        RECT 563.100 170.400 564.300 171.300 ;
        RECT 569.100 170.400 570.300 171.300 ;
        RECT 554.100 168.150 555.900 169.950 ;
        RECT 557.250 168.600 561.300 170.400 ;
        RECT 563.100 168.600 567.300 170.400 ;
        RECT 569.100 168.600 573.300 170.400 ;
        RECT 544.200 166.050 547.050 168.150 ;
        RECT 553.950 166.050 556.050 168.150 ;
        RECT 544.200 161.700 545.250 166.050 ;
        RECT 557.250 161.700 558.450 168.600 ;
        RECT 563.100 161.700 564.300 168.600 ;
        RECT 569.100 161.700 570.300 168.600 ;
        RECT 574.200 168.150 575.250 171.300 ;
        RECT 585.000 170.700 587.250 171.600 ;
        RECT 574.200 166.050 577.050 168.150 ;
        RECT 574.200 161.700 575.250 166.050 ;
        RECT 580.950 164.850 583.050 166.950 ;
        RECT 581.100 163.050 582.900 164.850 ;
        RECT 524.550 160.500 528.450 161.700 ;
        RECT 530.550 160.500 534.300 161.700 ;
        RECT 536.550 160.500 540.300 161.700 ;
        RECT 542.550 160.500 545.250 161.700 ;
        RECT 554.550 160.500 558.450 161.700 ;
        RECT 560.550 160.500 564.300 161.700 ;
        RECT 566.550 160.500 570.300 161.700 ;
        RECT 572.550 160.500 575.250 161.700 ;
        RECT 585.000 162.300 586.050 170.700 ;
        RECT 588.150 166.950 589.350 173.400 ;
        RECT 598.350 172.200 600.150 179.250 ;
        RECT 596.550 171.300 600.150 172.200 ;
        RECT 605.550 173.400 607.350 179.250 ;
        RECT 608.850 176.400 610.650 179.250 ;
        RECT 613.350 176.400 615.150 179.250 ;
        RECT 617.550 176.400 619.350 179.250 ;
        RECT 621.450 176.400 623.250 179.250 ;
        RECT 624.750 176.400 626.550 179.250 ;
        RECT 629.250 177.300 631.050 179.250 ;
        RECT 629.250 176.400 633.000 177.300 ;
        RECT 634.050 176.400 635.850 179.250 ;
        RECT 613.650 175.500 614.700 176.400 ;
        RECT 610.950 174.300 614.700 175.500 ;
        RECT 622.200 174.600 623.250 176.400 ;
        RECT 631.950 175.500 633.000 176.400 ;
        RECT 610.950 173.400 613.050 174.300 ;
        RECT 586.950 164.850 589.350 166.950 ;
        RECT 593.100 165.150 594.900 166.950 ;
        RECT 585.000 161.400 587.250 162.300 ;
        RECT 581.550 160.500 587.250 161.400 ;
        RECT 509.550 147.750 511.350 153.600 ;
        RECT 512.850 147.750 514.650 159.600 ;
        RECT 515.850 147.750 517.650 159.600 ;
        RECT 521.550 147.750 523.350 159.600 ;
        RECT 524.550 147.750 526.350 160.500 ;
        RECT 527.550 147.750 529.350 159.600 ;
        RECT 530.550 147.750 532.350 160.500 ;
        RECT 533.550 147.750 535.350 159.600 ;
        RECT 536.550 147.750 538.350 160.500 ;
        RECT 539.550 147.750 541.350 159.600 ;
        RECT 542.550 147.750 544.350 160.500 ;
        RECT 545.550 147.750 547.350 159.600 ;
        RECT 551.550 147.750 553.350 159.600 ;
        RECT 554.550 147.750 556.350 160.500 ;
        RECT 557.550 147.750 559.350 159.600 ;
        RECT 560.550 147.750 562.350 160.500 ;
        RECT 563.550 147.750 565.350 159.600 ;
        RECT 566.550 147.750 568.350 160.500 ;
        RECT 569.550 147.750 571.350 159.600 ;
        RECT 572.550 147.750 574.350 160.500 ;
        RECT 575.550 147.750 577.350 159.600 ;
        RECT 581.550 153.600 582.750 160.500 ;
        RECT 588.150 159.600 589.350 164.850 ;
        RECT 592.950 163.050 595.050 165.150 ;
        RECT 596.550 163.950 597.750 171.300 ;
        RECT 605.550 171.150 606.750 173.400 ;
        RECT 618.150 172.200 619.950 174.000 ;
        RECT 622.200 173.550 627.150 174.600 ;
        RECT 625.350 172.800 627.150 173.550 ;
        RECT 628.650 172.800 630.450 174.600 ;
        RECT 631.950 173.400 634.050 175.500 ;
        RECT 637.050 173.400 638.850 179.250 ;
        RECT 641.850 173.400 643.650 179.250 ;
        RECT 619.050 171.900 619.950 172.200 ;
        RECT 629.100 171.900 630.150 172.800 ;
        RECT 605.550 169.050 610.050 171.150 ;
        RECT 619.050 171.000 630.150 171.900 ;
        RECT 599.100 165.150 600.900 166.950 ;
        RECT 595.950 161.850 598.050 163.950 ;
        RECT 598.950 163.050 601.050 165.150 ;
        RECT 581.550 147.750 583.350 153.600 ;
        RECT 584.850 147.750 586.650 159.600 ;
        RECT 587.850 147.750 589.650 159.600 ;
        RECT 596.550 153.600 597.750 161.850 ;
        RECT 605.550 159.600 606.750 169.050 ;
        RECT 607.950 167.250 611.850 169.050 ;
        RECT 607.950 166.950 610.050 167.250 ;
        RECT 619.050 166.950 619.950 171.000 ;
        RECT 629.100 169.800 630.150 171.000 ;
        RECT 629.100 168.600 636.000 169.800 ;
        RECT 629.100 168.000 630.900 168.600 ;
        RECT 635.100 167.850 636.000 168.600 ;
        RECT 632.100 166.950 633.900 167.700 ;
        RECT 619.050 164.850 622.050 166.950 ;
        RECT 625.950 165.900 633.900 166.950 ;
        RECT 635.100 166.050 636.900 167.850 ;
        RECT 625.950 164.850 628.050 165.900 ;
        RECT 607.950 161.400 609.750 163.200 ;
        RECT 608.850 160.200 613.050 161.400 ;
        RECT 619.050 160.200 619.950 164.850 ;
        RECT 627.750 161.100 629.550 161.400 ;
        RECT 593.550 147.750 595.350 153.600 ;
        RECT 596.550 147.750 598.350 153.600 ;
        RECT 599.550 147.750 601.350 153.600 ;
        RECT 605.550 147.750 607.350 159.600 ;
        RECT 610.950 159.300 613.050 160.200 ;
        RECT 613.950 159.300 619.950 160.200 ;
        RECT 621.150 160.800 629.550 161.100 ;
        RECT 637.950 160.800 638.850 173.400 ;
        RECT 646.350 172.200 648.150 179.250 ;
        RECT 653.550 174.300 655.350 179.250 ;
        RECT 656.550 175.200 658.350 179.250 ;
        RECT 659.550 174.300 661.350 179.250 ;
        RECT 653.550 172.950 661.350 174.300 ;
        RECT 662.550 173.400 664.350 179.250 ;
        RECT 644.550 171.300 648.150 172.200 ;
        RECT 662.550 171.300 663.750 173.400 ;
        RECT 671.850 172.200 673.650 179.250 ;
        RECT 676.350 173.400 678.150 179.250 ;
        RECT 680.550 174.300 682.350 179.250 ;
        RECT 683.550 175.200 685.350 179.250 ;
        RECT 686.550 174.300 688.350 179.250 ;
        RECT 680.550 172.950 688.350 174.300 ;
        RECT 689.550 173.400 691.350 179.250 ;
        RECT 671.850 171.300 675.450 172.200 ;
        RECT 689.550 171.300 690.750 173.400 ;
        RECT 641.100 165.150 642.900 166.950 ;
        RECT 640.950 163.050 643.050 165.150 ;
        RECT 644.550 163.950 645.750 171.300 ;
        RECT 660.000 170.250 663.750 171.300 ;
        RECT 656.100 168.150 657.900 169.950 ;
        RECT 647.100 165.150 648.900 166.950 ;
        RECT 643.950 161.850 646.050 163.950 ;
        RECT 646.950 163.050 649.050 165.150 ;
        RECT 652.950 164.850 655.050 166.950 ;
        RECT 655.950 166.050 658.050 168.150 ;
        RECT 659.850 166.950 661.050 170.250 ;
        RECT 658.950 164.850 661.050 166.950 ;
        RECT 671.100 165.150 672.900 166.950 ;
        RECT 653.100 163.050 654.900 164.850 ;
        RECT 621.150 160.200 638.850 160.800 ;
        RECT 613.950 158.400 614.850 159.300 ;
        RECT 612.150 156.600 614.850 158.400 ;
        RECT 615.750 158.100 617.550 158.400 ;
        RECT 621.150 158.100 622.050 160.200 ;
        RECT 627.750 159.600 638.850 160.200 ;
        RECT 615.750 157.200 622.050 158.100 ;
        RECT 622.950 158.700 624.750 159.300 ;
        RECT 622.950 157.500 630.450 158.700 ;
        RECT 615.750 156.600 617.550 157.200 ;
        RECT 629.250 156.600 630.450 157.500 ;
        RECT 610.950 153.600 614.850 155.700 ;
        RECT 619.950 154.500 626.850 156.300 ;
        RECT 629.250 154.500 634.050 156.600 ;
        RECT 608.550 147.750 610.350 150.600 ;
        RECT 613.050 147.750 614.850 153.600 ;
        RECT 617.250 147.750 619.050 153.600 ;
        RECT 621.150 147.750 622.950 154.500 ;
        RECT 629.250 153.600 630.450 154.500 ;
        RECT 624.150 147.750 625.950 153.600 ;
        RECT 628.950 147.750 630.750 153.600 ;
        RECT 634.050 147.750 635.850 153.600 ;
        RECT 637.050 147.750 638.850 159.600 ;
        RECT 644.550 153.600 645.750 161.850 ;
        RECT 658.950 159.600 660.150 164.850 ;
        RECT 661.950 161.850 664.050 163.950 ;
        RECT 670.950 163.050 673.050 165.150 ;
        RECT 674.250 163.950 675.450 171.300 ;
        RECT 687.000 170.250 690.750 171.300 ;
        RECT 695.700 170.400 697.500 179.250 ;
        RECT 701.100 171.000 702.900 179.250 ;
        RECT 683.100 168.150 684.900 169.950 ;
        RECT 677.100 165.150 678.900 166.950 ;
        RECT 673.950 161.850 676.050 163.950 ;
        RECT 676.950 163.050 679.050 165.150 ;
        RECT 679.950 164.850 682.050 166.950 ;
        RECT 682.950 166.050 685.050 168.150 ;
        RECT 686.850 166.950 688.050 170.250 ;
        RECT 701.100 169.350 705.600 171.000 ;
        RECT 685.950 164.850 688.050 166.950 ;
        RECT 704.400 165.150 705.600 169.350 ;
        RECT 680.100 163.050 681.900 164.850 ;
        RECT 661.950 160.050 663.750 161.850 ;
        RECT 641.550 147.750 643.350 153.600 ;
        RECT 644.550 147.750 646.350 153.600 ;
        RECT 647.550 147.750 649.350 153.600 ;
        RECT 654.300 147.750 656.100 159.600 ;
        RECT 658.500 147.750 660.300 159.600 ;
        RECT 674.250 153.600 675.450 161.850 ;
        RECT 685.950 159.600 687.150 164.850 ;
        RECT 688.950 161.850 691.050 163.950 ;
        RECT 694.950 161.850 697.050 163.950 ;
        RECT 700.950 161.850 703.050 163.950 ;
        RECT 703.950 163.050 706.050 165.150 ;
        RECT 688.950 160.050 690.750 161.850 ;
        RECT 695.100 160.050 696.900 161.850 ;
        RECT 661.800 147.750 663.600 153.600 ;
        RECT 670.650 147.750 672.450 153.600 ;
        RECT 673.650 147.750 675.450 153.600 ;
        RECT 676.650 147.750 678.450 153.600 ;
        RECT 681.300 147.750 683.100 159.600 ;
        RECT 685.500 147.750 687.300 159.600 ;
        RECT 697.950 158.850 700.050 160.950 ;
        RECT 701.250 160.050 703.050 161.850 ;
        RECT 698.100 157.050 699.900 158.850 ;
        RECT 704.700 154.800 705.750 163.050 ;
        RECT 698.700 153.900 705.750 154.800 ;
        RECT 698.700 153.600 700.350 153.900 ;
        RECT 688.800 147.750 690.600 153.600 ;
        RECT 695.550 147.750 697.350 153.600 ;
        RECT 698.550 147.750 700.350 153.600 ;
        RECT 704.550 153.600 705.750 153.900 ;
        RECT 701.550 147.750 703.350 153.000 ;
        RECT 704.550 147.750 706.350 153.600 ;
        RECT 4.650 137.400 6.450 143.250 ;
        RECT 7.650 137.400 9.450 143.250 ;
        RECT 10.650 137.400 12.450 143.250 ;
        RECT 8.250 129.150 9.450 137.400 ;
        RECT 16.050 131.400 17.850 143.250 ;
        RECT 19.050 131.400 20.850 143.250 ;
        RECT 22.650 137.400 24.450 143.250 ;
        RECT 25.650 137.400 27.450 143.250 ;
        RECT 32.400 137.400 34.200 143.250 ;
        RECT 4.950 125.850 7.050 127.950 ;
        RECT 7.950 127.050 10.050 129.150 ;
        RECT 5.100 124.050 6.900 125.850 ;
        RECT 8.250 119.700 9.450 127.050 ;
        RECT 10.950 125.850 13.050 127.950 ;
        RECT 16.650 126.150 17.850 131.400 ;
        RECT 11.100 124.050 12.900 125.850 ;
        RECT 16.650 124.050 19.050 126.150 ;
        RECT 19.950 125.850 22.050 127.950 ;
        RECT 20.100 124.050 21.900 125.850 ;
        RECT 5.850 118.800 9.450 119.700 ;
        RECT 5.850 111.750 7.650 118.800 ;
        RECT 16.650 117.600 17.850 124.050 ;
        RECT 23.100 120.300 24.300 137.400 ;
        RECT 35.700 131.400 37.500 143.250 ;
        RECT 39.900 131.400 41.700 143.250 ;
        RECT 46.650 142.500 54.450 143.250 ;
        RECT 46.650 131.400 48.450 142.500 ;
        RECT 49.650 131.400 51.450 141.600 ;
        RECT 52.650 132.600 54.450 142.500 ;
        RECT 55.650 133.500 57.450 143.250 ;
        RECT 58.650 132.600 60.450 143.250 ;
        RECT 52.650 131.700 60.450 132.600 ;
        RECT 64.350 131.400 66.150 143.250 ;
        RECT 67.350 131.400 69.150 143.250 ;
        RECT 70.650 137.400 72.450 143.250 ;
        RECT 74.550 137.400 76.350 143.250 ;
        RECT 77.550 137.400 79.350 143.250 ;
        RECT 85.650 137.400 87.450 143.250 ;
        RECT 88.650 137.400 90.450 143.250 ;
        RECT 32.250 129.150 34.050 130.950 ;
        RECT 26.100 126.150 27.900 127.950 ;
        RECT 31.950 127.050 34.050 129.150 ;
        RECT 35.850 126.150 37.050 131.400 ;
        RECT 49.800 130.500 51.600 131.400 ;
        RECT 49.800 129.600 53.850 130.500 ;
        RECT 41.100 126.150 42.900 127.950 ;
        RECT 47.100 126.150 48.900 127.950 ;
        RECT 52.950 126.150 53.850 129.600 ;
        RECT 58.950 126.150 60.750 127.950 ;
        RECT 64.650 126.150 65.850 131.400 ;
        RECT 71.250 130.500 72.450 137.400 ;
        RECT 66.750 129.600 72.450 130.500 ;
        RECT 66.750 128.700 69.000 129.600 ;
        RECT 25.950 124.050 28.050 126.150 ;
        RECT 34.950 124.050 37.050 126.150 ;
        RECT 34.950 120.750 36.150 124.050 ;
        RECT 37.950 122.850 40.050 124.950 ;
        RECT 40.950 124.050 43.050 126.150 ;
        RECT 46.950 124.050 49.050 126.150 ;
        RECT 49.950 122.850 52.050 124.950 ;
        RECT 52.950 124.050 55.050 126.150 ;
        RECT 38.100 121.050 39.900 122.850 ;
        RECT 50.250 121.050 52.050 122.850 ;
        RECT 19.950 119.100 27.450 120.300 ;
        RECT 19.950 118.500 21.750 119.100 ;
        RECT 10.350 111.750 12.150 117.600 ;
        RECT 16.650 116.100 19.950 117.600 ;
        RECT 18.150 111.750 19.950 116.100 ;
        RECT 21.150 111.750 22.950 117.600 ;
        RECT 25.650 111.750 27.450 119.100 ;
        RECT 32.250 119.700 36.000 120.750 ;
        RECT 32.250 117.600 33.450 119.700 ;
        RECT 31.650 111.750 33.450 117.600 ;
        RECT 34.650 116.700 42.450 118.050 ;
        RECT 54.000 117.600 55.050 124.050 ;
        RECT 55.950 122.850 58.050 124.950 ;
        RECT 58.950 124.050 61.050 126.150 ;
        RECT 64.650 124.050 67.050 126.150 ;
        RECT 55.950 121.050 57.750 122.850 ;
        RECT 64.650 117.600 65.850 124.050 ;
        RECT 67.950 120.300 69.000 128.700 ;
        RECT 71.100 126.150 72.900 127.950 ;
        RECT 70.950 124.050 73.050 126.150 ;
        RECT 77.400 124.950 78.600 137.400 ;
        RECT 86.400 124.950 87.600 137.400 ;
        RECT 94.650 131.400 96.450 143.250 ;
        RECT 97.650 132.300 99.450 143.250 ;
        RECT 100.650 133.200 102.450 143.250 ;
        RECT 103.650 132.300 105.450 143.250 ;
        RECT 107.550 137.400 109.350 143.250 ;
        RECT 110.550 137.400 112.350 143.250 ;
        RECT 113.550 138.000 115.350 143.250 ;
        RECT 110.700 137.100 112.350 137.400 ;
        RECT 116.550 137.400 118.350 143.250 ;
        RECT 116.550 137.100 117.750 137.400 ;
        RECT 110.700 136.200 117.750 137.100 ;
        RECT 97.650 131.400 105.450 132.300 ;
        RECT 110.100 132.150 111.900 133.950 ;
        RECT 95.100 126.150 96.300 131.400 ;
        RECT 107.100 129.150 108.900 130.950 ;
        RECT 109.950 130.050 112.050 132.150 ;
        RECT 113.250 129.150 115.050 130.950 ;
        RECT 106.950 127.050 109.050 129.150 ;
        RECT 112.950 127.050 115.050 129.150 ;
        RECT 116.700 127.950 117.750 136.200 ;
        RECT 124.050 131.400 125.850 143.250 ;
        RECT 127.050 131.400 128.850 143.250 ;
        RECT 130.650 137.400 132.450 143.250 ;
        RECT 133.650 137.400 135.450 143.250 ;
        RECT 137.550 137.400 139.350 143.250 ;
        RECT 140.550 137.400 142.350 143.250 ;
        RECT 143.550 137.400 145.350 143.250 ;
        RECT 151.650 137.400 153.450 143.250 ;
        RECT 154.650 138.000 156.450 143.250 ;
        RECT 74.100 123.150 75.900 124.950 ;
        RECT 73.950 121.050 76.050 123.150 ;
        RECT 76.950 122.850 79.050 124.950 ;
        RECT 85.950 122.850 88.050 124.950 ;
        RECT 89.100 123.150 90.900 124.950 ;
        RECT 94.950 124.050 97.050 126.150 ;
        RECT 115.950 125.850 118.050 127.950 ;
        RECT 124.650 126.150 125.850 131.400 ;
        RECT 66.750 119.400 69.000 120.300 ;
        RECT 66.750 118.500 71.850 119.400 ;
        RECT 34.650 111.750 36.450 116.700 ;
        RECT 37.650 111.750 39.450 115.800 ;
        RECT 40.650 111.750 42.450 116.700 ;
        RECT 49.800 111.750 51.600 117.600 ;
        RECT 54.000 111.750 55.800 117.600 ;
        RECT 58.200 111.750 60.000 117.600 ;
        RECT 64.350 111.750 66.150 117.600 ;
        RECT 67.350 111.750 69.150 117.600 ;
        RECT 70.650 114.600 71.850 118.500 ;
        RECT 77.400 114.600 78.600 122.850 ;
        RECT 86.400 114.600 87.600 122.850 ;
        RECT 88.950 121.050 91.050 123.150 ;
        RECT 95.100 117.600 96.300 124.050 ;
        RECT 97.950 122.850 100.050 124.950 ;
        RECT 101.100 123.150 102.900 124.950 ;
        RECT 98.100 121.050 99.900 122.850 ;
        RECT 100.950 121.050 103.050 123.150 ;
        RECT 103.950 122.850 106.050 124.950 ;
        RECT 104.100 121.050 105.900 122.850 ;
        RECT 116.400 121.650 117.600 125.850 ;
        RECT 95.100 115.950 100.800 117.600 ;
        RECT 70.650 111.750 72.450 114.600 ;
        RECT 74.550 111.750 76.350 114.600 ;
        RECT 77.550 111.750 79.350 114.600 ;
        RECT 85.650 111.750 87.450 114.600 ;
        RECT 88.650 111.750 90.450 114.600 ;
        RECT 95.700 111.750 97.500 114.600 ;
        RECT 99.000 111.750 100.800 115.950 ;
        RECT 103.200 111.750 105.000 117.600 ;
        RECT 107.700 111.750 109.500 120.600 ;
        RECT 113.100 120.000 117.600 121.650 ;
        RECT 124.650 124.050 127.050 126.150 ;
        RECT 127.950 125.850 130.050 127.950 ;
        RECT 128.100 124.050 129.900 125.850 ;
        RECT 113.100 111.750 114.900 120.000 ;
        RECT 124.650 117.600 125.850 124.050 ;
        RECT 131.100 120.300 132.300 137.400 ;
        RECT 140.550 129.150 141.750 137.400 ;
        RECT 152.250 137.100 153.450 137.400 ;
        RECT 157.650 137.400 159.450 143.250 ;
        RECT 160.650 137.400 162.450 143.250 ;
        RECT 157.650 137.100 159.300 137.400 ;
        RECT 152.250 136.200 159.300 137.100 ;
        RECT 134.100 126.150 135.900 127.950 ;
        RECT 133.950 124.050 136.050 126.150 ;
        RECT 136.950 125.850 139.050 127.950 ;
        RECT 139.950 127.050 142.050 129.150 ;
        RECT 152.250 127.950 153.300 136.200 ;
        RECT 158.100 132.150 159.900 133.950 ;
        RECT 154.950 129.150 156.750 130.950 ;
        RECT 157.950 130.050 160.050 132.150 ;
        RECT 165.300 131.400 167.100 143.250 ;
        RECT 169.500 131.400 171.300 143.250 ;
        RECT 172.800 137.400 174.600 143.250 ;
        RECT 181.650 137.400 183.450 143.250 ;
        RECT 184.650 138.000 186.450 143.250 ;
        RECT 182.250 137.100 183.450 137.400 ;
        RECT 187.650 137.400 189.450 143.250 ;
        RECT 190.650 137.400 192.450 143.250 ;
        RECT 194.550 137.400 196.350 143.250 ;
        RECT 197.550 137.400 199.350 143.250 ;
        RECT 187.650 137.100 189.300 137.400 ;
        RECT 182.250 136.200 189.300 137.100 ;
        RECT 161.100 129.150 162.900 130.950 ;
        RECT 137.100 124.050 138.900 125.850 ;
        RECT 127.950 119.100 135.450 120.300 ;
        RECT 127.950 118.500 129.750 119.100 ;
        RECT 124.650 116.100 127.950 117.600 ;
        RECT 126.150 111.750 127.950 116.100 ;
        RECT 129.150 111.750 130.950 117.600 ;
        RECT 133.650 111.750 135.450 119.100 ;
        RECT 140.550 119.700 141.750 127.050 ;
        RECT 142.950 125.850 145.050 127.950 ;
        RECT 151.950 125.850 154.050 127.950 ;
        RECT 154.950 127.050 157.050 129.150 ;
        RECT 160.950 127.050 163.050 129.150 ;
        RECT 164.100 126.150 165.900 127.950 ;
        RECT 169.950 126.150 171.150 131.400 ;
        RECT 172.950 129.150 174.750 130.950 ;
        RECT 172.950 127.050 175.050 129.150 ;
        RECT 182.250 127.950 183.300 136.200 ;
        RECT 188.100 132.150 189.900 133.950 ;
        RECT 184.950 129.150 186.750 130.950 ;
        RECT 187.950 130.050 190.050 132.150 ;
        RECT 191.100 129.150 192.900 130.950 ;
        RECT 143.100 124.050 144.900 125.850 ;
        RECT 152.400 121.650 153.600 125.850 ;
        RECT 163.950 124.050 166.050 126.150 ;
        RECT 166.950 122.850 169.050 124.950 ;
        RECT 169.950 124.050 172.050 126.150 ;
        RECT 181.950 125.850 184.050 127.950 ;
        RECT 184.950 127.050 187.050 129.150 ;
        RECT 190.950 127.050 193.050 129.150 ;
        RECT 152.400 120.000 156.900 121.650 ;
        RECT 167.100 121.050 168.900 122.850 ;
        RECT 170.850 120.750 172.050 124.050 ;
        RECT 182.400 121.650 183.600 125.850 ;
        RECT 197.400 124.950 198.600 137.400 ;
        RECT 204.300 131.400 206.100 143.250 ;
        RECT 208.500 131.400 210.300 143.250 ;
        RECT 211.800 137.400 213.600 143.250 ;
        RECT 220.650 137.400 222.450 143.250 ;
        RECT 223.650 137.400 225.450 143.250 ;
        RECT 226.650 137.400 228.450 143.250 ;
        RECT 230.550 137.400 232.350 143.250 ;
        RECT 233.550 137.400 235.350 143.250 ;
        RECT 236.550 137.400 238.350 143.250 ;
        RECT 241.950 139.950 244.050 142.050 ;
        RECT 203.100 126.150 204.900 127.950 ;
        RECT 208.950 126.150 210.150 131.400 ;
        RECT 211.950 129.150 213.750 130.950 ;
        RECT 224.250 129.150 225.450 137.400 ;
        RECT 233.550 129.150 234.750 137.400 ;
        RECT 235.950 132.450 238.050 133.050 ;
        RECT 235.950 131.550 240.450 132.450 ;
        RECT 235.950 130.950 238.050 131.550 ;
        RECT 239.550 130.050 240.450 131.550 ;
        RECT 211.950 127.050 214.050 129.150 ;
        RECT 194.100 123.150 195.900 124.950 ;
        RECT 140.550 118.800 144.150 119.700 ;
        RECT 137.850 111.750 139.650 117.600 ;
        RECT 142.350 111.750 144.150 118.800 ;
        RECT 155.100 111.750 156.900 120.000 ;
        RECT 160.500 111.750 162.300 120.600 ;
        RECT 171.000 119.700 174.750 120.750 ;
        RECT 182.400 120.000 186.900 121.650 ;
        RECT 193.950 121.050 196.050 123.150 ;
        RECT 196.950 122.850 199.050 124.950 ;
        RECT 202.950 124.050 205.050 126.150 ;
        RECT 205.950 122.850 208.050 124.950 ;
        RECT 208.950 124.050 211.050 126.150 ;
        RECT 220.950 125.850 223.050 127.950 ;
        RECT 223.950 127.050 226.050 129.150 ;
        RECT 221.100 124.050 222.900 125.850 ;
        RECT 164.550 116.700 172.350 118.050 ;
        RECT 164.550 111.750 166.350 116.700 ;
        RECT 167.550 111.750 169.350 115.800 ;
        RECT 170.550 111.750 172.350 116.700 ;
        RECT 173.550 117.600 174.750 119.700 ;
        RECT 173.550 111.750 175.350 117.600 ;
        RECT 185.100 111.750 186.900 120.000 ;
        RECT 190.500 111.750 192.300 120.600 ;
        RECT 197.400 114.600 198.600 122.850 ;
        RECT 206.100 121.050 207.900 122.850 ;
        RECT 209.850 120.750 211.050 124.050 ;
        RECT 210.000 119.700 213.750 120.750 ;
        RECT 224.250 119.700 225.450 127.050 ;
        RECT 226.950 125.850 229.050 127.950 ;
        RECT 229.950 125.850 232.050 127.950 ;
        RECT 232.950 127.050 235.050 129.150 ;
        RECT 238.950 127.950 241.050 130.050 ;
        RECT 227.100 124.050 228.900 125.850 ;
        RECT 230.100 124.050 231.900 125.850 ;
        RECT 203.550 116.700 211.350 118.050 ;
        RECT 194.550 111.750 196.350 114.600 ;
        RECT 197.550 111.750 199.350 114.600 ;
        RECT 203.550 111.750 205.350 116.700 ;
        RECT 206.550 111.750 208.350 115.800 ;
        RECT 209.550 111.750 211.350 116.700 ;
        RECT 212.550 117.600 213.750 119.700 ;
        RECT 221.850 118.800 225.450 119.700 ;
        RECT 233.550 119.700 234.750 127.050 ;
        RECT 235.950 125.850 238.050 127.950 ;
        RECT 236.100 124.050 237.900 125.850 ;
        RECT 242.550 123.450 243.450 139.950 ;
        RECT 245.400 137.400 247.200 143.250 ;
        RECT 248.700 131.400 250.500 143.250 ;
        RECT 252.900 131.400 254.700 143.250 ;
        RECT 257.550 137.400 259.350 143.250 ;
        RECT 260.550 137.400 262.350 143.250 ;
        RECT 245.250 129.150 247.050 130.950 ;
        RECT 244.950 127.050 247.050 129.150 ;
        RECT 248.850 126.150 250.050 131.400 ;
        RECT 254.100 126.150 255.900 127.950 ;
        RECT 257.100 126.150 258.900 127.950 ;
        RECT 247.950 124.050 250.050 126.150 ;
        RECT 244.950 123.450 247.050 124.050 ;
        RECT 242.550 122.550 247.050 123.450 ;
        RECT 244.950 121.950 247.050 122.550 ;
        RECT 247.950 120.750 249.150 124.050 ;
        RECT 250.950 122.850 253.050 124.950 ;
        RECT 253.950 124.050 256.050 126.150 ;
        RECT 256.950 124.050 259.050 126.150 ;
        RECT 251.100 121.050 252.900 122.850 ;
        RECT 245.250 119.700 249.000 120.750 ;
        RECT 260.700 120.300 261.900 137.400 ;
        RECT 264.150 131.400 265.950 143.250 ;
        RECT 267.150 131.400 268.950 143.250 ;
        RECT 274.650 137.400 276.450 143.250 ;
        RECT 277.650 137.400 279.450 143.250 ;
        RECT 283.650 137.400 285.450 143.250 ;
        RECT 286.650 137.400 288.450 143.250 ;
        RECT 289.650 137.400 291.450 143.250 ;
        RECT 293.550 137.400 295.350 143.250 ;
        RECT 296.550 137.400 298.350 143.250 ;
        RECT 304.650 137.400 306.450 143.250 ;
        RECT 307.650 138.000 309.450 143.250 ;
        RECT 262.950 125.850 265.050 127.950 ;
        RECT 267.150 126.150 268.350 131.400 ;
        RECT 263.100 124.050 264.900 125.850 ;
        RECT 265.950 124.050 268.350 126.150 ;
        RECT 275.400 124.950 276.600 137.400 ;
        RECT 287.250 129.150 288.450 137.400 ;
        RECT 283.950 125.850 286.050 127.950 ;
        RECT 286.950 127.050 289.050 129.150 ;
        RECT 233.550 118.800 237.150 119.700 ;
        RECT 212.550 111.750 214.350 117.600 ;
        RECT 221.850 111.750 223.650 118.800 ;
        RECT 226.350 111.750 228.150 117.600 ;
        RECT 230.850 111.750 232.650 117.600 ;
        RECT 235.350 111.750 237.150 118.800 ;
        RECT 245.250 117.600 246.450 119.700 ;
        RECT 257.550 119.100 265.050 120.300 ;
        RECT 244.650 111.750 246.450 117.600 ;
        RECT 247.650 116.700 255.450 118.050 ;
        RECT 247.650 111.750 249.450 116.700 ;
        RECT 250.650 111.750 252.450 115.800 ;
        RECT 253.650 111.750 255.450 116.700 ;
        RECT 257.550 111.750 259.350 119.100 ;
        RECT 263.250 118.500 265.050 119.100 ;
        RECT 267.150 117.600 268.350 124.050 ;
        RECT 274.950 122.850 277.050 124.950 ;
        RECT 278.100 123.150 279.900 124.950 ;
        RECT 284.100 124.050 285.900 125.850 ;
        RECT 262.050 111.750 263.850 117.600 ;
        RECT 265.050 116.100 268.350 117.600 ;
        RECT 265.050 111.750 266.850 116.100 ;
        RECT 275.400 114.600 276.600 122.850 ;
        RECT 277.950 121.050 280.050 123.150 ;
        RECT 287.250 119.700 288.450 127.050 ;
        RECT 289.950 125.850 292.050 127.950 ;
        RECT 290.100 124.050 291.900 125.850 ;
        RECT 296.400 124.950 297.600 137.400 ;
        RECT 305.250 137.100 306.450 137.400 ;
        RECT 310.650 137.400 312.450 143.250 ;
        RECT 313.650 137.400 315.450 143.250 ;
        RECT 317.550 137.400 319.350 143.250 ;
        RECT 320.550 137.400 322.350 143.250 ;
        RECT 310.650 137.100 312.300 137.400 ;
        RECT 305.250 136.200 312.300 137.100 ;
        RECT 305.250 127.950 306.300 136.200 ;
        RECT 311.100 132.150 312.900 133.950 ;
        RECT 307.950 129.150 309.750 130.950 ;
        RECT 310.950 130.050 313.050 132.150 ;
        RECT 314.100 129.150 315.900 130.950 ;
        RECT 304.950 125.850 307.050 127.950 ;
        RECT 307.950 127.050 310.050 129.150 ;
        RECT 313.950 127.050 316.050 129.150 ;
        RECT 293.100 123.150 294.900 124.950 ;
        RECT 292.950 121.050 295.050 123.150 ;
        RECT 295.950 122.850 298.050 124.950 ;
        RECT 284.850 118.800 288.450 119.700 ;
        RECT 274.650 111.750 276.450 114.600 ;
        RECT 277.650 111.750 279.450 114.600 ;
        RECT 284.850 111.750 286.650 118.800 ;
        RECT 289.350 111.750 291.150 117.600 ;
        RECT 296.400 114.600 297.600 122.850 ;
        RECT 305.400 121.650 306.600 125.850 ;
        RECT 320.400 124.950 321.600 137.400 ;
        RECT 327.300 131.400 329.100 143.250 ;
        RECT 331.500 131.400 333.300 143.250 ;
        RECT 334.800 137.400 336.600 143.250 ;
        RECT 343.650 131.400 345.450 143.250 ;
        RECT 346.650 132.300 348.450 143.250 ;
        RECT 349.650 133.200 351.450 143.250 ;
        RECT 352.650 132.300 354.450 143.250 ;
        RECT 356.550 137.400 358.350 143.250 ;
        RECT 359.550 137.400 361.350 143.250 ;
        RECT 365.550 137.400 367.350 143.250 ;
        RECT 368.550 137.400 370.350 143.250 ;
        RECT 371.550 138.000 373.350 143.250 ;
        RECT 346.650 131.400 354.450 132.300 ;
        RECT 326.100 126.150 327.900 127.950 ;
        RECT 331.950 126.150 333.150 131.400 ;
        RECT 334.950 129.150 336.750 130.950 ;
        RECT 334.950 127.050 337.050 129.150 ;
        RECT 344.100 126.150 345.300 131.400 ;
        RECT 317.100 123.150 318.900 124.950 ;
        RECT 305.400 120.000 309.900 121.650 ;
        RECT 316.950 121.050 319.050 123.150 ;
        RECT 319.950 122.850 322.050 124.950 ;
        RECT 325.950 124.050 328.050 126.150 ;
        RECT 328.950 122.850 331.050 124.950 ;
        RECT 331.950 124.050 334.050 126.150 ;
        RECT 343.950 124.050 346.050 126.150 ;
        RECT 359.400 124.950 360.600 137.400 ;
        RECT 368.700 137.100 370.350 137.400 ;
        RECT 374.550 137.400 376.350 143.250 ;
        RECT 382.650 137.400 384.450 143.250 ;
        RECT 385.650 138.000 387.450 143.250 ;
        RECT 374.550 137.100 375.750 137.400 ;
        RECT 368.700 136.200 375.750 137.100 ;
        RECT 368.100 132.150 369.900 133.950 ;
        RECT 365.100 129.150 366.900 130.950 ;
        RECT 367.950 130.050 370.050 132.150 ;
        RECT 371.250 129.150 373.050 130.950 ;
        RECT 364.950 127.050 367.050 129.150 ;
        RECT 370.950 127.050 373.050 129.150 ;
        RECT 374.700 127.950 375.750 136.200 ;
        RECT 383.250 137.100 384.450 137.400 ;
        RECT 388.650 137.400 390.450 143.250 ;
        RECT 391.650 137.400 393.450 143.250 ;
        RECT 388.650 137.100 390.300 137.400 ;
        RECT 383.250 136.200 390.300 137.100 ;
        RECT 383.250 127.950 384.300 136.200 ;
        RECT 389.100 132.150 390.900 133.950 ;
        RECT 395.550 132.300 397.350 143.250 ;
        RECT 398.550 133.200 400.350 143.250 ;
        RECT 401.550 132.300 403.350 143.250 ;
        RECT 385.950 129.150 387.750 130.950 ;
        RECT 388.950 130.050 391.050 132.150 ;
        RECT 395.550 131.400 403.350 132.300 ;
        RECT 404.550 131.400 406.350 143.250 ;
        RECT 412.650 137.400 414.450 143.250 ;
        RECT 415.650 137.400 417.450 143.250 ;
        RECT 418.650 137.400 420.450 143.250 ;
        RECT 392.100 129.150 393.900 130.950 ;
        RECT 373.950 125.850 376.050 127.950 ;
        RECT 382.950 125.850 385.050 127.950 ;
        RECT 385.950 127.050 388.050 129.150 ;
        RECT 391.950 127.050 394.050 129.150 ;
        RECT 404.700 126.150 405.900 131.400 ;
        RECT 416.250 129.150 417.450 137.400 ;
        RECT 426.150 131.400 427.950 143.250 ;
        RECT 430.650 131.400 433.950 143.250 ;
        RECT 436.650 131.400 438.450 143.250 ;
        RECT 442.650 137.400 444.450 143.250 ;
        RECT 445.650 137.400 447.450 143.250 ;
        RECT 293.550 111.750 295.350 114.600 ;
        RECT 296.550 111.750 298.350 114.600 ;
        RECT 308.100 111.750 309.900 120.000 ;
        RECT 313.500 111.750 315.300 120.600 ;
        RECT 320.400 114.600 321.600 122.850 ;
        RECT 329.100 121.050 330.900 122.850 ;
        RECT 332.850 120.750 334.050 124.050 ;
        RECT 333.000 119.700 336.750 120.750 ;
        RECT 326.550 116.700 334.350 118.050 ;
        RECT 317.550 111.750 319.350 114.600 ;
        RECT 320.550 111.750 322.350 114.600 ;
        RECT 326.550 111.750 328.350 116.700 ;
        RECT 329.550 111.750 331.350 115.800 ;
        RECT 332.550 111.750 334.350 116.700 ;
        RECT 335.550 117.600 336.750 119.700 ;
        RECT 344.100 117.600 345.300 124.050 ;
        RECT 346.950 122.850 349.050 124.950 ;
        RECT 350.100 123.150 351.900 124.950 ;
        RECT 347.100 121.050 348.900 122.850 ;
        RECT 349.950 121.050 352.050 123.150 ;
        RECT 352.950 122.850 355.050 124.950 ;
        RECT 356.100 123.150 357.900 124.950 ;
        RECT 353.100 121.050 354.900 122.850 ;
        RECT 355.950 121.050 358.050 123.150 ;
        RECT 358.950 122.850 361.050 124.950 ;
        RECT 335.550 111.750 337.350 117.600 ;
        RECT 344.100 115.950 349.800 117.600 ;
        RECT 344.700 111.750 346.500 114.600 ;
        RECT 348.000 111.750 349.800 115.950 ;
        RECT 352.200 111.750 354.000 117.600 ;
        RECT 359.400 114.600 360.600 122.850 ;
        RECT 374.400 121.650 375.600 125.850 ;
        RECT 356.550 111.750 358.350 114.600 ;
        RECT 359.550 111.750 361.350 114.600 ;
        RECT 365.700 111.750 367.500 120.600 ;
        RECT 371.100 120.000 375.600 121.650 ;
        RECT 383.400 121.650 384.600 125.850 ;
        RECT 394.950 122.850 397.050 124.950 ;
        RECT 398.100 123.150 399.900 124.950 ;
        RECT 383.400 120.000 387.900 121.650 ;
        RECT 395.100 121.050 396.900 122.850 ;
        RECT 397.950 121.050 400.050 123.150 ;
        RECT 400.950 122.850 403.050 124.950 ;
        RECT 403.950 124.050 406.050 126.150 ;
        RECT 412.950 125.850 415.050 127.950 ;
        RECT 415.950 127.050 418.050 129.150 ;
        RECT 413.100 124.050 414.900 125.850 ;
        RECT 401.100 121.050 402.900 122.850 ;
        RECT 371.100 111.750 372.900 120.000 ;
        RECT 386.100 111.750 387.900 120.000 ;
        RECT 391.500 111.750 393.300 120.600 ;
        RECT 404.700 117.600 405.900 124.050 ;
        RECT 416.250 119.700 417.450 127.050 ;
        RECT 418.950 125.850 421.050 127.950 ;
        RECT 425.250 126.150 427.050 127.950 ;
        RECT 431.250 126.150 432.450 131.400 ;
        RECT 437.100 126.150 438.900 127.950 ;
        RECT 419.100 124.050 420.900 125.850 ;
        RECT 424.950 124.050 427.050 126.150 ;
        RECT 427.950 122.850 430.050 124.950 ;
        RECT 430.950 124.050 433.050 126.150 ;
        RECT 428.700 121.050 430.500 122.850 ;
        RECT 431.400 120.150 432.600 124.050 ;
        RECT 433.950 122.850 436.050 124.950 ;
        RECT 436.950 124.050 439.050 126.150 ;
        RECT 443.400 124.950 444.600 137.400 ;
        RECT 453.450 131.400 455.250 143.250 ;
        RECT 457.650 131.400 459.450 143.250 ;
        RECT 465.450 131.400 467.250 143.250 ;
        RECT 469.650 131.400 471.450 143.250 ;
        RECT 473.550 137.400 475.350 143.250 ;
        RECT 476.550 137.400 478.350 143.250 ;
        RECT 453.450 130.350 456.000 131.400 ;
        RECT 465.450 130.350 468.000 131.400 ;
        RECT 452.100 126.150 453.900 127.950 ;
        RECT 442.950 122.850 445.050 124.950 ;
        RECT 446.100 123.150 447.900 124.950 ;
        RECT 451.950 124.050 454.050 126.150 ;
        RECT 454.950 123.150 456.000 130.350 ;
        RECT 458.100 126.150 459.900 127.950 ;
        RECT 464.100 126.150 465.900 127.950 ;
        RECT 457.950 124.050 460.050 126.150 ;
        RECT 463.950 124.050 466.050 126.150 ;
        RECT 466.950 123.150 468.000 130.350 ;
        RECT 470.100 126.150 471.900 127.950 ;
        RECT 469.950 124.050 472.050 126.150 ;
        RECT 476.400 124.950 477.600 137.400 ;
        RECT 483.300 131.400 485.100 143.250 ;
        RECT 487.500 131.400 489.300 143.250 ;
        RECT 490.800 137.400 492.600 143.250 ;
        RECT 497.550 137.400 499.350 143.250 ;
        RECT 500.550 137.400 502.350 143.250 ;
        RECT 503.550 137.400 505.350 143.250 ;
        RECT 482.100 126.150 483.900 127.950 ;
        RECT 487.950 126.150 489.150 131.400 ;
        RECT 490.950 129.150 492.750 130.950 ;
        RECT 500.550 129.150 501.750 137.400 ;
        RECT 509.550 131.400 511.350 143.250 ;
        RECT 512.550 140.400 514.350 143.250 ;
        RECT 517.050 137.400 518.850 143.250 ;
        RECT 521.250 137.400 523.050 143.250 ;
        RECT 514.950 135.300 518.850 137.400 ;
        RECT 525.150 136.500 526.950 143.250 ;
        RECT 528.150 137.400 529.950 143.250 ;
        RECT 532.950 137.400 534.750 143.250 ;
        RECT 538.050 137.400 539.850 143.250 ;
        RECT 533.250 136.500 534.450 137.400 ;
        RECT 523.950 134.700 530.850 136.500 ;
        RECT 533.250 134.400 538.050 136.500 ;
        RECT 516.150 132.600 518.850 134.400 ;
        RECT 519.750 133.800 521.550 134.400 ;
        RECT 519.750 132.900 526.050 133.800 ;
        RECT 533.250 133.500 534.450 134.400 ;
        RECT 519.750 132.600 521.550 132.900 ;
        RECT 517.950 131.700 518.850 132.600 ;
        RECT 490.950 127.050 493.050 129.150 ;
        RECT 473.100 123.150 474.900 124.950 ;
        RECT 434.100 121.050 435.900 122.850 ;
        RECT 396.000 111.750 397.800 117.600 ;
        RECT 400.200 115.950 405.900 117.600 ;
        RECT 413.850 118.800 417.450 119.700 ;
        RECT 428.250 119.100 432.600 120.150 ;
        RECT 400.200 111.750 402.000 115.950 ;
        RECT 403.500 111.750 405.300 114.600 ;
        RECT 413.850 111.750 415.650 118.800 ;
        RECT 428.250 117.600 429.150 119.100 ;
        RECT 418.350 111.750 420.150 117.600 ;
        RECT 424.650 112.500 426.450 117.600 ;
        RECT 427.650 113.400 429.450 117.600 ;
        RECT 430.650 117.000 438.450 117.900 ;
        RECT 430.650 112.500 432.450 117.000 ;
        RECT 424.650 111.750 432.450 112.500 ;
        RECT 433.650 111.750 435.450 116.100 ;
        RECT 436.650 111.750 438.450 117.000 ;
        RECT 443.400 114.600 444.600 122.850 ;
        RECT 445.950 121.050 448.050 123.150 ;
        RECT 454.950 121.050 457.050 123.150 ;
        RECT 466.950 121.050 469.050 123.150 ;
        RECT 472.950 121.050 475.050 123.150 ;
        RECT 475.950 122.850 478.050 124.950 ;
        RECT 481.950 124.050 484.050 126.150 ;
        RECT 484.950 122.850 487.050 124.950 ;
        RECT 487.950 124.050 490.050 126.150 ;
        RECT 496.950 125.850 499.050 127.950 ;
        RECT 499.950 127.050 502.050 129.150 ;
        RECT 497.100 124.050 498.900 125.850 ;
        RECT 454.950 114.600 456.000 121.050 ;
        RECT 466.950 114.600 468.000 121.050 ;
        RECT 476.400 114.600 477.600 122.850 ;
        RECT 485.100 121.050 486.900 122.850 ;
        RECT 488.850 120.750 490.050 124.050 ;
        RECT 489.000 119.700 492.750 120.750 ;
        RECT 482.550 116.700 490.350 118.050 ;
        RECT 442.650 111.750 444.450 114.600 ;
        RECT 445.650 111.750 447.450 114.600 ;
        RECT 451.650 111.750 453.450 114.600 ;
        RECT 454.650 111.750 456.450 114.600 ;
        RECT 457.650 111.750 459.450 114.600 ;
        RECT 463.650 111.750 465.450 114.600 ;
        RECT 466.650 111.750 468.450 114.600 ;
        RECT 469.650 111.750 471.450 114.600 ;
        RECT 473.550 111.750 475.350 114.600 ;
        RECT 476.550 111.750 478.350 114.600 ;
        RECT 482.550 111.750 484.350 116.700 ;
        RECT 485.550 111.750 487.350 115.800 ;
        RECT 488.550 111.750 490.350 116.700 ;
        RECT 491.550 117.600 492.750 119.700 ;
        RECT 500.550 119.700 501.750 127.050 ;
        RECT 502.950 125.850 505.050 127.950 ;
        RECT 503.100 124.050 504.900 125.850 ;
        RECT 509.550 121.950 510.750 131.400 ;
        RECT 514.950 130.800 517.050 131.700 ;
        RECT 517.950 130.800 523.950 131.700 ;
        RECT 512.850 129.600 517.050 130.800 ;
        RECT 511.950 127.800 513.750 129.600 ;
        RECT 523.050 126.150 523.950 130.800 ;
        RECT 525.150 130.800 526.050 132.900 ;
        RECT 526.950 132.300 534.450 133.500 ;
        RECT 526.950 131.700 528.750 132.300 ;
        RECT 541.050 131.400 542.850 143.250 ;
        RECT 531.750 130.800 542.850 131.400 ;
        RECT 525.150 130.200 542.850 130.800 ;
        RECT 525.150 129.900 533.550 130.200 ;
        RECT 531.750 129.600 533.550 129.900 ;
        RECT 523.050 124.050 526.050 126.150 ;
        RECT 529.950 125.100 532.050 126.150 ;
        RECT 529.950 124.050 537.900 125.100 ;
        RECT 511.950 123.750 514.050 124.050 ;
        RECT 511.950 121.950 515.850 123.750 ;
        RECT 509.550 119.850 514.050 121.950 ;
        RECT 523.050 120.000 523.950 124.050 ;
        RECT 536.100 123.300 537.900 124.050 ;
        RECT 539.100 123.150 540.900 124.950 ;
        RECT 533.100 122.400 534.900 123.000 ;
        RECT 539.100 122.400 540.000 123.150 ;
        RECT 533.100 121.200 540.000 122.400 ;
        RECT 533.100 120.000 534.150 121.200 ;
        RECT 500.550 118.800 504.150 119.700 ;
        RECT 491.550 111.750 493.350 117.600 ;
        RECT 497.850 111.750 499.650 117.600 ;
        RECT 502.350 111.750 504.150 118.800 ;
        RECT 509.550 117.600 510.750 119.850 ;
        RECT 523.050 119.100 534.150 120.000 ;
        RECT 523.050 118.800 523.950 119.100 ;
        RECT 509.550 111.750 511.350 117.600 ;
        RECT 514.950 116.700 517.050 117.600 ;
        RECT 522.150 117.000 523.950 118.800 ;
        RECT 533.100 118.200 534.150 119.100 ;
        RECT 529.350 117.450 531.150 118.200 ;
        RECT 514.950 115.500 518.700 116.700 ;
        RECT 517.650 114.600 518.700 115.500 ;
        RECT 526.200 116.400 531.150 117.450 ;
        RECT 532.650 116.400 534.450 118.200 ;
        RECT 541.950 117.600 542.850 130.200 ;
        RECT 545.550 137.400 547.350 143.250 ;
        RECT 545.550 130.500 546.750 137.400 ;
        RECT 548.850 131.400 550.650 143.250 ;
        RECT 551.850 131.400 553.650 143.250 ;
        RECT 558.150 131.400 559.950 143.250 ;
        RECT 561.150 137.400 562.950 143.250 ;
        RECT 566.250 137.400 568.050 143.250 ;
        RECT 571.050 137.400 572.850 143.250 ;
        RECT 566.550 136.500 567.750 137.400 ;
        RECT 574.050 136.500 575.850 143.250 ;
        RECT 577.950 137.400 579.750 143.250 ;
        RECT 582.150 137.400 583.950 143.250 ;
        RECT 586.650 140.400 588.450 143.250 ;
        RECT 562.950 134.400 567.750 136.500 ;
        RECT 570.150 134.700 577.050 136.500 ;
        RECT 582.150 135.300 586.050 137.400 ;
        RECT 566.550 133.500 567.750 134.400 ;
        RECT 579.450 133.800 581.250 134.400 ;
        RECT 566.550 132.300 574.050 133.500 ;
        RECT 572.250 131.700 574.050 132.300 ;
        RECT 574.950 132.900 581.250 133.800 ;
        RECT 545.550 129.600 551.250 130.500 ;
        RECT 549.000 128.700 551.250 129.600 ;
        RECT 545.100 126.150 546.900 127.950 ;
        RECT 544.950 124.050 547.050 126.150 ;
        RECT 549.000 120.300 550.050 128.700 ;
        RECT 552.150 126.150 553.350 131.400 ;
        RECT 550.950 124.050 553.350 126.150 ;
        RECT 549.000 119.400 551.250 120.300 ;
        RECT 526.200 114.600 527.250 116.400 ;
        RECT 535.950 115.500 538.050 117.600 ;
        RECT 535.950 114.600 537.000 115.500 ;
        RECT 512.850 111.750 514.650 114.600 ;
        RECT 517.350 111.750 519.150 114.600 ;
        RECT 521.550 111.750 523.350 114.600 ;
        RECT 525.450 111.750 527.250 114.600 ;
        RECT 528.750 111.750 530.550 114.600 ;
        RECT 533.250 113.700 537.000 114.600 ;
        RECT 533.250 111.750 535.050 113.700 ;
        RECT 538.050 111.750 539.850 114.600 ;
        RECT 541.050 111.750 542.850 117.600 ;
        RECT 546.150 118.500 551.250 119.400 ;
        RECT 546.150 114.600 547.350 118.500 ;
        RECT 552.150 117.600 553.350 124.050 ;
        RECT 558.150 130.800 569.250 131.400 ;
        RECT 574.950 130.800 575.850 132.900 ;
        RECT 579.450 132.600 581.250 132.900 ;
        RECT 582.150 132.600 584.850 134.400 ;
        RECT 582.150 131.700 583.050 132.600 ;
        RECT 558.150 130.200 575.850 130.800 ;
        RECT 558.150 117.600 559.050 130.200 ;
        RECT 567.450 129.900 575.850 130.200 ;
        RECT 577.050 130.800 583.050 131.700 ;
        RECT 583.950 130.800 586.050 131.700 ;
        RECT 589.650 131.400 591.450 143.250 ;
        RECT 596.400 137.400 598.200 143.250 ;
        RECT 599.700 131.400 601.500 143.250 ;
        RECT 603.900 131.400 605.700 143.250 ;
        RECT 608.550 131.400 610.350 143.250 ;
        RECT 611.550 140.400 613.350 143.250 ;
        RECT 616.050 137.400 617.850 143.250 ;
        RECT 620.250 137.400 622.050 143.250 ;
        RECT 613.950 135.300 617.850 137.400 ;
        RECT 624.150 136.500 625.950 143.250 ;
        RECT 627.150 137.400 628.950 143.250 ;
        RECT 631.950 137.400 633.750 143.250 ;
        RECT 637.050 137.400 638.850 143.250 ;
        RECT 632.250 136.500 633.450 137.400 ;
        RECT 622.950 134.700 629.850 136.500 ;
        RECT 632.250 134.400 637.050 136.500 ;
        RECT 615.150 132.600 617.850 134.400 ;
        RECT 618.750 133.800 620.550 134.400 ;
        RECT 618.750 132.900 625.050 133.800 ;
        RECT 632.250 133.500 633.450 134.400 ;
        RECT 618.750 132.600 620.550 132.900 ;
        RECT 616.950 131.700 617.850 132.600 ;
        RECT 567.450 129.600 569.250 129.900 ;
        RECT 577.050 126.150 577.950 130.800 ;
        RECT 583.950 129.600 588.150 130.800 ;
        RECT 587.250 127.800 589.050 129.600 ;
        RECT 568.950 125.100 571.050 126.150 ;
        RECT 560.100 123.150 561.900 124.950 ;
        RECT 563.100 124.050 571.050 125.100 ;
        RECT 574.950 124.050 577.950 126.150 ;
        RECT 563.100 123.300 564.900 124.050 ;
        RECT 561.000 122.400 561.900 123.150 ;
        RECT 566.100 122.400 567.900 123.000 ;
        RECT 561.000 121.200 567.900 122.400 ;
        RECT 566.850 120.000 567.900 121.200 ;
        RECT 577.050 120.000 577.950 124.050 ;
        RECT 586.950 123.750 589.050 124.050 ;
        RECT 585.150 121.950 589.050 123.750 ;
        RECT 590.250 121.950 591.450 131.400 ;
        RECT 596.250 129.150 598.050 130.950 ;
        RECT 595.950 127.050 598.050 129.150 ;
        RECT 599.850 126.150 601.050 131.400 ;
        RECT 605.100 126.150 606.900 127.950 ;
        RECT 566.850 119.100 577.950 120.000 ;
        RECT 586.950 119.850 591.450 121.950 ;
        RECT 598.950 124.050 601.050 126.150 ;
        RECT 598.950 120.750 600.150 124.050 ;
        RECT 601.950 122.850 604.050 124.950 ;
        RECT 604.950 124.050 607.050 126.150 ;
        RECT 602.100 121.050 603.900 122.850 ;
        RECT 608.550 121.950 609.750 131.400 ;
        RECT 613.950 130.800 616.050 131.700 ;
        RECT 616.950 130.800 622.950 131.700 ;
        RECT 611.850 129.600 616.050 130.800 ;
        RECT 610.950 127.800 612.750 129.600 ;
        RECT 622.050 126.150 622.950 130.800 ;
        RECT 624.150 130.800 625.050 132.900 ;
        RECT 625.950 132.300 633.450 133.500 ;
        RECT 625.950 131.700 627.750 132.300 ;
        RECT 640.050 131.400 641.850 143.250 ;
        RECT 630.750 130.800 641.850 131.400 ;
        RECT 624.150 130.200 641.850 130.800 ;
        RECT 624.150 129.900 632.550 130.200 ;
        RECT 630.750 129.600 632.550 129.900 ;
        RECT 622.050 124.050 625.050 126.150 ;
        RECT 628.950 125.100 631.050 126.150 ;
        RECT 628.950 124.050 636.900 125.100 ;
        RECT 610.950 123.750 613.050 124.050 ;
        RECT 610.950 121.950 614.850 123.750 ;
        RECT 566.850 118.200 567.900 119.100 ;
        RECT 577.050 118.800 577.950 119.100 ;
        RECT 545.550 111.750 547.350 114.600 ;
        RECT 548.850 111.750 550.650 117.600 ;
        RECT 551.850 111.750 553.650 117.600 ;
        RECT 558.150 111.750 559.950 117.600 ;
        RECT 562.950 115.500 565.050 117.600 ;
        RECT 566.550 116.400 568.350 118.200 ;
        RECT 569.850 117.450 571.650 118.200 ;
        RECT 569.850 116.400 574.800 117.450 ;
        RECT 577.050 117.000 578.850 118.800 ;
        RECT 590.250 117.600 591.450 119.850 ;
        RECT 596.250 119.700 600.000 120.750 ;
        RECT 608.550 119.850 613.050 121.950 ;
        RECT 622.050 120.000 622.950 124.050 ;
        RECT 635.100 123.300 636.900 124.050 ;
        RECT 638.100 123.150 639.900 124.950 ;
        RECT 632.100 122.400 633.900 123.000 ;
        RECT 638.100 122.400 639.000 123.150 ;
        RECT 632.100 121.200 639.000 122.400 ;
        RECT 632.100 120.000 633.150 121.200 ;
        RECT 596.250 117.600 597.450 119.700 ;
        RECT 583.950 116.700 586.050 117.600 ;
        RECT 564.000 114.600 565.050 115.500 ;
        RECT 573.750 114.600 574.800 116.400 ;
        RECT 582.300 115.500 586.050 116.700 ;
        RECT 582.300 114.600 583.350 115.500 ;
        RECT 561.150 111.750 562.950 114.600 ;
        RECT 564.000 113.700 567.750 114.600 ;
        RECT 565.950 111.750 567.750 113.700 ;
        RECT 570.450 111.750 572.250 114.600 ;
        RECT 573.750 111.750 575.550 114.600 ;
        RECT 577.650 111.750 579.450 114.600 ;
        RECT 581.850 111.750 583.650 114.600 ;
        RECT 586.350 111.750 588.150 114.600 ;
        RECT 589.650 111.750 591.450 117.600 ;
        RECT 595.650 111.750 597.450 117.600 ;
        RECT 598.650 116.700 606.450 118.050 ;
        RECT 598.650 111.750 600.450 116.700 ;
        RECT 601.650 111.750 603.450 115.800 ;
        RECT 604.650 111.750 606.450 116.700 ;
        RECT 608.550 117.600 609.750 119.850 ;
        RECT 622.050 119.100 633.150 120.000 ;
        RECT 622.050 118.800 622.950 119.100 ;
        RECT 608.550 111.750 610.350 117.600 ;
        RECT 613.950 116.700 616.050 117.600 ;
        RECT 621.150 117.000 622.950 118.800 ;
        RECT 632.100 118.200 633.150 119.100 ;
        RECT 628.350 117.450 630.150 118.200 ;
        RECT 613.950 115.500 617.700 116.700 ;
        RECT 616.650 114.600 617.700 115.500 ;
        RECT 625.200 116.400 630.150 117.450 ;
        RECT 631.650 116.400 633.450 118.200 ;
        RECT 640.950 117.600 641.850 130.200 ;
        RECT 625.200 114.600 626.250 116.400 ;
        RECT 634.950 115.500 637.050 117.600 ;
        RECT 634.950 114.600 636.000 115.500 ;
        RECT 611.850 111.750 613.650 114.600 ;
        RECT 616.350 111.750 618.150 114.600 ;
        RECT 620.550 111.750 622.350 114.600 ;
        RECT 624.450 111.750 626.250 114.600 ;
        RECT 627.750 111.750 629.550 114.600 ;
        RECT 632.250 113.700 636.000 114.600 ;
        RECT 632.250 111.750 634.050 113.700 ;
        RECT 637.050 111.750 638.850 114.600 ;
        RECT 640.050 111.750 641.850 117.600 ;
        RECT 645.150 131.400 646.950 143.250 ;
        RECT 648.150 137.400 649.950 143.250 ;
        RECT 653.250 137.400 655.050 143.250 ;
        RECT 658.050 137.400 659.850 143.250 ;
        RECT 653.550 136.500 654.750 137.400 ;
        RECT 661.050 136.500 662.850 143.250 ;
        RECT 664.950 137.400 666.750 143.250 ;
        RECT 669.150 137.400 670.950 143.250 ;
        RECT 673.650 140.400 675.450 143.250 ;
        RECT 649.950 134.400 654.750 136.500 ;
        RECT 657.150 134.700 664.050 136.500 ;
        RECT 669.150 135.300 673.050 137.400 ;
        RECT 653.550 133.500 654.750 134.400 ;
        RECT 666.450 133.800 668.250 134.400 ;
        RECT 653.550 132.300 661.050 133.500 ;
        RECT 659.250 131.700 661.050 132.300 ;
        RECT 661.950 132.900 668.250 133.800 ;
        RECT 645.150 130.800 656.250 131.400 ;
        RECT 661.950 130.800 662.850 132.900 ;
        RECT 666.450 132.600 668.250 132.900 ;
        RECT 669.150 132.600 671.850 134.400 ;
        RECT 669.150 131.700 670.050 132.600 ;
        RECT 645.150 130.200 662.850 130.800 ;
        RECT 645.150 117.600 646.050 130.200 ;
        RECT 654.450 129.900 662.850 130.200 ;
        RECT 664.050 130.800 670.050 131.700 ;
        RECT 670.950 130.800 673.050 131.700 ;
        RECT 676.650 131.400 678.450 143.250 ;
        RECT 681.300 131.400 683.100 143.250 ;
        RECT 685.500 131.400 687.300 143.250 ;
        RECT 688.800 137.400 690.600 143.250 ;
        RECT 696.300 131.400 698.100 143.250 ;
        RECT 700.500 131.400 702.300 143.250 ;
        RECT 703.800 137.400 705.600 143.250 ;
        RECT 654.450 129.600 656.250 129.900 ;
        RECT 664.050 126.150 664.950 130.800 ;
        RECT 670.950 129.600 675.150 130.800 ;
        RECT 674.250 127.800 676.050 129.600 ;
        RECT 655.950 125.100 658.050 126.150 ;
        RECT 647.100 123.150 648.900 124.950 ;
        RECT 650.100 124.050 658.050 125.100 ;
        RECT 661.950 124.050 664.950 126.150 ;
        RECT 650.100 123.300 651.900 124.050 ;
        RECT 648.000 122.400 648.900 123.150 ;
        RECT 653.100 122.400 654.900 123.000 ;
        RECT 648.000 121.200 654.900 122.400 ;
        RECT 653.850 120.000 654.900 121.200 ;
        RECT 664.050 120.000 664.950 124.050 ;
        RECT 673.950 123.750 676.050 124.050 ;
        RECT 672.150 121.950 676.050 123.750 ;
        RECT 677.250 121.950 678.450 131.400 ;
        RECT 680.100 126.150 681.900 127.950 ;
        RECT 685.950 126.150 687.150 131.400 ;
        RECT 688.950 129.150 690.750 130.950 ;
        RECT 688.950 127.050 691.050 129.150 ;
        RECT 695.100 126.150 696.900 127.950 ;
        RECT 700.950 126.150 702.150 131.400 ;
        RECT 703.950 129.150 705.750 130.950 ;
        RECT 703.950 127.050 706.050 129.150 ;
        RECT 679.950 124.050 682.050 126.150 ;
        RECT 682.950 122.850 685.050 124.950 ;
        RECT 685.950 124.050 688.050 126.150 ;
        RECT 694.950 124.050 697.050 126.150 ;
        RECT 653.850 119.100 664.950 120.000 ;
        RECT 673.950 119.850 678.450 121.950 ;
        RECT 683.100 121.050 684.900 122.850 ;
        RECT 686.850 120.750 688.050 124.050 ;
        RECT 697.950 122.850 700.050 124.950 ;
        RECT 700.950 124.050 703.050 126.150 ;
        RECT 698.100 121.050 699.900 122.850 ;
        RECT 701.850 120.750 703.050 124.050 ;
        RECT 653.850 118.200 654.900 119.100 ;
        RECT 664.050 118.800 664.950 119.100 ;
        RECT 645.150 111.750 646.950 117.600 ;
        RECT 649.950 115.500 652.050 117.600 ;
        RECT 653.550 116.400 655.350 118.200 ;
        RECT 656.850 117.450 658.650 118.200 ;
        RECT 656.850 116.400 661.800 117.450 ;
        RECT 664.050 117.000 665.850 118.800 ;
        RECT 677.250 117.600 678.450 119.850 ;
        RECT 687.000 119.700 690.750 120.750 ;
        RECT 702.000 119.700 705.750 120.750 ;
        RECT 670.950 116.700 673.050 117.600 ;
        RECT 651.000 114.600 652.050 115.500 ;
        RECT 660.750 114.600 661.800 116.400 ;
        RECT 669.300 115.500 673.050 116.700 ;
        RECT 669.300 114.600 670.350 115.500 ;
        RECT 648.150 111.750 649.950 114.600 ;
        RECT 651.000 113.700 654.750 114.600 ;
        RECT 652.950 111.750 654.750 113.700 ;
        RECT 657.450 111.750 659.250 114.600 ;
        RECT 660.750 111.750 662.550 114.600 ;
        RECT 664.650 111.750 666.450 114.600 ;
        RECT 668.850 111.750 670.650 114.600 ;
        RECT 673.350 111.750 675.150 114.600 ;
        RECT 676.650 111.750 678.450 117.600 ;
        RECT 680.550 116.700 688.350 118.050 ;
        RECT 680.550 111.750 682.350 116.700 ;
        RECT 683.550 111.750 685.350 115.800 ;
        RECT 686.550 111.750 688.350 116.700 ;
        RECT 689.550 117.600 690.750 119.700 ;
        RECT 689.550 111.750 691.350 117.600 ;
        RECT 695.550 116.700 703.350 118.050 ;
        RECT 695.550 111.750 697.350 116.700 ;
        RECT 698.550 111.750 700.350 115.800 ;
        RECT 701.550 111.750 703.350 116.700 ;
        RECT 704.550 117.600 705.750 119.700 ;
        RECT 704.550 111.750 706.350 117.600 ;
        RECT 4.650 104.400 6.450 107.250 ;
        RECT 7.650 104.400 9.450 107.250 ;
        RECT 10.650 104.400 12.450 107.250 ;
        RECT 17.700 104.400 19.500 107.250 ;
        RECT 7.950 97.950 9.000 104.400 ;
        RECT 21.000 103.050 22.800 107.250 ;
        RECT 17.100 101.400 22.800 103.050 ;
        RECT 25.200 101.400 27.000 107.250 ;
        RECT 29.550 104.400 31.350 107.250 ;
        RECT 32.550 104.400 34.350 107.250 ;
        RECT 41.700 104.400 43.500 107.250 ;
        RECT 7.950 95.850 10.050 97.950 ;
        RECT 4.950 92.850 7.050 94.950 ;
        RECT 5.100 91.050 6.900 92.850 ;
        RECT 7.950 88.650 9.000 95.850 ;
        RECT 17.100 94.950 18.300 101.400 ;
        RECT 20.100 96.150 21.900 97.950 ;
        RECT 10.950 92.850 13.050 94.950 ;
        RECT 16.950 92.850 19.050 94.950 ;
        RECT 19.950 94.050 22.050 96.150 ;
        RECT 22.950 95.850 25.050 97.950 ;
        RECT 26.100 96.150 27.900 97.950 ;
        RECT 23.100 94.050 24.900 95.850 ;
        RECT 25.950 94.050 28.050 96.150 ;
        RECT 28.950 95.850 31.050 97.950 ;
        RECT 32.400 96.150 33.600 104.400 ;
        RECT 45.000 103.050 46.800 107.250 ;
        RECT 41.100 101.400 46.800 103.050 ;
        RECT 49.200 101.400 51.000 107.250 ;
        RECT 29.100 94.050 30.900 95.850 ;
        RECT 31.950 94.050 34.050 96.150 ;
        RECT 41.100 94.950 42.300 101.400 ;
        RECT 53.700 98.400 55.500 107.250 ;
        RECT 59.100 99.000 60.900 107.250 ;
        RECT 70.650 101.400 72.450 107.250 ;
        RECT 71.250 99.300 72.450 101.400 ;
        RECT 73.650 102.300 75.450 107.250 ;
        RECT 76.650 103.200 78.450 107.250 ;
        RECT 79.650 102.300 81.450 107.250 ;
        RECT 73.650 100.950 81.450 102.300 ;
        RECT 85.350 101.400 87.150 107.250 ;
        RECT 88.350 101.400 90.150 107.250 ;
        RECT 91.650 104.400 93.450 107.250 ;
        RECT 44.100 96.150 45.900 97.950 ;
        RECT 11.100 91.050 12.900 92.850 ;
        RECT 6.450 87.600 9.000 88.650 ;
        RECT 17.100 87.600 18.300 92.850 ;
        RECT 6.450 75.750 8.250 87.600 ;
        RECT 10.650 75.750 12.450 87.600 ;
        RECT 16.650 75.750 18.450 87.600 ;
        RECT 19.650 86.700 27.450 87.600 ;
        RECT 19.650 75.750 21.450 86.700 ;
        RECT 22.650 75.750 24.450 85.800 ;
        RECT 25.650 75.750 27.450 86.700 ;
        RECT 32.400 81.600 33.600 94.050 ;
        RECT 40.950 92.850 43.050 94.950 ;
        RECT 43.950 94.050 46.050 96.150 ;
        RECT 46.950 95.850 49.050 97.950 ;
        RECT 50.100 96.150 51.900 97.950 ;
        RECT 59.100 97.350 63.600 99.000 ;
        RECT 71.250 98.250 75.000 99.300 ;
        RECT 47.100 94.050 48.900 95.850 ;
        RECT 49.950 94.050 52.050 96.150 ;
        RECT 62.400 93.150 63.600 97.350 ;
        RECT 73.950 94.950 75.150 98.250 ;
        RECT 77.100 96.150 78.900 97.950 ;
        RECT 41.100 87.600 42.300 92.850 ;
        RECT 52.950 89.850 55.050 91.950 ;
        RECT 58.950 89.850 61.050 91.950 ;
        RECT 61.950 91.050 64.050 93.150 ;
        RECT 73.950 92.850 76.050 94.950 ;
        RECT 76.950 94.050 79.050 96.150 ;
        RECT 85.650 94.950 86.850 101.400 ;
        RECT 91.650 100.500 92.850 104.400 ;
        RECT 97.650 101.400 99.450 107.250 ;
        RECT 87.750 99.600 92.850 100.500 ;
        RECT 87.750 98.700 90.000 99.600 ;
        RECT 79.950 92.850 82.050 94.950 ;
        RECT 85.650 92.850 88.050 94.950 ;
        RECT 53.100 88.050 54.900 89.850 ;
        RECT 29.550 75.750 31.350 81.600 ;
        RECT 32.550 75.750 34.350 81.600 ;
        RECT 40.650 75.750 42.450 87.600 ;
        RECT 43.650 86.700 51.450 87.600 ;
        RECT 55.950 86.850 58.050 88.950 ;
        RECT 59.250 88.050 61.050 89.850 ;
        RECT 43.650 75.750 45.450 86.700 ;
        RECT 46.650 75.750 48.450 85.800 ;
        RECT 49.650 75.750 51.450 86.700 ;
        RECT 56.100 85.050 57.900 86.850 ;
        RECT 62.700 82.800 63.750 91.050 ;
        RECT 70.950 89.850 73.050 91.950 ;
        RECT 71.250 88.050 73.050 89.850 ;
        RECT 74.850 87.600 76.050 92.850 ;
        RECT 80.100 91.050 81.900 92.850 ;
        RECT 85.650 87.600 86.850 92.850 ;
        RECT 88.950 90.300 90.000 98.700 ;
        RECT 98.250 99.300 99.450 101.400 ;
        RECT 100.650 102.300 102.450 107.250 ;
        RECT 103.650 103.200 105.450 107.250 ;
        RECT 106.650 102.300 108.450 107.250 ;
        RECT 100.650 100.950 108.450 102.300 ;
        RECT 112.350 101.400 114.150 107.250 ;
        RECT 115.350 101.400 117.150 107.250 ;
        RECT 118.650 104.400 120.450 107.250 ;
        RECT 98.250 98.250 102.000 99.300 ;
        RECT 100.950 94.950 102.150 98.250 ;
        RECT 104.100 96.150 105.900 97.950 ;
        RECT 91.950 92.850 94.050 94.950 ;
        RECT 100.950 92.850 103.050 94.950 ;
        RECT 103.950 94.050 106.050 96.150 ;
        RECT 112.650 94.950 113.850 101.400 ;
        RECT 118.650 100.500 119.850 104.400 ;
        RECT 114.750 99.600 119.850 100.500 ;
        RECT 122.550 99.900 124.350 107.250 ;
        RECT 127.050 101.400 128.850 107.250 ;
        RECT 130.050 102.900 131.850 107.250 ;
        RECT 130.050 101.400 133.350 102.900 ;
        RECT 128.250 99.900 130.050 100.500 ;
        RECT 114.750 98.700 117.000 99.600 ;
        RECT 122.550 98.700 130.050 99.900 ;
        RECT 106.950 92.850 109.050 94.950 ;
        RECT 112.650 92.850 115.050 94.950 ;
        RECT 92.100 91.050 93.900 92.850 ;
        RECT 87.750 89.400 90.000 90.300 ;
        RECT 97.950 89.850 100.050 91.950 ;
        RECT 87.750 88.500 93.450 89.400 ;
        RECT 56.700 81.900 63.750 82.800 ;
        RECT 56.700 81.600 58.350 81.900 ;
        RECT 53.550 75.750 55.350 81.600 ;
        RECT 56.550 75.750 58.350 81.600 ;
        RECT 62.550 81.600 63.750 81.900 ;
        RECT 59.550 75.750 61.350 81.000 ;
        RECT 62.550 75.750 64.350 81.600 ;
        RECT 71.400 75.750 73.200 81.600 ;
        RECT 74.700 75.750 76.500 87.600 ;
        RECT 78.900 75.750 80.700 87.600 ;
        RECT 85.350 75.750 87.150 87.600 ;
        RECT 88.350 75.750 90.150 87.600 ;
        RECT 92.250 81.600 93.450 88.500 ;
        RECT 98.250 88.050 100.050 89.850 ;
        RECT 101.850 87.600 103.050 92.850 ;
        RECT 107.100 91.050 108.900 92.850 ;
        RECT 112.650 87.600 113.850 92.850 ;
        RECT 115.950 90.300 117.000 98.700 ;
        RECT 118.950 92.850 121.050 94.950 ;
        RECT 121.950 92.850 124.050 94.950 ;
        RECT 119.100 91.050 120.900 92.850 ;
        RECT 122.100 91.050 123.900 92.850 ;
        RECT 114.750 89.400 117.000 90.300 ;
        RECT 114.750 88.500 120.450 89.400 ;
        RECT 91.650 75.750 93.450 81.600 ;
        RECT 98.400 75.750 100.200 81.600 ;
        RECT 101.700 75.750 103.500 87.600 ;
        RECT 105.900 75.750 107.700 87.600 ;
        RECT 112.350 75.750 114.150 87.600 ;
        RECT 115.350 75.750 117.150 87.600 ;
        RECT 119.250 81.600 120.450 88.500 ;
        RECT 125.700 81.600 126.900 98.700 ;
        RECT 132.150 94.950 133.350 101.400 ;
        RECT 137.550 102.300 139.350 107.250 ;
        RECT 140.550 103.200 142.350 107.250 ;
        RECT 143.550 102.300 145.350 107.250 ;
        RECT 137.550 100.950 145.350 102.300 ;
        RECT 146.550 101.400 148.350 107.250 ;
        RECT 154.650 101.400 156.450 107.250 ;
        RECT 146.550 99.300 147.750 101.400 ;
        RECT 144.000 98.250 147.750 99.300 ;
        RECT 155.250 99.300 156.450 101.400 ;
        RECT 157.650 102.300 159.450 107.250 ;
        RECT 160.650 103.200 162.450 107.250 ;
        RECT 163.650 102.300 165.450 107.250 ;
        RECT 157.650 100.950 165.450 102.300 ;
        RECT 169.650 101.400 171.450 107.250 ;
        RECT 172.650 101.400 174.450 107.250 ;
        RECT 177.000 101.400 178.800 107.250 ;
        RECT 181.200 103.050 183.000 107.250 ;
        RECT 184.500 104.400 186.300 107.250 ;
        RECT 193.650 104.400 195.450 107.250 ;
        RECT 196.650 104.400 198.450 107.250 ;
        RECT 181.200 101.400 186.900 103.050 ;
        RECT 155.250 98.250 159.000 99.300 ;
        RECT 140.100 96.150 141.900 97.950 ;
        RECT 128.100 93.150 129.900 94.950 ;
        RECT 127.950 91.050 130.050 93.150 ;
        RECT 130.950 92.850 133.350 94.950 ;
        RECT 136.950 92.850 139.050 94.950 ;
        RECT 139.950 94.050 142.050 96.150 ;
        RECT 143.850 94.950 145.050 98.250 ;
        RECT 142.950 92.850 145.050 94.950 ;
        RECT 157.950 94.950 159.150 98.250 ;
        RECT 161.100 96.150 162.900 97.950 ;
        RECT 157.950 92.850 160.050 94.950 ;
        RECT 160.950 94.050 163.050 96.150 ;
        RECT 170.400 94.950 171.600 101.400 ;
        RECT 173.100 96.150 174.900 97.950 ;
        RECT 176.100 96.150 177.900 97.950 ;
        RECT 163.950 92.850 166.050 94.950 ;
        RECT 169.950 92.850 172.050 94.950 ;
        RECT 172.950 94.050 175.050 96.150 ;
        RECT 175.950 94.050 178.050 96.150 ;
        RECT 178.950 95.850 181.050 97.950 ;
        RECT 182.100 96.150 183.900 97.950 ;
        RECT 179.100 94.050 180.900 95.850 ;
        RECT 181.950 94.050 184.050 96.150 ;
        RECT 185.700 94.950 186.900 101.400 ;
        RECT 194.400 96.150 195.600 104.400 ;
        RECT 200.550 102.300 202.350 107.250 ;
        RECT 203.550 103.200 205.350 107.250 ;
        RECT 206.550 102.300 208.350 107.250 ;
        RECT 200.550 100.950 208.350 102.300 ;
        RECT 209.550 101.400 211.350 107.250 ;
        RECT 215.550 102.300 217.350 107.250 ;
        RECT 218.550 103.200 220.350 107.250 ;
        RECT 221.550 102.300 223.350 107.250 ;
        RECT 209.550 99.300 210.750 101.400 ;
        RECT 215.550 100.950 223.350 102.300 ;
        RECT 224.550 101.400 226.350 107.250 ;
        RECT 233.700 104.400 235.500 107.250 ;
        RECT 237.000 103.050 238.800 107.250 ;
        RECT 233.100 101.400 238.800 103.050 ;
        RECT 241.200 101.400 243.000 107.250 ;
        RECT 246.000 101.400 247.800 107.250 ;
        RECT 250.200 103.050 252.000 107.250 ;
        RECT 253.500 104.400 255.300 107.250 ;
        RECT 250.200 101.400 255.900 103.050 ;
        RECT 224.550 99.300 225.750 101.400 ;
        RECT 207.000 98.250 210.750 99.300 ;
        RECT 222.000 98.250 225.750 99.300 ;
        RECT 184.950 92.850 187.050 94.950 ;
        RECT 193.950 94.050 196.050 96.150 ;
        RECT 196.950 95.850 199.050 97.950 ;
        RECT 203.100 96.150 204.900 97.950 ;
        RECT 197.100 94.050 198.900 95.850 ;
        RECT 132.150 87.600 133.350 92.850 ;
        RECT 137.100 91.050 138.900 92.850 ;
        RECT 142.950 87.600 144.150 92.850 ;
        RECT 145.950 89.850 148.050 91.950 ;
        RECT 154.950 89.850 157.050 91.950 ;
        RECT 145.950 88.050 147.750 89.850 ;
        RECT 155.250 88.050 157.050 89.850 ;
        RECT 158.850 87.600 160.050 92.850 ;
        RECT 164.100 91.050 165.900 92.850 ;
        RECT 170.400 87.600 171.600 92.850 ;
        RECT 185.700 87.600 186.900 92.850 ;
        RECT 118.650 75.750 120.450 81.600 ;
        RECT 122.550 75.750 124.350 81.600 ;
        RECT 125.550 75.750 127.350 81.600 ;
        RECT 129.150 75.750 130.950 87.600 ;
        RECT 132.150 75.750 133.950 87.600 ;
        RECT 138.300 75.750 140.100 87.600 ;
        RECT 142.500 75.750 144.300 87.600 ;
        RECT 145.800 75.750 147.600 81.600 ;
        RECT 155.400 75.750 157.200 81.600 ;
        RECT 158.700 75.750 160.500 87.600 ;
        RECT 162.900 75.750 164.700 87.600 ;
        RECT 169.650 75.750 171.450 87.600 ;
        RECT 172.650 75.750 174.450 87.600 ;
        RECT 176.550 86.700 184.350 87.600 ;
        RECT 176.550 75.750 178.350 86.700 ;
        RECT 179.550 75.750 181.350 85.800 ;
        RECT 182.550 75.750 184.350 86.700 ;
        RECT 185.550 75.750 187.350 87.600 ;
        RECT 194.400 81.600 195.600 94.050 ;
        RECT 199.950 92.850 202.050 94.950 ;
        RECT 202.950 94.050 205.050 96.150 ;
        RECT 206.850 94.950 208.050 98.250 ;
        RECT 218.100 96.150 219.900 97.950 ;
        RECT 205.950 92.850 208.050 94.950 ;
        RECT 214.950 92.850 217.050 94.950 ;
        RECT 217.950 94.050 220.050 96.150 ;
        RECT 221.850 94.950 223.050 98.250 ;
        RECT 233.100 94.950 234.300 101.400 ;
        RECT 236.100 96.150 237.900 97.950 ;
        RECT 220.950 92.850 223.050 94.950 ;
        RECT 232.950 92.850 235.050 94.950 ;
        RECT 235.950 94.050 238.050 96.150 ;
        RECT 238.950 95.850 241.050 97.950 ;
        RECT 242.100 96.150 243.900 97.950 ;
        RECT 245.100 96.150 246.900 97.950 ;
        RECT 239.100 94.050 240.900 95.850 ;
        RECT 241.950 94.050 244.050 96.150 ;
        RECT 244.950 94.050 247.050 96.150 ;
        RECT 247.950 95.850 250.050 97.950 ;
        RECT 251.100 96.150 252.900 97.950 ;
        RECT 248.100 94.050 249.900 95.850 ;
        RECT 250.950 94.050 253.050 96.150 ;
        RECT 254.700 94.950 255.900 101.400 ;
        RECT 260.700 98.400 262.500 107.250 ;
        RECT 266.100 99.000 267.900 107.250 ;
        RECT 275.550 102.300 277.350 107.250 ;
        RECT 278.550 103.200 280.350 107.250 ;
        RECT 281.550 102.300 283.350 107.250 ;
        RECT 275.550 100.950 283.350 102.300 ;
        RECT 284.550 101.400 286.350 107.250 ;
        RECT 293.700 104.400 295.500 107.250 ;
        RECT 297.000 103.050 298.800 107.250 ;
        RECT 293.100 101.400 298.800 103.050 ;
        RECT 301.200 101.400 303.000 107.250 ;
        RECT 305.550 102.300 307.350 107.250 ;
        RECT 308.550 103.200 310.350 107.250 ;
        RECT 311.550 102.300 313.350 107.250 ;
        RECT 284.550 99.300 285.750 101.400 ;
        RECT 266.100 97.350 270.600 99.000 ;
        RECT 282.000 98.250 285.750 99.300 ;
        RECT 253.950 92.850 256.050 94.950 ;
        RECT 269.400 93.150 270.600 97.350 ;
        RECT 278.100 96.150 279.900 97.950 ;
        RECT 200.100 91.050 201.900 92.850 ;
        RECT 205.950 87.600 207.150 92.850 ;
        RECT 208.950 89.850 211.050 91.950 ;
        RECT 215.100 91.050 216.900 92.850 ;
        RECT 208.950 88.050 210.750 89.850 ;
        RECT 220.950 87.600 222.150 92.850 ;
        RECT 223.950 89.850 226.050 91.950 ;
        RECT 223.950 88.050 225.750 89.850 ;
        RECT 233.100 87.600 234.300 92.850 ;
        RECT 254.700 87.600 255.900 92.850 ;
        RECT 259.950 89.850 262.050 91.950 ;
        RECT 265.950 89.850 268.050 91.950 ;
        RECT 268.950 91.050 271.050 93.150 ;
        RECT 274.950 92.850 277.050 94.950 ;
        RECT 277.950 94.050 280.050 96.150 ;
        RECT 281.850 94.950 283.050 98.250 ;
        RECT 283.950 96.450 286.050 97.050 ;
        RECT 283.950 95.550 288.450 96.450 ;
        RECT 283.950 94.950 286.050 95.550 ;
        RECT 280.950 92.850 283.050 94.950 ;
        RECT 275.100 91.050 276.900 92.850 ;
        RECT 260.100 88.050 261.900 89.850 ;
        RECT 193.650 75.750 195.450 81.600 ;
        RECT 196.650 75.750 198.450 81.600 ;
        RECT 201.300 75.750 203.100 87.600 ;
        RECT 205.500 75.750 207.300 87.600 ;
        RECT 208.800 75.750 210.600 81.600 ;
        RECT 216.300 75.750 218.100 87.600 ;
        RECT 220.500 75.750 222.300 87.600 ;
        RECT 223.800 75.750 225.600 81.600 ;
        RECT 232.650 75.750 234.450 87.600 ;
        RECT 235.650 86.700 243.450 87.600 ;
        RECT 235.650 75.750 237.450 86.700 ;
        RECT 238.650 75.750 240.450 85.800 ;
        RECT 241.650 75.750 243.450 86.700 ;
        RECT 245.550 86.700 253.350 87.600 ;
        RECT 245.550 75.750 247.350 86.700 ;
        RECT 248.550 75.750 250.350 85.800 ;
        RECT 251.550 75.750 253.350 86.700 ;
        RECT 254.550 75.750 256.350 87.600 ;
        RECT 262.950 86.850 265.050 88.950 ;
        RECT 266.250 88.050 268.050 89.850 ;
        RECT 263.100 85.050 264.900 86.850 ;
        RECT 269.700 82.800 270.750 91.050 ;
        RECT 280.950 87.600 282.150 92.850 ;
        RECT 283.950 89.850 286.050 91.950 ;
        RECT 283.950 88.050 285.750 89.850 ;
        RECT 263.700 81.900 270.750 82.800 ;
        RECT 263.700 81.600 265.350 81.900 ;
        RECT 260.550 75.750 262.350 81.600 ;
        RECT 263.550 75.750 265.350 81.600 ;
        RECT 269.550 81.600 270.750 81.900 ;
        RECT 266.550 75.750 268.350 81.000 ;
        RECT 269.550 75.750 271.350 81.600 ;
        RECT 276.300 75.750 278.100 87.600 ;
        RECT 280.500 75.750 282.300 87.600 ;
        RECT 283.950 84.450 286.050 85.050 ;
        RECT 287.550 84.450 288.450 95.550 ;
        RECT 293.100 94.950 294.300 101.400 ;
        RECT 305.550 100.950 313.350 102.300 ;
        RECT 314.550 101.400 316.350 107.250 ;
        RECT 322.950 102.450 325.050 103.050 ;
        RECT 320.550 101.550 325.050 102.450 ;
        RECT 314.550 99.300 315.750 101.400 ;
        RECT 320.550 99.450 321.450 101.550 ;
        RECT 322.950 100.950 325.050 101.550 ;
        RECT 312.000 98.250 315.750 99.300 ;
        RECT 317.550 98.550 321.450 99.450 ;
        RECT 326.100 99.000 327.900 107.250 ;
        RECT 296.100 96.150 297.900 97.950 ;
        RECT 292.950 92.850 295.050 94.950 ;
        RECT 295.950 94.050 298.050 96.150 ;
        RECT 298.950 95.850 301.050 97.950 ;
        RECT 302.100 96.150 303.900 97.950 ;
        RECT 308.100 96.150 309.900 97.950 ;
        RECT 299.100 94.050 300.900 95.850 ;
        RECT 301.950 94.050 304.050 96.150 ;
        RECT 304.950 92.850 307.050 94.950 ;
        RECT 307.950 94.050 310.050 96.150 ;
        RECT 311.850 94.950 313.050 98.250 ;
        RECT 310.950 92.850 313.050 94.950 ;
        RECT 293.100 87.600 294.300 92.850 ;
        RECT 305.100 91.050 306.900 92.850 ;
        RECT 310.950 87.600 312.150 92.850 ;
        RECT 313.950 89.850 316.050 91.950 ;
        RECT 313.950 88.050 315.750 89.850 ;
        RECT 317.550 88.050 318.450 98.550 ;
        RECT 323.400 97.350 327.900 99.000 ;
        RECT 331.500 98.400 333.300 107.250 ;
        RECT 337.650 101.400 339.450 107.250 ;
        RECT 338.250 99.300 339.450 101.400 ;
        RECT 340.650 102.300 342.450 107.250 ;
        RECT 343.650 103.200 345.450 107.250 ;
        RECT 346.650 102.300 348.450 107.250 ;
        RECT 340.650 100.950 348.450 102.300 ;
        RECT 350.550 102.300 352.350 107.250 ;
        RECT 353.550 103.200 355.350 107.250 ;
        RECT 356.550 102.300 358.350 107.250 ;
        RECT 350.550 100.950 358.350 102.300 ;
        RECT 359.550 101.400 361.350 107.250 ;
        RECT 359.550 99.300 360.750 101.400 ;
        RECT 338.250 98.250 342.000 99.300 ;
        RECT 357.000 98.250 360.750 99.300 ;
        RECT 365.700 98.400 367.500 107.250 ;
        RECT 371.100 99.000 372.900 107.250 ;
        RECT 323.400 93.150 324.600 97.350 ;
        RECT 340.950 94.950 342.150 98.250 ;
        RECT 344.100 96.150 345.900 97.950 ;
        RECT 353.100 96.150 354.900 97.950 ;
        RECT 322.950 91.050 325.050 93.150 ;
        RECT 340.950 92.850 343.050 94.950 ;
        RECT 343.950 94.050 346.050 96.150 ;
        RECT 346.950 92.850 349.050 94.950 ;
        RECT 349.950 92.850 352.050 94.950 ;
        RECT 352.950 94.050 355.050 96.150 ;
        RECT 356.850 94.950 358.050 98.250 ;
        RECT 371.100 97.350 375.600 99.000 ;
        RECT 380.700 98.400 382.500 107.250 ;
        RECT 386.100 99.000 387.900 107.250 ;
        RECT 397.650 104.400 399.450 107.250 ;
        RECT 400.650 104.400 402.450 107.250 ;
        RECT 386.100 97.350 390.600 99.000 ;
        RECT 355.950 92.850 358.050 94.950 ;
        RECT 374.400 93.150 375.600 97.350 ;
        RECT 389.400 93.150 390.600 97.350 ;
        RECT 398.400 96.150 399.600 104.400 ;
        RECT 404.700 98.400 406.500 107.250 ;
        RECT 410.100 99.000 411.900 107.250 ;
        RECT 420.150 101.400 421.950 107.250 ;
        RECT 423.150 104.400 424.950 107.250 ;
        RECT 427.950 105.300 429.750 107.250 ;
        RECT 426.000 104.400 429.750 105.300 ;
        RECT 432.450 104.400 434.250 107.250 ;
        RECT 435.750 104.400 437.550 107.250 ;
        RECT 439.650 104.400 441.450 107.250 ;
        RECT 443.850 104.400 445.650 107.250 ;
        RECT 448.350 104.400 450.150 107.250 ;
        RECT 426.000 103.500 427.050 104.400 ;
        RECT 424.950 101.400 427.050 103.500 ;
        RECT 435.750 102.600 436.800 104.400 ;
        RECT 397.950 94.050 400.050 96.150 ;
        RECT 400.950 95.850 403.050 97.950 ;
        RECT 410.100 97.350 414.600 99.000 ;
        RECT 401.100 94.050 402.900 95.850 ;
        RECT 283.950 83.550 288.450 84.450 ;
        RECT 283.950 82.950 286.050 83.550 ;
        RECT 283.800 75.750 285.600 81.600 ;
        RECT 292.650 75.750 294.450 87.600 ;
        RECT 295.650 86.700 303.450 87.600 ;
        RECT 295.650 75.750 297.450 86.700 ;
        RECT 298.650 75.750 300.450 85.800 ;
        RECT 301.650 75.750 303.450 86.700 ;
        RECT 306.300 75.750 308.100 87.600 ;
        RECT 310.500 75.750 312.300 87.600 ;
        RECT 316.950 85.950 319.050 88.050 ;
        RECT 323.250 82.800 324.300 91.050 ;
        RECT 325.950 89.850 328.050 91.950 ;
        RECT 331.950 89.850 334.050 91.950 ;
        RECT 337.950 89.850 340.050 91.950 ;
        RECT 325.950 88.050 327.750 89.850 ;
        RECT 328.950 86.850 331.050 88.950 ;
        RECT 332.100 88.050 333.900 89.850 ;
        RECT 338.250 88.050 340.050 89.850 ;
        RECT 341.850 87.600 343.050 92.850 ;
        RECT 347.100 91.050 348.900 92.850 ;
        RECT 350.100 91.050 351.900 92.850 ;
        RECT 355.950 87.600 357.150 92.850 ;
        RECT 358.950 89.850 361.050 91.950 ;
        RECT 364.950 89.850 367.050 91.950 ;
        RECT 370.950 89.850 373.050 91.950 ;
        RECT 373.950 91.050 376.050 93.150 ;
        RECT 358.950 88.050 360.750 89.850 ;
        RECT 365.100 88.050 366.900 89.850 ;
        RECT 329.100 85.050 330.900 86.850 ;
        RECT 323.250 81.900 330.300 82.800 ;
        RECT 323.250 81.600 324.450 81.900 ;
        RECT 313.800 75.750 315.600 81.600 ;
        RECT 322.650 75.750 324.450 81.600 ;
        RECT 328.650 81.600 330.300 81.900 ;
        RECT 325.650 75.750 327.450 81.000 ;
        RECT 328.650 75.750 330.450 81.600 ;
        RECT 331.650 75.750 333.450 81.600 ;
        RECT 338.400 75.750 340.200 81.600 ;
        RECT 341.700 75.750 343.500 87.600 ;
        RECT 345.900 75.750 347.700 87.600 ;
        RECT 351.300 75.750 353.100 87.600 ;
        RECT 355.500 75.750 357.300 87.600 ;
        RECT 367.950 86.850 370.050 88.950 ;
        RECT 371.250 88.050 373.050 89.850 ;
        RECT 368.100 85.050 369.900 86.850 ;
        RECT 374.700 82.800 375.750 91.050 ;
        RECT 379.950 89.850 382.050 91.950 ;
        RECT 385.950 89.850 388.050 91.950 ;
        RECT 388.950 91.050 391.050 93.150 ;
        RECT 380.100 88.050 381.900 89.850 ;
        RECT 382.950 86.850 385.050 88.950 ;
        RECT 386.250 88.050 388.050 89.850 ;
        RECT 383.100 85.050 384.900 86.850 ;
        RECT 389.700 82.800 390.750 91.050 ;
        RECT 368.700 81.900 375.750 82.800 ;
        RECT 368.700 81.600 370.350 81.900 ;
        RECT 358.800 75.750 360.600 81.600 ;
        RECT 365.550 75.750 367.350 81.600 ;
        RECT 368.550 75.750 370.350 81.600 ;
        RECT 374.550 81.600 375.750 81.900 ;
        RECT 383.700 81.900 390.750 82.800 ;
        RECT 383.700 81.600 385.350 81.900 ;
        RECT 371.550 75.750 373.350 81.000 ;
        RECT 374.550 75.750 376.350 81.600 ;
        RECT 380.550 75.750 382.350 81.600 ;
        RECT 383.550 75.750 385.350 81.600 ;
        RECT 389.550 81.600 390.750 81.900 ;
        RECT 398.400 81.600 399.600 94.050 ;
        RECT 413.400 93.150 414.600 97.350 ;
        RECT 403.950 89.850 406.050 91.950 ;
        RECT 409.950 89.850 412.050 91.950 ;
        RECT 412.950 91.050 415.050 93.150 ;
        RECT 404.100 88.050 405.900 89.850 ;
        RECT 406.950 86.850 409.050 88.950 ;
        RECT 410.250 88.050 412.050 89.850 ;
        RECT 407.100 85.050 408.900 86.850 ;
        RECT 413.700 82.800 414.750 91.050 ;
        RECT 407.700 81.900 414.750 82.800 ;
        RECT 407.700 81.600 409.350 81.900 ;
        RECT 386.550 75.750 388.350 81.000 ;
        RECT 389.550 75.750 391.350 81.600 ;
        RECT 397.650 75.750 399.450 81.600 ;
        RECT 400.650 75.750 402.450 81.600 ;
        RECT 404.550 75.750 406.350 81.600 ;
        RECT 407.550 75.750 409.350 81.600 ;
        RECT 413.550 81.600 414.750 81.900 ;
        RECT 420.150 88.800 421.050 101.400 ;
        RECT 428.550 100.800 430.350 102.600 ;
        RECT 431.850 101.550 436.800 102.600 ;
        RECT 444.300 103.500 445.350 104.400 ;
        RECT 444.300 102.300 448.050 103.500 ;
        RECT 431.850 100.800 433.650 101.550 ;
        RECT 428.850 99.900 429.900 100.800 ;
        RECT 439.050 100.200 440.850 102.000 ;
        RECT 445.950 101.400 448.050 102.300 ;
        RECT 451.650 101.400 453.450 107.250 ;
        RECT 439.050 99.900 439.950 100.200 ;
        RECT 428.850 99.000 439.950 99.900 ;
        RECT 452.250 99.150 453.450 101.400 ;
        RECT 455.550 102.300 457.350 107.250 ;
        RECT 458.550 103.200 460.350 107.250 ;
        RECT 461.550 102.300 463.350 107.250 ;
        RECT 455.550 100.950 463.350 102.300 ;
        RECT 464.550 101.400 466.350 107.250 ;
        RECT 470.550 104.400 472.350 107.250 ;
        RECT 473.550 104.400 475.350 107.250 ;
        RECT 479.550 104.400 481.350 107.250 ;
        RECT 482.550 104.400 484.350 107.250 ;
        RECT 464.550 99.300 465.750 101.400 ;
        RECT 428.850 97.800 429.900 99.000 ;
        RECT 423.000 96.600 429.900 97.800 ;
        RECT 423.000 95.850 423.900 96.600 ;
        RECT 428.100 96.000 429.900 96.600 ;
        RECT 422.100 94.050 423.900 95.850 ;
        RECT 425.100 94.950 426.900 95.700 ;
        RECT 439.050 94.950 439.950 99.000 ;
        RECT 448.950 97.050 453.450 99.150 ;
        RECT 462.000 98.250 465.750 99.300 ;
        RECT 447.150 95.250 451.050 97.050 ;
        RECT 448.950 94.950 451.050 95.250 ;
        RECT 425.100 93.900 433.050 94.950 ;
        RECT 430.950 92.850 433.050 93.900 ;
        RECT 436.950 92.850 439.950 94.950 ;
        RECT 429.450 89.100 431.250 89.400 ;
        RECT 429.450 88.800 437.850 89.100 ;
        RECT 420.150 88.200 437.850 88.800 ;
        RECT 420.150 87.600 431.250 88.200 ;
        RECT 410.550 75.750 412.350 81.000 ;
        RECT 413.550 75.750 415.350 81.600 ;
        RECT 420.150 75.750 421.950 87.600 ;
        RECT 434.250 86.700 436.050 87.300 ;
        RECT 428.550 85.500 436.050 86.700 ;
        RECT 436.950 86.100 437.850 88.200 ;
        RECT 439.050 88.200 439.950 92.850 ;
        RECT 449.250 89.400 451.050 91.200 ;
        RECT 445.950 88.200 450.150 89.400 ;
        RECT 439.050 87.300 445.050 88.200 ;
        RECT 445.950 87.300 448.050 88.200 ;
        RECT 452.250 87.600 453.450 97.050 ;
        RECT 458.100 96.150 459.900 97.950 ;
        RECT 454.950 92.850 457.050 94.950 ;
        RECT 457.950 94.050 460.050 96.150 ;
        RECT 461.850 94.950 463.050 98.250 ;
        RECT 469.950 95.850 472.050 97.950 ;
        RECT 473.400 96.150 474.600 104.400 ;
        RECT 460.950 92.850 463.050 94.950 ;
        RECT 470.100 94.050 471.900 95.850 ;
        RECT 472.950 94.050 475.050 96.150 ;
        RECT 478.950 95.850 481.050 97.950 ;
        RECT 482.400 96.150 483.600 104.400 ;
        RECT 488.700 98.400 490.500 107.250 ;
        RECT 494.100 99.000 495.900 107.250 ;
        RECT 505.650 104.400 507.450 107.250 ;
        RECT 508.650 104.400 510.450 107.250 ;
        RECT 494.100 97.350 498.600 99.000 ;
        RECT 479.100 94.050 480.900 95.850 ;
        RECT 481.950 94.050 484.050 96.150 ;
        RECT 455.100 91.050 456.900 92.850 ;
        RECT 460.950 87.600 462.150 92.850 ;
        RECT 463.950 89.850 466.050 91.950 ;
        RECT 463.950 88.050 465.750 89.850 ;
        RECT 444.150 86.400 445.050 87.300 ;
        RECT 441.450 86.100 443.250 86.400 ;
        RECT 428.550 84.600 429.750 85.500 ;
        RECT 436.950 85.200 443.250 86.100 ;
        RECT 441.450 84.600 443.250 85.200 ;
        RECT 444.150 84.600 446.850 86.400 ;
        RECT 424.950 82.500 429.750 84.600 ;
        RECT 432.150 82.500 439.050 84.300 ;
        RECT 428.550 81.600 429.750 82.500 ;
        RECT 423.150 75.750 424.950 81.600 ;
        RECT 428.250 75.750 430.050 81.600 ;
        RECT 433.050 75.750 434.850 81.600 ;
        RECT 436.050 75.750 437.850 82.500 ;
        RECT 444.150 81.600 448.050 83.700 ;
        RECT 439.950 75.750 441.750 81.600 ;
        RECT 444.150 75.750 445.950 81.600 ;
        RECT 448.650 75.750 450.450 78.600 ;
        RECT 451.650 75.750 453.450 87.600 ;
        RECT 456.300 75.750 458.100 87.600 ;
        RECT 460.500 75.750 462.300 87.600 ;
        RECT 473.400 81.600 474.600 94.050 ;
        RECT 482.400 81.600 483.600 94.050 ;
        RECT 497.400 93.150 498.600 97.350 ;
        RECT 506.400 96.150 507.600 104.400 ;
        RECT 515.850 100.200 517.650 107.250 ;
        RECT 520.350 101.400 522.150 107.250 ;
        RECT 526.650 101.400 528.450 107.250 ;
        RECT 515.850 99.300 519.450 100.200 ;
        RECT 505.950 94.050 508.050 96.150 ;
        RECT 508.950 95.850 511.050 97.950 ;
        RECT 509.100 94.050 510.900 95.850 ;
        RECT 487.950 89.850 490.050 91.950 ;
        RECT 493.950 89.850 496.050 91.950 ;
        RECT 496.950 91.050 499.050 93.150 ;
        RECT 488.100 88.050 489.900 89.850 ;
        RECT 490.950 86.850 493.050 88.950 ;
        RECT 494.250 88.050 496.050 89.850 ;
        RECT 491.100 85.050 492.900 86.850 ;
        RECT 497.700 82.800 498.750 91.050 ;
        RECT 491.700 81.900 498.750 82.800 ;
        RECT 491.700 81.600 493.350 81.900 ;
        RECT 463.800 75.750 465.600 81.600 ;
        RECT 470.550 75.750 472.350 81.600 ;
        RECT 473.550 75.750 475.350 81.600 ;
        RECT 479.550 75.750 481.350 81.600 ;
        RECT 482.550 75.750 484.350 81.600 ;
        RECT 488.550 75.750 490.350 81.600 ;
        RECT 491.550 75.750 493.350 81.600 ;
        RECT 497.550 81.600 498.750 81.900 ;
        RECT 506.400 81.600 507.600 94.050 ;
        RECT 515.100 93.150 516.900 94.950 ;
        RECT 514.950 91.050 517.050 93.150 ;
        RECT 518.250 91.950 519.450 99.300 ;
        RECT 527.250 99.300 528.450 101.400 ;
        RECT 529.650 102.300 531.450 107.250 ;
        RECT 532.650 103.200 534.450 107.250 ;
        RECT 535.650 102.300 537.450 107.250 ;
        RECT 529.650 100.950 537.450 102.300 ;
        RECT 540.150 101.400 541.950 107.250 ;
        RECT 543.150 104.400 544.950 107.250 ;
        RECT 547.950 105.300 549.750 107.250 ;
        RECT 546.000 104.400 549.750 105.300 ;
        RECT 552.450 104.400 554.250 107.250 ;
        RECT 555.750 104.400 557.550 107.250 ;
        RECT 559.650 104.400 561.450 107.250 ;
        RECT 563.850 104.400 565.650 107.250 ;
        RECT 568.350 104.400 570.150 107.250 ;
        RECT 546.000 103.500 547.050 104.400 ;
        RECT 544.950 101.400 547.050 103.500 ;
        RECT 555.750 102.600 556.800 104.400 ;
        RECT 527.250 98.250 531.000 99.300 ;
        RECT 529.950 94.950 531.150 98.250 ;
        RECT 533.100 96.150 534.900 97.950 ;
        RECT 521.100 93.150 522.900 94.950 ;
        RECT 517.950 89.850 520.050 91.950 ;
        RECT 520.950 91.050 523.050 93.150 ;
        RECT 529.950 92.850 532.050 94.950 ;
        RECT 532.950 94.050 535.050 96.150 ;
        RECT 535.950 92.850 538.050 94.950 ;
        RECT 526.950 89.850 529.050 91.950 ;
        RECT 518.250 81.600 519.450 89.850 ;
        RECT 527.250 88.050 529.050 89.850 ;
        RECT 530.850 87.600 532.050 92.850 ;
        RECT 536.100 91.050 537.900 92.850 ;
        RECT 540.150 88.800 541.050 101.400 ;
        RECT 548.550 100.800 550.350 102.600 ;
        RECT 551.850 101.550 556.800 102.600 ;
        RECT 564.300 103.500 565.350 104.400 ;
        RECT 564.300 102.300 568.050 103.500 ;
        RECT 551.850 100.800 553.650 101.550 ;
        RECT 548.850 99.900 549.900 100.800 ;
        RECT 559.050 100.200 560.850 102.000 ;
        RECT 565.950 101.400 568.050 102.300 ;
        RECT 571.650 101.400 573.450 107.250 ;
        RECT 559.050 99.900 559.950 100.200 ;
        RECT 548.850 99.000 559.950 99.900 ;
        RECT 572.250 99.150 573.450 101.400 ;
        RECT 575.550 102.300 577.350 107.250 ;
        RECT 578.550 103.200 580.350 107.250 ;
        RECT 581.550 102.300 583.350 107.250 ;
        RECT 575.550 100.950 583.350 102.300 ;
        RECT 584.550 101.400 586.350 107.250 ;
        RECT 584.550 99.300 585.750 101.400 ;
        RECT 593.850 100.200 595.650 107.250 ;
        RECT 598.350 101.400 600.150 107.250 ;
        RECT 602.550 101.400 604.350 107.250 ;
        RECT 605.850 104.400 607.650 107.250 ;
        RECT 610.350 104.400 612.150 107.250 ;
        RECT 614.550 104.400 616.350 107.250 ;
        RECT 618.450 104.400 620.250 107.250 ;
        RECT 621.750 104.400 623.550 107.250 ;
        RECT 626.250 105.300 628.050 107.250 ;
        RECT 626.250 104.400 630.000 105.300 ;
        RECT 631.050 104.400 632.850 107.250 ;
        RECT 610.650 103.500 611.700 104.400 ;
        RECT 607.950 102.300 611.700 103.500 ;
        RECT 619.200 102.600 620.250 104.400 ;
        RECT 628.950 103.500 630.000 104.400 ;
        RECT 607.950 101.400 610.050 102.300 ;
        RECT 593.850 99.300 597.450 100.200 ;
        RECT 548.850 97.800 549.900 99.000 ;
        RECT 543.000 96.600 549.900 97.800 ;
        RECT 543.000 95.850 543.900 96.600 ;
        RECT 548.100 96.000 549.900 96.600 ;
        RECT 542.100 94.050 543.900 95.850 ;
        RECT 545.100 94.950 546.900 95.700 ;
        RECT 559.050 94.950 559.950 99.000 ;
        RECT 568.950 97.050 573.450 99.150 ;
        RECT 582.000 98.250 585.750 99.300 ;
        RECT 567.150 95.250 571.050 97.050 ;
        RECT 568.950 94.950 571.050 95.250 ;
        RECT 545.100 93.900 553.050 94.950 ;
        RECT 550.950 92.850 553.050 93.900 ;
        RECT 556.950 92.850 559.950 94.950 ;
        RECT 549.450 89.100 551.250 89.400 ;
        RECT 549.450 88.800 557.850 89.100 ;
        RECT 540.150 88.200 557.850 88.800 ;
        RECT 540.150 87.600 551.250 88.200 ;
        RECT 494.550 75.750 496.350 81.000 ;
        RECT 497.550 75.750 499.350 81.600 ;
        RECT 505.650 75.750 507.450 81.600 ;
        RECT 508.650 75.750 510.450 81.600 ;
        RECT 514.650 75.750 516.450 81.600 ;
        RECT 517.650 75.750 519.450 81.600 ;
        RECT 520.650 75.750 522.450 81.600 ;
        RECT 527.400 75.750 529.200 81.600 ;
        RECT 530.700 75.750 532.500 87.600 ;
        RECT 534.900 75.750 536.700 87.600 ;
        RECT 540.150 75.750 541.950 87.600 ;
        RECT 554.250 86.700 556.050 87.300 ;
        RECT 548.550 85.500 556.050 86.700 ;
        RECT 556.950 86.100 557.850 88.200 ;
        RECT 559.050 88.200 559.950 92.850 ;
        RECT 569.250 89.400 571.050 91.200 ;
        RECT 565.950 88.200 570.150 89.400 ;
        RECT 559.050 87.300 565.050 88.200 ;
        RECT 565.950 87.300 568.050 88.200 ;
        RECT 572.250 87.600 573.450 97.050 ;
        RECT 578.100 96.150 579.900 97.950 ;
        RECT 574.950 92.850 577.050 94.950 ;
        RECT 577.950 94.050 580.050 96.150 ;
        RECT 581.850 94.950 583.050 98.250 ;
        RECT 580.950 92.850 583.050 94.950 ;
        RECT 593.100 93.150 594.900 94.950 ;
        RECT 575.100 91.050 576.900 92.850 ;
        RECT 580.950 87.600 582.150 92.850 ;
        RECT 583.950 89.850 586.050 91.950 ;
        RECT 592.950 91.050 595.050 93.150 ;
        RECT 596.250 91.950 597.450 99.300 ;
        RECT 602.550 99.150 603.750 101.400 ;
        RECT 615.150 100.200 616.950 102.000 ;
        RECT 619.200 101.550 624.150 102.600 ;
        RECT 622.350 100.800 624.150 101.550 ;
        RECT 625.650 100.800 627.450 102.600 ;
        RECT 628.950 101.400 631.050 103.500 ;
        RECT 634.050 101.400 635.850 107.250 ;
        RECT 638.850 101.400 640.650 107.250 ;
        RECT 616.050 99.900 616.950 100.200 ;
        RECT 626.100 99.900 627.150 100.800 ;
        RECT 602.550 97.050 607.050 99.150 ;
        RECT 616.050 99.000 627.150 99.900 ;
        RECT 599.100 93.150 600.900 94.950 ;
        RECT 595.950 89.850 598.050 91.950 ;
        RECT 598.950 91.050 601.050 93.150 ;
        RECT 583.950 88.050 585.750 89.850 ;
        RECT 564.150 86.400 565.050 87.300 ;
        RECT 561.450 86.100 563.250 86.400 ;
        RECT 548.550 84.600 549.750 85.500 ;
        RECT 556.950 85.200 563.250 86.100 ;
        RECT 561.450 84.600 563.250 85.200 ;
        RECT 564.150 84.600 566.850 86.400 ;
        RECT 544.950 82.500 549.750 84.600 ;
        RECT 552.150 82.500 559.050 84.300 ;
        RECT 548.550 81.600 549.750 82.500 ;
        RECT 543.150 75.750 544.950 81.600 ;
        RECT 548.250 75.750 550.050 81.600 ;
        RECT 553.050 75.750 554.850 81.600 ;
        RECT 556.050 75.750 557.850 82.500 ;
        RECT 564.150 81.600 568.050 83.700 ;
        RECT 559.950 75.750 561.750 81.600 ;
        RECT 564.150 75.750 565.950 81.600 ;
        RECT 568.650 75.750 570.450 78.600 ;
        RECT 571.650 75.750 573.450 87.600 ;
        RECT 576.300 75.750 578.100 87.600 ;
        RECT 580.500 75.750 582.300 87.600 ;
        RECT 596.250 81.600 597.450 89.850 ;
        RECT 602.550 87.600 603.750 97.050 ;
        RECT 604.950 95.250 608.850 97.050 ;
        RECT 604.950 94.950 607.050 95.250 ;
        RECT 616.050 94.950 616.950 99.000 ;
        RECT 626.100 97.800 627.150 99.000 ;
        RECT 626.100 96.600 633.000 97.800 ;
        RECT 626.100 96.000 627.900 96.600 ;
        RECT 632.100 95.850 633.000 96.600 ;
        RECT 629.100 94.950 630.900 95.700 ;
        RECT 616.050 92.850 619.050 94.950 ;
        RECT 622.950 93.900 630.900 94.950 ;
        RECT 632.100 94.050 633.900 95.850 ;
        RECT 622.950 92.850 625.050 93.900 ;
        RECT 604.950 89.400 606.750 91.200 ;
        RECT 605.850 88.200 610.050 89.400 ;
        RECT 616.050 88.200 616.950 92.850 ;
        RECT 624.750 89.100 626.550 89.400 ;
        RECT 583.800 75.750 585.600 81.600 ;
        RECT 592.650 75.750 594.450 81.600 ;
        RECT 595.650 75.750 597.450 81.600 ;
        RECT 598.650 75.750 600.450 81.600 ;
        RECT 602.550 75.750 604.350 87.600 ;
        RECT 607.950 87.300 610.050 88.200 ;
        RECT 610.950 87.300 616.950 88.200 ;
        RECT 618.150 88.800 626.550 89.100 ;
        RECT 634.950 88.800 635.850 101.400 ;
        RECT 643.350 100.200 645.150 107.250 ;
        RECT 650.850 101.400 652.650 107.250 ;
        RECT 655.350 100.200 657.150 107.250 ;
        RECT 664.650 101.400 666.450 107.250 ;
        RECT 641.550 99.300 645.150 100.200 ;
        RECT 653.550 99.300 657.150 100.200 ;
        RECT 665.250 99.300 666.450 101.400 ;
        RECT 667.650 102.300 669.450 107.250 ;
        RECT 670.650 103.200 672.450 107.250 ;
        RECT 673.650 102.300 675.450 107.250 ;
        RECT 667.650 100.950 675.450 102.300 ;
        RECT 678.150 101.400 679.950 107.250 ;
        RECT 681.150 104.400 682.950 107.250 ;
        RECT 685.950 105.300 687.750 107.250 ;
        RECT 684.000 104.400 687.750 105.300 ;
        RECT 690.450 104.400 692.250 107.250 ;
        RECT 693.750 104.400 695.550 107.250 ;
        RECT 697.650 104.400 699.450 107.250 ;
        RECT 701.850 104.400 703.650 107.250 ;
        RECT 706.350 104.400 708.150 107.250 ;
        RECT 684.000 103.500 685.050 104.400 ;
        RECT 682.950 101.400 685.050 103.500 ;
        RECT 693.750 102.600 694.800 104.400 ;
        RECT 638.100 93.150 639.900 94.950 ;
        RECT 637.950 91.050 640.050 93.150 ;
        RECT 641.550 91.950 642.750 99.300 ;
        RECT 644.100 93.150 645.900 94.950 ;
        RECT 650.100 93.150 651.900 94.950 ;
        RECT 640.950 89.850 643.050 91.950 ;
        RECT 643.950 91.050 646.050 93.150 ;
        RECT 649.950 91.050 652.050 93.150 ;
        RECT 653.550 91.950 654.750 99.300 ;
        RECT 665.250 98.250 669.000 99.300 ;
        RECT 667.950 94.950 669.150 98.250 ;
        RECT 671.100 96.150 672.900 97.950 ;
        RECT 656.100 93.150 657.900 94.950 ;
        RECT 652.950 89.850 655.050 91.950 ;
        RECT 655.950 91.050 658.050 93.150 ;
        RECT 667.950 92.850 670.050 94.950 ;
        RECT 670.950 94.050 673.050 96.150 ;
        RECT 673.950 92.850 676.050 94.950 ;
        RECT 664.950 89.850 667.050 91.950 ;
        RECT 618.150 88.200 635.850 88.800 ;
        RECT 610.950 86.400 611.850 87.300 ;
        RECT 609.150 84.600 611.850 86.400 ;
        RECT 612.750 86.100 614.550 86.400 ;
        RECT 618.150 86.100 619.050 88.200 ;
        RECT 624.750 87.600 635.850 88.200 ;
        RECT 612.750 85.200 619.050 86.100 ;
        RECT 619.950 86.700 621.750 87.300 ;
        RECT 619.950 85.500 627.450 86.700 ;
        RECT 612.750 84.600 614.550 85.200 ;
        RECT 626.250 84.600 627.450 85.500 ;
        RECT 607.950 81.600 611.850 83.700 ;
        RECT 616.950 82.500 623.850 84.300 ;
        RECT 626.250 82.500 631.050 84.600 ;
        RECT 605.550 75.750 607.350 78.600 ;
        RECT 610.050 75.750 611.850 81.600 ;
        RECT 614.250 75.750 616.050 81.600 ;
        RECT 618.150 75.750 619.950 82.500 ;
        RECT 626.250 81.600 627.450 82.500 ;
        RECT 621.150 75.750 622.950 81.600 ;
        RECT 625.950 75.750 627.750 81.600 ;
        RECT 631.050 75.750 632.850 81.600 ;
        RECT 634.050 75.750 635.850 87.600 ;
        RECT 641.550 81.600 642.750 89.850 ;
        RECT 653.550 81.600 654.750 89.850 ;
        RECT 665.250 88.050 667.050 89.850 ;
        RECT 668.850 87.600 670.050 92.850 ;
        RECT 674.100 91.050 675.900 92.850 ;
        RECT 678.150 88.800 679.050 101.400 ;
        RECT 686.550 100.800 688.350 102.600 ;
        RECT 689.850 101.550 694.800 102.600 ;
        RECT 702.300 103.500 703.350 104.400 ;
        RECT 702.300 102.300 706.050 103.500 ;
        RECT 689.850 100.800 691.650 101.550 ;
        RECT 686.850 99.900 687.900 100.800 ;
        RECT 697.050 100.200 698.850 102.000 ;
        RECT 703.950 101.400 706.050 102.300 ;
        RECT 709.650 101.400 711.450 107.250 ;
        RECT 697.050 99.900 697.950 100.200 ;
        RECT 686.850 99.000 697.950 99.900 ;
        RECT 710.250 99.150 711.450 101.400 ;
        RECT 686.850 97.800 687.900 99.000 ;
        RECT 681.000 96.600 687.900 97.800 ;
        RECT 681.000 95.850 681.900 96.600 ;
        RECT 686.100 96.000 687.900 96.600 ;
        RECT 680.100 94.050 681.900 95.850 ;
        RECT 683.100 94.950 684.900 95.700 ;
        RECT 697.050 94.950 697.950 99.000 ;
        RECT 706.950 97.050 711.450 99.150 ;
        RECT 705.150 95.250 709.050 97.050 ;
        RECT 706.950 94.950 709.050 95.250 ;
        RECT 683.100 93.900 691.050 94.950 ;
        RECT 688.950 92.850 691.050 93.900 ;
        RECT 694.950 92.850 697.950 94.950 ;
        RECT 687.450 89.100 689.250 89.400 ;
        RECT 687.450 88.800 695.850 89.100 ;
        RECT 678.150 88.200 695.850 88.800 ;
        RECT 678.150 87.600 689.250 88.200 ;
        RECT 638.550 75.750 640.350 81.600 ;
        RECT 641.550 75.750 643.350 81.600 ;
        RECT 644.550 75.750 646.350 81.600 ;
        RECT 650.550 75.750 652.350 81.600 ;
        RECT 653.550 75.750 655.350 81.600 ;
        RECT 656.550 75.750 658.350 81.600 ;
        RECT 665.400 75.750 667.200 81.600 ;
        RECT 668.700 75.750 670.500 87.600 ;
        RECT 672.900 75.750 674.700 87.600 ;
        RECT 678.150 75.750 679.950 87.600 ;
        RECT 692.250 86.700 694.050 87.300 ;
        RECT 686.550 85.500 694.050 86.700 ;
        RECT 694.950 86.100 695.850 88.200 ;
        RECT 697.050 88.200 697.950 92.850 ;
        RECT 707.250 89.400 709.050 91.200 ;
        RECT 703.950 88.200 708.150 89.400 ;
        RECT 697.050 87.300 703.050 88.200 ;
        RECT 703.950 87.300 706.050 88.200 ;
        RECT 710.250 87.600 711.450 97.050 ;
        RECT 702.150 86.400 703.050 87.300 ;
        RECT 699.450 86.100 701.250 86.400 ;
        RECT 686.550 84.600 687.750 85.500 ;
        RECT 694.950 85.200 701.250 86.100 ;
        RECT 699.450 84.600 701.250 85.200 ;
        RECT 702.150 84.600 704.850 86.400 ;
        RECT 682.950 82.500 687.750 84.600 ;
        RECT 690.150 82.500 697.050 84.300 ;
        RECT 686.550 81.600 687.750 82.500 ;
        RECT 681.150 75.750 682.950 81.600 ;
        RECT 686.250 75.750 688.050 81.600 ;
        RECT 691.050 75.750 692.850 81.600 ;
        RECT 694.050 75.750 695.850 82.500 ;
        RECT 702.150 81.600 706.050 83.700 ;
        RECT 697.950 75.750 699.750 81.600 ;
        RECT 702.150 75.750 703.950 81.600 ;
        RECT 706.650 75.750 708.450 78.600 ;
        RECT 709.650 75.750 711.450 87.600 ;
        RECT 2.550 65.400 4.350 71.250 ;
        RECT 5.550 65.400 7.350 71.250 ;
        RECT 8.550 65.400 10.350 71.250 ;
        RECT 14.550 65.400 16.350 71.250 ;
        RECT 17.550 65.400 19.350 71.250 ;
        RECT 20.550 65.400 22.350 71.250 ;
        RECT 28.650 65.400 30.450 71.250 ;
        RECT 31.650 65.400 33.450 71.250 ;
        RECT 34.650 65.400 36.450 71.250 ;
        RECT 40.650 65.400 42.450 71.250 ;
        RECT 43.650 65.400 45.450 71.250 ;
        RECT 46.650 65.400 48.450 71.250 ;
        RECT 5.550 57.150 6.750 65.400 ;
        RECT 17.550 57.150 18.750 65.400 ;
        RECT 32.250 57.150 33.450 65.400 ;
        RECT 34.950 60.450 37.050 61.050 ;
        RECT 34.950 59.550 39.450 60.450 ;
        RECT 34.950 58.950 37.050 59.550 ;
        RECT 1.950 53.850 4.050 55.950 ;
        RECT 4.950 55.050 7.050 57.150 ;
        RECT 2.100 52.050 3.900 53.850 ;
        RECT 5.550 47.700 6.750 55.050 ;
        RECT 7.950 53.850 10.050 55.950 ;
        RECT 13.950 53.850 16.050 55.950 ;
        RECT 16.950 55.050 19.050 57.150 ;
        RECT 8.100 52.050 9.900 53.850 ;
        RECT 14.100 52.050 15.900 53.850 ;
        RECT 17.550 47.700 18.750 55.050 ;
        RECT 19.950 53.850 22.050 55.950 ;
        RECT 28.950 53.850 31.050 55.950 ;
        RECT 31.950 55.050 34.050 57.150 ;
        RECT 20.100 52.050 21.900 53.850 ;
        RECT 29.100 52.050 30.900 53.850 ;
        RECT 32.250 47.700 33.450 55.050 ;
        RECT 34.950 53.850 37.050 55.950 ;
        RECT 35.100 52.050 36.900 53.850 ;
        RECT 38.550 52.050 39.450 59.550 ;
        RECT 44.250 57.150 45.450 65.400 ;
        RECT 52.050 59.400 53.850 71.250 ;
        RECT 55.050 59.400 56.850 71.250 ;
        RECT 58.650 65.400 60.450 71.250 ;
        RECT 61.650 65.400 63.450 71.250 ;
        RECT 67.650 65.400 69.450 71.250 ;
        RECT 70.650 65.400 72.450 71.250 ;
        RECT 73.650 65.400 75.450 71.250 ;
        RECT 79.650 65.400 81.450 71.250 ;
        RECT 82.650 66.000 84.450 71.250 ;
        RECT 40.950 53.850 43.050 55.950 ;
        RECT 43.950 55.050 46.050 57.150 ;
        RECT 41.100 52.050 42.900 53.850 ;
        RECT 37.950 49.950 40.050 52.050 ;
        RECT 44.250 47.700 45.450 55.050 ;
        RECT 46.950 53.850 49.050 55.950 ;
        RECT 52.650 54.150 53.850 59.400 ;
        RECT 47.100 52.050 48.900 53.850 ;
        RECT 52.650 52.050 55.050 54.150 ;
        RECT 55.950 53.850 58.050 55.950 ;
        RECT 56.100 52.050 57.900 53.850 ;
        RECT 5.550 46.800 9.150 47.700 ;
        RECT 17.550 46.800 21.150 47.700 ;
        RECT 2.850 39.750 4.650 45.600 ;
        RECT 7.350 39.750 9.150 46.800 ;
        RECT 14.850 39.750 16.650 45.600 ;
        RECT 19.350 39.750 21.150 46.800 ;
        RECT 29.850 46.800 33.450 47.700 ;
        RECT 41.850 46.800 45.450 47.700 ;
        RECT 29.850 39.750 31.650 46.800 ;
        RECT 34.350 39.750 36.150 45.600 ;
        RECT 41.850 39.750 43.650 46.800 ;
        RECT 52.650 45.600 53.850 52.050 ;
        RECT 59.100 48.300 60.300 65.400 ;
        RECT 61.950 60.450 64.050 61.050 ;
        RECT 61.950 59.550 66.450 60.450 ;
        RECT 61.950 58.950 64.050 59.550 ;
        RECT 62.100 54.150 63.900 55.950 ;
        RECT 61.950 52.050 64.050 54.150 ;
        RECT 55.950 47.100 63.450 48.300 ;
        RECT 55.950 46.500 57.750 47.100 ;
        RECT 46.350 39.750 48.150 45.600 ;
        RECT 52.650 44.100 55.950 45.600 ;
        RECT 54.150 39.750 55.950 44.100 ;
        RECT 57.150 39.750 58.950 45.600 ;
        RECT 61.650 39.750 63.450 47.100 ;
        RECT 65.550 46.050 66.450 59.550 ;
        RECT 71.250 57.150 72.450 65.400 ;
        RECT 80.250 65.100 81.450 65.400 ;
        RECT 85.650 65.400 87.450 71.250 ;
        RECT 88.650 65.400 90.450 71.250 ;
        RECT 94.650 70.500 102.450 71.250 ;
        RECT 85.650 65.100 87.300 65.400 ;
        RECT 80.250 64.200 87.300 65.100 ;
        RECT 67.950 53.850 70.050 55.950 ;
        RECT 70.950 55.050 73.050 57.150 ;
        RECT 80.250 55.950 81.300 64.200 ;
        RECT 86.100 60.150 87.900 61.950 ;
        RECT 82.950 57.150 84.750 58.950 ;
        RECT 85.950 58.050 88.050 60.150 ;
        RECT 94.650 59.400 96.450 70.500 ;
        RECT 97.650 59.400 99.450 69.600 ;
        RECT 100.650 60.600 102.450 70.500 ;
        RECT 103.650 61.500 105.450 71.250 ;
        RECT 106.650 60.600 108.450 71.250 ;
        RECT 100.650 59.700 108.450 60.600 ;
        RECT 114.450 59.400 116.250 71.250 ;
        RECT 118.650 59.400 120.450 71.250 ;
        RECT 124.650 65.400 126.450 71.250 ;
        RECT 127.650 65.400 129.450 71.250 ;
        RECT 130.650 65.400 132.450 71.250 ;
        RECT 134.550 65.400 136.350 71.250 ;
        RECT 137.550 65.400 139.350 71.250 ;
        RECT 140.550 65.400 142.350 71.250 ;
        RECT 148.650 65.400 150.450 71.250 ;
        RECT 151.650 65.400 153.450 71.250 ;
        RECT 154.650 65.400 156.450 71.250 ;
        RECT 160.650 65.400 162.450 71.250 ;
        RECT 163.650 65.400 165.450 71.250 ;
        RECT 166.650 65.400 168.450 71.250 ;
        RECT 172.650 70.500 180.450 71.250 ;
        RECT 89.100 57.150 90.900 58.950 ;
        RECT 97.800 58.500 99.600 59.400 ;
        RECT 97.800 57.600 101.850 58.500 ;
        RECT 114.450 58.350 117.000 59.400 ;
        RECT 68.100 52.050 69.900 53.850 ;
        RECT 71.250 47.700 72.450 55.050 ;
        RECT 73.950 53.850 76.050 55.950 ;
        RECT 79.950 53.850 82.050 55.950 ;
        RECT 82.950 55.050 85.050 57.150 ;
        RECT 88.950 55.050 91.050 57.150 ;
        RECT 95.100 54.150 96.900 55.950 ;
        RECT 100.950 54.150 101.850 57.600 ;
        RECT 106.950 54.150 108.750 55.950 ;
        RECT 113.100 54.150 114.900 55.950 ;
        RECT 74.100 52.050 75.900 53.850 ;
        RECT 80.400 49.650 81.600 53.850 ;
        RECT 94.950 52.050 97.050 54.150 ;
        RECT 97.950 50.850 100.050 52.950 ;
        RECT 100.950 52.050 103.050 54.150 ;
        RECT 80.400 48.000 84.900 49.650 ;
        RECT 98.250 49.050 100.050 50.850 ;
        RECT 68.850 46.800 72.450 47.700 ;
        RECT 64.950 43.950 67.050 46.050 ;
        RECT 68.850 39.750 70.650 46.800 ;
        RECT 73.350 39.750 75.150 45.600 ;
        RECT 83.100 39.750 84.900 48.000 ;
        RECT 88.500 39.750 90.300 48.600 ;
        RECT 102.000 45.600 103.050 52.050 ;
        RECT 103.950 50.850 106.050 52.950 ;
        RECT 106.950 52.050 109.050 54.150 ;
        RECT 112.950 52.050 115.050 54.150 ;
        RECT 115.950 51.150 117.000 58.350 ;
        RECT 128.250 57.150 129.450 65.400 ;
        RECT 137.550 57.150 138.750 65.400 ;
        RECT 152.250 57.150 153.450 65.400 ;
        RECT 164.250 57.150 165.450 65.400 ;
        RECT 172.650 59.400 174.450 70.500 ;
        RECT 175.650 59.400 177.450 69.600 ;
        RECT 178.650 60.600 180.450 70.500 ;
        RECT 181.650 61.500 183.450 71.250 ;
        RECT 184.650 60.600 186.450 71.250 ;
        RECT 178.650 59.700 186.450 60.600 ;
        RECT 189.300 59.400 191.100 71.250 ;
        RECT 193.500 59.400 195.300 71.250 ;
        RECT 196.800 65.400 198.600 71.250 ;
        RECT 207.450 59.400 209.250 71.250 ;
        RECT 211.650 59.400 213.450 71.250 ;
        RECT 216.300 59.400 218.100 71.250 ;
        RECT 220.500 59.400 222.300 71.250 ;
        RECT 223.800 65.400 225.600 71.250 ;
        RECT 230.550 65.400 232.350 71.250 ;
        RECT 233.550 65.400 235.350 71.250 ;
        RECT 175.800 58.500 177.600 59.400 ;
        RECT 175.800 57.600 179.850 58.500 ;
        RECT 119.100 54.150 120.900 55.950 ;
        RECT 118.950 52.050 121.050 54.150 ;
        RECT 124.950 53.850 127.050 55.950 ;
        RECT 127.950 55.050 130.050 57.150 ;
        RECT 125.100 52.050 126.900 53.850 ;
        RECT 103.950 49.050 105.750 50.850 ;
        RECT 115.950 49.050 118.050 51.150 ;
        RECT 97.800 39.750 99.600 45.600 ;
        RECT 102.000 39.750 103.800 45.600 ;
        RECT 106.200 39.750 108.000 45.600 ;
        RECT 115.950 42.600 117.000 49.050 ;
        RECT 128.250 47.700 129.450 55.050 ;
        RECT 130.950 53.850 133.050 55.950 ;
        RECT 133.950 53.850 136.050 55.950 ;
        RECT 136.950 55.050 139.050 57.150 ;
        RECT 131.100 52.050 132.900 53.850 ;
        RECT 134.100 52.050 135.900 53.850 ;
        RECT 125.850 46.800 129.450 47.700 ;
        RECT 137.550 47.700 138.750 55.050 ;
        RECT 139.950 53.850 142.050 55.950 ;
        RECT 148.950 53.850 151.050 55.950 ;
        RECT 151.950 55.050 154.050 57.150 ;
        RECT 140.100 52.050 141.900 53.850 ;
        RECT 149.100 52.050 150.900 53.850 ;
        RECT 152.250 47.700 153.450 55.050 ;
        RECT 154.950 53.850 157.050 55.950 ;
        RECT 160.950 53.850 163.050 55.950 ;
        RECT 163.950 55.050 166.050 57.150 ;
        RECT 155.100 52.050 156.900 53.850 ;
        RECT 161.100 52.050 162.900 53.850 ;
        RECT 164.250 47.700 165.450 55.050 ;
        RECT 166.950 53.850 169.050 55.950 ;
        RECT 173.100 54.150 174.900 55.950 ;
        RECT 178.950 54.150 179.850 57.600 ;
        RECT 184.950 54.150 186.750 55.950 ;
        RECT 188.100 54.150 189.900 55.950 ;
        RECT 193.950 54.150 195.150 59.400 ;
        RECT 196.950 57.150 198.750 58.950 ;
        RECT 207.450 58.350 210.000 59.400 ;
        RECT 196.950 55.050 199.050 57.150 ;
        RECT 206.100 54.150 207.900 55.950 ;
        RECT 167.100 52.050 168.900 53.850 ;
        RECT 172.950 52.050 175.050 54.150 ;
        RECT 175.950 50.850 178.050 52.950 ;
        RECT 178.950 52.050 181.050 54.150 ;
        RECT 176.250 49.050 178.050 50.850 ;
        RECT 137.550 46.800 141.150 47.700 ;
        RECT 112.650 39.750 114.450 42.600 ;
        RECT 115.650 39.750 117.450 42.600 ;
        RECT 118.650 39.750 120.450 42.600 ;
        RECT 125.850 39.750 127.650 46.800 ;
        RECT 130.350 39.750 132.150 45.600 ;
        RECT 134.850 39.750 136.650 45.600 ;
        RECT 139.350 39.750 141.150 46.800 ;
        RECT 149.850 46.800 153.450 47.700 ;
        RECT 161.850 46.800 165.450 47.700 ;
        RECT 149.850 39.750 151.650 46.800 ;
        RECT 154.350 39.750 156.150 45.600 ;
        RECT 161.850 39.750 163.650 46.800 ;
        RECT 180.000 45.600 181.050 52.050 ;
        RECT 181.950 50.850 184.050 52.950 ;
        RECT 184.950 52.050 187.050 54.150 ;
        RECT 187.950 52.050 190.050 54.150 ;
        RECT 190.950 50.850 193.050 52.950 ;
        RECT 193.950 52.050 196.050 54.150 ;
        RECT 205.950 52.050 208.050 54.150 ;
        RECT 181.950 49.050 183.750 50.850 ;
        RECT 191.100 49.050 192.900 50.850 ;
        RECT 194.850 48.750 196.050 52.050 ;
        RECT 208.950 51.150 210.000 58.350 ;
        RECT 212.100 54.150 213.900 55.950 ;
        RECT 215.100 54.150 216.900 55.950 ;
        RECT 220.950 54.150 222.150 59.400 ;
        RECT 223.950 57.150 225.750 58.950 ;
        RECT 223.950 55.050 226.050 57.150 ;
        RECT 211.950 52.050 214.050 54.150 ;
        RECT 214.950 52.050 217.050 54.150 ;
        RECT 208.950 49.050 211.050 51.150 ;
        RECT 217.950 50.850 220.050 52.950 ;
        RECT 220.950 52.050 223.050 54.150 ;
        RECT 233.400 52.950 234.600 65.400 ;
        RECT 241.650 59.400 243.450 71.250 ;
        RECT 244.650 60.300 246.450 71.250 ;
        RECT 247.650 61.200 249.450 71.250 ;
        RECT 250.650 60.300 252.450 71.250 ;
        RECT 254.550 65.400 256.350 71.250 ;
        RECT 257.550 65.400 259.350 71.250 ;
        RECT 263.550 65.400 265.350 71.250 ;
        RECT 266.550 65.400 268.350 71.250 ;
        RECT 269.550 66.000 271.350 71.250 ;
        RECT 244.650 59.400 252.450 60.300 ;
        RECT 242.100 54.150 243.300 59.400 ;
        RECT 218.100 49.050 219.900 50.850 ;
        RECT 195.000 47.700 198.750 48.750 ;
        RECT 166.350 39.750 168.150 45.600 ;
        RECT 175.800 39.750 177.600 45.600 ;
        RECT 180.000 39.750 181.800 45.600 ;
        RECT 184.200 39.750 186.000 45.600 ;
        RECT 188.550 44.700 196.350 46.050 ;
        RECT 188.550 39.750 190.350 44.700 ;
        RECT 191.550 39.750 193.350 43.800 ;
        RECT 194.550 39.750 196.350 44.700 ;
        RECT 197.550 45.600 198.750 47.700 ;
        RECT 197.550 39.750 199.350 45.600 ;
        RECT 208.950 42.600 210.000 49.050 ;
        RECT 221.850 48.750 223.050 52.050 ;
        RECT 230.100 51.150 231.900 52.950 ;
        RECT 229.950 49.050 232.050 51.150 ;
        RECT 232.950 50.850 235.050 52.950 ;
        RECT 241.950 52.050 244.050 54.150 ;
        RECT 257.400 52.950 258.600 65.400 ;
        RECT 266.700 65.100 268.350 65.400 ;
        RECT 272.550 65.400 274.350 71.250 ;
        RECT 272.550 65.100 273.750 65.400 ;
        RECT 266.700 64.200 273.750 65.100 ;
        RECT 266.100 60.150 267.900 61.950 ;
        RECT 263.100 57.150 264.900 58.950 ;
        RECT 265.950 58.050 268.050 60.150 ;
        RECT 269.250 57.150 271.050 58.950 ;
        RECT 262.950 55.050 265.050 57.150 ;
        RECT 268.950 55.050 271.050 57.150 ;
        RECT 272.700 55.950 273.750 64.200 ;
        RECT 278.550 60.300 280.350 71.250 ;
        RECT 281.550 61.200 283.350 71.250 ;
        RECT 284.550 60.300 286.350 71.250 ;
        RECT 278.550 59.400 286.350 60.300 ;
        RECT 287.550 59.400 289.350 71.250 ;
        RECT 293.550 65.400 295.350 71.250 ;
        RECT 296.550 65.400 298.350 71.250 ;
        RECT 299.550 65.400 301.350 71.250 ;
        RECT 305.550 65.400 307.350 71.250 ;
        RECT 308.550 65.400 310.350 71.250 ;
        RECT 311.550 65.400 313.350 71.250 ;
        RECT 317.550 65.400 319.350 71.250 ;
        RECT 320.550 65.400 322.350 71.250 ;
        RECT 323.550 65.400 325.350 71.250 ;
        RECT 259.950 52.950 262.050 55.050 ;
        RECT 271.950 53.850 274.050 55.950 ;
        RECT 287.700 54.150 288.900 59.400 ;
        RECT 296.550 57.150 297.750 65.400 ;
        RECT 222.000 47.700 225.750 48.750 ;
        RECT 215.550 44.700 223.350 46.050 ;
        RECT 205.650 39.750 207.450 42.600 ;
        RECT 208.650 39.750 210.450 42.600 ;
        RECT 211.650 39.750 213.450 42.600 ;
        RECT 215.550 39.750 217.350 44.700 ;
        RECT 218.550 39.750 220.350 43.800 ;
        RECT 221.550 39.750 223.350 44.700 ;
        RECT 224.550 45.600 225.750 47.700 ;
        RECT 224.550 39.750 226.350 45.600 ;
        RECT 233.400 42.600 234.600 50.850 ;
        RECT 242.100 45.600 243.300 52.050 ;
        RECT 244.950 50.850 247.050 52.950 ;
        RECT 248.100 51.150 249.900 52.950 ;
        RECT 245.100 49.050 246.900 50.850 ;
        RECT 247.950 49.050 250.050 51.150 ;
        RECT 250.950 50.850 253.050 52.950 ;
        RECT 254.100 51.150 255.900 52.950 ;
        RECT 251.100 49.050 252.900 50.850 ;
        RECT 253.950 49.050 256.050 51.150 ;
        RECT 256.950 50.850 259.050 52.950 ;
        RECT 260.550 51.450 261.450 52.950 ;
        RECT 262.950 51.450 265.050 52.050 ;
        RECT 242.100 43.950 247.800 45.600 ;
        RECT 230.550 39.750 232.350 42.600 ;
        RECT 233.550 39.750 235.350 42.600 ;
        RECT 242.700 39.750 244.500 42.600 ;
        RECT 246.000 39.750 247.800 43.950 ;
        RECT 250.200 39.750 252.000 45.600 ;
        RECT 257.400 42.600 258.600 50.850 ;
        RECT 260.550 50.550 265.050 51.450 ;
        RECT 262.950 49.950 265.050 50.550 ;
        RECT 272.400 49.650 273.600 53.850 ;
        RECT 277.950 50.850 280.050 52.950 ;
        RECT 281.100 51.150 282.900 52.950 ;
        RECT 254.550 39.750 256.350 42.600 ;
        RECT 257.550 39.750 259.350 42.600 ;
        RECT 263.700 39.750 265.500 48.600 ;
        RECT 269.100 48.000 273.600 49.650 ;
        RECT 278.100 49.050 279.900 50.850 ;
        RECT 280.950 49.050 283.050 51.150 ;
        RECT 283.950 50.850 286.050 52.950 ;
        RECT 286.950 52.050 289.050 54.150 ;
        RECT 292.950 53.850 295.050 55.950 ;
        RECT 295.950 55.050 298.050 57.150 ;
        RECT 301.950 55.950 304.050 58.050 ;
        RECT 308.550 57.150 309.750 65.400 ;
        RECT 320.550 57.150 321.750 65.400 ;
        RECT 325.950 60.450 328.050 61.050 ;
        RECT 325.950 59.550 330.450 60.450 ;
        RECT 325.950 58.950 328.050 59.550 ;
        RECT 293.100 52.050 294.900 53.850 ;
        RECT 284.100 49.050 285.900 50.850 ;
        RECT 269.100 39.750 270.900 48.000 ;
        RECT 287.700 45.600 288.900 52.050 ;
        RECT 296.550 47.700 297.750 55.050 ;
        RECT 298.950 53.850 301.050 55.950 ;
        RECT 299.100 52.050 300.900 53.850 ;
        RECT 302.550 48.450 303.450 55.950 ;
        RECT 304.950 53.850 307.050 55.950 ;
        RECT 307.950 55.050 310.050 57.150 ;
        RECT 305.100 52.050 306.900 53.850 ;
        RECT 304.950 48.450 307.050 49.050 ;
        RECT 296.550 46.800 300.150 47.700 ;
        RECT 302.550 47.550 307.050 48.450 ;
        RECT 304.950 46.950 307.050 47.550 ;
        RECT 308.550 47.700 309.750 55.050 ;
        RECT 310.950 53.850 313.050 55.950 ;
        RECT 316.950 53.850 319.050 55.950 ;
        RECT 319.950 55.050 322.050 57.150 ;
        RECT 311.100 52.050 312.900 53.850 ;
        RECT 317.100 52.050 318.900 53.850 ;
        RECT 320.550 47.700 321.750 55.050 ;
        RECT 322.950 53.850 325.050 55.950 ;
        RECT 323.100 52.050 324.900 53.850 ;
        RECT 329.550 52.050 330.450 59.550 ;
        RECT 333.450 59.400 335.250 71.250 ;
        RECT 337.650 59.400 339.450 71.250 ;
        RECT 343.650 65.400 345.450 71.250 ;
        RECT 346.650 65.400 348.450 71.250 ;
        RECT 349.650 65.400 351.450 71.250 ;
        RECT 333.450 58.350 336.000 59.400 ;
        RECT 332.100 54.150 333.900 55.950 ;
        RECT 331.950 52.050 334.050 54.150 ;
        RECT 328.950 49.950 331.050 52.050 ;
        RECT 334.950 51.150 336.000 58.350 ;
        RECT 347.250 57.150 348.450 65.400 ;
        RECT 353.550 59.400 355.350 71.250 ;
        RECT 357.750 59.400 359.550 71.250 ;
        RECT 365.550 65.400 367.350 71.250 ;
        RECT 368.550 65.400 370.350 71.250 ;
        RECT 371.550 66.000 373.350 71.250 ;
        RECT 368.700 65.100 370.350 65.400 ;
        RECT 374.550 65.400 376.350 71.250 ;
        RECT 382.650 65.400 384.450 71.250 ;
        RECT 385.650 65.400 387.450 71.250 ;
        RECT 391.650 65.400 393.450 71.250 ;
        RECT 394.650 66.000 396.450 71.250 ;
        RECT 374.550 65.100 375.750 65.400 ;
        RECT 368.700 64.200 375.750 65.100 ;
        RECT 368.100 60.150 369.900 61.950 ;
        RECT 357.000 58.350 359.550 59.400 ;
        RECT 338.100 54.150 339.900 55.950 ;
        RECT 337.950 52.050 340.050 54.150 ;
        RECT 343.950 53.850 346.050 55.950 ;
        RECT 346.950 55.050 349.050 57.150 ;
        RECT 344.100 52.050 345.900 53.850 ;
        RECT 334.950 49.050 337.050 51.150 ;
        RECT 308.550 46.800 312.150 47.700 ;
        RECT 320.550 46.800 324.150 47.700 ;
        RECT 279.000 39.750 280.800 45.600 ;
        RECT 283.200 43.950 288.900 45.600 ;
        RECT 283.200 39.750 285.000 43.950 ;
        RECT 286.500 39.750 288.300 42.600 ;
        RECT 293.850 39.750 295.650 45.600 ;
        RECT 298.350 39.750 300.150 46.800 ;
        RECT 305.850 39.750 307.650 45.600 ;
        RECT 310.350 39.750 312.150 46.800 ;
        RECT 317.850 39.750 319.650 45.600 ;
        RECT 322.350 39.750 324.150 46.800 ;
        RECT 334.950 42.600 336.000 49.050 ;
        RECT 347.250 47.700 348.450 55.050 ;
        RECT 349.950 53.850 352.050 55.950 ;
        RECT 353.100 54.150 354.900 55.950 ;
        RECT 350.100 52.050 351.900 53.850 ;
        RECT 352.950 52.050 355.050 54.150 ;
        RECT 357.000 51.150 358.050 58.350 ;
        RECT 365.100 57.150 366.900 58.950 ;
        RECT 367.950 58.050 370.050 60.150 ;
        RECT 371.250 57.150 373.050 58.950 ;
        RECT 359.100 54.150 360.900 55.950 ;
        RECT 364.950 55.050 367.050 57.150 ;
        RECT 370.950 55.050 373.050 57.150 ;
        RECT 374.700 55.950 375.750 64.200 ;
        RECT 358.950 52.050 361.050 54.150 ;
        RECT 373.950 53.850 376.050 55.950 ;
        RECT 355.950 49.050 358.050 51.150 ;
        RECT 374.400 49.650 375.600 53.850 ;
        RECT 383.400 52.950 384.600 65.400 ;
        RECT 392.250 65.100 393.450 65.400 ;
        RECT 397.650 65.400 399.450 71.250 ;
        RECT 400.650 65.400 402.450 71.250 ;
        RECT 397.650 65.100 399.300 65.400 ;
        RECT 392.250 64.200 399.300 65.100 ;
        RECT 392.250 55.950 393.300 64.200 ;
        RECT 398.100 60.150 399.900 61.950 ;
        RECT 404.550 60.300 406.350 71.250 ;
        RECT 407.550 61.200 409.350 71.250 ;
        RECT 410.550 60.300 412.350 71.250 ;
        RECT 394.950 57.150 396.750 58.950 ;
        RECT 397.950 58.050 400.050 60.150 ;
        RECT 404.550 59.400 412.350 60.300 ;
        RECT 413.550 59.400 415.350 71.250 ;
        RECT 419.550 59.400 421.350 71.250 ;
        RECT 423.750 59.400 425.550 71.250 ;
        RECT 433.650 65.400 435.450 71.250 ;
        RECT 436.650 65.400 438.450 71.250 ;
        RECT 439.650 65.400 441.450 71.250 ;
        RECT 446.400 65.400 448.200 71.250 ;
        RECT 401.100 57.150 402.900 58.950 ;
        RECT 391.950 53.850 394.050 55.950 ;
        RECT 394.950 55.050 397.050 57.150 ;
        RECT 400.950 55.050 403.050 57.150 ;
        RECT 413.700 54.150 414.900 59.400 ;
        RECT 423.000 58.350 425.550 59.400 ;
        RECT 419.100 54.150 420.900 55.950 ;
        RECT 382.950 50.850 385.050 52.950 ;
        RECT 386.100 51.150 387.900 52.950 ;
        RECT 344.850 46.800 348.450 47.700 ;
        RECT 331.650 39.750 333.450 42.600 ;
        RECT 334.650 39.750 336.450 42.600 ;
        RECT 337.650 39.750 339.450 42.600 ;
        RECT 344.850 39.750 346.650 46.800 ;
        RECT 349.350 39.750 351.150 45.600 ;
        RECT 357.000 42.600 358.050 49.050 ;
        RECT 353.550 39.750 355.350 42.600 ;
        RECT 356.550 39.750 358.350 42.600 ;
        RECT 359.550 39.750 361.350 42.600 ;
        RECT 365.700 39.750 367.500 48.600 ;
        RECT 371.100 48.000 375.600 49.650 ;
        RECT 371.100 39.750 372.900 48.000 ;
        RECT 383.400 42.600 384.600 50.850 ;
        RECT 385.950 49.050 388.050 51.150 ;
        RECT 392.400 49.650 393.600 53.850 ;
        RECT 403.950 50.850 406.050 52.950 ;
        RECT 407.100 51.150 408.900 52.950 ;
        RECT 392.400 48.000 396.900 49.650 ;
        RECT 404.100 49.050 405.900 50.850 ;
        RECT 406.950 49.050 409.050 51.150 ;
        RECT 409.950 50.850 412.050 52.950 ;
        RECT 412.950 52.050 415.050 54.150 ;
        RECT 418.950 52.050 421.050 54.150 ;
        RECT 410.100 49.050 411.900 50.850 ;
        RECT 382.650 39.750 384.450 42.600 ;
        RECT 385.650 39.750 387.450 42.600 ;
        RECT 395.100 39.750 396.900 48.000 ;
        RECT 400.500 39.750 402.300 48.600 ;
        RECT 413.700 45.600 414.900 52.050 ;
        RECT 423.000 51.150 424.050 58.350 ;
        RECT 437.250 57.150 438.450 65.400 ;
        RECT 449.700 59.400 451.500 71.250 ;
        RECT 453.900 59.400 455.700 71.250 ;
        RECT 461.400 65.400 463.200 71.250 ;
        RECT 464.700 59.400 466.500 71.250 ;
        RECT 468.900 59.400 470.700 71.250 ;
        RECT 477.450 59.400 479.250 71.250 ;
        RECT 481.650 59.400 483.450 71.250 ;
        RECT 487.650 65.400 489.450 71.250 ;
        RECT 490.650 65.400 492.450 71.250 ;
        RECT 497.400 65.400 499.200 71.250 ;
        RECT 446.250 57.150 448.050 58.950 ;
        RECT 425.100 54.150 426.900 55.950 ;
        RECT 424.950 52.050 427.050 54.150 ;
        RECT 433.950 53.850 436.050 55.950 ;
        RECT 436.950 55.050 439.050 57.150 ;
        RECT 434.100 52.050 435.900 53.850 ;
        RECT 421.950 49.050 424.050 51.150 ;
        RECT 405.000 39.750 406.800 45.600 ;
        RECT 409.200 43.950 414.900 45.600 ;
        RECT 409.200 39.750 411.000 43.950 ;
        RECT 423.000 42.600 424.050 49.050 ;
        RECT 437.250 47.700 438.450 55.050 ;
        RECT 439.950 53.850 442.050 55.950 ;
        RECT 445.950 55.050 448.050 57.150 ;
        RECT 449.850 54.150 451.050 59.400 ;
        RECT 461.250 57.150 463.050 58.950 ;
        RECT 455.100 54.150 456.900 55.950 ;
        RECT 460.950 55.050 463.050 57.150 ;
        RECT 464.850 54.150 466.050 59.400 ;
        RECT 477.450 58.350 480.000 59.400 ;
        RECT 470.100 54.150 471.900 55.950 ;
        RECT 476.100 54.150 477.900 55.950 ;
        RECT 440.100 52.050 441.900 53.850 ;
        RECT 448.950 52.050 451.050 54.150 ;
        RECT 448.950 48.750 450.150 52.050 ;
        RECT 451.950 50.850 454.050 52.950 ;
        RECT 454.950 52.050 457.050 54.150 ;
        RECT 463.950 52.050 466.050 54.150 ;
        RECT 452.100 49.050 453.900 50.850 ;
        RECT 463.950 48.750 465.150 52.050 ;
        RECT 466.950 50.850 469.050 52.950 ;
        RECT 469.950 52.050 472.050 54.150 ;
        RECT 475.950 52.050 478.050 54.150 ;
        RECT 478.950 51.150 480.000 58.350 ;
        RECT 482.100 54.150 483.900 55.950 ;
        RECT 481.950 52.050 484.050 54.150 ;
        RECT 488.400 52.950 489.600 65.400 ;
        RECT 500.700 59.400 502.500 71.250 ;
        RECT 504.900 59.400 506.700 71.250 ;
        RECT 511.650 59.400 513.450 71.250 ;
        RECT 514.650 60.300 516.450 71.250 ;
        RECT 517.650 61.200 519.450 71.250 ;
        RECT 520.650 60.300 522.450 71.250 ;
        RECT 514.650 59.400 522.450 60.300 ;
        RECT 528.450 59.400 530.250 71.250 ;
        RECT 532.650 59.400 534.450 71.250 ;
        RECT 536.550 59.400 538.350 71.250 ;
        RECT 541.050 59.550 542.850 71.250 ;
        RECT 544.050 60.900 545.850 71.250 ;
        RECT 551.550 65.400 553.350 71.250 ;
        RECT 554.550 65.400 556.350 71.250 ;
        RECT 557.550 65.400 559.350 71.250 ;
        RECT 563.550 65.400 565.350 71.250 ;
        RECT 566.550 65.400 568.350 71.250 ;
        RECT 569.550 65.400 571.350 71.250 ;
        RECT 578.400 65.400 580.200 71.250 ;
        RECT 544.050 59.550 546.450 60.900 ;
        RECT 497.250 57.150 499.050 58.950 ;
        RECT 496.950 55.050 499.050 57.150 ;
        RECT 500.850 54.150 502.050 59.400 ;
        RECT 506.100 54.150 507.900 55.950 ;
        RECT 512.100 54.150 513.300 59.400 ;
        RECT 528.450 58.350 531.000 59.400 ;
        RECT 527.100 54.150 528.900 55.950 ;
        RECT 467.100 49.050 468.900 50.850 ;
        RECT 478.950 49.050 481.050 51.150 ;
        RECT 487.950 50.850 490.050 52.950 ;
        RECT 491.100 51.150 492.900 52.950 ;
        RECT 499.950 52.050 502.050 54.150 ;
        RECT 434.850 46.800 438.450 47.700 ;
        RECT 446.250 47.700 450.000 48.750 ;
        RECT 461.250 47.700 465.000 48.750 ;
        RECT 412.500 39.750 414.300 42.600 ;
        RECT 419.550 39.750 421.350 42.600 ;
        RECT 422.550 39.750 424.350 42.600 ;
        RECT 425.550 39.750 427.350 42.600 ;
        RECT 434.850 39.750 436.650 46.800 ;
        RECT 446.250 45.600 447.450 47.700 ;
        RECT 439.350 39.750 441.150 45.600 ;
        RECT 445.650 39.750 447.450 45.600 ;
        RECT 448.650 44.700 456.450 46.050 ;
        RECT 461.250 45.600 462.450 47.700 ;
        RECT 448.650 39.750 450.450 44.700 ;
        RECT 451.650 39.750 453.450 43.800 ;
        RECT 454.650 39.750 456.450 44.700 ;
        RECT 460.650 39.750 462.450 45.600 ;
        RECT 463.650 44.700 471.450 46.050 ;
        RECT 463.650 39.750 465.450 44.700 ;
        RECT 466.650 39.750 468.450 43.800 ;
        RECT 469.650 39.750 471.450 44.700 ;
        RECT 478.950 42.600 480.000 49.050 ;
        RECT 488.400 42.600 489.600 50.850 ;
        RECT 490.950 49.050 493.050 51.150 ;
        RECT 499.950 48.750 501.150 52.050 ;
        RECT 502.950 50.850 505.050 52.950 ;
        RECT 505.950 52.050 508.050 54.150 ;
        RECT 511.950 52.050 514.050 54.150 ;
        RECT 503.100 49.050 504.900 50.850 ;
        RECT 497.250 47.700 501.000 48.750 ;
        RECT 497.250 45.600 498.450 47.700 ;
        RECT 475.650 39.750 477.450 42.600 ;
        RECT 478.650 39.750 480.450 42.600 ;
        RECT 481.650 39.750 483.450 42.600 ;
        RECT 487.650 39.750 489.450 42.600 ;
        RECT 490.650 39.750 492.450 42.600 ;
        RECT 496.650 39.750 498.450 45.600 ;
        RECT 499.650 44.700 507.450 46.050 ;
        RECT 499.650 39.750 501.450 44.700 ;
        RECT 502.650 39.750 504.450 43.800 ;
        RECT 505.650 39.750 507.450 44.700 ;
        RECT 512.100 45.600 513.300 52.050 ;
        RECT 514.950 50.850 517.050 52.950 ;
        RECT 518.100 51.150 519.900 52.950 ;
        RECT 515.100 49.050 516.900 50.850 ;
        RECT 517.950 49.050 520.050 51.150 ;
        RECT 520.950 50.850 523.050 52.950 ;
        RECT 526.950 52.050 529.050 54.150 ;
        RECT 529.950 51.150 531.000 58.350 ;
        RECT 536.550 58.200 537.750 59.400 ;
        RECT 541.950 58.200 543.750 58.650 ;
        RECT 536.550 57.000 543.750 58.200 ;
        RECT 541.950 56.850 543.750 57.000 ;
        RECT 533.100 54.150 534.900 55.950 ;
        RECT 539.100 54.150 540.900 55.950 ;
        RECT 532.950 52.050 535.050 54.150 ;
        RECT 536.100 51.150 537.900 52.950 ;
        RECT 538.950 52.050 541.050 54.150 ;
        RECT 521.100 49.050 522.900 50.850 ;
        RECT 529.950 49.050 532.050 51.150 ;
        RECT 535.950 49.050 538.050 51.150 ;
        RECT 512.100 43.950 517.800 45.600 ;
        RECT 512.700 39.750 514.500 42.600 ;
        RECT 516.000 39.750 517.800 43.950 ;
        RECT 520.200 39.750 522.000 45.600 ;
        RECT 529.950 42.600 531.000 49.050 ;
        RECT 542.700 48.600 543.600 56.850 ;
        RECT 545.100 52.950 546.450 59.550 ;
        RECT 554.550 57.150 555.750 65.400 ;
        RECT 566.550 57.150 567.750 65.400 ;
        RECT 581.700 59.400 583.500 71.250 ;
        RECT 585.900 59.400 587.700 71.250 ;
        RECT 592.650 65.400 594.450 71.250 ;
        RECT 595.650 65.400 597.450 71.250 ;
        RECT 601.650 65.400 603.450 71.250 ;
        RECT 604.650 65.400 606.450 71.250 ;
        RECT 578.250 57.150 580.050 58.950 ;
        RECT 550.950 53.850 553.050 55.950 ;
        RECT 553.950 55.050 556.050 57.150 ;
        RECT 544.950 50.850 547.050 52.950 ;
        RECT 551.100 52.050 552.900 53.850 ;
        RECT 541.950 47.700 543.750 48.600 ;
        RECT 540.450 46.800 543.750 47.700 ;
        RECT 540.450 42.600 541.350 46.800 ;
        RECT 546.000 45.600 547.050 50.850 ;
        RECT 554.550 47.700 555.750 55.050 ;
        RECT 556.950 53.850 559.050 55.950 ;
        RECT 562.950 53.850 565.050 55.950 ;
        RECT 565.950 55.050 568.050 57.150 ;
        RECT 557.100 52.050 558.900 53.850 ;
        RECT 563.100 52.050 564.900 53.850 ;
        RECT 566.550 47.700 567.750 55.050 ;
        RECT 568.950 53.850 571.050 55.950 ;
        RECT 577.950 55.050 580.050 57.150 ;
        RECT 581.850 54.150 583.050 59.400 ;
        RECT 587.100 54.150 588.900 55.950 ;
        RECT 569.100 52.050 570.900 53.850 ;
        RECT 580.950 52.050 583.050 54.150 ;
        RECT 580.950 48.750 582.150 52.050 ;
        RECT 583.950 50.850 586.050 52.950 ;
        RECT 586.950 52.050 589.050 54.150 ;
        RECT 593.400 52.950 594.600 65.400 ;
        RECT 602.400 52.950 603.600 65.400 ;
        RECT 608.550 59.400 610.350 71.250 ;
        RECT 611.550 68.400 613.350 71.250 ;
        RECT 616.050 65.400 617.850 71.250 ;
        RECT 620.250 65.400 622.050 71.250 ;
        RECT 613.950 63.300 617.850 65.400 ;
        RECT 624.150 64.500 625.950 71.250 ;
        RECT 627.150 65.400 628.950 71.250 ;
        RECT 631.950 65.400 633.750 71.250 ;
        RECT 637.050 65.400 638.850 71.250 ;
        RECT 632.250 64.500 633.450 65.400 ;
        RECT 622.950 62.700 629.850 64.500 ;
        RECT 632.250 62.400 637.050 64.500 ;
        RECT 615.150 60.600 617.850 62.400 ;
        RECT 618.750 61.800 620.550 62.400 ;
        RECT 618.750 60.900 625.050 61.800 ;
        RECT 632.250 61.500 633.450 62.400 ;
        RECT 618.750 60.600 620.550 60.900 ;
        RECT 616.950 59.700 617.850 60.600 ;
        RECT 592.950 50.850 595.050 52.950 ;
        RECT 596.100 51.150 597.900 52.950 ;
        RECT 584.100 49.050 585.900 50.850 ;
        RECT 578.250 47.700 582.000 48.750 ;
        RECT 554.550 46.800 558.150 47.700 ;
        RECT 566.550 46.800 570.150 47.700 ;
        RECT 526.650 39.750 528.450 42.600 ;
        RECT 529.650 39.750 531.450 42.600 ;
        RECT 532.650 39.750 534.450 42.600 ;
        RECT 536.550 39.750 538.350 42.600 ;
        RECT 539.550 39.750 541.350 42.600 ;
        RECT 542.550 39.750 544.350 42.600 ;
        RECT 545.550 39.750 547.350 45.600 ;
        RECT 551.850 39.750 553.650 45.600 ;
        RECT 556.350 39.750 558.150 46.800 ;
        RECT 563.850 39.750 565.650 45.600 ;
        RECT 568.350 39.750 570.150 46.800 ;
        RECT 578.250 45.600 579.450 47.700 ;
        RECT 577.650 39.750 579.450 45.600 ;
        RECT 580.650 44.700 588.450 46.050 ;
        RECT 580.650 39.750 582.450 44.700 ;
        RECT 583.650 39.750 585.450 43.800 ;
        RECT 586.650 39.750 588.450 44.700 ;
        RECT 593.400 42.600 594.600 50.850 ;
        RECT 595.950 49.050 598.050 51.150 ;
        RECT 601.950 50.850 604.050 52.950 ;
        RECT 605.100 51.150 606.900 52.950 ;
        RECT 602.400 42.600 603.600 50.850 ;
        RECT 604.950 49.050 607.050 51.150 ;
        RECT 608.550 49.950 609.750 59.400 ;
        RECT 613.950 58.800 616.050 59.700 ;
        RECT 616.950 58.800 622.950 59.700 ;
        RECT 611.850 57.600 616.050 58.800 ;
        RECT 610.950 55.800 612.750 57.600 ;
        RECT 622.050 54.150 622.950 58.800 ;
        RECT 624.150 58.800 625.050 60.900 ;
        RECT 625.950 60.300 633.450 61.500 ;
        RECT 625.950 59.700 627.750 60.300 ;
        RECT 640.050 59.400 641.850 71.250 ;
        RECT 646.650 65.400 648.450 71.250 ;
        RECT 649.650 65.400 651.450 71.250 ;
        RECT 652.650 65.400 654.450 71.250 ;
        RECT 659.400 65.400 661.200 71.250 ;
        RECT 630.750 58.800 641.850 59.400 ;
        RECT 624.150 58.200 641.850 58.800 ;
        RECT 624.150 57.900 632.550 58.200 ;
        RECT 630.750 57.600 632.550 57.900 ;
        RECT 622.050 52.050 625.050 54.150 ;
        RECT 628.950 53.100 631.050 54.150 ;
        RECT 628.950 52.050 636.900 53.100 ;
        RECT 610.950 51.750 613.050 52.050 ;
        RECT 610.950 49.950 614.850 51.750 ;
        RECT 608.550 47.850 613.050 49.950 ;
        RECT 622.050 48.000 622.950 52.050 ;
        RECT 635.100 51.300 636.900 52.050 ;
        RECT 638.100 51.150 639.900 52.950 ;
        RECT 632.100 50.400 633.900 51.000 ;
        RECT 638.100 50.400 639.000 51.150 ;
        RECT 632.100 49.200 639.000 50.400 ;
        RECT 632.100 48.000 633.150 49.200 ;
        RECT 608.550 45.600 609.750 47.850 ;
        RECT 622.050 47.100 633.150 48.000 ;
        RECT 622.050 46.800 622.950 47.100 ;
        RECT 592.650 39.750 594.450 42.600 ;
        RECT 595.650 39.750 597.450 42.600 ;
        RECT 601.650 39.750 603.450 42.600 ;
        RECT 604.650 39.750 606.450 42.600 ;
        RECT 608.550 39.750 610.350 45.600 ;
        RECT 613.950 44.700 616.050 45.600 ;
        RECT 621.150 45.000 622.950 46.800 ;
        RECT 632.100 46.200 633.150 47.100 ;
        RECT 628.350 45.450 630.150 46.200 ;
        RECT 613.950 43.500 617.700 44.700 ;
        RECT 616.650 42.600 617.700 43.500 ;
        RECT 625.200 44.400 630.150 45.450 ;
        RECT 631.650 44.400 633.450 46.200 ;
        RECT 640.950 45.600 641.850 58.200 ;
        RECT 650.250 57.150 651.450 65.400 ;
        RECT 662.700 59.400 664.500 71.250 ;
        RECT 666.900 59.400 668.700 71.250 ;
        RECT 673.650 65.400 675.450 71.250 ;
        RECT 676.650 65.400 678.450 71.250 ;
        RECT 659.250 57.150 661.050 58.950 ;
        RECT 646.950 53.850 649.050 55.950 ;
        RECT 649.950 55.050 652.050 57.150 ;
        RECT 647.100 52.050 648.900 53.850 ;
        RECT 650.250 47.700 651.450 55.050 ;
        RECT 652.950 53.850 655.050 55.950 ;
        RECT 658.950 55.050 661.050 57.150 ;
        RECT 662.850 54.150 664.050 59.400 ;
        RECT 668.100 54.150 669.900 55.950 ;
        RECT 653.100 52.050 654.900 53.850 ;
        RECT 661.950 52.050 664.050 54.150 ;
        RECT 661.950 48.750 663.150 52.050 ;
        RECT 664.950 50.850 667.050 52.950 ;
        RECT 667.950 52.050 670.050 54.150 ;
        RECT 674.400 52.950 675.600 65.400 ;
        RECT 680.550 59.400 682.350 71.250 ;
        RECT 683.550 68.400 685.350 71.250 ;
        RECT 688.050 65.400 689.850 71.250 ;
        RECT 692.250 65.400 694.050 71.250 ;
        RECT 685.950 63.300 689.850 65.400 ;
        RECT 696.150 64.500 697.950 71.250 ;
        RECT 699.150 65.400 700.950 71.250 ;
        RECT 703.950 65.400 705.750 71.250 ;
        RECT 709.050 65.400 710.850 71.250 ;
        RECT 704.250 64.500 705.450 65.400 ;
        RECT 694.950 62.700 701.850 64.500 ;
        RECT 704.250 62.400 709.050 64.500 ;
        RECT 687.150 60.600 689.850 62.400 ;
        RECT 690.750 61.800 692.550 62.400 ;
        RECT 690.750 60.900 697.050 61.800 ;
        RECT 704.250 61.500 705.450 62.400 ;
        RECT 690.750 60.600 692.550 60.900 ;
        RECT 688.950 59.700 689.850 60.600 ;
        RECT 673.950 50.850 676.050 52.950 ;
        RECT 677.100 51.150 678.900 52.950 ;
        RECT 665.100 49.050 666.900 50.850 ;
        RECT 625.200 42.600 626.250 44.400 ;
        RECT 634.950 43.500 637.050 45.600 ;
        RECT 634.950 42.600 636.000 43.500 ;
        RECT 611.850 39.750 613.650 42.600 ;
        RECT 616.350 39.750 618.150 42.600 ;
        RECT 620.550 39.750 622.350 42.600 ;
        RECT 624.450 39.750 626.250 42.600 ;
        RECT 627.750 39.750 629.550 42.600 ;
        RECT 632.250 41.700 636.000 42.600 ;
        RECT 632.250 39.750 634.050 41.700 ;
        RECT 637.050 39.750 638.850 42.600 ;
        RECT 640.050 39.750 641.850 45.600 ;
        RECT 647.850 46.800 651.450 47.700 ;
        RECT 659.250 47.700 663.000 48.750 ;
        RECT 647.850 39.750 649.650 46.800 ;
        RECT 659.250 45.600 660.450 47.700 ;
        RECT 652.350 39.750 654.150 45.600 ;
        RECT 658.650 39.750 660.450 45.600 ;
        RECT 661.650 44.700 669.450 46.050 ;
        RECT 661.650 39.750 663.450 44.700 ;
        RECT 664.650 39.750 666.450 43.800 ;
        RECT 667.650 39.750 669.450 44.700 ;
        RECT 674.400 42.600 675.600 50.850 ;
        RECT 676.950 49.050 679.050 51.150 ;
        RECT 680.550 49.950 681.750 59.400 ;
        RECT 685.950 58.800 688.050 59.700 ;
        RECT 688.950 58.800 694.950 59.700 ;
        RECT 683.850 57.600 688.050 58.800 ;
        RECT 682.950 55.800 684.750 57.600 ;
        RECT 694.050 54.150 694.950 58.800 ;
        RECT 696.150 58.800 697.050 60.900 ;
        RECT 697.950 60.300 705.450 61.500 ;
        RECT 697.950 59.700 699.750 60.300 ;
        RECT 712.050 59.400 713.850 71.250 ;
        RECT 702.750 58.800 713.850 59.400 ;
        RECT 696.150 58.200 713.850 58.800 ;
        RECT 696.150 57.900 704.550 58.200 ;
        RECT 702.750 57.600 704.550 57.900 ;
        RECT 694.050 52.050 697.050 54.150 ;
        RECT 700.950 53.100 703.050 54.150 ;
        RECT 700.950 52.050 708.900 53.100 ;
        RECT 682.950 51.750 685.050 52.050 ;
        RECT 682.950 49.950 686.850 51.750 ;
        RECT 680.550 47.850 685.050 49.950 ;
        RECT 694.050 48.000 694.950 52.050 ;
        RECT 707.100 51.300 708.900 52.050 ;
        RECT 710.100 51.150 711.900 52.950 ;
        RECT 704.100 50.400 705.900 51.000 ;
        RECT 710.100 50.400 711.000 51.150 ;
        RECT 704.100 49.200 711.000 50.400 ;
        RECT 704.100 48.000 705.150 49.200 ;
        RECT 680.550 45.600 681.750 47.850 ;
        RECT 694.050 47.100 705.150 48.000 ;
        RECT 694.050 46.800 694.950 47.100 ;
        RECT 673.650 39.750 675.450 42.600 ;
        RECT 676.650 39.750 678.450 42.600 ;
        RECT 680.550 39.750 682.350 45.600 ;
        RECT 685.950 44.700 688.050 45.600 ;
        RECT 693.150 45.000 694.950 46.800 ;
        RECT 704.100 46.200 705.150 47.100 ;
        RECT 700.350 45.450 702.150 46.200 ;
        RECT 685.950 43.500 689.700 44.700 ;
        RECT 688.650 42.600 689.700 43.500 ;
        RECT 697.200 44.400 702.150 45.450 ;
        RECT 703.650 44.400 705.450 46.200 ;
        RECT 712.950 45.600 713.850 58.200 ;
        RECT 697.200 42.600 698.250 44.400 ;
        RECT 706.950 43.500 709.050 45.600 ;
        RECT 706.950 42.600 708.000 43.500 ;
        RECT 683.850 39.750 685.650 42.600 ;
        RECT 688.350 39.750 690.150 42.600 ;
        RECT 692.550 39.750 694.350 42.600 ;
        RECT 696.450 39.750 698.250 42.600 ;
        RECT 699.750 39.750 701.550 42.600 ;
        RECT 704.250 41.700 708.000 42.600 ;
        RECT 704.250 39.750 706.050 41.700 ;
        RECT 709.050 39.750 710.850 42.600 ;
        RECT 712.050 39.750 713.850 45.600 ;
        RECT 8.100 27.000 9.900 35.250 ;
        RECT 5.400 25.350 9.900 27.000 ;
        RECT 13.500 26.400 15.300 35.250 ;
        RECT 18.000 29.400 19.800 35.250 ;
        RECT 22.200 31.050 24.000 35.250 ;
        RECT 25.500 32.400 27.300 35.250 ;
        RECT 22.200 29.400 27.900 31.050 ;
        RECT 34.650 29.400 36.450 35.250 ;
        RECT 5.400 21.150 6.600 25.350 ;
        RECT 17.100 24.150 18.900 25.950 ;
        RECT 16.950 22.050 19.050 24.150 ;
        RECT 19.950 23.850 22.050 25.950 ;
        RECT 23.100 24.150 24.900 25.950 ;
        RECT 20.100 22.050 21.900 23.850 ;
        RECT 22.950 22.050 25.050 24.150 ;
        RECT 26.700 22.950 27.900 29.400 ;
        RECT 35.250 27.300 36.450 29.400 ;
        RECT 37.650 30.300 39.450 35.250 ;
        RECT 40.650 31.200 42.450 35.250 ;
        RECT 43.650 30.300 45.450 35.250 ;
        RECT 37.650 28.950 45.450 30.300 ;
        RECT 47.550 30.300 49.350 35.250 ;
        RECT 50.550 31.200 52.350 35.250 ;
        RECT 53.550 30.300 55.350 35.250 ;
        RECT 47.550 28.950 55.350 30.300 ;
        RECT 56.550 29.400 58.350 35.250 ;
        RECT 56.550 27.300 57.750 29.400 ;
        RECT 35.250 26.250 39.000 27.300 ;
        RECT 54.000 26.250 57.750 27.300 ;
        RECT 68.100 27.000 69.900 35.250 ;
        RECT 37.950 22.950 39.150 26.250 ;
        RECT 41.100 24.150 42.900 25.950 ;
        RECT 50.100 24.150 51.900 25.950 ;
        RECT 4.950 19.050 7.050 21.150 ;
        RECT 25.950 20.850 28.050 22.950 ;
        RECT 37.950 20.850 40.050 22.950 ;
        RECT 40.950 22.050 43.050 24.150 ;
        RECT 43.950 20.850 46.050 22.950 ;
        RECT 46.950 20.850 49.050 22.950 ;
        RECT 49.950 22.050 52.050 24.150 ;
        RECT 53.850 22.950 55.050 26.250 ;
        RECT 52.950 20.850 55.050 22.950 ;
        RECT 65.400 25.350 69.900 27.000 ;
        RECT 73.500 26.400 75.300 35.250 ;
        RECT 77.700 26.400 79.500 35.250 ;
        RECT 83.100 27.000 84.900 35.250 ;
        RECT 93.000 29.400 94.800 35.250 ;
        RECT 97.200 31.050 99.000 35.250 ;
        RECT 100.500 32.400 102.300 35.250 ;
        RECT 110.700 32.400 112.500 35.250 ;
        RECT 114.000 31.050 115.800 35.250 ;
        RECT 97.200 29.400 102.900 31.050 ;
        RECT 83.100 25.350 87.600 27.000 ;
        RECT 88.950 25.950 91.050 28.050 ;
        RECT 65.400 21.150 66.600 25.350 ;
        RECT 86.400 21.150 87.600 25.350 ;
        RECT 5.250 10.800 6.300 19.050 ;
        RECT 7.950 17.850 10.050 19.950 ;
        RECT 13.950 17.850 16.050 19.950 ;
        RECT 7.950 16.050 9.750 17.850 ;
        RECT 10.950 14.850 13.050 16.950 ;
        RECT 14.100 16.050 15.900 17.850 ;
        RECT 26.700 15.600 27.900 20.850 ;
        RECT 34.950 17.850 37.050 19.950 ;
        RECT 35.250 16.050 37.050 17.850 ;
        RECT 38.850 15.600 40.050 20.850 ;
        RECT 44.100 19.050 45.900 20.850 ;
        RECT 47.100 19.050 48.900 20.850 ;
        RECT 52.950 15.600 54.150 20.850 ;
        RECT 55.950 17.850 58.050 19.950 ;
        RECT 64.950 19.050 67.050 21.150 ;
        RECT 55.950 16.050 57.750 17.850 ;
        RECT 11.100 13.050 12.900 14.850 ;
        RECT 17.550 14.700 25.350 15.600 ;
        RECT 5.250 9.900 12.300 10.800 ;
        RECT 5.250 9.600 6.450 9.900 ;
        RECT 4.650 3.750 6.450 9.600 ;
        RECT 10.650 9.600 12.300 9.900 ;
        RECT 7.650 3.750 9.450 9.000 ;
        RECT 10.650 3.750 12.450 9.600 ;
        RECT 13.650 3.750 15.450 9.600 ;
        RECT 17.550 3.750 19.350 14.700 ;
        RECT 20.550 3.750 22.350 13.800 ;
        RECT 23.550 3.750 25.350 14.700 ;
        RECT 26.550 3.750 28.350 15.600 ;
        RECT 35.400 3.750 37.200 9.600 ;
        RECT 38.700 3.750 40.500 15.600 ;
        RECT 42.900 3.750 44.700 15.600 ;
        RECT 48.300 3.750 50.100 15.600 ;
        RECT 52.500 3.750 54.300 15.600 ;
        RECT 65.250 10.800 66.300 19.050 ;
        RECT 67.950 17.850 70.050 19.950 ;
        RECT 73.950 17.850 76.050 19.950 ;
        RECT 76.950 17.850 79.050 19.950 ;
        RECT 82.950 17.850 85.050 19.950 ;
        RECT 85.950 19.050 88.050 21.150 ;
        RECT 67.950 16.050 69.750 17.850 ;
        RECT 70.950 14.850 73.050 16.950 ;
        RECT 74.100 16.050 75.900 17.850 ;
        RECT 77.100 16.050 78.900 17.850 ;
        RECT 79.950 14.850 82.050 16.950 ;
        RECT 83.250 16.050 85.050 17.850 ;
        RECT 71.100 13.050 72.900 14.850 ;
        RECT 80.100 13.050 81.900 14.850 ;
        RECT 86.700 10.800 87.750 19.050 ;
        RECT 89.550 16.050 90.450 25.950 ;
        RECT 92.100 24.150 93.900 25.950 ;
        RECT 91.950 22.050 94.050 24.150 ;
        RECT 94.950 23.850 97.050 25.950 ;
        RECT 98.100 24.150 99.900 25.950 ;
        RECT 95.100 22.050 96.900 23.850 ;
        RECT 97.950 22.050 100.050 24.150 ;
        RECT 101.700 22.950 102.900 29.400 ;
        RECT 110.100 29.400 115.800 31.050 ;
        RECT 118.200 29.400 120.000 35.250 ;
        RECT 122.550 32.400 124.350 35.250 ;
        RECT 125.550 32.400 127.350 35.250 ;
        RECT 110.100 22.950 111.300 29.400 ;
        RECT 113.100 24.150 114.900 25.950 ;
        RECT 100.950 20.850 103.050 22.950 ;
        RECT 109.950 20.850 112.050 22.950 ;
        RECT 112.950 22.050 115.050 24.150 ;
        RECT 115.950 23.850 118.050 25.950 ;
        RECT 119.100 24.150 120.900 25.950 ;
        RECT 116.100 22.050 117.900 23.850 ;
        RECT 118.950 22.050 121.050 24.150 ;
        RECT 121.950 23.850 124.050 25.950 ;
        RECT 125.400 24.150 126.600 32.400 ;
        RECT 133.650 29.400 135.450 35.250 ;
        RECT 134.250 27.300 135.450 29.400 ;
        RECT 136.650 30.300 138.450 35.250 ;
        RECT 139.650 31.200 141.450 35.250 ;
        RECT 142.650 30.300 144.450 35.250 ;
        RECT 148.650 32.400 150.450 35.250 ;
        RECT 151.650 32.400 153.450 35.250 ;
        RECT 136.650 28.950 144.450 30.300 ;
        RECT 134.250 26.250 138.000 27.300 ;
        RECT 122.100 22.050 123.900 23.850 ;
        RECT 124.950 22.050 127.050 24.150 ;
        RECT 136.950 22.950 138.150 26.250 ;
        RECT 140.100 24.150 141.900 25.950 ;
        RECT 149.400 24.150 150.600 32.400 ;
        RECT 155.550 30.300 157.350 35.250 ;
        RECT 158.550 31.200 160.350 35.250 ;
        RECT 161.550 30.300 163.350 35.250 ;
        RECT 155.550 28.950 163.350 30.300 ;
        RECT 164.550 29.400 166.350 35.250 ;
        RECT 170.550 30.300 172.350 35.250 ;
        RECT 173.550 31.200 175.350 35.250 ;
        RECT 176.550 30.300 178.350 35.250 ;
        RECT 164.550 27.300 165.750 29.400 ;
        RECT 170.550 28.950 178.350 30.300 ;
        RECT 179.550 29.400 181.350 35.250 ;
        RECT 179.550 27.300 180.750 29.400 ;
        RECT 162.000 26.250 165.750 27.300 ;
        RECT 177.000 26.250 180.750 27.300 ;
        RECT 185.700 26.400 187.500 35.250 ;
        RECT 191.100 27.000 192.900 35.250 ;
        RECT 88.950 13.950 91.050 16.050 ;
        RECT 101.700 15.600 102.900 20.850 ;
        RECT 110.100 15.600 111.300 20.850 ;
        RECT 92.550 14.700 100.350 15.600 ;
        RECT 65.250 9.900 72.300 10.800 ;
        RECT 65.250 9.600 66.450 9.900 ;
        RECT 55.800 3.750 57.600 9.600 ;
        RECT 64.650 3.750 66.450 9.600 ;
        RECT 70.650 9.600 72.300 9.900 ;
        RECT 80.700 9.900 87.750 10.800 ;
        RECT 80.700 9.600 82.350 9.900 ;
        RECT 67.650 3.750 69.450 9.000 ;
        RECT 70.650 3.750 72.450 9.600 ;
        RECT 73.650 3.750 75.450 9.600 ;
        RECT 77.550 3.750 79.350 9.600 ;
        RECT 80.550 3.750 82.350 9.600 ;
        RECT 86.550 9.600 87.750 9.900 ;
        RECT 83.550 3.750 85.350 9.000 ;
        RECT 86.550 3.750 88.350 9.600 ;
        RECT 92.550 3.750 94.350 14.700 ;
        RECT 95.550 3.750 97.350 13.800 ;
        RECT 98.550 3.750 100.350 14.700 ;
        RECT 101.550 3.750 103.350 15.600 ;
        RECT 109.650 3.750 111.450 15.600 ;
        RECT 112.650 14.700 120.450 15.600 ;
        RECT 112.650 3.750 114.450 14.700 ;
        RECT 115.650 3.750 117.450 13.800 ;
        RECT 118.650 3.750 120.450 14.700 ;
        RECT 125.400 9.600 126.600 22.050 ;
        RECT 136.950 20.850 139.050 22.950 ;
        RECT 139.950 22.050 142.050 24.150 ;
        RECT 142.950 20.850 145.050 22.950 ;
        RECT 148.950 22.050 151.050 24.150 ;
        RECT 151.950 23.850 154.050 25.950 ;
        RECT 158.100 24.150 159.900 25.950 ;
        RECT 152.100 22.050 153.900 23.850 ;
        RECT 133.950 17.850 136.050 19.950 ;
        RECT 134.250 16.050 136.050 17.850 ;
        RECT 137.850 15.600 139.050 20.850 ;
        RECT 143.100 19.050 144.900 20.850 ;
        RECT 122.550 3.750 124.350 9.600 ;
        RECT 125.550 3.750 127.350 9.600 ;
        RECT 134.400 3.750 136.200 9.600 ;
        RECT 137.700 3.750 139.500 15.600 ;
        RECT 141.900 3.750 143.700 15.600 ;
        RECT 149.400 9.600 150.600 22.050 ;
        RECT 154.950 20.850 157.050 22.950 ;
        RECT 157.950 22.050 160.050 24.150 ;
        RECT 161.850 22.950 163.050 26.250 ;
        RECT 173.100 24.150 174.900 25.950 ;
        RECT 160.950 20.850 163.050 22.950 ;
        RECT 169.950 20.850 172.050 22.950 ;
        RECT 172.950 22.050 175.050 24.150 ;
        RECT 176.850 22.950 178.050 26.250 ;
        RECT 191.100 25.350 195.600 27.000 ;
        RECT 200.700 26.400 202.500 35.250 ;
        RECT 206.100 27.000 207.900 35.250 ;
        RECT 218.700 32.400 220.500 35.250 ;
        RECT 222.000 31.050 223.800 35.250 ;
        RECT 218.100 29.400 223.800 31.050 ;
        RECT 226.200 29.400 228.000 35.250 ;
        RECT 206.100 25.350 210.600 27.000 ;
        RECT 175.950 20.850 178.050 22.950 ;
        RECT 194.400 21.150 195.600 25.350 ;
        RECT 209.400 21.150 210.600 25.350 ;
        RECT 218.100 22.950 219.300 29.400 ;
        RECT 230.700 26.400 232.500 35.250 ;
        RECT 236.100 27.000 237.900 35.250 ;
        RECT 248.700 32.400 250.500 35.250 ;
        RECT 252.000 31.050 253.800 35.250 ;
        RECT 248.100 29.400 253.800 31.050 ;
        RECT 256.200 29.400 258.000 35.250 ;
        RECT 221.100 24.150 222.900 25.950 ;
        RECT 155.100 19.050 156.900 20.850 ;
        RECT 160.950 15.600 162.150 20.850 ;
        RECT 163.950 17.850 166.050 19.950 ;
        RECT 170.100 19.050 171.900 20.850 ;
        RECT 163.950 16.050 165.750 17.850 ;
        RECT 175.950 15.600 177.150 20.850 ;
        RECT 178.950 17.850 181.050 19.950 ;
        RECT 184.950 17.850 187.050 19.950 ;
        RECT 190.950 17.850 193.050 19.950 ;
        RECT 193.950 19.050 196.050 21.150 ;
        RECT 178.950 16.050 180.750 17.850 ;
        RECT 185.100 16.050 186.900 17.850 ;
        RECT 148.650 3.750 150.450 9.600 ;
        RECT 151.650 3.750 153.450 9.600 ;
        RECT 156.300 3.750 158.100 15.600 ;
        RECT 160.500 3.750 162.300 15.600 ;
        RECT 163.800 3.750 165.600 9.600 ;
        RECT 171.300 3.750 173.100 15.600 ;
        RECT 175.500 3.750 177.300 15.600 ;
        RECT 187.950 14.850 190.050 16.950 ;
        RECT 191.250 16.050 193.050 17.850 ;
        RECT 188.100 13.050 189.900 14.850 ;
        RECT 194.700 10.800 195.750 19.050 ;
        RECT 199.950 17.850 202.050 19.950 ;
        RECT 205.950 17.850 208.050 19.950 ;
        RECT 208.950 19.050 211.050 21.150 ;
        RECT 217.950 20.850 220.050 22.950 ;
        RECT 220.950 22.050 223.050 24.150 ;
        RECT 223.950 23.850 226.050 25.950 ;
        RECT 227.100 24.150 228.900 25.950 ;
        RECT 236.100 25.350 240.600 27.000 ;
        RECT 224.100 22.050 225.900 23.850 ;
        RECT 226.950 22.050 229.050 24.150 ;
        RECT 239.400 21.150 240.600 25.350 ;
        RECT 248.100 22.950 249.300 29.400 ;
        RECT 260.700 26.400 262.500 35.250 ;
        RECT 266.100 27.000 267.900 35.250 ;
        RECT 275.850 29.400 277.650 35.250 ;
        RECT 280.350 28.200 282.150 35.250 ;
        RECT 287.550 32.400 289.350 35.250 ;
        RECT 278.550 27.300 282.150 28.200 ;
        RECT 288.150 28.500 289.350 32.400 ;
        RECT 290.850 29.400 292.650 35.250 ;
        RECT 293.850 29.400 295.650 35.250 ;
        RECT 303.150 30.900 304.950 35.250 ;
        RECT 301.650 29.400 304.950 30.900 ;
        RECT 306.150 29.400 307.950 35.250 ;
        RECT 288.150 27.600 293.250 28.500 ;
        RECT 251.100 24.150 252.900 25.950 ;
        RECT 200.100 16.050 201.900 17.850 ;
        RECT 202.950 14.850 205.050 16.950 ;
        RECT 206.250 16.050 208.050 17.850 ;
        RECT 203.100 13.050 204.900 14.850 ;
        RECT 209.700 10.800 210.750 19.050 ;
        RECT 218.100 15.600 219.300 20.850 ;
        RECT 229.950 17.850 232.050 19.950 ;
        RECT 235.950 17.850 238.050 19.950 ;
        RECT 238.950 19.050 241.050 21.150 ;
        RECT 247.950 20.850 250.050 22.950 ;
        RECT 250.950 22.050 253.050 24.150 ;
        RECT 253.950 23.850 256.050 25.950 ;
        RECT 257.100 24.150 258.900 25.950 ;
        RECT 266.100 25.350 270.600 27.000 ;
        RECT 254.100 22.050 255.900 23.850 ;
        RECT 256.950 22.050 259.050 24.150 ;
        RECT 269.400 21.150 270.600 25.350 ;
        RECT 275.100 21.150 276.900 22.950 ;
        RECT 230.100 16.050 231.900 17.850 ;
        RECT 188.700 9.900 195.750 10.800 ;
        RECT 188.700 9.600 190.350 9.900 ;
        RECT 178.800 3.750 180.600 9.600 ;
        RECT 185.550 3.750 187.350 9.600 ;
        RECT 188.550 3.750 190.350 9.600 ;
        RECT 194.550 9.600 195.750 9.900 ;
        RECT 203.700 9.900 210.750 10.800 ;
        RECT 203.700 9.600 205.350 9.900 ;
        RECT 191.550 3.750 193.350 9.000 ;
        RECT 194.550 3.750 196.350 9.600 ;
        RECT 200.550 3.750 202.350 9.600 ;
        RECT 203.550 3.750 205.350 9.600 ;
        RECT 209.550 9.600 210.750 9.900 ;
        RECT 206.550 3.750 208.350 9.000 ;
        RECT 209.550 3.750 211.350 9.600 ;
        RECT 217.650 3.750 219.450 15.600 ;
        RECT 220.650 14.700 228.450 15.600 ;
        RECT 232.950 14.850 235.050 16.950 ;
        RECT 236.250 16.050 238.050 17.850 ;
        RECT 220.650 3.750 222.450 14.700 ;
        RECT 223.650 3.750 225.450 13.800 ;
        RECT 226.650 3.750 228.450 14.700 ;
        RECT 233.100 13.050 234.900 14.850 ;
        RECT 239.700 10.800 240.750 19.050 ;
        RECT 248.100 15.600 249.300 20.850 ;
        RECT 259.950 17.850 262.050 19.950 ;
        RECT 265.950 17.850 268.050 19.950 ;
        RECT 268.950 19.050 271.050 21.150 ;
        RECT 274.950 19.050 277.050 21.150 ;
        RECT 278.550 19.950 279.750 27.300 ;
        RECT 291.000 26.700 293.250 27.600 ;
        RECT 281.100 21.150 282.900 22.950 ;
        RECT 260.100 16.050 261.900 17.850 ;
        RECT 233.700 9.900 240.750 10.800 ;
        RECT 233.700 9.600 235.350 9.900 ;
        RECT 230.550 3.750 232.350 9.600 ;
        RECT 233.550 3.750 235.350 9.600 ;
        RECT 239.550 9.600 240.750 9.900 ;
        RECT 236.550 3.750 238.350 9.000 ;
        RECT 239.550 3.750 241.350 9.600 ;
        RECT 247.650 3.750 249.450 15.600 ;
        RECT 250.650 14.700 258.450 15.600 ;
        RECT 262.950 14.850 265.050 16.950 ;
        RECT 266.250 16.050 268.050 17.850 ;
        RECT 250.650 3.750 252.450 14.700 ;
        RECT 253.650 3.750 255.450 13.800 ;
        RECT 256.650 3.750 258.450 14.700 ;
        RECT 263.100 13.050 264.900 14.850 ;
        RECT 269.700 10.800 270.750 19.050 ;
        RECT 277.950 17.850 280.050 19.950 ;
        RECT 280.950 19.050 283.050 21.150 ;
        RECT 286.950 20.850 289.050 22.950 ;
        RECT 287.100 19.050 288.900 20.850 ;
        RECT 291.000 18.300 292.050 26.700 ;
        RECT 294.150 22.950 295.350 29.400 ;
        RECT 292.950 20.850 295.350 22.950 ;
        RECT 263.700 9.900 270.750 10.800 ;
        RECT 263.700 9.600 265.350 9.900 ;
        RECT 260.550 3.750 262.350 9.600 ;
        RECT 263.550 3.750 265.350 9.600 ;
        RECT 269.550 9.600 270.750 9.900 ;
        RECT 278.550 9.600 279.750 17.850 ;
        RECT 291.000 17.400 293.250 18.300 ;
        RECT 287.550 16.500 293.250 17.400 ;
        RECT 287.550 9.600 288.750 16.500 ;
        RECT 294.150 15.600 295.350 20.850 ;
        RECT 301.650 22.950 302.850 29.400 ;
        RECT 304.950 27.900 306.750 28.500 ;
        RECT 310.650 27.900 312.450 35.250 ;
        RECT 314.550 32.400 316.350 35.250 ;
        RECT 304.950 26.700 312.450 27.900 ;
        RECT 315.150 28.500 316.350 32.400 ;
        RECT 317.850 29.400 319.650 35.250 ;
        RECT 320.850 29.400 322.650 35.250 ;
        RECT 315.150 27.600 320.250 28.500 ;
        RECT 318.000 26.700 320.250 27.600 ;
        RECT 301.650 20.850 304.050 22.950 ;
        RECT 305.100 21.150 306.900 22.950 ;
        RECT 301.650 15.600 302.850 20.850 ;
        RECT 304.950 19.050 307.050 21.150 ;
        RECT 266.550 3.750 268.350 9.000 ;
        RECT 269.550 3.750 271.350 9.600 ;
        RECT 275.550 3.750 277.350 9.600 ;
        RECT 278.550 3.750 280.350 9.600 ;
        RECT 281.550 3.750 283.350 9.600 ;
        RECT 287.550 3.750 289.350 9.600 ;
        RECT 290.850 3.750 292.650 15.600 ;
        RECT 293.850 3.750 295.650 15.600 ;
        RECT 301.050 3.750 302.850 15.600 ;
        RECT 304.050 3.750 305.850 15.600 ;
        RECT 308.100 9.600 309.300 26.700 ;
        RECT 310.950 20.850 313.050 22.950 ;
        RECT 313.950 20.850 316.050 22.950 ;
        RECT 311.100 19.050 312.900 20.850 ;
        RECT 314.100 19.050 315.900 20.850 ;
        RECT 318.000 18.300 319.050 26.700 ;
        RECT 321.150 22.950 322.350 29.400 ;
        RECT 326.700 26.400 328.500 35.250 ;
        RECT 332.100 27.000 333.900 35.250 ;
        RECT 342.000 29.400 343.800 35.250 ;
        RECT 346.200 29.400 348.000 35.250 ;
        RECT 350.400 29.400 352.200 35.250 ;
        RECT 359.550 30.300 361.350 35.250 ;
        RECT 362.550 31.200 364.350 35.250 ;
        RECT 365.550 30.300 367.350 35.250 ;
        RECT 332.100 25.350 336.600 27.000 ;
        RECT 319.950 20.850 322.350 22.950 ;
        RECT 335.400 21.150 336.600 25.350 ;
        RECT 344.250 24.150 346.050 25.950 ;
        RECT 318.000 17.400 320.250 18.300 ;
        RECT 314.550 16.500 320.250 17.400 ;
        RECT 314.550 9.600 315.750 16.500 ;
        RECT 321.150 15.600 322.350 20.850 ;
        RECT 325.950 17.850 328.050 19.950 ;
        RECT 331.950 17.850 334.050 19.950 ;
        RECT 334.950 19.050 337.050 21.150 ;
        RECT 340.950 20.850 343.050 22.950 ;
        RECT 343.950 22.050 346.050 24.150 ;
        RECT 346.950 22.950 348.000 29.400 ;
        RECT 359.550 28.950 367.350 30.300 ;
        RECT 368.550 29.400 370.350 35.250 ;
        RECT 377.700 32.400 379.500 35.250 ;
        RECT 381.000 31.050 382.800 35.250 ;
        RECT 377.100 29.400 382.800 31.050 ;
        RECT 385.200 29.400 387.000 35.250 ;
        RECT 389.550 30.300 391.350 35.250 ;
        RECT 392.550 31.200 394.350 35.250 ;
        RECT 395.550 30.300 397.350 35.250 ;
        RECT 368.550 27.300 369.750 29.400 ;
        RECT 366.000 26.250 369.750 27.300 ;
        RECT 349.950 24.150 351.750 25.950 ;
        RECT 362.100 24.150 363.900 25.950 ;
        RECT 346.950 20.850 349.050 22.950 ;
        RECT 349.950 22.050 352.050 24.150 ;
        RECT 352.950 20.850 355.050 22.950 ;
        RECT 358.950 20.850 361.050 22.950 ;
        RECT 361.950 22.050 364.050 24.150 ;
        RECT 365.850 22.950 367.050 26.250 ;
        RECT 377.100 22.950 378.300 29.400 ;
        RECT 389.550 28.950 397.350 30.300 ;
        RECT 398.550 29.400 400.350 35.250 ;
        RECT 404.550 32.400 406.350 35.250 ;
        RECT 407.550 32.400 409.350 35.250 ;
        RECT 398.550 27.300 399.750 29.400 ;
        RECT 396.000 26.250 399.750 27.300 ;
        RECT 380.100 24.150 381.900 25.950 ;
        RECT 364.950 20.850 367.050 22.950 ;
        RECT 376.950 20.850 379.050 22.950 ;
        RECT 379.950 22.050 382.050 24.150 ;
        RECT 382.950 23.850 385.050 25.950 ;
        RECT 386.100 24.150 387.900 25.950 ;
        RECT 392.100 24.150 393.900 25.950 ;
        RECT 383.100 22.050 384.900 23.850 ;
        RECT 385.950 22.050 388.050 24.150 ;
        RECT 388.950 20.850 391.050 22.950 ;
        RECT 391.950 22.050 394.050 24.150 ;
        RECT 395.850 22.950 397.050 26.250 ;
        RECT 403.950 23.850 406.050 25.950 ;
        RECT 407.400 24.150 408.600 32.400 ;
        RECT 413.700 26.400 415.500 35.250 ;
        RECT 419.100 27.000 420.900 35.250 ;
        RECT 428.550 32.400 430.350 35.250 ;
        RECT 431.550 32.400 433.350 35.250 ;
        RECT 419.100 25.350 423.600 27.000 ;
        RECT 394.950 20.850 397.050 22.950 ;
        RECT 404.100 22.050 405.900 23.850 ;
        RECT 406.950 22.050 409.050 24.150 ;
        RECT 341.250 19.050 343.050 20.850 ;
        RECT 326.100 16.050 327.900 17.850 ;
        RECT 307.650 3.750 309.450 9.600 ;
        RECT 310.650 3.750 312.450 9.600 ;
        RECT 314.550 3.750 316.350 9.600 ;
        RECT 317.850 3.750 319.650 15.600 ;
        RECT 320.850 3.750 322.650 15.600 ;
        RECT 328.950 14.850 331.050 16.950 ;
        RECT 332.250 16.050 334.050 17.850 ;
        RECT 329.100 13.050 330.900 14.850 ;
        RECT 335.700 10.800 336.750 19.050 ;
        RECT 348.150 17.400 349.050 20.850 ;
        RECT 353.100 19.050 354.900 20.850 ;
        RECT 359.100 19.050 360.900 20.850 ;
        RECT 348.150 16.500 352.200 17.400 ;
        RECT 350.400 15.600 352.200 16.500 ;
        RECT 364.950 15.600 366.150 20.850 ;
        RECT 367.950 17.850 370.050 19.950 ;
        RECT 367.950 16.050 369.750 17.850 ;
        RECT 377.100 15.600 378.300 20.850 ;
        RECT 389.100 19.050 390.900 20.850 ;
        RECT 394.950 15.600 396.150 20.850 ;
        RECT 397.950 17.850 400.050 19.950 ;
        RECT 397.950 16.050 399.750 17.850 ;
        RECT 329.700 9.900 336.750 10.800 ;
        RECT 329.700 9.600 331.350 9.900 ;
        RECT 326.550 3.750 328.350 9.600 ;
        RECT 329.550 3.750 331.350 9.600 ;
        RECT 335.550 9.600 336.750 9.900 ;
        RECT 341.550 14.400 349.350 15.300 ;
        RECT 332.550 3.750 334.350 9.000 ;
        RECT 335.550 3.750 337.350 9.600 ;
        RECT 341.550 3.750 343.350 14.400 ;
        RECT 344.550 3.750 346.350 13.500 ;
        RECT 347.550 4.500 349.350 14.400 ;
        RECT 350.550 5.400 352.350 15.600 ;
        RECT 353.550 4.500 355.350 15.600 ;
        RECT 347.550 3.750 355.350 4.500 ;
        RECT 360.300 3.750 362.100 15.600 ;
        RECT 364.500 3.750 366.300 15.600 ;
        RECT 367.800 3.750 369.600 9.600 ;
        RECT 376.650 3.750 378.450 15.600 ;
        RECT 379.650 14.700 387.450 15.600 ;
        RECT 379.650 3.750 381.450 14.700 ;
        RECT 382.650 3.750 384.450 13.800 ;
        RECT 385.650 3.750 387.450 14.700 ;
        RECT 390.300 3.750 392.100 15.600 ;
        RECT 394.500 3.750 396.300 15.600 ;
        RECT 407.400 9.600 408.600 22.050 ;
        RECT 422.400 21.150 423.600 25.350 ;
        RECT 427.950 23.850 430.050 25.950 ;
        RECT 431.400 24.150 432.600 32.400 ;
        RECT 438.150 29.400 439.950 35.250 ;
        RECT 441.150 32.400 442.950 35.250 ;
        RECT 445.950 33.300 447.750 35.250 ;
        RECT 444.000 32.400 447.750 33.300 ;
        RECT 450.450 32.400 452.250 35.250 ;
        RECT 453.750 32.400 455.550 35.250 ;
        RECT 457.650 32.400 459.450 35.250 ;
        RECT 461.850 32.400 463.650 35.250 ;
        RECT 466.350 32.400 468.150 35.250 ;
        RECT 444.000 31.500 445.050 32.400 ;
        RECT 442.950 29.400 445.050 31.500 ;
        RECT 453.750 30.600 454.800 32.400 ;
        RECT 428.100 22.050 429.900 23.850 ;
        RECT 430.950 22.050 433.050 24.150 ;
        RECT 412.950 17.850 415.050 19.950 ;
        RECT 418.950 17.850 421.050 19.950 ;
        RECT 421.950 19.050 424.050 21.150 ;
        RECT 413.100 16.050 414.900 17.850 ;
        RECT 415.950 14.850 418.050 16.950 ;
        RECT 419.250 16.050 421.050 17.850 ;
        RECT 416.100 13.050 417.900 14.850 ;
        RECT 422.700 10.800 423.750 19.050 ;
        RECT 416.700 9.900 423.750 10.800 ;
        RECT 416.700 9.600 418.350 9.900 ;
        RECT 397.800 3.750 399.600 9.600 ;
        RECT 404.550 3.750 406.350 9.600 ;
        RECT 407.550 3.750 409.350 9.600 ;
        RECT 413.550 3.750 415.350 9.600 ;
        RECT 416.550 3.750 418.350 9.600 ;
        RECT 422.550 9.600 423.750 9.900 ;
        RECT 431.400 9.600 432.600 22.050 ;
        RECT 438.150 16.800 439.050 29.400 ;
        RECT 446.550 28.800 448.350 30.600 ;
        RECT 449.850 29.550 454.800 30.600 ;
        RECT 462.300 31.500 463.350 32.400 ;
        RECT 462.300 30.300 466.050 31.500 ;
        RECT 449.850 28.800 451.650 29.550 ;
        RECT 446.850 27.900 447.900 28.800 ;
        RECT 457.050 28.200 458.850 30.000 ;
        RECT 463.950 29.400 466.050 30.300 ;
        RECT 469.650 29.400 471.450 35.250 ;
        RECT 473.550 32.400 475.350 35.250 ;
        RECT 476.550 32.400 478.350 35.250 ;
        RECT 484.650 32.400 486.450 35.250 ;
        RECT 487.650 32.400 489.450 35.250 ;
        RECT 457.050 27.900 457.950 28.200 ;
        RECT 446.850 27.000 457.950 27.900 ;
        RECT 470.250 27.150 471.450 29.400 ;
        RECT 446.850 25.800 447.900 27.000 ;
        RECT 441.000 24.600 447.900 25.800 ;
        RECT 441.000 23.850 441.900 24.600 ;
        RECT 446.100 24.000 447.900 24.600 ;
        RECT 440.100 22.050 441.900 23.850 ;
        RECT 443.100 22.950 444.900 23.700 ;
        RECT 457.050 22.950 457.950 27.000 ;
        RECT 466.950 25.050 471.450 27.150 ;
        RECT 465.150 23.250 469.050 25.050 ;
        RECT 466.950 22.950 469.050 23.250 ;
        RECT 443.100 21.900 451.050 22.950 ;
        RECT 448.950 20.850 451.050 21.900 ;
        RECT 454.950 20.850 457.950 22.950 ;
        RECT 447.450 17.100 449.250 17.400 ;
        RECT 447.450 16.800 455.850 17.100 ;
        RECT 438.150 16.200 455.850 16.800 ;
        RECT 438.150 15.600 449.250 16.200 ;
        RECT 419.550 3.750 421.350 9.000 ;
        RECT 422.550 3.750 424.350 9.600 ;
        RECT 428.550 3.750 430.350 9.600 ;
        RECT 431.550 3.750 433.350 9.600 ;
        RECT 438.150 3.750 439.950 15.600 ;
        RECT 452.250 14.700 454.050 15.300 ;
        RECT 446.550 13.500 454.050 14.700 ;
        RECT 454.950 14.100 455.850 16.200 ;
        RECT 457.050 16.200 457.950 20.850 ;
        RECT 467.250 17.400 469.050 19.200 ;
        RECT 463.950 16.200 468.150 17.400 ;
        RECT 457.050 15.300 463.050 16.200 ;
        RECT 463.950 15.300 466.050 16.200 ;
        RECT 470.250 15.600 471.450 25.050 ;
        RECT 472.950 23.850 475.050 25.950 ;
        RECT 476.400 24.150 477.600 32.400 ;
        RECT 485.400 24.150 486.600 32.400 ;
        RECT 492.150 29.400 493.950 35.250 ;
        RECT 495.150 32.400 496.950 35.250 ;
        RECT 499.950 33.300 501.750 35.250 ;
        RECT 498.000 32.400 501.750 33.300 ;
        RECT 504.450 32.400 506.250 35.250 ;
        RECT 507.750 32.400 509.550 35.250 ;
        RECT 511.650 32.400 513.450 35.250 ;
        RECT 515.850 32.400 517.650 35.250 ;
        RECT 520.350 32.400 522.150 35.250 ;
        RECT 498.000 31.500 499.050 32.400 ;
        RECT 496.950 29.400 499.050 31.500 ;
        RECT 507.750 30.600 508.800 32.400 ;
        RECT 473.100 22.050 474.900 23.850 ;
        RECT 475.950 22.050 478.050 24.150 ;
        RECT 484.950 22.050 487.050 24.150 ;
        RECT 487.950 23.850 490.050 25.950 ;
        RECT 488.100 22.050 489.900 23.850 ;
        RECT 462.150 14.400 463.050 15.300 ;
        RECT 459.450 14.100 461.250 14.400 ;
        RECT 446.550 12.600 447.750 13.500 ;
        RECT 454.950 13.200 461.250 14.100 ;
        RECT 459.450 12.600 461.250 13.200 ;
        RECT 462.150 12.600 464.850 14.400 ;
        RECT 442.950 10.500 447.750 12.600 ;
        RECT 450.150 10.500 457.050 12.300 ;
        RECT 446.550 9.600 447.750 10.500 ;
        RECT 441.150 3.750 442.950 9.600 ;
        RECT 446.250 3.750 448.050 9.600 ;
        RECT 451.050 3.750 452.850 9.600 ;
        RECT 454.050 3.750 455.850 10.500 ;
        RECT 462.150 9.600 466.050 11.700 ;
        RECT 457.950 3.750 459.750 9.600 ;
        RECT 462.150 3.750 463.950 9.600 ;
        RECT 466.650 3.750 468.450 6.600 ;
        RECT 469.650 3.750 471.450 15.600 ;
        RECT 476.400 9.600 477.600 22.050 ;
        RECT 485.400 9.600 486.600 22.050 ;
        RECT 492.150 16.800 493.050 29.400 ;
        RECT 500.550 28.800 502.350 30.600 ;
        RECT 503.850 29.550 508.800 30.600 ;
        RECT 516.300 31.500 517.350 32.400 ;
        RECT 516.300 30.300 520.050 31.500 ;
        RECT 503.850 28.800 505.650 29.550 ;
        RECT 500.850 27.900 501.900 28.800 ;
        RECT 511.050 28.200 512.850 30.000 ;
        RECT 517.950 29.400 520.050 30.300 ;
        RECT 523.650 29.400 525.450 35.250 ;
        RECT 529.650 32.400 531.450 35.250 ;
        RECT 532.650 32.400 534.450 35.250 ;
        RECT 535.650 32.400 537.450 35.250 ;
        RECT 511.050 27.900 511.950 28.200 ;
        RECT 500.850 27.000 511.950 27.900 ;
        RECT 524.250 27.150 525.450 29.400 ;
        RECT 500.850 25.800 501.900 27.000 ;
        RECT 495.000 24.600 501.900 25.800 ;
        RECT 495.000 23.850 495.900 24.600 ;
        RECT 500.100 24.000 501.900 24.600 ;
        RECT 494.100 22.050 495.900 23.850 ;
        RECT 497.100 22.950 498.900 23.700 ;
        RECT 511.050 22.950 511.950 27.000 ;
        RECT 520.950 25.050 525.450 27.150 ;
        RECT 519.150 23.250 523.050 25.050 ;
        RECT 520.950 22.950 523.050 23.250 ;
        RECT 497.100 21.900 505.050 22.950 ;
        RECT 502.950 20.850 505.050 21.900 ;
        RECT 508.950 20.850 511.950 22.950 ;
        RECT 501.450 17.100 503.250 17.400 ;
        RECT 501.450 16.800 509.850 17.100 ;
        RECT 492.150 16.200 509.850 16.800 ;
        RECT 492.150 15.600 503.250 16.200 ;
        RECT 473.550 3.750 475.350 9.600 ;
        RECT 476.550 3.750 478.350 9.600 ;
        RECT 484.650 3.750 486.450 9.600 ;
        RECT 487.650 3.750 489.450 9.600 ;
        RECT 492.150 3.750 493.950 15.600 ;
        RECT 506.250 14.700 508.050 15.300 ;
        RECT 500.550 13.500 508.050 14.700 ;
        RECT 508.950 14.100 509.850 16.200 ;
        RECT 511.050 16.200 511.950 20.850 ;
        RECT 521.250 17.400 523.050 19.200 ;
        RECT 517.950 16.200 522.150 17.400 ;
        RECT 511.050 15.300 517.050 16.200 ;
        RECT 517.950 15.300 520.050 16.200 ;
        RECT 524.250 15.600 525.450 25.050 ;
        RECT 532.950 25.950 534.000 32.400 ;
        RECT 539.550 29.400 541.350 35.250 ;
        RECT 542.850 32.400 544.650 35.250 ;
        RECT 547.350 32.400 549.150 35.250 ;
        RECT 551.550 32.400 553.350 35.250 ;
        RECT 555.450 32.400 557.250 35.250 ;
        RECT 558.750 32.400 560.550 35.250 ;
        RECT 563.250 33.300 565.050 35.250 ;
        RECT 563.250 32.400 567.000 33.300 ;
        RECT 568.050 32.400 569.850 35.250 ;
        RECT 547.650 31.500 548.700 32.400 ;
        RECT 544.950 30.300 548.700 31.500 ;
        RECT 556.200 30.600 557.250 32.400 ;
        RECT 565.950 31.500 567.000 32.400 ;
        RECT 544.950 29.400 547.050 30.300 ;
        RECT 539.550 27.150 540.750 29.400 ;
        RECT 552.150 28.200 553.950 30.000 ;
        RECT 556.200 29.550 561.150 30.600 ;
        RECT 559.350 28.800 561.150 29.550 ;
        RECT 562.650 28.800 564.450 30.600 ;
        RECT 565.950 29.400 568.050 31.500 ;
        RECT 571.050 29.400 572.850 35.250 ;
        RECT 575.550 32.400 577.350 35.250 ;
        RECT 578.550 32.400 580.350 35.250 ;
        RECT 553.050 27.900 553.950 28.200 ;
        RECT 563.100 27.900 564.150 28.800 ;
        RECT 532.950 23.850 535.050 25.950 ;
        RECT 539.550 25.050 544.050 27.150 ;
        RECT 553.050 27.000 564.150 27.900 ;
        RECT 529.950 20.850 532.050 22.950 ;
        RECT 530.100 19.050 531.900 20.850 ;
        RECT 532.950 16.650 534.000 23.850 ;
        RECT 535.950 20.850 538.050 22.950 ;
        RECT 536.100 19.050 537.900 20.850 ;
        RECT 516.150 14.400 517.050 15.300 ;
        RECT 513.450 14.100 515.250 14.400 ;
        RECT 500.550 12.600 501.750 13.500 ;
        RECT 508.950 13.200 515.250 14.100 ;
        RECT 513.450 12.600 515.250 13.200 ;
        RECT 516.150 12.600 518.850 14.400 ;
        RECT 496.950 10.500 501.750 12.600 ;
        RECT 504.150 10.500 511.050 12.300 ;
        RECT 500.550 9.600 501.750 10.500 ;
        RECT 495.150 3.750 496.950 9.600 ;
        RECT 500.250 3.750 502.050 9.600 ;
        RECT 505.050 3.750 506.850 9.600 ;
        RECT 508.050 3.750 509.850 10.500 ;
        RECT 516.150 9.600 520.050 11.700 ;
        RECT 511.950 3.750 513.750 9.600 ;
        RECT 516.150 3.750 517.950 9.600 ;
        RECT 520.650 3.750 522.450 6.600 ;
        RECT 523.650 3.750 525.450 15.600 ;
        RECT 531.450 15.600 534.000 16.650 ;
        RECT 539.550 15.600 540.750 25.050 ;
        RECT 541.950 23.250 545.850 25.050 ;
        RECT 541.950 22.950 544.050 23.250 ;
        RECT 553.050 22.950 553.950 27.000 ;
        RECT 563.100 25.800 564.150 27.000 ;
        RECT 563.100 24.600 570.000 25.800 ;
        RECT 563.100 24.000 564.900 24.600 ;
        RECT 569.100 23.850 570.000 24.600 ;
        RECT 566.100 22.950 567.900 23.700 ;
        RECT 553.050 20.850 556.050 22.950 ;
        RECT 559.950 21.900 567.900 22.950 ;
        RECT 569.100 22.050 570.900 23.850 ;
        RECT 559.950 20.850 562.050 21.900 ;
        RECT 541.950 17.400 543.750 19.200 ;
        RECT 542.850 16.200 547.050 17.400 ;
        RECT 553.050 16.200 553.950 20.850 ;
        RECT 561.750 17.100 563.550 17.400 ;
        RECT 531.450 3.750 533.250 15.600 ;
        RECT 535.650 3.750 537.450 15.600 ;
        RECT 539.550 3.750 541.350 15.600 ;
        RECT 544.950 15.300 547.050 16.200 ;
        RECT 547.950 15.300 553.950 16.200 ;
        RECT 555.150 16.800 563.550 17.100 ;
        RECT 571.950 16.800 572.850 29.400 ;
        RECT 574.950 23.850 577.050 25.950 ;
        RECT 578.400 24.150 579.600 32.400 ;
        RECT 584.550 30.300 586.350 35.250 ;
        RECT 587.550 31.200 589.350 35.250 ;
        RECT 590.550 30.300 592.350 35.250 ;
        RECT 584.550 28.950 592.350 30.300 ;
        RECT 593.550 29.400 595.350 35.250 ;
        RECT 599.550 32.400 601.350 35.250 ;
        RECT 602.550 32.400 604.350 35.250 ;
        RECT 605.550 32.400 607.350 35.250 ;
        RECT 611.550 32.400 613.350 35.250 ;
        RECT 614.550 32.400 616.350 35.250 ;
        RECT 617.550 32.400 619.350 35.250 ;
        RECT 625.650 32.400 627.450 35.250 ;
        RECT 628.650 32.400 630.450 35.250 ;
        RECT 631.650 32.400 633.450 35.250 ;
        RECT 593.550 27.300 594.750 29.400 ;
        RECT 591.000 26.250 594.750 27.300 ;
        RECT 587.100 24.150 588.900 25.950 ;
        RECT 575.100 22.050 576.900 23.850 ;
        RECT 577.950 22.050 580.050 24.150 ;
        RECT 555.150 16.200 572.850 16.800 ;
        RECT 547.950 14.400 548.850 15.300 ;
        RECT 546.150 12.600 548.850 14.400 ;
        RECT 549.750 14.100 551.550 14.400 ;
        RECT 555.150 14.100 556.050 16.200 ;
        RECT 561.750 15.600 572.850 16.200 ;
        RECT 549.750 13.200 556.050 14.100 ;
        RECT 556.950 14.700 558.750 15.300 ;
        RECT 556.950 13.500 564.450 14.700 ;
        RECT 549.750 12.600 551.550 13.200 ;
        RECT 563.250 12.600 564.450 13.500 ;
        RECT 544.950 9.600 548.850 11.700 ;
        RECT 553.950 10.500 560.850 12.300 ;
        RECT 563.250 10.500 568.050 12.600 ;
        RECT 542.550 3.750 544.350 6.600 ;
        RECT 547.050 3.750 548.850 9.600 ;
        RECT 551.250 3.750 553.050 9.600 ;
        RECT 555.150 3.750 556.950 10.500 ;
        RECT 563.250 9.600 564.450 10.500 ;
        RECT 558.150 3.750 559.950 9.600 ;
        RECT 562.950 3.750 564.750 9.600 ;
        RECT 568.050 3.750 569.850 9.600 ;
        RECT 571.050 3.750 572.850 15.600 ;
        RECT 578.400 9.600 579.600 22.050 ;
        RECT 583.950 20.850 586.050 22.950 ;
        RECT 586.950 22.050 589.050 24.150 ;
        RECT 590.850 22.950 592.050 26.250 ;
        RECT 603.000 25.950 604.050 32.400 ;
        RECT 615.000 25.950 616.050 32.400 ;
        RECT 601.950 23.850 604.050 25.950 ;
        RECT 613.950 23.850 616.050 25.950 ;
        RECT 589.950 20.850 592.050 22.950 ;
        RECT 598.950 20.850 601.050 22.950 ;
        RECT 584.100 19.050 585.900 20.850 ;
        RECT 589.950 15.600 591.150 20.850 ;
        RECT 592.950 17.850 595.050 19.950 ;
        RECT 599.100 19.050 600.900 20.850 ;
        RECT 592.950 16.050 594.750 17.850 ;
        RECT 603.000 16.650 604.050 23.850 ;
        RECT 604.950 20.850 607.050 22.950 ;
        RECT 610.950 20.850 613.050 22.950 ;
        RECT 605.100 19.050 606.900 20.850 ;
        RECT 611.100 19.050 612.900 20.850 ;
        RECT 615.000 16.650 616.050 23.850 ;
        RECT 628.950 25.950 630.000 32.400 ;
        RECT 635.550 30.300 637.350 35.250 ;
        RECT 638.550 31.200 640.350 35.250 ;
        RECT 641.550 30.300 643.350 35.250 ;
        RECT 635.550 28.950 643.350 30.300 ;
        RECT 644.550 29.400 646.350 35.250 ;
        RECT 644.550 27.300 645.750 29.400 ;
        RECT 653.850 28.200 655.650 35.250 ;
        RECT 658.350 29.400 660.150 35.250 ;
        RECT 664.650 32.400 666.450 35.250 ;
        RECT 667.650 32.400 669.450 35.250 ;
        RECT 671.550 32.400 673.350 35.250 ;
        RECT 674.550 32.400 676.350 35.250 ;
        RECT 677.550 32.400 679.350 35.250 ;
        RECT 653.850 27.300 657.450 28.200 ;
        RECT 642.000 26.250 645.750 27.300 ;
        RECT 628.950 23.850 631.050 25.950 ;
        RECT 638.100 24.150 639.900 25.950 ;
        RECT 616.950 20.850 619.050 22.950 ;
        RECT 625.950 20.850 628.050 22.950 ;
        RECT 617.100 19.050 618.900 20.850 ;
        RECT 626.100 19.050 627.900 20.850 ;
        RECT 628.950 16.650 630.000 23.850 ;
        RECT 631.950 20.850 634.050 22.950 ;
        RECT 634.950 20.850 637.050 22.950 ;
        RECT 637.950 22.050 640.050 24.150 ;
        RECT 641.850 22.950 643.050 26.250 ;
        RECT 640.950 20.850 643.050 22.950 ;
        RECT 653.100 21.150 654.900 22.950 ;
        RECT 632.100 19.050 633.900 20.850 ;
        RECT 635.100 19.050 636.900 20.850 ;
        RECT 603.000 15.600 605.550 16.650 ;
        RECT 615.000 15.600 617.550 16.650 ;
        RECT 575.550 3.750 577.350 9.600 ;
        RECT 578.550 3.750 580.350 9.600 ;
        RECT 585.300 3.750 587.100 15.600 ;
        RECT 589.500 3.750 591.300 15.600 ;
        RECT 592.800 3.750 594.600 9.600 ;
        RECT 599.550 3.750 601.350 15.600 ;
        RECT 603.750 3.750 605.550 15.600 ;
        RECT 611.550 3.750 613.350 15.600 ;
        RECT 615.750 3.750 617.550 15.600 ;
        RECT 627.450 15.600 630.000 16.650 ;
        RECT 640.950 15.600 642.150 20.850 ;
        RECT 643.950 17.850 646.050 19.950 ;
        RECT 652.950 19.050 655.050 21.150 ;
        RECT 656.250 19.950 657.450 27.300 ;
        RECT 665.400 24.150 666.600 32.400 ;
        RECT 675.000 25.950 676.050 32.400 ;
        RECT 683.850 29.400 685.650 35.250 ;
        RECT 688.350 28.200 690.150 35.250 ;
        RECT 697.650 32.400 699.450 35.250 ;
        RECT 700.650 32.400 702.450 35.250 ;
        RECT 659.100 21.150 660.900 22.950 ;
        RECT 664.950 22.050 667.050 24.150 ;
        RECT 667.950 23.850 670.050 25.950 ;
        RECT 673.950 23.850 676.050 25.950 ;
        RECT 668.100 22.050 669.900 23.850 ;
        RECT 655.950 17.850 658.050 19.950 ;
        RECT 658.950 19.050 661.050 21.150 ;
        RECT 643.950 16.050 645.750 17.850 ;
        RECT 627.450 3.750 629.250 15.600 ;
        RECT 631.650 3.750 633.450 15.600 ;
        RECT 636.300 3.750 638.100 15.600 ;
        RECT 640.500 3.750 642.300 15.600 ;
        RECT 656.250 9.600 657.450 17.850 ;
        RECT 665.400 9.600 666.600 22.050 ;
        RECT 670.950 20.850 673.050 22.950 ;
        RECT 671.100 19.050 672.900 20.850 ;
        RECT 675.000 16.650 676.050 23.850 ;
        RECT 686.550 27.300 690.150 28.200 ;
        RECT 676.950 20.850 679.050 22.950 ;
        RECT 683.100 21.150 684.900 22.950 ;
        RECT 677.100 19.050 678.900 20.850 ;
        RECT 682.950 19.050 685.050 21.150 ;
        RECT 686.550 19.950 687.750 27.300 ;
        RECT 698.400 24.150 699.600 32.400 ;
        RECT 704.850 29.400 706.650 35.250 ;
        RECT 709.350 28.200 711.150 35.250 ;
        RECT 707.550 27.300 711.150 28.200 ;
        RECT 689.100 21.150 690.900 22.950 ;
        RECT 697.950 22.050 700.050 24.150 ;
        RECT 700.950 23.850 703.050 25.950 ;
        RECT 701.100 22.050 702.900 23.850 ;
        RECT 685.950 17.850 688.050 19.950 ;
        RECT 688.950 19.050 691.050 21.150 ;
        RECT 675.000 15.600 677.550 16.650 ;
        RECT 643.800 3.750 645.600 9.600 ;
        RECT 652.650 3.750 654.450 9.600 ;
        RECT 655.650 3.750 657.450 9.600 ;
        RECT 658.650 3.750 660.450 9.600 ;
        RECT 664.650 3.750 666.450 9.600 ;
        RECT 667.650 3.750 669.450 9.600 ;
        RECT 671.550 3.750 673.350 15.600 ;
        RECT 675.750 3.750 677.550 15.600 ;
        RECT 686.550 9.600 687.750 17.850 ;
        RECT 698.400 9.600 699.600 22.050 ;
        RECT 704.100 21.150 705.900 22.950 ;
        RECT 703.950 19.050 706.050 21.150 ;
        RECT 707.550 19.950 708.750 27.300 ;
        RECT 710.100 21.150 711.900 22.950 ;
        RECT 706.950 17.850 709.050 19.950 ;
        RECT 709.950 19.050 712.050 21.150 ;
        RECT 707.550 9.600 708.750 17.850 ;
        RECT 683.550 3.750 685.350 9.600 ;
        RECT 686.550 3.750 688.350 9.600 ;
        RECT 689.550 3.750 691.350 9.600 ;
        RECT 697.650 3.750 699.450 9.600 ;
        RECT 700.650 3.750 702.450 9.600 ;
        RECT 704.550 3.750 706.350 9.600 ;
        RECT 707.550 3.750 709.350 9.600 ;
        RECT 710.550 3.750 712.350 9.600 ;
      LAYER metal2 ;
        RECT 184.950 682.950 187.050 685.050 ;
        RECT 229.950 682.950 232.050 685.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 28.950 679.950 31.050 682.050 ;
        RECT 133.950 679.950 136.050 682.050 ;
        RECT 4.950 676.950 7.050 679.050 ;
        RECT 5.400 673.050 6.450 676.950 ;
        RECT 10.950 673.950 13.050 676.050 ;
        RECT 4.950 670.950 7.050 673.050 ;
        RECT 8.250 671.250 10.050 672.150 ;
        RECT 10.950 671.850 13.050 672.750 ;
        RECT 13.950 671.250 16.050 672.150 ;
        RECT 4.950 668.850 6.750 669.750 ;
        RECT 7.950 667.950 10.050 670.050 ;
        RECT 13.950 667.950 16.050 670.050 ;
        RECT 8.400 661.050 9.450 667.950 ;
        RECT 14.400 664.050 15.450 667.950 ;
        RECT 13.950 661.950 16.050 664.050 ;
        RECT 17.400 661.050 18.450 679.950 ;
        RECT 25.950 673.950 28.050 676.050 ;
        RECT 26.400 673.050 27.450 673.950 ;
        RECT 25.950 670.950 28.050 673.050 ;
        RECT 19.950 668.250 21.750 669.150 ;
        RECT 22.950 667.950 25.050 670.050 ;
        RECT 26.400 667.050 27.450 670.950 ;
        RECT 29.400 670.050 30.450 679.950 ;
        RECT 73.950 676.950 76.050 679.050 ;
        RECT 106.950 676.950 109.050 679.050 ;
        RECT 74.400 676.050 75.450 676.950 ;
        RECT 55.950 673.950 58.050 676.050 ;
        RECT 64.950 673.950 67.050 676.050 ;
        RECT 73.950 673.950 76.050 676.050 ;
        RECT 82.950 673.950 85.050 676.050 ;
        RECT 97.950 673.950 100.050 676.050 ;
        RECT 31.950 670.950 34.050 673.050 ;
        RECT 32.400 670.050 33.450 670.950 ;
        RECT 28.950 667.950 31.050 670.050 ;
        RECT 31.950 667.950 34.050 670.050 ;
        RECT 34.950 667.950 37.050 670.050 ;
        RECT 37.950 667.950 40.050 670.050 ;
        RECT 41.250 668.250 43.050 669.150 ;
        RECT 46.950 667.950 49.050 670.050 ;
        RECT 49.950 668.250 51.750 669.150 ;
        RECT 52.950 667.950 55.050 670.050 ;
        RECT 35.400 667.050 36.450 667.950 ;
        RECT 19.950 664.950 22.050 667.050 ;
        RECT 23.250 665.850 24.750 666.750 ;
        RECT 25.950 664.950 28.050 667.050 ;
        RECT 29.250 665.850 31.050 666.750 ;
        RECT 31.950 665.850 33.750 666.750 ;
        RECT 34.950 664.950 37.050 667.050 ;
        RECT 38.250 665.850 39.750 666.750 ;
        RECT 40.950 664.950 43.050 667.050 ;
        RECT 7.950 658.950 10.050 661.050 ;
        RECT 16.950 658.950 19.050 661.050 ;
        RECT 20.400 655.050 21.450 664.950 ;
        RECT 22.950 661.950 25.050 664.050 ;
        RECT 25.950 662.850 28.050 663.750 ;
        RECT 28.950 661.950 31.050 664.050 ;
        RECT 34.950 662.850 37.050 663.750 ;
        RECT 19.950 652.950 22.050 655.050 ;
        RECT 4.950 634.950 7.050 637.050 ;
        RECT 13.950 634.950 16.050 637.050 ;
        RECT 5.400 634.050 6.450 634.950 ;
        RECT 4.950 631.950 7.050 634.050 ;
        RECT 8.250 632.250 9.750 633.150 ;
        RECT 10.950 631.950 13.050 634.050 ;
        RECT 14.400 631.050 15.450 634.950 ;
        RECT 23.400 634.050 24.450 661.950 ;
        RECT 25.950 658.950 28.050 661.050 ;
        RECT 22.950 631.950 25.050 634.050 ;
        RECT 4.950 629.850 6.750 630.750 ;
        RECT 7.950 628.950 10.050 631.050 ;
        RECT 11.250 629.850 13.050 630.750 ;
        RECT 13.950 628.950 16.050 631.050 ;
        RECT 19.950 628.950 22.050 631.050 ;
        RECT 23.250 629.250 25.050 630.150 ;
        RECT 8.400 622.050 9.450 628.950 ;
        RECT 10.950 625.950 13.050 628.050 ;
        RECT 13.950 626.850 16.050 627.750 ;
        RECT 16.950 626.250 19.050 627.150 ;
        RECT 19.950 626.850 21.750 627.750 ;
        RECT 22.950 625.950 25.050 628.050 ;
        RECT 7.950 619.950 10.050 622.050 ;
        RECT 7.950 604.950 10.050 607.050 ;
        RECT 8.400 598.050 9.450 604.950 ;
        RECT 11.400 604.050 12.450 625.950 ;
        RECT 16.950 622.950 19.050 625.050 ;
        RECT 10.950 601.950 13.050 604.050 ;
        RECT 17.400 598.050 18.450 622.950 ;
        RECT 23.400 616.050 24.450 625.950 ;
        RECT 26.400 619.050 27.450 658.950 ;
        RECT 25.950 616.950 28.050 619.050 ;
        RECT 22.950 613.950 25.050 616.050 ;
        RECT 22.950 610.950 25.050 613.050 ;
        RECT 4.950 596.250 6.750 597.150 ;
        RECT 7.950 595.950 10.050 598.050 ;
        RECT 11.250 596.250 13.050 597.150 ;
        RECT 13.950 596.250 15.750 597.150 ;
        RECT 16.950 595.950 19.050 598.050 ;
        RECT 20.250 596.250 22.050 597.150 ;
        RECT 4.950 594.450 7.050 595.050 ;
        RECT 2.400 593.400 7.050 594.450 ;
        RECT 8.250 593.850 9.750 594.750 ;
        RECT 10.950 594.450 13.050 595.050 ;
        RECT 13.950 594.450 16.050 595.050 ;
        RECT 2.400 555.450 3.450 593.400 ;
        RECT 4.950 592.950 7.050 593.400 ;
        RECT 10.950 593.400 16.050 594.450 ;
        RECT 17.250 593.850 18.750 594.750 ;
        RECT 10.950 592.950 13.050 593.400 ;
        RECT 13.950 592.950 16.050 593.400 ;
        RECT 19.950 592.950 22.050 595.050 ;
        RECT 7.950 583.950 10.050 586.050 ;
        RECT 8.400 559.050 9.450 583.950 ;
        RECT 11.400 562.050 12.450 592.950 ;
        RECT 20.400 592.050 21.450 592.950 ;
        RECT 19.950 589.950 22.050 592.050 ;
        RECT 20.400 562.050 21.450 589.950 ;
        RECT 23.400 583.050 24.450 610.950 ;
        RECT 26.400 591.450 27.450 616.950 ;
        RECT 29.400 610.050 30.450 661.950 ;
        RECT 47.400 634.050 48.450 667.950 ;
        RECT 56.400 667.050 57.450 673.950 ;
        RECT 83.400 673.050 84.450 673.950 ;
        RECT 98.400 673.050 99.450 673.950 ;
        RECT 58.950 670.950 61.050 673.050 ;
        RECT 61.950 671.250 64.050 672.150 ;
        RECT 64.950 671.850 67.050 672.750 ;
        RECT 67.950 671.250 69.750 672.150 ;
        RECT 70.950 670.950 73.050 673.050 ;
        RECT 76.950 672.450 79.050 673.050 ;
        RECT 74.400 671.400 79.050 672.450 ;
        RECT 59.400 670.050 60.450 670.950 ;
        RECT 74.400 670.050 75.450 671.400 ;
        RECT 76.950 670.950 79.050 671.400 ;
        RECT 80.250 671.250 81.750 672.150 ;
        RECT 82.950 670.950 85.050 673.050 ;
        RECT 91.950 670.950 94.050 673.050 ;
        RECT 95.250 671.250 96.750 672.150 ;
        RECT 97.950 670.950 100.050 673.050 ;
        RECT 58.950 667.950 61.050 670.050 ;
        RECT 61.950 667.950 64.050 670.050 ;
        RECT 67.950 667.950 70.050 670.050 ;
        RECT 71.250 668.850 73.050 669.750 ;
        RECT 73.950 667.950 76.050 670.050 ;
        RECT 76.950 668.850 78.750 669.750 ;
        RECT 79.950 667.950 82.050 670.050 ;
        RECT 83.250 668.850 84.750 669.750 ;
        RECT 85.950 669.450 88.050 670.050 ;
        RECT 85.950 668.400 90.450 669.450 ;
        RECT 91.950 668.850 93.750 669.750 ;
        RECT 85.950 667.950 88.050 668.400 ;
        RECT 49.950 664.950 52.050 667.050 ;
        RECT 53.250 665.850 54.750 666.750 ;
        RECT 55.950 664.950 58.050 667.050 ;
        RECT 59.250 665.850 61.050 666.750 ;
        RECT 50.400 661.050 51.450 664.950 ;
        RECT 55.950 662.850 58.050 663.750 ;
        RECT 49.950 658.950 52.050 661.050 ;
        RECT 62.400 643.050 63.450 667.950 ;
        RECT 68.400 649.050 69.450 667.950 ;
        RECT 80.400 667.050 81.450 667.950 ;
        RECT 73.950 666.450 76.050 667.050 ;
        RECT 76.950 666.450 79.050 667.050 ;
        RECT 73.950 665.400 79.050 666.450 ;
        RECT 73.950 664.950 76.050 665.400 ;
        RECT 76.950 664.950 79.050 665.400 ;
        RECT 79.950 664.950 82.050 667.050 ;
        RECT 85.950 665.850 88.050 666.750 ;
        RECT 89.400 655.050 90.450 668.400 ;
        RECT 94.950 667.950 97.050 670.050 ;
        RECT 98.250 668.850 99.750 669.750 ;
        RECT 100.950 667.950 103.050 670.050 ;
        RECT 103.950 667.950 106.050 670.050 ;
        RECT 91.950 664.950 94.050 667.050 ;
        RECT 82.950 652.950 85.050 655.050 ;
        RECT 88.950 652.950 91.050 655.050 ;
        RECT 67.950 646.950 70.050 649.050 ;
        RECT 52.950 640.950 55.050 643.050 ;
        RECT 61.950 640.950 64.050 643.050 ;
        RECT 31.950 631.950 34.050 634.050 ;
        RECT 37.950 633.450 40.050 634.050 ;
        RECT 35.250 632.250 36.750 633.150 ;
        RECT 37.950 632.400 42.450 633.450 ;
        RECT 37.950 631.950 40.050 632.400 ;
        RECT 31.950 629.850 33.750 630.750 ;
        RECT 34.950 628.950 37.050 631.050 ;
        RECT 38.250 629.850 40.050 630.750 ;
        RECT 37.950 625.950 40.050 628.050 ;
        RECT 28.950 607.950 31.050 610.050 ;
        RECT 31.950 601.950 34.050 604.050 ;
        RECT 32.400 598.050 33.450 601.950 ;
        RECT 38.400 598.050 39.450 625.950 ;
        RECT 41.400 613.050 42.450 632.400 ;
        RECT 46.950 631.950 49.050 634.050 ;
        RECT 43.950 629.250 46.050 630.150 ;
        RECT 49.950 629.250 52.050 630.150 ;
        RECT 53.400 628.050 54.450 640.950 ;
        RECT 55.950 632.250 58.050 633.150 ;
        RECT 76.950 632.250 79.050 633.150 ;
        RECT 55.950 628.950 58.050 631.050 ;
        RECT 59.250 629.250 60.750 630.150 ;
        RECT 61.950 628.950 64.050 631.050 ;
        RECT 65.250 629.250 67.050 630.150 ;
        RECT 67.950 629.250 69.750 630.150 ;
        RECT 70.950 628.950 73.050 631.050 ;
        RECT 74.250 629.250 75.750 630.150 ;
        RECT 76.950 628.950 79.050 631.050 ;
        RECT 43.950 625.950 46.050 628.050 ;
        RECT 47.250 626.250 48.750 627.150 ;
        RECT 49.950 625.950 52.050 628.050 ;
        RECT 52.950 625.950 55.050 628.050 ;
        RECT 44.400 622.050 45.450 625.950 ;
        RECT 46.950 622.950 49.050 625.050 ;
        RECT 43.950 619.950 46.050 622.050 ;
        RECT 50.400 613.050 51.450 625.950 ;
        RECT 56.400 619.050 57.450 628.950 ;
        RECT 58.950 625.950 61.050 628.050 ;
        RECT 62.250 626.850 63.750 627.750 ;
        RECT 64.950 627.450 67.050 628.050 ;
        RECT 67.950 627.450 70.050 628.050 ;
        RECT 64.950 626.400 70.050 627.450 ;
        RECT 71.250 626.850 72.750 627.750 ;
        RECT 64.950 625.950 67.050 626.400 ;
        RECT 67.950 625.950 70.050 626.400 ;
        RECT 73.950 625.950 76.050 628.050 ;
        RECT 55.950 616.950 58.050 619.050 ;
        RECT 65.400 616.050 66.450 625.950 ;
        RECT 77.400 619.050 78.450 628.950 ;
        RECT 83.400 625.050 84.450 652.950 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 86.400 631.050 87.450 646.950 ;
        RECT 85.950 628.950 88.050 631.050 ;
        RECT 85.950 626.850 88.050 627.750 ;
        RECT 92.400 627.450 93.450 664.950 ;
        RECT 95.400 664.050 96.450 667.950 ;
        RECT 97.950 664.950 100.050 667.050 ;
        RECT 100.950 665.850 103.050 666.750 ;
        RECT 94.950 661.950 97.050 664.050 ;
        RECT 98.400 658.050 99.450 664.950 ;
        RECT 104.400 661.050 105.450 667.950 ;
        RECT 107.400 666.450 108.450 676.950 ;
        RECT 113.400 674.400 129.450 675.450 ;
        RECT 113.400 673.050 114.450 674.400 ;
        RECT 128.400 673.050 129.450 674.400 ;
        RECT 112.950 670.950 115.050 673.050 ;
        RECT 115.950 670.950 118.050 673.050 ;
        RECT 124.950 670.950 127.050 673.050 ;
        RECT 127.950 670.950 130.050 673.050 ;
        RECT 109.950 668.250 111.750 669.150 ;
        RECT 112.950 667.950 115.050 670.050 ;
        RECT 116.400 667.050 117.450 670.950 ;
        RECT 118.950 667.950 121.050 670.050 ;
        RECT 121.950 667.950 124.050 670.050 ;
        RECT 125.400 667.050 126.450 670.950 ;
        RECT 127.950 667.950 130.050 670.050 ;
        RECT 131.250 668.250 133.050 669.150 ;
        RECT 109.950 666.450 112.050 667.050 ;
        RECT 107.400 665.400 112.050 666.450 ;
        RECT 113.250 665.850 114.750 666.750 ;
        RECT 109.950 664.950 112.050 665.400 ;
        RECT 115.950 664.950 118.050 667.050 ;
        RECT 119.250 665.850 121.050 666.750 ;
        RECT 121.950 665.850 123.750 666.750 ;
        RECT 124.950 664.950 127.050 667.050 ;
        RECT 128.250 665.850 129.750 666.750 ;
        RECT 130.950 664.950 133.050 667.050 ;
        RECT 106.950 661.950 109.050 664.050 ;
        RECT 115.950 662.850 118.050 663.750 ;
        RECT 121.950 661.950 124.050 664.050 ;
        RECT 124.950 662.850 127.050 663.750 ;
        RECT 127.950 661.950 130.050 664.050 ;
        RECT 134.400 663.450 135.450 679.950 ;
        RECT 158.400 677.400 171.450 678.450 ;
        RECT 158.400 676.050 159.450 677.400 ;
        RECT 170.400 676.050 171.450 677.400 ;
        RECT 157.950 673.950 160.050 676.050 ;
        RECT 160.950 673.950 163.050 676.050 ;
        RECT 166.950 673.950 169.050 676.050 ;
        RECT 169.950 673.950 172.050 676.050 ;
        RECT 148.950 670.950 151.050 673.050 ;
        RECT 149.400 670.050 150.450 670.950 ;
        RECT 136.950 668.250 138.750 669.150 ;
        RECT 139.950 667.950 142.050 670.050 ;
        RECT 143.250 668.250 145.050 669.150 ;
        RECT 148.950 667.950 151.050 670.050 ;
        RECT 154.950 667.950 157.050 670.050 ;
        RECT 158.250 668.250 160.050 669.150 ;
        RECT 136.950 664.950 139.050 667.050 ;
        RECT 140.250 665.850 141.750 666.750 ;
        RECT 142.950 664.950 145.050 667.050 ;
        RECT 148.950 665.850 150.750 666.750 ;
        RECT 151.950 664.950 154.050 667.050 ;
        RECT 155.250 665.850 156.750 666.750 ;
        RECT 157.950 664.950 160.050 667.050 ;
        RECT 137.400 664.050 138.450 664.950 ;
        RECT 131.400 662.400 135.450 663.450 ;
        RECT 103.950 658.950 106.050 661.050 ;
        RECT 97.950 655.950 100.050 658.050 ;
        RECT 97.950 631.950 100.050 634.050 ;
        RECT 98.400 631.050 99.450 631.950 ;
        RECT 94.950 629.250 96.750 630.150 ;
        RECT 97.950 628.950 100.050 631.050 ;
        RECT 103.950 628.950 106.050 631.050 ;
        RECT 94.950 627.450 97.050 628.050 ;
        RECT 88.950 626.250 91.050 627.150 ;
        RECT 92.400 626.400 97.050 627.450 ;
        RECT 98.250 626.850 100.050 627.750 ;
        RECT 94.950 625.950 97.050 626.400 ;
        RECT 100.950 626.250 103.050 627.150 ;
        RECT 103.950 626.850 106.050 627.750 ;
        RECT 107.400 625.050 108.450 661.950 ;
        RECT 109.950 655.950 112.050 658.050 ;
        RECT 110.400 631.050 111.450 655.950 ;
        RECT 122.400 655.050 123.450 661.950 ;
        RECT 121.950 652.950 124.050 655.050 ;
        RECT 118.950 635.250 121.050 636.150 ;
        RECT 115.950 632.250 117.750 633.150 ;
        RECT 118.950 631.950 121.050 634.050 ;
        RECT 124.950 633.450 127.050 634.050 ;
        RECT 128.400 633.450 129.450 661.950 ;
        RECT 122.250 632.250 123.750 633.150 ;
        RECT 124.950 632.400 129.450 633.450 ;
        RECT 124.950 631.950 127.050 632.400 ;
        RECT 109.950 628.950 112.050 631.050 ;
        RECT 115.950 628.950 118.050 631.050 ;
        RECT 121.950 628.950 124.050 631.050 ;
        RECT 125.250 629.850 127.050 630.750 ;
        RECT 109.950 626.850 112.050 627.750 ;
        RECT 112.950 626.250 115.050 627.150 ;
        RECT 82.950 622.950 85.050 625.050 ;
        RECT 88.950 622.950 91.050 625.050 ;
        RECT 100.950 622.950 103.050 625.050 ;
        RECT 103.950 622.950 106.050 625.050 ;
        RECT 106.950 622.950 109.050 625.050 ;
        RECT 112.950 622.950 115.050 625.050 ;
        RECT 89.400 622.050 90.450 622.950 ;
        RECT 88.950 619.950 91.050 622.050 ;
        RECT 76.950 616.950 79.050 619.050 ;
        RECT 88.950 616.950 91.050 619.050 ;
        RECT 64.950 613.950 67.050 616.050 ;
        RECT 40.950 610.950 43.050 613.050 ;
        RECT 49.950 610.950 52.050 613.050 ;
        RECT 43.950 607.950 46.050 610.050 ;
        RECT 44.400 601.050 45.450 607.950 ;
        RECT 55.950 604.950 58.050 607.050 ;
        RECT 61.950 604.950 64.050 607.050 ;
        RECT 56.400 604.050 57.450 604.950 ;
        RECT 49.950 601.950 52.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 50.400 601.050 51.450 601.950 ;
        RECT 62.400 601.050 63.450 604.950 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 43.950 598.950 46.050 601.050 ;
        RECT 47.250 599.250 48.750 600.150 ;
        RECT 49.950 598.950 52.050 601.050 ;
        RECT 52.950 599.250 55.050 600.150 ;
        RECT 55.950 599.850 58.050 600.750 ;
        RECT 58.950 599.250 60.750 600.150 ;
        RECT 61.950 598.950 64.050 601.050 ;
        RECT 64.950 598.950 67.050 601.050 ;
        RECT 70.950 600.450 73.050 601.050 ;
        RECT 68.400 599.400 73.050 600.450 ;
        RECT 74.250 599.850 75.750 600.750 ;
        RECT 28.950 596.250 30.750 597.150 ;
        RECT 31.950 595.950 34.050 598.050 ;
        RECT 35.250 596.250 37.050 597.150 ;
        RECT 37.950 595.950 40.050 598.050 ;
        RECT 40.950 595.950 43.050 598.050 ;
        RECT 44.250 596.850 45.750 597.750 ;
        RECT 46.950 595.950 49.050 598.050 ;
        RECT 50.250 596.850 52.050 597.750 ;
        RECT 52.950 597.450 55.050 598.050 ;
        RECT 52.950 596.400 57.450 597.450 ;
        RECT 52.950 595.950 55.050 596.400 ;
        RECT 28.950 592.950 31.050 595.050 ;
        RECT 32.250 593.850 33.750 594.750 ;
        RECT 34.950 592.950 37.050 595.050 ;
        RECT 40.950 593.850 43.050 594.750 ;
        RECT 26.400 590.400 30.450 591.450 ;
        RECT 22.950 580.950 25.050 583.050 ;
        RECT 25.950 580.950 28.050 583.050 ;
        RECT 10.950 559.950 13.050 562.050 ;
        RECT 19.950 559.950 22.050 562.050 ;
        RECT 22.950 560.250 25.050 561.150 ;
        RECT 4.950 557.250 7.050 558.150 ;
        RECT 7.950 556.950 10.050 559.050 ;
        RECT 10.950 557.250 13.050 558.150 ;
        RECT 13.950 557.250 15.750 558.150 ;
        RECT 16.950 556.950 19.050 559.050 ;
        RECT 20.250 557.250 21.750 558.150 ;
        RECT 22.950 556.950 25.050 559.050 ;
        RECT 4.950 555.450 7.050 556.050 ;
        RECT 2.400 554.400 7.050 555.450 ;
        RECT 4.950 553.950 7.050 554.400 ;
        RECT 8.250 554.250 9.750 555.150 ;
        RECT 10.950 553.950 13.050 556.050 ;
        RECT 13.950 553.950 16.050 556.050 ;
        RECT 17.250 554.850 18.750 555.750 ;
        RECT 19.950 553.950 22.050 556.050 ;
        RECT 22.950 553.950 25.050 556.050 ;
        RECT 5.400 544.050 6.450 553.950 ;
        RECT 7.950 550.950 10.050 553.050 ;
        RECT 11.400 550.050 12.450 553.950 ;
        RECT 10.950 547.950 13.050 550.050 ;
        RECT 14.400 547.050 15.450 553.950 ;
        RECT 16.950 550.950 19.050 553.050 ;
        RECT 7.950 544.950 10.050 547.050 ;
        RECT 13.950 544.950 16.050 547.050 ;
        RECT 4.950 541.950 7.050 544.050 ;
        RECT 8.400 526.050 9.450 544.950 ;
        RECT 17.400 544.050 18.450 550.950 ;
        RECT 20.400 550.050 21.450 553.950 ;
        RECT 19.950 547.950 22.050 550.050 ;
        RECT 13.950 541.950 16.050 544.050 ;
        RECT 16.950 541.950 19.050 544.050 ;
        RECT 4.950 524.250 6.750 525.150 ;
        RECT 7.950 523.950 10.050 526.050 ;
        RECT 11.250 524.250 13.050 525.150 ;
        RECT 4.950 520.950 7.050 523.050 ;
        RECT 8.250 521.850 9.750 522.750 ;
        RECT 10.950 520.950 13.050 523.050 ;
        RECT 1.950 508.950 4.050 511.050 ;
        RECT 2.400 481.050 3.450 508.950 ;
        RECT 5.400 493.050 6.450 520.950 ;
        RECT 14.400 519.450 15.450 541.950 ;
        RECT 16.950 538.950 19.050 541.050 ;
        RECT 17.400 523.050 18.450 538.950 ;
        RECT 19.950 533.400 22.050 535.500 ;
        RECT 16.950 520.950 19.050 523.050 ;
        RECT 11.400 518.400 15.450 519.450 ;
        RECT 7.950 494.400 10.050 496.500 ;
        RECT 4.950 490.950 7.050 493.050 ;
        RECT 1.950 478.950 4.050 481.050 ;
        RECT 5.400 477.450 6.450 490.950 ;
        RECT 8.400 477.600 9.600 494.400 ;
        RECT 2.400 476.400 6.450 477.450 ;
        RECT 2.400 442.050 3.450 476.400 ;
        RECT 7.950 475.500 10.050 477.600 ;
        RECT 11.400 457.050 12.450 518.400 ;
        RECT 17.400 490.050 18.450 520.950 ;
        RECT 20.400 516.600 21.600 533.400 ;
        RECT 19.950 514.500 22.050 516.600 ;
        RECT 16.950 487.950 19.050 490.050 ;
        RECT 13.950 485.250 16.050 486.150 ;
        RECT 13.950 478.950 16.050 481.050 ;
        RECT 14.400 475.050 15.450 478.950 ;
        RECT 13.950 472.950 16.050 475.050 ;
        RECT 17.400 468.450 18.450 487.950 ;
        RECT 19.950 485.250 22.050 486.150 ;
        RECT 19.950 481.950 22.050 484.050 ;
        RECT 20.400 481.050 21.450 481.950 ;
        RECT 19.950 478.950 22.050 481.050 ;
        RECT 23.400 478.050 24.450 553.950 ;
        RECT 26.400 550.050 27.450 580.950 ;
        RECT 25.950 547.950 28.050 550.050 ;
        RECT 25.950 529.950 28.050 532.050 ;
        RECT 26.400 529.050 27.450 529.950 ;
        RECT 25.950 526.950 28.050 529.050 ;
        RECT 25.950 524.850 28.050 525.750 ;
        RECT 29.400 522.450 30.450 590.400 ;
        RECT 35.400 585.450 36.450 592.950 ;
        RECT 37.950 586.950 40.050 589.050 ;
        RECT 38.400 585.450 39.450 586.950 ;
        RECT 47.400 586.050 48.450 595.950 ;
        RECT 52.950 592.950 55.050 595.050 ;
        RECT 35.400 584.400 39.450 585.450 ;
        RECT 31.950 556.950 34.050 559.050 ;
        RECT 31.950 554.850 34.050 555.750 ;
        RECT 38.400 555.450 39.450 584.400 ;
        RECT 46.950 583.950 49.050 586.050 ;
        RECT 53.400 559.050 54.450 592.950 ;
        RECT 56.400 583.050 57.450 596.400 ;
        RECT 58.950 595.950 61.050 598.050 ;
        RECT 62.250 596.850 64.050 597.750 ;
        RECT 59.400 586.050 60.450 595.950 ;
        RECT 65.400 589.050 66.450 598.950 ;
        RECT 68.400 592.050 69.450 599.400 ;
        RECT 70.950 598.950 73.050 599.400 ;
        RECT 76.950 598.950 79.050 601.050 ;
        RECT 70.950 596.850 73.050 597.750 ;
        RECT 76.950 596.850 79.050 597.750 ;
        RECT 79.950 596.250 81.750 597.150 ;
        RECT 82.950 595.950 85.050 598.050 ;
        RECT 86.250 596.250 88.050 597.150 ;
        RECT 79.950 592.950 82.050 595.050 ;
        RECT 83.250 593.850 84.750 594.750 ;
        RECT 85.950 592.950 88.050 595.050 ;
        RECT 67.950 589.950 70.050 592.050 ;
        RECT 80.400 589.050 81.450 592.950 ;
        RECT 86.400 592.050 87.450 592.950 ;
        RECT 85.950 589.950 88.050 592.050 ;
        RECT 64.950 586.950 67.050 589.050 ;
        RECT 79.950 586.950 82.050 589.050 ;
        RECT 89.400 586.050 90.450 616.950 ;
        RECT 97.950 607.950 100.050 610.050 ;
        RECT 98.400 601.050 99.450 607.950 ;
        RECT 91.950 598.950 94.050 601.050 ;
        RECT 95.250 599.250 96.750 600.150 ;
        RECT 97.950 598.950 100.050 601.050 ;
        RECT 91.950 596.850 93.750 597.750 ;
        RECT 94.950 595.950 97.050 598.050 ;
        RECT 98.250 596.850 99.750 597.750 ;
        RECT 100.950 595.950 103.050 598.050 ;
        RECT 100.950 593.850 103.050 594.750 ;
        RECT 97.950 589.950 100.050 592.050 ;
        RECT 58.950 583.950 61.050 586.050 ;
        RECT 79.950 583.950 82.050 586.050 ;
        RECT 88.950 583.950 91.050 586.050 ;
        RECT 55.950 580.950 58.050 583.050 ;
        RECT 61.950 562.950 64.050 565.050 ;
        RECT 58.950 559.950 61.050 562.050 ;
        RECT 40.950 557.250 42.750 558.150 ;
        RECT 43.950 556.950 46.050 559.050 ;
        RECT 49.950 556.950 52.050 559.050 ;
        RECT 52.950 556.950 55.050 559.050 ;
        RECT 55.950 557.250 58.050 558.150 ;
        RECT 58.950 557.850 61.050 558.750 ;
        RECT 40.950 555.450 43.050 556.050 ;
        RECT 34.950 554.250 37.050 555.150 ;
        RECT 38.400 554.400 43.050 555.450 ;
        RECT 44.250 554.850 46.050 555.750 ;
        RECT 40.950 553.950 43.050 554.400 ;
        RECT 46.950 554.250 49.050 555.150 ;
        RECT 49.950 554.850 52.050 555.750 ;
        RECT 52.950 553.950 55.050 556.050 ;
        RECT 55.950 553.950 58.050 556.050 ;
        RECT 34.950 550.950 37.050 553.050 ;
        RECT 37.950 550.950 40.050 553.050 ;
        RECT 46.950 550.950 49.050 553.050 ;
        RECT 35.400 547.050 36.450 550.950 ;
        RECT 34.950 544.950 37.050 547.050 ;
        RECT 31.950 528.450 34.050 529.050 ;
        RECT 31.950 527.400 36.450 528.450 ;
        RECT 31.950 526.950 34.050 527.400 ;
        RECT 31.950 524.850 34.050 525.750 ;
        RECT 26.400 521.400 30.450 522.450 ;
        RECT 26.400 487.050 27.450 521.400 ;
        RECT 28.950 495.300 31.050 497.400 ;
        RECT 29.250 491.700 30.450 495.300 ;
        RECT 28.950 489.600 31.050 491.700 ;
        RECT 25.950 484.950 28.050 487.050 ;
        RECT 25.950 481.950 28.050 484.050 ;
        RECT 19.950 475.950 22.050 478.050 ;
        RECT 22.950 475.950 25.050 478.050 ;
        RECT 20.400 472.050 21.450 475.950 ;
        RECT 19.950 469.950 22.050 472.050 ;
        RECT 26.400 471.450 27.450 481.950 ;
        RECT 29.250 477.600 30.450 489.600 ;
        RECT 31.950 481.950 34.050 484.050 ;
        RECT 35.400 481.050 36.450 527.400 ;
        RECT 38.400 505.050 39.450 550.950 ;
        RECT 46.950 544.950 49.050 547.050 ;
        RECT 40.950 533.400 43.050 535.500 ;
        RECT 41.250 521.400 42.450 533.400 ;
        RECT 43.950 530.250 46.050 531.150 ;
        RECT 43.950 526.950 46.050 529.050 ;
        RECT 40.950 519.300 43.050 521.400 ;
        RECT 41.250 515.700 42.450 519.300 ;
        RECT 44.400 517.050 45.450 526.950 ;
        RECT 40.950 513.600 43.050 515.700 ;
        RECT 43.950 514.950 46.050 517.050 ;
        RECT 44.400 511.050 45.450 514.950 ;
        RECT 43.950 508.950 46.050 511.050 ;
        RECT 37.950 502.950 40.050 505.050 ;
        RECT 37.950 499.950 40.050 502.050 ;
        RECT 31.950 479.850 34.050 480.750 ;
        RECT 34.950 478.950 37.050 481.050 ;
        RECT 28.950 475.500 31.050 477.600 ;
        RECT 26.400 470.400 30.450 471.450 ;
        RECT 17.400 467.400 21.450 468.450 ;
        RECT 4.950 454.950 7.050 457.050 ;
        RECT 8.250 455.250 9.750 456.150 ;
        RECT 10.950 454.950 13.050 457.050 ;
        RECT 14.250 455.250 15.750 456.150 ;
        RECT 16.950 454.950 19.050 457.050 ;
        RECT 4.950 452.850 6.750 453.750 ;
        RECT 7.950 451.950 10.050 454.050 ;
        RECT 11.250 452.850 12.750 453.750 ;
        RECT 13.950 451.950 16.050 454.050 ;
        RECT 17.250 452.850 19.050 453.750 ;
        RECT 4.950 448.950 7.050 451.050 ;
        RECT 1.950 439.950 4.050 442.050 ;
        RECT 1.950 415.950 4.050 418.050 ;
        RECT 2.400 406.050 3.450 415.950 ;
        RECT 5.400 415.050 6.450 448.950 ;
        RECT 8.400 448.050 9.450 451.950 ;
        RECT 10.950 448.950 13.050 451.050 ;
        RECT 20.400 450.450 21.450 467.400 ;
        RECT 22.950 457.950 25.050 460.050 ;
        RECT 23.400 457.050 24.450 457.950 ;
        RECT 22.950 454.950 25.050 457.050 ;
        RECT 22.950 452.850 25.050 453.750 ;
        RECT 25.950 452.250 28.050 453.150 ;
        RECT 20.400 449.400 24.450 450.450 ;
        RECT 7.950 445.950 10.050 448.050 ;
        RECT 7.950 436.950 10.050 439.050 ;
        RECT 8.400 415.050 9.450 436.950 ;
        RECT 11.400 427.050 12.450 448.950 ;
        RECT 13.950 445.950 16.050 448.050 ;
        RECT 10.950 424.950 13.050 427.050 ;
        RECT 14.400 423.450 15.450 445.950 ;
        RECT 11.400 422.400 15.450 423.450 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 7.950 412.950 10.050 415.050 ;
        RECT 4.950 410.850 7.050 411.750 ;
        RECT 7.950 410.250 10.050 411.150 ;
        RECT 4.950 406.950 7.050 409.050 ;
        RECT 7.950 406.950 10.050 409.050 ;
        RECT 1.950 403.950 4.050 406.050 ;
        RECT 5.400 388.050 6.450 406.950 ;
        RECT 8.400 406.050 9.450 406.950 ;
        RECT 7.950 403.950 10.050 406.050 ;
        RECT 7.950 397.950 10.050 400.050 ;
        RECT 4.950 385.950 7.050 388.050 ;
        RECT 1.950 382.950 4.050 385.050 ;
        RECT 2.400 382.050 3.450 382.950 ;
        RECT 1.950 379.950 4.050 382.050 ;
        RECT 5.400 379.050 6.450 385.950 ;
        RECT 8.400 382.050 9.450 397.950 ;
        RECT 11.400 385.050 12.450 422.400 ;
        RECT 23.400 418.050 24.450 449.400 ;
        RECT 25.950 448.950 28.050 451.050 ;
        RECT 26.400 442.050 27.450 448.950 ;
        RECT 25.950 439.950 28.050 442.050 ;
        RECT 26.400 426.450 27.450 439.950 ;
        RECT 29.400 430.050 30.450 470.400 ;
        RECT 34.950 466.950 37.050 469.050 ;
        RECT 31.950 456.450 34.050 457.050 ;
        RECT 35.400 456.450 36.450 466.950 ;
        RECT 38.400 463.050 39.450 499.950 ;
        RECT 47.400 499.050 48.450 544.950 ;
        RECT 53.400 538.050 54.450 553.950 ;
        RECT 56.400 550.050 57.450 553.950 ;
        RECT 62.400 553.050 63.450 562.950 ;
        RECT 70.950 561.450 73.050 562.050 ;
        RECT 68.400 560.400 73.050 561.450 ;
        RECT 64.950 557.250 67.050 558.150 ;
        RECT 64.950 553.950 67.050 556.050 ;
        RECT 61.950 550.950 64.050 553.050 ;
        RECT 55.950 547.950 58.050 550.050 ;
        RECT 65.400 547.050 66.450 553.950 ;
        RECT 68.400 547.050 69.450 560.400 ;
        RECT 70.950 559.950 73.050 560.400 ;
        RECT 74.250 560.250 75.750 561.150 ;
        RECT 76.950 559.950 79.050 562.050 ;
        RECT 70.950 557.850 72.750 558.750 ;
        RECT 73.950 556.950 76.050 559.050 ;
        RECT 77.250 557.850 79.050 558.750 ;
        RECT 80.400 556.050 81.450 583.950 ;
        RECT 82.950 562.950 85.050 565.050 ;
        RECT 88.950 562.950 91.050 565.050 ;
        RECT 94.950 562.950 97.050 565.050 ;
        RECT 83.400 562.050 84.450 562.950 ;
        RECT 89.400 562.050 90.450 562.950 ;
        RECT 82.950 559.950 85.050 562.050 ;
        RECT 86.250 560.250 87.750 561.150 ;
        RECT 88.950 559.950 91.050 562.050 ;
        RECT 95.400 559.050 96.450 562.950 ;
        RECT 82.950 557.850 84.750 558.750 ;
        RECT 85.950 556.950 88.050 559.050 ;
        RECT 89.250 557.850 91.050 558.750 ;
        RECT 94.950 556.950 97.050 559.050 ;
        RECT 76.950 553.950 79.050 556.050 ;
        RECT 79.950 553.950 82.050 556.050 ;
        RECT 85.950 553.950 88.050 556.050 ;
        RECT 91.950 554.250 94.050 555.150 ;
        RECT 94.950 554.850 97.050 555.750 ;
        RECT 77.400 550.050 78.450 553.950 ;
        RECT 79.950 550.950 82.050 553.050 ;
        RECT 76.950 547.950 79.050 550.050 ;
        RECT 64.950 544.950 67.050 547.050 ;
        RECT 67.950 544.950 70.050 547.050 ;
        RECT 55.950 541.950 58.050 544.050 ;
        RECT 49.950 535.950 52.050 538.050 ;
        RECT 52.950 535.950 55.050 538.050 ;
        RECT 50.400 525.450 51.450 535.950 ;
        RECT 56.400 532.050 57.450 541.950 ;
        RECT 80.400 538.050 81.450 550.950 ;
        RECT 79.950 535.950 82.050 538.050 ;
        RECT 55.950 531.450 58.050 532.050 ;
        RECT 55.950 530.400 60.450 531.450 ;
        RECT 55.950 529.950 58.050 530.400 ;
        RECT 52.950 527.250 55.050 528.150 ;
        RECT 55.950 527.850 58.050 528.750 ;
        RECT 52.950 525.450 55.050 526.050 ;
        RECT 50.400 524.400 55.050 525.450 ;
        RECT 52.950 523.950 55.050 524.400 ;
        RECT 59.400 501.450 60.450 530.400 ;
        RECT 76.950 529.950 79.050 532.050 ;
        RECT 77.400 529.050 78.450 529.950 ;
        RECT 70.950 526.950 73.050 529.050 ;
        RECT 76.950 526.950 79.050 529.050 ;
        RECT 80.250 527.250 81.750 528.150 ;
        RECT 82.950 526.950 85.050 529.050 ;
        RECT 61.950 524.250 63.750 525.150 ;
        RECT 64.950 523.950 67.050 526.050 ;
        RECT 68.250 524.250 70.050 525.150 ;
        RECT 65.250 521.850 66.750 522.750 ;
        RECT 67.950 522.450 70.050 523.050 ;
        RECT 71.400 522.450 72.450 526.950 ;
        RECT 73.950 523.950 76.050 526.050 ;
        RECT 77.250 524.850 78.750 525.750 ;
        RECT 79.950 523.950 82.050 526.050 ;
        RECT 83.250 524.850 85.050 525.750 ;
        RECT 67.950 521.400 72.450 522.450 ;
        RECT 73.950 521.850 76.050 522.750 ;
        RECT 67.950 520.950 70.050 521.400 ;
        RECT 82.950 520.950 85.050 523.050 ;
        RECT 56.400 500.400 60.450 501.450 ;
        RECT 46.950 496.950 49.050 499.050 ;
        RECT 43.950 490.950 46.050 493.050 ;
        RECT 44.400 487.050 45.450 490.950 ;
        RECT 56.400 487.050 57.450 500.400 ;
        RECT 68.400 499.050 69.450 520.950 ;
        RECT 79.950 502.950 82.050 505.050 ;
        RECT 58.950 496.950 61.050 499.050 ;
        RECT 67.950 496.950 70.050 499.050 ;
        RECT 59.400 496.050 60.450 496.950 ;
        RECT 58.950 493.950 61.050 496.050 ;
        RECT 67.950 493.950 70.050 496.050 ;
        RECT 73.950 495.300 76.050 497.400 ;
        RECT 76.950 496.950 79.050 499.050 ;
        RECT 62.250 488.250 63.750 489.150 ;
        RECT 64.950 487.950 67.050 490.050 ;
        RECT 40.950 485.250 42.750 486.150 ;
        RECT 43.950 484.950 46.050 487.050 ;
        RECT 47.250 485.250 48.750 486.150 ;
        RECT 53.250 485.250 55.050 486.150 ;
        RECT 55.950 484.950 58.050 487.050 ;
        RECT 58.950 485.850 60.750 486.750 ;
        RECT 61.950 484.950 64.050 487.050 ;
        RECT 65.250 485.850 67.050 486.750 ;
        RECT 40.950 481.950 43.050 484.050 ;
        RECT 44.250 482.850 45.750 483.750 ;
        RECT 46.950 481.950 49.050 484.050 ;
        RECT 50.250 482.850 51.750 483.750 ;
        RECT 52.950 481.950 55.050 484.050 ;
        RECT 55.950 481.950 58.050 484.050 ;
        RECT 64.950 481.950 67.050 484.050 ;
        RECT 41.400 469.050 42.450 481.950 ;
        RECT 47.400 480.450 48.450 481.950 ;
        RECT 47.400 479.400 51.450 480.450 ;
        RECT 50.400 478.050 51.450 479.400 ;
        RECT 52.950 478.950 55.050 481.050 ;
        RECT 46.950 475.950 49.050 478.050 ;
        RECT 49.950 475.950 52.050 478.050 ;
        RECT 43.950 469.950 46.050 472.050 ;
        RECT 40.950 466.950 43.050 469.050 ;
        RECT 37.950 460.950 40.050 463.050 ;
        RECT 40.950 461.400 43.050 463.500 ;
        RECT 37.950 458.250 40.050 459.150 ;
        RECT 31.950 455.400 36.450 456.450 ;
        RECT 31.950 454.950 34.050 455.400 ;
        RECT 31.950 452.850 34.050 453.750 ;
        RECT 31.950 448.950 34.050 451.050 ;
        RECT 28.950 427.950 31.050 430.050 ;
        RECT 26.400 425.400 30.450 426.450 ;
        RECT 13.950 416.250 16.050 417.150 ;
        RECT 19.950 415.950 22.050 418.050 ;
        RECT 22.950 415.950 25.050 418.050 ;
        RECT 20.400 415.050 21.450 415.950 ;
        RECT 29.400 415.050 30.450 425.400 ;
        RECT 32.400 418.050 33.450 448.950 ;
        RECT 35.400 424.050 36.450 455.400 ;
        RECT 37.950 454.950 40.050 457.050 ;
        RECT 38.400 436.050 39.450 454.950 ;
        RECT 41.550 449.400 42.750 461.400 ;
        RECT 44.400 454.050 45.450 469.950 ;
        RECT 43.950 451.950 46.050 454.050 ;
        RECT 40.950 447.300 43.050 449.400 ;
        RECT 43.950 448.950 46.050 451.050 ;
        RECT 41.550 443.700 42.750 447.300 ;
        RECT 40.950 441.600 43.050 443.700 ;
        RECT 37.950 433.950 40.050 436.050 ;
        RECT 34.950 421.950 37.050 424.050 ;
        RECT 40.950 421.950 43.050 424.050 ;
        RECT 31.950 415.950 34.050 418.050 ;
        RECT 13.950 412.950 16.050 415.050 ;
        RECT 17.250 413.250 18.750 414.150 ;
        RECT 19.950 412.950 22.050 415.050 ;
        RECT 23.250 413.250 25.050 414.150 ;
        RECT 25.950 413.250 27.750 414.150 ;
        RECT 28.950 412.950 31.050 415.050 ;
        RECT 32.250 413.250 33.750 414.150 ;
        RECT 34.950 412.950 37.050 415.050 ;
        RECT 38.250 413.250 40.050 414.150 ;
        RECT 14.400 400.050 15.450 412.950 ;
        RECT 41.400 412.050 42.450 421.950 ;
        RECT 44.400 418.050 45.450 448.950 ;
        RECT 47.400 439.050 48.450 475.950 ;
        RECT 49.950 456.450 52.050 457.050 ;
        RECT 53.400 456.450 54.450 478.950 ;
        RECT 56.400 478.050 57.450 481.950 ;
        RECT 55.950 475.950 58.050 478.050 ;
        RECT 58.950 472.950 61.050 475.050 ;
        RECT 49.950 455.400 54.450 456.450 ;
        RECT 49.950 454.950 52.050 455.400 ;
        RECT 49.950 452.850 52.050 453.750 ;
        RECT 46.950 436.950 49.050 439.050 ;
        RECT 53.400 433.050 54.450 455.400 ;
        RECT 55.950 454.950 58.050 457.050 ;
        RECT 55.950 452.850 58.050 453.750 ;
        RECT 59.400 441.450 60.450 472.950 ;
        RECT 65.400 469.050 66.450 481.950 ;
        RECT 68.400 478.050 69.450 493.950 ;
        RECT 74.550 491.700 75.750 495.300 ;
        RECT 70.950 487.950 73.050 490.050 ;
        RECT 73.950 489.600 76.050 491.700 ;
        RECT 71.400 484.050 72.450 487.950 ;
        RECT 70.950 481.950 73.050 484.050 ;
        RECT 70.950 479.850 73.050 480.750 ;
        RECT 67.950 475.950 70.050 478.050 ;
        RECT 74.550 477.600 75.750 489.600 ;
        RECT 73.950 475.500 76.050 477.600 ;
        RECT 67.950 472.950 70.050 475.050 ;
        RECT 64.950 466.950 67.050 469.050 ;
        RECT 61.950 461.400 64.050 463.500 ;
        RECT 62.400 444.600 63.600 461.400 ;
        RECT 65.400 445.050 66.450 466.950 ;
        RECT 61.950 442.500 64.050 444.600 ;
        RECT 64.950 442.950 67.050 445.050 ;
        RECT 56.400 440.400 60.450 441.450 ;
        RECT 52.950 430.950 55.050 433.050 ;
        RECT 49.950 418.950 52.050 421.050 ;
        RECT 50.400 418.050 51.450 418.950 ;
        RECT 56.400 418.050 57.450 440.400 ;
        RECT 43.950 415.950 46.050 418.050 ;
        RECT 47.250 416.250 48.750 417.150 ;
        RECT 49.950 415.950 52.050 418.050 ;
        RECT 52.950 415.950 55.050 418.050 ;
        RECT 55.950 415.950 58.050 418.050 ;
        RECT 61.950 417.450 64.050 418.050 ;
        RECT 59.400 416.400 64.050 417.450 ;
        RECT 43.950 413.850 45.750 414.750 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 50.250 413.850 52.050 414.750 ;
        RECT 16.950 409.950 19.050 412.050 ;
        RECT 20.250 410.850 21.750 411.750 ;
        RECT 22.950 409.950 25.050 412.050 ;
        RECT 25.950 409.950 28.050 412.050 ;
        RECT 29.250 410.850 30.750 411.750 ;
        RECT 31.950 409.950 34.050 412.050 ;
        RECT 35.250 410.850 36.750 411.750 ;
        RECT 37.950 409.950 40.050 412.050 ;
        RECT 40.950 409.950 43.050 412.050 ;
        RECT 13.950 397.950 16.050 400.050 ;
        RECT 13.950 391.950 16.050 394.050 ;
        RECT 10.950 382.950 13.050 385.050 ;
        RECT 7.950 379.950 10.050 382.050 ;
        RECT 11.250 380.250 13.050 381.150 ;
        RECT 1.950 377.850 3.750 378.750 ;
        RECT 4.950 376.950 7.050 379.050 ;
        RECT 8.250 377.850 9.750 378.750 ;
        RECT 10.950 376.950 13.050 379.050 ;
        RECT 1.950 373.950 4.050 376.050 ;
        RECT 4.950 374.850 7.050 375.750 ;
        RECT 2.400 349.050 3.450 373.950 ;
        RECT 4.950 358.950 7.050 361.050 ;
        RECT 5.400 349.050 6.450 358.950 ;
        RECT 11.400 351.450 12.450 376.950 ;
        RECT 14.400 354.450 15.450 391.950 ;
        RECT 23.400 391.050 24.450 409.950 ;
        RECT 26.400 394.050 27.450 409.950 ;
        RECT 28.950 406.950 31.050 409.050 ;
        RECT 29.400 402.450 30.450 406.950 ;
        RECT 32.400 406.050 33.450 409.950 ;
        RECT 43.950 406.950 46.050 409.050 ;
        RECT 31.950 403.950 34.050 406.050 ;
        RECT 29.400 401.400 33.450 402.450 ;
        RECT 25.950 391.950 28.050 394.050 ;
        RECT 22.950 388.950 25.050 391.050 ;
        RECT 19.950 385.950 22.050 388.050 ;
        RECT 16.950 383.250 19.050 384.150 ;
        RECT 19.950 383.850 22.050 384.750 ;
        RECT 25.950 384.450 28.050 385.050 ;
        RECT 22.950 383.250 24.750 384.150 ;
        RECT 25.950 383.400 30.450 384.450 ;
        RECT 25.950 382.950 28.050 383.400 ;
        RECT 16.950 379.950 19.050 382.050 ;
        RECT 22.950 379.950 25.050 382.050 ;
        RECT 26.250 380.850 28.050 381.750 ;
        RECT 14.400 353.400 18.450 354.450 ;
        RECT 11.400 350.400 15.450 351.450 ;
        RECT 14.400 349.050 15.450 350.400 ;
        RECT 1.950 346.950 4.050 349.050 ;
        RECT 4.950 346.950 7.050 349.050 ;
        RECT 10.950 347.250 13.050 348.150 ;
        RECT 13.950 346.950 16.050 349.050 ;
        RECT 4.950 345.450 7.050 346.050 ;
        RECT 2.400 344.400 7.050 345.450 ;
        RECT 2.400 328.050 3.450 344.400 ;
        RECT 4.950 343.950 7.050 344.400 ;
        RECT 8.250 344.250 9.750 345.150 ;
        RECT 10.950 343.950 13.050 346.050 ;
        RECT 14.250 344.250 16.050 345.150 ;
        RECT 4.950 341.850 6.750 342.750 ;
        RECT 7.950 340.950 10.050 343.050 ;
        RECT 11.400 340.050 12.450 343.950 ;
        RECT 13.950 340.950 16.050 343.050 ;
        RECT 4.950 337.950 7.050 340.050 ;
        RECT 10.950 339.450 13.050 340.050 ;
        RECT 8.400 338.400 13.050 339.450 ;
        RECT 1.950 325.950 4.050 328.050 ;
        RECT 2.400 301.050 3.450 325.950 ;
        RECT 5.400 313.050 6.450 337.950 ;
        RECT 8.400 316.050 9.450 338.400 ;
        RECT 10.950 337.950 13.050 338.400 ;
        RECT 13.950 337.950 16.050 340.050 ;
        RECT 7.950 313.950 10.050 316.050 ;
        RECT 4.950 310.950 7.050 313.050 ;
        RECT 7.950 310.950 10.050 313.050 ;
        RECT 4.950 308.850 7.050 309.750 ;
        RECT 1.950 298.950 4.050 301.050 ;
        RECT 1.950 280.950 4.050 283.050 ;
        RECT 2.400 259.050 3.450 280.950 ;
        RECT 4.950 277.950 7.050 280.050 ;
        RECT 5.400 273.450 6.450 277.950 ;
        RECT 8.400 277.050 9.450 310.950 ;
        RECT 10.950 308.850 13.050 309.750 ;
        RECT 14.400 309.450 15.450 337.950 ;
        RECT 17.400 313.050 18.450 353.400 ;
        RECT 19.950 352.950 22.050 355.050 ;
        RECT 20.400 352.050 21.450 352.950 ;
        RECT 19.950 349.950 22.050 352.050 ;
        RECT 29.400 346.050 30.450 383.400 ;
        RECT 32.400 361.050 33.450 401.400 ;
        RECT 37.950 388.950 40.050 391.050 ;
        RECT 38.400 388.050 39.450 388.950 ;
        RECT 37.950 385.950 40.050 388.050 ;
        RECT 44.400 385.050 45.450 406.950 ;
        RECT 47.400 400.050 48.450 412.950 ;
        RECT 53.400 409.050 54.450 415.950 ;
        RECT 59.400 415.050 60.450 416.400 ;
        RECT 61.950 415.950 64.050 416.400 ;
        RECT 55.950 413.250 58.050 414.150 ;
        RECT 58.950 412.950 61.050 415.050 ;
        RECT 61.950 413.850 64.050 414.750 ;
        RECT 64.950 413.250 67.050 414.150 ;
        RECT 55.950 409.950 58.050 412.050 ;
        RECT 52.950 406.950 55.050 409.050 ;
        RECT 59.400 408.450 60.450 412.950 ;
        RECT 61.950 409.950 64.050 412.050 ;
        RECT 64.950 409.950 67.050 412.050 ;
        RECT 56.400 407.400 60.450 408.450 ;
        RECT 49.950 403.950 52.050 406.050 ;
        RECT 46.950 397.950 49.050 400.050 ;
        RECT 34.950 383.250 37.050 384.150 ;
        RECT 37.950 383.850 40.050 384.750 ;
        RECT 43.950 384.450 46.050 385.050 ;
        RECT 41.400 383.400 46.050 384.450 ;
        RECT 34.950 379.950 37.050 382.050 ;
        RECT 37.950 379.950 40.050 382.050 ;
        RECT 31.950 358.950 34.050 361.050 ;
        RECT 19.950 344.250 22.050 345.150 ;
        RECT 28.950 343.950 31.050 346.050 ;
        RECT 38.400 345.450 39.450 379.950 ;
        RECT 41.400 355.050 42.450 383.400 ;
        RECT 43.950 382.950 46.050 383.400 ;
        RECT 43.950 380.850 46.050 381.750 ;
        RECT 46.950 380.250 49.050 381.150 ;
        RECT 46.950 376.950 49.050 379.050 ;
        RECT 50.400 370.050 51.450 403.950 ;
        RECT 52.950 391.950 55.050 394.050 ;
        RECT 53.400 385.050 54.450 391.950 ;
        RECT 52.950 382.950 55.050 385.050 ;
        RECT 52.950 380.850 55.050 381.750 ;
        RECT 56.400 379.050 57.450 407.400 ;
        RECT 62.400 400.050 63.450 409.950 ;
        RECT 61.950 397.950 64.050 400.050 ;
        RECT 64.950 391.950 67.050 394.050 ;
        RECT 65.400 388.050 66.450 391.950 ;
        RECT 68.400 388.050 69.450 472.950 ;
        RECT 70.950 463.950 73.050 466.050 ;
        RECT 71.400 457.050 72.450 463.950 ;
        RECT 77.400 463.050 78.450 496.950 ;
        RECT 76.950 460.950 79.050 463.050 ;
        RECT 80.400 460.050 81.450 502.950 ;
        RECT 83.400 496.050 84.450 520.950 ;
        RECT 82.950 493.950 85.050 496.050 ;
        RECT 82.950 485.250 85.050 486.150 ;
        RECT 82.950 481.950 85.050 484.050 ;
        RECT 83.400 481.050 84.450 481.950 ;
        RECT 82.950 478.950 85.050 481.050 ;
        RECT 86.400 475.050 87.450 553.950 ;
        RECT 91.950 550.950 94.050 553.050 ;
        RECT 98.400 552.450 99.450 589.950 ;
        RECT 104.400 589.050 105.450 622.950 ;
        RECT 116.400 622.050 117.450 628.950 ;
        RECT 122.400 628.050 123.450 628.950 ;
        RECT 128.400 628.050 129.450 632.400 ;
        RECT 121.950 625.950 124.050 628.050 ;
        RECT 127.950 625.950 130.050 628.050 ;
        RECT 131.400 625.050 132.450 662.400 ;
        RECT 136.950 661.950 139.050 664.050 ;
        RECT 143.400 655.050 144.450 664.950 ;
        RECT 151.950 662.850 154.050 663.750 ;
        RECT 158.400 661.050 159.450 664.950 ;
        RECT 157.950 658.950 160.050 661.050 ;
        RECT 161.400 655.050 162.450 673.950 ;
        RECT 163.950 671.250 166.050 672.150 ;
        RECT 166.950 671.850 169.050 672.750 ;
        RECT 169.950 671.250 171.750 672.150 ;
        RECT 172.950 670.950 175.050 673.050 ;
        RECT 175.950 670.950 178.050 673.050 ;
        RECT 163.950 667.950 166.050 670.050 ;
        RECT 169.950 667.950 172.050 670.050 ;
        RECT 173.250 668.850 175.050 669.750 ;
        RECT 164.400 664.050 165.450 667.950 ;
        RECT 170.400 667.050 171.450 667.950 ;
        RECT 169.950 664.950 172.050 667.050 ;
        RECT 176.400 664.050 177.450 670.950 ;
        RECT 185.400 670.050 186.450 682.950 ;
        RECT 193.950 679.950 196.050 682.050 ;
        RECT 217.950 679.950 220.050 682.050 ;
        RECT 190.950 673.950 193.050 676.050 ;
        RECT 191.400 670.050 192.450 673.950 ;
        RECT 194.400 673.050 195.450 679.950 ;
        RECT 214.950 676.950 217.050 679.050 ;
        RECT 196.950 673.950 199.050 676.050 ;
        RECT 202.950 673.950 205.050 676.050 ;
        RECT 193.950 670.950 196.050 673.050 ;
        RECT 197.250 671.850 198.750 672.750 ;
        RECT 199.950 670.950 202.050 673.050 ;
        RECT 178.950 667.950 181.050 670.050 ;
        RECT 181.950 668.250 183.750 669.150 ;
        RECT 184.950 667.950 187.050 670.050 ;
        RECT 188.250 668.250 190.050 669.150 ;
        RECT 190.950 667.950 193.050 670.050 ;
        RECT 193.950 668.850 196.050 669.750 ;
        RECT 199.950 668.850 202.050 669.750 ;
        RECT 163.950 661.950 166.050 664.050 ;
        RECT 175.950 661.950 178.050 664.050 ;
        RECT 136.950 652.950 139.050 655.050 ;
        RECT 142.950 652.950 145.050 655.050 ;
        RECT 160.950 652.950 163.050 655.050 ;
        RECT 172.950 652.950 175.050 655.050 ;
        RECT 137.400 634.050 138.450 652.950 ;
        RECT 157.950 635.250 160.050 636.150 ;
        RECT 166.950 635.250 169.050 636.150 ;
        RECT 173.400 634.050 174.450 652.950 ;
        RECT 136.950 631.950 139.050 634.050 ;
        RECT 151.950 633.450 154.050 634.050 ;
        RECT 149.400 632.400 154.050 633.450 ;
        RECT 137.400 631.050 138.450 631.950 ;
        RECT 133.950 629.250 135.750 630.150 ;
        RECT 136.950 628.950 139.050 631.050 ;
        RECT 140.250 629.250 141.750 630.150 ;
        RECT 142.950 628.950 145.050 631.050 ;
        RECT 146.250 629.250 148.050 630.150 ;
        RECT 133.950 625.950 136.050 628.050 ;
        RECT 137.250 626.850 138.750 627.750 ;
        RECT 139.950 625.950 142.050 628.050 ;
        RECT 143.250 626.850 144.750 627.750 ;
        RECT 145.950 627.450 148.050 628.050 ;
        RECT 149.400 627.450 150.450 632.400 ;
        RECT 151.950 631.950 154.050 632.400 ;
        RECT 155.250 632.250 156.750 633.150 ;
        RECT 157.950 631.950 160.050 634.050 ;
        RECT 161.250 632.250 163.050 633.150 ;
        RECT 163.950 632.250 165.750 633.150 ;
        RECT 166.950 631.950 169.050 634.050 ;
        RECT 170.250 632.250 171.750 633.150 ;
        RECT 172.950 631.950 175.050 634.050 ;
        RECT 179.400 633.450 180.450 667.950 ;
        RECT 181.950 664.950 184.050 667.050 ;
        RECT 185.250 665.850 186.750 666.750 ;
        RECT 187.950 664.950 190.050 667.050 ;
        RECT 182.400 658.050 183.450 664.950 ;
        RECT 188.400 661.050 189.450 664.950 ;
        RECT 203.400 664.050 204.450 673.950 ;
        RECT 215.400 673.050 216.450 676.950 ;
        RECT 218.400 676.050 219.450 679.950 ;
        RECT 217.950 673.950 220.050 676.050 ;
        RECT 208.950 670.950 211.050 673.050 ;
        RECT 212.250 671.250 213.750 672.150 ;
        RECT 214.950 670.950 217.050 673.050 ;
        RECT 205.950 667.950 208.050 670.050 ;
        RECT 209.250 668.850 210.750 669.750 ;
        RECT 211.950 667.950 214.050 670.050 ;
        RECT 215.250 668.850 217.050 669.750 ;
        RECT 205.950 665.850 208.050 666.750 ;
        RECT 202.950 661.950 205.050 664.050 ;
        RECT 212.400 661.050 213.450 667.950 ;
        RECT 218.400 666.450 219.450 673.950 ;
        RECT 230.400 673.050 231.450 682.950 ;
        RECT 244.950 679.950 247.050 682.050 ;
        RECT 340.950 679.950 343.050 682.050 ;
        RECT 349.950 679.950 352.050 682.050 ;
        RECT 499.950 679.950 502.050 682.050 ;
        RECT 514.950 679.950 517.050 682.050 ;
        RECT 241.950 676.950 244.050 679.050 ;
        RECT 232.950 673.950 235.050 676.050 ;
        RECT 223.950 670.950 226.050 673.050 ;
        RECT 229.950 670.950 232.050 673.050 ;
        RECT 233.250 671.850 234.750 672.750 ;
        RECT 235.950 670.950 238.050 673.050 ;
        RECT 224.400 670.050 225.450 670.950 ;
        RECT 242.400 670.050 243.450 676.950 ;
        RECT 220.950 668.250 222.750 669.150 ;
        RECT 223.950 667.950 226.050 670.050 ;
        RECT 227.250 668.250 229.050 669.150 ;
        RECT 229.950 668.850 232.050 669.750 ;
        RECT 232.950 667.950 235.050 670.050 ;
        RECT 235.950 668.850 238.050 669.750 ;
        RECT 238.950 667.950 241.050 670.050 ;
        RECT 241.950 667.950 244.050 670.050 ;
        RECT 220.950 666.450 223.050 667.050 ;
        RECT 218.400 665.400 223.050 666.450 ;
        RECT 224.250 665.850 225.750 666.750 ;
        RECT 220.950 664.950 223.050 665.400 ;
        RECT 226.950 664.950 229.050 667.050 ;
        RECT 233.400 661.050 234.450 667.950 ;
        RECT 239.400 664.050 240.450 667.950 ;
        RECT 245.400 667.050 246.450 679.950 ;
        RECT 253.950 676.950 256.050 679.050 ;
        RECT 271.950 676.950 274.050 679.050 ;
        RECT 292.950 676.950 295.050 679.050 ;
        RECT 301.950 676.950 304.050 679.050 ;
        RECT 307.950 676.950 310.050 679.050 ;
        RECT 247.950 667.950 250.050 670.050 ;
        RECT 251.250 668.250 253.050 669.150 ;
        RECT 254.400 667.050 255.450 676.950 ;
        RECT 272.400 676.050 273.450 676.950 ;
        RECT 293.400 676.050 294.450 676.950 ;
        RECT 265.950 673.950 268.050 676.050 ;
        RECT 271.950 673.950 274.050 676.050 ;
        RECT 286.950 673.950 289.050 676.050 ;
        RECT 292.950 673.950 295.050 676.050 ;
        RECT 259.950 672.450 262.050 673.050 ;
        RECT 257.400 671.400 262.050 672.450 ;
        RECT 241.950 665.850 243.750 666.750 ;
        RECT 244.950 664.950 247.050 667.050 ;
        RECT 248.250 665.850 249.750 666.750 ;
        RECT 250.950 664.950 253.050 667.050 ;
        RECT 253.950 664.950 256.050 667.050 ;
        RECT 238.950 661.950 241.050 664.050 ;
        RECT 244.950 662.850 247.050 663.750 ;
        RECT 187.950 658.950 190.050 661.050 ;
        RECT 211.950 658.950 214.050 661.050 ;
        RECT 232.950 658.950 235.050 661.050 ;
        RECT 181.950 655.950 184.050 658.050 ;
        RECT 251.400 640.050 252.450 664.950 ;
        RECT 250.950 637.950 253.050 640.050 ;
        RECT 199.950 635.250 202.050 636.150 ;
        RECT 208.950 634.950 211.050 637.050 ;
        RECT 220.950 635.250 223.050 636.150 ;
        RECT 232.950 634.950 235.050 637.050 ;
        RECT 209.400 634.050 210.450 634.950 ;
        RECT 181.950 633.450 184.050 634.050 ;
        RECT 179.400 632.400 184.050 633.450 ;
        RECT 187.950 633.450 190.050 634.050 ;
        RECT 151.950 629.850 153.750 630.750 ;
        RECT 154.950 628.950 157.050 631.050 ;
        RECT 145.950 626.400 150.450 627.450 ;
        RECT 145.950 625.950 148.050 626.400 ;
        RECT 140.400 625.050 141.450 625.950 ;
        RECT 130.950 622.950 133.050 625.050 ;
        RECT 139.950 622.950 142.050 625.050 ;
        RECT 155.400 622.050 156.450 628.950 ;
        RECT 115.950 619.950 118.050 622.050 ;
        RECT 133.950 619.950 136.050 622.050 ;
        RECT 154.950 619.950 157.050 622.050 ;
        RECT 106.950 601.950 109.050 604.050 ;
        RECT 107.400 594.450 108.450 601.950 ;
        RECT 116.400 601.050 117.450 619.950 ;
        RECT 118.950 607.950 121.050 610.050 ;
        RECT 115.950 598.950 118.050 601.050 ;
        RECT 119.400 598.050 120.450 607.950 ;
        RECT 127.950 604.950 130.050 607.050 ;
        RECT 128.400 598.050 129.450 604.950 ;
        RECT 109.950 596.250 111.750 597.150 ;
        RECT 112.950 595.950 115.050 598.050 ;
        RECT 118.950 595.950 121.050 598.050 ;
        RECT 121.950 595.950 124.050 598.050 ;
        RECT 127.950 595.950 130.050 598.050 ;
        RECT 131.250 596.250 133.050 597.150 ;
        RECT 109.950 594.450 112.050 595.050 ;
        RECT 107.400 593.400 112.050 594.450 ;
        RECT 113.250 593.850 114.750 594.750 ;
        RECT 109.950 592.950 112.050 593.400 ;
        RECT 115.950 592.950 118.050 595.050 ;
        RECT 119.250 593.850 121.050 594.750 ;
        RECT 121.950 593.850 123.750 594.750 ;
        RECT 124.950 592.950 127.050 595.050 ;
        RECT 128.250 593.850 129.750 594.750 ;
        RECT 130.950 594.450 133.050 595.050 ;
        RECT 134.400 594.450 135.450 619.950 ;
        RECT 139.950 604.950 142.050 607.050 ;
        RECT 142.950 604.950 145.050 607.050 ;
        RECT 140.400 598.050 141.450 604.950 ;
        RECT 143.400 601.050 144.450 604.950 ;
        RECT 158.400 601.050 159.450 631.950 ;
        RECT 160.950 628.950 163.050 631.050 ;
        RECT 163.950 630.450 166.050 631.050 ;
        RECT 163.950 629.400 168.450 630.450 ;
        RECT 163.950 628.950 166.050 629.400 ;
        RECT 161.400 619.050 162.450 628.950 ;
        RECT 163.950 625.950 166.050 628.050 ;
        RECT 160.950 616.950 163.050 619.050 ;
        RECT 160.950 607.950 163.050 610.050 ;
        RECT 142.950 598.950 145.050 601.050 ;
        RECT 146.250 599.250 147.750 600.150 ;
        RECT 148.950 598.950 151.050 601.050 ;
        RECT 151.950 598.950 154.050 601.050 ;
        RECT 155.250 599.250 156.750 600.150 ;
        RECT 157.950 598.950 160.050 601.050 ;
        RECT 161.400 598.050 162.450 607.950 ;
        RECT 139.950 595.950 142.050 598.050 ;
        RECT 143.250 596.850 144.750 597.750 ;
        RECT 145.950 595.950 148.050 598.050 ;
        RECT 149.250 596.850 151.050 597.750 ;
        RECT 151.950 596.850 153.750 597.750 ;
        RECT 154.950 595.950 157.050 598.050 ;
        RECT 158.250 596.850 159.750 597.750 ;
        RECT 160.950 595.950 163.050 598.050 ;
        RECT 130.950 593.400 135.450 594.450 ;
        RECT 139.950 593.850 142.050 594.750 ;
        RECT 130.950 592.950 133.050 593.400 ;
        RECT 145.950 592.950 148.050 595.050 ;
        RECT 112.950 589.950 115.050 592.050 ;
        RECT 115.950 590.850 118.050 591.750 ;
        RECT 124.950 590.850 127.050 591.750 ;
        RECT 130.950 589.950 133.050 592.050 ;
        RECT 103.950 586.950 106.050 589.050 ;
        RECT 113.400 565.050 114.450 589.950 ;
        RECT 127.950 586.950 130.050 589.050 ;
        RECT 124.950 565.950 127.050 568.050 ;
        RECT 112.950 562.950 115.050 565.050 ;
        RECT 115.950 561.450 118.050 562.050 ;
        RECT 109.950 560.250 112.050 561.150 ;
        RECT 113.400 560.400 118.050 561.450 ;
        RECT 121.950 561.450 124.050 562.050 ;
        RECT 125.400 561.450 126.450 565.950 ;
        RECT 100.950 557.250 102.750 558.150 ;
        RECT 103.950 556.950 106.050 559.050 ;
        RECT 107.250 557.250 108.750 558.150 ;
        RECT 109.950 556.950 112.050 559.050 ;
        RECT 113.400 556.050 114.450 560.400 ;
        RECT 115.950 559.950 118.050 560.400 ;
        RECT 119.250 560.250 120.750 561.150 ;
        RECT 121.950 560.400 126.450 561.450 ;
        RECT 121.950 559.950 124.050 560.400 ;
        RECT 115.950 557.850 117.750 558.750 ;
        RECT 118.950 556.950 121.050 559.050 ;
        RECT 122.250 557.850 124.050 558.750 ;
        RECT 100.950 553.950 103.050 556.050 ;
        RECT 104.250 554.850 105.750 555.750 ;
        RECT 106.950 555.450 109.050 556.050 ;
        RECT 109.950 555.450 112.050 556.050 ;
        RECT 106.950 554.400 112.050 555.450 ;
        RECT 106.950 553.950 109.050 554.400 ;
        RECT 109.950 553.950 112.050 554.400 ;
        RECT 112.950 553.950 115.050 556.050 ;
        RECT 125.400 553.050 126.450 560.400 ;
        RECT 98.400 551.400 102.450 552.450 ;
        RECT 88.950 535.950 91.050 538.050 ;
        RECT 89.400 526.050 90.450 535.950 ;
        RECT 92.400 529.050 93.450 550.950 ;
        RECT 97.950 538.950 100.050 541.050 ;
        RECT 98.400 529.050 99.450 538.950 ;
        RECT 101.400 535.050 102.450 551.400 ;
        RECT 103.950 550.950 106.050 553.050 ;
        RECT 124.950 550.950 127.050 553.050 ;
        RECT 104.400 544.050 105.450 550.950 ;
        RECT 118.950 544.950 121.050 547.050 ;
        RECT 103.950 541.950 106.050 544.050 ;
        RECT 112.950 541.950 115.050 544.050 ;
        RECT 100.950 532.950 103.050 535.050 ;
        RECT 109.950 532.950 112.050 535.050 ;
        RECT 91.950 526.950 94.050 529.050 ;
        RECT 95.250 527.250 96.750 528.150 ;
        RECT 97.950 526.950 100.050 529.050 ;
        RECT 88.950 523.950 91.050 526.050 ;
        RECT 92.250 524.850 93.750 525.750 ;
        RECT 94.950 523.950 97.050 526.050 ;
        RECT 98.250 524.850 100.050 525.750 ;
        RECT 100.950 524.250 102.750 525.150 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 107.250 524.250 109.050 525.150 ;
        RECT 88.950 521.850 91.050 522.750 ;
        RECT 91.950 508.950 94.050 511.050 ;
        RECT 88.950 493.950 91.050 496.050 ;
        RECT 89.400 490.050 90.450 493.950 ;
        RECT 88.950 487.950 91.050 490.050 ;
        RECT 88.950 485.250 91.050 486.150 ;
        RECT 88.950 481.950 91.050 484.050 ;
        RECT 88.950 475.950 91.050 478.050 ;
        RECT 85.950 472.950 88.050 475.050 ;
        RECT 89.400 466.050 90.450 475.950 ;
        RECT 92.400 475.050 93.450 508.950 ;
        RECT 95.400 502.050 96.450 523.950 ;
        RECT 104.250 521.850 105.750 522.750 ;
        RECT 106.950 520.950 109.050 523.050 ;
        RECT 103.950 517.950 106.050 520.050 ;
        RECT 100.950 502.950 103.050 505.050 ;
        RECT 94.950 499.950 97.050 502.050 ;
        RECT 94.950 494.400 97.050 496.500 ;
        RECT 95.400 477.600 96.600 494.400 ;
        RECT 97.950 487.950 100.050 490.050 ;
        RECT 98.400 478.050 99.450 487.950 ;
        RECT 94.950 475.500 97.050 477.600 ;
        RECT 97.950 475.950 100.050 478.050 ;
        RECT 91.950 472.950 94.050 475.050 ;
        RECT 97.950 472.950 100.050 475.050 ;
        RECT 94.950 469.950 97.050 472.050 ;
        RECT 82.950 463.950 85.050 466.050 ;
        RECT 85.950 463.950 88.050 466.050 ;
        RECT 88.950 463.950 91.050 466.050 ;
        RECT 79.950 457.950 82.050 460.050 ;
        RECT 70.950 454.950 73.050 457.050 ;
        RECT 74.250 455.250 75.750 456.150 ;
        RECT 76.950 454.950 79.050 457.050 ;
        RECT 70.950 452.850 72.750 453.750 ;
        RECT 73.950 451.950 76.050 454.050 ;
        RECT 77.250 452.850 78.750 453.750 ;
        RECT 79.950 451.950 82.050 454.050 ;
        RECT 70.950 445.950 73.050 448.050 ;
        RECT 64.950 385.950 67.050 388.050 ;
        RECT 67.950 385.950 70.050 388.050 ;
        RECT 58.950 382.950 61.050 385.050 ;
        RECT 62.250 383.250 64.050 384.150 ;
        RECT 64.950 383.850 67.050 384.750 ;
        RECT 67.950 383.250 70.050 384.150 ;
        RECT 58.950 380.850 60.750 381.750 ;
        RECT 61.950 379.950 64.050 382.050 ;
        RECT 64.950 379.950 67.050 382.050 ;
        RECT 67.950 379.950 70.050 382.050 ;
        RECT 52.950 376.950 55.050 379.050 ;
        RECT 55.950 376.950 58.050 379.050 ;
        RECT 49.950 367.950 52.050 370.050 ;
        RECT 40.950 352.950 43.050 355.050 ;
        RECT 46.950 352.950 49.050 355.050 ;
        RECT 47.400 349.050 48.450 352.950 ;
        RECT 53.400 349.050 54.450 376.950 ;
        RECT 61.950 361.950 64.050 364.050 ;
        RECT 62.400 352.050 63.450 361.950 ;
        RECT 61.950 349.950 64.050 352.050 ;
        RECT 46.950 346.950 49.050 349.050 ;
        RECT 49.950 347.250 52.050 348.150 ;
        RECT 52.950 346.950 55.050 349.050 ;
        RECT 35.400 344.400 39.450 345.450 ;
        RECT 35.400 343.050 36.450 344.400 ;
        RECT 40.950 344.250 43.050 345.150 ;
        RECT 43.950 343.950 46.050 346.050 ;
        RECT 46.950 344.250 48.750 345.150 ;
        RECT 49.950 343.950 52.050 346.050 ;
        RECT 55.950 345.450 58.050 346.050 ;
        RECT 53.250 344.250 54.750 345.150 ;
        RECT 55.950 344.400 60.450 345.450 ;
        RECT 55.950 343.950 58.050 344.400 ;
        RECT 19.950 340.950 22.050 343.050 ;
        RECT 23.250 341.250 24.750 342.150 ;
        RECT 25.950 340.950 28.050 343.050 ;
        RECT 29.250 341.250 31.050 342.150 ;
        RECT 31.950 341.250 33.750 342.150 ;
        RECT 34.950 340.950 37.050 343.050 ;
        RECT 38.250 341.250 39.750 342.150 ;
        RECT 40.950 340.950 43.050 343.050 ;
        RECT 20.400 340.050 21.450 340.950 ;
        RECT 19.950 337.950 22.050 340.050 ;
        RECT 22.950 337.950 25.050 340.050 ;
        RECT 26.250 338.850 27.750 339.750 ;
        RECT 28.950 337.950 31.050 340.050 ;
        RECT 31.950 337.950 34.050 340.050 ;
        RECT 35.250 338.850 36.750 339.750 ;
        RECT 37.950 337.950 40.050 340.050 ;
        RECT 23.400 331.050 24.450 337.950 ;
        RECT 29.400 337.050 30.450 337.950 ;
        RECT 32.400 337.050 33.450 337.950 ;
        RECT 28.950 334.950 31.050 337.050 ;
        RECT 31.950 334.950 34.050 337.050 ;
        RECT 31.950 331.950 34.050 334.050 ;
        RECT 34.950 331.950 37.050 334.050 ;
        RECT 22.950 328.950 25.050 331.050 ;
        RECT 25.950 319.950 28.050 322.050 ;
        RECT 26.400 313.050 27.450 319.950 ;
        RECT 32.400 313.050 33.450 331.950 ;
        RECT 35.400 313.050 36.450 331.950 ;
        RECT 38.400 313.050 39.450 337.950 ;
        RECT 41.400 334.050 42.450 340.950 ;
        RECT 44.400 337.050 45.450 343.950 ;
        RECT 46.950 340.950 49.050 343.050 ;
        RECT 50.400 340.050 51.450 343.950 ;
        RECT 52.950 340.950 55.050 343.050 ;
        RECT 56.250 341.850 58.050 342.750 ;
        RECT 49.950 337.950 52.050 340.050 ;
        RECT 55.950 337.950 58.050 340.050 ;
        RECT 50.400 337.050 51.450 337.950 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 49.950 334.950 52.050 337.050 ;
        RECT 40.950 331.950 43.050 334.050 ;
        RECT 52.950 328.950 55.050 331.050 ;
        RECT 46.950 325.950 49.050 328.050 ;
        RECT 40.950 322.950 43.050 325.050 ;
        RECT 16.950 310.950 19.050 313.050 ;
        RECT 19.950 310.950 22.050 313.050 ;
        RECT 23.250 311.250 24.750 312.150 ;
        RECT 25.950 310.950 28.050 313.050 ;
        RECT 31.950 310.950 34.050 313.050 ;
        RECT 34.950 310.950 37.050 313.050 ;
        RECT 37.950 310.950 40.050 313.050 ;
        RECT 16.950 309.450 19.050 310.050 ;
        RECT 14.400 308.400 19.050 309.450 ;
        RECT 20.250 308.850 21.750 309.750 ;
        RECT 16.950 307.950 19.050 308.400 ;
        RECT 22.950 307.950 25.050 310.050 ;
        RECT 26.250 308.850 28.050 309.750 ;
        RECT 34.950 309.450 37.050 310.050 ;
        RECT 38.400 309.450 39.450 310.950 ;
        RECT 41.400 310.050 42.450 322.950 ;
        RECT 47.400 316.050 48.450 325.950 ;
        RECT 53.400 316.050 54.450 328.950 ;
        RECT 46.950 313.950 49.050 316.050 ;
        RECT 52.950 313.950 55.050 316.050 ;
        RECT 43.950 311.250 46.050 312.150 ;
        RECT 46.950 311.850 49.050 312.750 ;
        RECT 49.950 311.250 51.750 312.150 ;
        RECT 52.950 310.950 55.050 313.050 ;
        RECT 31.950 308.250 33.750 309.150 ;
        RECT 34.950 308.400 39.450 309.450 ;
        RECT 34.950 307.950 37.050 308.400 ;
        RECT 40.950 307.950 43.050 310.050 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 49.950 307.950 52.050 310.050 ;
        RECT 53.250 308.850 55.050 309.750 ;
        RECT 10.950 304.950 13.050 307.050 ;
        RECT 13.950 304.950 16.050 307.050 ;
        RECT 16.950 305.850 19.050 306.750 ;
        RECT 7.950 274.950 10.050 277.050 ;
        RECT 11.400 274.050 12.450 304.950 ;
        RECT 14.400 283.050 15.450 304.950 ;
        RECT 16.950 298.950 19.050 301.050 ;
        RECT 13.950 280.950 16.050 283.050 ;
        RECT 17.400 277.050 18.450 298.950 ;
        RECT 16.950 274.950 19.050 277.050 ;
        RECT 5.400 272.400 9.450 273.450 ;
        RECT 8.400 271.050 9.450 272.400 ;
        RECT 10.950 271.950 13.050 274.050 ;
        RECT 13.950 271.950 16.050 274.050 ;
        RECT 14.400 271.050 15.450 271.950 ;
        RECT 23.400 271.050 24.450 307.950 ;
        RECT 50.400 307.050 51.450 307.950 ;
        RECT 25.950 304.950 28.050 307.050 ;
        RECT 31.950 304.950 34.050 307.050 ;
        RECT 35.250 305.850 36.750 306.750 ;
        RECT 37.950 304.950 40.050 307.050 ;
        RECT 41.250 305.850 43.050 306.750 ;
        RECT 49.950 304.950 52.050 307.050 ;
        RECT 26.400 298.050 27.450 304.950 ;
        RECT 25.950 295.950 28.050 298.050 ;
        RECT 32.400 295.050 33.450 304.950 ;
        RECT 34.950 301.950 37.050 304.050 ;
        RECT 37.950 302.850 40.050 303.750 ;
        RECT 31.950 292.950 34.050 295.050 ;
        RECT 35.400 292.050 36.450 301.950 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 43.950 289.950 46.050 292.050 ;
        RECT 34.950 286.950 37.050 289.050 ;
        RECT 31.950 277.950 34.050 280.050 ;
        RECT 32.400 277.050 33.450 277.950 ;
        RECT 35.400 277.050 36.450 286.950 ;
        RECT 44.400 282.450 45.450 289.950 ;
        RECT 44.400 281.400 48.450 282.450 ;
        RECT 43.950 277.950 46.050 280.050 ;
        RECT 31.950 274.950 34.050 277.050 ;
        RECT 34.950 274.950 37.050 277.050 ;
        RECT 35.400 274.050 36.450 274.950 ;
        RECT 28.950 272.250 31.050 273.150 ;
        RECT 31.950 271.950 34.050 274.050 ;
        RECT 34.950 271.950 37.050 274.050 ;
        RECT 40.950 273.450 43.050 274.050 ;
        RECT 44.400 273.450 45.450 277.950 ;
        RECT 38.250 272.250 39.750 273.150 ;
        RECT 40.950 272.400 45.450 273.450 ;
        RECT 40.950 271.950 43.050 272.400 ;
        RECT 4.950 269.250 6.750 270.150 ;
        RECT 7.950 268.950 10.050 271.050 ;
        RECT 11.250 269.250 12.750 270.150 ;
        RECT 13.950 268.950 16.050 271.050 ;
        RECT 17.250 269.250 19.050 270.150 ;
        RECT 19.950 269.250 21.750 270.150 ;
        RECT 22.950 268.950 25.050 271.050 ;
        RECT 26.250 269.250 27.750 270.150 ;
        RECT 28.950 268.950 31.050 271.050 ;
        RECT 4.950 265.950 7.050 268.050 ;
        RECT 8.250 266.850 9.750 267.750 ;
        RECT 10.950 265.950 13.050 268.050 ;
        RECT 14.250 266.850 15.750 267.750 ;
        RECT 16.950 265.950 19.050 268.050 ;
        RECT 19.950 265.950 22.050 268.050 ;
        RECT 23.250 266.850 24.750 267.750 ;
        RECT 25.950 265.950 28.050 268.050 ;
        RECT 28.950 265.950 31.050 268.050 ;
        RECT 5.400 262.050 6.450 265.950 ;
        RECT 13.950 262.950 16.050 265.050 ;
        RECT 4.950 259.950 7.050 262.050 ;
        RECT 1.950 256.950 4.050 259.050 ;
        RECT 14.400 244.050 15.450 262.950 ;
        RECT 17.400 256.050 18.450 265.950 ;
        RECT 20.400 259.050 21.450 265.950 ;
        RECT 26.400 262.050 27.450 265.950 ;
        RECT 25.950 259.950 28.050 262.050 ;
        RECT 19.950 256.950 22.050 259.050 ;
        RECT 16.950 253.950 19.050 256.050 ;
        RECT 20.400 253.050 21.450 256.950 ;
        RECT 19.950 250.950 22.050 253.050 ;
        RECT 26.400 244.050 27.450 259.950 ;
        RECT 7.950 243.450 10.050 244.050 ;
        RECT 7.950 242.400 12.450 243.450 ;
        RECT 7.950 241.950 10.050 242.400 ;
        RECT 1.950 238.950 4.050 241.050 ;
        RECT 4.950 239.250 7.050 240.150 ;
        RECT 7.950 239.850 10.050 240.750 ;
        RECT 2.400 172.050 3.450 238.950 ;
        RECT 4.950 235.950 7.050 238.050 ;
        RECT 11.400 211.050 12.450 242.400 ;
        RECT 13.950 241.950 16.050 244.050 ;
        RECT 19.950 241.950 22.050 244.050 ;
        RECT 25.950 241.950 28.050 244.050 ;
        RECT 13.950 238.950 16.050 241.050 ;
        RECT 17.250 239.250 19.050 240.150 ;
        RECT 19.950 239.850 22.050 240.750 ;
        RECT 22.950 239.250 25.050 240.150 ;
        RECT 26.400 238.050 27.450 241.950 ;
        RECT 13.950 236.850 15.750 237.750 ;
        RECT 16.950 235.950 19.050 238.050 ;
        RECT 19.950 235.950 22.050 238.050 ;
        RECT 22.950 235.950 25.050 238.050 ;
        RECT 25.950 235.950 28.050 238.050 ;
        RECT 17.400 235.050 18.450 235.950 ;
        RECT 16.950 232.950 19.050 235.050 ;
        RECT 7.950 208.950 10.050 211.050 ;
        RECT 10.950 208.950 13.050 211.050 ;
        RECT 8.400 202.050 9.450 208.950 ;
        RECT 20.400 208.050 21.450 235.950 ;
        RECT 29.400 235.050 30.450 265.950 ;
        RECT 32.400 262.050 33.450 271.950 ;
        RECT 34.950 269.850 36.750 270.750 ;
        RECT 37.950 268.950 40.050 271.050 ;
        RECT 41.250 269.850 43.050 270.750 ;
        RECT 38.400 265.050 39.450 268.950 ;
        RECT 40.950 265.950 43.050 268.050 ;
        RECT 37.950 262.950 40.050 265.050 ;
        RECT 31.950 259.950 34.050 262.050 ;
        RECT 41.400 256.050 42.450 265.950 ;
        RECT 37.950 253.950 40.050 256.050 ;
        RECT 40.950 253.950 43.050 256.050 ;
        RECT 31.950 235.950 34.050 238.050 ;
        RECT 35.250 236.250 37.050 237.150 ;
        RECT 25.950 233.850 27.750 234.750 ;
        RECT 28.950 232.950 31.050 235.050 ;
        RECT 32.250 233.850 33.750 234.750 ;
        RECT 34.950 232.950 37.050 235.050 ;
        RECT 38.400 234.450 39.450 253.950 ;
        RECT 40.950 244.950 43.050 247.050 ;
        RECT 41.400 244.050 42.450 244.950 ;
        RECT 44.400 244.050 45.450 272.400 ;
        RECT 47.400 259.050 48.450 281.400 ;
        RECT 56.400 280.050 57.450 337.950 ;
        RECT 59.400 334.050 60.450 344.400 ;
        RECT 62.400 343.050 63.450 349.950 ;
        RECT 65.400 343.050 66.450 379.950 ;
        RECT 68.400 379.050 69.450 379.950 ;
        RECT 67.950 376.950 70.050 379.050 ;
        RECT 71.400 373.050 72.450 445.950 ;
        RECT 74.400 442.050 75.450 451.950 ;
        RECT 79.950 449.850 82.050 450.750 ;
        RECT 79.950 442.950 82.050 445.050 ;
        RECT 73.950 439.950 76.050 442.050 ;
        RECT 80.400 421.050 81.450 442.950 ;
        RECT 83.400 439.050 84.450 463.950 ;
        RECT 86.400 460.050 87.450 463.950 ;
        RECT 88.950 460.950 91.050 463.050 ;
        RECT 85.950 457.950 88.050 460.050 ;
        RECT 89.400 457.050 90.450 460.950 ;
        RECT 88.950 454.950 91.050 457.050 ;
        RECT 85.950 452.250 87.750 453.150 ;
        RECT 88.950 451.950 91.050 454.050 ;
        RECT 92.250 452.250 94.050 453.150 ;
        RECT 89.250 449.850 90.750 450.750 ;
        RECT 91.950 448.950 94.050 451.050 ;
        RECT 92.400 442.050 93.450 448.950 ;
        RECT 91.950 439.950 94.050 442.050 ;
        RECT 82.950 436.950 85.050 439.050 ;
        RECT 85.950 433.950 88.050 436.050 ;
        RECT 82.950 424.950 85.050 427.050 ;
        RECT 83.400 424.050 84.450 424.950 ;
        RECT 82.950 421.950 85.050 424.050 ;
        RECT 79.950 418.950 82.050 421.050 ;
        RECT 83.400 417.450 84.450 421.950 ;
        RECT 86.400 418.050 87.450 433.950 ;
        RECT 95.400 432.450 96.450 469.950 ;
        RECT 98.400 436.050 99.450 472.950 ;
        RECT 101.400 472.050 102.450 502.950 ;
        RECT 104.400 486.450 105.450 517.950 ;
        RECT 107.400 508.050 108.450 520.950 ;
        RECT 106.950 505.950 109.050 508.050 ;
        RECT 110.400 505.050 111.450 532.950 ;
        RECT 113.400 532.050 114.450 541.950 ;
        RECT 112.950 529.950 115.050 532.050 ;
        RECT 113.400 529.050 114.450 529.950 ;
        RECT 119.400 529.050 120.450 544.950 ;
        RECT 124.950 529.950 127.050 532.050 ;
        RECT 125.400 529.050 126.450 529.950 ;
        RECT 112.950 526.950 115.050 529.050 ;
        RECT 116.250 527.250 117.750 528.150 ;
        RECT 118.950 526.950 121.050 529.050 ;
        RECT 122.250 527.250 123.750 528.150 ;
        RECT 124.950 526.950 127.050 529.050 ;
        RECT 112.950 524.850 114.750 525.750 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 119.250 524.850 120.750 525.750 ;
        RECT 121.950 523.950 124.050 526.050 ;
        RECT 125.250 524.850 127.050 525.750 ;
        RECT 112.950 505.950 115.050 508.050 ;
        RECT 109.950 502.950 112.050 505.050 ;
        RECT 106.950 488.250 109.050 489.150 ;
        RECT 113.400 487.050 114.450 505.950 ;
        RECT 116.400 502.050 117.450 523.950 ;
        RECT 122.400 517.050 123.450 523.950 ;
        RECT 121.950 514.950 124.050 517.050 ;
        RECT 115.950 499.950 118.050 502.050 ;
        RECT 122.400 490.050 123.450 514.950 ;
        RECT 128.400 511.050 129.450 586.950 ;
        RECT 131.400 571.050 132.450 589.950 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 131.400 562.050 132.450 568.950 ;
        RECT 142.950 565.950 145.050 568.050 ;
        RECT 136.950 563.250 139.050 564.150 ;
        RECT 130.950 559.950 133.050 562.050 ;
        RECT 134.250 560.250 135.750 561.150 ;
        RECT 136.950 559.950 139.050 562.050 ;
        RECT 140.250 560.250 142.050 561.150 ;
        RECT 143.400 559.050 144.450 565.950 ;
        RECT 146.400 559.050 147.450 592.950 ;
        RECT 155.400 592.050 156.450 595.950 ;
        RECT 164.400 595.050 165.450 625.950 ;
        RECT 160.950 593.850 163.050 594.750 ;
        RECT 163.950 592.950 166.050 595.050 ;
        RECT 154.950 589.950 157.050 592.050 ;
        RECT 167.400 586.050 168.450 629.400 ;
        RECT 169.950 628.950 172.050 631.050 ;
        RECT 173.250 629.850 175.050 630.750 ;
        RECT 170.400 622.050 171.450 628.950 ;
        RECT 179.400 622.050 180.450 632.400 ;
        RECT 181.950 631.950 184.050 632.400 ;
        RECT 185.250 632.250 186.750 633.150 ;
        RECT 187.950 632.400 192.450 633.450 ;
        RECT 187.950 631.950 190.050 632.400 ;
        RECT 181.950 629.850 183.750 630.750 ;
        RECT 184.950 628.950 187.050 631.050 ;
        RECT 188.250 629.850 190.050 630.750 ;
        RECT 191.400 628.050 192.450 632.400 ;
        RECT 193.950 631.950 196.050 634.050 ;
        RECT 197.250 632.250 198.750 633.150 ;
        RECT 199.950 631.950 202.050 634.050 ;
        RECT 203.250 632.250 205.050 633.150 ;
        RECT 208.950 631.950 211.050 634.050 ;
        RECT 212.250 632.250 213.750 633.150 ;
        RECT 214.950 631.950 217.050 634.050 ;
        RECT 217.950 632.250 219.750 633.150 ;
        RECT 220.950 631.950 223.050 634.050 ;
        RECT 226.950 633.450 229.050 634.050 ;
        RECT 224.250 632.250 225.750 633.150 ;
        RECT 226.950 632.400 231.450 633.450 ;
        RECT 226.950 631.950 229.050 632.400 ;
        RECT 193.950 629.850 195.750 630.750 ;
        RECT 196.950 628.950 199.050 631.050 ;
        RECT 200.400 628.050 201.450 631.950 ;
        RECT 202.950 628.950 205.050 631.050 ;
        RECT 208.950 629.850 210.750 630.750 ;
        RECT 211.950 628.950 214.050 631.050 ;
        RECT 215.250 629.850 217.050 630.750 ;
        RECT 217.950 628.950 220.050 631.050 ;
        RECT 184.950 625.950 187.050 628.050 ;
        RECT 190.950 625.950 193.050 628.050 ;
        RECT 199.950 625.950 202.050 628.050 ;
        RECT 169.950 619.950 172.050 622.050 ;
        RECT 178.950 619.950 181.050 622.050 ;
        RECT 181.950 604.950 184.050 607.050 ;
        RECT 172.950 603.450 175.050 604.050 ;
        RECT 172.950 602.400 177.450 603.450 ;
        RECT 172.950 601.950 175.050 602.400 ;
        RECT 169.950 599.250 172.050 600.150 ;
        RECT 172.950 599.850 175.050 600.750 ;
        RECT 169.950 595.950 172.050 598.050 ;
        RECT 166.950 583.950 169.050 586.050 ;
        RECT 176.400 571.050 177.450 602.400 ;
        RECT 182.400 598.050 183.450 604.950 ;
        RECT 185.400 604.050 186.450 625.950 ;
        RECT 199.950 616.950 202.050 619.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 190.950 603.450 193.050 604.050 ;
        RECT 188.400 602.400 193.050 603.450 ;
        RECT 178.950 596.250 180.750 597.150 ;
        RECT 181.950 595.950 184.050 598.050 ;
        RECT 185.400 595.050 186.450 601.950 ;
        RECT 188.400 598.050 189.450 602.400 ;
        RECT 190.950 601.950 193.050 602.400 ;
        RECT 190.950 599.850 193.050 600.750 ;
        RECT 193.950 599.250 196.050 600.150 ;
        RECT 200.400 598.050 201.450 616.950 ;
        RECT 203.400 616.050 204.450 628.950 ;
        RECT 208.950 625.950 211.050 628.050 ;
        RECT 202.950 613.950 205.050 616.050 ;
        RECT 205.950 604.950 208.050 607.050 ;
        RECT 202.950 601.950 205.050 604.050 ;
        RECT 187.950 597.450 190.050 598.050 ;
        RECT 187.950 596.400 192.450 597.450 ;
        RECT 187.950 595.950 190.050 596.400 ;
        RECT 178.950 592.950 181.050 595.050 ;
        RECT 182.250 593.850 183.750 594.750 ;
        RECT 184.950 592.950 187.050 595.050 ;
        RECT 188.250 593.850 190.050 594.750 ;
        RECT 184.950 590.850 187.050 591.750 ;
        RECT 191.400 586.050 192.450 596.400 ;
        RECT 193.950 595.950 196.050 598.050 ;
        RECT 199.950 595.950 202.050 598.050 ;
        RECT 203.400 595.050 204.450 601.950 ;
        RECT 206.400 598.050 207.450 604.950 ;
        RECT 209.400 601.050 210.450 625.950 ;
        RECT 212.400 619.050 213.450 628.950 ;
        RECT 217.950 619.950 220.050 622.050 ;
        RECT 211.950 616.950 214.050 619.050 ;
        RECT 211.950 613.950 214.050 616.050 ;
        RECT 208.950 598.950 211.050 601.050 ;
        RECT 205.950 595.950 208.050 598.050 ;
        RECT 209.250 596.250 211.050 597.150 ;
        RECT 199.950 593.850 201.750 594.750 ;
        RECT 202.950 592.950 205.050 595.050 ;
        RECT 206.250 593.850 207.750 594.750 ;
        RECT 208.950 592.950 211.050 595.050 ;
        RECT 212.400 592.050 213.450 613.950 ;
        RECT 214.950 601.950 217.050 604.050 ;
        RECT 215.400 598.050 216.450 601.950 ;
        RECT 214.950 595.950 217.050 598.050 ;
        RECT 218.400 595.050 219.450 619.950 ;
        RECT 221.400 604.050 222.450 631.950 ;
        RECT 223.950 628.950 226.050 631.050 ;
        RECT 227.250 629.850 229.050 630.750 ;
        RECT 224.400 625.050 225.450 628.950 ;
        RECT 223.950 622.950 226.050 625.050 ;
        RECT 230.400 613.050 231.450 632.400 ;
        RECT 233.400 631.050 234.450 634.950 ;
        RECT 257.400 633.450 258.450 671.400 ;
        RECT 259.950 670.950 262.050 671.400 ;
        RECT 263.250 671.250 265.050 672.150 ;
        RECT 265.950 671.850 268.050 672.750 ;
        RECT 268.950 671.250 271.050 672.150 ;
        RECT 271.950 671.850 274.050 672.750 ;
        RECT 274.950 671.250 277.050 672.150 ;
        RECT 283.950 671.250 286.050 672.150 ;
        RECT 286.950 671.850 289.050 672.750 ;
        RECT 289.950 671.250 292.050 672.150 ;
        RECT 292.950 671.850 295.050 672.750 ;
        RECT 295.950 671.250 297.750 672.150 ;
        RECT 298.950 670.950 301.050 673.050 ;
        RECT 302.400 672.450 303.450 676.950 ;
        RECT 308.400 676.050 309.450 676.950 ;
        RECT 307.950 673.950 310.050 676.050 ;
        RECT 316.950 675.450 319.050 676.050 ;
        RECT 314.400 674.400 319.050 675.450 ;
        RECT 304.950 672.450 307.050 673.050 ;
        RECT 302.400 671.400 307.050 672.450 ;
        RECT 308.250 671.850 309.750 672.750 ;
        RECT 310.950 672.450 313.050 673.050 ;
        RECT 314.400 672.450 315.450 674.400 ;
        RECT 316.950 673.950 319.050 674.400 ;
        RECT 325.950 673.950 328.050 676.050 ;
        RECT 326.400 673.050 327.450 673.950 ;
        RECT 302.400 670.050 303.450 671.400 ;
        RECT 304.950 670.950 307.050 671.400 ;
        RECT 310.950 671.400 315.450 672.450 ;
        RECT 316.950 671.850 319.050 672.750 ;
        RECT 310.950 670.950 313.050 671.400 ;
        RECT 259.950 668.850 261.750 669.750 ;
        RECT 262.950 667.950 265.050 670.050 ;
        RECT 268.950 667.950 271.050 670.050 ;
        RECT 274.950 667.950 277.050 670.050 ;
        RECT 283.950 667.950 286.050 670.050 ;
        RECT 289.950 667.950 292.050 670.050 ;
        RECT 295.950 667.950 298.050 670.050 ;
        RECT 299.250 668.850 301.050 669.750 ;
        RECT 301.950 667.950 304.050 670.050 ;
        RECT 304.950 668.850 307.050 669.750 ;
        RECT 310.950 668.850 313.050 669.750 ;
        RECT 263.400 661.050 264.450 667.950 ;
        RECT 262.950 658.950 265.050 661.050 ;
        RECT 269.400 649.050 270.450 667.950 ;
        RECT 275.400 667.050 276.450 667.950 ;
        RECT 274.950 664.950 277.050 667.050 ;
        RECT 290.400 649.050 291.450 667.950 ;
        RECT 296.400 667.050 297.450 667.950 ;
        RECT 295.950 664.950 298.050 667.050 ;
        RECT 304.950 658.950 307.050 661.050 ;
        RECT 268.950 646.950 271.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 268.950 634.950 271.050 637.050 ;
        RECT 257.400 632.400 261.450 633.450 ;
        RECT 260.400 631.050 261.450 632.400 ;
        RECT 265.950 632.250 268.050 633.150 ;
        RECT 232.950 628.950 235.050 631.050 ;
        RECT 235.950 629.250 238.050 630.150 ;
        RECT 241.950 629.250 244.050 630.150 ;
        RECT 247.950 629.250 250.050 630.150 ;
        RECT 253.950 629.250 256.050 630.150 ;
        RECT 256.950 629.250 258.750 630.150 ;
        RECT 259.950 628.950 262.050 631.050 ;
        RECT 265.950 630.450 268.050 631.050 ;
        RECT 269.400 630.450 270.450 634.950 ;
        RECT 274.950 631.950 277.050 634.050 ;
        RECT 278.250 632.250 279.750 633.150 ;
        RECT 280.950 631.950 283.050 634.050 ;
        RECT 284.400 631.050 285.450 646.950 ;
        RECT 289.950 634.950 292.050 637.050 ;
        RECT 295.950 635.250 298.050 636.150 ;
        RECT 286.950 631.950 289.050 634.050 ;
        RECT 287.400 631.050 288.450 631.950 ;
        RECT 263.250 629.250 264.750 630.150 ;
        RECT 265.950 629.400 270.450 630.450 ;
        RECT 265.950 628.950 268.050 629.400 ;
        RECT 271.950 628.950 274.050 631.050 ;
        RECT 274.950 629.850 276.750 630.750 ;
        RECT 277.950 628.950 280.050 631.050 ;
        RECT 281.250 629.850 283.050 630.750 ;
        RECT 283.950 628.950 286.050 631.050 ;
        RECT 286.950 628.950 289.050 631.050 ;
        RECT 290.400 630.450 291.450 634.950 ;
        RECT 292.950 632.250 294.750 633.150 ;
        RECT 295.950 631.950 298.050 634.050 ;
        RECT 299.250 632.250 300.750 633.150 ;
        RECT 301.950 631.950 304.050 634.050 ;
        RECT 292.950 630.450 295.050 631.050 ;
        RECT 290.400 629.400 295.050 630.450 ;
        RECT 292.950 628.950 295.050 629.400 ;
        RECT 298.950 628.950 301.050 631.050 ;
        RECT 302.250 629.850 304.050 630.750 ;
        RECT 233.400 627.450 234.450 628.950 ;
        RECT 235.950 627.450 238.050 628.050 ;
        RECT 233.400 626.400 238.050 627.450 ;
        RECT 235.950 625.950 238.050 626.400 ;
        RECT 239.250 626.250 240.750 627.150 ;
        RECT 241.950 625.950 244.050 628.050 ;
        RECT 247.950 625.950 250.050 628.050 ;
        RECT 251.250 626.250 252.750 627.150 ;
        RECT 253.950 625.950 256.050 628.050 ;
        RECT 256.950 625.950 259.050 628.050 ;
        RECT 260.250 626.850 261.750 627.750 ;
        RECT 262.950 625.950 265.050 628.050 ;
        RECT 238.950 622.950 241.050 625.050 ;
        RECT 229.950 610.950 232.050 613.050 ;
        RECT 220.950 601.950 223.050 604.050 ;
        RECT 224.400 602.400 234.450 603.450 ;
        RECT 224.400 600.450 225.450 602.400 ;
        RECT 221.400 599.400 225.450 600.450 ;
        RECT 221.400 598.050 222.450 599.400 ;
        RECT 226.950 598.950 229.050 601.050 ;
        RECT 220.950 595.950 223.050 598.050 ;
        RECT 224.250 596.250 226.050 597.150 ;
        RECT 214.950 593.850 216.750 594.750 ;
        RECT 217.950 592.950 220.050 595.050 ;
        RECT 221.250 593.850 222.750 594.750 ;
        RECT 223.950 592.950 226.050 595.050 ;
        RECT 202.950 590.850 205.050 591.750 ;
        RECT 211.950 589.950 214.050 592.050 ;
        RECT 217.950 590.850 220.050 591.750 ;
        RECT 220.950 589.950 223.050 592.050 ;
        RECT 184.950 583.950 187.050 586.050 ;
        RECT 190.950 583.950 193.050 586.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 175.950 568.950 178.050 571.050 ;
        RECT 148.950 562.950 151.050 565.050 ;
        RECT 149.400 559.050 150.450 562.950 ;
        RECT 155.400 562.050 156.450 568.950 ;
        RECT 160.950 563.250 163.050 564.150 ;
        RECT 154.950 559.950 157.050 562.050 ;
        RECT 157.950 560.250 159.750 561.150 ;
        RECT 160.950 559.950 163.050 562.050 ;
        RECT 164.250 560.250 165.750 561.150 ;
        RECT 166.950 559.950 169.050 562.050 ;
        RECT 130.950 557.850 132.750 558.750 ;
        RECT 133.950 558.450 136.050 559.050 ;
        RECT 133.950 557.400 138.450 558.450 ;
        RECT 133.950 556.950 136.050 557.400 ;
        RECT 137.400 553.050 138.450 557.400 ;
        RECT 139.950 556.950 142.050 559.050 ;
        RECT 142.950 556.950 145.050 559.050 ;
        RECT 145.950 556.950 148.050 559.050 ;
        RECT 148.950 556.950 151.050 559.050 ;
        RECT 152.250 557.250 154.050 558.150 ;
        RECT 157.950 556.950 160.050 559.050 ;
        RECT 140.400 556.050 141.450 556.950 ;
        RECT 158.400 556.050 159.450 556.950 ;
        RECT 139.950 553.950 142.050 556.050 ;
        RECT 142.950 554.850 145.050 555.750 ;
        RECT 145.950 554.250 148.050 555.150 ;
        RECT 148.950 554.850 150.750 555.750 ;
        RECT 151.950 553.950 154.050 556.050 ;
        RECT 157.950 553.950 160.050 556.050 ;
        RECT 140.400 553.050 141.450 553.950 ;
        RECT 161.400 553.050 162.450 559.950 ;
        RECT 163.950 556.950 166.050 559.050 ;
        RECT 167.250 557.850 169.050 558.750 ;
        RECT 172.950 558.450 175.050 559.050 ;
        RECT 170.400 557.400 175.050 558.450 ;
        RECT 136.950 550.950 139.050 553.050 ;
        RECT 139.950 550.950 142.050 553.050 ;
        RECT 145.950 550.950 148.050 553.050 ;
        RECT 160.950 550.950 163.050 553.050 ;
        RECT 130.950 529.950 133.050 532.050 ;
        RECT 130.950 527.850 133.050 528.750 ;
        RECT 133.950 527.250 136.050 528.150 ;
        RECT 130.950 523.950 133.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 127.950 508.950 130.050 511.050 ;
        RECT 131.400 490.050 132.450 523.950 ;
        RECT 137.400 505.050 138.450 550.950 ;
        RECT 139.950 547.950 142.050 550.050 ;
        RECT 140.400 522.450 141.450 547.950 ;
        RECT 146.400 535.050 147.450 550.950 ;
        RECT 160.950 544.950 163.050 547.050 ;
        RECT 161.400 541.050 162.450 544.950 ;
        RECT 164.400 541.050 165.450 556.950 ;
        RECT 170.400 556.050 171.450 557.400 ;
        RECT 172.950 556.950 175.050 557.400 ;
        RECT 178.950 556.950 181.050 559.050 ;
        RECT 182.250 557.250 184.050 558.150 ;
        RECT 169.950 553.950 172.050 556.050 ;
        RECT 172.950 554.850 175.050 555.750 ;
        RECT 175.950 554.250 178.050 555.150 ;
        RECT 178.950 554.850 180.750 555.750 ;
        RECT 181.950 553.950 184.050 556.050 ;
        RECT 182.400 553.050 183.450 553.950 ;
        RECT 175.950 550.950 178.050 553.050 ;
        RECT 181.950 550.950 184.050 553.050 ;
        RECT 169.950 541.950 172.050 544.050 ;
        RECT 160.950 538.950 163.050 541.050 ;
        RECT 163.950 538.950 166.050 541.050 ;
        RECT 148.950 535.950 151.050 538.050 ;
        RECT 166.950 535.950 169.050 538.050 ;
        RECT 142.950 532.950 145.050 535.050 ;
        RECT 145.950 532.950 148.050 535.050 ;
        RECT 143.400 528.450 144.450 532.950 ;
        RECT 149.400 529.050 150.450 535.950 ;
        RECT 151.950 529.950 154.050 532.050 ;
        RECT 157.950 529.950 160.050 532.050 ;
        RECT 163.950 529.950 166.050 532.050 ;
        RECT 143.400 527.400 147.450 528.450 ;
        RECT 146.400 526.050 147.450 527.400 ;
        RECT 148.950 526.950 151.050 529.050 ;
        RECT 152.400 526.050 153.450 529.950 ;
        RECT 164.400 529.050 165.450 529.950 ;
        RECT 154.950 527.250 157.050 528.150 ;
        RECT 157.950 527.850 160.050 528.750 ;
        RECT 160.950 527.250 162.750 528.150 ;
        RECT 163.950 526.950 166.050 529.050 ;
        RECT 167.400 526.050 168.450 535.950 ;
        RECT 170.400 529.050 171.450 541.950 ;
        RECT 172.950 535.950 175.050 538.050 ;
        RECT 173.400 532.050 174.450 535.950 ;
        RECT 185.400 532.050 186.450 583.950 ;
        RECT 199.950 577.950 202.050 580.050 ;
        RECT 200.400 562.050 201.450 577.950 ;
        RECT 205.950 563.250 208.050 564.150 ;
        RECT 211.950 562.950 214.050 565.050 ;
        RECT 199.950 559.950 202.050 562.050 ;
        RECT 203.250 560.250 204.750 561.150 ;
        RECT 205.950 559.950 208.050 562.050 ;
        RECT 209.250 560.250 211.050 561.150 ;
        RECT 190.950 556.950 193.050 559.050 ;
        RECT 199.950 557.850 201.750 558.750 ;
        RECT 202.950 556.950 205.050 559.050 ;
        RECT 208.950 556.950 211.050 559.050 ;
        RECT 187.950 554.250 190.050 555.150 ;
        RECT 190.950 554.850 193.050 555.750 ;
        RECT 209.400 553.050 210.450 556.950 ;
        RECT 212.400 553.050 213.450 562.950 ;
        RECT 214.950 556.950 217.050 559.050 ;
        RECT 221.400 556.050 222.450 589.950 ;
        RECT 227.400 580.050 228.450 598.950 ;
        RECT 233.400 598.050 234.450 602.400 ;
        RECT 239.400 601.050 240.450 622.950 ;
        RECT 242.400 616.050 243.450 625.950 ;
        RECT 248.400 616.050 249.450 625.950 ;
        RECT 250.950 622.950 253.050 625.050 ;
        RECT 241.950 613.950 244.050 616.050 ;
        RECT 247.950 613.950 250.050 616.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 254.400 601.050 255.450 625.950 ;
        RECT 257.400 619.050 258.450 625.950 ;
        RECT 256.950 616.950 259.050 619.050 ;
        RECT 256.950 613.950 259.050 616.050 ;
        RECT 257.400 601.050 258.450 613.950 ;
        RECT 272.400 610.050 273.450 628.950 ;
        RECT 278.400 622.050 279.450 628.950 ;
        RECT 283.950 626.250 286.050 627.150 ;
        RECT 286.950 626.850 289.050 627.750 ;
        RECT 289.950 625.950 292.050 628.050 ;
        RECT 283.950 622.950 286.050 625.050 ;
        RECT 277.950 619.950 280.050 622.050 ;
        RECT 280.950 610.950 283.050 613.050 ;
        RECT 271.950 607.950 274.050 610.050 ;
        RECT 268.950 604.950 271.050 607.050 ;
        RECT 238.950 598.950 241.050 601.050 ;
        RECT 244.950 598.950 247.050 601.050 ;
        RECT 248.250 599.850 249.750 600.750 ;
        RECT 250.950 598.950 253.050 601.050 ;
        RECT 253.950 598.950 256.050 601.050 ;
        RECT 256.950 598.950 259.050 601.050 ;
        RECT 262.950 598.950 265.050 601.050 ;
        RECT 265.950 598.950 268.050 601.050 ;
        RECT 229.950 596.250 231.750 597.150 ;
        RECT 232.950 595.950 235.050 598.050 ;
        RECT 236.250 596.250 238.050 597.150 ;
        RECT 244.950 596.850 247.050 597.750 ;
        RECT 250.950 596.850 253.050 597.750 ;
        RECT 256.950 596.850 259.050 597.750 ;
        RECT 259.950 596.250 262.050 597.150 ;
        RECT 229.950 592.950 232.050 595.050 ;
        RECT 233.250 593.850 234.750 594.750 ;
        RECT 235.950 592.950 238.050 595.050 ;
        RECT 259.950 594.450 262.050 595.050 ;
        RECT 257.400 593.400 262.050 594.450 ;
        RECT 230.400 592.050 231.450 592.950 ;
        RECT 229.950 589.950 232.050 592.050 ;
        RECT 236.400 580.050 237.450 592.950 ;
        RECT 226.950 577.950 229.050 580.050 ;
        RECT 235.950 577.950 238.050 580.050 ;
        RECT 244.950 562.950 247.050 565.050 ;
        RECT 223.950 560.250 226.050 561.150 ;
        RECT 235.950 559.950 238.050 562.050 ;
        RECT 223.950 556.950 226.050 559.050 ;
        RECT 227.250 557.250 228.750 558.150 ;
        RECT 229.950 556.950 232.050 559.050 ;
        RECT 233.250 557.250 235.050 558.150 ;
        RECT 214.950 554.850 217.050 555.750 ;
        RECT 217.950 554.250 220.050 555.150 ;
        RECT 220.950 553.950 223.050 556.050 ;
        RECT 226.950 553.950 229.050 556.050 ;
        RECT 230.250 554.850 231.750 555.750 ;
        RECT 232.950 553.950 235.050 556.050 ;
        RECT 187.950 550.950 190.050 553.050 ;
        RECT 208.950 550.950 211.050 553.050 ;
        RECT 211.950 550.950 214.050 553.050 ;
        RECT 217.950 550.950 220.050 553.050 ;
        RECT 188.400 550.050 189.450 550.950 ;
        RECT 187.950 547.950 190.050 550.050 ;
        RECT 205.950 544.950 208.050 547.050 ;
        RECT 190.950 532.950 193.050 535.050 ;
        RECT 172.950 529.950 175.050 532.050 ;
        RECT 184.950 529.950 187.050 532.050 ;
        RECT 169.950 526.950 172.050 529.050 ;
        RECT 173.250 527.850 174.750 528.750 ;
        RECT 175.950 528.450 178.050 529.050 ;
        RECT 175.950 527.400 180.450 528.450 ;
        RECT 175.950 526.950 178.050 527.400 ;
        RECT 142.950 524.250 144.750 525.150 ;
        RECT 145.950 523.950 148.050 526.050 ;
        RECT 151.950 523.950 154.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 164.250 524.850 166.050 525.750 ;
        RECT 166.950 523.950 169.050 526.050 ;
        RECT 169.950 524.850 172.050 525.750 ;
        RECT 172.950 523.950 175.050 526.050 ;
        RECT 175.950 524.850 178.050 525.750 ;
        RECT 155.400 523.050 156.450 523.950 ;
        RECT 142.950 522.450 145.050 523.050 ;
        RECT 140.400 521.400 145.050 522.450 ;
        RECT 146.250 521.850 147.750 522.750 ;
        RECT 142.950 520.950 145.050 521.400 ;
        RECT 148.950 520.950 151.050 523.050 ;
        RECT 152.250 521.850 154.050 522.750 ;
        RECT 154.950 520.950 157.050 523.050 ;
        RECT 139.950 517.950 142.050 520.050 ;
        RECT 148.950 518.850 151.050 519.750 ;
        RECT 140.400 511.050 141.450 517.950 ;
        RECT 161.400 517.050 162.450 523.950 ;
        RECT 163.950 520.950 166.050 523.050 ;
        RECT 160.950 514.950 163.050 517.050 ;
        RECT 139.950 508.950 142.050 511.050 ;
        RECT 151.950 508.950 154.050 511.050 ;
        RECT 136.950 502.950 139.050 505.050 ;
        RECT 145.950 502.950 148.050 505.050 ;
        RECT 136.950 490.950 139.050 493.050 ;
        RECT 137.400 490.050 138.450 490.950 ;
        RECT 121.950 487.950 124.050 490.050 ;
        RECT 130.950 487.950 133.050 490.050 ;
        RECT 136.950 487.950 139.050 490.050 ;
        RECT 140.250 488.250 141.750 489.150 ;
        RECT 106.950 486.450 109.050 487.050 ;
        RECT 104.400 485.400 109.050 486.450 ;
        RECT 106.950 484.950 109.050 485.400 ;
        RECT 110.250 485.250 111.750 486.150 ;
        RECT 112.950 484.950 115.050 487.050 ;
        RECT 116.250 485.250 118.050 486.150 ;
        RECT 121.950 485.250 123.750 486.150 ;
        RECT 128.250 485.250 129.750 486.150 ;
        RECT 134.250 485.250 136.050 486.150 ;
        RECT 136.950 485.850 138.750 486.750 ;
        RECT 139.950 484.950 142.050 487.050 ;
        RECT 143.250 485.850 145.050 486.750 ;
        RECT 109.950 481.950 112.050 484.050 ;
        RECT 113.250 482.850 114.750 483.750 ;
        RECT 115.950 481.950 118.050 484.050 ;
        RECT 121.950 481.950 124.050 484.050 ;
        RECT 125.250 482.850 126.750 483.750 ;
        RECT 127.950 481.950 130.050 484.050 ;
        RECT 131.250 482.850 132.750 483.750 ;
        RECT 133.950 481.950 136.050 484.050 ;
        RECT 116.400 480.450 117.450 481.950 ;
        RECT 122.400 481.050 123.450 481.950 ;
        RECT 113.400 479.400 117.450 480.450 ;
        RECT 113.400 475.050 114.450 479.400 ;
        RECT 121.950 478.950 124.050 481.050 ;
        RECT 124.950 478.950 127.050 481.050 ;
        RECT 115.950 475.950 118.050 478.050 ;
        RECT 112.950 472.950 115.050 475.050 ;
        RECT 100.950 469.950 103.050 472.050 ;
        RECT 116.400 460.050 117.450 475.950 ;
        RECT 118.950 463.950 121.050 466.050 ;
        RECT 115.950 457.950 118.050 460.050 ;
        RECT 119.400 457.050 120.450 463.950 ;
        RECT 125.400 462.450 126.450 478.950 ;
        RECT 130.950 475.950 133.050 478.050 ;
        RECT 131.400 475.050 132.450 475.950 ;
        RECT 130.950 472.950 133.050 475.050 ;
        RECT 125.400 461.400 129.450 462.450 ;
        RECT 124.950 457.950 127.050 460.050 ;
        RECT 125.400 457.050 126.450 457.950 ;
        RECT 128.400 457.050 129.450 461.400 ;
        RECT 112.950 454.950 115.050 457.050 ;
        RECT 116.250 455.850 117.750 456.750 ;
        RECT 118.950 454.950 121.050 457.050 ;
        RECT 124.950 454.950 127.050 457.050 ;
        RECT 127.950 454.950 130.050 457.050 ;
        RECT 125.400 454.050 126.450 454.950 ;
        RECT 100.950 452.250 102.750 453.150 ;
        RECT 103.950 451.950 106.050 454.050 ;
        RECT 107.250 452.250 109.050 453.150 ;
        RECT 112.950 452.850 115.050 453.750 ;
        RECT 118.950 452.850 121.050 453.750 ;
        RECT 121.950 452.250 123.750 453.150 ;
        RECT 124.950 451.950 127.050 454.050 ;
        RECT 128.250 452.250 130.050 453.150 ;
        RECT 104.250 449.850 105.750 450.750 ;
        RECT 106.950 448.950 109.050 451.050 ;
        RECT 121.950 448.950 124.050 451.050 ;
        RECT 125.250 449.850 126.750 450.750 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 115.950 445.950 118.050 448.050 ;
        RECT 97.950 433.950 100.050 436.050 ;
        RECT 95.400 431.400 99.450 432.450 ;
        RECT 73.950 416.250 76.050 417.150 ;
        RECT 80.400 416.400 84.450 417.450 ;
        RECT 80.400 415.050 81.450 416.400 ;
        RECT 85.950 415.950 88.050 418.050 ;
        RECT 89.250 416.250 90.750 417.150 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 77.250 413.250 78.750 414.150 ;
        RECT 79.950 412.950 82.050 415.050 ;
        RECT 83.250 413.250 85.050 414.150 ;
        RECT 85.950 413.850 87.750 414.750 ;
        RECT 88.950 412.950 91.050 415.050 ;
        RECT 92.250 413.850 94.050 414.750 ;
        RECT 74.400 412.050 75.450 412.950 ;
        RECT 73.950 409.950 76.050 412.050 ;
        RECT 76.950 409.950 79.050 412.050 ;
        RECT 80.250 410.850 81.750 411.750 ;
        RECT 82.950 409.950 85.050 412.050 ;
        RECT 85.950 409.950 88.050 412.050 ;
        RECT 73.950 390.450 76.050 391.050 ;
        RECT 77.400 390.450 78.450 409.950 ;
        RECT 79.950 406.950 82.050 409.050 ;
        RECT 73.950 389.400 78.450 390.450 ;
        RECT 73.950 388.950 76.050 389.400 ;
        RECT 76.950 385.950 79.050 388.050 ;
        RECT 77.400 382.050 78.450 385.950 ;
        RECT 80.400 385.050 81.450 406.950 ;
        RECT 82.950 388.950 85.050 391.050 ;
        RECT 79.950 382.950 82.050 385.050 ;
        RECT 80.400 382.050 81.450 382.950 ;
        RECT 83.400 382.050 84.450 388.950 ;
        RECT 73.950 380.250 75.750 381.150 ;
        RECT 76.950 379.950 79.050 382.050 ;
        RECT 79.950 379.950 82.050 382.050 ;
        RECT 82.950 379.950 85.050 382.050 ;
        RECT 73.950 376.950 76.050 379.050 ;
        RECT 77.250 377.850 78.750 378.750 ;
        RECT 79.950 376.950 82.050 379.050 ;
        RECT 83.250 377.850 85.050 378.750 ;
        RECT 70.950 370.950 73.050 373.050 ;
        RECT 74.400 364.050 75.450 376.950 ;
        RECT 86.400 376.050 87.450 409.950 ;
        RECT 89.400 391.050 90.450 412.950 ;
        RECT 91.950 409.950 94.050 412.050 ;
        RECT 92.400 406.050 93.450 409.950 ;
        RECT 98.400 406.050 99.450 431.400 ;
        RECT 101.400 424.050 102.450 445.950 ;
        RECT 103.950 442.950 106.050 445.050 ;
        RECT 106.950 442.950 109.050 445.050 ;
        RECT 100.950 421.950 103.050 424.050 ;
        RECT 104.400 415.050 105.450 442.950 ;
        RECT 107.400 421.050 108.450 442.950 ;
        RECT 112.950 439.950 115.050 442.050 ;
        RECT 113.400 421.050 114.450 439.950 ;
        RECT 106.950 418.950 109.050 421.050 ;
        RECT 112.950 418.950 115.050 421.050 ;
        RECT 116.400 418.050 117.450 445.950 ;
        RECT 131.400 445.050 132.450 472.950 ;
        RECT 134.400 448.050 135.450 481.950 ;
        RECT 146.400 475.050 147.450 502.950 ;
        RECT 148.950 490.950 151.050 493.050 ;
        RECT 149.400 487.050 150.450 490.950 ;
        RECT 152.400 490.050 153.450 508.950 ;
        RECT 164.400 508.050 165.450 520.950 ;
        RECT 163.950 505.950 166.050 508.050 ;
        RECT 164.400 502.050 165.450 505.950 ;
        RECT 163.950 499.950 166.050 502.050 ;
        RECT 157.950 491.250 160.050 492.150 ;
        RECT 151.950 487.950 154.050 490.050 ;
        RECT 155.250 488.250 156.750 489.150 ;
        RECT 161.250 488.250 163.050 489.150 ;
        RECT 148.950 484.950 151.050 487.050 ;
        RECT 151.950 485.850 153.750 486.750 ;
        RECT 154.950 486.450 157.050 487.050 ;
        RECT 154.950 485.400 159.450 486.450 ;
        RECT 154.950 484.950 157.050 485.400 ;
        RECT 158.400 483.450 159.450 485.400 ;
        RECT 160.950 484.950 163.050 487.050 ;
        RECT 160.950 483.450 163.050 484.050 ;
        RECT 158.400 482.400 163.050 483.450 ;
        RECT 160.950 481.950 163.050 482.400 ;
        RECT 139.950 472.950 142.050 475.050 ;
        RECT 145.950 472.950 148.050 475.050 ;
        RECT 136.950 466.950 139.050 469.050 ;
        RECT 137.400 454.050 138.450 466.950 ;
        RECT 140.400 457.050 141.450 472.950 ;
        RECT 148.950 463.950 151.050 466.050 ;
        RECT 160.950 463.950 163.050 466.050 ;
        RECT 139.950 454.950 142.050 457.050 ;
        RECT 143.250 455.250 144.750 456.150 ;
        RECT 145.950 454.950 148.050 457.050 ;
        RECT 136.950 451.950 139.050 454.050 ;
        RECT 140.250 452.850 141.750 453.750 ;
        RECT 142.950 451.950 145.050 454.050 ;
        RECT 146.250 452.850 148.050 453.750 ;
        RECT 136.950 449.850 139.050 450.750 ;
        RECT 139.950 448.950 142.050 451.050 ;
        RECT 133.950 445.950 136.050 448.050 ;
        RECT 130.950 442.950 133.050 445.050 ;
        RECT 130.950 433.950 133.050 436.050 ;
        RECT 124.950 421.950 127.050 424.050 ;
        RECT 115.950 417.450 118.050 418.050 ;
        RECT 113.400 416.400 118.050 417.450 ;
        RECT 113.400 415.050 114.450 416.400 ;
        RECT 115.950 415.950 118.050 416.400 ;
        RECT 119.250 416.250 120.750 417.150 ;
        RECT 125.400 415.050 126.450 421.950 ;
        RECT 100.950 413.250 102.750 414.150 ;
        RECT 103.950 412.950 106.050 415.050 ;
        RECT 109.950 413.250 111.750 414.150 ;
        RECT 112.950 412.950 115.050 415.050 ;
        RECT 115.950 413.850 117.750 414.750 ;
        RECT 118.950 412.950 121.050 415.050 ;
        RECT 122.250 413.850 124.050 414.750 ;
        RECT 124.950 412.950 127.050 415.050 ;
        RECT 127.950 413.250 130.050 414.150 ;
        RECT 100.950 409.950 103.050 412.050 ;
        RECT 104.250 410.850 106.050 411.750 ;
        RECT 109.950 409.950 112.050 412.050 ;
        RECT 113.250 410.850 115.050 411.750 ;
        RECT 91.950 403.950 94.050 406.050 ;
        RECT 97.950 403.950 100.050 406.050 ;
        RECT 101.400 402.450 102.450 409.950 ;
        RECT 115.950 403.950 118.050 406.050 ;
        RECT 98.400 401.400 102.450 402.450 ;
        RECT 91.950 391.950 94.050 394.050 ;
        RECT 88.950 388.950 91.050 391.050 ;
        RECT 92.400 388.050 93.450 391.950 ;
        RECT 91.950 385.950 94.050 388.050 ;
        RECT 92.400 385.050 93.450 385.950 ;
        RECT 98.400 385.050 99.450 401.400 ;
        RECT 88.950 382.950 91.050 385.050 ;
        RECT 91.950 382.950 94.050 385.050 ;
        RECT 95.250 383.250 96.750 384.150 ;
        RECT 97.950 382.950 100.050 385.050 ;
        RECT 103.950 384.450 106.050 385.050 ;
        RECT 101.400 383.400 106.050 384.450 ;
        RECT 89.400 382.050 90.450 382.950 ;
        RECT 88.950 379.950 91.050 382.050 ;
        RECT 92.250 380.850 93.750 381.750 ;
        RECT 94.950 379.950 97.050 382.050 ;
        RECT 98.250 380.850 100.050 381.750 ;
        RECT 88.950 377.850 91.050 378.750 ;
        RECT 91.950 376.950 94.050 379.050 ;
        RECT 79.950 374.850 82.050 375.750 ;
        RECT 85.950 373.950 88.050 376.050 ;
        RECT 86.400 364.050 87.450 373.950 ;
        RECT 88.950 370.950 91.050 373.050 ;
        RECT 73.950 361.950 76.050 364.050 ;
        RECT 85.950 361.950 88.050 364.050 ;
        RECT 67.950 352.950 70.050 355.050 ;
        RECT 68.400 343.050 69.450 352.950 ;
        RECT 76.950 346.950 79.050 349.050 ;
        RECT 77.400 345.450 78.450 346.950 ;
        RECT 74.400 344.400 78.450 345.450 ;
        RECT 61.950 340.950 64.050 343.050 ;
        RECT 64.950 340.950 67.050 343.050 ;
        RECT 67.950 340.950 70.050 343.050 ;
        RECT 71.250 341.250 73.050 342.150 ;
        RECT 61.950 338.850 64.050 339.750 ;
        RECT 64.950 338.250 67.050 339.150 ;
        RECT 67.950 338.850 69.750 339.750 ;
        RECT 70.950 337.950 73.050 340.050 ;
        RECT 64.950 334.950 67.050 337.050 ;
        RECT 70.950 334.950 73.050 337.050 ;
        RECT 58.950 331.950 61.050 334.050 ;
        RECT 59.400 315.450 60.450 331.950 ;
        RECT 67.950 316.950 70.050 319.050 ;
        RECT 61.950 315.450 64.050 316.050 ;
        RECT 59.400 314.400 64.050 315.450 ;
        RECT 61.950 313.950 64.050 314.400 ;
        RECT 68.400 313.050 69.450 316.950 ;
        RECT 71.400 316.050 72.450 334.950 ;
        RECT 70.950 313.950 73.050 316.050 ;
        RECT 58.950 311.250 61.050 312.150 ;
        RECT 61.950 311.850 64.050 312.750 ;
        RECT 64.950 311.250 66.750 312.150 ;
        RECT 67.950 310.950 70.050 313.050 ;
        RECT 74.400 312.450 75.450 344.400 ;
        RECT 85.950 344.250 88.050 345.150 ;
        RECT 76.950 341.250 78.750 342.150 ;
        RECT 79.950 340.950 82.050 343.050 ;
        RECT 83.250 341.250 84.750 342.150 ;
        RECT 85.950 340.950 88.050 343.050 ;
        RECT 76.950 337.950 79.050 340.050 ;
        RECT 80.250 338.850 81.750 339.750 ;
        RECT 82.950 337.950 85.050 340.050 ;
        RECT 77.400 336.450 78.450 337.950 ;
        RECT 77.400 335.400 81.450 336.450 ;
        RECT 76.950 331.950 79.050 334.050 ;
        RECT 71.400 311.400 75.450 312.450 ;
        RECT 58.950 307.950 61.050 310.050 ;
        RECT 61.950 307.950 64.050 310.050 ;
        RECT 64.950 307.950 67.050 310.050 ;
        RECT 68.250 308.850 70.050 309.750 ;
        RECT 58.950 304.950 61.050 307.050 ;
        RECT 59.400 283.050 60.450 304.950 ;
        RECT 58.950 280.950 61.050 283.050 ;
        RECT 55.950 277.950 58.050 280.050 ;
        RECT 62.400 277.050 63.450 307.950 ;
        RECT 65.400 307.050 66.450 307.950 ;
        RECT 64.950 304.950 67.050 307.050 ;
        RECT 67.950 277.950 70.050 280.050 ;
        RECT 55.950 275.250 58.050 276.150 ;
        RECT 61.950 274.950 64.050 277.050 ;
        RECT 49.950 271.950 52.050 274.050 ;
        RECT 53.250 272.250 54.750 273.150 ;
        RECT 55.950 271.950 58.050 274.050 ;
        RECT 59.250 272.250 61.050 273.150 ;
        RECT 64.950 271.950 67.050 274.050 ;
        RECT 68.400 273.450 69.450 277.950 ;
        RECT 71.400 277.050 72.450 311.400 ;
        RECT 73.950 309.450 76.050 310.050 ;
        RECT 77.400 309.450 78.450 331.950 ;
        RECT 80.400 325.050 81.450 335.400 ;
        RECT 86.400 334.050 87.450 340.950 ;
        RECT 89.400 340.050 90.450 370.950 ;
        RECT 88.950 337.950 91.050 340.050 ;
        RECT 92.400 339.450 93.450 376.950 ;
        RECT 95.400 349.050 96.450 379.950 ;
        RECT 101.400 358.050 102.450 383.400 ;
        RECT 103.950 382.950 106.050 383.400 ;
        RECT 107.250 383.250 109.050 384.150 ;
        RECT 116.400 382.050 117.450 403.950 ;
        RECT 119.400 397.050 120.450 412.950 ;
        RECT 121.950 409.950 124.050 412.050 ;
        RECT 127.950 409.950 130.050 412.050 ;
        RECT 122.400 400.050 123.450 409.950 ;
        RECT 121.950 397.950 124.050 400.050 ;
        RECT 124.950 397.950 127.050 400.050 ;
        RECT 118.950 394.950 121.050 397.050 ;
        RECT 118.950 391.950 121.050 394.050 ;
        RECT 119.400 388.050 120.450 391.950 ;
        RECT 118.950 385.950 121.050 388.050 ;
        RECT 103.950 380.850 105.750 381.750 ;
        RECT 106.950 379.950 109.050 382.050 ;
        RECT 112.950 380.250 114.750 381.150 ;
        RECT 115.950 379.950 118.050 382.050 ;
        RECT 119.250 380.250 121.050 381.150 ;
        RECT 107.400 373.050 108.450 379.950 ;
        RECT 112.950 376.950 115.050 379.050 ;
        RECT 116.250 377.850 117.750 378.750 ;
        RECT 118.950 376.950 121.050 379.050 ;
        RECT 106.950 370.950 109.050 373.050 ;
        RECT 113.400 361.050 114.450 376.950 ;
        RECT 119.400 376.050 120.450 376.950 ;
        RECT 118.950 373.950 121.050 376.050 ;
        RECT 122.400 373.050 123.450 397.950 ;
        RECT 125.400 385.050 126.450 397.950 ;
        RECT 127.950 391.950 130.050 394.050 ;
        RECT 124.950 382.950 127.050 385.050 ;
        RECT 128.400 382.050 129.450 391.950 ;
        RECT 131.400 382.050 132.450 433.950 ;
        RECT 133.950 413.850 136.050 414.750 ;
        RECT 136.950 413.250 139.050 414.150 ;
        RECT 133.950 409.950 136.050 412.050 ;
        RECT 136.950 409.950 139.050 412.050 ;
        RECT 134.400 385.050 135.450 409.950 ;
        RECT 140.400 397.050 141.450 448.950 ;
        RECT 143.400 442.050 144.450 451.950 ;
        RECT 149.400 451.050 150.450 463.950 ;
        RECT 154.950 460.950 157.050 463.050 ;
        RECT 151.950 457.950 154.050 460.050 ;
        RECT 152.400 454.050 153.450 457.950 ;
        RECT 155.400 457.050 156.450 460.950 ;
        RECT 161.400 457.050 162.450 463.950 ;
        RECT 154.950 454.950 157.050 457.050 ;
        RECT 158.250 455.250 159.750 456.150 ;
        RECT 160.950 454.950 163.050 457.050 ;
        RECT 164.400 456.450 165.450 499.950 ;
        RECT 166.950 485.250 169.050 486.150 ;
        RECT 169.950 485.850 172.050 486.750 ;
        RECT 166.950 481.950 169.050 484.050 ;
        RECT 169.950 472.950 172.050 475.050 ;
        RECT 166.950 469.950 169.050 472.050 ;
        RECT 167.400 457.050 168.450 469.950 ;
        RECT 170.400 460.050 171.450 472.950 ;
        RECT 173.400 460.050 174.450 523.950 ;
        RECT 179.400 523.050 180.450 527.400 ;
        RECT 181.950 524.250 183.750 525.150 ;
        RECT 184.950 523.950 187.050 526.050 ;
        RECT 188.250 524.250 190.050 525.150 ;
        RECT 178.950 520.950 181.050 523.050 ;
        RECT 181.950 520.950 184.050 523.050 ;
        RECT 185.250 521.850 186.750 522.750 ;
        RECT 182.400 511.050 183.450 520.950 ;
        RECT 181.950 508.950 184.050 511.050 ;
        RECT 182.400 499.050 183.450 508.950 ;
        RECT 181.950 496.950 184.050 499.050 ;
        RECT 181.950 491.250 184.050 492.150 ;
        RECT 191.400 490.050 192.450 532.950 ;
        RECT 206.400 529.050 207.450 544.950 ;
        RECT 205.950 526.950 208.050 529.050 ;
        RECT 209.250 527.250 210.750 528.150 ;
        RECT 211.950 526.950 214.050 529.050 ;
        RECT 193.950 524.250 195.750 525.150 ;
        RECT 196.950 523.950 199.050 526.050 ;
        RECT 200.250 524.250 202.050 525.150 ;
        RECT 205.950 524.850 207.750 525.750 ;
        RECT 208.950 523.950 211.050 526.050 ;
        RECT 212.250 524.850 213.750 525.750 ;
        RECT 214.950 523.950 217.050 526.050 ;
        RECT 197.250 521.850 198.750 522.750 ;
        RECT 199.950 520.950 202.050 523.050 ;
        RECT 205.950 522.450 208.050 523.050 ;
        RECT 209.400 522.450 210.450 523.950 ;
        RECT 205.950 521.400 210.450 522.450 ;
        RECT 214.950 521.850 217.050 522.750 ;
        RECT 205.950 520.950 208.050 521.400 ;
        RECT 206.400 505.050 207.450 520.950 ;
        RECT 205.950 502.950 208.050 505.050 ;
        RECT 178.950 488.250 180.750 489.150 ;
        RECT 181.950 487.950 184.050 490.050 ;
        RECT 185.250 488.250 186.750 489.150 ;
        RECT 187.950 487.950 190.050 490.050 ;
        RECT 190.950 487.950 193.050 490.050 ;
        RECT 202.950 488.250 205.050 489.150 ;
        RECT 175.950 485.250 178.050 486.150 ;
        RECT 178.950 484.950 181.050 487.050 ;
        RECT 175.950 481.950 178.050 484.050 ;
        RECT 176.400 481.050 177.450 481.950 ;
        RECT 175.950 478.950 178.050 481.050 ;
        RECT 176.400 466.050 177.450 478.950 ;
        RECT 175.950 463.950 178.050 466.050 ;
        RECT 179.400 463.050 180.450 484.950 ;
        RECT 182.400 475.050 183.450 487.950 ;
        RECT 184.950 484.950 187.050 487.050 ;
        RECT 188.250 485.850 190.050 486.750 ;
        RECT 190.950 484.950 193.050 487.050 ;
        RECT 193.950 485.250 195.750 486.150 ;
        RECT 196.950 484.950 199.050 487.050 ;
        RECT 200.250 485.250 201.750 486.150 ;
        RECT 202.950 484.950 205.050 487.050 ;
        RECT 185.400 475.050 186.450 484.950 ;
        RECT 181.950 472.950 184.050 475.050 ;
        RECT 184.950 472.950 187.050 475.050 ;
        RECT 181.950 466.950 184.050 469.050 ;
        RECT 178.950 460.950 181.050 463.050 ;
        RECT 169.950 457.950 172.050 460.050 ;
        RECT 172.950 457.950 175.050 460.050 ;
        RECT 175.950 457.950 178.050 460.050 ;
        RECT 166.950 456.450 169.050 457.050 ;
        RECT 164.400 455.400 169.050 456.450 ;
        RECT 170.250 455.850 171.750 456.750 ;
        RECT 172.950 456.450 175.050 457.050 ;
        RECT 176.400 456.450 177.450 457.950 ;
        RECT 151.950 451.950 154.050 454.050 ;
        RECT 155.250 452.850 156.750 453.750 ;
        RECT 157.950 451.950 160.050 454.050 ;
        RECT 161.250 452.850 163.050 453.750 ;
        RECT 148.950 448.950 151.050 451.050 ;
        RECT 151.950 449.850 154.050 450.750 ;
        RECT 158.400 445.050 159.450 451.950 ;
        RECT 151.950 442.950 154.050 445.050 ;
        RECT 157.950 442.950 160.050 445.050 ;
        RECT 142.950 439.950 145.050 442.050 ;
        RECT 145.950 416.250 148.050 417.150 ;
        RECT 152.400 415.050 153.450 442.950 ;
        RECT 164.400 442.050 165.450 455.400 ;
        RECT 166.950 454.950 169.050 455.400 ;
        RECT 172.950 455.400 177.450 456.450 ;
        RECT 172.950 454.950 175.050 455.400 ;
        RECT 176.400 454.050 177.450 455.400 ;
        RECT 179.400 454.050 180.450 460.950 ;
        RECT 182.400 457.050 183.450 466.950 ;
        RECT 187.950 460.950 190.050 463.050 ;
        RECT 188.400 457.050 189.450 460.950 ;
        RECT 191.400 457.050 192.450 484.950 ;
        RECT 193.950 481.950 196.050 484.050 ;
        RECT 197.250 482.850 198.750 483.750 ;
        RECT 199.950 481.950 202.050 484.050 ;
        RECT 194.400 463.050 195.450 481.950 ;
        RECT 200.400 481.050 201.450 481.950 ;
        RECT 199.950 478.950 202.050 481.050 ;
        RECT 206.400 468.450 207.450 502.950 ;
        RECT 214.950 499.950 217.050 502.050 ;
        RECT 215.400 490.050 216.450 499.950 ;
        RECT 208.950 487.950 211.050 490.050 ;
        RECT 212.250 488.250 213.750 489.150 ;
        RECT 214.950 487.950 217.050 490.050 ;
        RECT 208.950 485.850 210.750 486.750 ;
        RECT 211.950 484.950 214.050 487.050 ;
        RECT 215.250 485.850 217.050 486.750 ;
        RECT 212.400 475.050 213.450 484.950 ;
        RECT 214.950 481.950 217.050 484.050 ;
        RECT 211.950 472.950 214.050 475.050 ;
        RECT 208.950 469.950 211.050 472.050 ;
        RECT 203.400 467.400 207.450 468.450 ;
        RECT 193.950 460.950 196.050 463.050 ;
        RECT 181.950 454.950 184.050 457.050 ;
        RECT 185.250 455.250 186.750 456.150 ;
        RECT 187.950 454.950 190.050 457.050 ;
        RECT 190.950 454.950 193.050 457.050 ;
        RECT 194.400 454.050 195.450 460.950 ;
        RECT 166.950 452.850 169.050 453.750 ;
        RECT 172.950 452.850 175.050 453.750 ;
        RECT 175.950 451.950 178.050 454.050 ;
        RECT 178.950 451.950 181.050 454.050 ;
        RECT 182.250 452.850 183.750 453.750 ;
        RECT 184.950 451.950 187.050 454.050 ;
        RECT 188.250 452.850 190.050 453.750 ;
        RECT 190.950 452.250 192.750 453.150 ;
        RECT 193.950 451.950 196.050 454.050 ;
        RECT 197.250 452.250 199.050 453.150 ;
        RECT 163.950 439.950 166.050 442.050 ;
        RECT 176.400 433.050 177.450 451.950 ;
        RECT 178.950 449.850 181.050 450.750 ;
        RECT 187.950 448.950 190.050 451.050 ;
        RECT 190.950 448.950 193.050 451.050 ;
        RECT 194.250 449.850 195.750 450.750 ;
        RECT 203.400 450.450 204.450 467.400 ;
        RECT 209.400 465.450 210.450 469.950 ;
        RECT 206.400 464.400 210.450 465.450 ;
        RECT 206.400 457.050 207.450 464.400 ;
        RECT 205.950 454.950 208.050 457.050 ;
        RECT 209.250 455.250 211.050 456.150 ;
        RECT 215.400 454.050 216.450 481.950 ;
        RECT 218.400 481.050 219.450 550.950 ;
        RECT 233.400 550.050 234.450 553.950 ;
        RECT 236.400 553.050 237.450 559.950 ;
        RECT 245.400 559.050 246.450 562.950 ;
        RECT 238.950 556.950 241.050 559.050 ;
        RECT 244.950 556.950 247.050 559.050 ;
        RECT 250.950 556.950 253.050 559.050 ;
        RECT 254.250 557.250 256.050 558.150 ;
        RECT 257.400 556.050 258.450 593.400 ;
        RECT 259.950 592.950 262.050 593.400 ;
        RECT 263.400 559.050 264.450 598.950 ;
        RECT 265.950 596.850 268.050 597.750 ;
        RECT 259.950 557.250 262.050 558.150 ;
        RECT 262.950 556.950 265.050 559.050 ;
        RECT 265.950 557.250 268.050 558.150 ;
        RECT 238.950 554.850 241.050 555.750 ;
        RECT 241.950 554.250 244.050 555.150 ;
        RECT 244.950 554.850 247.050 555.750 ;
        RECT 247.950 554.250 250.050 555.150 ;
        RECT 250.950 554.850 252.750 555.750 ;
        RECT 253.950 553.950 256.050 556.050 ;
        RECT 256.950 553.950 259.050 556.050 ;
        RECT 259.950 553.950 262.050 556.050 ;
        RECT 263.250 554.250 264.750 555.150 ;
        RECT 265.950 553.950 268.050 556.050 ;
        RECT 235.950 550.950 238.050 553.050 ;
        RECT 241.950 550.950 244.050 553.050 ;
        RECT 247.950 550.950 250.050 553.050 ;
        RECT 262.950 550.950 265.050 553.050 ;
        RECT 232.950 547.950 235.050 550.050 ;
        RECT 244.950 544.950 247.050 547.050 ;
        RECT 235.950 541.950 238.050 544.050 ;
        RECT 229.950 538.950 232.050 541.050 ;
        RECT 226.950 533.400 229.050 535.500 ;
        RECT 227.400 516.600 228.600 533.400 ;
        RECT 230.400 519.450 231.450 538.950 ;
        RECT 232.950 526.950 235.050 529.050 ;
        RECT 232.950 524.850 235.050 525.750 ;
        RECT 230.400 518.400 234.450 519.450 ;
        RECT 226.950 514.500 229.050 516.600 ;
        RECT 220.950 508.950 223.050 511.050 ;
        RECT 217.950 478.950 220.050 481.050 ;
        RECT 221.400 475.050 222.450 508.950 ;
        RECT 223.950 487.950 226.050 490.050 ;
        RECT 226.950 487.950 229.050 490.050 ;
        RECT 224.400 487.050 225.450 487.950 ;
        RECT 223.950 484.950 226.050 487.050 ;
        RECT 223.950 482.850 226.050 483.750 ;
        RECT 227.400 478.050 228.450 487.950 ;
        RECT 233.400 487.050 234.450 518.400 ;
        RECT 229.950 485.250 232.050 486.150 ;
        RECT 232.950 484.950 235.050 487.050 ;
        RECT 229.950 481.950 232.050 484.050 ;
        RECT 233.250 482.250 235.050 483.150 ;
        RECT 232.950 478.950 235.050 481.050 ;
        RECT 223.950 475.950 226.050 478.050 ;
        RECT 226.950 475.950 229.050 478.050 ;
        RECT 232.950 475.950 235.050 478.050 ;
        RECT 220.950 472.950 223.050 475.050 ;
        RECT 224.400 466.050 225.450 475.950 ;
        RECT 223.950 463.950 226.050 466.050 ;
        RECT 220.950 460.950 223.050 463.050 ;
        RECT 226.950 460.950 229.050 463.050 ;
        RECT 205.950 452.850 207.750 453.750 ;
        RECT 211.950 452.250 213.750 453.150 ;
        RECT 214.950 451.950 217.050 454.050 ;
        RECT 218.250 452.250 220.050 453.150 ;
        RECT 221.400 451.050 222.450 460.950 ;
        RECT 227.400 454.050 228.450 460.950 ;
        RECT 233.400 454.050 234.450 475.950 ;
        RECT 236.400 468.450 237.450 541.950 ;
        RECT 238.950 532.950 241.050 535.050 ;
        RECT 239.400 529.050 240.450 532.950 ;
        RECT 238.950 526.950 241.050 529.050 ;
        RECT 238.950 524.850 241.050 525.750 ;
        RECT 238.950 520.950 241.050 523.050 ;
        RECT 239.400 493.050 240.450 520.950 ;
        RECT 245.400 499.050 246.450 544.950 ;
        RECT 247.950 533.400 250.050 535.500 ;
        RECT 248.250 521.400 249.450 533.400 ;
        RECT 269.400 532.050 270.450 604.950 ;
        RECT 271.950 601.950 274.050 604.050 ;
        RECT 272.400 598.050 273.450 601.950 ;
        RECT 281.400 601.050 282.450 610.950 ;
        RECT 290.400 607.050 291.450 625.950 ;
        RECT 295.950 622.950 298.050 625.050 ;
        RECT 289.950 604.950 292.050 607.050 ;
        RECT 286.950 601.950 289.050 604.050 ;
        RECT 290.400 601.050 291.450 604.950 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 274.950 598.950 277.050 601.050 ;
        RECT 280.950 600.450 283.050 601.050 ;
        RECT 283.950 600.450 286.050 601.050 ;
        RECT 278.250 599.250 279.750 600.150 ;
        RECT 280.950 599.400 286.050 600.450 ;
        RECT 287.250 599.850 288.750 600.750 ;
        RECT 280.950 598.950 283.050 599.400 ;
        RECT 283.950 598.950 286.050 599.400 ;
        RECT 289.950 598.950 292.050 601.050 ;
        RECT 271.950 595.950 274.050 598.050 ;
        RECT 275.250 596.850 276.750 597.750 ;
        RECT 277.950 595.950 280.050 598.050 ;
        RECT 281.250 596.850 283.050 597.750 ;
        RECT 283.950 596.850 286.050 597.750 ;
        RECT 286.950 595.950 289.050 598.050 ;
        RECT 289.950 596.850 292.050 597.750 ;
        RECT 278.400 595.050 279.450 595.950 ;
        RECT 271.950 593.850 274.050 594.750 ;
        RECT 274.950 592.950 277.050 595.050 ;
        RECT 277.950 592.950 280.050 595.050 ;
        RECT 271.950 589.950 274.050 592.050 ;
        RECT 272.400 556.050 273.450 589.950 ;
        RECT 275.400 561.450 276.450 592.950 ;
        RECT 283.950 562.950 286.050 565.050 ;
        RECT 275.400 560.400 279.450 561.450 ;
        RECT 278.400 559.050 279.450 560.400 ;
        RECT 284.400 559.050 285.450 562.950 ;
        RECT 274.950 557.250 276.750 558.150 ;
        RECT 277.950 556.950 280.050 559.050 ;
        RECT 283.950 556.950 286.050 559.050 ;
        RECT 271.950 553.950 274.050 556.050 ;
        RECT 274.950 553.950 277.050 556.050 ;
        RECT 278.250 554.850 280.050 555.750 ;
        RECT 280.950 554.250 283.050 555.150 ;
        RECT 283.950 554.850 286.050 555.750 ;
        RECT 275.400 550.050 276.450 553.950 ;
        RECT 287.400 553.050 288.450 595.950 ;
        RECT 293.400 565.050 294.450 601.950 ;
        RECT 296.400 598.050 297.450 622.950 ;
        RECT 299.400 616.050 300.450 628.950 ;
        RECT 298.950 613.950 301.050 616.050 ;
        RECT 301.950 603.450 304.050 604.050 ;
        RECT 305.400 603.450 306.450 658.950 ;
        RECT 314.400 649.050 315.450 671.400 ;
        RECT 319.950 671.250 322.050 672.150 ;
        RECT 325.950 670.950 328.050 673.050 ;
        RECT 329.250 671.250 330.750 672.150 ;
        RECT 331.950 670.950 334.050 673.050 ;
        RECT 319.950 667.950 322.050 670.050 ;
        RECT 325.950 668.850 327.750 669.750 ;
        RECT 328.950 667.950 331.050 670.050 ;
        RECT 332.250 668.850 333.750 669.750 ;
        RECT 334.950 669.450 337.050 670.050 ;
        RECT 334.950 668.400 339.450 669.450 ;
        RECT 334.950 667.950 337.050 668.400 ;
        RECT 338.400 667.050 339.450 668.400 ;
        RECT 334.950 665.850 337.050 666.750 ;
        RECT 337.950 664.950 340.050 667.050 ;
        RECT 313.950 646.950 316.050 649.050 ;
        RECT 316.950 640.950 319.050 643.050 ;
        RECT 310.950 635.250 313.050 636.150 ;
        RECT 317.400 634.050 318.450 640.950 ;
        RECT 328.950 638.400 331.050 640.500 ;
        RECT 307.950 632.250 309.750 633.150 ;
        RECT 310.950 631.950 313.050 634.050 ;
        RECT 314.250 632.250 315.750 633.150 ;
        RECT 316.950 631.950 319.050 634.050 ;
        RECT 307.950 628.950 310.050 631.050 ;
        RECT 308.400 607.050 309.450 628.950 ;
        RECT 311.400 622.050 312.450 631.950 ;
        RECT 313.950 628.950 316.050 631.050 ;
        RECT 317.250 629.850 319.050 630.750 ;
        RECT 310.950 619.950 313.050 622.050 ;
        RECT 329.400 621.600 330.600 638.400 ;
        RECT 341.400 633.450 342.450 679.950 ;
        RECT 343.950 676.950 346.050 679.050 ;
        RECT 344.400 673.050 345.450 676.950 ;
        RECT 350.400 673.050 351.450 679.950 ;
        RECT 412.950 677.400 415.050 679.500 ;
        RECT 433.950 677.400 436.050 679.500 ;
        RECT 358.950 673.950 361.050 676.050 ;
        RECT 370.950 673.950 373.050 676.050 ;
        RECT 376.950 673.950 379.050 676.050 ;
        RECT 343.950 670.950 346.050 673.050 ;
        RECT 347.250 671.250 348.750 672.150 ;
        RECT 349.950 670.950 352.050 673.050 ;
        RECT 353.250 671.250 354.750 672.150 ;
        RECT 355.950 670.950 358.050 673.050 ;
        RECT 358.950 671.850 360.750 672.750 ;
        RECT 361.950 672.450 364.050 673.050 ;
        RECT 364.950 672.450 367.050 673.050 ;
        RECT 361.950 671.400 367.050 672.450 ;
        RECT 361.950 670.950 364.050 671.400 ;
        RECT 364.950 670.950 367.050 671.400 ;
        RECT 367.950 671.250 370.050 672.150 ;
        RECT 343.950 668.850 345.750 669.750 ;
        RECT 346.950 667.950 349.050 670.050 ;
        RECT 350.250 668.850 351.750 669.750 ;
        RECT 352.950 667.950 355.050 670.050 ;
        RECT 356.250 668.850 358.050 669.750 ;
        RECT 361.950 668.850 364.050 669.750 ;
        RECT 353.400 667.050 354.450 667.950 ;
        RECT 352.950 666.450 355.050 667.050 ;
        RECT 352.950 665.400 357.450 666.450 ;
        RECT 352.950 664.950 355.050 665.400 ;
        RECT 349.950 639.300 352.050 641.400 ;
        RECT 350.250 635.700 351.450 639.300 ;
        RECT 349.950 633.600 352.050 635.700 ;
        RECT 338.400 632.400 342.450 633.450 ;
        RECT 334.950 629.250 337.050 630.150 ;
        RECT 334.950 627.450 337.050 628.050 ;
        RECT 338.400 627.450 339.450 632.400 ;
        RECT 340.950 629.250 343.050 630.150 ;
        RECT 334.950 626.400 339.450 627.450 ;
        RECT 334.950 625.950 337.050 626.400 ;
        RECT 340.950 625.950 343.050 628.050 ;
        RECT 328.950 619.500 331.050 621.600 ;
        RECT 319.950 616.950 322.050 619.050 ;
        RECT 325.950 616.950 328.050 619.050 ;
        RECT 310.950 613.950 313.050 616.050 ;
        RECT 307.950 604.950 310.050 607.050 ;
        RECT 301.950 602.400 306.450 603.450 ;
        RECT 301.950 601.950 304.050 602.400 ;
        RECT 305.400 601.050 306.450 602.400 ;
        RECT 311.400 601.050 312.450 613.950 ;
        RECT 320.400 604.050 321.450 616.950 ;
        RECT 319.950 601.950 322.050 604.050 ;
        RECT 298.950 599.250 301.050 600.150 ;
        RECT 301.950 599.850 304.050 600.750 ;
        RECT 304.950 598.950 307.050 601.050 ;
        RECT 308.250 599.250 309.750 600.150 ;
        RECT 310.950 598.950 313.050 601.050 ;
        RECT 319.950 599.850 322.050 600.750 ;
        RECT 322.950 599.250 325.050 600.150 ;
        RECT 295.950 595.950 298.050 598.050 ;
        RECT 298.950 595.950 301.050 598.050 ;
        RECT 304.950 596.850 306.750 597.750 ;
        RECT 307.950 595.950 310.050 598.050 ;
        RECT 311.250 596.850 312.750 597.750 ;
        RECT 313.950 595.950 316.050 598.050 ;
        RECT 322.950 595.950 325.050 598.050 ;
        RECT 299.400 595.050 300.450 595.950 ;
        RECT 298.950 592.950 301.050 595.050 ;
        RECT 308.400 594.450 309.450 595.950 ;
        RECT 308.400 593.400 312.450 594.450 ;
        RECT 313.950 593.850 316.050 594.750 ;
        RECT 326.400 594.450 327.450 616.950 ;
        RECT 341.400 613.050 342.450 625.950 ;
        RECT 350.250 621.600 351.450 633.600 ;
        RECT 352.950 625.950 355.050 628.050 ;
        RECT 352.950 623.850 355.050 624.750 ;
        RECT 349.950 619.500 352.050 621.600 ;
        RECT 346.950 613.950 349.050 616.050 ;
        RECT 340.950 610.950 343.050 613.050 ;
        RECT 337.950 607.950 340.050 610.050 ;
        RECT 328.950 596.250 330.750 597.150 ;
        RECT 331.950 595.950 334.050 598.050 ;
        RECT 335.250 596.250 337.050 597.150 ;
        RECT 328.950 594.450 331.050 595.050 ;
        RECT 326.400 593.400 331.050 594.450 ;
        RECT 332.250 593.850 333.750 594.750 ;
        RECT 334.950 594.450 337.050 595.050 ;
        RECT 338.400 594.450 339.450 607.950 ;
        RECT 340.950 604.950 343.050 607.050 ;
        RECT 341.400 601.050 342.450 604.950 ;
        RECT 340.950 598.950 343.050 601.050 ;
        RECT 341.400 598.050 342.450 598.950 ;
        RECT 347.400 598.050 348.450 613.950 ;
        RECT 356.400 607.050 357.450 665.400 ;
        RECT 365.400 664.050 366.450 670.950 ;
        RECT 367.950 667.950 370.050 670.050 ;
        RECT 371.400 669.450 372.450 673.950 ;
        RECT 373.950 671.250 376.050 672.150 ;
        RECT 376.950 671.850 379.050 672.750 ;
        RECT 382.950 672.450 385.050 673.050 ;
        RECT 379.950 671.250 381.750 672.150 ;
        RECT 382.950 671.400 387.450 672.450 ;
        RECT 382.950 670.950 385.050 671.400 ;
        RECT 373.950 669.450 376.050 670.050 ;
        RECT 371.400 668.400 376.050 669.450 ;
        RECT 373.950 667.950 376.050 668.400 ;
        RECT 379.950 667.950 382.050 670.050 ;
        RECT 383.250 668.850 385.050 669.750 ;
        RECT 380.400 667.050 381.450 667.950 ;
        RECT 373.950 664.950 376.050 667.050 ;
        RECT 379.950 664.950 382.050 667.050 ;
        RECT 364.950 661.950 367.050 664.050 ;
        RECT 374.400 631.050 375.450 664.950 ;
        RECT 386.400 664.050 387.450 671.400 ;
        RECT 391.950 670.950 394.050 673.050 ;
        RECT 395.250 671.250 396.750 672.150 ;
        RECT 397.950 670.950 400.050 673.050 ;
        RECT 403.950 672.450 406.050 673.050 ;
        RECT 401.250 671.250 402.750 672.150 ;
        RECT 403.950 671.400 408.450 672.450 ;
        RECT 403.950 670.950 406.050 671.400 ;
        RECT 407.400 670.050 408.450 671.400 ;
        RECT 391.950 668.850 393.750 669.750 ;
        RECT 394.950 667.950 397.050 670.050 ;
        RECT 398.250 668.850 399.750 669.750 ;
        RECT 400.950 667.950 403.050 670.050 ;
        RECT 404.250 668.850 406.050 669.750 ;
        RECT 406.950 667.950 409.050 670.050 ;
        RECT 395.400 664.050 396.450 667.950 ;
        RECT 401.400 667.050 402.450 667.950 ;
        RECT 400.950 664.950 403.050 667.050 ;
        RECT 385.950 661.950 388.050 664.050 ;
        RECT 394.950 661.950 397.050 664.050 ;
        RECT 397.950 639.300 400.050 641.400 ;
        RECT 398.550 635.700 399.750 639.300 ;
        RECT 401.400 637.050 402.450 664.950 ;
        RECT 413.400 660.600 414.600 677.400 ;
        RECT 418.950 670.950 421.050 673.050 ;
        RECT 424.950 672.450 427.050 673.050 ;
        RECT 422.400 671.400 427.050 672.450 ;
        RECT 418.950 668.850 421.050 669.750 ;
        RECT 412.950 658.500 415.050 660.600 ;
        RECT 418.950 638.400 421.050 640.500 ;
        RECT 397.950 633.600 400.050 635.700 ;
        RECT 400.950 634.950 403.050 637.050 ;
        RECT 358.950 629.250 361.050 630.150 ;
        RECT 364.950 629.250 367.050 630.150 ;
        RECT 373.950 628.950 376.050 631.050 ;
        RECT 382.950 629.250 385.050 630.150 ;
        RECT 388.950 629.250 391.050 630.150 ;
        RECT 358.950 625.950 361.050 628.050 ;
        RECT 373.950 626.850 376.050 627.750 ;
        RECT 376.950 626.250 379.050 627.150 ;
        RECT 382.950 625.950 385.050 628.050 ;
        RECT 386.250 626.250 387.750 627.150 ;
        RECT 388.950 625.950 391.050 628.050 ;
        RECT 394.950 625.950 397.050 628.050 ;
        RECT 355.950 604.950 358.050 607.050 ;
        RECT 359.400 604.050 360.450 625.950 ;
        RECT 383.400 625.050 384.450 625.950 ;
        RECT 389.400 625.050 390.450 625.950 ;
        RECT 376.950 622.950 379.050 625.050 ;
        RECT 382.950 622.950 385.050 625.050 ;
        RECT 385.950 622.950 388.050 625.050 ;
        RECT 388.950 622.950 391.050 625.050 ;
        RECT 394.950 623.850 397.050 624.750 ;
        RECT 386.400 604.050 387.450 622.950 ;
        RECT 398.550 621.600 399.750 633.600 ;
        RECT 397.950 619.500 400.050 621.600 ;
        RECT 358.950 601.950 361.050 604.050 ;
        RECT 364.950 601.950 367.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 352.950 598.950 355.050 601.050 ;
        RECT 355.950 600.450 358.050 601.050 ;
        RECT 355.950 599.400 360.450 600.450 ;
        RECT 355.950 598.950 358.050 599.400 ;
        RECT 340.950 595.950 343.050 598.050 ;
        RECT 343.950 595.950 346.050 598.050 ;
        RECT 346.950 595.950 349.050 598.050 ;
        RECT 350.250 596.250 352.050 597.150 ;
        RECT 344.400 595.050 345.450 595.950 ;
        RECT 292.950 562.950 295.050 565.050 ;
        RECT 289.950 559.950 292.050 562.050 ;
        RECT 293.250 560.250 294.750 561.150 ;
        RECT 295.950 559.950 298.050 562.050 ;
        RECT 289.950 557.850 291.750 558.750 ;
        RECT 292.950 556.950 295.050 559.050 ;
        RECT 296.250 557.850 298.050 558.750 ;
        RECT 301.950 557.250 304.050 558.150 ;
        RECT 307.950 556.950 310.050 559.050 ;
        RECT 293.400 556.050 294.450 556.950 ;
        RECT 292.950 553.950 295.050 556.050 ;
        RECT 301.950 555.450 304.050 556.050 ;
        RECT 298.950 554.250 300.750 555.150 ;
        RECT 301.950 554.400 306.450 555.450 ;
        RECT 307.950 554.850 310.050 555.750 ;
        RECT 301.950 553.950 304.050 554.400 ;
        RECT 280.950 550.950 283.050 553.050 ;
        RECT 286.950 550.950 289.050 553.050 ;
        RECT 292.950 550.950 295.050 553.050 ;
        RECT 298.950 550.950 301.050 553.050 ;
        RECT 274.950 547.950 277.050 550.050 ;
        RECT 250.950 530.250 253.050 531.150 ;
        RECT 253.950 529.950 256.050 532.050 ;
        RECT 268.950 529.950 271.050 532.050 ;
        RECT 274.950 529.950 277.050 532.050 ;
        RECT 250.950 526.950 253.050 529.050 ;
        RECT 251.400 523.050 252.450 526.950 ;
        RECT 247.950 519.300 250.050 521.400 ;
        RECT 250.950 520.950 253.050 523.050 ;
        RECT 248.250 515.700 249.450 519.300 ;
        RECT 247.950 513.600 250.050 515.700 ;
        RECT 250.950 511.950 253.050 514.050 ;
        RECT 251.400 508.050 252.450 511.950 ;
        RECT 250.950 505.950 253.050 508.050 ;
        RECT 244.950 496.950 247.050 499.050 ;
        RECT 238.950 490.950 241.050 493.050 ;
        RECT 238.950 487.950 241.050 490.050 ;
        RECT 242.250 488.250 243.750 489.150 ;
        RECT 244.950 487.950 247.050 490.050 ;
        RECT 251.400 487.050 252.450 505.950 ;
        RECT 254.400 490.050 255.450 529.950 ;
        RECT 275.400 529.050 276.450 529.950 ;
        RECT 256.950 526.950 259.050 529.050 ;
        RECT 268.950 526.950 271.050 529.050 ;
        RECT 272.250 527.250 273.750 528.150 ;
        RECT 274.950 526.950 277.050 529.050 ;
        RECT 257.400 511.050 258.450 526.950 ;
        RECT 259.950 524.250 261.750 525.150 ;
        RECT 262.950 523.950 265.050 526.050 ;
        RECT 266.250 524.250 268.050 525.150 ;
        RECT 268.950 524.850 270.750 525.750 ;
        RECT 271.950 523.950 274.050 526.050 ;
        RECT 275.250 524.850 276.750 525.750 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 259.950 520.950 262.050 523.050 ;
        RECT 263.250 521.850 264.750 522.750 ;
        RECT 265.950 520.950 268.050 523.050 ;
        RECT 260.400 520.050 261.450 520.950 ;
        RECT 259.950 517.950 262.050 520.050 ;
        RECT 262.950 517.950 265.050 520.050 ;
        RECT 256.950 508.950 259.050 511.050 ;
        RECT 259.950 502.950 262.050 505.050 ;
        RECT 253.950 487.950 256.050 490.050 ;
        RECT 256.950 488.250 259.050 489.150 ;
        RECT 238.950 485.850 240.750 486.750 ;
        RECT 241.950 484.950 244.050 487.050 ;
        RECT 245.250 485.850 247.050 486.750 ;
        RECT 247.950 485.250 249.750 486.150 ;
        RECT 250.950 484.950 253.050 487.050 ;
        RECT 254.250 485.250 255.750 486.150 ;
        RECT 256.950 484.950 259.050 487.050 ;
        RECT 257.400 484.050 258.450 484.950 ;
        RECT 247.950 483.450 250.050 484.050 ;
        RECT 245.400 482.400 250.050 483.450 ;
        RECT 251.250 482.850 252.750 483.750 ;
        RECT 241.950 472.950 244.050 475.050 ;
        RECT 236.400 467.400 240.450 468.450 ;
        RECT 235.950 454.950 238.050 457.050 ;
        RECT 223.950 452.250 225.750 453.150 ;
        RECT 226.950 451.950 229.050 454.050 ;
        RECT 230.250 452.250 232.050 453.150 ;
        RECT 232.950 451.950 235.050 454.050 ;
        RECT 235.950 452.850 238.050 453.750 ;
        RECT 203.400 449.400 207.450 450.450 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 166.950 430.950 169.050 433.050 ;
        RECT 175.950 430.950 178.050 433.050 ;
        RECT 161.250 416.250 162.750 417.150 ;
        RECT 163.950 415.950 166.050 418.050 ;
        RECT 145.950 412.950 148.050 415.050 ;
        RECT 149.250 413.250 150.750 414.150 ;
        RECT 151.950 412.950 154.050 415.050 ;
        RECT 155.250 413.250 157.050 414.150 ;
        RECT 157.950 413.850 159.750 414.750 ;
        RECT 160.950 412.950 163.050 415.050 ;
        RECT 164.250 413.850 166.050 414.750 ;
        RECT 146.400 412.050 147.450 412.950 ;
        RECT 161.400 412.050 162.450 412.950 ;
        RECT 145.950 409.950 148.050 412.050 ;
        RECT 148.950 409.950 151.050 412.050 ;
        RECT 152.250 410.850 153.750 411.750 ;
        RECT 154.950 409.950 157.050 412.050 ;
        RECT 157.950 409.950 160.050 412.050 ;
        RECT 160.950 409.950 163.050 412.050 ;
        RECT 145.950 397.950 148.050 400.050 ;
        RECT 139.950 394.950 142.050 397.050 ;
        RECT 136.950 385.950 139.050 388.050 ;
        RECT 133.950 382.950 136.050 385.050 ;
        RECT 124.950 380.250 126.750 381.150 ;
        RECT 127.950 379.950 130.050 382.050 ;
        RECT 130.950 379.950 133.050 382.050 ;
        RECT 133.950 381.450 136.050 382.050 ;
        RECT 137.400 381.450 138.450 385.950 ;
        RECT 140.400 382.050 141.450 394.950 ;
        RECT 146.400 388.050 147.450 397.950 ;
        RECT 149.400 397.050 150.450 409.950 ;
        RECT 151.950 406.950 154.050 409.050 ;
        RECT 148.950 394.950 151.050 397.050 ;
        RECT 142.950 385.950 145.050 388.050 ;
        RECT 145.950 385.950 148.050 388.050 ;
        RECT 143.400 385.050 144.450 385.950 ;
        RECT 152.400 385.050 153.450 406.950 ;
        RECT 155.400 406.050 156.450 409.950 ;
        RECT 154.950 403.950 157.050 406.050 ;
        RECT 154.950 391.950 157.050 394.050 ;
        RECT 142.950 382.950 145.050 385.050 ;
        RECT 146.250 383.250 147.750 384.150 ;
        RECT 148.950 382.950 151.050 385.050 ;
        RECT 151.950 382.950 154.050 385.050 ;
        RECT 155.400 382.050 156.450 391.950 ;
        RECT 158.400 385.050 159.450 409.950 ;
        RECT 167.400 406.050 168.450 430.950 ;
        RECT 178.950 418.950 181.050 421.050 ;
        RECT 179.400 418.050 180.450 418.950 ;
        RECT 172.950 416.250 175.050 417.150 ;
        RECT 178.950 415.950 181.050 418.050 ;
        RECT 179.400 415.050 180.450 415.950 ;
        RECT 172.950 412.950 175.050 415.050 ;
        RECT 176.250 413.250 177.750 414.150 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 182.250 413.250 184.050 414.150 ;
        RECT 173.400 412.050 174.450 412.950 ;
        RECT 172.950 409.950 175.050 412.050 ;
        RECT 175.950 409.950 178.050 412.050 ;
        RECT 179.250 410.850 180.750 411.750 ;
        RECT 181.950 409.950 184.050 412.050 ;
        RECT 185.400 411.450 186.450 445.950 ;
        RECT 188.400 418.050 189.450 448.950 ;
        RECT 193.950 442.950 196.050 445.050 ;
        RECT 190.950 423.300 193.050 425.400 ;
        RECT 191.550 419.700 192.750 423.300 ;
        RECT 187.950 415.950 190.050 418.050 ;
        RECT 190.950 417.600 193.050 419.700 ;
        RECT 187.950 411.450 190.050 412.050 ;
        RECT 185.400 410.400 190.050 411.450 ;
        RECT 182.400 406.050 183.450 409.950 ;
        RECT 166.950 403.950 169.050 406.050 ;
        RECT 181.950 403.950 184.050 406.050 ;
        RECT 185.400 397.050 186.450 410.400 ;
        RECT 187.950 409.950 190.050 410.400 ;
        RECT 187.950 407.850 190.050 408.750 ;
        RECT 187.950 403.950 190.050 406.050 ;
        RECT 191.550 405.600 192.750 417.600 ;
        RECT 194.400 409.050 195.450 442.950 ;
        RECT 202.950 430.950 205.050 433.050 ;
        RECT 203.400 415.050 204.450 430.950 ;
        RECT 206.400 421.050 207.450 449.400 ;
        RECT 211.950 448.950 214.050 451.050 ;
        RECT 215.250 449.850 216.750 450.750 ;
        RECT 220.950 448.950 223.050 451.050 ;
        RECT 223.950 448.950 226.050 451.050 ;
        RECT 227.250 449.850 228.750 450.750 ;
        RECT 232.950 448.950 235.050 451.050 ;
        RECT 212.400 447.450 213.450 448.950 ;
        RECT 212.400 446.400 216.450 447.450 ;
        RECT 211.950 422.400 214.050 424.500 ;
        RECT 205.950 418.950 208.050 421.050 ;
        RECT 199.950 413.250 202.050 414.150 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 205.950 413.250 208.050 414.150 ;
        RECT 199.950 409.950 202.050 412.050 ;
        RECT 193.950 406.950 196.050 409.050 ;
        RECT 169.950 394.950 172.050 397.050 ;
        RECT 172.950 394.950 175.050 397.050 ;
        RECT 184.950 394.950 187.050 397.050 ;
        RECT 157.950 382.950 160.050 385.050 ;
        RECT 170.400 382.050 171.450 394.950 ;
        RECT 173.400 382.050 174.450 394.950 ;
        RECT 175.950 388.950 178.050 391.050 ;
        RECT 184.950 388.950 187.050 391.050 ;
        RECT 176.400 382.050 177.450 388.950 ;
        RECT 185.400 388.050 186.450 388.950 ;
        RECT 178.950 385.950 181.050 388.050 ;
        RECT 184.950 385.950 187.050 388.050 ;
        RECT 133.950 380.400 138.450 381.450 ;
        RECT 133.950 379.950 136.050 380.400 ;
        RECT 139.950 379.950 142.050 382.050 ;
        RECT 143.250 380.850 144.750 381.750 ;
        RECT 145.950 379.950 148.050 382.050 ;
        RECT 149.250 380.850 151.050 381.750 ;
        RECT 151.950 380.250 153.750 381.150 ;
        RECT 154.950 379.950 157.050 382.050 ;
        RECT 158.250 380.250 160.050 381.150 ;
        RECT 166.950 380.250 168.750 381.150 ;
        RECT 169.950 379.950 172.050 382.050 ;
        RECT 172.950 379.950 175.050 382.050 ;
        RECT 175.950 379.950 178.050 382.050 ;
        RECT 179.400 381.450 180.450 385.950 ;
        RECT 181.950 383.250 184.050 384.150 ;
        RECT 184.950 383.850 187.050 384.750 ;
        RECT 181.950 381.450 184.050 382.050 ;
        RECT 179.400 380.400 184.050 381.450 ;
        RECT 181.950 379.950 184.050 380.400 ;
        RECT 124.950 376.950 127.050 379.050 ;
        RECT 128.250 377.850 129.750 378.750 ;
        RECT 130.950 376.950 133.050 379.050 ;
        RECT 134.250 377.850 136.050 378.750 ;
        RECT 139.950 377.850 142.050 378.750 ;
        RECT 142.950 376.950 145.050 379.050 ;
        RECT 130.950 374.850 133.050 375.750 ;
        RECT 139.950 373.950 142.050 376.050 ;
        RECT 121.950 370.950 124.050 373.050 ;
        RECT 124.950 370.950 127.050 373.050 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 112.950 358.950 115.050 361.050 ;
        RECT 100.950 355.950 103.050 358.050 ;
        RECT 112.950 352.950 115.050 355.050 ;
        RECT 94.950 346.950 97.050 349.050 ;
        RECT 97.950 343.950 100.050 346.050 ;
        RECT 109.950 343.950 112.050 346.050 ;
        RECT 98.400 343.050 99.450 343.950 ;
        RECT 110.400 343.050 111.450 343.950 ;
        RECT 94.950 341.250 96.750 342.150 ;
        RECT 97.950 340.950 100.050 343.050 ;
        RECT 103.950 340.950 106.050 343.050 ;
        RECT 109.950 340.950 112.050 343.050 ;
        RECT 94.950 339.450 97.050 340.050 ;
        RECT 92.400 338.400 97.050 339.450 ;
        RECT 98.250 338.850 100.050 339.750 ;
        RECT 94.950 337.950 97.050 338.400 ;
        RECT 100.950 338.250 103.050 339.150 ;
        RECT 103.950 338.850 106.050 339.750 ;
        RECT 106.950 338.250 109.050 339.150 ;
        RECT 109.950 338.850 112.050 339.750 ;
        RECT 100.950 336.450 103.050 337.050 ;
        RECT 98.400 335.400 103.050 336.450 ;
        RECT 85.950 331.950 88.050 334.050 ;
        RECT 82.950 328.950 85.050 331.050 ;
        RECT 79.950 322.950 82.050 325.050 ;
        RECT 83.400 312.450 84.450 328.950 ;
        RECT 86.400 328.050 87.450 331.950 ;
        RECT 98.400 331.050 99.450 335.400 ;
        RECT 100.950 334.950 103.050 335.400 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 97.950 328.950 100.050 331.050 ;
        RECT 107.400 328.050 108.450 334.950 ;
        RECT 85.950 325.950 88.050 328.050 ;
        RECT 106.950 325.950 109.050 328.050 ;
        RECT 113.400 322.050 114.450 352.950 ;
        RECT 92.400 320.400 99.450 321.450 ;
        RECT 85.950 316.950 88.050 319.050 ;
        RECT 80.400 311.400 84.450 312.450 ;
        RECT 80.400 310.050 81.450 311.400 ;
        RECT 73.950 308.400 78.450 309.450 ;
        RECT 73.950 307.950 76.050 308.400 ;
        RECT 79.950 307.950 82.050 310.050 ;
        RECT 83.250 308.250 85.050 309.150 ;
        RECT 73.950 305.850 75.750 306.750 ;
        RECT 76.950 304.950 79.050 307.050 ;
        RECT 80.250 305.850 81.750 306.750 ;
        RECT 82.950 304.950 85.050 307.050 ;
        RECT 76.950 302.850 79.050 303.750 ;
        RECT 76.950 298.950 79.050 301.050 ;
        RECT 70.950 274.950 73.050 277.050 ;
        RECT 68.400 272.400 72.450 273.450 ;
        RECT 65.400 271.050 66.450 271.950 ;
        RECT 71.400 271.050 72.450 272.400 ;
        RECT 49.950 269.850 51.750 270.750 ;
        RECT 52.950 268.950 55.050 271.050 ;
        RECT 58.950 268.950 61.050 271.050 ;
        RECT 61.950 269.250 63.750 270.150 ;
        RECT 64.950 268.950 67.050 271.050 ;
        RECT 68.250 269.250 69.750 270.150 ;
        RECT 70.950 268.950 73.050 271.050 ;
        RECT 74.250 269.250 76.050 270.150 ;
        RECT 49.950 265.950 52.050 268.050 ;
        RECT 46.950 256.950 49.050 259.050 ;
        RECT 40.950 241.950 43.050 244.050 ;
        RECT 43.950 241.950 46.050 244.050 ;
        RECT 40.950 236.250 42.750 237.150 ;
        RECT 43.950 235.950 46.050 238.050 ;
        RECT 47.250 236.250 49.050 237.150 ;
        RECT 40.950 234.450 43.050 235.050 ;
        RECT 38.400 233.400 43.050 234.450 ;
        RECT 44.250 233.850 45.750 234.750 ;
        RECT 28.950 230.850 31.050 231.750 ;
        RECT 28.950 217.950 31.050 220.050 ;
        RECT 13.950 205.950 16.050 208.050 ;
        RECT 19.950 205.950 22.050 208.050 ;
        RECT 7.950 199.950 10.050 202.050 ;
        RECT 8.400 199.050 9.450 199.950 ;
        RECT 14.400 199.050 15.450 205.950 ;
        RECT 29.400 205.050 30.450 217.950 ;
        RECT 35.400 208.050 36.450 232.950 ;
        RECT 34.950 205.950 37.050 208.050 ;
        RECT 38.400 205.050 39.450 233.400 ;
        RECT 40.950 232.950 43.050 233.400 ;
        RECT 46.950 232.950 49.050 235.050 ;
        RECT 47.400 232.050 48.450 232.950 ;
        RECT 40.950 229.950 43.050 232.050 ;
        RECT 46.950 229.950 49.050 232.050 ;
        RECT 41.400 205.050 42.450 229.950 ;
        RECT 43.950 214.950 46.050 217.050 ;
        RECT 44.400 205.050 45.450 214.950 ;
        RECT 19.950 203.250 22.050 204.150 ;
        RECT 28.950 202.950 31.050 205.050 ;
        RECT 34.950 203.250 37.050 204.150 ;
        RECT 37.950 202.950 40.050 205.050 ;
        RECT 40.950 202.950 43.050 205.050 ;
        RECT 43.950 202.950 46.050 205.050 ;
        RECT 50.400 204.450 51.450 265.950 ;
        RECT 53.400 265.050 54.450 268.950 ;
        RECT 55.950 265.950 58.050 268.050 ;
        RECT 59.400 267.450 60.450 268.950 ;
        RECT 61.950 267.450 64.050 268.050 ;
        RECT 59.400 266.400 64.050 267.450 ;
        RECT 65.250 266.850 66.750 267.750 ;
        RECT 61.950 265.950 64.050 266.400 ;
        RECT 67.950 265.950 70.050 268.050 ;
        RECT 71.250 266.850 72.750 267.750 ;
        RECT 73.950 265.950 76.050 268.050 ;
        RECT 52.950 262.950 55.050 265.050 ;
        RECT 52.950 247.950 55.050 250.050 ;
        RECT 53.400 214.050 54.450 247.950 ;
        RECT 56.400 241.050 57.450 265.950 ;
        RECT 62.400 262.050 63.450 265.950 ;
        RECT 77.400 262.050 78.450 298.950 ;
        RECT 82.950 286.950 85.050 289.050 ;
        RECT 79.950 269.250 82.050 270.150 ;
        RECT 79.950 267.450 82.050 268.050 ;
        RECT 83.400 267.450 84.450 286.950 ;
        RECT 86.400 280.050 87.450 316.950 ;
        RECT 88.950 307.950 91.050 310.050 ;
        RECT 92.400 307.050 93.450 320.400 ;
        RECT 94.950 316.950 97.050 319.050 ;
        RECT 95.400 310.050 96.450 316.950 ;
        RECT 98.400 313.050 99.450 320.400 ;
        RECT 112.950 319.950 115.050 322.050 ;
        RECT 106.950 316.950 109.050 319.050 ;
        RECT 107.400 316.050 108.450 316.950 ;
        RECT 116.400 316.050 117.450 367.950 ;
        RECT 121.950 358.950 124.050 361.050 ;
        RECT 122.400 346.050 123.450 358.950 ;
        RECT 121.950 343.950 124.050 346.050 ;
        RECT 118.950 341.250 121.050 342.150 ;
        RECT 121.950 341.850 124.050 342.750 ;
        RECT 118.950 337.950 121.050 340.050 ;
        RECT 119.400 319.050 120.450 337.950 ;
        RECT 125.400 337.050 126.450 370.950 ;
        RECT 136.950 367.950 139.050 370.050 ;
        RECT 130.950 358.950 133.050 361.050 ;
        RECT 131.400 346.050 132.450 358.950 ;
        RECT 137.400 346.050 138.450 367.950 ;
        RECT 130.950 343.950 133.050 346.050 ;
        RECT 134.250 344.250 135.750 345.150 ;
        RECT 136.950 343.950 139.050 346.050 ;
        RECT 127.950 341.250 130.050 342.150 ;
        RECT 130.950 341.850 132.750 342.750 ;
        RECT 133.950 340.950 136.050 343.050 ;
        RECT 137.250 341.850 139.050 342.750 ;
        RECT 127.950 337.950 130.050 340.050 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 124.950 331.950 127.050 334.050 ;
        RECT 121.950 328.950 124.050 331.050 ;
        RECT 118.950 316.950 121.050 319.050 ;
        RECT 106.950 313.950 109.050 316.050 ;
        RECT 115.950 313.950 118.050 316.050 ;
        RECT 118.950 313.950 121.050 316.050 ;
        RECT 97.950 310.950 100.050 313.050 ;
        RECT 103.950 311.250 106.050 312.150 ;
        RECT 106.950 311.850 109.050 312.750 ;
        RECT 112.950 312.450 115.050 313.050 ;
        RECT 109.950 311.250 111.750 312.150 ;
        RECT 112.950 311.400 117.450 312.450 ;
        RECT 112.950 310.950 115.050 311.400 ;
        RECT 94.950 307.950 97.050 310.050 ;
        RECT 98.250 308.250 100.050 309.150 ;
        RECT 103.950 307.950 106.050 310.050 ;
        RECT 109.950 307.950 112.050 310.050 ;
        RECT 113.250 308.850 115.050 309.750 ;
        RECT 88.950 305.850 90.750 306.750 ;
        RECT 91.950 304.950 94.050 307.050 ;
        RECT 95.250 305.850 96.750 306.750 ;
        RECT 97.950 304.950 100.050 307.050 ;
        RECT 91.950 302.850 94.050 303.750 ;
        RECT 94.950 301.950 97.050 304.050 ;
        RECT 85.950 277.950 88.050 280.050 ;
        RECT 85.950 271.950 88.050 274.050 ;
        RECT 85.950 269.850 88.050 270.750 ;
        RECT 88.950 269.250 91.050 270.150 ;
        RECT 79.950 266.400 84.450 267.450 ;
        RECT 79.950 265.950 82.050 266.400 ;
        RECT 88.950 265.950 91.050 268.050 ;
        RECT 89.400 265.050 90.450 265.950 ;
        RECT 95.400 265.050 96.450 301.950 ;
        RECT 98.400 298.050 99.450 304.950 ;
        RECT 97.950 295.950 100.050 298.050 ;
        RECT 104.400 295.050 105.450 307.950 ;
        RECT 106.950 304.950 109.050 307.050 ;
        RECT 103.950 292.950 106.050 295.050 ;
        RECT 107.400 286.050 108.450 304.950 ;
        RECT 110.400 301.050 111.450 307.950 ;
        RECT 112.950 304.950 115.050 307.050 ;
        RECT 109.950 298.950 112.050 301.050 ;
        RECT 106.950 283.950 109.050 286.050 ;
        RECT 106.950 274.950 109.050 277.050 ;
        RECT 100.950 271.950 103.050 274.050 ;
        RECT 101.400 271.050 102.450 271.950 ;
        RECT 97.950 269.250 99.750 270.150 ;
        RECT 100.950 268.950 103.050 271.050 ;
        RECT 103.950 269.250 106.050 270.150 ;
        RECT 97.950 265.950 100.050 268.050 ;
        RECT 101.250 266.850 103.050 267.750 ;
        RECT 79.950 262.950 82.050 265.050 ;
        RECT 88.950 262.950 91.050 265.050 ;
        RECT 94.950 262.950 97.050 265.050 ;
        RECT 61.950 259.950 64.050 262.050 ;
        RECT 76.950 259.950 79.050 262.050 ;
        RECT 58.950 256.950 61.050 259.050 ;
        RECT 59.400 241.050 60.450 256.950 ;
        RECT 62.400 247.050 63.450 259.950 ;
        RECT 67.950 253.950 70.050 256.050 ;
        RECT 61.950 244.950 64.050 247.050 ;
        RECT 55.950 238.950 58.050 241.050 ;
        RECT 58.950 238.950 61.050 241.050 ;
        RECT 62.250 239.250 63.750 240.150 ;
        RECT 64.950 238.950 67.050 241.050 ;
        RECT 55.950 235.950 58.050 238.050 ;
        RECT 59.250 236.850 60.750 237.750 ;
        RECT 61.950 235.950 64.050 238.050 ;
        RECT 65.250 236.850 67.050 237.750 ;
        RECT 55.950 233.850 58.050 234.750 ;
        RECT 64.950 232.950 67.050 235.050 ;
        RECT 55.950 214.950 58.050 217.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 52.950 208.950 55.050 211.050 ;
        RECT 53.400 205.050 54.450 208.950 ;
        RECT 47.400 203.400 51.450 204.450 ;
        RECT 16.950 200.250 18.750 201.150 ;
        RECT 19.950 199.950 22.050 202.050 ;
        RECT 23.250 200.250 24.750 201.150 ;
        RECT 25.950 199.950 28.050 202.050 ;
        RECT 31.950 200.250 33.750 201.150 ;
        RECT 34.950 199.950 37.050 202.050 ;
        RECT 40.950 201.450 43.050 202.050 ;
        RECT 38.250 200.250 39.750 201.150 ;
        RECT 40.950 200.400 45.450 201.450 ;
        RECT 40.950 199.950 43.050 200.400 ;
        RECT 4.950 197.250 6.750 198.150 ;
        RECT 7.950 196.950 10.050 199.050 ;
        RECT 13.950 196.950 16.050 199.050 ;
        RECT 16.950 196.950 19.050 199.050 ;
        RECT 4.950 193.950 7.050 196.050 ;
        RECT 8.250 194.850 10.050 195.750 ;
        RECT 10.950 194.250 13.050 195.150 ;
        RECT 13.950 194.850 16.050 195.750 ;
        RECT 1.950 169.950 4.050 172.050 ;
        RECT 5.400 169.050 6.450 193.950 ;
        RECT 20.400 193.050 21.450 199.950 ;
        RECT 22.950 196.950 25.050 199.050 ;
        RECT 26.250 197.850 28.050 198.750 ;
        RECT 31.950 198.450 34.050 199.050 ;
        RECT 29.400 197.400 34.050 198.450 ;
        RECT 23.400 196.050 24.450 196.950 ;
        RECT 22.950 193.950 25.050 196.050 ;
        RECT 25.950 193.950 28.050 196.050 ;
        RECT 10.950 190.950 13.050 193.050 ;
        RECT 19.950 190.950 22.050 193.050 ;
        RECT 7.950 187.950 10.050 190.050 ;
        RECT 8.400 169.050 9.450 187.950 ;
        RECT 22.950 172.950 25.050 175.050 ;
        RECT 13.950 169.950 16.050 172.050 ;
        RECT 16.950 169.950 19.050 172.050 ;
        RECT 14.400 169.050 15.450 169.950 ;
        RECT 17.400 169.050 18.450 169.950 ;
        RECT 23.400 169.050 24.450 172.950 ;
        RECT 26.400 169.050 27.450 193.950 ;
        RECT 1.950 166.950 4.050 169.050 ;
        RECT 4.950 166.950 7.050 169.050 ;
        RECT 7.950 166.950 10.050 169.050 ;
        RECT 11.250 167.250 12.750 168.150 ;
        RECT 13.950 166.950 16.050 169.050 ;
        RECT 16.950 166.950 19.050 169.050 ;
        RECT 20.250 167.250 21.750 168.150 ;
        RECT 22.950 166.950 25.050 169.050 ;
        RECT 25.950 166.950 28.050 169.050 ;
        RECT 2.400 142.050 3.450 166.950 ;
        RECT 4.950 163.950 7.050 166.050 ;
        RECT 8.250 164.850 9.750 165.750 ;
        RECT 10.950 163.950 13.050 166.050 ;
        RECT 14.250 164.850 16.050 165.750 ;
        RECT 16.950 164.850 18.750 165.750 ;
        RECT 19.950 163.950 22.050 166.050 ;
        RECT 23.250 164.850 24.750 165.750 ;
        RECT 25.950 165.450 28.050 166.050 ;
        RECT 29.400 165.450 30.450 197.400 ;
        RECT 31.950 196.950 34.050 197.400 ;
        RECT 31.950 193.950 34.050 196.050 ;
        RECT 32.400 178.050 33.450 193.950 ;
        RECT 31.950 175.950 34.050 178.050 ;
        RECT 35.400 172.050 36.450 199.950 ;
        RECT 37.950 196.950 40.050 199.050 ;
        RECT 41.250 197.850 43.050 198.750 ;
        RECT 34.950 169.950 37.050 172.050 ;
        RECT 31.950 166.950 34.050 169.050 ;
        RECT 32.400 166.050 33.450 166.950 ;
        RECT 25.950 164.400 30.450 165.450 ;
        RECT 25.950 163.950 28.050 164.400 ;
        RECT 4.950 161.850 7.050 162.750 ;
        RECT 13.950 160.950 16.050 163.050 ;
        RECT 25.950 161.850 28.050 162.750 ;
        RECT 1.950 139.950 4.050 142.050 ;
        RECT 10.950 130.950 13.050 133.050 ;
        RECT 11.400 130.050 12.450 130.950 ;
        RECT 4.950 129.450 7.050 130.050 ;
        RECT 2.400 128.400 7.050 129.450 ;
        RECT 2.400 121.050 3.450 128.400 ;
        RECT 4.950 127.950 7.050 128.400 ;
        RECT 8.250 128.250 9.750 129.150 ;
        RECT 10.950 127.950 13.050 130.050 ;
        RECT 4.950 125.850 6.750 126.750 ;
        RECT 7.950 124.950 10.050 127.050 ;
        RECT 11.250 125.850 13.050 126.750 ;
        RECT 8.400 123.450 9.450 124.950 ;
        RECT 5.400 122.400 9.450 123.450 ;
        RECT 1.950 118.950 4.050 121.050 ;
        RECT 5.400 97.050 6.450 122.400 ;
        RECT 14.400 120.450 15.450 160.950 ;
        RECT 29.400 160.050 30.450 164.400 ;
        RECT 31.950 163.950 34.050 166.050 ;
        RECT 35.400 163.050 36.450 169.950 ;
        RECT 38.400 169.050 39.450 196.950 ;
        RECT 44.400 195.450 45.450 200.400 ;
        RECT 41.400 194.400 45.450 195.450 ;
        RECT 41.400 184.050 42.450 194.400 ;
        RECT 47.400 193.050 48.450 203.400 ;
        RECT 52.950 202.950 55.050 205.050 ;
        RECT 56.400 202.050 57.450 214.950 ;
        RECT 61.950 211.950 64.050 214.050 ;
        RECT 62.400 202.050 63.450 211.950 ;
        RECT 65.400 211.050 66.450 232.950 ;
        RECT 68.400 220.050 69.450 253.950 ;
        RECT 73.950 244.950 76.050 247.050 ;
        RECT 70.950 241.950 73.050 244.050 ;
        RECT 71.400 241.050 72.450 241.950 ;
        RECT 70.950 238.950 73.050 241.050 ;
        RECT 70.950 236.850 73.050 237.750 ;
        RECT 70.950 223.950 73.050 226.050 ;
        RECT 67.950 217.950 70.050 220.050 ;
        RECT 64.950 208.950 67.050 211.050 ;
        RECT 71.400 205.050 72.450 223.950 ;
        RECT 70.950 202.950 73.050 205.050 ;
        RECT 53.250 200.250 54.750 201.150 ;
        RECT 55.950 199.950 58.050 202.050 ;
        RECT 61.950 199.950 64.050 202.050 ;
        RECT 74.400 201.450 75.450 244.950 ;
        RECT 80.400 244.050 81.450 262.950 ;
        RECT 98.400 262.050 99.450 265.950 ;
        RECT 97.950 259.950 100.050 262.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 94.950 247.950 97.050 250.050 ;
        RECT 85.950 244.950 88.050 247.050 ;
        RECT 88.950 244.950 91.050 247.050 ;
        RECT 86.400 244.050 87.450 244.950 ;
        RECT 79.950 241.950 82.050 244.050 ;
        RECT 85.950 241.950 88.050 244.050 ;
        RECT 82.950 239.250 85.050 240.150 ;
        RECT 85.950 239.850 88.050 240.750 ;
        RECT 89.400 238.050 90.450 244.950 ;
        RECT 95.400 244.050 96.450 247.950 ;
        RECT 94.950 241.950 97.050 244.050 ;
        RECT 95.400 238.050 96.450 241.950 ;
        RECT 98.400 241.050 99.450 256.950 ;
        RECT 107.400 247.050 108.450 274.950 ;
        RECT 110.400 274.050 111.450 298.950 ;
        RECT 109.950 271.950 112.050 274.050 ;
        RECT 109.950 269.250 112.050 270.150 ;
        RECT 109.950 265.950 112.050 268.050 ;
        RECT 113.400 262.050 114.450 304.950 ;
        RECT 116.400 301.050 117.450 311.400 ;
        RECT 119.400 304.050 120.450 313.950 ;
        RECT 122.400 313.050 123.450 328.950 ;
        RECT 125.400 313.050 126.450 331.950 ;
        RECT 134.400 325.050 135.450 340.950 ;
        RECT 136.950 337.950 139.050 340.050 ;
        RECT 137.400 331.050 138.450 337.950 ;
        RECT 140.400 334.050 141.450 373.950 ;
        RECT 143.400 373.050 144.450 376.950 ;
        RECT 146.400 376.050 147.450 379.950 ;
        RECT 148.950 376.950 151.050 379.050 ;
        RECT 151.950 376.950 154.050 379.050 ;
        RECT 155.250 377.850 156.750 378.750 ;
        RECT 157.950 376.950 160.050 379.050 ;
        RECT 160.950 376.950 163.050 379.050 ;
        RECT 166.950 376.950 169.050 379.050 ;
        RECT 170.250 377.850 171.750 378.750 ;
        RECT 172.950 376.950 175.050 379.050 ;
        RECT 176.250 377.850 178.050 378.750 ;
        RECT 178.950 376.950 181.050 379.050 ;
        RECT 145.950 373.950 148.050 376.050 ;
        RECT 142.950 370.950 145.050 373.050 ;
        RECT 145.950 364.950 148.050 367.050 ;
        RECT 142.950 349.950 145.050 352.050 ;
        RECT 143.400 346.050 144.450 349.950 ;
        RECT 142.950 343.950 145.050 346.050 ;
        RECT 142.950 341.250 145.050 342.150 ;
        RECT 142.950 337.950 145.050 340.050 ;
        RECT 146.400 337.050 147.450 364.950 ;
        RECT 149.400 358.050 150.450 376.950 ;
        RECT 152.400 373.050 153.450 376.950 ;
        RECT 151.950 370.950 154.050 373.050 ;
        RECT 154.950 358.950 157.050 361.050 ;
        RECT 148.950 355.950 151.050 358.050 ;
        RECT 155.400 343.050 156.450 358.950 ;
        RECT 148.950 341.850 151.050 342.750 ;
        RECT 151.950 341.250 154.050 342.150 ;
        RECT 154.950 340.950 157.050 343.050 ;
        RECT 158.400 340.050 159.450 376.950 ;
        RECT 161.400 367.050 162.450 376.950 ;
        RECT 167.400 370.050 168.450 376.950 ;
        RECT 169.950 373.950 172.050 376.050 ;
        RECT 172.950 374.850 175.050 375.750 ;
        RECT 166.950 367.950 169.050 370.050 ;
        RECT 160.950 364.950 163.050 367.050 ;
        RECT 170.400 349.050 171.450 373.950 ;
        RECT 172.950 355.950 175.050 358.050 ;
        RECT 166.950 346.950 169.050 349.050 ;
        RECT 169.950 346.950 172.050 349.050 ;
        RECT 160.950 344.250 163.050 345.150 ;
        RECT 167.400 343.050 168.450 346.950 ;
        RECT 160.950 340.950 163.050 343.050 ;
        RECT 164.250 341.250 165.750 342.150 ;
        RECT 166.950 340.950 169.050 343.050 ;
        RECT 170.250 341.250 172.050 342.150 ;
        RECT 161.400 340.050 162.450 340.950 ;
        RECT 151.950 337.950 154.050 340.050 ;
        RECT 157.950 337.950 160.050 340.050 ;
        RECT 160.950 337.950 163.050 340.050 ;
        RECT 163.950 337.950 166.050 340.050 ;
        RECT 167.250 338.850 168.750 339.750 ;
        RECT 169.950 339.450 172.050 340.050 ;
        RECT 173.400 339.450 174.450 355.950 ;
        RECT 179.400 352.050 180.450 376.950 ;
        RECT 188.400 361.050 189.450 403.950 ;
        RECT 190.950 403.500 193.050 405.600 ;
        RECT 200.400 400.050 201.450 409.950 ;
        RECT 199.950 397.950 202.050 400.050 ;
        RECT 193.950 391.950 196.050 394.050 ;
        RECT 194.400 385.050 195.450 391.950 ;
        RECT 199.950 388.950 202.050 391.050 ;
        RECT 200.400 385.050 201.450 388.950 ;
        RECT 203.400 385.050 204.450 412.950 ;
        RECT 205.950 409.950 208.050 412.050 ;
        RECT 212.400 405.600 213.600 422.400 ;
        RECT 211.950 403.500 214.050 405.600 ;
        RECT 215.400 388.050 216.450 446.400 ;
        RECT 224.400 439.050 225.450 448.950 ;
        RECT 217.950 436.950 220.050 439.050 ;
        RECT 223.950 436.950 226.050 439.050 ;
        RECT 218.400 415.050 219.450 436.950 ;
        RECT 233.400 430.050 234.450 448.950 ;
        RECT 239.400 445.050 240.450 467.400 ;
        RECT 242.400 457.050 243.450 472.950 ;
        RECT 241.950 454.950 244.050 457.050 ;
        RECT 241.950 452.850 244.050 453.750 ;
        RECT 238.950 442.950 241.050 445.050 ;
        RECT 232.950 427.950 235.050 430.050 ;
        RECT 217.950 412.950 220.050 415.050 ;
        RECT 223.950 413.250 226.050 414.150 ;
        RECT 229.950 413.250 232.050 414.150 ;
        RECT 218.400 388.050 219.450 412.950 ;
        RECT 223.950 409.950 226.050 412.050 ;
        RECT 229.950 411.450 232.050 412.050 ;
        RECT 233.400 411.450 234.450 427.950 ;
        RECT 238.950 422.400 241.050 424.500 ;
        RECT 229.950 410.400 234.450 411.450 ;
        RECT 229.950 409.950 232.050 410.400 ;
        RECT 224.400 391.050 225.450 409.950 ;
        RECT 239.400 405.600 240.600 422.400 ;
        RECT 245.400 418.050 246.450 482.400 ;
        RECT 247.950 481.950 250.050 482.400 ;
        RECT 253.950 481.950 256.050 484.050 ;
        RECT 256.950 481.950 259.050 484.050 ;
        RECT 257.400 481.050 258.450 481.950 ;
        RECT 256.950 478.950 259.050 481.050 ;
        RECT 253.950 472.950 256.050 475.050 ;
        RECT 247.950 463.950 250.050 466.050 ;
        RECT 248.400 457.050 249.450 463.950 ;
        RECT 254.400 457.050 255.450 472.950 ;
        RECT 260.400 472.050 261.450 502.950 ;
        RECT 259.950 469.950 262.050 472.050 ;
        RECT 259.950 466.950 262.050 469.050 ;
        RECT 256.950 460.950 259.050 463.050 ;
        RECT 247.950 454.950 250.050 457.050 ;
        RECT 251.250 455.250 252.750 456.150 ;
        RECT 253.950 454.950 256.050 457.050 ;
        RECT 257.400 454.050 258.450 460.950 ;
        RECT 247.950 452.850 249.750 453.750 ;
        RECT 250.950 451.950 253.050 454.050 ;
        RECT 254.250 452.850 255.750 453.750 ;
        RECT 256.950 451.950 259.050 454.050 ;
        RECT 247.950 445.950 250.050 448.050 ;
        RECT 244.950 415.950 247.050 418.050 ;
        RECT 244.950 413.250 247.050 414.150 ;
        RECT 244.950 409.950 247.050 412.050 ;
        RECT 245.400 406.050 246.450 409.950 ;
        RECT 238.950 403.500 241.050 405.600 ;
        RECT 244.950 403.950 247.050 406.050 ;
        RECT 248.400 400.050 249.450 445.950 ;
        RECT 251.400 433.050 252.450 451.950 ;
        RECT 253.950 448.950 256.050 451.050 ;
        RECT 256.950 449.850 259.050 450.750 ;
        RECT 254.400 439.050 255.450 448.950 ;
        RECT 260.400 447.450 261.450 466.950 ;
        RECT 263.400 466.050 264.450 517.950 ;
        RECT 266.400 511.050 267.450 520.950 ;
        RECT 272.400 520.050 273.450 523.950 ;
        RECT 277.950 521.850 280.050 522.750 ;
        RECT 271.950 517.950 274.050 520.050 ;
        RECT 277.950 514.950 280.050 517.050 ;
        RECT 265.950 508.950 268.050 511.050 ;
        RECT 271.950 490.950 274.050 493.050 ;
        RECT 265.950 488.250 268.050 489.150 ;
        RECT 272.400 487.050 273.450 490.950 ;
        RECT 278.400 490.050 279.450 514.950 ;
        RECT 281.400 513.450 282.450 550.950 ;
        RECT 286.950 544.950 289.050 547.050 ;
        RECT 287.400 529.050 288.450 544.950 ;
        RECT 289.950 541.950 292.050 544.050 ;
        RECT 283.950 527.250 285.750 528.150 ;
        RECT 286.950 526.950 289.050 529.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 287.250 524.850 289.050 525.750 ;
        RECT 284.400 523.050 285.450 523.950 ;
        RECT 283.950 520.950 286.050 523.050 ;
        RECT 286.950 520.950 289.050 523.050 ;
        RECT 284.400 517.050 285.450 520.950 ;
        RECT 283.950 514.950 286.050 517.050 ;
        RECT 281.400 512.400 285.450 513.450 ;
        RECT 284.400 493.050 285.450 512.400 ;
        RECT 283.950 490.950 286.050 493.050 ;
        RECT 277.950 487.950 280.050 490.050 ;
        RECT 281.250 488.250 282.750 489.150 ;
        RECT 265.950 484.950 268.050 487.050 ;
        RECT 269.250 485.250 270.750 486.150 ;
        RECT 271.950 484.950 274.050 487.050 ;
        RECT 275.250 485.250 277.050 486.150 ;
        RECT 277.950 485.850 279.750 486.750 ;
        RECT 280.950 484.950 283.050 487.050 ;
        RECT 284.250 485.850 286.050 486.750 ;
        RECT 266.400 475.050 267.450 484.950 ;
        RECT 281.400 484.050 282.450 484.950 ;
        RECT 268.950 481.950 271.050 484.050 ;
        RECT 272.250 482.850 273.750 483.750 ;
        RECT 274.950 481.950 277.050 484.050 ;
        RECT 280.950 481.950 283.050 484.050 ;
        RECT 281.400 481.050 282.450 481.950 ;
        RECT 274.950 478.950 277.050 481.050 ;
        RECT 280.950 478.950 283.050 481.050 ;
        RECT 265.950 472.950 268.050 475.050 ;
        RECT 268.950 472.950 271.050 475.050 ;
        RECT 262.950 463.950 265.050 466.050 ;
        RECT 269.400 457.050 270.450 472.950 ;
        RECT 271.950 469.950 274.050 472.050 ;
        RECT 272.400 457.050 273.450 469.950 ;
        RECT 262.950 454.950 265.050 457.050 ;
        RECT 266.250 455.250 267.750 456.150 ;
        RECT 268.950 454.950 271.050 457.050 ;
        RECT 271.950 454.950 274.050 457.050 ;
        RECT 262.950 452.850 264.750 453.750 ;
        RECT 265.950 451.950 268.050 454.050 ;
        RECT 269.250 452.850 270.750 453.750 ;
        RECT 271.950 451.950 274.050 454.050 ;
        RECT 275.400 451.050 276.450 478.950 ;
        RECT 287.400 472.050 288.450 520.950 ;
        RECT 290.400 505.050 291.450 541.950 ;
        RECT 293.400 523.050 294.450 550.950 ;
        RECT 298.950 538.950 301.050 541.050 ;
        RECT 299.400 526.050 300.450 538.950 ;
        RECT 305.400 528.450 306.450 554.400 ;
        RECT 311.400 552.450 312.450 593.400 ;
        RECT 328.950 592.950 331.050 593.400 ;
        RECT 334.950 593.400 339.450 594.450 ;
        RECT 340.950 593.850 342.750 594.750 ;
        RECT 334.950 592.950 337.050 593.400 ;
        RECT 343.950 592.950 346.050 595.050 ;
        RECT 347.250 593.850 348.750 594.750 ;
        RECT 349.950 592.950 352.050 595.050 ;
        RECT 343.950 590.850 346.050 591.750 ;
        RECT 350.400 564.450 351.450 592.950 ;
        RECT 347.400 563.400 351.450 564.450 ;
        RECT 322.950 559.950 325.050 562.050 ;
        RECT 313.950 557.250 316.050 558.150 ;
        RECT 319.950 557.250 322.050 558.150 ;
        RECT 313.950 555.450 316.050 556.050 ;
        RECT 313.950 554.400 318.450 555.450 ;
        RECT 313.950 553.950 316.050 554.400 ;
        RECT 311.400 551.400 315.450 552.450 ;
        RECT 307.950 528.450 310.050 529.050 ;
        RECT 305.400 527.400 310.050 528.450 ;
        RECT 295.950 524.250 297.750 525.150 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 302.250 524.250 304.050 525.150 ;
        RECT 292.950 520.950 295.050 523.050 ;
        RECT 295.950 520.950 298.050 523.050 ;
        RECT 299.250 521.850 300.750 522.750 ;
        RECT 301.950 522.450 304.050 523.050 ;
        RECT 305.400 522.450 306.450 527.400 ;
        RECT 307.950 526.950 310.050 527.400 ;
        RECT 307.950 524.850 310.050 525.750 ;
        RECT 310.950 524.250 313.050 525.150 ;
        RECT 301.950 521.400 306.450 522.450 ;
        RECT 301.950 520.950 304.050 521.400 ;
        RECT 310.950 520.950 313.050 523.050 ;
        RECT 301.950 517.950 304.050 520.050 ;
        RECT 289.950 502.950 292.050 505.050 ;
        RECT 292.950 490.950 295.050 493.050 ;
        RECT 293.400 487.050 294.450 490.950 ;
        RECT 298.950 488.250 301.050 489.150 ;
        RECT 289.950 485.250 291.750 486.150 ;
        RECT 292.950 484.950 295.050 487.050 ;
        RECT 296.250 485.250 297.750 486.150 ;
        RECT 298.950 484.950 301.050 487.050 ;
        RECT 289.950 481.950 292.050 484.050 ;
        RECT 293.250 482.850 294.750 483.750 ;
        RECT 295.950 481.950 298.050 484.050 ;
        RECT 289.950 478.950 292.050 481.050 ;
        RECT 286.950 469.950 289.050 472.050 ;
        RECT 277.950 463.950 280.050 466.050 ;
        RECT 280.950 463.950 283.050 466.050 ;
        RECT 278.400 457.050 279.450 463.950 ;
        RECT 281.400 460.050 282.450 463.950 ;
        RECT 290.400 460.050 291.450 478.950 ;
        RECT 296.400 472.050 297.450 481.950 ;
        RECT 299.400 478.050 300.450 484.950 ;
        RECT 298.950 475.950 301.050 478.050 ;
        RECT 302.400 474.450 303.450 517.950 ;
        RECT 304.950 490.950 307.050 493.050 ;
        RECT 305.400 486.450 306.450 490.950 ;
        RECT 311.400 490.050 312.450 520.950 ;
        RECT 314.400 520.050 315.450 551.400 ;
        RECT 317.400 532.050 318.450 554.400 ;
        RECT 323.400 541.050 324.450 559.950 ;
        RECT 347.400 559.050 348.450 563.400 ;
        RECT 328.950 558.450 331.050 559.050 ;
        RECT 326.400 557.400 331.050 558.450 ;
        RECT 322.950 538.950 325.050 541.050 ;
        RECT 326.400 538.050 327.450 557.400 ;
        RECT 328.950 556.950 331.050 557.400 ;
        RECT 346.950 556.950 349.050 559.050 ;
        RECT 328.950 554.850 331.050 555.750 ;
        RECT 349.950 554.850 352.050 555.750 ;
        RECT 346.950 538.950 349.050 541.050 ;
        RECT 325.950 535.950 328.050 538.050 ;
        RECT 326.400 535.050 327.450 535.950 ;
        RECT 325.950 532.950 328.050 535.050 ;
        RECT 343.950 532.950 346.050 535.050 ;
        RECT 316.950 529.950 319.050 532.050 ;
        RECT 316.950 526.950 319.050 529.050 ;
        RECT 322.950 526.950 325.050 529.050 ;
        RECT 334.950 526.950 337.050 529.050 ;
        RECT 323.400 526.050 324.450 526.950 ;
        RECT 316.950 524.850 319.050 525.750 ;
        RECT 319.950 524.250 321.750 525.150 ;
        RECT 322.950 523.950 325.050 526.050 ;
        RECT 331.950 525.450 334.050 526.050 ;
        RECT 326.250 524.250 328.050 525.150 ;
        RECT 329.400 524.400 334.050 525.450 ;
        RECT 316.950 520.950 319.050 523.050 ;
        RECT 319.950 520.950 322.050 523.050 ;
        RECT 323.250 521.850 324.750 522.750 ;
        RECT 325.950 522.450 328.050 523.050 ;
        RECT 329.400 522.450 330.450 524.400 ;
        RECT 331.950 523.950 334.050 524.400 ;
        RECT 335.400 523.050 336.450 526.950 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 341.250 524.250 343.050 525.150 ;
        RECT 325.950 521.400 330.450 522.450 ;
        RECT 331.950 521.850 333.750 522.750 ;
        RECT 325.950 520.950 328.050 521.400 ;
        RECT 334.950 520.950 337.050 523.050 ;
        RECT 338.250 521.850 339.750 522.750 ;
        RECT 340.950 520.950 343.050 523.050 ;
        RECT 313.950 517.950 316.050 520.050 ;
        RECT 313.950 511.950 316.050 514.050 ;
        RECT 307.950 488.250 310.050 489.150 ;
        RECT 310.950 487.950 313.050 490.050 ;
        RECT 314.400 487.050 315.450 511.950 ;
        RECT 317.400 490.050 318.450 520.950 ;
        RECT 320.400 519.450 321.450 520.950 ;
        RECT 320.400 518.400 324.450 519.450 ;
        RECT 323.400 502.050 324.450 518.400 ;
        RECT 322.950 499.950 325.050 502.050 ;
        RECT 319.950 496.950 322.050 499.050 ;
        RECT 316.950 487.950 319.050 490.050 ;
        RECT 320.400 487.050 321.450 496.950 ;
        RECT 323.400 487.050 324.450 499.950 ;
        RECT 307.950 486.450 310.050 487.050 ;
        RECT 305.400 485.400 310.050 486.450 ;
        RECT 307.950 484.950 310.050 485.400 ;
        RECT 311.250 485.250 312.750 486.150 ;
        RECT 313.950 484.950 316.050 487.050 ;
        RECT 317.250 485.250 319.050 486.150 ;
        RECT 319.950 484.950 322.050 487.050 ;
        RECT 322.950 484.950 325.050 487.050 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 314.250 482.850 315.750 483.750 ;
        RECT 316.950 481.950 319.050 484.050 ;
        RECT 319.950 482.250 322.050 483.150 ;
        RECT 322.950 482.850 325.050 483.750 ;
        RECT 310.950 478.950 313.050 481.050 ;
        RECT 299.400 473.400 303.450 474.450 ;
        RECT 295.950 469.950 298.050 472.050 ;
        RECT 292.950 466.950 295.050 469.050 ;
        RECT 293.400 460.050 294.450 466.950 ;
        RECT 280.950 457.950 283.050 460.050 ;
        RECT 289.950 457.950 292.050 460.050 ;
        RECT 292.950 457.950 295.050 460.050 ;
        RECT 299.400 457.050 300.450 473.400 ;
        RECT 304.950 463.950 307.050 466.050 ;
        RECT 305.400 460.050 306.450 463.950 ;
        RECT 304.950 457.950 307.050 460.050 ;
        RECT 277.950 454.950 280.050 457.050 ;
        RECT 281.250 455.850 282.750 456.750 ;
        RECT 283.950 454.950 286.050 457.050 ;
        RECT 289.950 455.250 292.050 456.150 ;
        RECT 292.950 455.850 295.050 456.750 ;
        RECT 295.950 455.250 297.750 456.150 ;
        RECT 298.950 454.950 301.050 457.050 ;
        RECT 304.950 455.850 307.050 456.750 ;
        RECT 307.950 455.250 310.050 456.150 ;
        RECT 311.400 454.050 312.450 478.950 ;
        RECT 313.950 460.950 316.050 463.050 ;
        RECT 314.400 457.050 315.450 460.950 ;
        RECT 317.400 460.050 318.450 481.950 ;
        RECT 319.950 478.950 322.050 481.050 ;
        RECT 320.400 463.050 321.450 478.950 ;
        RECT 322.950 466.950 325.050 469.050 ;
        RECT 319.950 460.950 322.050 463.050 ;
        RECT 316.950 457.950 319.050 460.050 ;
        RECT 313.950 454.950 316.050 457.050 ;
        RECT 317.250 455.250 318.750 456.150 ;
        RECT 319.950 454.950 322.050 457.050 ;
        RECT 323.400 454.050 324.450 466.950 ;
        RECT 326.400 466.050 327.450 520.950 ;
        RECT 334.950 518.850 337.050 519.750 ;
        RECT 341.400 496.050 342.450 520.950 ;
        RECT 340.950 493.950 343.050 496.050 ;
        RECT 340.950 490.950 343.050 493.050 ;
        RECT 337.950 488.250 340.050 489.150 ;
        RECT 328.950 485.250 330.750 486.150 ;
        RECT 331.950 484.950 334.050 487.050 ;
        RECT 335.250 485.250 336.750 486.150 ;
        RECT 337.950 484.950 340.050 487.050 ;
        RECT 341.400 484.050 342.450 490.950 ;
        RECT 344.400 490.050 345.450 532.950 ;
        RECT 347.400 532.050 348.450 538.950 ;
        RECT 346.950 529.950 349.050 532.050 ;
        RECT 346.950 527.850 349.050 528.750 ;
        RECT 349.950 527.250 352.050 528.150 ;
        RECT 349.950 523.950 352.050 526.050 ;
        RECT 353.400 505.050 354.450 598.950 ;
        RECT 355.950 596.850 358.050 597.750 ;
        RECT 359.400 552.450 360.450 599.400 ;
        RECT 361.950 596.850 364.050 597.750 ;
        RECT 361.950 566.400 364.050 568.500 ;
        RECT 356.400 551.400 360.450 552.450 ;
        RECT 356.400 544.050 357.450 551.400 ;
        RECT 358.950 547.950 361.050 550.050 ;
        RECT 362.400 549.600 363.600 566.400 ;
        RECT 355.950 541.950 358.050 544.050 ;
        RECT 355.950 529.950 358.050 532.050 ;
        RECT 359.400 531.450 360.450 547.950 ;
        RECT 361.950 547.500 364.050 549.600 ;
        RECT 365.400 535.050 366.450 601.950 ;
        RECT 370.950 599.250 373.050 600.150 ;
        RECT 391.950 599.250 394.050 600.150 ;
        RECT 391.950 595.950 394.050 598.050 ;
        RECT 382.950 567.300 385.050 569.400 ;
        RECT 383.250 563.700 384.450 567.300 ;
        RECT 382.950 561.600 385.050 563.700 ;
        RECT 367.950 557.250 370.050 558.150 ;
        RECT 373.950 557.250 376.050 558.150 ;
        RECT 367.950 553.950 370.050 556.050 ;
        RECT 373.950 553.950 376.050 556.050 ;
        RECT 379.950 553.950 382.050 556.050 ;
        RECT 368.400 553.050 369.450 553.950 ;
        RECT 367.950 550.950 370.050 553.050 ;
        RECT 373.950 535.950 376.050 538.050 ;
        RECT 364.950 532.950 367.050 535.050 ;
        RECT 370.950 533.400 373.050 535.500 ;
        RECT 359.400 530.400 363.450 531.450 ;
        RECT 355.950 527.850 358.050 528.750 ;
        RECT 358.950 527.250 361.050 528.150 ;
        RECT 358.950 523.950 361.050 526.050 ;
        RECT 352.950 502.950 355.050 505.050 ;
        RECT 349.950 493.950 352.050 496.050 ;
        RECT 358.950 493.950 361.050 496.050 ;
        RECT 343.950 487.950 346.050 490.050 ;
        RECT 350.400 487.050 351.450 493.950 ;
        RECT 352.950 490.950 355.050 493.050 ;
        RECT 353.400 490.050 354.450 490.950 ;
        RECT 359.400 490.050 360.450 493.950 ;
        RECT 352.950 487.950 355.050 490.050 ;
        RECT 356.250 488.250 357.750 489.150 ;
        RECT 358.950 487.950 361.050 490.050 ;
        RECT 346.950 486.450 349.050 487.050 ;
        RECT 344.400 485.400 349.050 486.450 ;
        RECT 328.950 481.950 331.050 484.050 ;
        RECT 332.250 482.850 333.750 483.750 ;
        RECT 334.950 481.950 337.050 484.050 ;
        RECT 340.950 481.950 343.050 484.050 ;
        RECT 325.950 463.950 328.050 466.050 ;
        RECT 340.950 460.950 343.050 463.050 ;
        RECT 331.950 459.450 334.050 460.050 ;
        RECT 331.950 458.400 339.450 459.450 ;
        RECT 331.950 457.950 334.050 458.400 ;
        RECT 328.950 454.950 331.050 457.050 ;
        RECT 332.250 455.850 333.750 456.750 ;
        RECT 334.950 454.950 337.050 457.050 ;
        RECT 277.950 452.850 280.050 453.750 ;
        RECT 280.950 451.950 283.050 454.050 ;
        RECT 283.950 452.850 286.050 453.750 ;
        RECT 289.950 451.950 292.050 454.050 ;
        RECT 295.950 451.950 298.050 454.050 ;
        RECT 299.250 452.850 301.050 453.750 ;
        RECT 307.950 451.950 310.050 454.050 ;
        RECT 310.950 451.950 313.050 454.050 ;
        RECT 313.950 452.850 315.750 453.750 ;
        RECT 316.950 451.950 319.050 454.050 ;
        RECT 320.250 452.850 321.750 453.750 ;
        RECT 322.950 451.950 325.050 454.050 ;
        RECT 328.950 452.850 331.050 453.750 ;
        RECT 331.950 451.950 334.050 454.050 ;
        RECT 334.950 452.850 337.050 453.750 ;
        RECT 268.950 448.950 271.050 451.050 ;
        RECT 271.950 449.850 274.050 450.750 ;
        RECT 274.950 448.950 277.050 451.050 ;
        RECT 257.400 446.400 261.450 447.450 ;
        RECT 253.950 436.950 256.050 439.050 ;
        RECT 253.950 433.950 256.050 436.050 ;
        RECT 250.950 430.950 253.050 433.050 ;
        RECT 254.400 424.050 255.450 433.950 ;
        RECT 253.950 421.950 256.050 424.050 ;
        RECT 250.950 413.250 253.050 414.150 ;
        RECT 250.950 411.450 253.050 412.050 ;
        RECT 254.400 411.450 255.450 421.950 ;
        RECT 250.950 410.400 255.450 411.450 ;
        RECT 250.950 409.950 253.050 410.400 ;
        RECT 254.400 403.050 255.450 410.400 ;
        RECT 253.950 400.950 256.050 403.050 ;
        RECT 247.950 397.950 250.050 400.050 ;
        RECT 250.950 394.950 253.050 397.050 ;
        RECT 247.950 391.950 250.050 394.050 ;
        RECT 223.950 388.950 226.050 391.050 ;
        RECT 238.950 388.950 241.050 391.050 ;
        RECT 241.950 389.400 244.050 391.500 ;
        RECT 205.950 385.950 208.050 388.050 ;
        RECT 214.950 385.950 217.050 388.050 ;
        RECT 217.950 385.950 220.050 388.050 ;
        RECT 223.950 385.950 226.050 388.050 ;
        RECT 190.950 382.950 193.050 385.050 ;
        RECT 193.950 382.950 196.050 385.050 ;
        RECT 197.250 383.250 198.750 384.150 ;
        RECT 199.950 382.950 202.050 385.050 ;
        RECT 202.950 382.950 205.050 385.050 ;
        RECT 191.400 382.050 192.450 382.950 ;
        RECT 206.400 382.050 207.450 385.950 ;
        RECT 218.400 385.050 219.450 385.950 ;
        RECT 214.950 383.250 216.750 384.150 ;
        RECT 217.950 382.950 220.050 385.050 ;
        RECT 190.950 379.950 193.050 382.050 ;
        RECT 194.250 380.850 195.750 381.750 ;
        RECT 196.950 379.950 199.050 382.050 ;
        RECT 200.250 380.850 202.050 381.750 ;
        RECT 202.950 380.250 204.750 381.150 ;
        RECT 205.950 379.950 208.050 382.050 ;
        RECT 209.250 380.250 211.050 381.150 ;
        RECT 214.950 379.950 217.050 382.050 ;
        RECT 218.250 380.850 220.050 381.750 ;
        RECT 224.400 381.450 225.450 385.950 ;
        RECT 221.400 380.400 225.450 381.450 ;
        RECT 190.950 377.850 193.050 378.750 ;
        RECT 190.950 373.950 193.050 376.050 ;
        RECT 187.950 358.950 190.050 361.050 ;
        RECT 178.950 349.950 181.050 352.050 ;
        RECT 175.950 344.250 178.050 345.150 ;
        RECT 175.950 340.950 178.050 343.050 ;
        RECT 179.250 341.250 180.750 342.150 ;
        RECT 181.950 340.950 184.050 343.050 ;
        RECT 185.250 341.250 187.050 342.150 ;
        RECT 169.950 338.400 174.450 339.450 ;
        RECT 169.950 337.950 172.050 338.400 ;
        RECT 175.950 337.950 178.050 340.050 ;
        RECT 178.950 337.950 181.050 340.050 ;
        RECT 182.250 338.850 183.750 339.750 ;
        RECT 184.950 337.950 187.050 340.050 ;
        RECT 164.400 337.050 165.450 337.950 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 145.950 334.950 148.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 139.950 331.950 142.050 334.050 ;
        RECT 136.950 328.950 139.050 331.050 ;
        RECT 133.950 322.950 136.050 325.050 ;
        RECT 139.950 316.950 142.050 319.050 ;
        RECT 133.950 313.950 136.050 316.050 ;
        RECT 121.950 310.950 124.050 313.050 ;
        RECT 124.950 310.950 127.050 313.050 ;
        RECT 130.950 312.450 133.050 313.050 ;
        RECT 134.400 312.450 135.450 313.950 ;
        RECT 140.400 313.050 141.450 316.950 ;
        RECT 143.400 313.050 144.450 334.950 ;
        RECT 170.400 334.050 171.450 337.950 ;
        RECT 145.950 331.950 148.050 334.050 ;
        RECT 169.950 331.950 172.050 334.050 ;
        RECT 128.250 311.250 129.750 312.150 ;
        RECT 130.950 311.400 135.450 312.450 ;
        RECT 130.950 310.950 133.050 311.400 ;
        RECT 134.400 310.050 135.450 311.400 ;
        RECT 139.950 310.950 142.050 313.050 ;
        RECT 142.950 310.950 145.050 313.050 ;
        RECT 140.400 310.050 141.450 310.950 ;
        RECT 121.950 307.950 124.050 310.050 ;
        RECT 125.250 308.850 126.750 309.750 ;
        RECT 127.950 307.950 130.050 310.050 ;
        RECT 131.250 308.850 133.050 309.750 ;
        RECT 133.950 307.950 136.050 310.050 ;
        RECT 136.950 307.950 139.050 310.050 ;
        RECT 139.950 307.950 142.050 310.050 ;
        RECT 143.250 308.250 145.050 309.150 ;
        RECT 121.950 305.850 124.050 306.750 ;
        RECT 118.950 301.950 121.050 304.050 ;
        RECT 128.400 301.050 129.450 307.950 ;
        RECT 137.400 307.050 138.450 307.950 ;
        RECT 130.950 304.950 133.050 307.050 ;
        RECT 133.950 305.850 135.750 306.750 ;
        RECT 136.950 304.950 139.050 307.050 ;
        RECT 140.250 305.850 141.750 306.750 ;
        RECT 142.950 304.950 145.050 307.050 ;
        RECT 115.950 298.950 118.050 301.050 ;
        RECT 127.950 298.950 130.050 301.050 ;
        RECT 127.950 292.950 130.050 295.050 ;
        RECT 124.950 280.950 127.050 283.050 ;
        RECT 121.950 277.950 124.050 280.050 ;
        RECT 122.400 274.050 123.450 277.950 ;
        RECT 118.950 272.250 121.050 273.150 ;
        RECT 121.950 271.950 124.050 274.050 ;
        RECT 125.400 271.050 126.450 280.950 ;
        RECT 128.400 277.050 129.450 292.950 ;
        RECT 131.400 280.050 132.450 304.950 ;
        RECT 133.950 301.950 136.050 304.050 ;
        RECT 136.950 302.850 139.050 303.750 ;
        RECT 139.950 301.950 142.050 304.050 ;
        RECT 134.400 298.050 135.450 301.950 ;
        RECT 133.950 295.950 136.050 298.050 ;
        RECT 133.950 280.950 136.050 283.050 ;
        RECT 130.950 277.950 133.050 280.050 ;
        RECT 127.950 274.950 130.050 277.050 ;
        RECT 134.400 271.050 135.450 280.950 ;
        RECT 140.400 279.450 141.450 301.950 ;
        RECT 143.400 283.050 144.450 304.950 ;
        RECT 146.400 301.050 147.450 331.950 ;
        RECT 154.950 316.950 157.050 319.050 ;
        RECT 151.950 313.950 154.050 316.050 ;
        RECT 148.950 310.950 151.050 313.050 ;
        RECT 149.400 310.050 150.450 310.950 ;
        RECT 152.400 310.050 153.450 313.950 ;
        RECT 155.400 310.050 156.450 316.950 ;
        RECT 166.950 313.950 169.050 316.050 ;
        RECT 167.400 313.050 168.450 313.950 ;
        RECT 160.950 310.950 163.050 313.050 ;
        RECT 166.950 310.950 169.050 313.050 ;
        RECT 148.950 307.950 151.050 310.050 ;
        RECT 151.950 307.950 154.050 310.050 ;
        RECT 154.950 307.950 157.050 310.050 ;
        RECT 158.250 308.250 160.050 309.150 ;
        RECT 148.950 305.850 150.750 306.750 ;
        RECT 151.950 304.950 154.050 307.050 ;
        RECT 155.250 305.850 156.750 306.750 ;
        RECT 157.950 306.450 160.050 307.050 ;
        RECT 161.400 306.450 162.450 310.950 ;
        RECT 163.950 307.950 166.050 310.050 ;
        RECT 167.400 307.050 168.450 310.950 ;
        RECT 169.950 307.950 172.050 310.050 ;
        RECT 173.250 308.250 175.050 309.150 ;
        RECT 157.950 305.400 162.450 306.450 ;
        RECT 163.950 305.850 165.750 306.750 ;
        RECT 157.950 304.950 160.050 305.400 ;
        RECT 166.950 304.950 169.050 307.050 ;
        RECT 170.250 305.850 171.750 306.750 ;
        RECT 172.950 304.950 175.050 307.050 ;
        RECT 148.950 301.950 151.050 304.050 ;
        RECT 151.950 302.850 154.050 303.750 ;
        RECT 154.950 301.950 157.050 304.050 ;
        RECT 157.950 301.950 160.050 304.050 ;
        RECT 163.950 301.950 166.050 304.050 ;
        RECT 166.950 302.850 169.050 303.750 ;
        RECT 145.950 298.950 148.050 301.050 ;
        RECT 149.400 298.050 150.450 301.950 ;
        RECT 148.950 295.950 151.050 298.050 ;
        RECT 151.950 283.950 154.050 286.050 ;
        RECT 142.950 280.950 145.050 283.050 ;
        RECT 137.400 278.400 141.450 279.450 ;
        RECT 137.400 274.050 138.450 278.400 ;
        RECT 142.950 277.950 145.050 280.050 ;
        RECT 136.950 271.950 139.050 274.050 ;
        RECT 139.950 272.250 142.050 273.150 ;
        RECT 118.950 268.950 121.050 271.050 ;
        RECT 122.250 269.250 123.750 270.150 ;
        RECT 124.950 268.950 127.050 271.050 ;
        RECT 128.250 269.250 130.050 270.150 ;
        RECT 130.950 269.250 132.750 270.150 ;
        RECT 133.950 268.950 136.050 271.050 ;
        RECT 137.250 269.250 138.750 270.150 ;
        RECT 139.950 268.950 142.050 271.050 ;
        RECT 140.400 268.050 141.450 268.950 ;
        RECT 121.950 265.950 124.050 268.050 ;
        RECT 125.250 266.850 126.750 267.750 ;
        RECT 127.950 265.950 130.050 268.050 ;
        RECT 130.950 265.950 133.050 268.050 ;
        RECT 134.250 266.850 135.750 267.750 ;
        RECT 136.950 265.950 139.050 268.050 ;
        RECT 139.950 265.950 142.050 268.050 ;
        RECT 121.950 262.950 124.050 265.050 ;
        RECT 127.950 262.950 130.050 265.050 ;
        RECT 130.950 262.950 133.050 265.050 ;
        RECT 112.950 259.950 115.050 262.050 ;
        RECT 122.400 259.050 123.450 262.950 ;
        RECT 128.400 259.050 129.450 262.950 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 127.950 256.950 130.050 259.050 ;
        RECT 112.950 253.950 115.050 256.050 ;
        RECT 106.950 244.950 109.050 247.050 ;
        RECT 106.950 241.950 109.050 244.050 ;
        RECT 113.400 241.050 114.450 253.950 ;
        RECT 115.950 244.950 118.050 247.050 ;
        RECT 97.950 238.950 100.050 241.050 ;
        RECT 103.950 239.250 106.050 240.150 ;
        RECT 106.950 239.850 109.050 240.750 ;
        RECT 109.950 239.250 111.750 240.150 ;
        RECT 112.950 238.950 115.050 241.050 ;
        RECT 76.950 236.850 79.050 237.750 ;
        RECT 82.950 235.950 85.050 238.050 ;
        RECT 85.950 235.950 88.050 238.050 ;
        RECT 88.950 235.950 91.050 238.050 ;
        RECT 91.950 235.950 94.050 238.050 ;
        RECT 94.950 235.950 97.050 238.050 ;
        RECT 98.250 236.250 100.050 237.150 ;
        RECT 103.950 235.950 106.050 238.050 ;
        RECT 109.950 235.950 112.050 238.050 ;
        RECT 113.250 236.850 115.050 237.750 ;
        RECT 79.950 229.950 82.050 232.050 ;
        RECT 67.950 200.250 70.050 201.150 ;
        RECT 71.400 200.400 75.450 201.450 ;
        RECT 49.950 197.850 51.750 198.750 ;
        RECT 52.950 196.950 55.050 199.050 ;
        RECT 56.250 197.850 58.050 198.750 ;
        RECT 58.950 197.250 60.750 198.150 ;
        RECT 61.950 196.950 64.050 199.050 ;
        RECT 67.950 198.450 70.050 199.050 ;
        RECT 71.400 198.450 72.450 200.400 ;
        RECT 80.400 199.050 81.450 229.950 ;
        RECT 83.400 229.050 84.450 235.950 ;
        RECT 82.950 226.950 85.050 229.050 ;
        RECT 65.250 197.250 66.750 198.150 ;
        RECT 67.950 197.400 72.450 198.450 ;
        RECT 67.950 196.950 70.050 197.400 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 79.950 196.950 82.050 199.050 ;
        RECT 83.250 197.250 85.050 198.150 ;
        RECT 49.950 193.950 52.050 196.050 ;
        RECT 58.950 193.950 61.050 196.050 ;
        RECT 62.250 194.850 63.750 195.750 ;
        RECT 64.950 193.950 67.050 196.050 ;
        RECT 43.950 190.950 46.050 193.050 ;
        RECT 46.950 190.950 49.050 193.050 ;
        RECT 40.950 181.950 43.050 184.050 ;
        RECT 44.400 181.050 45.450 190.950 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 50.400 178.050 51.450 193.950 ;
        RECT 52.950 190.950 55.050 193.050 ;
        RECT 43.950 175.950 46.050 178.050 ;
        RECT 49.950 175.950 52.050 178.050 ;
        RECT 44.400 172.050 45.450 175.950 ;
        RECT 53.400 172.050 54.450 190.950 ;
        RECT 59.400 175.050 60.450 193.950 ;
        RECT 65.400 187.050 66.450 193.950 ;
        RECT 64.950 184.950 67.050 187.050 ;
        RECT 68.400 184.050 69.450 196.950 ;
        RECT 70.950 193.950 73.050 196.050 ;
        RECT 73.950 194.850 76.050 195.750 ;
        RECT 76.950 194.250 79.050 195.150 ;
        RECT 79.950 194.850 81.750 195.750 ;
        RECT 82.950 193.950 85.050 196.050 ;
        RECT 67.950 181.950 70.050 184.050 ;
        RECT 71.400 175.050 72.450 193.950 ;
        RECT 83.400 193.050 84.450 193.950 ;
        RECT 76.950 190.950 79.050 193.050 ;
        RECT 82.950 190.950 85.050 193.050 ;
        RECT 77.400 184.050 78.450 190.950 ;
        RECT 86.400 187.050 87.450 235.950 ;
        RECT 92.400 235.050 93.450 235.950 ;
        RECT 88.950 233.850 90.750 234.750 ;
        RECT 91.950 232.950 94.050 235.050 ;
        RECT 95.250 233.850 96.750 234.750 ;
        RECT 97.950 232.950 100.050 235.050 ;
        RECT 103.950 232.950 106.050 235.050 ;
        RECT 98.400 232.050 99.450 232.950 ;
        RECT 91.950 230.850 94.050 231.750 ;
        RECT 97.950 229.950 100.050 232.050 ;
        RECT 104.400 226.050 105.450 232.950 ;
        RECT 110.400 229.050 111.450 235.950 ;
        RECT 109.950 226.950 112.050 229.050 ;
        RECT 103.950 223.950 106.050 226.050 ;
        RECT 109.950 217.950 112.050 220.050 ;
        RECT 110.400 202.050 111.450 217.950 ;
        RECT 97.950 200.250 100.050 201.150 ;
        RECT 109.950 199.950 112.050 202.050 ;
        RECT 112.950 200.250 115.050 201.150 ;
        RECT 88.950 197.250 90.750 198.150 ;
        RECT 91.950 196.950 94.050 199.050 ;
        RECT 95.250 197.250 96.750 198.150 ;
        RECT 97.950 196.950 100.050 199.050 ;
        RECT 103.950 197.250 105.750 198.150 ;
        RECT 106.950 196.950 109.050 199.050 ;
        RECT 110.250 197.250 111.750 198.150 ;
        RECT 112.950 196.950 115.050 199.050 ;
        RECT 88.950 193.950 91.050 196.050 ;
        RECT 92.250 194.850 93.750 195.750 ;
        RECT 94.950 193.950 97.050 196.050 ;
        RECT 89.400 193.050 90.450 193.950 ;
        RECT 88.950 190.950 91.050 193.050 ;
        RECT 91.950 190.950 94.050 193.050 ;
        RECT 89.400 190.050 90.450 190.950 ;
        RECT 88.950 187.950 91.050 190.050 ;
        RECT 85.950 184.950 88.050 187.050 ;
        RECT 76.950 181.950 79.050 184.050 ;
        RECT 85.950 181.950 88.050 184.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 55.950 172.950 58.050 175.050 ;
        RECT 58.950 172.950 61.050 175.050 ;
        RECT 61.950 172.950 64.050 175.050 ;
        RECT 70.950 172.950 73.050 175.050 ;
        RECT 43.950 169.950 46.050 172.050 ;
        RECT 49.950 169.950 52.050 172.050 ;
        RECT 52.950 169.950 55.050 172.050 ;
        RECT 56.400 171.450 57.450 172.950 ;
        RECT 56.400 170.400 60.450 171.450 ;
        RECT 37.950 166.950 40.050 169.050 ;
        RECT 43.950 166.950 46.050 169.050 ;
        RECT 46.950 167.250 49.050 168.150 ;
        RECT 49.950 167.850 52.050 168.750 ;
        RECT 52.950 167.250 54.750 168.150 ;
        RECT 55.950 166.950 58.050 169.050 ;
        RECT 37.950 163.950 40.050 166.050 ;
        RECT 44.400 165.450 45.450 166.950 ;
        RECT 46.950 165.450 49.050 166.050 ;
        RECT 41.250 164.250 43.050 165.150 ;
        RECT 44.400 164.400 49.050 165.450 ;
        RECT 46.950 163.950 49.050 164.400 ;
        RECT 52.950 163.950 55.050 166.050 ;
        RECT 56.250 164.850 58.050 165.750 ;
        RECT 31.950 161.850 33.750 162.750 ;
        RECT 34.950 160.950 37.050 163.050 ;
        RECT 38.250 161.850 39.750 162.750 ;
        RECT 40.950 160.950 43.050 163.050 ;
        RECT 43.950 160.950 46.050 163.050 ;
        RECT 25.950 157.950 28.050 160.050 ;
        RECT 28.950 157.950 31.050 160.050 ;
        RECT 34.950 158.850 37.050 159.750 ;
        RECT 37.950 157.950 40.050 160.050 ;
        RECT 19.950 129.450 22.050 130.050 ;
        RECT 26.400 129.450 27.450 157.950 ;
        RECT 38.400 130.050 39.450 157.950 ;
        RECT 44.400 133.050 45.450 160.950 ;
        RECT 53.400 160.050 54.450 163.950 ;
        RECT 59.400 163.050 60.450 170.400 ;
        RECT 62.400 169.050 63.450 172.950 ;
        RECT 83.400 172.050 84.450 178.950 ;
        RECT 64.950 169.950 67.050 172.050 ;
        RECT 79.950 169.950 82.050 172.050 ;
        RECT 82.950 169.950 85.050 172.050 ;
        RECT 61.950 166.950 64.050 169.050 ;
        RECT 62.400 166.050 63.450 166.950 ;
        RECT 65.400 166.050 66.450 169.950 ;
        RECT 86.400 169.050 87.450 181.950 ;
        RECT 92.400 181.050 93.450 190.950 ;
        RECT 95.400 187.050 96.450 193.950 ;
        RECT 94.950 184.950 97.050 187.050 ;
        RECT 91.950 178.950 94.050 181.050 ;
        RECT 98.400 178.050 99.450 196.950 ;
        RECT 103.950 193.950 106.050 196.050 ;
        RECT 107.250 194.850 108.750 195.750 ;
        RECT 109.950 193.950 112.050 196.050 ;
        RECT 104.400 190.050 105.450 193.950 ;
        RECT 113.400 193.050 114.450 196.950 ;
        RECT 106.950 190.950 109.050 193.050 ;
        RECT 112.950 190.950 115.050 193.050 ;
        RECT 103.950 187.950 106.050 190.050 ;
        RECT 107.400 184.050 108.450 190.950 ;
        RECT 106.950 181.950 109.050 184.050 ;
        RECT 106.950 178.950 109.050 181.050 ;
        RECT 91.950 175.950 94.050 178.050 ;
        RECT 97.950 175.950 100.050 178.050 ;
        RECT 76.950 167.250 79.050 168.150 ;
        RECT 79.950 167.850 82.050 168.750 ;
        RECT 82.950 167.250 84.750 168.150 ;
        RECT 85.950 166.950 88.050 169.050 ;
        RECT 61.950 163.950 64.050 166.050 ;
        RECT 64.950 163.950 67.050 166.050 ;
        RECT 67.950 163.950 70.050 166.050 ;
        RECT 71.250 164.250 73.050 165.150 ;
        RECT 76.950 163.950 79.050 166.050 ;
        RECT 82.950 163.950 85.050 166.050 ;
        RECT 86.250 164.850 88.050 165.750 ;
        RECT 65.400 163.050 66.450 163.950 ;
        RECT 58.950 160.950 61.050 163.050 ;
        RECT 61.950 161.850 63.750 162.750 ;
        RECT 64.950 160.950 67.050 163.050 ;
        RECT 68.250 161.850 69.750 162.750 ;
        RECT 70.950 160.950 73.050 163.050 ;
        RECT 76.950 162.450 79.050 163.050 ;
        RECT 79.950 162.450 82.050 163.050 ;
        RECT 76.950 161.400 82.050 162.450 ;
        RECT 76.950 160.950 79.050 161.400 ;
        RECT 79.950 160.950 82.050 161.400 ;
        RECT 85.950 160.950 88.050 163.050 ;
        RECT 52.950 157.950 55.050 160.050 ;
        RECT 64.950 158.850 67.050 159.750 ;
        RECT 82.950 154.950 85.050 157.050 ;
        RECT 76.950 136.950 79.050 139.050 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 43.950 130.950 46.050 133.050 ;
        RECT 19.950 128.400 24.450 129.450 ;
        RECT 26.400 128.400 30.450 129.450 ;
        RECT 19.950 127.950 22.050 128.400 ;
        RECT 16.950 125.250 19.050 126.150 ;
        RECT 19.950 125.850 22.050 126.750 ;
        RECT 16.950 121.950 19.050 124.050 ;
        RECT 19.950 121.950 22.050 124.050 ;
        RECT 14.400 119.400 18.450 120.450 ;
        RECT 7.950 97.950 10.050 100.050 ;
        RECT 17.400 97.050 18.450 119.400 ;
        RECT 20.400 100.050 21.450 121.950 ;
        RECT 23.400 121.050 24.450 128.400 ;
        RECT 25.950 125.250 28.050 126.150 ;
        RECT 29.400 124.050 30.450 128.400 ;
        RECT 31.950 128.250 34.050 129.150 ;
        RECT 37.950 127.950 40.050 130.050 ;
        RECT 31.950 124.950 34.050 127.050 ;
        RECT 35.250 125.250 36.750 126.150 ;
        RECT 37.950 124.950 40.050 127.050 ;
        RECT 41.250 125.250 43.050 126.150 ;
        RECT 25.950 121.950 28.050 124.050 ;
        RECT 28.950 121.950 31.050 124.050 ;
        RECT 22.950 118.950 25.050 121.050 ;
        RECT 26.400 118.050 27.450 121.950 ;
        RECT 25.950 115.950 28.050 118.050 ;
        RECT 32.400 106.050 33.450 124.950 ;
        RECT 34.950 121.950 37.050 124.050 ;
        RECT 38.250 122.850 39.750 123.750 ;
        RECT 40.950 121.950 43.050 124.050 ;
        RECT 44.400 123.450 45.450 130.950 ;
        RECT 55.950 127.950 58.050 130.050 ;
        RECT 67.950 127.950 70.050 130.050 ;
        RECT 56.400 127.050 57.450 127.950 ;
        RECT 46.950 125.250 48.750 126.150 ;
        RECT 49.950 124.950 52.050 127.050 ;
        RECT 53.250 125.250 54.750 126.150 ;
        RECT 55.950 124.950 58.050 127.050 ;
        RECT 59.250 125.250 61.050 126.150 ;
        RECT 64.950 125.250 67.050 126.150 ;
        RECT 46.950 123.450 49.050 124.050 ;
        RECT 44.400 122.400 49.050 123.450 ;
        RECT 50.250 122.850 51.750 123.750 ;
        RECT 31.950 103.950 34.050 106.050 ;
        RECT 37.950 103.950 40.050 106.050 ;
        RECT 22.950 100.950 25.050 103.050 ;
        RECT 23.400 100.050 24.450 100.950 ;
        RECT 19.950 97.950 22.050 100.050 ;
        RECT 22.950 97.950 25.050 100.050 ;
        RECT 28.950 97.950 31.050 100.050 ;
        RECT 4.950 96.450 7.050 97.050 ;
        RECT 2.400 95.400 7.050 96.450 ;
        RECT 8.250 95.850 9.750 96.750 ;
        RECT 10.950 96.450 13.050 97.050 ;
        RECT 2.400 58.050 3.450 95.400 ;
        RECT 4.950 94.950 7.050 95.400 ;
        RECT 10.950 95.400 15.450 96.450 ;
        RECT 10.950 94.950 13.050 95.400 ;
        RECT 4.950 92.850 7.050 93.750 ;
        RECT 10.950 92.850 13.050 93.750 ;
        RECT 14.400 61.050 15.450 95.400 ;
        RECT 16.950 94.950 19.050 97.050 ;
        RECT 20.250 95.250 22.050 96.150 ;
        RECT 22.950 95.850 25.050 96.750 ;
        RECT 25.950 95.250 28.050 96.150 ;
        RECT 28.950 95.850 31.050 96.750 ;
        RECT 31.950 95.250 34.050 96.150 ;
        RECT 34.950 94.950 37.050 97.050 ;
        RECT 16.950 92.850 18.750 93.750 ;
        RECT 19.950 91.950 22.050 94.050 ;
        RECT 22.950 91.950 25.050 94.050 ;
        RECT 25.950 91.950 28.050 94.050 ;
        RECT 28.950 91.950 31.050 94.050 ;
        RECT 31.950 91.950 34.050 94.050 ;
        RECT 13.950 58.950 16.050 61.050 ;
        RECT 14.400 58.050 15.450 58.950 ;
        RECT 23.400 58.050 24.450 91.950 ;
        RECT 26.400 91.050 27.450 91.950 ;
        RECT 25.950 88.950 28.050 91.050 ;
        RECT 29.400 60.450 30.450 91.950 ;
        RECT 32.400 91.050 33.450 91.950 ;
        RECT 31.950 88.950 34.050 91.050 ;
        RECT 35.400 64.050 36.450 94.950 ;
        RECT 34.950 61.950 37.050 64.050 ;
        RECT 26.400 59.400 30.450 60.450 ;
        RECT 1.950 55.950 4.050 58.050 ;
        RECT 7.950 57.450 10.050 58.050 ;
        RECT 5.250 56.250 6.750 57.150 ;
        RECT 7.950 56.400 12.450 57.450 ;
        RECT 7.950 55.950 10.050 56.400 ;
        RECT 1.950 53.850 3.750 54.750 ;
        RECT 4.950 52.950 7.050 55.050 ;
        RECT 8.250 53.850 10.050 54.750 ;
        RECT 5.400 31.050 6.450 52.950 ;
        RECT 11.400 49.050 12.450 56.400 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 19.950 57.450 22.050 58.050 ;
        RECT 22.950 57.450 25.050 58.050 ;
        RECT 17.250 56.250 18.750 57.150 ;
        RECT 19.950 56.400 25.050 57.450 ;
        RECT 19.950 55.950 22.050 56.400 ;
        RECT 22.950 55.950 25.050 56.400 ;
        RECT 13.950 53.850 15.750 54.750 ;
        RECT 16.950 52.950 19.050 55.050 ;
        RECT 20.250 53.850 22.050 54.750 ;
        RECT 13.950 49.950 16.050 52.050 ;
        RECT 10.950 46.950 13.050 49.050 ;
        RECT 4.950 28.950 7.050 31.050 ;
        RECT 5.400 24.450 6.450 28.950 ;
        RECT 10.950 25.950 13.050 28.050 ;
        RECT 5.400 23.400 9.450 24.450 ;
        RECT 8.400 22.050 9.450 23.400 ;
        RECT 11.400 22.050 12.450 25.950 ;
        RECT 14.400 25.050 15.450 49.950 ;
        RECT 17.400 28.050 18.450 52.950 ;
        RECT 26.400 52.050 27.450 59.400 ;
        RECT 34.950 58.950 37.050 61.050 ;
        RECT 35.400 58.050 36.450 58.950 ;
        RECT 28.950 55.950 31.050 58.050 ;
        RECT 32.250 56.250 33.750 57.150 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 38.400 55.050 39.450 103.950 ;
        RECT 41.400 100.050 42.450 121.950 ;
        RECT 44.400 118.050 45.450 122.400 ;
        RECT 46.950 121.950 49.050 122.400 ;
        RECT 52.950 121.950 55.050 124.050 ;
        RECT 56.250 122.850 57.750 123.750 ;
        RECT 58.950 121.950 61.050 124.050 ;
        RECT 64.950 121.950 67.050 124.050 ;
        RECT 43.950 115.950 46.050 118.050 ;
        RECT 59.400 108.450 60.450 121.950 ;
        RECT 65.400 121.050 66.450 121.950 ;
        RECT 64.950 118.950 67.050 121.050 ;
        RECT 56.400 107.400 60.450 108.450 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 47.400 100.050 48.450 100.950 ;
        RECT 40.950 97.950 43.050 100.050 ;
        RECT 46.950 97.950 49.050 100.050 ;
        RECT 53.400 97.050 54.450 100.950 ;
        RECT 56.400 100.050 57.450 107.400 ;
        RECT 58.950 103.950 61.050 106.050 ;
        RECT 55.950 97.950 58.050 100.050 ;
        RECT 40.950 94.950 43.050 97.050 ;
        RECT 44.250 95.250 46.050 96.150 ;
        RECT 46.950 95.850 49.050 96.750 ;
        RECT 49.950 95.250 52.050 96.150 ;
        RECT 52.950 94.950 55.050 97.050 ;
        RECT 53.400 94.050 54.450 94.950 ;
        RECT 59.400 94.050 60.450 103.950 ;
        RECT 64.950 100.950 67.050 103.050 ;
        RECT 40.950 92.850 42.750 93.750 ;
        RECT 43.950 91.950 46.050 94.050 ;
        RECT 46.950 91.950 49.050 94.050 ;
        RECT 49.950 91.950 52.050 94.050 ;
        RECT 52.950 91.950 55.050 94.050 ;
        RECT 58.950 91.950 61.050 94.050 ;
        RECT 62.250 92.250 64.050 93.150 ;
        RECT 44.400 91.050 45.450 91.950 ;
        RECT 43.950 88.950 46.050 91.050 ;
        RECT 47.400 79.050 48.450 91.950 ;
        RECT 52.950 89.850 54.750 90.750 ;
        RECT 55.950 88.950 58.050 91.050 ;
        RECT 59.250 89.850 60.750 90.750 ;
        RECT 61.950 88.950 64.050 91.050 ;
        RECT 55.950 86.850 58.050 87.750 ;
        RECT 46.950 76.950 49.050 79.050 ;
        RECT 52.950 73.950 55.050 76.050 ;
        RECT 46.950 67.950 49.050 70.050 ;
        RECT 47.400 58.050 48.450 67.950 ;
        RECT 49.950 61.950 52.050 64.050 ;
        RECT 44.250 56.250 45.750 57.150 ;
        RECT 46.950 55.950 49.050 58.050 ;
        RECT 28.950 53.850 30.750 54.750 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 35.250 53.850 37.050 54.750 ;
        RECT 37.950 52.950 40.050 55.050 ;
        RECT 40.950 53.850 42.750 54.750 ;
        RECT 43.950 52.950 46.050 55.050 ;
        RECT 47.250 53.850 49.050 54.750 ;
        RECT 44.400 52.050 45.450 52.950 ;
        RECT 25.950 49.950 28.050 52.050 ;
        RECT 37.950 49.950 40.050 52.050 ;
        RECT 43.950 49.950 46.050 52.050 ;
        RECT 46.950 49.950 49.050 52.050 ;
        RECT 38.400 49.050 39.450 49.950 ;
        RECT 37.950 46.950 40.050 49.050 ;
        RECT 19.950 28.950 22.050 31.050 ;
        RECT 34.950 28.950 37.050 31.050 ;
        RECT 20.400 28.050 21.450 28.950 ;
        RECT 16.950 25.950 19.050 28.050 ;
        RECT 19.950 25.950 22.050 28.050 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 23.250 19.050 24.150 ;
        RECT 19.950 23.850 22.050 24.750 ;
        RECT 22.950 23.250 24.750 24.150 ;
        RECT 25.950 22.950 28.050 25.050 ;
        RECT 14.400 22.050 15.450 22.950 ;
        RECT 35.400 22.050 36.450 28.950 ;
        RECT 47.400 28.050 48.450 49.950 ;
        RECT 50.400 28.050 51.450 61.950 ;
        RECT 53.400 58.050 54.450 73.950 ;
        RECT 58.950 64.950 61.050 67.050 ;
        RECT 52.950 55.950 55.050 58.050 ;
        RECT 55.950 55.950 58.050 58.050 ;
        RECT 59.400 55.050 60.450 64.950 ;
        RECT 62.400 61.050 63.450 88.950 ;
        RECT 65.400 76.050 66.450 100.950 ;
        RECT 68.400 100.050 69.450 127.950 ;
        RECT 74.400 127.050 75.450 133.950 ;
        RECT 77.400 127.050 78.450 136.950 ;
        RECT 70.950 125.250 73.050 126.150 ;
        RECT 73.950 124.950 76.050 127.050 ;
        RECT 76.950 124.950 79.050 127.050 ;
        RECT 73.950 122.250 76.050 123.150 ;
        RECT 76.950 122.850 79.050 123.750 ;
        RECT 73.950 118.950 76.050 121.050 ;
        RECT 83.400 114.450 84.450 154.950 ;
        RECT 86.400 136.050 87.450 160.950 ;
        RECT 85.950 133.950 88.050 136.050 ;
        RECT 85.950 127.950 88.050 130.050 ;
        RECT 86.400 127.050 87.450 127.950 ;
        RECT 85.950 124.950 88.050 127.050 ;
        RECT 85.950 122.850 88.050 123.750 ;
        RECT 92.400 123.450 93.450 175.950 ;
        RECT 97.950 172.950 100.050 175.050 ;
        RECT 98.400 166.050 99.450 172.950 ;
        RECT 107.400 169.050 108.450 178.950 ;
        RECT 109.950 175.950 112.050 178.050 ;
        RECT 110.400 169.050 111.450 175.950 ;
        RECT 116.400 171.450 117.450 244.950 ;
        RECT 121.950 241.950 124.050 244.050 ;
        RECT 122.400 238.050 123.450 241.950 ;
        RECT 131.400 241.050 132.450 262.950 ;
        RECT 137.400 262.050 138.450 265.950 ;
        RECT 136.950 259.950 139.050 262.050 ;
        RECT 140.400 256.050 141.450 265.950 ;
        RECT 143.400 262.050 144.450 277.950 ;
        RECT 152.400 277.050 153.450 283.950 ;
        RECT 155.400 280.050 156.450 301.950 ;
        RECT 154.950 277.950 157.050 280.050 ;
        RECT 155.400 277.050 156.450 277.950 ;
        RECT 148.950 275.250 151.050 276.150 ;
        RECT 151.950 274.950 154.050 277.050 ;
        RECT 154.950 274.950 157.050 277.050 ;
        RECT 158.400 274.050 159.450 301.950 ;
        RECT 160.950 298.950 163.050 301.050 ;
        RECT 145.950 272.250 147.750 273.150 ;
        RECT 148.950 271.950 151.050 274.050 ;
        RECT 152.250 272.250 153.750 273.150 ;
        RECT 154.950 271.950 157.050 274.050 ;
        RECT 157.950 271.950 160.050 274.050 ;
        RECT 145.950 268.950 148.050 271.050 ;
        RECT 151.950 268.950 154.050 271.050 ;
        RECT 155.250 269.850 157.050 270.750 ;
        RECT 161.400 270.450 162.450 298.950 ;
        RECT 164.400 277.050 165.450 301.950 ;
        RECT 176.400 301.050 177.450 337.950 ;
        RECT 179.400 337.050 180.450 337.950 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 313.950 184.050 316.050 ;
        RECT 178.950 311.250 181.050 312.150 ;
        RECT 181.950 311.850 184.050 312.750 ;
        RECT 184.950 311.250 186.750 312.150 ;
        RECT 187.950 310.950 190.050 313.050 ;
        RECT 191.400 310.050 192.450 373.950 ;
        RECT 193.950 350.400 196.050 352.500 ;
        RECT 197.400 352.050 198.450 379.950 ;
        RECT 202.950 376.950 205.050 379.050 ;
        RECT 206.250 377.850 207.750 378.750 ;
        RECT 203.400 373.050 204.450 376.950 ;
        RECT 202.950 370.950 205.050 373.050 ;
        RECT 211.950 370.950 214.050 373.050 ;
        RECT 194.400 333.600 195.600 350.400 ;
        RECT 196.950 349.950 199.050 352.050 ;
        RECT 202.950 349.950 205.050 352.050 ;
        RECT 196.950 346.950 199.050 349.050 ;
        RECT 193.950 331.500 196.050 333.600 ;
        RECT 197.400 327.450 198.450 346.950 ;
        RECT 199.950 341.250 202.050 342.150 ;
        RECT 199.950 337.950 202.050 340.050 ;
        RECT 200.400 337.050 201.450 337.950 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 194.400 326.400 198.450 327.450 ;
        RECT 194.400 316.050 195.450 326.400 ;
        RECT 196.950 319.950 199.050 322.050 ;
        RECT 197.400 316.050 198.450 319.950 ;
        RECT 193.950 313.950 196.050 316.050 ;
        RECT 196.950 313.950 199.050 316.050 ;
        RECT 193.950 310.950 196.050 313.050 ;
        RECT 197.250 311.850 198.750 312.750 ;
        RECT 199.950 310.950 202.050 313.050 ;
        RECT 178.950 307.950 181.050 310.050 ;
        RECT 181.950 307.950 184.050 310.050 ;
        RECT 184.950 307.950 187.050 310.050 ;
        RECT 188.250 308.850 190.050 309.750 ;
        RECT 190.950 307.950 193.050 310.050 ;
        RECT 193.950 308.850 196.050 309.750 ;
        RECT 196.950 307.950 199.050 310.050 ;
        RECT 199.950 308.850 202.050 309.750 ;
        RECT 166.950 298.950 169.050 301.050 ;
        RECT 175.950 298.950 178.050 301.050 ;
        RECT 163.950 274.950 166.050 277.050 ;
        RECT 163.950 271.950 166.050 274.050 ;
        RECT 164.400 271.050 165.450 271.950 ;
        RECT 158.400 269.400 162.450 270.450 ;
        RECT 152.400 268.050 153.450 268.950 ;
        RECT 151.950 265.950 154.050 268.050 ;
        RECT 154.950 265.950 157.050 268.050 ;
        RECT 155.400 262.050 156.450 265.950 ;
        RECT 142.950 259.950 145.050 262.050 ;
        RECT 151.950 259.950 154.050 262.050 ;
        RECT 154.950 259.950 157.050 262.050 ;
        RECT 139.950 253.950 142.050 256.050 ;
        RECT 145.950 250.950 148.050 253.050 ;
        RECT 136.950 244.950 139.050 247.050 ;
        RECT 137.400 244.050 138.450 244.950 ;
        RECT 136.950 241.950 139.050 244.050 ;
        RECT 142.950 241.950 145.050 244.050 ;
        RECT 143.400 241.050 144.450 241.950 ;
        RECT 130.950 238.950 133.050 241.050 ;
        RECT 133.950 239.250 136.050 240.150 ;
        RECT 136.950 239.850 139.050 240.750 ;
        RECT 139.950 239.250 141.750 240.150 ;
        RECT 142.950 238.950 145.050 241.050 ;
        RECT 118.950 235.950 121.050 238.050 ;
        RECT 121.950 235.950 124.050 238.050 ;
        RECT 124.950 235.950 127.050 238.050 ;
        RECT 128.250 236.250 130.050 237.150 ;
        RECT 130.950 235.950 133.050 238.050 ;
        RECT 133.950 235.950 136.050 238.050 ;
        RECT 136.950 235.950 139.050 238.050 ;
        RECT 139.950 235.950 142.050 238.050 ;
        RECT 143.250 236.850 145.050 237.750 ;
        RECT 118.950 233.850 120.750 234.750 ;
        RECT 121.950 232.950 124.050 235.050 ;
        RECT 125.250 233.850 126.750 234.750 ;
        RECT 127.950 232.950 130.050 235.050 ;
        RECT 121.950 230.850 124.050 231.750 ;
        RECT 131.400 231.450 132.450 235.950 ;
        RECT 134.400 235.050 135.450 235.950 ;
        RECT 133.950 232.950 136.050 235.050 ;
        RECT 128.400 230.400 132.450 231.450 ;
        RECT 118.950 223.950 121.050 226.050 ;
        RECT 119.400 202.050 120.450 223.950 ;
        RECT 124.950 220.950 127.050 223.050 ;
        RECT 121.950 211.950 124.050 214.050 ;
        RECT 118.950 199.950 121.050 202.050 ;
        RECT 118.950 197.250 121.050 198.150 ;
        RECT 118.950 193.950 121.050 196.050 ;
        RECT 119.400 184.050 120.450 193.950 ;
        RECT 122.400 193.050 123.450 211.950 ;
        RECT 125.400 205.050 126.450 220.950 ;
        RECT 128.400 220.050 129.450 230.400 ;
        RECT 134.400 229.050 135.450 232.950 ;
        RECT 133.950 226.950 136.050 229.050 ;
        RECT 137.400 226.050 138.450 235.950 ;
        RECT 136.950 223.950 139.050 226.050 ;
        RECT 127.950 217.950 130.050 220.050 ;
        RECT 130.950 217.950 133.050 220.050 ;
        RECT 124.950 202.950 127.050 205.050 ;
        RECT 124.950 197.850 127.050 198.750 ;
        RECT 127.950 197.250 130.050 198.150 ;
        RECT 127.950 193.950 130.050 196.050 ;
        RECT 128.400 193.050 129.450 193.950 ;
        RECT 121.950 190.950 124.050 193.050 ;
        RECT 127.950 190.950 130.050 193.050 ;
        RECT 118.950 181.950 121.050 184.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 113.400 170.400 117.450 171.450 ;
        RECT 106.950 166.950 109.050 169.050 ;
        RECT 109.950 166.950 112.050 169.050 ;
        RECT 94.950 164.250 96.750 165.150 ;
        RECT 97.950 163.950 100.050 166.050 ;
        RECT 101.250 164.250 103.050 165.150 ;
        RECT 106.950 164.850 109.050 165.750 ;
        RECT 109.950 164.250 112.050 165.150 ;
        RECT 94.950 160.950 97.050 163.050 ;
        RECT 98.250 161.850 99.750 162.750 ;
        RECT 100.950 160.950 103.050 163.050 ;
        RECT 109.950 160.950 112.050 163.050 ;
        RECT 95.400 154.050 96.450 160.950 ;
        RECT 94.950 151.950 97.050 154.050 ;
        RECT 113.400 139.050 114.450 170.400 ;
        RECT 115.950 166.950 118.050 169.050 ;
        RECT 115.950 164.850 118.050 165.750 ;
        RECT 115.950 160.950 118.050 163.050 ;
        RECT 116.400 154.050 117.450 160.950 ;
        RECT 115.950 151.950 118.050 154.050 ;
        RECT 115.950 148.950 118.050 151.050 ;
        RECT 112.950 136.950 115.050 139.050 ;
        RECT 109.950 131.250 112.050 132.150 ;
        RECT 116.400 130.050 117.450 148.950 ;
        RECT 97.950 127.950 100.050 130.050 ;
        RECT 103.950 127.950 106.050 130.050 ;
        RECT 106.950 128.250 108.750 129.150 ;
        RECT 109.950 127.950 112.050 130.050 ;
        RECT 113.250 128.250 114.750 129.150 ;
        RECT 115.950 127.950 118.050 130.050 ;
        RECT 98.400 127.050 99.450 127.950 ;
        RECT 104.400 127.050 105.450 127.950 ;
        RECT 94.950 125.250 96.750 126.150 ;
        RECT 97.950 124.950 100.050 127.050 ;
        RECT 103.950 124.950 106.050 127.050 ;
        RECT 106.950 126.450 109.050 127.050 ;
        RECT 106.950 125.400 111.450 126.450 ;
        RECT 106.950 124.950 109.050 125.400 ;
        RECT 94.950 123.450 97.050 124.050 ;
        RECT 88.950 122.250 91.050 123.150 ;
        RECT 92.400 122.400 97.050 123.450 ;
        RECT 98.250 122.850 100.050 123.750 ;
        RECT 94.950 121.950 97.050 122.400 ;
        RECT 100.950 122.250 103.050 123.150 ;
        RECT 103.950 122.850 106.050 123.750 ;
        RECT 88.950 118.950 91.050 121.050 ;
        RECT 100.950 118.950 103.050 121.050 ;
        RECT 106.950 118.950 109.050 121.050 ;
        RECT 89.400 115.050 90.450 118.950 ;
        RECT 83.400 113.400 87.450 114.450 ;
        RECT 79.950 106.950 82.050 109.050 ;
        RECT 67.950 97.950 70.050 100.050 ;
        RECT 64.950 73.950 67.050 76.050 ;
        RECT 64.950 70.950 67.050 73.050 ;
        RECT 65.400 61.050 66.450 70.950 ;
        RECT 68.400 61.050 69.450 97.950 ;
        RECT 80.400 97.050 81.450 106.950 ;
        RECT 86.400 99.450 87.450 113.400 ;
        RECT 88.950 112.950 91.050 115.050 ;
        RECT 97.950 112.950 100.050 115.050 ;
        RECT 86.400 98.400 90.450 99.450 ;
        RECT 73.950 94.950 76.050 97.050 ;
        RECT 77.250 95.250 78.750 96.150 ;
        RECT 79.950 94.950 82.050 97.050 ;
        RECT 85.950 94.950 88.050 97.050 ;
        RECT 70.950 91.950 73.050 94.050 ;
        RECT 74.250 92.850 75.750 93.750 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 80.250 92.850 82.050 93.750 ;
        RECT 85.950 92.850 88.050 93.750 ;
        RECT 70.950 89.850 73.050 90.750 ;
        RECT 73.950 88.950 76.050 91.050 ;
        RECT 77.400 90.450 78.450 91.950 ;
        RECT 77.400 89.400 81.450 90.450 ;
        RECT 70.950 76.950 73.050 79.050 ;
        RECT 61.950 58.950 64.050 61.050 ;
        RECT 64.950 58.950 67.050 61.050 ;
        RECT 67.950 58.950 70.050 61.050 ;
        RECT 71.400 60.450 72.450 76.950 ;
        RECT 74.400 73.050 75.450 88.950 ;
        RECT 80.400 88.050 81.450 89.400 ;
        RECT 79.950 85.950 82.050 88.050 ;
        RECT 73.950 70.950 76.050 73.050 ;
        RECT 76.950 67.950 79.050 70.050 ;
        RECT 71.400 59.400 75.450 60.450 ;
        RECT 52.950 53.250 55.050 54.150 ;
        RECT 55.950 53.850 58.050 54.750 ;
        RECT 58.950 52.950 61.050 55.050 ;
        RECT 61.950 53.250 64.050 54.150 ;
        RECT 52.950 49.950 55.050 52.050 ;
        RECT 61.950 49.950 64.050 52.050 ;
        RECT 53.400 49.050 54.450 49.950 ;
        RECT 65.400 49.050 66.450 58.950 ;
        RECT 68.400 58.050 69.450 58.950 ;
        RECT 74.400 58.050 75.450 59.400 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 71.250 56.250 72.750 57.150 ;
        RECT 73.950 55.950 76.050 58.050 ;
        RECT 67.950 53.850 69.750 54.750 ;
        RECT 70.950 52.950 73.050 55.050 ;
        RECT 74.250 53.850 76.050 54.750 ;
        RECT 71.400 49.050 72.450 52.950 ;
        RECT 77.400 49.050 78.450 67.950 ;
        RECT 89.400 64.050 90.450 98.400 ;
        RECT 98.400 94.050 99.450 112.950 ;
        RECT 101.400 103.050 102.450 118.950 ;
        RECT 103.950 115.950 106.050 118.050 ;
        RECT 100.950 100.950 103.050 103.050 ;
        RECT 104.400 99.450 105.450 115.950 ;
        RECT 101.400 98.400 105.450 99.450 ;
        RECT 101.400 97.050 102.450 98.400 ;
        RECT 107.400 97.050 108.450 118.950 ;
        RECT 110.400 115.050 111.450 125.400 ;
        RECT 112.950 124.950 115.050 127.050 ;
        RECT 116.250 125.850 118.050 126.750 ;
        RECT 113.400 124.050 114.450 124.950 ;
        RECT 112.950 121.950 115.050 124.050 ;
        RECT 109.950 112.950 112.050 115.050 ;
        RECT 100.950 94.950 103.050 97.050 ;
        RECT 104.250 95.250 105.750 96.150 ;
        RECT 106.950 94.950 109.050 97.050 ;
        RECT 91.950 92.850 94.050 93.750 ;
        RECT 94.950 91.950 97.050 94.050 ;
        RECT 97.950 91.950 100.050 94.050 ;
        RECT 101.250 92.850 102.750 93.750 ;
        RECT 103.950 91.950 106.050 94.050 ;
        RECT 107.250 92.850 109.050 93.750 ;
        RECT 95.400 67.050 96.450 91.950 ;
        RECT 97.950 89.850 100.050 90.750 ;
        RECT 104.400 82.050 105.450 91.950 ;
        RECT 103.950 79.950 106.050 82.050 ;
        RECT 94.950 64.950 97.050 67.050 ;
        RECT 79.950 61.950 82.050 64.050 ;
        RECT 88.950 61.950 91.050 64.050 ;
        RECT 80.400 58.050 81.450 61.950 ;
        RECT 85.950 59.250 88.050 60.150 ;
        RECT 97.950 58.950 100.050 61.050 ;
        RECT 103.950 58.950 106.050 61.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 83.250 56.250 84.750 57.150 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 89.250 56.250 91.050 57.150 ;
        RECT 79.950 53.850 81.750 54.750 ;
        RECT 82.950 52.950 85.050 55.050 ;
        RECT 52.950 46.950 55.050 49.050 ;
        RECT 64.950 46.950 67.050 49.050 ;
        RECT 70.950 46.950 73.050 49.050 ;
        RECT 76.950 46.950 79.050 49.050 ;
        RECT 53.400 43.050 54.450 46.950 ;
        RECT 71.400 46.050 72.450 46.950 ;
        RECT 64.950 43.950 67.050 46.050 ;
        RECT 70.950 43.950 73.050 46.050 ;
        RECT 52.950 40.950 55.050 43.050 ;
        RECT 52.950 37.950 55.050 40.050 ;
        RECT 37.950 25.950 40.050 28.050 ;
        RECT 46.950 25.950 49.050 28.050 ;
        RECT 49.950 25.950 52.050 28.050 ;
        RECT 38.400 25.050 39.450 25.950 ;
        RECT 53.400 25.050 54.450 37.950 ;
        RECT 61.950 34.950 64.050 37.050 ;
        RECT 37.950 22.950 40.050 25.050 ;
        RECT 41.250 23.250 42.750 24.150 ;
        RECT 43.950 22.950 46.050 25.050 ;
        RECT 46.950 22.950 49.050 25.050 ;
        RECT 50.250 23.250 51.750 24.150 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 55.950 22.950 58.050 25.050 ;
        RECT 56.400 22.050 57.450 22.950 ;
        RECT 4.950 20.250 6.750 21.150 ;
        RECT 7.950 19.950 10.050 22.050 ;
        RECT 10.950 19.950 13.050 22.050 ;
        RECT 13.950 19.950 16.050 22.050 ;
        RECT 16.950 19.950 19.050 22.050 ;
        RECT 22.950 19.950 25.050 22.050 ;
        RECT 26.250 20.850 28.050 21.750 ;
        RECT 34.950 19.950 37.050 22.050 ;
        RECT 38.250 20.850 39.750 21.750 ;
        RECT 40.950 19.950 43.050 22.050 ;
        RECT 44.250 20.850 46.050 21.750 ;
        RECT 46.950 20.850 48.750 21.750 ;
        RECT 49.950 19.950 52.050 22.050 ;
        RECT 53.250 20.850 54.750 21.750 ;
        RECT 55.950 19.950 58.050 22.050 ;
        RECT 11.400 19.050 12.450 19.950 ;
        RECT 4.950 16.950 7.050 19.050 ;
        RECT 8.250 17.850 9.750 18.750 ;
        RECT 10.950 16.950 13.050 19.050 ;
        RECT 14.250 17.850 16.050 18.750 ;
        RECT 34.950 17.850 37.050 18.750 ;
        RECT 55.950 17.850 58.050 18.750 ;
        RECT 62.400 18.450 63.450 34.950 ;
        RECT 65.400 28.050 66.450 43.950 ;
        RECT 83.400 40.050 84.450 52.950 ;
        RECT 86.400 51.450 87.450 55.950 ;
        RECT 98.400 55.050 99.450 58.950 ;
        RECT 104.400 55.050 105.450 58.950 ;
        RECT 88.950 52.950 91.050 55.050 ;
        RECT 94.950 53.250 96.750 54.150 ;
        RECT 97.950 52.950 100.050 55.050 ;
        RECT 101.250 53.250 102.750 54.150 ;
        RECT 103.950 52.950 106.050 55.050 ;
        RECT 107.250 53.250 109.050 54.150 ;
        RECT 86.400 50.400 90.450 51.450 ;
        RECT 82.950 37.950 85.050 40.050 ;
        RECT 82.950 28.950 85.050 31.050 ;
        RECT 64.950 25.950 67.050 28.050 ;
        RECT 70.950 25.950 73.050 28.050 ;
        RECT 79.950 25.950 82.050 28.050 ;
        RECT 64.950 20.250 66.750 21.150 ;
        RECT 67.950 19.950 70.050 22.050 ;
        RECT 71.400 19.050 72.450 25.950 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 74.400 22.050 75.450 22.950 ;
        RECT 73.950 19.950 76.050 22.050 ;
        RECT 76.950 19.950 79.050 22.050 ;
        RECT 80.400 19.050 81.450 25.950 ;
        RECT 83.400 22.050 84.450 28.950 ;
        RECT 89.400 28.050 90.450 50.400 ;
        RECT 94.950 49.950 97.050 52.050 ;
        RECT 98.250 50.850 99.750 51.750 ;
        RECT 100.950 49.950 103.050 52.050 ;
        RECT 104.250 50.850 105.750 51.750 ;
        RECT 106.950 49.950 109.050 52.050 ;
        RECT 95.400 49.050 96.450 49.950 ;
        RECT 94.950 46.950 97.050 49.050 ;
        RECT 101.400 34.050 102.450 49.950 ;
        RECT 103.950 46.950 106.050 49.050 ;
        RECT 100.950 31.950 103.050 34.050 ;
        RECT 104.400 30.450 105.450 46.950 ;
        RECT 110.400 37.050 111.450 112.950 ;
        RECT 119.400 103.050 120.450 178.950 ;
        RECT 122.400 169.050 123.450 190.950 ;
        RECT 131.400 189.450 132.450 217.950 ;
        RECT 140.400 214.050 141.450 235.950 ;
        RECT 139.950 211.950 142.050 214.050 ;
        RECT 142.950 205.950 145.050 208.050 ;
        RECT 133.950 202.950 136.050 205.050 ;
        RECT 128.400 188.400 132.450 189.450 ;
        RECT 128.400 187.050 129.450 188.400 ;
        RECT 127.950 184.950 130.050 187.050 ;
        RECT 130.950 184.950 133.050 187.050 ;
        RECT 127.950 181.950 130.050 184.050 ;
        RECT 124.950 169.950 127.050 172.050 ;
        RECT 121.950 166.950 124.050 169.050 ;
        RECT 125.400 166.050 126.450 169.950 ;
        RECT 128.400 169.050 129.450 181.950 ;
        RECT 127.950 166.950 130.050 169.050 ;
        RECT 131.400 166.050 132.450 184.950 ;
        RECT 134.400 184.050 135.450 202.950 ;
        RECT 143.400 202.050 144.450 205.950 ;
        RECT 146.400 205.050 147.450 250.950 ;
        RECT 148.950 244.950 151.050 247.050 ;
        RECT 149.400 238.050 150.450 244.950 ;
        RECT 152.400 241.050 153.450 259.950 ;
        RECT 151.950 238.950 154.050 241.050 ;
        RECT 158.400 240.450 159.450 269.400 ;
        RECT 163.950 268.950 166.050 271.050 ;
        RECT 160.950 266.250 163.050 267.150 ;
        RECT 163.950 266.850 166.050 267.750 ;
        RECT 160.950 262.950 163.050 265.050 ;
        RECT 167.400 264.450 168.450 298.950 ;
        RECT 169.950 279.450 172.050 280.050 ;
        RECT 172.950 279.450 175.050 280.050 ;
        RECT 169.950 278.400 175.050 279.450 ;
        RECT 169.950 277.950 172.050 278.400 ;
        RECT 172.950 277.950 175.050 278.400 ;
        RECT 172.950 275.250 175.050 276.150 ;
        RECT 179.400 274.050 180.450 307.950 ;
        RECT 169.950 272.250 171.750 273.150 ;
        RECT 172.950 271.950 175.050 274.050 ;
        RECT 176.250 272.250 177.750 273.150 ;
        RECT 178.950 271.950 181.050 274.050 ;
        RECT 169.950 270.450 172.050 271.050 ;
        RECT 169.950 269.400 174.450 270.450 ;
        RECT 169.950 268.950 172.050 269.400 ;
        RECT 173.400 268.050 174.450 269.400 ;
        RECT 175.950 268.950 178.050 271.050 ;
        RECT 179.250 269.850 181.050 270.750 ;
        RECT 169.950 265.950 172.050 268.050 ;
        RECT 172.950 265.950 175.050 268.050 ;
        RECT 164.400 263.400 168.450 264.450 ;
        RECT 161.400 244.050 162.450 262.950 ;
        RECT 160.950 241.950 163.050 244.050 ;
        RECT 158.400 239.400 162.450 240.450 ;
        RECT 148.950 235.950 151.050 238.050 ;
        RECT 151.950 237.450 154.050 238.050 ;
        RECT 154.950 237.450 157.050 238.050 ;
        RECT 151.950 236.400 157.050 237.450 ;
        RECT 151.950 235.950 154.050 236.400 ;
        RECT 154.950 235.950 157.050 236.400 ;
        RECT 158.250 236.250 160.050 237.150 ;
        RECT 148.950 233.850 150.750 234.750 ;
        RECT 151.950 232.950 154.050 235.050 ;
        RECT 155.250 233.850 156.750 234.750 ;
        RECT 157.950 232.950 160.050 235.050 ;
        RECT 148.950 229.950 151.050 232.050 ;
        RECT 151.950 230.850 154.050 231.750 ;
        RECT 154.950 229.950 157.050 232.050 ;
        RECT 161.400 231.450 162.450 239.400 ;
        RECT 164.400 235.050 165.450 263.400 ;
        RECT 170.400 250.050 171.450 265.950 ;
        RECT 176.400 262.050 177.450 268.950 ;
        RECT 175.950 259.950 178.050 262.050 ;
        RECT 169.950 247.950 172.050 250.050 ;
        RECT 166.950 244.950 169.050 247.050 ;
        RECT 167.400 238.050 168.450 244.950 ;
        RECT 170.400 241.050 171.450 247.950 ;
        RECT 169.950 238.950 172.050 241.050 ;
        RECT 173.250 239.250 174.750 240.150 ;
        RECT 175.950 238.950 178.050 241.050 ;
        RECT 178.950 238.950 181.050 241.050 ;
        RECT 179.400 238.050 180.450 238.950 ;
        RECT 182.400 238.050 183.450 307.950 ;
        RECT 185.400 277.050 186.450 307.950 ;
        RECT 190.950 304.950 193.050 307.050 ;
        RECT 191.400 277.050 192.450 304.950 ;
        RECT 184.950 274.950 187.050 277.050 ;
        RECT 187.950 275.250 190.050 276.150 ;
        RECT 190.950 274.950 193.050 277.050 ;
        RECT 184.950 272.250 186.750 273.150 ;
        RECT 187.950 271.950 190.050 274.050 ;
        RECT 191.250 272.250 192.750 273.150 ;
        RECT 193.950 271.950 196.050 274.050 ;
        RECT 184.950 268.950 187.050 271.050 ;
        RECT 185.400 265.050 186.450 268.950 ;
        RECT 184.950 262.950 187.050 265.050 ;
        RECT 188.400 259.050 189.450 271.950 ;
        RECT 190.950 268.950 193.050 271.050 ;
        RECT 194.250 269.850 196.050 270.750 ;
        RECT 191.400 262.050 192.450 268.950 ;
        RECT 193.950 265.950 196.050 268.050 ;
        RECT 190.950 259.950 193.050 262.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 253.950 193.050 256.050 ;
        RECT 187.950 250.950 190.050 253.050 ;
        RECT 188.400 247.050 189.450 250.950 ;
        RECT 187.950 244.950 190.050 247.050 ;
        RECT 166.950 235.950 169.050 238.050 ;
        RECT 170.250 236.850 171.750 237.750 ;
        RECT 172.950 235.950 175.050 238.050 ;
        RECT 176.250 236.850 178.050 237.750 ;
        RECT 178.950 235.950 181.050 238.050 ;
        RECT 181.950 235.950 184.050 238.050 ;
        RECT 184.950 235.950 187.050 238.050 ;
        RECT 188.250 236.250 190.050 237.150 ;
        RECT 191.400 235.050 192.450 253.950 ;
        RECT 194.400 253.050 195.450 265.950 ;
        RECT 197.400 256.050 198.450 307.950 ;
        RECT 203.400 306.450 204.450 349.950 ;
        RECT 205.950 341.250 208.050 342.150 ;
        RECT 212.400 340.050 213.450 370.950 ;
        RECT 215.400 364.050 216.450 379.950 ;
        RECT 214.950 361.950 217.050 364.050 ;
        RECT 221.400 355.050 222.450 380.400 ;
        RECT 226.950 380.250 228.750 381.150 ;
        RECT 229.950 379.950 232.050 382.050 ;
        RECT 233.250 380.250 235.050 381.150 ;
        RECT 239.400 379.050 240.450 388.950 ;
        RECT 230.250 377.850 231.750 378.750 ;
        RECT 232.950 376.950 235.050 379.050 ;
        RECT 238.950 376.950 241.050 379.050 ;
        RECT 242.400 372.600 243.600 389.400 ;
        RECT 248.400 385.050 249.450 391.950 ;
        RECT 247.950 382.950 250.050 385.050 ;
        RECT 244.950 379.950 247.050 382.050 ;
        RECT 247.950 380.850 250.050 381.750 ;
        RECT 241.950 370.500 244.050 372.600 ;
        RECT 245.400 358.050 246.450 379.950 ;
        RECT 247.950 376.950 250.050 379.050 ;
        RECT 223.950 355.950 226.050 358.050 ;
        RECT 244.950 355.950 247.050 358.050 ;
        RECT 214.950 351.300 217.050 353.400 ;
        RECT 220.950 352.950 223.050 355.050 ;
        RECT 215.250 347.700 216.450 351.300 ;
        RECT 214.950 345.600 217.050 347.700 ;
        RECT 205.950 337.950 208.050 340.050 ;
        RECT 211.950 337.950 214.050 340.050 ;
        RECT 206.400 331.050 207.450 337.950 ;
        RECT 205.950 328.950 208.050 331.050 ;
        RECT 212.400 316.050 213.450 337.950 ;
        RECT 215.250 333.600 216.450 345.600 ;
        RECT 224.400 342.450 225.450 355.950 ;
        RECT 244.950 350.400 247.050 352.500 ;
        RECT 226.950 344.250 229.050 345.150 ;
        RECT 226.950 342.450 229.050 343.050 ;
        RECT 224.400 341.400 229.050 342.450 ;
        RECT 226.950 340.950 229.050 341.400 ;
        RECT 230.250 341.250 231.750 342.150 ;
        RECT 232.950 340.950 235.050 343.050 ;
        RECT 236.250 341.250 238.050 342.150 ;
        RECT 241.950 340.950 244.050 343.050 ;
        RECT 217.950 337.950 220.050 340.050 ;
        RECT 229.950 337.950 232.050 340.050 ;
        RECT 233.250 338.850 234.750 339.750 ;
        RECT 235.950 337.950 238.050 340.050 ;
        RECT 217.950 335.850 220.050 336.750 ;
        RECT 230.400 334.050 231.450 337.950 ;
        RECT 236.400 337.050 237.450 337.950 ;
        RECT 235.950 334.950 238.050 337.050 ;
        RECT 214.950 331.500 217.050 333.600 ;
        RECT 229.950 331.950 232.050 334.050 ;
        RECT 211.950 313.950 214.050 316.050 ;
        RECT 214.950 313.950 217.050 316.050 ;
        RECT 205.950 310.950 208.050 313.050 ;
        RECT 215.400 312.450 216.450 313.950 ;
        RECT 212.400 311.400 216.450 312.450 ;
        RECT 206.400 310.050 207.450 310.950 ;
        RECT 212.400 310.050 213.450 311.400 ;
        RECT 232.950 310.950 235.050 313.050 ;
        RECT 233.400 310.050 234.450 310.950 ;
        RECT 205.950 307.950 208.050 310.050 ;
        RECT 208.950 308.250 210.750 309.150 ;
        RECT 211.950 307.950 214.050 310.050 ;
        RECT 215.250 308.250 217.050 309.150 ;
        RECT 220.950 308.250 222.750 309.150 ;
        RECT 223.950 307.950 226.050 310.050 ;
        RECT 227.250 308.250 229.050 309.150 ;
        RECT 229.950 308.250 231.750 309.150 ;
        RECT 232.950 307.950 235.050 310.050 ;
        RECT 236.250 308.250 238.050 309.150 ;
        RECT 203.400 305.400 207.450 306.450 ;
        RECT 202.950 301.950 205.050 304.050 ;
        RECT 203.400 298.050 204.450 301.950 ;
        RECT 202.950 295.950 205.050 298.050 ;
        RECT 202.950 270.450 205.050 271.050 ;
        RECT 206.400 270.450 207.450 305.400 ;
        RECT 208.950 304.950 211.050 307.050 ;
        RECT 212.250 305.850 213.750 306.750 ;
        RECT 214.950 304.950 217.050 307.050 ;
        RECT 220.950 304.950 223.050 307.050 ;
        RECT 224.250 305.850 225.750 306.750 ;
        RECT 226.950 304.950 229.050 307.050 ;
        RECT 229.950 304.950 232.050 307.050 ;
        RECT 233.250 305.850 234.750 306.750 ;
        RECT 235.950 304.950 238.050 307.050 ;
        RECT 209.400 304.050 210.450 304.950 ;
        RECT 221.400 304.050 222.450 304.950 ;
        RECT 208.950 301.950 211.050 304.050 ;
        RECT 220.950 301.950 223.050 304.050 ;
        RECT 227.400 301.050 228.450 304.950 ;
        RECT 236.400 301.050 237.450 304.950 ;
        RECT 226.950 298.950 229.050 301.050 ;
        RECT 235.950 298.950 238.050 301.050 ;
        RECT 214.950 280.950 217.050 283.050 ;
        RECT 215.400 274.050 216.450 280.950 ;
        RECT 229.950 275.250 232.050 276.150 ;
        RECT 236.400 274.050 237.450 298.950 ;
        RECT 242.400 274.050 243.450 340.950 ;
        RECT 245.400 333.600 246.600 350.400 ;
        RECT 248.400 340.050 249.450 376.950 ;
        RECT 251.400 373.050 252.450 394.950 ;
        RECT 254.400 385.050 255.450 400.950 ;
        RECT 253.950 382.950 256.050 385.050 ;
        RECT 253.950 380.850 256.050 381.750 ;
        RECT 250.950 370.950 253.050 373.050 ;
        RECT 257.400 372.450 258.450 446.400 ;
        RECT 269.400 442.050 270.450 448.950 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 268.950 439.950 271.050 442.050 ;
        RECT 262.950 430.950 265.050 433.050 ;
        RECT 259.950 423.300 262.050 425.400 ;
        RECT 260.250 419.700 261.450 423.300 ;
        RECT 263.400 421.050 264.450 430.950 ;
        RECT 259.950 417.600 262.050 419.700 ;
        RECT 262.950 418.950 265.050 421.050 ;
        RECT 265.950 418.950 268.050 421.050 ;
        RECT 260.250 405.600 261.450 417.600 ;
        RECT 262.950 409.950 265.050 412.050 ;
        RECT 262.950 407.850 265.050 408.750 ;
        RECT 259.950 403.500 262.050 405.600 ;
        RECT 266.400 403.050 267.450 418.950 ;
        RECT 275.400 418.050 276.450 445.950 ;
        RECT 274.950 415.950 277.050 418.050 ;
        RECT 277.950 416.250 280.050 417.150 ;
        RECT 268.950 413.250 270.750 414.150 ;
        RECT 271.950 412.950 274.050 415.050 ;
        RECT 275.250 413.250 276.750 414.150 ;
        RECT 277.950 412.950 280.050 415.050 ;
        RECT 268.950 409.950 271.050 412.050 ;
        RECT 272.250 410.850 273.750 411.750 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 277.950 409.950 280.050 412.050 ;
        RECT 265.950 400.950 268.050 403.050 ;
        RECT 262.950 389.400 265.050 391.500 ;
        RECT 269.400 391.050 270.450 409.950 ;
        RECT 278.400 406.050 279.450 409.950 ;
        RECT 277.950 403.950 280.050 406.050 ;
        RECT 274.950 397.950 277.050 400.050 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 254.400 371.400 258.450 372.450 ;
        RECT 250.950 341.250 253.050 342.150 ;
        RECT 247.950 337.950 250.050 340.050 ;
        RECT 250.950 337.950 253.050 340.050 ;
        RECT 251.400 334.050 252.450 337.950 ;
        RECT 244.950 331.500 247.050 333.600 ;
        RECT 250.950 331.950 253.050 334.050 ;
        RECT 254.400 328.050 255.450 371.400 ;
        RECT 256.950 341.250 259.050 342.150 ;
        RECT 256.950 339.450 259.050 340.050 ;
        RECT 260.400 339.450 261.450 382.950 ;
        RECT 263.250 377.400 264.450 389.400 ;
        RECT 268.950 388.950 271.050 391.050 ;
        RECT 265.950 386.250 268.050 387.150 ;
        RECT 265.950 382.950 268.050 385.050 ;
        RECT 262.950 375.300 265.050 377.400 ;
        RECT 263.250 371.700 264.450 375.300 ;
        RECT 262.950 369.600 265.050 371.700 ;
        RECT 266.400 364.050 267.450 382.950 ;
        RECT 275.400 382.050 276.450 397.950 ;
        RECT 271.950 380.250 273.750 381.150 ;
        RECT 274.950 379.950 277.050 382.050 ;
        RECT 278.250 380.250 280.050 381.150 ;
        RECT 271.950 376.950 274.050 379.050 ;
        RECT 275.250 377.850 276.750 378.750 ;
        RECT 277.950 376.950 280.050 379.050 ;
        RECT 272.400 376.050 273.450 376.950 ;
        RECT 271.950 373.950 274.050 376.050 ;
        RECT 278.400 373.050 279.450 376.950 ;
        RECT 268.950 370.950 271.050 373.050 ;
        RECT 277.950 370.950 280.050 373.050 ;
        RECT 281.400 372.450 282.450 451.950 ;
        RECT 283.950 418.950 286.050 421.050 ;
        RECT 284.400 415.050 285.450 418.950 ;
        RECT 290.400 418.050 291.450 451.950 ;
        RECT 296.400 451.050 297.450 451.950 ;
        RECT 295.950 448.950 298.050 451.050 ;
        RECT 310.950 448.950 313.050 451.050 ;
        RECT 322.950 449.850 325.050 450.750 ;
        RECT 301.950 418.950 304.050 421.050 ;
        RECT 307.950 418.950 310.050 421.050 ;
        RECT 289.950 415.950 292.050 418.050 ;
        RECT 295.950 415.950 298.050 418.050 ;
        RECT 296.400 415.050 297.450 415.950 ;
        RECT 302.400 415.050 303.450 418.950 ;
        RECT 283.950 412.950 286.050 415.050 ;
        RECT 286.950 414.450 289.050 415.050 ;
        RECT 289.950 414.450 292.050 415.050 ;
        RECT 286.950 413.400 292.050 414.450 ;
        RECT 286.950 412.950 289.050 413.400 ;
        RECT 289.950 412.950 292.050 413.400 ;
        RECT 292.950 413.250 294.750 414.150 ;
        RECT 295.950 412.950 298.050 415.050 ;
        RECT 299.250 413.250 300.750 414.150 ;
        RECT 301.950 412.950 304.050 415.050 ;
        RECT 305.250 413.250 307.050 414.150 ;
        RECT 283.950 410.250 286.050 411.150 ;
        RECT 286.950 410.850 289.050 411.750 ;
        RECT 290.400 411.450 291.450 412.950 ;
        RECT 292.950 411.450 295.050 412.050 ;
        RECT 290.400 410.400 295.050 411.450 ;
        RECT 296.250 410.850 297.750 411.750 ;
        RECT 292.950 409.950 295.050 410.400 ;
        RECT 298.950 409.950 301.050 412.050 ;
        RECT 302.250 410.850 303.750 411.750 ;
        RECT 304.950 409.950 307.050 412.050 ;
        RECT 283.950 406.950 286.050 409.050 ;
        RECT 289.950 406.950 292.050 409.050 ;
        RECT 286.950 400.950 289.050 403.050 ;
        RECT 287.400 382.050 288.450 400.950 ;
        RECT 290.400 385.050 291.450 406.950 ;
        RECT 292.950 403.950 295.050 406.050 ;
        RECT 289.950 382.950 292.050 385.050 ;
        RECT 283.950 380.250 285.750 381.150 ;
        RECT 286.950 379.950 289.050 382.050 ;
        RECT 290.250 380.250 292.050 381.150 ;
        RECT 283.950 376.950 286.050 379.050 ;
        RECT 287.250 377.850 288.750 378.750 ;
        RECT 289.950 376.950 292.050 379.050 ;
        RECT 284.400 376.050 285.450 376.950 ;
        RECT 283.950 373.950 286.050 376.050 ;
        RECT 281.400 371.400 285.450 372.450 ;
        RECT 265.950 361.950 268.050 364.050 ;
        RECT 265.950 351.300 268.050 353.400 ;
        RECT 266.250 347.700 267.450 351.300 ;
        RECT 265.950 345.600 268.050 347.700 ;
        RECT 256.950 338.400 261.450 339.450 ;
        RECT 256.950 337.950 259.050 338.400 ;
        RECT 257.400 331.050 258.450 337.950 ;
        RECT 266.250 333.600 267.450 345.600 ;
        RECT 269.400 340.050 270.450 370.950 ;
        RECT 271.950 367.950 274.050 370.050 ;
        RECT 268.950 337.950 271.050 340.050 ;
        RECT 268.950 335.850 271.050 336.750 ;
        RECT 265.950 331.500 268.050 333.600 ;
        RECT 272.400 331.050 273.450 367.950 ;
        RECT 277.950 342.450 280.050 343.050 ;
        RECT 275.400 341.400 280.050 342.450 ;
        RECT 275.400 337.050 276.450 341.400 ;
        RECT 277.950 340.950 280.050 341.400 ;
        RECT 277.950 338.850 280.050 339.750 ;
        RECT 280.950 338.250 283.050 339.150 ;
        RECT 274.950 334.950 277.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 281.400 334.050 282.450 334.950 ;
        RECT 280.950 331.950 283.050 334.050 ;
        RECT 256.950 328.950 259.050 331.050 ;
        RECT 271.950 328.950 274.050 331.050 ;
        RECT 244.950 325.950 247.050 328.050 ;
        RECT 253.950 325.950 256.050 328.050 ;
        RECT 265.950 325.950 268.050 328.050 ;
        RECT 245.400 310.050 246.450 325.950 ;
        RECT 253.950 322.950 256.050 325.050 ;
        RECT 247.950 316.950 250.050 319.050 ;
        RECT 248.400 313.050 249.450 316.950 ;
        RECT 254.400 313.050 255.450 322.950 ;
        RECT 262.950 319.950 265.050 322.050 ;
        RECT 263.400 316.050 264.450 319.950 ;
        RECT 259.950 313.950 262.050 316.050 ;
        RECT 262.950 313.950 265.050 316.050 ;
        RECT 266.400 313.050 267.450 325.950 ;
        RECT 271.950 322.950 274.050 325.050 ;
        RECT 274.950 322.950 277.050 325.050 ;
        RECT 280.950 322.950 283.050 325.050 ;
        RECT 272.400 313.050 273.450 322.950 ;
        RECT 275.400 316.050 276.450 322.950 ;
        RECT 274.950 313.950 277.050 316.050 ;
        RECT 277.950 313.950 280.050 316.050 ;
        RECT 278.400 313.050 279.450 313.950 ;
        RECT 247.950 310.950 250.050 313.050 ;
        RECT 251.250 311.250 252.750 312.150 ;
        RECT 253.950 310.950 256.050 313.050 ;
        RECT 256.950 311.250 259.050 312.150 ;
        RECT 259.950 311.850 262.050 312.750 ;
        RECT 262.950 311.250 264.750 312.150 ;
        RECT 265.950 310.950 268.050 313.050 ;
        RECT 271.950 310.950 274.050 313.050 ;
        RECT 275.250 311.850 276.750 312.750 ;
        RECT 277.950 310.950 280.050 313.050 ;
        RECT 244.950 307.950 247.050 310.050 ;
        RECT 248.250 308.850 249.750 309.750 ;
        RECT 250.950 307.950 253.050 310.050 ;
        RECT 254.250 308.850 256.050 309.750 ;
        RECT 256.950 307.950 259.050 310.050 ;
        RECT 259.950 307.950 262.050 310.050 ;
        RECT 262.950 307.950 265.050 310.050 ;
        RECT 266.250 308.850 268.050 309.750 ;
        RECT 271.950 308.850 274.050 309.750 ;
        RECT 277.950 308.850 280.050 309.750 ;
        RECT 244.950 305.850 247.050 306.750 ;
        RECT 247.950 295.950 250.050 298.050 ;
        RECT 214.950 271.950 217.050 274.050 ;
        RECT 226.950 272.250 228.750 273.150 ;
        RECT 229.950 271.950 232.050 274.050 ;
        RECT 233.250 272.250 234.750 273.150 ;
        RECT 235.950 271.950 238.050 274.050 ;
        RECT 241.950 271.950 244.050 274.050 ;
        RECT 215.400 271.050 216.450 271.950 ;
        RECT 200.400 269.400 207.450 270.450 ;
        RECT 196.950 253.950 199.050 256.050 ;
        RECT 193.950 250.950 196.050 253.050 ;
        RECT 200.400 244.050 201.450 269.400 ;
        RECT 202.950 268.950 205.050 269.400 ;
        RECT 211.950 269.250 213.750 270.150 ;
        RECT 214.950 268.950 217.050 271.050 ;
        RECT 218.250 269.250 219.750 270.150 ;
        RECT 220.950 268.950 223.050 271.050 ;
        RECT 224.250 269.250 226.050 270.150 ;
        RECT 226.950 268.950 229.050 271.050 ;
        RECT 229.950 268.950 232.050 271.050 ;
        RECT 232.950 268.950 235.050 271.050 ;
        RECT 236.250 269.850 238.050 270.750 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 227.400 268.050 228.450 268.950 ;
        RECT 202.950 266.850 205.050 267.750 ;
        RECT 205.950 266.250 208.050 267.150 ;
        RECT 211.950 265.950 214.050 268.050 ;
        RECT 215.250 266.850 216.750 267.750 ;
        RECT 217.950 265.950 220.050 268.050 ;
        RECT 221.250 266.850 222.750 267.750 ;
        RECT 223.950 265.950 226.050 268.050 ;
        RECT 226.950 265.950 229.050 268.050 ;
        RECT 205.950 262.950 208.050 265.050 ;
        RECT 206.400 259.050 207.450 262.950 ;
        RECT 218.400 262.050 219.450 265.950 ;
        RECT 224.400 265.050 225.450 265.950 ;
        RECT 223.950 262.950 226.050 265.050 ;
        RECT 217.950 259.950 220.050 262.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 202.950 247.950 205.050 250.050 ;
        RECT 196.950 241.950 199.050 244.050 ;
        RECT 199.950 241.950 202.050 244.050 ;
        RECT 203.400 241.050 204.450 247.950 ;
        RECT 230.400 247.050 231.450 268.950 ;
        RECT 241.950 266.250 244.050 267.150 ;
        RECT 244.950 266.850 247.050 267.750 ;
        RECT 241.950 262.950 244.050 265.050 ;
        RECT 244.950 262.950 247.050 265.050 ;
        RECT 242.400 253.050 243.450 262.950 ;
        RECT 241.950 250.950 244.050 253.050 ;
        RECT 220.950 244.950 223.050 247.050 ;
        RECT 229.950 244.950 232.050 247.050 ;
        RECT 235.950 244.950 238.050 247.050 ;
        RECT 205.950 241.950 208.050 244.050 ;
        RECT 214.950 243.450 217.050 244.050 ;
        RECT 214.950 242.400 219.450 243.450 ;
        RECT 214.950 241.950 217.050 242.400 ;
        RECT 193.950 239.250 196.050 240.150 ;
        RECT 196.950 239.850 199.050 240.750 ;
        RECT 199.950 239.250 201.750 240.150 ;
        RECT 202.950 238.950 205.050 241.050 ;
        RECT 193.950 237.450 196.050 238.050 ;
        RECT 193.950 236.400 198.450 237.450 ;
        RECT 193.950 235.950 196.050 236.400 ;
        RECT 163.950 232.950 166.050 235.050 ;
        RECT 166.950 233.850 169.050 234.750 ;
        RECT 172.950 232.950 175.050 235.050 ;
        RECT 175.950 232.950 178.050 235.050 ;
        RECT 178.950 233.850 180.750 234.750 ;
        RECT 181.950 232.950 184.050 235.050 ;
        RECT 185.250 233.850 186.750 234.750 ;
        RECT 187.950 232.950 190.050 235.050 ;
        RECT 190.950 232.950 193.050 235.050 ;
        RECT 193.950 232.950 196.050 235.050 ;
        RECT 158.400 230.400 162.450 231.450 ;
        RECT 149.400 226.050 150.450 229.950 ;
        RECT 148.950 223.950 151.050 226.050 ;
        RECT 155.400 217.050 156.450 229.950 ;
        RECT 154.950 214.950 157.050 217.050 ;
        RECT 145.950 202.950 148.050 205.050 ;
        RECT 136.950 199.950 139.050 202.050 ;
        RECT 140.250 200.250 141.750 201.150 ;
        RECT 142.950 199.950 145.050 202.050 ;
        RECT 145.950 199.950 148.050 202.050 ;
        RECT 149.250 200.250 150.750 201.150 ;
        RECT 151.950 199.950 154.050 202.050 ;
        RECT 154.950 199.950 157.050 202.050 ;
        RECT 136.950 197.850 138.750 198.750 ;
        RECT 139.950 196.950 142.050 199.050 ;
        RECT 143.250 197.850 145.050 198.750 ;
        RECT 145.950 197.850 147.750 198.750 ;
        RECT 148.950 196.950 151.050 199.050 ;
        RECT 152.250 197.850 154.050 198.750 ;
        RECT 136.950 193.950 139.050 196.050 ;
        RECT 137.400 193.050 138.450 193.950 ;
        RECT 149.400 193.050 150.450 196.950 ;
        RECT 136.950 190.950 139.050 193.050 ;
        RECT 148.950 190.950 151.050 193.050 ;
        RECT 133.950 181.950 136.050 184.050 ;
        RECT 137.400 166.050 138.450 190.950 ;
        RECT 148.950 187.950 151.050 190.050 ;
        RECT 149.400 181.050 150.450 187.950 ;
        RECT 148.950 178.950 151.050 181.050 ;
        RECT 145.950 172.950 148.050 175.050 ;
        RECT 146.400 169.050 147.450 172.950 ;
        RECT 149.400 169.050 150.450 178.950 ;
        RECT 155.400 178.050 156.450 199.950 ;
        RECT 158.400 190.050 159.450 230.400 ;
        RECT 163.950 229.950 166.050 232.050 ;
        RECT 164.400 205.050 165.450 229.950 ;
        RECT 163.950 202.950 166.050 205.050 ;
        RECT 166.950 203.250 169.050 204.150 ;
        RECT 160.950 199.950 163.050 202.050 ;
        RECT 164.250 200.250 165.750 201.150 ;
        RECT 166.950 199.950 169.050 202.050 ;
        RECT 170.250 200.250 172.050 201.150 ;
        RECT 160.950 197.850 162.750 198.750 ;
        RECT 163.950 196.950 166.050 199.050 ;
        RECT 166.950 196.950 169.050 199.050 ;
        RECT 169.950 196.950 172.050 199.050 ;
        RECT 163.950 193.950 166.050 196.050 ;
        RECT 157.950 187.950 160.050 190.050 ;
        RECT 157.950 178.950 160.050 181.050 ;
        RECT 154.950 175.950 157.050 178.050 ;
        RECT 154.950 169.950 157.050 172.050 ;
        RECT 155.400 169.050 156.450 169.950 ;
        RECT 139.950 166.950 142.050 169.050 ;
        RECT 143.250 167.250 144.750 168.150 ;
        RECT 145.950 166.950 148.050 169.050 ;
        RECT 148.950 166.950 151.050 169.050 ;
        RECT 152.250 167.250 153.750 168.150 ;
        RECT 154.950 166.950 157.050 169.050 ;
        RECT 158.400 168.450 159.450 178.950 ;
        RECT 164.400 175.050 165.450 193.950 ;
        RECT 163.950 172.950 166.050 175.050 ;
        RECT 158.400 167.400 162.450 168.450 ;
        RECT 121.950 164.250 123.750 165.150 ;
        RECT 124.950 163.950 127.050 166.050 ;
        RECT 127.950 163.950 130.050 166.050 ;
        RECT 130.950 163.950 133.050 166.050 ;
        RECT 136.950 163.950 139.050 166.050 ;
        RECT 140.250 164.850 141.750 165.750 ;
        RECT 142.950 163.950 145.050 166.050 ;
        RECT 146.250 164.850 148.050 165.750 ;
        RECT 148.950 164.850 150.750 165.750 ;
        RECT 151.950 163.950 154.050 166.050 ;
        RECT 155.250 164.850 156.750 165.750 ;
        RECT 157.950 163.950 160.050 166.050 ;
        RECT 128.400 163.050 129.450 163.950 ;
        RECT 143.400 163.050 144.450 163.950 ;
        RECT 121.950 160.950 124.050 163.050 ;
        RECT 125.250 161.850 126.750 162.750 ;
        RECT 127.950 160.950 130.050 163.050 ;
        RECT 131.250 161.850 133.050 162.750 ;
        RECT 136.950 161.850 139.050 162.750 ;
        RECT 142.950 160.950 145.050 163.050 ;
        RECT 122.400 154.050 123.450 160.950 ;
        RECT 127.950 158.850 130.050 159.750 ;
        RECT 130.950 157.950 133.050 160.050 ;
        RECT 121.950 151.950 124.050 154.050 ;
        RECT 124.950 145.950 127.050 148.050 ;
        RECT 121.950 136.950 124.050 139.050 ;
        RECT 122.400 106.050 123.450 136.950 ;
        RECT 125.400 130.050 126.450 145.950 ;
        RECT 127.950 133.950 130.050 136.050 ;
        RECT 128.400 130.050 129.450 133.950 ;
        RECT 124.950 127.950 127.050 130.050 ;
        RECT 127.950 127.950 130.050 130.050 ;
        RECT 124.950 125.250 127.050 126.150 ;
        RECT 127.950 125.850 130.050 126.750 ;
        RECT 124.950 121.950 127.050 124.050 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 121.950 103.950 124.050 106.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 128.400 97.050 129.450 121.950 ;
        RECT 131.400 118.050 132.450 157.950 ;
        RECT 133.950 154.950 136.050 157.050 ;
        RECT 134.400 148.050 135.450 154.950 ;
        RECT 133.950 145.950 136.050 148.050 ;
        RECT 148.950 142.950 151.050 145.050 ;
        RECT 133.950 139.950 136.050 142.050 ;
        RECT 134.400 130.050 135.450 139.950 ;
        RECT 136.950 133.950 139.050 136.050 ;
        RECT 137.400 130.050 138.450 133.950 ;
        RECT 133.950 127.950 136.050 130.050 ;
        RECT 136.950 127.950 139.050 130.050 ;
        RECT 140.250 128.250 141.750 129.150 ;
        RECT 142.950 127.950 145.050 130.050 ;
        RECT 145.950 127.950 148.050 130.050 ;
        RECT 133.950 125.250 136.050 126.150 ;
        RECT 136.950 125.850 138.750 126.750 ;
        RECT 139.950 124.950 142.050 127.050 ;
        RECT 143.250 125.850 145.050 126.750 ;
        RECT 133.950 121.950 136.050 124.050 ;
        RECT 140.400 121.050 141.450 124.950 ;
        RECT 146.400 124.050 147.450 127.950 ;
        RECT 145.950 121.950 148.050 124.050 ;
        RECT 139.950 118.950 142.050 121.050 ;
        RECT 130.950 115.950 133.050 118.050 ;
        RECT 149.400 109.050 150.450 142.950 ;
        RECT 152.400 139.050 153.450 163.950 ;
        RECT 157.950 161.850 160.050 162.750 ;
        RECT 161.400 145.050 162.450 167.400 ;
        RECT 160.950 142.950 163.050 145.050 ;
        RECT 160.950 139.950 163.050 142.050 ;
        RECT 151.950 136.950 154.050 139.050 ;
        RECT 161.400 133.050 162.450 139.950 ;
        RECT 157.950 131.250 160.050 132.150 ;
        RECT 160.950 130.950 163.050 133.050 ;
        RECT 164.400 130.050 165.450 172.950 ;
        RECT 167.400 172.050 168.450 196.950 ;
        RECT 170.400 181.050 171.450 196.950 ;
        RECT 173.400 196.050 174.450 232.950 ;
        RECT 176.400 217.050 177.450 232.950 ;
        RECT 188.400 232.050 189.450 232.950 ;
        RECT 178.950 229.950 181.050 232.050 ;
        RECT 181.950 230.850 184.050 231.750 ;
        RECT 184.950 229.950 187.050 232.050 ;
        RECT 187.950 229.950 190.050 232.050 ;
        RECT 179.400 223.050 180.450 229.950 ;
        RECT 185.400 226.050 186.450 229.950 ;
        RECT 194.400 229.050 195.450 232.950 ;
        RECT 193.950 226.950 196.050 229.050 ;
        RECT 197.400 226.050 198.450 236.400 ;
        RECT 199.950 235.950 202.050 238.050 ;
        RECT 203.250 236.850 205.050 237.750 ;
        RECT 199.950 232.950 202.050 235.050 ;
        RECT 184.950 223.950 187.050 226.050 ;
        RECT 196.950 223.950 199.050 226.050 ;
        RECT 178.950 220.950 181.050 223.050 ;
        RECT 175.950 214.950 178.050 217.050 ;
        RECT 178.950 205.950 181.050 208.050 ;
        RECT 175.950 199.950 178.050 202.050 ;
        RECT 176.400 199.050 177.450 199.950 ;
        RECT 179.400 199.050 180.450 205.950 ;
        RECT 181.950 202.950 184.050 205.050 ;
        RECT 175.950 196.950 178.050 199.050 ;
        RECT 178.950 196.950 181.050 199.050 ;
        RECT 172.950 193.950 175.050 196.050 ;
        RECT 175.950 194.850 178.050 195.750 ;
        RECT 178.950 194.250 181.050 195.150 ;
        RECT 178.950 190.950 181.050 193.050 ;
        RECT 179.400 187.050 180.450 190.950 ;
        RECT 178.950 184.950 181.050 187.050 ;
        RECT 179.400 184.050 180.450 184.950 ;
        RECT 178.950 181.950 181.050 184.050 ;
        RECT 169.950 178.950 172.050 181.050 ;
        RECT 182.400 178.050 183.450 202.950 ;
        RECT 190.950 199.950 193.050 202.050 ;
        RECT 184.950 197.250 187.050 198.150 ;
        RECT 187.950 197.850 190.050 198.750 ;
        RECT 184.950 193.950 187.050 196.050 ;
        RECT 187.950 193.950 190.050 196.050 ;
        RECT 175.950 175.950 178.050 178.050 ;
        RECT 181.950 175.950 184.050 178.050 ;
        RECT 169.950 172.950 172.050 175.050 ;
        RECT 166.950 169.950 169.050 172.050 ;
        RECT 170.400 169.050 171.450 172.950 ;
        RECT 176.400 169.050 177.450 175.950 ;
        RECT 178.950 172.950 181.050 175.050 ;
        RECT 166.950 166.950 169.050 169.050 ;
        RECT 169.950 166.950 172.050 169.050 ;
        RECT 173.250 167.250 174.750 168.150 ;
        RECT 175.950 166.950 178.050 169.050 ;
        RECT 167.400 166.050 168.450 166.950 ;
        RECT 166.950 163.950 169.050 166.050 ;
        RECT 170.250 164.850 171.750 165.750 ;
        RECT 172.950 163.950 175.050 166.050 ;
        RECT 176.250 164.850 178.050 165.750 ;
        RECT 173.400 163.050 174.450 163.950 ;
        RECT 166.950 161.850 169.050 162.750 ;
        RECT 172.950 160.950 175.050 163.050 ;
        RECT 173.400 148.050 174.450 160.950 ;
        RECT 172.950 145.950 175.050 148.050 ;
        RECT 175.950 142.950 178.050 145.050 ;
        RECT 166.950 136.950 169.050 139.050 ;
        RECT 167.400 130.050 168.450 136.950 ;
        RECT 151.950 127.950 154.050 130.050 ;
        RECT 155.250 128.250 156.750 129.150 ;
        RECT 157.950 127.950 160.050 130.050 ;
        RECT 161.250 128.250 163.050 129.150 ;
        RECT 163.950 127.950 166.050 130.050 ;
        RECT 166.950 127.950 169.050 130.050 ;
        RECT 172.950 128.250 175.050 129.150 ;
        RECT 167.400 127.050 168.450 127.950 ;
        RECT 151.950 125.850 153.750 126.750 ;
        RECT 154.950 124.950 157.050 127.050 ;
        RECT 157.950 124.950 160.050 127.050 ;
        RECT 160.950 124.950 163.050 127.050 ;
        RECT 163.950 125.250 165.750 126.150 ;
        RECT 166.950 124.950 169.050 127.050 ;
        RECT 172.950 126.450 175.050 127.050 ;
        RECT 176.400 126.450 177.450 142.950 ;
        RECT 179.400 142.050 180.450 172.950 ;
        RECT 185.400 172.050 186.450 193.950 ;
        RECT 188.400 190.050 189.450 193.950 ;
        RECT 187.950 187.950 190.050 190.050 ;
        RECT 184.950 169.950 187.050 172.050 ;
        RECT 181.950 164.250 183.750 165.150 ;
        RECT 184.950 163.950 187.050 166.050 ;
        RECT 188.250 164.250 190.050 165.150 ;
        RECT 181.950 160.950 184.050 163.050 ;
        RECT 185.250 161.850 186.750 162.750 ;
        RECT 187.950 160.950 190.050 163.050 ;
        RECT 188.400 145.050 189.450 160.950 ;
        RECT 187.950 142.950 190.050 145.050 ;
        RECT 178.950 139.950 181.050 142.050 ;
        RECT 178.950 136.950 181.050 139.050 ;
        RECT 179.400 127.050 180.450 136.950 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 182.400 133.050 183.450 133.950 ;
        RECT 191.400 133.050 192.450 199.950 ;
        RECT 200.400 199.050 201.450 232.950 ;
        RECT 206.400 205.050 207.450 241.950 ;
        RECT 211.950 239.250 214.050 240.150 ;
        RECT 214.950 239.850 217.050 240.750 ;
        RECT 218.400 238.050 219.450 242.400 ;
        RECT 211.950 235.950 214.050 238.050 ;
        RECT 217.950 237.450 220.050 238.050 ;
        RECT 215.400 236.400 220.050 237.450 ;
        RECT 211.950 232.950 214.050 235.050 ;
        RECT 212.400 223.050 213.450 232.950 ;
        RECT 215.400 226.050 216.450 236.400 ;
        RECT 217.950 235.950 220.050 236.400 ;
        RECT 221.400 235.050 222.450 244.950 ;
        RECT 236.400 244.050 237.450 244.950 ;
        RECT 235.950 241.950 238.050 244.050 ;
        RECT 232.950 239.250 235.050 240.150 ;
        RECT 235.950 239.850 238.050 240.750 ;
        RECT 238.950 239.250 240.750 240.150 ;
        RECT 241.950 238.950 244.050 241.050 ;
        RECT 223.950 235.950 226.050 238.050 ;
        RECT 227.250 236.250 229.050 237.150 ;
        RECT 232.950 235.950 235.050 238.050 ;
        RECT 235.950 235.950 238.050 238.050 ;
        RECT 238.950 235.950 241.050 238.050 ;
        RECT 242.250 236.850 244.050 237.750 ;
        RECT 245.400 237.450 246.450 262.950 ;
        RECT 248.400 262.050 249.450 295.950 ;
        RECT 257.400 286.050 258.450 307.950 ;
        RECT 260.400 304.050 261.450 307.950 ;
        RECT 259.950 301.950 262.050 304.050 ;
        RECT 281.400 301.050 282.450 322.950 ;
        RECT 284.400 319.050 285.450 371.400 ;
        RECT 290.400 364.050 291.450 376.950 ;
        RECT 293.400 373.050 294.450 403.950 ;
        RECT 305.400 403.050 306.450 409.950 ;
        RECT 308.400 406.050 309.450 418.950 ;
        RECT 307.950 403.950 310.050 406.050 ;
        RECT 304.950 400.950 307.050 403.050 ;
        RECT 311.400 397.050 312.450 448.950 ;
        RECT 332.400 418.050 333.450 451.950 ;
        RECT 338.400 427.050 339.450 458.400 ;
        RECT 337.950 424.950 340.050 427.050 ;
        RECT 334.950 418.950 337.050 421.050 ;
        RECT 331.950 415.950 334.050 418.050 ;
        RECT 313.950 413.250 316.050 414.150 ;
        RECT 319.950 413.250 322.050 414.150 ;
        RECT 322.950 412.950 325.050 415.050 ;
        RECT 325.950 413.250 328.050 414.150 ;
        RECT 331.950 413.250 334.050 414.150 ;
        RECT 313.950 409.950 316.050 412.050 ;
        RECT 317.250 410.250 318.750 411.150 ;
        RECT 319.950 409.950 322.050 412.050 ;
        RECT 323.400 411.450 324.450 412.950 ;
        RECT 325.950 411.450 328.050 412.050 ;
        RECT 323.400 410.400 328.050 411.450 ;
        RECT 331.950 411.450 334.050 412.050 ;
        RECT 335.400 411.450 336.450 418.950 ;
        RECT 341.400 415.050 342.450 460.950 ;
        RECT 344.400 457.050 345.450 485.400 ;
        RECT 346.950 484.950 349.050 485.400 ;
        RECT 349.950 484.950 352.050 487.050 ;
        RECT 352.950 485.850 354.750 486.750 ;
        RECT 355.950 484.950 358.050 487.050 ;
        RECT 359.250 485.850 361.050 486.750 ;
        RECT 346.950 482.850 349.050 483.750 ;
        RECT 349.950 482.250 352.050 483.150 ;
        RECT 349.950 478.950 352.050 481.050 ;
        RECT 356.400 472.050 357.450 484.950 ;
        RECT 358.950 481.950 361.050 484.050 ;
        RECT 355.950 469.950 358.050 472.050 ;
        RECT 352.950 463.950 355.050 466.050 ;
        RECT 353.400 457.050 354.450 463.950 ;
        RECT 359.400 457.050 360.450 481.950 ;
        RECT 343.950 454.950 346.050 457.050 ;
        RECT 352.950 454.950 355.050 457.050 ;
        RECT 356.250 455.250 357.750 456.150 ;
        RECT 358.950 454.950 361.050 457.050 ;
        RECT 362.400 456.450 363.450 530.400 ;
        RECT 364.950 529.950 367.050 532.050 ;
        RECT 367.950 530.250 370.050 531.150 ;
        RECT 365.400 528.450 366.450 529.950 ;
        RECT 367.950 528.450 370.050 529.050 ;
        RECT 365.400 527.400 370.050 528.450 ;
        RECT 365.400 460.050 366.450 527.400 ;
        RECT 367.950 526.950 370.050 527.400 ;
        RECT 371.550 521.400 372.750 533.400 ;
        RECT 370.950 519.300 373.050 521.400 ;
        RECT 371.550 515.700 372.750 519.300 ;
        RECT 370.950 513.600 373.050 515.700 ;
        RECT 370.950 495.300 373.050 497.400 ;
        RECT 371.550 491.700 372.750 495.300 ;
        RECT 370.950 489.600 373.050 491.700 ;
        RECT 367.950 481.950 370.050 484.050 ;
        RECT 367.950 479.850 370.050 480.750 ;
        RECT 367.950 475.950 370.050 478.050 ;
        RECT 371.550 477.600 372.750 489.600 ;
        RECT 368.400 463.050 369.450 475.950 ;
        RECT 370.950 475.500 373.050 477.600 ;
        RECT 367.950 460.950 370.050 463.050 ;
        RECT 368.400 460.050 369.450 460.950 ;
        RECT 364.950 457.950 367.050 460.050 ;
        RECT 367.950 457.950 370.050 460.050 ;
        RECT 362.400 455.400 366.450 456.450 ;
        RECT 367.950 455.850 370.050 456.750 ;
        RECT 343.950 452.250 345.750 453.150 ;
        RECT 346.950 451.950 349.050 454.050 ;
        RECT 350.250 452.250 352.050 453.150 ;
        RECT 352.950 452.850 354.750 453.750 ;
        RECT 355.950 451.950 358.050 454.050 ;
        RECT 359.250 452.850 360.750 453.750 ;
        RECT 361.950 451.950 364.050 454.050 ;
        RECT 343.950 448.950 346.050 451.050 ;
        RECT 347.250 449.850 348.750 450.750 ;
        RECT 349.950 448.950 352.050 451.050 ;
        RECT 358.950 448.950 361.050 451.050 ;
        RECT 361.950 449.850 364.050 450.750 ;
        RECT 359.400 447.450 360.450 448.950 ;
        RECT 359.400 446.400 363.450 447.450 ;
        RECT 352.950 415.950 355.050 418.050 ;
        RECT 337.950 413.250 340.050 414.150 ;
        RECT 340.950 412.950 343.050 415.050 ;
        RECT 343.950 413.250 346.050 414.150 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 325.950 409.950 328.050 410.400 ;
        RECT 329.250 410.250 330.750 411.150 ;
        RECT 331.950 410.400 336.450 411.450 ;
        RECT 331.950 409.950 334.050 410.400 ;
        RECT 337.950 409.950 340.050 412.050 ;
        RECT 341.250 410.250 342.750 411.150 ;
        RECT 343.950 409.950 346.050 412.050 ;
        RECT 346.950 410.250 349.050 411.150 ;
        RECT 349.950 410.850 352.050 411.750 ;
        RECT 314.400 409.050 315.450 409.950 ;
        RECT 338.400 409.050 339.450 409.950 ;
        RECT 313.950 406.950 316.050 409.050 ;
        RECT 316.950 406.950 319.050 409.050 ;
        RECT 328.950 406.950 331.050 409.050 ;
        RECT 337.950 406.950 340.050 409.050 ;
        RECT 340.950 406.950 343.050 409.050 ;
        RECT 317.400 403.050 318.450 406.950 ;
        RECT 341.400 406.050 342.450 406.950 ;
        RECT 340.950 403.950 343.050 406.050 ;
        RECT 344.400 403.050 345.450 409.950 ;
        RECT 346.950 406.950 349.050 409.050 ;
        RECT 313.950 400.950 316.050 403.050 ;
        RECT 316.950 400.950 319.050 403.050 ;
        RECT 343.950 400.950 346.050 403.050 ;
        RECT 310.950 394.950 313.050 397.050 ;
        RECT 314.400 388.050 315.450 400.950 ;
        RECT 340.950 397.950 343.050 400.050 ;
        RECT 328.950 394.950 331.050 397.050 ;
        RECT 329.400 388.050 330.450 394.950 ;
        RECT 295.950 385.950 298.050 388.050 ;
        RECT 310.950 385.950 313.050 388.050 ;
        RECT 313.950 385.950 316.050 388.050 ;
        RECT 319.950 385.950 322.050 388.050 ;
        RECT 328.950 385.950 331.050 388.050 ;
        RECT 337.950 385.950 340.050 388.050 ;
        RECT 296.400 382.050 297.450 385.950 ;
        RECT 311.400 385.050 312.450 385.950 ;
        RECT 310.950 382.950 313.050 385.050 ;
        RECT 314.250 383.850 315.750 384.750 ;
        RECT 316.950 382.950 319.050 385.050 ;
        RECT 295.950 379.950 298.050 382.050 ;
        RECT 301.950 379.950 304.050 382.050 ;
        RECT 305.250 380.250 307.050 381.150 ;
        RECT 310.950 380.850 313.050 381.750 ;
        RECT 313.950 379.950 316.050 382.050 ;
        RECT 316.950 380.850 319.050 381.750 ;
        RECT 295.950 377.850 297.750 378.750 ;
        RECT 298.950 376.950 301.050 379.050 ;
        RECT 302.250 377.850 303.750 378.750 ;
        RECT 304.950 376.950 307.050 379.050 ;
        RECT 307.950 376.950 310.050 379.050 ;
        RECT 305.400 376.050 306.450 376.950 ;
        RECT 298.950 374.850 301.050 375.750 ;
        RECT 304.950 373.950 307.050 376.050 ;
        RECT 292.950 370.950 295.050 373.050 ;
        RECT 304.950 370.950 307.050 373.050 ;
        RECT 289.950 361.950 292.050 364.050 ;
        RECT 295.950 343.950 298.050 346.050 ;
        RECT 301.950 344.250 304.050 345.150 ;
        RECT 296.400 343.050 297.450 343.950 ;
        RECT 286.950 340.950 289.050 343.050 ;
        RECT 292.950 341.250 294.750 342.150 ;
        RECT 295.950 340.950 298.050 343.050 ;
        RECT 299.250 341.250 300.750 342.150 ;
        RECT 301.950 340.950 304.050 343.050 ;
        RECT 286.950 338.850 289.050 339.750 ;
        RECT 289.950 338.250 292.050 339.150 ;
        RECT 292.950 337.950 295.050 340.050 ;
        RECT 296.250 338.850 297.750 339.750 ;
        RECT 298.950 339.450 301.050 340.050 ;
        RECT 305.400 339.450 306.450 370.950 ;
        RECT 298.950 338.400 306.450 339.450 ;
        RECT 298.950 337.950 301.050 338.400 ;
        RECT 286.950 334.950 289.050 337.050 ;
        RECT 289.950 334.950 292.050 337.050 ;
        RECT 293.400 336.450 294.450 337.950 ;
        RECT 293.400 335.400 297.450 336.450 ;
        RECT 287.400 319.050 288.450 334.950 ;
        RECT 290.400 331.050 291.450 334.950 ;
        RECT 292.950 331.950 295.050 334.050 ;
        RECT 289.950 328.950 292.050 331.050 ;
        RECT 290.400 325.050 291.450 328.950 ;
        RECT 289.950 322.950 292.050 325.050 ;
        RECT 283.950 316.950 286.050 319.050 ;
        RECT 286.950 316.950 289.050 319.050 ;
        RECT 287.400 313.050 288.450 316.950 ;
        RECT 293.400 316.050 294.450 331.950 ;
        RECT 296.400 319.050 297.450 335.400 ;
        RECT 298.950 325.950 301.050 328.050 ;
        RECT 295.950 316.950 298.050 319.050 ;
        RECT 289.950 313.950 292.050 316.050 ;
        RECT 292.950 313.950 295.050 316.050 ;
        RECT 290.400 313.050 291.450 313.950 ;
        RECT 296.400 313.050 297.450 316.950 ;
        RECT 299.400 313.050 300.450 325.950 ;
        RECT 308.400 322.050 309.450 376.950 ;
        RECT 314.400 370.050 315.450 379.950 ;
        RECT 320.400 378.450 321.450 385.950 ;
        RECT 341.400 385.050 342.450 397.950 ;
        RECT 343.950 394.950 346.050 397.050 ;
        RECT 325.950 383.250 328.050 384.150 ;
        RECT 328.950 383.850 331.050 384.750 ;
        RECT 334.950 384.450 337.050 385.050 ;
        RECT 332.400 383.400 337.050 384.450 ;
        RECT 338.250 383.850 339.750 384.750 ;
        RECT 332.400 382.050 333.450 383.400 ;
        RECT 334.950 382.950 337.050 383.400 ;
        RECT 340.950 382.950 343.050 385.050 ;
        RECT 325.950 379.950 328.050 382.050 ;
        RECT 328.950 379.950 331.050 382.050 ;
        RECT 331.950 379.950 334.050 382.050 ;
        RECT 334.950 380.850 337.050 381.750 ;
        RECT 340.950 380.850 343.050 381.750 ;
        RECT 317.400 377.400 321.450 378.450 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 313.950 350.400 316.050 352.500 ;
        RECT 310.950 343.950 313.050 346.050 ;
        RECT 307.950 319.950 310.050 322.050 ;
        RECT 307.950 316.950 310.050 319.050 ;
        RECT 286.950 310.950 289.050 313.050 ;
        RECT 289.950 310.950 292.050 313.050 ;
        RECT 293.250 311.250 294.750 312.150 ;
        RECT 295.950 310.950 298.050 313.050 ;
        RECT 298.950 310.950 301.050 313.050 ;
        RECT 302.250 311.250 303.750 312.150 ;
        RECT 304.950 310.950 307.050 313.050 ;
        RECT 308.400 310.050 309.450 316.950 ;
        RECT 311.400 312.450 312.450 343.950 ;
        RECT 314.400 333.600 315.600 350.400 ;
        RECT 317.400 334.050 318.450 377.400 ;
        RECT 322.950 361.950 325.050 364.050 ;
        RECT 319.950 341.250 322.050 342.150 ;
        RECT 319.950 337.950 322.050 340.050 ;
        RECT 313.950 331.500 316.050 333.600 ;
        RECT 316.950 331.950 319.050 334.050 ;
        RECT 320.400 313.050 321.450 337.950 ;
        RECT 323.400 322.050 324.450 361.950 ;
        RECT 325.950 341.250 328.050 342.150 ;
        RECT 325.950 337.950 328.050 340.050 ;
        RECT 326.400 330.450 327.450 337.950 ;
        RECT 329.400 334.050 330.450 379.950 ;
        RECT 334.950 351.300 337.050 353.400 ;
        RECT 337.950 352.950 340.050 355.050 ;
        RECT 335.250 347.700 336.450 351.300 ;
        RECT 334.950 345.600 337.050 347.700 ;
        RECT 331.950 340.950 334.050 343.050 ;
        RECT 328.950 331.950 331.050 334.050 ;
        RECT 326.400 329.400 330.450 330.450 ;
        RECT 325.950 325.950 328.050 328.050 ;
        RECT 322.950 319.950 325.050 322.050 ;
        RECT 326.400 313.050 327.450 325.950 ;
        RECT 311.400 311.400 315.450 312.450 ;
        RECT 314.400 310.050 315.450 311.400 ;
        RECT 316.950 310.950 319.050 313.050 ;
        RECT 319.950 310.950 322.050 313.050 ;
        RECT 323.250 311.250 324.750 312.150 ;
        RECT 325.950 310.950 328.050 313.050 ;
        RECT 317.400 310.050 318.450 310.950 ;
        RECT 286.950 309.450 289.050 310.050 ;
        RECT 284.400 308.400 289.050 309.450 ;
        RECT 290.250 308.850 291.750 309.750 ;
        RECT 284.400 304.050 285.450 308.400 ;
        RECT 286.950 307.950 289.050 308.400 ;
        RECT 292.950 307.950 295.050 310.050 ;
        RECT 296.250 308.850 298.050 309.750 ;
        RECT 298.950 308.850 300.750 309.750 ;
        RECT 301.950 307.950 304.050 310.050 ;
        RECT 305.250 308.850 306.750 309.750 ;
        RECT 307.950 309.450 310.050 310.050 ;
        RECT 307.950 308.400 312.450 309.450 ;
        RECT 307.950 307.950 310.050 308.400 ;
        RECT 286.950 305.850 289.050 306.750 ;
        RECT 289.950 304.950 292.050 307.050 ;
        RECT 283.950 301.950 286.050 304.050 ;
        RECT 280.950 298.950 283.050 301.050 ;
        RECT 284.400 297.450 285.450 301.950 ;
        RECT 281.400 296.400 285.450 297.450 ;
        RECT 256.950 283.950 259.050 286.050 ;
        RECT 262.950 283.950 265.050 286.050 ;
        RECT 263.400 274.050 264.450 283.950 ;
        RECT 268.950 275.250 271.050 276.150 ;
        RECT 281.400 274.050 282.450 296.400 ;
        RECT 286.950 295.950 289.050 298.050 ;
        RECT 250.950 271.950 253.050 274.050 ;
        RECT 262.950 271.950 265.050 274.050 ;
        RECT 266.250 272.250 267.750 273.150 ;
        RECT 268.950 271.950 271.050 274.050 ;
        RECT 280.950 273.450 283.050 274.050 ;
        RECT 272.250 272.250 274.050 273.150 ;
        RECT 278.400 272.400 283.050 273.450 ;
        RECT 247.950 259.950 250.050 262.050 ;
        RECT 251.400 244.050 252.450 271.950 ;
        RECT 253.950 269.250 255.750 270.150 ;
        RECT 262.950 269.850 264.750 270.750 ;
        RECT 265.950 268.950 268.050 271.050 ;
        RECT 271.950 268.950 274.050 271.050 ;
        RECT 274.950 269.250 277.050 270.150 ;
        RECT 253.950 265.950 256.050 268.050 ;
        RECT 257.250 266.850 259.050 267.750 ;
        RECT 259.950 265.950 262.050 268.050 ;
        RECT 254.400 256.050 255.450 265.950 ;
        RECT 253.950 253.950 256.050 256.050 ;
        RECT 250.950 241.950 253.050 244.050 ;
        RECT 247.950 237.450 250.050 238.050 ;
        RECT 245.400 236.400 250.050 237.450 ;
        RECT 217.950 233.850 219.750 234.750 ;
        RECT 220.950 232.950 223.050 235.050 ;
        RECT 224.250 233.850 225.750 234.750 ;
        RECT 226.950 232.950 229.050 235.050 ;
        RECT 220.950 230.850 223.050 231.750 ;
        RECT 214.950 223.950 217.050 226.050 ;
        RECT 217.950 223.950 220.050 226.050 ;
        RECT 211.950 220.950 214.050 223.050 ;
        RECT 205.950 202.950 208.050 205.050 ;
        RECT 208.950 202.950 211.050 205.050 ;
        RECT 205.950 200.250 208.050 201.150 ;
        RECT 193.950 197.250 196.050 198.150 ;
        RECT 196.950 197.250 198.750 198.150 ;
        RECT 199.950 196.950 202.050 199.050 ;
        RECT 203.250 197.250 204.750 198.150 ;
        RECT 205.950 196.950 208.050 199.050 ;
        RECT 193.950 193.950 196.050 196.050 ;
        RECT 196.950 193.950 199.050 196.050 ;
        RECT 200.250 194.850 201.750 195.750 ;
        RECT 202.950 193.950 205.050 196.050 ;
        RECT 194.400 172.050 195.450 193.950 ;
        RECT 197.400 193.050 198.450 193.950 ;
        RECT 196.950 190.950 199.050 193.050 ;
        RECT 199.950 187.950 202.050 190.050 ;
        RECT 193.950 169.950 196.050 172.050 ;
        RECT 193.950 166.950 196.050 169.050 ;
        RECT 193.950 164.850 196.050 165.750 ;
        RECT 196.950 164.250 199.050 165.150 ;
        RECT 193.950 151.950 196.050 154.050 ;
        RECT 181.950 130.950 184.050 133.050 ;
        RECT 187.950 131.250 190.050 132.150 ;
        RECT 190.950 130.950 193.050 133.050 ;
        RECT 182.400 130.050 183.450 130.950 ;
        RECT 181.950 127.950 184.050 130.050 ;
        RECT 185.250 128.250 186.750 129.150 ;
        RECT 187.950 127.950 190.050 130.050 ;
        RECT 191.250 128.250 193.050 129.150 ;
        RECT 188.400 127.050 189.450 127.950 ;
        RECT 194.400 127.050 195.450 151.950 ;
        RECT 196.950 136.950 199.050 139.050 ;
        RECT 197.400 127.050 198.450 136.950 ;
        RECT 200.400 130.050 201.450 187.950 ;
        RECT 203.400 181.050 204.450 193.950 ;
        RECT 206.400 190.050 207.450 196.950 ;
        RECT 205.950 187.950 208.050 190.050 ;
        RECT 209.400 186.450 210.450 202.950 ;
        RECT 218.400 202.050 219.450 223.950 ;
        RECT 223.950 220.950 226.050 223.050 ;
        RECT 220.950 205.950 223.050 208.050 ;
        RECT 214.950 200.250 217.050 201.150 ;
        RECT 217.950 199.950 220.050 202.050 ;
        RECT 221.400 199.050 222.450 205.950 ;
        RECT 224.400 205.050 225.450 220.950 ;
        RECT 233.400 220.050 234.450 235.950 ;
        RECT 232.950 217.950 235.050 220.050 ;
        RECT 226.950 214.950 229.050 217.050 ;
        RECT 223.950 202.950 226.050 205.050 ;
        RECT 227.400 202.050 228.450 214.950 ;
        RECT 226.950 199.950 229.050 202.050 ;
        RECT 230.250 200.250 231.750 201.150 ;
        RECT 214.950 196.950 217.050 199.050 ;
        RECT 218.250 197.250 219.750 198.150 ;
        RECT 220.950 196.950 223.050 199.050 ;
        RECT 224.250 197.250 226.050 198.150 ;
        RECT 226.950 197.850 228.750 198.750 ;
        RECT 229.950 196.950 232.050 199.050 ;
        RECT 233.250 197.850 235.050 198.750 ;
        RECT 217.950 193.950 220.050 196.050 ;
        RECT 221.250 194.850 222.750 195.750 ;
        RECT 223.950 193.950 226.050 196.050 ;
        RECT 224.400 193.050 225.450 193.950 ;
        RECT 223.950 190.950 226.050 193.050 ;
        RECT 230.400 190.050 231.450 196.950 ;
        RECT 229.950 187.950 232.050 190.050 ;
        RECT 232.950 187.950 235.050 190.050 ;
        RECT 206.400 185.400 210.450 186.450 ;
        RECT 202.950 178.950 205.050 181.050 ;
        RECT 202.950 169.950 205.050 172.050 ;
        RECT 203.400 169.050 204.450 169.950 ;
        RECT 206.400 169.050 207.450 185.400 ;
        RECT 208.950 181.950 211.050 184.050 ;
        RECT 202.950 166.950 205.050 169.050 ;
        RECT 205.950 166.950 208.050 169.050 ;
        RECT 209.400 166.050 210.450 181.950 ;
        RECT 226.950 172.950 229.050 175.050 ;
        RECT 214.950 166.950 217.050 169.050 ;
        RECT 220.950 166.950 223.050 169.050 ;
        RECT 224.250 167.250 226.050 168.150 ;
        RECT 202.950 164.850 205.050 165.750 ;
        RECT 205.950 164.250 207.750 165.150 ;
        RECT 208.950 163.950 211.050 166.050 ;
        RECT 212.250 164.250 214.050 165.150 ;
        RECT 202.950 160.950 205.050 163.050 ;
        RECT 205.950 160.950 208.050 163.050 ;
        RECT 209.250 161.850 210.750 162.750 ;
        RECT 203.400 139.050 204.450 160.950 ;
        RECT 202.950 136.950 205.050 139.050 ;
        RECT 206.400 133.050 207.450 160.950 ;
        RECT 215.400 148.050 216.450 166.950 ;
        RECT 220.950 164.850 222.750 165.750 ;
        RECT 227.400 162.450 228.450 172.950 ;
        RECT 233.400 169.050 234.450 187.950 ;
        RECT 236.400 187.050 237.450 235.950 ;
        RECT 239.400 226.050 240.450 235.950 ;
        RECT 245.400 235.050 246.450 236.400 ;
        RECT 247.950 235.950 250.050 236.400 ;
        RECT 250.950 235.950 253.050 238.050 ;
        RECT 253.950 235.950 256.050 238.050 ;
        RECT 257.250 236.250 259.050 237.150 ;
        RECT 251.400 235.050 252.450 235.950 ;
        RECT 244.950 232.950 247.050 235.050 ;
        RECT 247.950 233.850 249.750 234.750 ;
        RECT 250.950 232.950 253.050 235.050 ;
        RECT 254.250 233.850 255.750 234.750 ;
        RECT 256.950 234.450 259.050 235.050 ;
        RECT 260.400 234.450 261.450 265.950 ;
        RECT 266.400 265.050 267.450 268.950 ;
        RECT 272.400 268.050 273.450 268.950 ;
        RECT 278.400 268.050 279.450 272.400 ;
        RECT 280.950 271.950 283.050 272.400 ;
        RECT 280.950 269.850 283.050 270.750 ;
        RECT 283.950 269.250 286.050 270.150 ;
        RECT 271.950 265.950 274.050 268.050 ;
        RECT 274.950 265.950 277.050 268.050 ;
        RECT 277.950 265.950 280.050 268.050 ;
        RECT 283.950 267.450 286.050 268.050 ;
        RECT 287.400 267.450 288.450 295.950 ;
        RECT 290.400 274.050 291.450 304.950 ;
        RECT 298.950 301.950 301.050 304.050 ;
        RECT 295.950 278.400 298.050 280.500 ;
        RECT 289.950 271.950 292.050 274.050 ;
        RECT 283.950 266.400 288.450 267.450 ;
        RECT 283.950 265.950 286.050 266.400 ;
        RECT 275.400 265.050 276.450 265.950 ;
        RECT 265.950 262.950 268.050 265.050 ;
        RECT 274.950 262.950 277.050 265.050 ;
        RECT 266.400 261.450 267.450 262.950 ;
        RECT 266.400 260.400 270.450 261.450 ;
        RECT 269.400 241.050 270.450 260.400 ;
        RECT 274.950 256.950 277.050 259.050 ;
        RECT 275.400 244.050 276.450 256.950 ;
        RECT 277.950 247.950 280.050 250.050 ;
        RECT 274.950 241.950 277.050 244.050 ;
        RECT 262.950 238.950 265.050 241.050 ;
        RECT 266.250 239.250 267.750 240.150 ;
        RECT 268.950 238.950 271.050 241.050 ;
        RECT 274.950 238.950 277.050 241.050 ;
        RECT 262.950 236.850 264.750 237.750 ;
        RECT 265.950 235.950 268.050 238.050 ;
        RECT 269.250 236.850 270.750 237.750 ;
        RECT 271.950 237.450 274.050 238.050 ;
        RECT 275.400 237.450 276.450 238.950 ;
        RECT 271.950 236.400 276.450 237.450 ;
        RECT 271.950 235.950 274.050 236.400 ;
        RECT 256.950 233.400 261.450 234.450 ;
        RECT 256.950 232.950 259.050 233.400 ;
        RECT 262.950 232.950 265.050 235.050 ;
        RECT 250.950 230.850 253.050 231.750 ;
        RECT 241.950 226.950 244.050 229.050 ;
        RECT 238.950 223.950 241.050 226.050 ;
        RECT 242.400 199.050 243.450 226.950 ;
        RECT 253.950 220.950 256.050 223.050 ;
        RECT 250.950 202.950 253.050 205.050 ;
        RECT 247.950 200.250 250.050 201.150 ;
        RECT 238.950 197.250 240.750 198.150 ;
        RECT 241.950 196.950 244.050 199.050 ;
        RECT 245.250 197.250 246.750 198.150 ;
        RECT 247.950 196.950 250.050 199.050 ;
        RECT 238.950 193.950 241.050 196.050 ;
        RECT 242.250 194.850 243.750 195.750 ;
        RECT 244.950 193.950 247.050 196.050 ;
        RECT 235.950 184.950 238.050 187.050 ;
        RECT 235.950 175.950 238.050 178.050 ;
        RECT 236.400 172.050 237.450 175.950 ;
        RECT 235.950 169.950 238.050 172.050 ;
        RECT 232.950 166.950 235.050 169.050 ;
        RECT 229.950 164.250 231.750 165.150 ;
        RECT 232.950 163.950 235.050 166.050 ;
        RECT 236.250 164.250 238.050 165.150 ;
        RECT 229.950 162.450 232.050 163.050 ;
        RECT 227.400 161.400 232.050 162.450 ;
        RECT 233.250 161.850 234.750 162.750 ;
        RECT 229.950 160.950 232.050 161.400 ;
        RECT 235.950 160.950 238.050 163.050 ;
        RECT 230.400 151.050 231.450 160.950 ;
        RECT 236.400 157.050 237.450 160.950 ;
        RECT 235.950 154.950 238.050 157.050 ;
        RECT 229.950 148.950 232.050 151.050 ;
        RECT 214.950 145.950 217.050 148.050 ;
        RECT 229.950 139.950 232.050 142.050 ;
        RECT 214.950 136.950 217.050 139.050 ;
        RECT 205.950 130.950 208.050 133.050 ;
        RECT 199.950 127.950 202.050 130.050 ;
        RECT 205.950 127.950 208.050 130.050 ;
        RECT 211.950 128.250 214.050 129.150 ;
        RECT 206.400 127.050 207.450 127.950 ;
        RECT 170.250 125.250 171.750 126.150 ;
        RECT 172.950 125.400 177.450 126.450 ;
        RECT 172.950 124.950 175.050 125.400 ;
        RECT 178.950 124.950 181.050 127.050 ;
        RECT 181.950 125.850 183.750 126.750 ;
        RECT 184.950 124.950 187.050 127.050 ;
        RECT 187.950 124.950 190.050 127.050 ;
        RECT 190.950 124.950 193.050 127.050 ;
        RECT 193.950 124.950 196.050 127.050 ;
        RECT 196.950 124.950 199.050 127.050 ;
        RECT 202.950 125.250 204.750 126.150 ;
        RECT 205.950 124.950 208.050 127.050 ;
        RECT 209.250 125.250 210.750 126.150 ;
        RECT 211.950 124.950 214.050 127.050 ;
        RECT 155.400 115.050 156.450 124.950 ;
        RECT 154.950 112.950 157.050 115.050 ;
        RECT 148.950 106.950 151.050 109.050 ;
        RECT 133.950 103.950 136.050 106.050 ;
        RECT 142.950 103.950 145.050 106.050 ;
        RECT 130.950 97.950 133.050 100.050 ;
        RECT 131.400 97.050 132.450 97.950 ;
        RECT 112.950 96.450 115.050 97.050 ;
        RECT 112.950 95.400 117.450 96.450 ;
        RECT 112.950 94.950 115.050 95.400 ;
        RECT 112.950 92.850 115.050 93.750 ;
        RECT 116.400 91.050 117.450 95.400 ;
        RECT 121.950 94.950 124.050 97.050 ;
        RECT 127.950 94.950 130.050 97.050 ;
        RECT 130.950 94.950 133.050 97.050 ;
        RECT 134.400 94.050 135.450 103.950 ;
        RECT 136.950 100.950 139.050 103.050 ;
        RECT 137.400 97.050 138.450 100.950 ;
        RECT 143.400 97.050 144.450 103.950 ;
        RECT 151.950 100.950 154.050 103.050 ;
        RECT 148.950 97.950 151.050 100.050 ;
        RECT 136.950 94.950 139.050 97.050 ;
        RECT 140.250 95.250 141.750 96.150 ;
        RECT 142.950 94.950 145.050 97.050 ;
        RECT 118.950 92.850 121.050 93.750 ;
        RECT 121.950 92.850 124.050 93.750 ;
        RECT 127.950 92.250 130.050 93.150 ;
        RECT 130.950 92.850 133.050 93.750 ;
        RECT 133.950 91.950 136.050 94.050 ;
        RECT 136.950 92.850 138.750 93.750 ;
        RECT 139.950 91.950 142.050 94.050 ;
        RECT 143.250 92.850 144.750 93.750 ;
        RECT 145.950 91.950 148.050 94.050 ;
        RECT 115.950 88.950 118.050 91.050 ;
        RECT 127.950 88.950 130.050 91.050 ;
        RECT 130.950 88.950 133.050 91.050 ;
        RECT 115.950 79.950 118.050 82.050 ;
        RECT 116.400 55.050 117.450 79.950 ;
        RECT 128.400 61.050 129.450 88.950 ;
        RECT 131.400 70.050 132.450 88.950 ;
        RECT 134.400 88.050 135.450 91.950 ;
        RECT 145.950 89.850 148.050 90.750 ;
        RECT 133.950 85.950 136.050 88.050 ;
        RECT 130.950 67.950 133.050 70.050 ;
        RECT 131.400 66.450 132.450 67.950 ;
        RECT 131.400 65.400 135.450 66.450 ;
        RECT 130.950 61.950 133.050 64.050 ;
        RECT 127.950 58.950 130.050 61.050 ;
        RECT 131.400 58.050 132.450 61.950 ;
        RECT 134.400 58.050 135.450 65.400 ;
        RECT 149.400 64.050 150.450 97.950 ;
        RECT 152.400 97.050 153.450 100.950 ;
        RECT 158.400 100.050 159.450 124.950 ;
        RECT 161.400 118.050 162.450 124.950 ;
        RECT 163.950 121.950 166.050 124.050 ;
        RECT 167.250 122.850 168.750 123.750 ;
        RECT 169.950 121.950 172.050 124.050 ;
        RECT 164.400 121.050 165.450 121.950 ;
        RECT 163.950 118.950 166.050 121.050 ;
        RECT 160.950 115.950 163.050 118.050 ;
        RECT 154.950 97.950 157.050 100.050 ;
        RECT 157.950 97.950 160.050 100.050 ;
        RECT 151.950 94.950 154.050 97.050 ;
        RECT 155.400 94.050 156.450 97.950 ;
        RECT 164.400 97.050 165.450 118.950 ;
        RECT 170.400 115.050 171.450 121.950 ;
        RECT 169.950 112.950 172.050 115.050 ;
        RECT 185.400 112.050 186.450 124.950 ;
        RECT 191.400 115.050 192.450 124.950 ;
        RECT 193.950 122.250 196.050 123.150 ;
        RECT 196.950 122.850 199.050 123.750 ;
        RECT 202.950 121.950 205.050 124.050 ;
        RECT 206.250 122.850 207.750 123.750 ;
        RECT 208.950 121.950 211.050 124.050 ;
        RECT 203.400 121.050 204.450 121.950 ;
        RECT 193.950 118.950 196.050 121.050 ;
        RECT 202.950 118.950 205.050 121.050 ;
        RECT 194.400 118.050 195.450 118.950 ;
        RECT 193.950 115.950 196.050 118.050 ;
        RECT 209.400 115.050 210.450 121.950 ;
        RECT 190.950 112.950 193.050 115.050 ;
        RECT 208.950 112.950 211.050 115.050 ;
        RECT 211.950 112.950 214.050 115.050 ;
        RECT 184.950 109.950 187.050 112.050 ;
        RECT 184.950 106.950 187.050 109.050 ;
        RECT 178.950 103.950 181.050 106.050 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 157.950 94.950 160.050 97.050 ;
        RECT 161.250 95.250 162.750 96.150 ;
        RECT 163.950 94.950 166.050 97.050 ;
        RECT 167.400 94.050 168.450 100.950 ;
        RECT 179.400 100.050 180.450 103.950 ;
        RECT 178.950 97.950 181.050 100.050 ;
        RECT 185.400 97.050 186.450 106.950 ;
        RECT 196.950 103.950 199.050 106.050 ;
        RECT 199.950 103.950 202.050 106.050 ;
        RECT 197.400 100.050 198.450 103.950 ;
        RECT 196.950 97.950 199.050 100.050 ;
        RECT 200.400 97.050 201.450 103.950 ;
        RECT 212.400 97.050 213.450 112.950 ;
        RECT 215.400 112.050 216.450 136.950 ;
        RECT 230.400 132.450 231.450 139.950 ;
        RECT 239.400 133.050 240.450 193.950 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 242.400 172.050 243.450 178.950 ;
        RECT 245.400 178.050 246.450 193.950 ;
        RECT 248.400 193.050 249.450 196.950 ;
        RECT 247.950 190.950 250.050 193.050 ;
        RECT 244.950 175.950 247.050 178.050 ;
        RECT 251.400 172.050 252.450 202.950 ;
        RECT 254.400 202.050 255.450 220.950 ;
        RECT 263.400 202.050 264.450 232.950 ;
        RECT 266.400 232.050 267.450 235.950 ;
        RECT 268.950 232.950 271.050 235.050 ;
        RECT 271.950 233.850 274.050 234.750 ;
        RECT 265.950 229.950 268.050 232.050 ;
        RECT 269.400 223.050 270.450 232.950 ;
        RECT 278.400 232.050 279.450 247.950 ;
        RECT 290.400 244.050 291.450 271.950 ;
        RECT 296.400 261.600 297.600 278.400 ;
        RECT 295.950 259.500 298.050 261.600 ;
        RECT 292.950 244.950 295.050 247.050 ;
        RECT 293.400 244.050 294.450 244.950 ;
        RECT 286.950 241.950 289.050 244.050 ;
        RECT 289.950 241.950 292.050 244.050 ;
        RECT 292.950 241.950 295.050 244.050 ;
        RECT 280.950 238.950 283.050 241.050 ;
        RECT 284.250 239.250 286.050 240.150 ;
        RECT 286.950 239.850 289.050 240.750 ;
        RECT 289.950 239.250 292.050 240.150 ;
        RECT 292.950 239.850 295.050 240.750 ;
        RECT 295.950 239.250 298.050 240.150 ;
        RECT 280.950 236.850 282.750 237.750 ;
        RECT 283.950 235.950 286.050 238.050 ;
        RECT 286.950 235.950 289.050 238.050 ;
        RECT 289.950 235.950 292.050 238.050 ;
        RECT 292.950 235.950 295.050 238.050 ;
        RECT 295.950 235.950 298.050 238.050 ;
        RECT 284.400 235.050 285.450 235.950 ;
        RECT 283.950 232.950 286.050 235.050 ;
        RECT 277.950 229.950 280.050 232.050 ;
        RECT 268.950 220.950 271.050 223.050 ;
        RECT 287.400 205.050 288.450 235.950 ;
        RECT 290.400 208.050 291.450 235.950 ;
        RECT 289.950 205.950 292.050 208.050 ;
        RECT 283.950 203.250 286.050 204.150 ;
        RECT 286.950 202.950 289.050 205.050 ;
        RECT 253.950 199.950 256.050 202.050 ;
        RECT 257.250 200.250 258.750 201.150 ;
        RECT 262.950 199.950 265.050 202.050 ;
        RECT 280.950 200.250 282.750 201.150 ;
        RECT 283.950 199.950 286.050 202.050 ;
        RECT 287.250 200.250 288.750 201.150 ;
        RECT 289.950 199.950 292.050 202.050 ;
        RECT 253.950 197.850 255.750 198.750 ;
        RECT 256.950 196.950 259.050 199.050 ;
        RECT 260.250 197.850 262.050 198.750 ;
        RECT 265.950 196.950 268.050 199.050 ;
        RECT 271.950 196.950 274.050 199.050 ;
        RECT 275.250 197.250 277.050 198.150 ;
        RECT 280.950 196.950 283.050 199.050 ;
        RECT 253.950 193.950 256.050 196.050 ;
        RECT 254.400 190.050 255.450 193.950 ;
        RECT 257.400 193.050 258.450 196.950 ;
        RECT 281.400 196.050 282.450 196.950 ;
        RECT 265.950 194.850 268.050 195.750 ;
        RECT 268.950 194.250 271.050 195.150 ;
        RECT 271.950 194.850 273.750 195.750 ;
        RECT 274.950 193.950 277.050 196.050 ;
        RECT 280.950 193.950 283.050 196.050 ;
        RECT 256.950 190.950 259.050 193.050 ;
        RECT 268.950 190.950 271.050 193.050 ;
        RECT 253.950 187.950 256.050 190.050 ;
        RECT 265.950 178.950 268.050 181.050 ;
        RECT 253.950 172.950 256.050 175.050 ;
        RECT 254.400 172.050 255.450 172.950 ;
        RECT 241.950 169.950 244.050 172.050 ;
        RECT 244.950 169.950 247.050 172.050 ;
        RECT 250.950 169.950 253.050 172.050 ;
        RECT 253.950 169.950 256.050 172.050 ;
        RECT 245.400 166.050 246.450 169.950 ;
        RECT 250.950 166.950 253.050 169.050 ;
        RECT 251.400 166.050 252.450 166.950 ;
        RECT 241.950 164.250 243.750 165.150 ;
        RECT 244.950 163.950 247.050 166.050 ;
        RECT 248.250 164.250 250.050 165.150 ;
        RECT 250.950 163.950 253.050 166.050 ;
        RECT 254.400 163.050 255.450 169.950 ;
        RECT 262.950 166.950 265.050 169.050 ;
        RECT 256.950 163.950 259.050 166.050 ;
        RECT 260.250 164.250 262.050 165.150 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 245.250 161.850 246.750 162.750 ;
        RECT 247.950 160.950 250.050 163.050 ;
        RECT 250.950 161.850 252.750 162.750 ;
        RECT 253.950 160.950 256.050 163.050 ;
        RECT 257.250 161.850 258.750 162.750 ;
        RECT 259.950 160.950 262.050 163.050 ;
        RECT 242.400 160.050 243.450 160.950 ;
        RECT 241.950 157.950 244.050 160.050 ;
        RECT 241.950 154.950 244.050 157.050 ;
        RECT 242.400 142.050 243.450 154.950 ;
        RECT 248.400 151.050 249.450 160.950 ;
        RECT 253.950 158.850 256.050 159.750 ;
        RECT 263.400 157.050 264.450 166.950 ;
        RECT 262.950 154.950 265.050 157.050 ;
        RECT 247.950 148.950 250.050 151.050 ;
        RECT 266.400 142.050 267.450 178.950 ;
        RECT 269.400 172.050 270.450 190.950 ;
        RECT 275.400 190.050 276.450 193.950 ;
        RECT 274.950 187.950 277.050 190.050 ;
        RECT 268.950 169.950 271.050 172.050 ;
        RECT 277.950 169.950 280.050 172.050 ;
        RECT 278.400 166.050 279.450 169.950 ;
        RECT 281.400 169.050 282.450 193.950 ;
        RECT 284.400 193.050 285.450 199.950 ;
        RECT 286.950 196.950 289.050 199.050 ;
        RECT 290.250 197.850 292.050 198.750 ;
        RECT 283.950 190.950 286.050 193.050 ;
        RECT 280.950 166.950 283.050 169.050 ;
        RECT 287.400 168.450 288.450 196.950 ;
        RECT 289.950 193.950 292.050 196.050 ;
        RECT 290.400 190.050 291.450 193.950 ;
        RECT 293.400 190.050 294.450 235.950 ;
        RECT 296.400 235.050 297.450 235.950 ;
        RECT 299.400 235.050 300.450 301.950 ;
        RECT 302.400 301.050 303.450 307.950 ;
        RECT 307.950 305.850 310.050 306.750 ;
        RECT 301.950 298.950 304.050 301.050 ;
        RECT 311.400 292.050 312.450 308.400 ;
        RECT 313.950 307.950 316.050 310.050 ;
        RECT 316.950 307.950 319.050 310.050 ;
        RECT 320.250 308.850 321.750 309.750 ;
        RECT 322.950 307.950 325.050 310.050 ;
        RECT 326.250 308.850 328.050 309.750 ;
        RECT 329.400 309.450 330.450 329.400 ;
        RECT 332.400 319.050 333.450 340.950 ;
        RECT 335.250 333.600 336.450 345.600 ;
        RECT 338.400 343.050 339.450 352.950 ;
        RECT 340.950 346.950 343.050 349.050 ;
        RECT 337.950 340.950 340.050 343.050 ;
        RECT 337.950 337.950 340.050 340.050 ;
        RECT 341.400 337.050 342.450 346.950 ;
        RECT 344.400 340.050 345.450 394.950 ;
        RECT 349.950 385.950 352.050 388.050 ;
        RECT 346.950 383.250 349.050 384.150 ;
        RECT 349.950 383.850 352.050 384.750 ;
        RECT 346.950 379.950 349.050 382.050 ;
        RECT 349.950 376.950 352.050 379.050 ;
        RECT 350.400 343.050 351.450 376.950 ;
        RECT 353.400 346.050 354.450 415.950 ;
        RECT 362.400 415.050 363.450 446.400 ;
        RECT 365.400 418.050 366.450 455.400 ;
        RECT 370.950 455.250 373.050 456.150 ;
        RECT 367.950 451.950 370.050 454.050 ;
        RECT 370.950 451.950 373.050 454.050 ;
        RECT 368.400 448.050 369.450 451.950 ;
        RECT 367.950 445.950 370.050 448.050 ;
        RECT 371.400 421.050 372.450 451.950 ;
        RECT 374.400 424.050 375.450 535.950 ;
        RECT 380.400 532.050 381.450 553.950 ;
        RECT 383.250 549.600 384.450 561.600 ;
        RECT 392.400 556.050 393.450 595.950 ;
        RECT 401.400 595.050 402.450 634.950 ;
        RECT 406.950 629.250 409.050 630.150 ;
        RECT 412.950 629.250 415.050 630.150 ;
        RECT 406.950 625.950 409.050 628.050 ;
        RECT 412.950 625.950 415.050 628.050 ;
        RECT 407.400 613.050 408.450 625.950 ;
        RECT 413.400 619.050 414.450 625.950 ;
        RECT 419.400 621.600 420.600 638.400 ;
        RECT 418.950 619.500 421.050 621.600 ;
        RECT 412.950 616.950 415.050 619.050 ;
        RECT 422.400 613.050 423.450 671.400 ;
        RECT 424.950 670.950 427.050 671.400 ;
        RECT 424.950 668.850 427.050 669.750 ;
        RECT 434.250 665.400 435.450 677.400 ;
        RECT 451.950 676.950 454.050 679.050 ;
        RECT 457.950 676.950 460.050 679.050 ;
        RECT 463.950 676.950 466.050 679.050 ;
        RECT 469.950 678.450 472.050 679.050 ;
        RECT 469.950 677.400 474.450 678.450 ;
        RECT 469.950 676.950 472.050 677.400 ;
        RECT 436.950 674.250 439.050 675.150 ;
        RECT 439.950 673.950 442.050 676.050 ;
        RECT 448.950 673.950 451.050 676.050 ;
        RECT 436.950 672.450 439.050 673.050 ;
        RECT 440.400 672.450 441.450 673.950 ;
        RECT 436.950 671.400 441.450 672.450 ;
        RECT 436.950 670.950 439.050 671.400 ;
        RECT 445.950 671.250 448.050 672.150 ;
        RECT 448.950 671.850 451.050 672.750 ;
        RECT 445.950 667.950 448.050 670.050 ;
        RECT 433.950 663.300 436.050 665.400 ;
        RECT 452.400 664.050 453.450 676.950 ;
        RECT 458.400 673.050 459.450 676.950 ;
        RECT 464.400 673.050 465.450 676.950 ;
        RECT 473.400 676.050 474.450 677.400 ;
        RECT 475.950 676.950 478.050 679.050 ;
        RECT 484.950 676.950 487.050 679.050 ;
        RECT 476.400 676.050 477.450 676.950 ;
        RECT 466.950 673.950 469.050 676.050 ;
        RECT 469.950 673.950 472.050 676.050 ;
        RECT 472.950 673.950 475.050 676.050 ;
        RECT 475.950 673.950 478.050 676.050 ;
        RECT 457.950 670.950 460.050 673.050 ;
        RECT 461.250 671.250 462.750 672.150 ;
        RECT 463.950 670.950 466.050 673.050 ;
        RECT 467.400 670.050 468.450 673.950 ;
        RECT 470.400 673.050 471.450 673.950 ;
        RECT 476.400 673.050 477.450 673.950 ;
        RECT 485.400 673.050 486.450 676.950 ;
        RECT 500.400 676.050 501.450 679.950 ;
        RECT 499.950 673.950 502.050 676.050 ;
        RECT 511.950 673.950 514.050 676.050 ;
        RECT 469.950 670.950 472.050 673.050 ;
        RECT 473.250 671.850 474.750 672.750 ;
        RECT 475.950 670.950 478.050 673.050 ;
        RECT 484.950 670.950 487.050 673.050 ;
        RECT 488.250 671.250 489.750 672.150 ;
        RECT 490.950 670.950 493.050 673.050 ;
        RECT 496.950 672.450 499.050 673.050 ;
        RECT 494.400 671.400 499.050 672.450 ;
        RECT 500.250 671.850 501.750 672.750 ;
        RECT 494.400 670.050 495.450 671.400 ;
        RECT 496.950 670.950 499.050 671.400 ;
        RECT 502.950 670.950 505.050 673.050 ;
        RECT 505.950 670.950 508.050 673.050 ;
        RECT 508.950 671.250 511.050 672.150 ;
        RECT 511.950 671.850 514.050 672.750 ;
        RECT 454.950 667.950 457.050 670.050 ;
        RECT 458.250 668.850 459.750 669.750 ;
        RECT 460.950 667.950 463.050 670.050 ;
        RECT 464.250 668.850 466.050 669.750 ;
        RECT 466.950 667.950 469.050 670.050 ;
        RECT 469.950 668.850 472.050 669.750 ;
        RECT 475.950 668.850 478.050 669.750 ;
        RECT 481.950 669.450 484.050 670.050 ;
        RECT 479.400 668.400 484.050 669.450 ;
        RECT 485.250 668.850 486.750 669.750 ;
        RECT 454.950 665.850 457.050 666.750 ;
        RECT 460.950 664.950 463.050 667.050 ;
        RECT 466.950 664.950 469.050 667.050 ;
        RECT 434.250 659.700 435.450 663.300 ;
        RECT 451.950 661.950 454.050 664.050 ;
        RECT 433.950 657.600 436.050 659.700 ;
        RECT 436.950 631.950 439.050 634.050 ;
        RECT 457.950 632.250 460.050 633.150 ;
        RECT 430.950 628.950 433.050 631.050 ;
        RECT 427.950 626.250 430.050 627.150 ;
        RECT 430.950 626.850 433.050 627.750 ;
        RECT 427.950 622.950 430.050 625.050 ;
        RECT 437.400 622.050 438.450 631.950 ;
        RECT 439.950 629.250 442.050 630.150 ;
        RECT 445.950 629.250 448.050 630.150 ;
        RECT 448.950 629.250 450.750 630.150 ;
        RECT 451.950 628.950 454.050 631.050 ;
        RECT 455.250 629.250 456.750 630.150 ;
        RECT 457.950 628.950 460.050 631.050 ;
        RECT 439.950 625.950 442.050 628.050 ;
        RECT 443.250 626.250 444.750 627.150 ;
        RECT 445.950 625.950 448.050 628.050 ;
        RECT 448.950 625.950 451.050 628.050 ;
        RECT 452.250 626.850 453.750 627.750 ;
        RECT 454.950 625.950 457.050 628.050 ;
        RECT 442.950 622.950 445.050 625.050 ;
        RECT 449.400 622.050 450.450 625.950 ;
        RECT 436.950 619.950 439.050 622.050 ;
        RECT 442.950 619.950 445.050 622.050 ;
        RECT 448.950 619.950 451.050 622.050 ;
        RECT 406.950 610.950 409.050 613.050 ;
        RECT 421.950 610.950 424.050 613.050 ;
        RECT 403.950 605.400 406.050 607.500 ;
        RECT 400.950 592.950 403.050 595.050 ;
        RECT 404.400 588.600 405.600 605.400 ;
        RECT 409.950 604.950 412.050 607.050 ;
        RECT 424.950 605.400 427.050 607.500 ;
        RECT 410.400 601.050 411.450 604.950 ;
        RECT 409.950 598.950 412.050 601.050 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 409.950 596.850 412.050 597.750 ;
        RECT 415.950 596.850 418.050 597.750 ;
        RECT 415.950 592.950 418.050 595.050 ;
        RECT 425.250 593.400 426.450 605.400 ;
        RECT 433.950 603.450 436.050 604.050 ;
        RECT 427.950 602.250 430.050 603.150 ;
        RECT 431.400 602.400 436.050 603.450 ;
        RECT 427.950 600.450 430.050 601.050 ;
        RECT 431.400 600.450 432.450 602.400 ;
        RECT 433.950 601.950 436.050 602.400 ;
        RECT 443.400 601.050 444.450 619.950 ;
        RECT 455.400 619.050 456.450 625.950 ;
        RECT 461.400 625.050 462.450 664.950 ;
        RECT 467.400 640.050 468.450 664.950 ;
        RECT 479.400 664.050 480.450 668.400 ;
        RECT 481.950 667.950 484.050 668.400 ;
        RECT 487.950 667.950 490.050 670.050 ;
        RECT 491.250 668.850 493.050 669.750 ;
        RECT 493.950 667.950 496.050 670.050 ;
        RECT 496.950 668.850 499.050 669.750 ;
        RECT 502.950 668.850 505.050 669.750 ;
        RECT 506.400 669.450 507.450 670.950 ;
        RECT 508.950 669.450 511.050 670.050 ;
        RECT 506.400 668.400 511.050 669.450 ;
        RECT 508.950 667.950 511.050 668.400 ;
        RECT 481.950 665.850 484.050 666.750 ;
        RECT 478.950 661.950 481.050 664.050 ;
        RECT 478.950 640.950 481.050 643.050 ;
        RECT 466.950 637.950 469.050 640.050 ;
        RECT 479.400 634.050 480.450 640.950 ;
        RECT 487.950 637.950 490.050 640.050 ;
        RECT 463.950 631.950 466.050 634.050 ;
        RECT 469.950 633.450 472.050 634.050 ;
        RECT 467.250 632.250 468.750 633.150 ;
        RECT 469.950 632.400 474.450 633.450 ;
        RECT 469.950 631.950 472.050 632.400 ;
        RECT 463.950 629.850 465.750 630.750 ;
        RECT 466.950 628.950 469.050 631.050 ;
        RECT 470.250 629.850 472.050 630.750 ;
        RECT 460.950 622.950 463.050 625.050 ;
        RECT 463.950 622.950 466.050 625.050 ;
        RECT 454.950 616.950 457.050 619.050 ;
        RECT 448.950 604.950 451.050 607.050 ;
        RECT 449.400 601.050 450.450 604.950 ;
        RECT 457.950 601.950 460.050 604.050 ;
        RECT 460.950 601.950 463.050 604.050 ;
        RECT 458.400 601.050 459.450 601.950 ;
        RECT 464.400 601.050 465.450 622.950 ;
        RECT 473.400 619.050 474.450 632.400 ;
        RECT 478.950 631.950 481.050 634.050 ;
        RECT 482.250 632.250 483.750 633.150 ;
        RECT 484.950 631.950 487.050 634.050 ;
        RECT 478.950 629.850 480.750 630.750 ;
        RECT 481.950 628.950 484.050 631.050 ;
        RECT 485.250 629.850 487.050 630.750 ;
        RECT 482.400 628.050 483.450 628.950 ;
        RECT 481.950 625.950 484.050 628.050 ;
        RECT 488.400 625.050 489.450 637.950 ;
        RECT 490.950 634.950 493.050 637.050 ;
        RECT 508.950 634.950 511.050 637.050 ;
        RECT 491.400 634.050 492.450 634.950 ;
        RECT 490.950 631.950 493.050 634.050 ;
        RECT 494.250 632.250 495.750 633.150 ;
        RECT 496.950 631.950 499.050 634.050 ;
        RECT 490.950 629.850 492.750 630.750 ;
        RECT 493.950 628.950 496.050 631.050 ;
        RECT 497.250 629.850 499.050 630.750 ;
        RECT 499.950 629.250 502.050 630.150 ;
        RECT 505.950 629.250 508.050 630.150 ;
        RECT 499.950 625.950 502.050 628.050 ;
        RECT 503.250 626.250 504.750 627.150 ;
        RECT 505.950 625.950 508.050 628.050 ;
        RECT 500.400 625.050 501.450 625.950 ;
        RECT 506.400 625.050 507.450 625.950 ;
        RECT 487.950 622.950 490.050 625.050 ;
        RECT 499.950 622.950 502.050 625.050 ;
        RECT 502.950 622.950 505.050 625.050 ;
        RECT 505.950 622.950 508.050 625.050 ;
        RECT 472.950 616.950 475.050 619.050 ;
        RECT 503.400 610.050 504.450 622.950 ;
        RECT 502.950 607.950 505.050 610.050 ;
        RECT 484.950 604.950 487.050 607.050 ;
        RECT 481.950 601.950 484.050 604.050 ;
        RECT 427.950 599.400 432.450 600.450 ;
        RECT 433.950 599.850 436.050 600.750 ;
        RECT 442.950 600.450 445.050 601.050 ;
        RECT 427.950 598.950 430.050 599.400 ;
        RECT 436.950 599.250 439.050 600.150 ;
        RECT 440.400 599.400 445.050 600.450 ;
        RECT 403.950 586.500 406.050 588.600 ;
        RECT 394.950 560.250 397.050 561.150 ;
        RECT 394.950 556.950 397.050 559.050 ;
        RECT 398.250 557.250 399.750 558.150 ;
        RECT 400.950 556.950 403.050 559.050 ;
        RECT 409.950 558.450 412.050 559.050 ;
        RECT 404.250 557.250 406.050 558.150 ;
        RECT 407.400 557.400 412.050 558.450 ;
        RECT 407.400 556.050 408.450 557.400 ;
        RECT 409.950 556.950 412.050 557.400 ;
        RECT 385.950 555.450 388.050 556.050 ;
        RECT 385.950 554.400 390.450 555.450 ;
        RECT 385.950 553.950 388.050 554.400 ;
        RECT 385.950 551.850 388.050 552.750 ;
        RECT 389.400 550.050 390.450 554.400 ;
        RECT 391.950 553.950 394.050 556.050 ;
        RECT 397.950 553.950 400.050 556.050 ;
        RECT 401.250 554.850 402.750 555.750 ;
        RECT 403.950 555.450 406.050 556.050 ;
        RECT 406.950 555.450 409.050 556.050 ;
        RECT 403.950 554.400 409.050 555.450 ;
        RECT 409.950 554.850 412.050 555.750 ;
        RECT 403.950 553.950 406.050 554.400 ;
        RECT 406.950 553.950 409.050 554.400 ;
        RECT 412.950 554.250 415.050 555.150 ;
        RECT 398.400 553.050 399.450 553.950 ;
        RECT 397.950 550.950 400.050 553.050 ;
        RECT 400.950 550.950 403.050 553.050 ;
        RECT 412.950 550.950 415.050 553.050 ;
        RECT 382.950 547.500 385.050 549.600 ;
        RECT 388.950 547.950 391.050 550.050 ;
        RECT 385.950 532.950 388.050 535.050 ;
        RECT 391.950 533.400 394.050 535.500 ;
        RECT 379.950 529.950 382.050 532.050 ;
        RECT 380.400 529.050 381.450 529.950 ;
        RECT 386.400 529.050 387.450 532.950 ;
        RECT 379.950 528.450 382.050 529.050 ;
        RECT 379.950 527.400 384.450 528.450 ;
        RECT 379.950 526.950 382.050 527.400 ;
        RECT 379.950 524.850 382.050 525.750 ;
        RECT 376.950 502.950 379.050 505.050 ;
        RECT 377.400 469.050 378.450 502.950 ;
        RECT 379.950 485.250 382.050 486.150 ;
        RECT 379.950 483.450 382.050 484.050 ;
        RECT 383.400 483.450 384.450 527.400 ;
        RECT 385.950 526.950 388.050 529.050 ;
        RECT 385.950 524.850 388.050 525.750 ;
        RECT 392.400 516.600 393.600 533.400 ;
        RECT 401.400 529.050 402.450 550.950 ;
        RECT 413.400 550.050 414.450 550.950 ;
        RECT 412.950 547.950 415.050 550.050 ;
        RECT 416.400 544.050 417.450 592.950 ;
        RECT 424.950 591.300 427.050 593.400 ;
        RECT 425.250 587.700 426.450 591.300 ;
        RECT 424.950 585.600 427.050 587.700 ;
        RECT 418.950 557.250 421.050 558.150 ;
        RECT 424.950 557.250 427.050 558.150 ;
        RECT 418.950 553.950 421.050 556.050 ;
        RECT 424.950 555.450 427.050 556.050 ;
        RECT 428.400 555.450 429.450 598.950 ;
        RECT 436.950 595.950 439.050 598.050 ;
        RECT 440.400 595.050 441.450 599.400 ;
        RECT 442.950 598.950 445.050 599.400 ;
        RECT 446.250 599.250 447.750 600.150 ;
        RECT 448.950 598.950 451.050 601.050 ;
        RECT 457.950 598.950 460.050 601.050 ;
        RECT 461.250 599.850 462.750 600.750 ;
        RECT 463.950 598.950 466.050 601.050 ;
        RECT 442.950 596.850 444.750 597.750 ;
        RECT 445.950 595.950 448.050 598.050 ;
        RECT 449.250 596.850 450.750 597.750 ;
        RECT 451.950 595.950 454.050 598.050 ;
        RECT 457.950 596.850 460.050 597.750 ;
        RECT 463.950 596.850 466.050 597.750 ;
        RECT 469.950 596.250 471.750 597.150 ;
        RECT 472.950 595.950 475.050 598.050 ;
        RECT 476.250 596.250 478.050 597.150 ;
        RECT 439.950 592.950 442.050 595.050 ;
        RECT 430.950 557.250 433.050 558.150 ;
        RECT 436.950 557.250 439.050 558.150 ;
        RECT 422.250 554.250 423.750 555.150 ;
        RECT 424.950 554.400 429.450 555.450 ;
        RECT 424.950 553.950 427.050 554.400 ;
        RECT 430.950 553.950 433.050 556.050 ;
        RECT 434.250 554.250 435.750 555.150 ;
        RECT 436.950 553.950 439.050 556.050 ;
        RECT 419.400 553.050 420.450 553.950 ;
        RECT 418.950 550.950 421.050 553.050 ;
        RECT 421.950 550.950 424.050 553.050 ;
        RECT 433.950 550.950 436.050 553.050 ;
        RECT 422.400 547.050 423.450 550.950 ;
        RECT 421.950 544.950 424.050 547.050 ;
        RECT 415.950 541.950 418.050 544.050 ;
        RECT 436.950 541.950 439.050 544.050 ;
        RECT 406.950 532.950 409.050 535.050 ;
        RECT 407.400 529.050 408.450 532.950 ;
        RECT 400.950 526.950 403.050 529.050 ;
        RECT 404.250 527.250 405.750 528.150 ;
        RECT 406.950 526.950 409.050 529.050 ;
        RECT 415.950 528.450 418.050 529.050 ;
        RECT 413.400 527.400 418.050 528.450 ;
        RECT 400.950 524.850 402.750 525.750 ;
        RECT 403.950 523.950 406.050 526.050 ;
        RECT 407.250 524.850 408.750 525.750 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 391.950 514.500 394.050 516.600 ;
        RECT 391.950 494.400 394.050 496.500 ;
        RECT 385.950 485.250 388.050 486.150 ;
        RECT 379.950 482.400 384.450 483.450 ;
        RECT 379.950 481.950 382.050 482.400 ;
        RECT 383.400 481.050 384.450 482.400 ;
        RECT 385.950 481.950 388.050 484.050 ;
        RECT 382.950 478.950 385.050 481.050 ;
        RECT 376.950 466.950 379.050 469.050 ;
        RECT 377.400 457.050 378.450 466.950 ;
        RECT 376.950 454.950 379.050 457.050 ;
        RECT 382.950 456.450 385.050 457.050 ;
        RECT 386.400 456.450 387.450 481.950 ;
        RECT 392.400 477.600 393.600 494.400 ;
        RECT 400.950 485.250 403.050 486.150 ;
        RECT 400.950 481.950 403.050 484.050 ;
        RECT 391.950 475.500 394.050 477.600 ;
        RECT 401.400 475.050 402.450 481.950 ;
        RECT 400.950 472.950 403.050 475.050 ;
        RECT 394.950 469.950 397.050 472.050 ;
        RECT 391.950 457.950 394.050 460.050 ;
        RECT 392.400 457.050 393.450 457.950 ;
        RECT 380.250 455.250 381.750 456.150 ;
        RECT 382.950 455.400 387.450 456.450 ;
        RECT 382.950 454.950 385.050 455.400 ;
        RECT 391.950 454.950 394.050 457.050 ;
        RECT 376.950 452.850 378.750 453.750 ;
        RECT 379.950 451.950 382.050 454.050 ;
        RECT 383.250 452.850 384.750 453.750 ;
        RECT 385.950 453.450 388.050 454.050 ;
        RECT 385.950 452.400 390.450 453.450 ;
        RECT 391.950 452.850 394.050 453.750 ;
        RECT 385.950 451.950 388.050 452.400 ;
        RECT 379.950 448.950 382.050 451.050 ;
        RECT 385.950 449.850 388.050 450.750 ;
        RECT 373.950 421.950 376.050 424.050 ;
        RECT 370.950 418.950 373.050 421.050 ;
        RECT 373.950 418.950 376.050 421.050 ;
        RECT 364.950 415.950 367.050 418.050 ;
        RECT 370.950 415.950 373.050 418.050 ;
        RECT 371.400 415.050 372.450 415.950 ;
        RECT 355.950 412.950 358.050 415.050 ;
        RECT 358.950 413.250 361.050 414.150 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 364.950 413.250 367.050 414.150 ;
        RECT 370.950 412.950 373.050 415.050 ;
        RECT 356.400 391.050 357.450 412.950 ;
        RECT 358.950 409.950 361.050 412.050 ;
        RECT 362.250 410.250 363.750 411.150 ;
        RECT 364.950 409.950 367.050 412.050 ;
        RECT 367.950 410.250 370.050 411.150 ;
        RECT 370.950 410.850 373.050 411.750 ;
        RECT 359.400 397.050 360.450 409.950 ;
        RECT 361.950 406.950 364.050 409.050 ;
        RECT 367.950 406.950 370.050 409.050 ;
        RECT 358.950 394.950 361.050 397.050 ;
        RECT 355.950 388.950 358.050 391.050 ;
        RECT 362.400 387.450 363.450 406.950 ;
        RECT 368.400 406.050 369.450 406.950 ;
        RECT 367.950 403.950 370.050 406.050 ;
        RECT 362.400 386.400 366.450 387.450 ;
        RECT 365.400 385.050 366.450 386.400 ;
        RECT 370.950 385.950 373.050 388.050 ;
        RECT 374.400 387.450 375.450 418.950 ;
        RECT 376.950 413.250 379.050 414.150 ;
        RECT 376.950 409.950 379.050 412.050 ;
        RECT 380.400 408.450 381.450 448.950 ;
        RECT 389.400 448.050 390.450 452.400 ;
        RECT 388.950 445.950 391.050 448.050 ;
        RECT 395.400 421.050 396.450 469.950 ;
        RECT 404.400 457.050 405.450 523.950 ;
        RECT 409.950 521.850 412.050 522.750 ;
        RECT 413.400 514.050 414.450 527.400 ;
        RECT 415.950 526.950 418.050 527.400 ;
        RECT 421.950 526.950 424.050 529.050 ;
        RECT 424.950 526.950 427.050 529.050 ;
        RECT 415.950 524.850 418.050 525.750 ;
        RECT 421.950 524.850 424.050 525.750 ;
        RECT 425.400 522.450 426.450 526.950 ;
        RECT 427.950 524.250 429.750 525.150 ;
        RECT 430.950 523.950 433.050 526.050 ;
        RECT 434.250 524.250 436.050 525.150 ;
        RECT 427.950 522.450 430.050 523.050 ;
        RECT 425.400 521.400 430.050 522.450 ;
        RECT 431.250 521.850 432.750 522.750 ;
        RECT 427.950 520.950 430.050 521.400 ;
        RECT 433.950 520.950 436.050 523.050 ;
        RECT 412.950 511.950 415.050 514.050 ;
        RECT 406.950 485.250 409.050 486.150 ;
        RECT 406.950 481.950 409.050 484.050 ;
        RECT 407.400 478.050 408.450 481.950 ;
        RECT 406.950 475.950 409.050 478.050 ;
        RECT 407.400 466.050 408.450 475.950 ;
        RECT 406.950 463.950 409.050 466.050 ;
        RECT 413.400 460.050 414.450 511.950 ;
        RECT 418.950 495.300 421.050 497.400 ;
        RECT 419.550 491.700 420.750 495.300 ;
        RECT 418.950 489.600 421.050 491.700 ;
        RECT 415.950 481.950 418.050 484.050 ;
        RECT 415.950 479.850 418.050 480.750 ;
        RECT 419.550 477.600 420.750 489.600 ;
        RECT 427.950 485.250 430.050 486.150 ;
        RECT 433.950 485.250 436.050 486.150 ;
        RECT 424.950 481.950 427.050 484.050 ;
        RECT 427.950 481.950 430.050 484.050 ;
        RECT 433.950 481.950 436.050 484.050 ;
        RECT 418.950 475.500 421.050 477.600 ;
        RECT 415.950 472.950 418.050 475.050 ;
        RECT 412.950 457.950 415.050 460.050 ;
        RECT 397.950 454.950 400.050 457.050 ;
        RECT 400.950 454.950 403.050 457.050 ;
        RECT 403.950 454.950 406.050 457.050 ;
        RECT 397.950 452.850 400.050 453.750 ;
        RECT 401.400 450.450 402.450 454.950 ;
        RECT 403.950 452.250 405.750 453.150 ;
        RECT 406.950 451.950 409.050 454.050 ;
        RECT 410.250 452.250 412.050 453.150 ;
        RECT 403.950 450.450 406.050 451.050 ;
        RECT 401.400 449.400 406.050 450.450 ;
        RECT 407.250 449.850 408.750 450.750 ;
        RECT 403.950 448.950 406.050 449.400 ;
        RECT 409.950 448.950 412.050 451.050 ;
        RECT 394.950 418.950 397.050 421.050 ;
        RECT 382.950 415.950 385.050 418.050 ;
        RECT 388.950 415.950 391.050 418.050 ;
        RECT 400.950 416.250 403.050 417.150 ;
        RECT 382.950 413.850 385.050 414.750 ;
        RECT 385.950 413.250 388.050 414.150 ;
        RECT 382.950 409.950 385.050 412.050 ;
        RECT 385.950 409.950 388.050 412.050 ;
        RECT 389.400 411.450 390.450 415.950 ;
        RECT 391.950 413.250 393.750 414.150 ;
        RECT 394.950 412.950 397.050 415.050 ;
        RECT 400.950 414.450 403.050 415.050 ;
        RECT 404.400 414.450 405.450 448.950 ;
        RECT 416.400 430.050 417.450 472.950 ;
        RECT 421.950 461.400 424.050 463.500 ;
        RECT 418.950 457.950 421.050 460.050 ;
        RECT 415.950 427.950 418.050 430.050 ;
        RECT 415.950 416.250 418.050 417.150 ;
        RECT 398.250 413.250 399.750 414.150 ;
        RECT 400.950 413.400 405.450 414.450 ;
        RECT 400.950 412.950 403.050 413.400 ;
        RECT 406.950 413.250 408.750 414.150 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 413.250 413.250 414.750 414.150 ;
        RECT 415.950 412.950 418.050 415.050 ;
        RECT 391.950 411.450 394.050 412.050 ;
        RECT 389.400 410.400 394.050 411.450 ;
        RECT 395.250 410.850 396.750 411.750 ;
        RECT 391.950 409.950 394.050 410.400 ;
        RECT 397.950 409.950 400.050 412.050 ;
        RECT 406.950 409.950 409.050 412.050 ;
        RECT 410.250 410.850 411.750 411.750 ;
        RECT 412.950 409.950 415.050 412.050 ;
        RECT 377.400 407.400 381.450 408.450 ;
        RECT 377.400 400.050 378.450 407.400 ;
        RECT 379.950 403.950 382.050 406.050 ;
        RECT 376.950 397.950 379.050 400.050 ;
        RECT 374.400 386.400 378.450 387.450 ;
        RECT 358.950 382.950 361.050 385.050 ;
        RECT 364.950 384.450 367.050 385.050 ;
        RECT 367.950 384.450 370.050 385.050 ;
        RECT 362.250 383.250 363.750 384.150 ;
        RECT 364.950 383.400 370.050 384.450 ;
        RECT 371.250 383.850 372.750 384.750 ;
        RECT 364.950 382.950 367.050 383.400 ;
        RECT 367.950 382.950 370.050 383.400 ;
        RECT 373.950 382.950 376.050 385.050 ;
        RECT 355.950 379.950 358.050 382.050 ;
        RECT 359.250 380.850 360.750 381.750 ;
        RECT 361.950 379.950 364.050 382.050 ;
        RECT 365.250 380.850 367.050 381.750 ;
        RECT 367.950 380.850 370.050 381.750 ;
        RECT 373.950 380.850 376.050 381.750 ;
        RECT 355.950 377.850 358.050 378.750 ;
        RECT 377.400 352.050 378.450 386.400 ;
        RECT 380.400 385.050 381.450 403.950 ;
        RECT 379.950 382.950 382.050 385.050 ;
        RECT 379.950 380.850 382.050 381.750 ;
        RECT 383.400 376.050 384.450 409.950 ;
        RECT 398.400 409.050 399.450 409.950 ;
        RECT 407.400 409.050 408.450 409.950 ;
        RECT 397.950 406.950 400.050 409.050 ;
        RECT 406.950 406.950 409.050 409.050 ;
        RECT 419.400 406.050 420.450 457.950 ;
        RECT 422.400 444.600 423.600 461.400 ;
        RECT 425.400 451.050 426.450 481.950 ;
        RECT 428.400 481.050 429.450 481.950 ;
        RECT 427.950 478.950 430.050 481.050 ;
        RECT 428.400 466.050 429.450 478.950 ;
        RECT 434.400 475.050 435.450 481.950 ;
        RECT 433.950 472.950 436.050 475.050 ;
        RECT 427.950 463.950 430.050 466.050 ;
        RECT 430.950 463.950 433.050 466.050 ;
        RECT 433.950 463.950 436.050 466.050 ;
        RECT 427.950 460.950 430.050 463.050 ;
        RECT 428.400 457.050 429.450 460.950 ;
        RECT 427.950 454.950 430.050 457.050 ;
        RECT 427.950 452.850 430.050 453.750 ;
        RECT 424.950 448.950 427.050 451.050 ;
        RECT 421.950 442.500 424.050 444.600 ;
        RECT 421.950 418.950 424.050 421.050 ;
        RECT 422.400 418.050 423.450 418.950 ;
        RECT 421.950 415.950 424.050 418.050 ;
        RECT 425.250 416.250 426.750 417.150 ;
        RECT 427.950 415.950 430.050 418.050 ;
        RECT 421.950 413.850 423.750 414.750 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 428.250 413.850 430.050 414.750 ;
        RECT 431.400 409.050 432.450 463.950 ;
        RECT 434.400 457.050 435.450 463.950 ;
        RECT 433.950 454.950 436.050 457.050 ;
        RECT 433.950 452.850 436.050 453.750 ;
        RECT 437.400 418.050 438.450 541.950 ;
        RECT 440.400 529.050 441.450 592.950 ;
        RECT 446.400 559.050 447.450 595.950 ;
        RECT 451.950 593.850 454.050 594.750 ;
        RECT 469.950 592.950 472.050 595.050 ;
        RECT 473.250 593.850 474.750 594.750 ;
        RECT 475.950 592.950 478.050 595.050 ;
        RECT 476.400 592.050 477.450 592.950 ;
        RECT 475.950 589.950 478.050 592.050 ;
        RECT 472.950 562.950 475.050 565.050 ;
        RECT 473.400 559.050 474.450 562.950 ;
        RECT 482.400 561.450 483.450 601.950 ;
        RECT 485.400 601.050 486.450 604.950 ;
        RECT 490.950 601.950 493.050 604.050 ;
        RECT 496.950 601.950 499.050 604.050 ;
        RECT 499.950 601.950 502.050 604.050 ;
        RECT 497.400 601.050 498.450 601.950 ;
        RECT 484.950 598.950 487.050 601.050 ;
        RECT 488.250 599.250 490.050 600.150 ;
        RECT 490.950 599.850 493.050 600.750 ;
        RECT 493.950 599.250 496.050 600.150 ;
        RECT 496.950 598.950 499.050 601.050 ;
        RECT 484.950 596.850 486.750 597.750 ;
        RECT 487.950 595.950 490.050 598.050 ;
        RECT 493.950 595.950 496.050 598.050 ;
        RECT 496.950 596.850 499.050 597.750 ;
        RECT 478.950 560.250 481.050 561.150 ;
        RECT 482.400 560.400 486.450 561.450 ;
        RECT 442.950 557.250 445.050 558.150 ;
        RECT 445.950 556.950 448.050 559.050 ;
        RECT 454.950 558.450 457.050 559.050 ;
        RECT 463.950 558.450 466.050 559.050 ;
        RECT 448.950 557.250 451.050 558.150 ;
        RECT 454.950 557.400 459.450 558.450 ;
        RECT 454.950 556.950 457.050 557.400 ;
        RECT 442.950 553.950 445.050 556.050 ;
        RECT 446.250 554.250 447.750 555.150 ;
        RECT 448.950 553.950 451.050 556.050 ;
        RECT 451.950 554.250 454.050 555.150 ;
        RECT 454.950 554.850 457.050 555.750 ;
        RECT 443.400 553.050 444.450 553.950 ;
        RECT 442.950 550.950 445.050 553.050 ;
        RECT 445.950 550.950 448.050 553.050 ;
        RECT 443.400 550.050 444.450 550.950 ;
        RECT 442.950 547.950 445.050 550.050 ;
        RECT 446.400 543.450 447.450 550.950 ;
        RECT 449.400 547.050 450.450 553.950 ;
        RECT 451.950 550.950 454.050 553.050 ;
        RECT 448.950 544.950 451.050 547.050 ;
        RECT 452.400 543.450 453.450 550.950 ;
        RECT 446.400 542.400 453.450 543.450 ;
        RECT 458.400 541.050 459.450 557.400 ;
        RECT 461.400 557.400 466.050 558.450 ;
        RECT 461.400 553.050 462.450 557.400 ;
        RECT 463.950 556.950 466.050 557.400 ;
        RECT 469.950 557.250 471.750 558.150 ;
        RECT 472.950 556.950 475.050 559.050 ;
        RECT 476.250 557.250 477.750 558.150 ;
        RECT 478.950 556.950 481.050 559.050 ;
        RECT 481.950 556.950 484.050 559.050 ;
        RECT 463.950 554.850 466.050 555.750 ;
        RECT 466.950 554.250 469.050 555.150 ;
        RECT 469.950 553.950 472.050 556.050 ;
        RECT 473.250 554.850 474.750 555.750 ;
        RECT 475.950 553.950 478.050 556.050 ;
        RECT 460.950 550.950 463.050 553.050 ;
        RECT 466.950 550.950 469.050 553.050 ;
        RECT 467.400 550.050 468.450 550.950 ;
        RECT 466.950 547.950 469.050 550.050 ;
        RECT 470.400 547.050 471.450 553.950 ;
        RECT 469.950 544.950 472.050 547.050 ;
        RECT 457.950 538.950 460.050 541.050 ;
        RECT 476.400 538.050 477.450 553.950 ;
        RECT 479.400 553.050 480.450 556.950 ;
        RECT 478.950 550.950 481.050 553.050 ;
        RECT 475.950 535.950 478.050 538.050 ;
        RECT 445.950 533.400 448.050 535.500 ;
        RECT 466.950 533.400 469.050 535.500 ;
        RECT 482.400 535.050 483.450 556.950 ;
        RECT 442.950 530.250 445.050 531.150 ;
        RECT 439.950 526.950 442.050 529.050 ;
        RECT 442.950 526.950 445.050 529.050 ;
        RECT 443.400 523.050 444.450 526.950 ;
        RECT 442.950 520.950 445.050 523.050 ;
        RECT 446.550 521.400 447.750 533.400 ;
        RECT 454.950 529.950 457.050 532.050 ;
        RECT 455.400 529.050 456.450 529.950 ;
        RECT 454.950 526.950 457.050 529.050 ;
        RECT 460.950 526.950 463.050 529.050 ;
        RECT 454.950 524.850 457.050 525.750 ;
        RECT 460.950 524.850 463.050 525.750 ;
        RECT 439.950 494.400 442.050 496.500 ;
        RECT 440.400 477.600 441.600 494.400 ;
        RECT 443.400 487.050 444.450 520.950 ;
        RECT 445.950 519.300 448.050 521.400 ;
        RECT 446.550 515.700 447.750 519.300 ;
        RECT 448.950 517.950 451.050 520.050 ;
        RECT 445.950 513.600 448.050 515.700 ;
        RECT 442.950 484.950 445.050 487.050 ;
        RECT 445.950 481.950 448.050 484.050 ;
        RECT 439.950 475.500 442.050 477.600 ;
        RECT 446.400 469.050 447.450 481.950 ;
        RECT 445.950 466.950 448.050 469.050 ;
        RECT 442.950 461.400 445.050 463.500 ;
        RECT 443.250 449.400 444.450 461.400 ;
        RECT 445.950 458.250 448.050 459.150 ;
        RECT 445.950 454.950 448.050 457.050 ;
        RECT 442.950 447.300 445.050 449.400 ;
        RECT 446.400 448.050 447.450 454.950 ;
        RECT 449.400 451.050 450.450 517.950 ;
        RECT 467.400 516.600 468.600 533.400 ;
        RECT 481.950 532.950 484.050 535.050 ;
        RECT 485.400 532.050 486.450 560.400 ;
        RECT 490.950 559.950 493.050 562.050 ;
        RECT 491.400 559.050 492.450 559.950 ;
        RECT 494.400 559.050 495.450 595.950 ;
        RECT 500.400 559.050 501.450 601.950 ;
        RECT 503.400 601.050 504.450 607.950 ;
        RECT 502.950 598.950 505.050 601.050 ;
        RECT 505.950 598.950 508.050 601.050 ;
        RECT 502.950 596.250 505.050 597.150 ;
        RECT 505.950 596.850 508.050 597.750 ;
        RECT 502.950 592.950 505.050 595.050 ;
        RECT 505.950 592.950 508.050 595.050 ;
        RECT 506.400 559.050 507.450 592.950 ;
        RECT 509.400 562.050 510.450 634.950 ;
        RECT 515.400 625.050 516.450 679.950 ;
        RECT 520.950 677.400 523.050 679.500 ;
        RECT 517.950 674.250 520.050 675.150 ;
        RECT 517.950 670.950 520.050 673.050 ;
        RECT 521.550 665.400 522.750 677.400 ;
        RECT 523.950 676.950 526.050 679.050 ;
        RECT 541.950 677.400 544.050 679.500 ;
        RECT 520.950 663.300 523.050 665.400 ;
        RECT 521.550 659.700 522.750 663.300 ;
        RECT 520.950 657.600 523.050 659.700 ;
        RECT 517.950 638.400 520.050 640.500 ;
        RECT 514.950 622.950 517.050 625.050 ;
        RECT 518.400 621.600 519.600 638.400 ;
        RECT 524.400 637.050 525.450 676.950 ;
        RECT 529.950 672.450 532.050 673.050 ;
        RECT 527.400 671.400 532.050 672.450 ;
        RECT 523.950 634.950 526.050 637.050 ;
        RECT 523.950 629.250 526.050 630.150 ;
        RECT 523.950 625.950 526.050 628.050 ;
        RECT 527.400 627.450 528.450 671.400 ;
        RECT 529.950 670.950 532.050 671.400 ;
        RECT 535.950 670.950 538.050 673.050 ;
        RECT 529.950 668.850 532.050 669.750 ;
        RECT 535.950 668.850 538.050 669.750 ;
        RECT 542.400 660.600 543.600 677.400 ;
        RECT 595.950 676.950 598.050 679.050 ;
        RECT 661.950 677.400 664.050 679.500 ;
        RECT 682.950 677.400 685.050 679.500 ;
        RECT 550.950 672.450 553.050 673.050 ;
        RECT 548.400 671.400 553.050 672.450 ;
        RECT 548.400 667.050 549.450 671.400 ;
        RECT 550.950 670.950 553.050 671.400 ;
        RECT 554.250 671.250 555.750 672.150 ;
        RECT 556.950 670.950 559.050 673.050 ;
        RECT 580.950 671.250 583.050 672.150 ;
        RECT 550.950 668.850 552.750 669.750 ;
        RECT 553.950 667.950 556.050 670.050 ;
        RECT 557.250 668.850 558.750 669.750 ;
        RECT 559.950 667.950 562.050 670.050 ;
        RECT 565.950 668.250 567.750 669.150 ;
        RECT 568.950 667.950 571.050 670.050 ;
        RECT 572.250 668.250 574.050 669.150 ;
        RECT 580.950 667.950 583.050 670.050 ;
        RECT 547.950 664.950 550.050 667.050 ;
        RECT 559.950 665.850 562.050 666.750 ;
        RECT 565.950 664.950 568.050 667.050 ;
        RECT 569.250 665.850 570.750 666.750 ;
        RECT 571.950 664.950 574.050 667.050 ;
        RECT 541.950 658.500 544.050 660.600 ;
        RECT 538.950 639.300 541.050 641.400 ;
        RECT 539.250 635.700 540.450 639.300 ;
        RECT 538.950 633.600 541.050 635.700 ;
        RECT 547.950 634.950 550.050 637.050 ;
        RECT 556.950 634.950 559.050 637.050 ;
        RECT 529.950 629.250 532.050 630.150 ;
        RECT 529.950 627.450 532.050 628.050 ;
        RECT 527.400 626.400 532.050 627.450 ;
        RECT 529.950 625.950 532.050 626.400 ;
        RECT 517.950 619.500 520.050 621.600 ;
        RECT 530.400 613.050 531.450 625.950 ;
        RECT 539.250 621.600 540.450 633.600 ;
        RECT 541.950 631.950 544.050 634.050 ;
        RECT 542.400 628.050 543.450 631.950 ;
        RECT 541.950 625.950 544.050 628.050 ;
        RECT 548.400 625.050 549.450 634.950 ;
        RECT 557.400 634.050 558.450 634.950 ;
        RECT 550.950 631.950 553.050 634.050 ;
        RECT 554.250 632.250 555.750 633.150 ;
        RECT 556.950 631.950 559.050 634.050 ;
        RECT 572.400 631.050 573.450 664.950 ;
        RECT 577.950 639.300 580.050 641.400 ;
        RECT 578.550 635.700 579.750 639.300 ;
        RECT 577.950 633.600 580.050 635.700 ;
        RECT 550.950 629.850 552.750 630.750 ;
        RECT 553.950 628.950 556.050 631.050 ;
        RECT 557.250 629.850 559.050 630.750 ;
        RECT 559.950 629.250 562.050 630.150 ;
        RECT 565.950 629.250 568.050 630.150 ;
        RECT 571.950 628.950 574.050 631.050 ;
        RECT 574.950 628.950 577.050 631.050 ;
        RECT 541.950 623.850 544.050 624.750 ;
        RECT 547.950 622.950 550.050 625.050 ;
        RECT 538.950 619.500 541.050 621.600 ;
        RECT 554.400 616.050 555.450 628.950 ;
        RECT 575.400 628.050 576.450 628.950 ;
        RECT 559.950 625.950 562.050 628.050 ;
        RECT 563.250 626.250 564.750 627.150 ;
        RECT 565.950 625.950 568.050 628.050 ;
        RECT 574.950 625.950 577.050 628.050 ;
        RECT 560.400 625.050 561.450 625.950 ;
        RECT 559.950 622.950 562.050 625.050 ;
        RECT 562.950 622.950 565.050 625.050 ;
        RECT 574.950 623.850 577.050 624.750 ;
        RECT 532.950 613.950 535.050 616.050 ;
        RECT 553.950 613.950 556.050 616.050 ;
        RECT 529.950 610.950 532.050 613.050 ;
        RECT 517.950 601.950 520.050 604.050 ;
        RECT 520.950 601.950 523.050 604.050 ;
        RECT 529.950 603.450 532.050 604.050 ;
        RECT 533.400 603.450 534.450 613.950 ;
        RECT 547.950 610.950 550.050 613.050 ;
        RECT 538.950 605.400 541.050 607.500 ;
        RECT 529.950 602.400 534.450 603.450 ;
        RECT 529.950 601.950 532.050 602.400 ;
        RECT 535.950 602.250 538.050 603.150 ;
        RECT 521.400 601.050 522.450 601.950 ;
        RECT 511.950 598.950 514.050 601.050 ;
        RECT 514.950 598.950 517.050 601.050 ;
        RECT 518.250 599.850 519.750 600.750 ;
        RECT 520.950 598.950 523.050 601.050 ;
        RECT 526.950 599.250 529.050 600.150 ;
        RECT 529.950 599.850 532.050 600.750 ;
        RECT 535.950 598.950 538.050 601.050 ;
        RECT 508.950 559.950 511.050 562.050 ;
        RECT 487.950 557.250 489.750 558.150 ;
        RECT 490.950 556.950 493.050 559.050 ;
        RECT 493.950 556.950 496.050 559.050 ;
        RECT 496.950 556.950 499.050 559.050 ;
        RECT 499.950 556.950 502.050 559.050 ;
        RECT 505.950 556.950 508.050 559.050 ;
        RECT 509.250 557.250 511.050 558.150 ;
        RECT 487.950 553.950 490.050 556.050 ;
        RECT 491.250 554.850 493.050 555.750 ;
        RECT 493.950 554.250 496.050 555.150 ;
        RECT 496.950 554.850 499.050 555.750 ;
        RECT 499.950 554.850 502.050 555.750 ;
        RECT 502.950 554.250 505.050 555.150 ;
        RECT 505.950 554.850 507.750 555.750 ;
        RECT 508.950 553.950 511.050 556.050 ;
        RECT 493.950 550.950 496.050 553.050 ;
        RECT 502.950 550.950 505.050 553.050 ;
        RECT 505.950 550.950 508.050 553.050 ;
        RECT 494.400 544.050 495.450 550.950 ;
        RECT 503.400 550.050 504.450 550.950 ;
        RECT 502.950 547.950 505.050 550.050 ;
        RECT 493.950 541.950 496.050 544.050 ;
        RECT 490.950 532.950 493.050 535.050 ;
        RECT 502.950 532.950 505.050 535.050 ;
        RECT 472.950 529.950 475.050 532.050 ;
        RECT 481.950 529.950 484.050 532.050 ;
        RECT 484.950 529.950 487.050 532.050 ;
        RECT 469.950 526.950 472.050 529.050 ;
        RECT 466.950 514.500 469.050 516.600 ;
        RECT 463.950 490.950 466.050 493.050 ;
        RECT 451.950 488.250 454.050 489.150 ;
        RECT 464.400 487.050 465.450 490.950 ;
        RECT 470.400 490.050 471.450 526.950 ;
        RECT 473.400 499.050 474.450 529.950 ;
        RECT 482.400 529.050 483.450 529.950 ;
        RECT 475.950 526.950 478.050 529.050 ;
        RECT 481.950 526.950 484.050 529.050 ;
        RECT 485.250 527.250 486.750 528.150 ;
        RECT 487.950 526.950 490.050 529.050 ;
        RECT 476.400 523.050 477.450 526.950 ;
        RECT 478.950 523.950 481.050 526.050 ;
        RECT 482.250 524.850 483.750 525.750 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 488.250 524.850 490.050 525.750 ;
        RECT 475.950 520.950 478.050 523.050 ;
        RECT 478.950 521.850 481.050 522.750 ;
        RECT 485.400 520.050 486.450 523.950 ;
        RECT 484.950 517.950 487.050 520.050 ;
        RECT 472.950 496.950 475.050 499.050 ;
        RECT 491.400 496.050 492.450 532.950 ;
        RECT 503.400 532.050 504.450 532.950 ;
        RECT 496.950 529.950 499.050 532.050 ;
        RECT 499.950 529.950 502.050 532.050 ;
        RECT 502.950 529.950 505.050 532.050 ;
        RECT 500.400 529.050 501.450 529.950 ;
        RECT 506.400 529.050 507.450 550.950 ;
        RECT 509.400 547.050 510.450 553.950 ;
        RECT 508.950 544.950 511.050 547.050 ;
        RECT 512.400 544.050 513.450 598.950 ;
        RECT 514.950 596.850 517.050 597.750 ;
        RECT 520.950 596.850 523.050 597.750 ;
        RECT 526.950 595.950 529.050 598.050 ;
        RECT 536.400 592.050 537.450 598.950 ;
        RECT 539.550 593.400 540.750 605.400 ;
        RECT 548.400 601.050 549.450 610.950 ;
        RECT 550.950 604.950 553.050 607.050 ;
        RECT 559.950 605.400 562.050 607.500 ;
        RECT 547.950 598.950 550.050 601.050 ;
        RECT 547.950 596.850 550.050 597.750 ;
        RECT 551.400 595.050 552.450 604.950 ;
        RECT 553.950 598.950 556.050 601.050 ;
        RECT 553.950 596.850 556.050 597.750 ;
        RECT 535.950 589.950 538.050 592.050 ;
        RECT 538.950 591.300 541.050 593.400 ;
        RECT 550.950 592.950 553.050 595.050 ;
        RECT 539.550 587.700 540.750 591.300 ;
        RECT 560.400 588.600 561.600 605.400 ;
        RECT 563.400 604.050 564.450 622.950 ;
        RECT 578.550 621.600 579.750 633.600 ;
        RECT 581.400 628.050 582.450 667.950 ;
        RECT 589.950 631.950 592.050 634.050 ;
        RECT 586.950 629.250 589.050 630.150 ;
        RECT 580.950 625.950 583.050 628.050 ;
        RECT 586.950 625.950 589.050 628.050 ;
        RECT 590.400 627.450 591.450 631.950 ;
        RECT 592.950 629.250 595.050 630.150 ;
        RECT 592.950 627.450 595.050 628.050 ;
        RECT 590.400 626.400 595.050 627.450 ;
        RECT 592.950 625.950 595.050 626.400 ;
        RECT 577.950 619.500 580.050 621.600 ;
        RECT 581.400 613.050 582.450 625.950 ;
        RECT 587.400 622.050 588.450 625.950 ;
        RECT 586.950 619.950 589.050 622.050 ;
        RECT 580.950 610.950 583.050 613.050 ;
        RECT 577.950 604.950 580.050 607.050 ;
        RECT 589.950 604.950 592.050 607.050 ;
        RECT 578.400 604.050 579.450 604.950 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 577.950 601.950 580.050 604.050 ;
        RECT 586.950 601.950 589.050 604.050 ;
        RECT 590.400 601.050 591.450 604.950 ;
        RECT 596.400 603.450 597.450 676.950 ;
        RECT 622.950 673.950 625.050 676.050 ;
        RECT 631.950 675.450 634.050 676.050 ;
        RECT 629.400 674.400 634.050 675.450 ;
        RECT 616.950 672.450 619.050 673.050 ;
        RECT 601.950 671.250 604.050 672.150 ;
        RECT 614.400 671.400 619.050 672.450 ;
        RECT 610.950 668.850 613.050 669.750 ;
        RECT 614.400 667.050 615.450 671.400 ;
        RECT 616.950 670.950 619.050 671.400 ;
        RECT 623.400 670.050 624.450 673.950 ;
        RECT 616.950 668.850 619.050 669.750 ;
        RECT 619.950 668.250 621.750 669.150 ;
        RECT 622.950 667.950 625.050 670.050 ;
        RECT 626.250 668.250 628.050 669.150 ;
        RECT 613.950 664.950 616.050 667.050 ;
        RECT 619.950 664.950 622.050 667.050 ;
        RECT 623.250 665.850 624.750 666.750 ;
        RECT 625.950 664.950 628.050 667.050 ;
        RECT 614.400 646.050 615.450 664.950 ;
        RECT 620.400 646.050 621.450 664.950 ;
        RECT 629.400 661.050 630.450 674.400 ;
        RECT 631.950 673.950 634.050 674.400 ;
        RECT 649.950 673.950 652.050 676.050 ;
        RECT 658.950 674.250 661.050 675.150 ;
        RECT 631.950 671.850 634.050 672.750 ;
        RECT 634.950 671.250 637.050 672.150 ;
        RECT 640.950 670.950 643.050 673.050 ;
        RECT 644.250 671.250 645.750 672.150 ;
        RECT 646.950 670.950 649.050 673.050 ;
        RECT 650.400 670.050 651.450 673.950 ;
        RECT 658.950 670.950 661.050 673.050 ;
        RECT 634.950 667.950 637.050 670.050 ;
        RECT 640.950 668.850 642.750 669.750 ;
        RECT 643.950 667.950 646.050 670.050 ;
        RECT 647.250 668.850 648.750 669.750 ;
        RECT 649.950 667.950 652.050 670.050 ;
        RECT 643.950 664.950 646.050 667.050 ;
        RECT 649.950 665.850 652.050 666.750 ;
        RECT 628.950 658.950 631.050 661.050 ;
        RECT 604.950 643.950 607.050 646.050 ;
        RECT 613.950 643.950 616.050 646.050 ;
        RECT 619.950 643.950 622.050 646.050 ;
        RECT 598.950 638.400 601.050 640.500 ;
        RECT 599.400 621.600 600.600 638.400 ;
        RECT 598.950 619.500 601.050 621.600 ;
        RECT 605.400 616.050 606.450 643.950 ;
        RECT 629.400 637.050 630.450 658.950 ;
        RECT 628.950 634.950 631.050 637.050 ;
        RECT 631.950 634.950 634.050 637.050 ;
        RECT 619.950 631.950 622.050 634.050 ;
        RECT 607.950 629.250 610.050 630.150 ;
        RECT 613.950 629.250 616.050 630.150 ;
        RECT 607.950 625.950 610.050 628.050 ;
        RECT 611.250 626.250 612.750 627.150 ;
        RECT 613.950 625.950 616.050 628.050 ;
        RECT 620.400 627.450 621.450 631.950 ;
        RECT 632.400 631.050 633.450 634.950 ;
        RECT 622.950 629.250 624.750 630.150 ;
        RECT 625.950 628.950 628.050 631.050 ;
        RECT 631.950 628.950 634.050 631.050 ;
        RECT 634.950 629.250 637.050 630.150 ;
        RECT 640.950 629.250 643.050 630.150 ;
        RECT 622.950 627.450 625.050 628.050 ;
        RECT 620.400 626.400 625.050 627.450 ;
        RECT 626.250 626.850 628.050 627.750 ;
        RECT 622.950 625.950 625.050 626.400 ;
        RECT 628.950 626.250 631.050 627.150 ;
        RECT 631.950 626.850 634.050 627.750 ;
        RECT 634.950 625.950 637.050 628.050 ;
        RECT 610.950 622.950 613.050 625.050 ;
        RECT 604.950 613.950 607.050 616.050 ;
        RECT 614.400 610.050 615.450 625.950 ;
        RECT 628.950 622.950 631.050 625.050 ;
        RECT 629.400 610.050 630.450 622.950 ;
        RECT 635.400 618.450 636.450 625.950 ;
        RECT 635.400 617.400 639.450 618.450 ;
        RECT 631.950 613.950 634.050 616.050 ;
        RECT 634.950 613.950 637.050 616.050 ;
        RECT 604.950 607.950 607.050 610.050 ;
        RECT 610.950 607.950 613.050 610.050 ;
        RECT 613.950 607.950 616.050 610.050 ;
        RECT 619.950 607.950 622.050 610.050 ;
        RECT 628.950 607.950 631.050 610.050 ;
        RECT 593.400 602.400 597.450 603.450 ;
        RECT 571.950 598.950 574.050 601.050 ;
        RECT 575.250 599.250 577.050 600.150 ;
        RECT 577.950 599.850 580.050 600.750 ;
        RECT 580.950 599.250 583.050 600.150 ;
        RECT 583.950 598.950 586.050 601.050 ;
        RECT 587.250 599.850 588.750 600.750 ;
        RECT 589.950 598.950 592.050 601.050 ;
        RECT 571.950 596.850 573.750 597.750 ;
        RECT 574.950 595.950 577.050 598.050 ;
        RECT 577.950 595.950 580.050 598.050 ;
        RECT 580.950 595.950 583.050 598.050 ;
        RECT 583.950 596.850 586.050 597.750 ;
        RECT 589.950 596.850 592.050 597.750 ;
        RECT 578.400 592.050 579.450 595.950 ;
        RECT 577.950 589.950 580.050 592.050 ;
        RECT 581.400 589.050 582.450 595.950 ;
        RECT 538.950 585.600 541.050 587.700 ;
        RECT 559.950 586.500 562.050 588.600 ;
        RECT 571.950 586.950 574.050 589.050 ;
        RECT 580.950 586.950 583.050 589.050 ;
        RECT 550.950 574.950 553.050 577.050 ;
        RECT 526.950 562.950 529.050 565.050 ;
        RECT 541.950 562.950 544.050 565.050 ;
        RECT 517.950 558.450 520.050 559.050 ;
        RECT 517.950 557.400 522.450 558.450 ;
        RECT 517.950 556.950 520.050 557.400 ;
        RECT 514.950 554.250 517.050 555.150 ;
        RECT 517.950 554.850 520.050 555.750 ;
        RECT 514.950 550.950 517.050 553.050 ;
        RECT 517.950 547.950 520.050 550.050 ;
        RECT 511.950 541.950 514.050 544.050 ;
        RECT 514.950 541.950 517.050 544.050 ;
        RECT 508.950 532.950 511.050 535.050 ;
        RECT 509.400 532.050 510.450 532.950 ;
        RECT 515.400 532.050 516.450 541.950 ;
        RECT 508.950 529.950 511.050 532.050 ;
        RECT 511.950 529.950 514.050 532.050 ;
        RECT 514.950 529.950 517.050 532.050 ;
        RECT 493.950 527.250 496.050 528.150 ;
        RECT 496.950 527.850 499.050 528.750 ;
        RECT 499.950 526.950 502.050 529.050 ;
        RECT 503.250 527.850 504.750 528.750 ;
        RECT 505.950 528.450 508.050 529.050 ;
        RECT 505.950 527.400 510.450 528.450 ;
        RECT 511.950 527.850 514.050 528.750 ;
        RECT 505.950 526.950 508.050 527.400 ;
        RECT 509.400 526.050 510.450 527.400 ;
        RECT 514.950 527.250 517.050 528.150 ;
        RECT 493.950 523.950 496.050 526.050 ;
        RECT 499.950 524.850 502.050 525.750 ;
        RECT 505.950 524.850 508.050 525.750 ;
        RECT 508.950 523.950 511.050 526.050 ;
        RECT 514.950 523.950 517.050 526.050 ;
        RECT 494.400 523.050 495.450 523.950 ;
        RECT 493.950 520.950 496.050 523.050 ;
        RECT 511.950 520.950 514.050 523.050 ;
        RECT 493.950 508.950 496.050 511.050 ;
        RECT 490.950 493.950 493.050 496.050 ;
        RECT 481.950 490.950 484.050 493.050 ;
        RECT 494.400 492.450 495.450 508.950 ;
        RECT 491.400 491.400 495.450 492.450 ;
        RECT 466.950 488.250 469.050 489.150 ;
        RECT 469.950 487.950 472.050 490.050 ;
        RECT 482.400 487.050 483.450 490.950 ;
        RECT 487.950 488.250 490.050 489.150 ;
        RECT 451.950 484.950 454.050 487.050 ;
        RECT 455.250 485.250 456.750 486.150 ;
        RECT 457.950 484.950 460.050 487.050 ;
        RECT 461.250 485.250 463.050 486.150 ;
        RECT 463.950 484.950 466.050 487.050 ;
        RECT 466.950 484.950 469.050 487.050 ;
        RECT 470.250 485.250 471.750 486.150 ;
        RECT 472.950 484.950 475.050 487.050 ;
        RECT 476.250 485.250 478.050 486.150 ;
        RECT 478.950 485.250 480.750 486.150 ;
        RECT 481.950 484.950 484.050 487.050 ;
        RECT 485.250 485.250 486.750 486.150 ;
        RECT 487.950 484.950 490.050 487.050 ;
        RECT 454.950 481.950 457.050 484.050 ;
        RECT 458.250 482.850 459.750 483.750 ;
        RECT 460.950 481.950 463.050 484.050 ;
        RECT 454.950 478.950 457.050 481.050 ;
        RECT 455.400 457.050 456.450 478.950 ;
        RECT 461.400 478.050 462.450 481.950 ;
        RECT 464.400 481.050 465.450 484.950 ;
        RECT 467.400 484.050 468.450 484.950 ;
        RECT 466.950 481.950 469.050 484.050 ;
        RECT 469.950 481.950 472.050 484.050 ;
        RECT 473.250 482.850 474.750 483.750 ;
        RECT 475.950 481.950 478.050 484.050 ;
        RECT 478.950 481.950 481.050 484.050 ;
        RECT 482.250 482.850 483.750 483.750 ;
        RECT 484.950 481.950 487.050 484.050 ;
        RECT 476.400 481.050 477.450 481.950 ;
        RECT 463.950 478.950 466.050 481.050 ;
        RECT 475.950 478.950 478.050 481.050 ;
        RECT 460.950 475.950 463.050 478.050 ;
        RECT 457.950 457.950 460.050 460.050 ;
        RECT 461.400 457.050 462.450 475.950 ;
        RECT 466.950 460.950 469.050 463.050 ;
        RECT 472.950 460.950 475.050 463.050 ;
        RECT 463.950 457.950 466.050 460.050 ;
        RECT 454.950 454.950 457.050 457.050 ;
        RECT 458.250 455.850 459.750 456.750 ;
        RECT 460.950 454.950 463.050 457.050 ;
        RECT 454.950 452.850 457.050 453.750 ;
        RECT 460.950 452.850 463.050 453.750 ;
        RECT 448.950 448.950 451.050 451.050 ;
        RECT 454.950 448.950 457.050 451.050 ;
        RECT 443.250 443.700 444.450 447.300 ;
        RECT 445.950 445.950 448.050 448.050 ;
        RECT 442.950 441.600 445.050 443.700 ;
        RECT 448.950 427.950 451.050 430.050 ;
        RECT 442.950 424.950 445.050 427.050 ;
        RECT 439.950 422.400 442.050 424.500 ;
        RECT 436.950 415.950 439.050 418.050 ;
        RECT 430.950 406.950 433.050 409.050 ;
        RECT 406.950 403.950 409.050 406.050 ;
        RECT 418.950 403.950 421.050 406.050 ;
        RECT 394.950 400.950 397.050 403.050 ;
        RECT 395.400 385.050 396.450 400.950 ;
        RECT 403.950 388.950 406.050 391.050 ;
        RECT 388.950 384.450 391.050 385.050 ;
        RECT 388.950 383.400 393.450 384.450 ;
        RECT 388.950 382.950 391.050 383.400 ;
        RECT 385.950 380.250 388.050 381.150 ;
        RECT 388.950 380.850 391.050 381.750 ;
        RECT 385.950 376.950 388.050 379.050 ;
        RECT 382.950 373.950 385.050 376.050 ;
        RECT 385.950 373.950 388.050 376.050 ;
        RECT 376.950 349.950 379.050 352.050 ;
        RECT 376.950 347.250 379.050 348.150 ;
        RECT 352.950 343.950 355.050 346.050 ;
        RECT 358.950 343.950 361.050 346.050 ;
        RECT 373.950 344.250 375.750 345.150 ;
        RECT 376.950 343.950 379.050 346.050 ;
        RECT 380.250 344.250 381.750 345.150 ;
        RECT 382.950 343.950 385.050 346.050 ;
        RECT 346.950 341.250 348.750 342.150 ;
        RECT 349.950 340.950 352.050 343.050 ;
        RECT 355.950 340.950 358.050 343.050 ;
        RECT 343.950 337.950 346.050 340.050 ;
        RECT 346.950 337.950 349.050 340.050 ;
        RECT 350.250 338.850 352.050 339.750 ;
        RECT 352.950 338.250 355.050 339.150 ;
        RECT 355.950 338.850 358.050 339.750 ;
        RECT 337.950 335.850 340.050 336.750 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 352.950 334.950 355.050 337.050 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 334.950 331.500 337.050 333.600 ;
        RECT 337.950 331.950 340.050 334.050 ;
        RECT 334.950 322.950 337.050 325.050 ;
        RECT 331.950 316.950 334.050 319.050 ;
        RECT 331.950 311.250 334.050 312.150 ;
        RECT 331.950 309.450 334.050 310.050 ;
        RECT 329.400 308.400 334.050 309.450 ;
        RECT 316.950 305.850 319.050 306.750 ;
        RECT 323.400 292.050 324.450 307.950 ;
        RECT 310.950 289.950 313.050 292.050 ;
        RECT 313.950 289.950 316.050 292.050 ;
        RECT 322.950 289.950 325.050 292.050 ;
        RECT 310.950 271.950 313.050 274.050 ;
        RECT 301.950 269.250 304.050 270.150 ;
        RECT 307.950 269.250 310.050 270.150 ;
        RECT 301.950 265.950 304.050 268.050 ;
        RECT 307.950 267.450 310.050 268.050 ;
        RECT 311.400 267.450 312.450 271.950 ;
        RECT 307.950 266.400 312.450 267.450 ;
        RECT 307.950 265.950 310.050 266.400 ;
        RECT 302.400 244.050 303.450 265.950 ;
        RECT 304.950 244.950 307.050 247.050 ;
        RECT 301.950 241.950 304.050 244.050 ;
        RECT 305.400 241.050 306.450 244.950 ;
        RECT 314.400 241.050 315.450 289.950 ;
        RECT 316.950 279.300 319.050 281.400 ;
        RECT 329.400 280.050 330.450 308.400 ;
        RECT 331.950 307.950 334.050 308.400 ;
        RECT 335.400 298.050 336.450 322.950 ;
        RECT 334.950 295.950 337.050 298.050 ;
        RECT 317.250 275.700 318.450 279.300 ;
        RECT 328.950 277.950 331.050 280.050 ;
        RECT 316.950 273.600 319.050 275.700 ;
        RECT 322.950 274.950 325.050 277.050 ;
        RECT 317.250 261.600 318.450 273.600 ;
        RECT 319.950 265.950 322.050 268.050 ;
        RECT 319.950 263.850 322.050 264.750 ;
        RECT 316.950 259.500 319.050 261.600 ;
        RECT 323.400 247.050 324.450 274.950 ;
        RECT 329.400 274.050 330.450 277.950 ;
        RECT 328.950 271.950 331.050 274.050 ;
        RECT 338.400 271.050 339.450 331.950 ;
        RECT 343.950 319.950 346.050 322.050 ;
        RECT 340.950 313.950 343.050 316.050 ;
        RECT 341.400 277.050 342.450 313.950 ;
        RECT 340.950 274.950 343.050 277.050 ;
        RECT 325.950 268.950 328.050 271.050 ;
        RECT 328.950 269.250 331.050 270.150 ;
        RECT 334.950 269.250 337.050 270.150 ;
        RECT 337.950 268.950 340.050 271.050 ;
        RECT 340.950 268.950 343.050 271.050 ;
        RECT 322.950 244.950 325.050 247.050 ;
        RECT 326.400 244.050 327.450 268.950 ;
        RECT 328.950 265.950 331.050 268.050 ;
        RECT 332.250 266.250 333.750 267.150 ;
        RECT 334.950 265.950 337.050 268.050 ;
        RECT 337.950 266.250 340.050 267.150 ;
        RECT 340.950 266.850 343.050 267.750 ;
        RECT 322.950 241.950 325.050 244.050 ;
        RECT 325.950 241.950 328.050 244.050 ;
        RECT 329.400 243.450 330.450 265.950 ;
        RECT 331.950 262.950 334.050 265.050 ;
        RECT 335.400 264.450 336.450 265.950 ;
        RECT 337.950 264.450 340.050 265.050 ;
        RECT 335.400 263.400 342.450 264.450 ;
        RECT 337.950 262.950 340.050 263.400 ;
        RECT 331.950 243.450 334.050 244.050 ;
        RECT 329.400 242.400 334.050 243.450 ;
        RECT 331.950 241.950 334.050 242.400 ;
        RECT 323.400 241.050 324.450 241.950 ;
        RECT 301.950 238.950 304.050 241.050 ;
        RECT 304.950 238.950 307.050 241.050 ;
        RECT 313.950 238.950 316.050 241.050 ;
        RECT 319.950 238.950 322.050 241.050 ;
        RECT 322.950 238.950 325.050 241.050 ;
        RECT 326.250 239.250 327.750 240.150 ;
        RECT 328.950 238.950 331.050 241.050 ;
        RECT 331.950 239.850 334.050 240.750 ;
        RECT 341.400 240.450 342.450 263.400 ;
        RECT 344.400 259.050 345.450 319.950 ;
        RECT 352.950 311.250 355.050 312.150 ;
        RECT 349.950 307.950 352.050 310.050 ;
        RECT 350.400 274.050 351.450 307.950 ;
        RECT 356.400 298.050 357.450 334.950 ;
        RECT 359.400 316.050 360.450 343.950 ;
        RECT 361.950 341.250 363.750 342.150 ;
        RECT 364.950 340.950 367.050 343.050 ;
        RECT 370.950 340.950 373.050 343.050 ;
        RECT 373.950 340.950 376.050 343.050 ;
        RECT 379.950 340.950 382.050 343.050 ;
        RECT 383.250 341.850 385.050 342.750 ;
        RECT 361.950 337.950 364.050 340.050 ;
        RECT 365.250 338.850 367.050 339.750 ;
        RECT 367.950 338.250 370.050 339.150 ;
        RECT 370.950 338.850 373.050 339.750 ;
        RECT 367.950 336.450 370.050 337.050 ;
        RECT 374.400 336.450 375.450 340.950 ;
        RECT 380.400 337.050 381.450 340.950 ;
        RECT 386.400 340.050 387.450 373.950 ;
        RECT 392.400 349.050 393.450 383.400 ;
        RECT 394.950 382.950 397.050 385.050 ;
        RECT 398.250 383.250 399.750 384.150 ;
        RECT 400.950 382.950 403.050 385.050 ;
        RECT 404.400 382.050 405.450 388.950 ;
        RECT 394.950 380.850 396.750 381.750 ;
        RECT 397.950 379.950 400.050 382.050 ;
        RECT 401.250 380.850 402.750 381.750 ;
        RECT 403.950 379.950 406.050 382.050 ;
        RECT 398.400 376.050 399.450 379.950 ;
        RECT 403.950 377.850 406.050 378.750 ;
        RECT 407.400 376.050 408.450 403.950 ;
        RECT 421.950 387.450 424.050 388.050 ;
        RECT 419.400 386.400 424.050 387.450 ;
        RECT 419.400 385.050 420.450 386.400 ;
        RECT 421.950 385.950 424.050 386.400 ;
        RECT 424.950 385.950 427.050 388.050 ;
        RECT 427.950 385.950 430.050 388.050 ;
        RECT 433.950 385.950 436.050 388.050 ;
        RECT 425.400 385.050 426.450 385.950 ;
        RECT 409.950 382.950 412.050 385.050 ;
        RECT 418.950 382.950 421.050 385.050 ;
        RECT 421.950 383.850 423.750 384.750 ;
        RECT 424.950 382.950 427.050 385.050 ;
        RECT 410.400 378.450 411.450 382.950 ;
        RECT 412.950 380.250 414.750 381.150 ;
        RECT 415.950 379.950 418.050 382.050 ;
        RECT 419.250 380.250 421.050 381.150 ;
        RECT 424.950 380.850 427.050 381.750 ;
        RECT 428.400 379.050 429.450 385.950 ;
        RECT 430.950 383.250 433.050 384.150 ;
        RECT 430.950 379.950 433.050 382.050 ;
        RECT 412.950 378.450 415.050 379.050 ;
        RECT 410.400 377.400 415.050 378.450 ;
        RECT 416.250 377.850 417.750 378.750 ;
        RECT 412.950 376.950 415.050 377.400 ;
        RECT 418.950 376.950 421.050 379.050 ;
        RECT 427.950 376.950 430.050 379.050 ;
        RECT 431.400 376.050 432.450 379.950 ;
        RECT 397.950 373.950 400.050 376.050 ;
        RECT 406.950 373.950 409.050 376.050 ;
        RECT 421.950 373.950 424.050 376.050 ;
        RECT 430.950 373.950 433.050 376.050 ;
        RECT 394.950 352.950 397.050 355.050 ;
        RECT 391.950 346.950 394.050 349.050 ;
        RECT 395.400 346.050 396.450 352.950 ;
        RECT 400.950 349.950 403.050 352.050 ;
        RECT 409.950 351.300 412.050 353.400 ;
        RECT 391.950 343.950 394.050 346.050 ;
        RECT 394.950 343.950 397.050 346.050 ;
        RECT 388.950 341.250 391.050 342.150 ;
        RECT 385.950 337.950 388.050 340.050 ;
        RECT 388.950 339.450 391.050 340.050 ;
        RECT 392.400 339.450 393.450 343.950 ;
        RECT 394.950 341.850 397.050 342.750 ;
        RECT 397.950 341.250 400.050 342.150 ;
        RECT 388.950 338.400 393.450 339.450 ;
        RECT 388.950 337.950 391.050 338.400 ;
        RECT 397.950 337.950 400.050 340.050 ;
        RECT 367.950 335.400 375.450 336.450 ;
        RECT 367.950 334.950 370.050 335.400 ;
        RECT 367.950 328.950 370.050 331.050 ;
        RECT 358.950 313.950 361.050 316.050 ;
        RECT 358.950 308.250 360.750 309.150 ;
        RECT 361.950 307.950 364.050 310.050 ;
        RECT 365.250 308.250 367.050 309.150 ;
        RECT 358.950 304.950 361.050 307.050 ;
        RECT 362.250 305.850 363.750 306.750 ;
        RECT 364.950 306.450 367.050 307.050 ;
        RECT 368.400 306.450 369.450 328.950 ;
        RECT 374.400 313.050 375.450 335.400 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 391.950 334.950 394.050 337.050 ;
        RECT 379.950 322.950 382.050 325.050 ;
        RECT 388.950 322.950 391.050 325.050 ;
        RECT 373.950 310.950 376.050 313.050 ;
        RECT 373.950 308.850 376.050 309.750 ;
        RECT 376.950 308.250 379.050 309.150 ;
        RECT 364.950 305.400 369.450 306.450 ;
        RECT 364.950 304.950 367.050 305.400 ;
        RECT 376.950 304.950 379.050 307.050 ;
        RECT 355.950 295.950 358.050 298.050 ;
        RECT 359.400 292.050 360.450 304.950 ;
        RECT 377.400 295.050 378.450 304.950 ;
        RECT 376.950 292.950 379.050 295.050 ;
        RECT 358.950 289.950 361.050 292.050 ;
        RECT 358.950 277.950 361.050 280.050 ;
        RECT 349.950 271.950 352.050 274.050 ;
        RECT 355.950 272.250 358.050 273.150 ;
        RECT 346.950 269.250 348.750 270.150 ;
        RECT 349.950 268.950 352.050 271.050 ;
        RECT 353.250 269.250 354.750 270.150 ;
        RECT 355.950 268.950 358.050 271.050 ;
        RECT 346.950 265.950 349.050 268.050 ;
        RECT 350.250 266.850 351.750 267.750 ;
        RECT 352.950 265.950 355.050 268.050 ;
        RECT 347.400 264.450 348.450 265.950 ;
        RECT 347.400 263.400 351.450 264.450 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 346.950 245.400 349.050 247.500 ;
        RECT 343.950 242.250 346.050 243.150 ;
        RECT 343.950 240.450 346.050 241.050 ;
        RECT 334.950 239.250 337.050 240.150 ;
        RECT 341.400 239.400 346.050 240.450 ;
        RECT 343.950 238.950 346.050 239.400 ;
        RECT 302.400 238.050 303.450 238.950 ;
        RECT 301.950 235.950 304.050 238.050 ;
        RECT 307.950 235.950 310.050 238.050 ;
        RECT 311.250 236.250 313.050 237.150 ;
        RECT 314.400 235.050 315.450 238.950 ;
        RECT 320.400 238.050 321.450 238.950 ;
        RECT 316.950 235.950 319.050 238.050 ;
        RECT 319.950 235.950 322.050 238.050 ;
        RECT 323.250 236.850 324.750 237.750 ;
        RECT 325.950 235.950 328.050 238.050 ;
        RECT 329.250 236.850 331.050 237.750 ;
        RECT 334.950 235.950 337.050 238.050 ;
        RECT 295.950 232.950 298.050 235.050 ;
        RECT 298.950 232.950 301.050 235.050 ;
        RECT 301.950 233.850 303.750 234.750 ;
        RECT 304.950 232.950 307.050 235.050 ;
        RECT 308.250 233.850 309.750 234.750 ;
        RECT 310.950 232.950 313.050 235.050 ;
        RECT 313.950 232.950 316.050 235.050 ;
        RECT 298.950 229.950 301.050 232.050 ;
        RECT 304.950 230.850 307.050 231.750 ;
        RECT 311.400 231.450 312.450 232.950 ;
        RECT 317.400 232.050 318.450 235.950 ;
        RECT 326.400 235.050 327.450 235.950 ;
        RECT 319.950 233.850 322.050 234.750 ;
        RECT 325.950 232.950 328.050 235.050 ;
        RECT 347.550 233.400 348.750 245.400 ;
        RECT 350.400 235.050 351.450 263.400 ;
        RECT 353.400 262.050 354.450 265.950 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 352.950 244.950 355.050 247.050 ;
        RECT 313.950 231.450 316.050 232.050 ;
        RECT 311.400 230.400 316.050 231.450 ;
        RECT 313.950 229.950 316.050 230.400 ;
        RECT 316.950 229.950 319.050 232.050 ;
        RECT 346.950 231.300 349.050 233.400 ;
        RECT 349.950 232.950 352.050 235.050 ;
        RECT 299.400 202.050 300.450 229.950 ;
        RECT 347.550 227.700 348.750 231.300 ;
        RECT 346.950 225.600 349.050 227.700 ;
        RECT 307.950 205.950 310.050 208.050 ;
        RECT 313.950 205.950 316.050 208.050 ;
        RECT 298.950 199.950 301.050 202.050 ;
        RECT 304.950 200.250 307.050 201.150 ;
        RECT 295.950 197.250 297.750 198.150 ;
        RECT 298.950 196.950 301.050 199.050 ;
        RECT 302.250 197.250 303.750 198.150 ;
        RECT 304.950 196.950 307.050 199.050 ;
        RECT 295.950 193.950 298.050 196.050 ;
        RECT 299.250 194.850 300.750 195.750 ;
        RECT 301.950 193.950 304.050 196.050 ;
        RECT 296.400 193.050 297.450 193.950 ;
        RECT 295.950 190.950 298.050 193.050 ;
        RECT 289.950 187.950 292.050 190.050 ;
        RECT 292.950 187.950 295.050 190.050 ;
        RECT 287.400 167.400 291.450 168.450 ;
        RECT 268.950 164.250 270.750 165.150 ;
        RECT 271.950 163.950 274.050 166.050 ;
        RECT 275.250 164.250 277.050 165.150 ;
        RECT 277.950 163.950 280.050 166.050 ;
        RECT 283.950 163.950 286.050 166.050 ;
        RECT 287.250 164.250 289.050 165.150 ;
        RECT 268.950 160.950 271.050 163.050 ;
        RECT 272.250 161.850 273.750 162.750 ;
        RECT 274.950 160.950 277.050 163.050 ;
        RECT 277.950 161.850 279.750 162.750 ;
        RECT 280.950 160.950 283.050 163.050 ;
        RECT 284.250 161.850 285.750 162.750 ;
        RECT 286.950 160.950 289.050 163.050 ;
        RECT 269.400 160.050 270.450 160.950 ;
        RECT 275.400 160.050 276.450 160.950 ;
        RECT 290.400 160.050 291.450 167.400 ;
        RECT 296.400 166.050 297.450 190.950 ;
        RECT 302.400 187.050 303.450 193.950 ;
        RECT 301.950 184.950 304.050 187.050 ;
        RECT 308.400 172.050 309.450 205.950 ;
        RECT 314.400 199.050 315.450 205.950 ;
        RECT 322.950 203.250 325.050 204.150 ;
        RECT 353.400 202.050 354.450 244.950 ;
        RECT 355.950 240.450 358.050 241.050 ;
        RECT 359.400 240.450 360.450 277.950 ;
        RECT 380.400 273.450 381.450 322.950 ;
        RECT 385.950 313.950 388.050 316.050 ;
        RECT 389.400 313.050 390.450 322.950 ;
        RECT 382.950 310.950 385.050 313.050 ;
        RECT 385.950 311.850 387.750 312.750 ;
        RECT 388.950 310.950 391.050 313.050 ;
        RECT 382.950 308.850 385.050 309.750 ;
        RECT 388.950 308.850 391.050 309.750 ;
        RECT 392.400 301.050 393.450 334.950 ;
        RECT 398.400 334.050 399.450 337.950 ;
        RECT 397.950 331.950 400.050 334.050 ;
        RECT 401.400 325.050 402.450 349.950 ;
        RECT 410.550 347.700 411.750 351.300 ;
        RECT 409.950 345.600 412.050 347.700 ;
        RECT 406.950 339.450 409.050 340.050 ;
        RECT 404.400 338.400 409.050 339.450 ;
        RECT 404.400 331.050 405.450 338.400 ;
        RECT 406.950 337.950 409.050 338.400 ;
        RECT 406.950 335.850 409.050 336.750 ;
        RECT 410.550 333.600 411.750 345.600 ;
        RECT 418.950 341.250 421.050 342.150 ;
        RECT 418.950 337.950 421.050 340.050 ;
        RECT 409.950 331.500 412.050 333.600 ;
        RECT 403.950 328.950 406.050 331.050 ;
        RECT 400.950 322.950 403.050 325.050 ;
        RECT 397.950 319.950 400.050 322.050 ;
        RECT 394.950 311.250 397.050 312.150 ;
        RECT 394.950 309.450 397.050 310.050 ;
        RECT 398.400 309.450 399.450 319.950 ;
        RECT 400.950 310.950 403.050 313.050 ;
        RECT 394.950 308.400 399.450 309.450 ;
        RECT 394.950 307.950 397.050 308.400 ;
        RECT 401.400 307.050 402.450 310.950 ;
        RECT 403.950 308.250 405.750 309.150 ;
        RECT 406.950 307.950 409.050 310.050 ;
        RECT 410.250 308.250 412.050 309.150 ;
        RECT 412.950 308.250 414.750 309.150 ;
        RECT 415.950 307.950 418.050 310.050 ;
        RECT 419.250 308.250 421.050 309.150 ;
        RECT 400.950 304.950 403.050 307.050 ;
        RECT 403.950 304.950 406.050 307.050 ;
        RECT 407.250 305.850 408.750 306.750 ;
        RECT 409.950 304.950 412.050 307.050 ;
        RECT 412.950 304.950 415.050 307.050 ;
        RECT 416.250 305.850 417.750 306.750 ;
        RECT 418.950 304.950 421.050 307.050 ;
        RECT 404.400 301.050 405.450 304.950 ;
        RECT 391.950 298.950 394.050 301.050 ;
        RECT 403.950 298.950 406.050 301.050 ;
        RECT 397.950 295.950 400.050 298.050 ;
        RECT 380.400 272.400 384.450 273.450 ;
        RECT 361.950 269.250 364.050 270.150 ;
        RECT 367.950 269.250 370.050 270.150 ;
        RECT 373.950 269.250 376.050 270.150 ;
        RECT 379.950 269.250 382.050 270.150 ;
        RECT 361.950 265.950 364.050 268.050 ;
        RECT 365.250 266.250 366.750 267.150 ;
        RECT 367.950 265.950 370.050 268.050 ;
        RECT 373.950 265.950 376.050 268.050 ;
        RECT 377.250 266.250 378.750 267.150 ;
        RECT 379.950 265.950 382.050 268.050 ;
        RECT 362.400 265.050 363.450 265.950 ;
        RECT 361.950 262.950 364.050 265.050 ;
        RECT 364.950 262.950 367.050 265.050 ;
        RECT 361.950 259.950 364.050 262.050 ;
        RECT 362.400 241.050 363.450 259.950 ;
        RECT 365.400 247.050 366.450 262.950 ;
        RECT 368.400 262.050 369.450 265.950 ;
        RECT 374.400 265.050 375.450 265.950 ;
        RECT 373.950 262.950 376.050 265.050 ;
        RECT 376.950 262.950 379.050 265.050 ;
        RECT 377.400 262.050 378.450 262.950 ;
        RECT 367.950 259.950 370.050 262.050 ;
        RECT 376.950 259.950 379.050 262.050 ;
        RECT 370.950 250.950 373.050 253.050 ;
        RECT 364.950 244.950 367.050 247.050 ;
        RECT 367.950 245.400 370.050 247.500 ;
        RECT 364.950 241.950 367.050 244.050 ;
        RECT 355.950 239.400 360.450 240.450 ;
        RECT 355.950 238.950 358.050 239.400 ;
        RECT 361.950 238.950 364.050 241.050 ;
        RECT 355.950 236.850 358.050 237.750 ;
        RECT 361.950 236.850 364.050 237.750 ;
        RECT 355.950 229.950 358.050 232.050 ;
        RECT 319.950 200.250 321.750 201.150 ;
        RECT 322.950 199.950 325.050 202.050 ;
        RECT 326.250 200.250 327.750 201.150 ;
        RECT 328.950 199.950 331.050 202.050 ;
        RECT 334.950 201.450 337.050 202.050 ;
        RECT 332.400 200.400 337.050 201.450 ;
        RECT 323.400 199.050 324.450 199.950 ;
        RECT 313.950 196.950 316.050 199.050 ;
        RECT 319.950 196.950 322.050 199.050 ;
        RECT 322.950 196.950 325.050 199.050 ;
        RECT 325.950 196.950 328.050 199.050 ;
        RECT 329.250 197.850 331.050 198.750 ;
        RECT 310.950 194.250 313.050 195.150 ;
        RECT 313.950 194.850 316.050 195.750 ;
        RECT 320.400 193.050 321.450 196.950 ;
        RECT 322.950 193.950 325.050 196.050 ;
        RECT 310.950 190.950 313.050 193.050 ;
        RECT 319.950 190.950 322.050 193.050 ;
        RECT 313.950 187.950 316.050 190.050 ;
        RECT 307.950 169.950 310.050 172.050 ;
        RECT 314.400 169.050 315.450 187.950 ;
        RECT 319.950 184.950 322.050 187.050 ;
        RECT 320.400 169.050 321.450 184.950 ;
        RECT 307.950 168.450 310.050 169.050 ;
        RECT 305.400 167.400 310.050 168.450 ;
        RECT 292.950 164.250 294.750 165.150 ;
        RECT 295.950 163.950 298.050 166.050 ;
        RECT 299.250 164.250 301.050 165.150 ;
        RECT 292.950 160.950 295.050 163.050 ;
        RECT 296.250 161.850 297.750 162.750 ;
        RECT 298.950 160.950 301.050 163.050 ;
        RECT 268.950 157.950 271.050 160.050 ;
        RECT 274.950 157.950 277.050 160.050 ;
        RECT 280.950 158.850 283.050 159.750 ;
        RECT 289.950 157.950 292.050 160.050 ;
        RECT 271.950 154.950 274.050 157.050 ;
        RECT 268.950 145.950 271.050 148.050 ;
        RECT 241.950 139.950 244.050 142.050 ;
        RECT 247.950 139.950 250.050 142.050 ;
        RECT 265.950 139.950 268.050 142.050 ;
        RECT 241.950 136.950 244.050 139.050 ;
        RECT 227.400 131.400 231.450 132.450 ;
        RECT 232.950 132.450 235.050 133.050 ;
        RECT 235.950 132.450 238.050 133.050 ;
        RECT 232.950 131.400 238.050 132.450 ;
        RECT 227.400 130.050 228.450 131.400 ;
        RECT 232.950 130.950 235.050 131.400 ;
        RECT 235.950 130.950 238.050 131.400 ;
        RECT 238.950 130.950 241.050 133.050 ;
        RECT 224.250 128.250 225.750 129.150 ;
        RECT 226.950 127.950 229.050 130.050 ;
        RECT 229.950 127.950 232.050 130.050 ;
        RECT 233.250 128.250 234.750 129.150 ;
        RECT 238.950 127.950 241.050 130.050 ;
        RECT 220.950 125.850 222.750 126.750 ;
        RECT 223.950 124.950 226.050 127.050 ;
        RECT 227.250 125.850 229.050 126.750 ;
        RECT 229.950 125.850 231.750 126.750 ;
        RECT 232.950 124.950 235.050 127.050 ;
        RECT 236.250 125.850 238.050 126.750 ;
        RECT 224.400 118.050 225.450 124.950 ;
        RECT 239.400 124.050 240.450 127.950 ;
        RECT 232.950 121.950 235.050 124.050 ;
        RECT 238.950 121.950 241.050 124.050 ;
        RECT 223.950 115.950 226.050 118.050 ;
        RECT 214.950 109.950 217.050 112.050 ;
        RECT 220.950 109.950 223.050 112.050 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 215.400 97.050 216.450 100.950 ;
        RECT 221.400 97.050 222.450 109.950 ;
        RECT 223.950 103.950 226.050 106.050 ;
        RECT 169.950 94.950 172.050 97.050 ;
        RECT 173.250 95.250 175.050 96.150 ;
        RECT 175.950 95.250 178.050 96.150 ;
        RECT 178.950 95.850 181.050 96.750 ;
        RECT 181.950 95.250 183.750 96.150 ;
        RECT 184.950 94.950 187.050 97.050 ;
        RECT 193.950 95.250 196.050 96.150 ;
        RECT 196.950 95.850 199.050 96.750 ;
        RECT 199.950 94.950 202.050 97.050 ;
        RECT 203.250 95.250 204.750 96.150 ;
        RECT 205.950 94.950 208.050 97.050 ;
        RECT 211.950 94.950 214.050 97.050 ;
        RECT 214.950 94.950 217.050 97.050 ;
        RECT 218.250 95.250 219.750 96.150 ;
        RECT 220.950 94.950 223.050 97.050 ;
        RECT 224.400 94.050 225.450 103.950 ;
        RECT 229.950 100.950 232.050 103.050 ;
        RECT 151.950 91.950 154.050 94.050 ;
        RECT 154.950 91.950 157.050 94.050 ;
        RECT 158.250 92.850 159.750 93.750 ;
        RECT 160.950 91.950 163.050 94.050 ;
        RECT 164.250 92.850 166.050 93.750 ;
        RECT 166.950 91.950 169.050 94.050 ;
        RECT 169.950 92.850 171.750 93.750 ;
        RECT 172.950 91.950 175.050 94.050 ;
        RECT 175.950 91.950 178.050 94.050 ;
        RECT 181.950 91.950 184.050 94.050 ;
        RECT 185.250 92.850 187.050 93.750 ;
        RECT 187.950 91.950 190.050 94.050 ;
        RECT 193.950 91.950 196.050 94.050 ;
        RECT 199.950 92.850 201.750 93.750 ;
        RECT 202.950 91.950 205.050 94.050 ;
        RECT 206.250 92.850 207.750 93.750 ;
        RECT 208.950 93.450 211.050 94.050 ;
        RECT 208.950 92.400 213.450 93.450 ;
        RECT 214.950 92.850 216.750 93.750 ;
        RECT 208.950 91.950 211.050 92.400 ;
        RECT 152.400 87.450 153.450 91.950 ;
        RECT 161.400 91.050 162.450 91.950 ;
        RECT 154.950 89.850 157.050 90.750 ;
        RECT 160.950 88.950 163.050 91.050 ;
        RECT 152.400 86.400 156.450 87.450 ;
        RECT 148.950 61.950 151.050 64.050 ;
        RECT 139.950 58.950 142.050 61.050 ;
        RECT 140.400 58.050 141.450 58.950 ;
        RECT 149.400 58.050 150.450 61.950 ;
        RECT 155.400 58.050 156.450 86.400 ;
        RECT 173.400 82.050 174.450 91.950 ;
        RECT 166.950 79.950 169.050 82.050 ;
        RECT 172.950 79.950 175.050 82.050 ;
        RECT 167.400 58.050 168.450 79.950 ;
        RECT 181.950 73.950 184.050 76.050 ;
        RECT 169.950 61.950 172.050 64.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 128.250 56.250 129.750 57.150 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 133.950 55.950 136.050 58.050 ;
        RECT 137.250 56.250 138.750 57.150 ;
        RECT 139.950 55.950 142.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 154.950 57.450 157.050 58.050 ;
        RECT 152.250 56.250 153.750 57.150 ;
        RECT 154.950 56.400 159.450 57.450 ;
        RECT 154.950 55.950 157.050 56.400 ;
        RECT 112.950 53.250 115.050 54.150 ;
        RECT 115.950 52.950 118.050 55.050 ;
        RECT 118.950 53.250 121.050 54.150 ;
        RECT 124.950 53.850 126.750 54.750 ;
        RECT 127.950 52.950 130.050 55.050 ;
        RECT 131.250 53.850 133.050 54.750 ;
        RECT 133.950 53.850 135.750 54.750 ;
        RECT 136.950 52.950 139.050 55.050 ;
        RECT 140.250 53.850 142.050 54.750 ;
        RECT 142.950 52.950 145.050 55.050 ;
        RECT 148.950 53.850 150.750 54.750 ;
        RECT 151.950 52.950 154.050 55.050 ;
        RECT 155.250 53.850 157.050 54.750 ;
        RECT 112.950 49.950 115.050 52.050 ;
        RECT 116.250 50.250 117.750 51.150 ;
        RECT 118.950 49.950 121.050 52.050 ;
        RECT 113.400 46.050 114.450 49.950 ;
        RECT 119.400 49.050 120.450 49.950 ;
        RECT 115.950 46.950 118.050 49.050 ;
        RECT 118.950 46.950 121.050 49.050 ;
        RECT 112.950 43.950 115.050 46.050 ;
        RECT 109.950 34.950 112.050 37.050 ;
        RECT 116.400 30.450 117.450 46.950 ;
        RECT 121.950 43.950 124.050 46.050 ;
        RECT 122.400 34.050 123.450 43.950 ;
        RECT 128.400 34.050 129.450 52.950 ;
        RECT 137.400 49.050 138.450 52.950 ;
        RECT 136.950 46.950 139.050 49.050 ;
        RECT 137.400 40.050 138.450 46.950 ;
        RECT 143.400 43.050 144.450 52.950 ;
        RECT 158.400 49.050 159.450 56.400 ;
        RECT 164.250 56.250 165.750 57.150 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 170.400 55.050 171.450 61.950 ;
        RECT 175.950 58.950 178.050 61.050 ;
        RECT 176.400 55.050 177.450 58.950 ;
        RECT 182.400 55.050 183.450 73.950 ;
        RECT 188.400 58.050 189.450 91.950 ;
        RECT 203.400 79.050 204.450 91.950 ;
        RECT 205.950 88.950 208.050 91.050 ;
        RECT 208.950 89.850 211.050 90.750 ;
        RECT 202.950 76.950 205.050 79.050 ;
        RECT 202.950 64.950 205.050 67.050 ;
        RECT 203.400 64.050 204.450 64.950 ;
        RECT 206.400 64.050 207.450 88.950 ;
        RECT 212.400 88.050 213.450 92.400 ;
        RECT 217.950 91.950 220.050 94.050 ;
        RECT 221.250 92.850 222.750 93.750 ;
        RECT 223.950 91.950 226.050 94.050 ;
        RECT 218.400 91.050 219.450 91.950 ;
        RECT 217.950 88.950 220.050 91.050 ;
        RECT 223.950 89.850 226.050 90.750 ;
        RECT 211.950 85.950 214.050 88.050 ;
        RECT 223.950 79.950 226.050 82.050 ;
        RECT 224.400 78.450 225.450 79.950 ;
        RECT 230.400 79.050 231.450 100.950 ;
        RECT 233.400 97.050 234.450 121.950 ;
        RECT 242.400 115.050 243.450 136.950 ;
        RECT 248.400 136.050 249.450 139.950 ;
        RECT 247.950 133.950 250.050 136.050 ;
        RECT 259.950 130.950 262.050 133.050 ;
        RECT 244.950 128.250 247.050 129.150 ;
        RECT 244.950 124.950 247.050 127.050 ;
        RECT 248.250 125.250 249.750 126.150 ;
        RECT 250.950 124.950 253.050 127.050 ;
        RECT 254.250 125.250 256.050 126.150 ;
        RECT 256.950 125.250 259.050 126.150 ;
        RECT 245.400 124.050 246.450 124.950 ;
        RECT 244.950 121.950 247.050 124.050 ;
        RECT 247.950 121.950 250.050 124.050 ;
        RECT 251.250 122.850 252.750 123.750 ;
        RECT 253.950 121.950 256.050 124.050 ;
        RECT 256.950 121.950 259.050 124.050 ;
        RECT 241.950 112.950 244.050 115.050 ;
        RECT 248.400 106.050 249.450 121.950 ;
        RECT 254.400 109.050 255.450 121.950 ;
        RECT 257.400 121.050 258.450 121.950 ;
        RECT 256.950 118.950 259.050 121.050 ;
        RECT 256.950 115.950 259.050 118.050 ;
        RECT 253.950 106.950 256.050 109.050 ;
        RECT 247.950 103.950 250.050 106.050 ;
        RECT 257.400 105.450 258.450 115.950 ;
        RECT 260.400 115.050 261.450 130.950 ;
        RECT 262.950 125.850 265.050 126.750 ;
        RECT 265.950 125.250 268.050 126.150 ;
        RECT 262.950 121.950 265.050 124.050 ;
        RECT 265.950 121.950 268.050 124.050 ;
        RECT 259.950 112.950 262.050 115.050 ;
        RECT 263.400 112.050 264.450 121.950 ;
        RECT 269.400 121.050 270.450 145.950 ;
        RECT 272.400 145.050 273.450 154.950 ;
        RECT 271.950 142.950 274.050 145.050 ;
        RECT 272.400 124.050 273.450 142.950 ;
        RECT 275.400 139.050 276.450 157.950 ;
        RECT 293.400 157.050 294.450 160.950 ;
        RECT 299.400 159.450 300.450 160.950 ;
        RECT 305.400 160.050 306.450 167.400 ;
        RECT 307.950 166.950 310.050 167.400 ;
        RECT 311.250 167.250 312.750 168.150 ;
        RECT 313.950 166.950 316.050 169.050 ;
        RECT 317.250 167.250 318.750 168.150 ;
        RECT 319.950 166.950 322.050 169.050 ;
        RECT 323.400 166.050 324.450 193.950 ;
        RECT 332.400 187.050 333.450 200.400 ;
        RECT 334.950 199.950 337.050 200.400 ;
        RECT 338.250 200.250 339.750 201.150 ;
        RECT 340.950 199.950 343.050 202.050 ;
        RECT 352.950 199.950 355.050 202.050 ;
        RECT 356.400 199.050 357.450 229.950 ;
        RECT 365.400 204.450 366.450 241.950 ;
        RECT 368.400 228.600 369.600 245.400 ;
        RECT 367.950 226.500 370.050 228.600 ;
        RECT 362.400 203.400 366.450 204.450 ;
        RECT 334.950 197.850 336.750 198.750 ;
        RECT 337.950 196.950 340.050 199.050 ;
        RECT 341.250 197.850 343.050 198.750 ;
        RECT 349.950 197.250 352.050 198.150 ;
        RECT 355.950 196.950 358.050 199.050 ;
        RECT 338.400 196.050 339.450 196.950 ;
        RECT 337.950 193.950 340.050 196.050 ;
        RECT 346.950 194.250 348.750 195.150 ;
        RECT 349.950 193.950 352.050 196.050 ;
        RECT 355.950 194.850 358.050 195.750 ;
        RECT 346.950 192.450 349.050 193.050 ;
        RECT 344.400 191.400 349.050 192.450 ;
        RECT 331.950 184.950 334.050 187.050 ;
        RECT 331.950 169.950 334.050 172.050 ;
        RECT 332.400 169.050 333.450 169.950 ;
        RECT 331.950 166.950 334.050 169.050 ;
        RECT 307.950 164.850 309.750 165.750 ;
        RECT 310.950 163.950 313.050 166.050 ;
        RECT 314.250 164.850 315.750 165.750 ;
        RECT 316.950 163.950 319.050 166.050 ;
        RECT 320.250 164.850 322.050 165.750 ;
        RECT 322.950 163.950 325.050 166.050 ;
        RECT 325.950 164.250 327.750 165.150 ;
        RECT 328.950 163.950 331.050 166.050 ;
        RECT 311.400 163.050 312.450 163.950 ;
        RECT 332.400 163.050 333.450 166.950 ;
        RECT 344.400 166.050 345.450 191.400 ;
        RECT 346.950 190.950 349.050 191.400 ;
        RECT 352.950 169.950 355.050 172.050 ;
        RECT 349.950 167.250 352.050 168.150 ;
        RECT 352.950 167.850 355.050 168.750 ;
        RECT 355.950 167.250 357.750 168.150 ;
        RECT 358.950 166.950 361.050 169.050 ;
        RECT 334.950 165.450 337.050 166.050 ;
        RECT 334.950 164.400 339.450 165.450 ;
        RECT 334.950 163.950 337.050 164.400 ;
        RECT 310.950 160.950 313.050 163.050 ;
        RECT 325.950 160.950 328.050 163.050 ;
        RECT 329.250 161.850 330.750 162.750 ;
        RECT 331.950 160.950 334.050 163.050 ;
        RECT 335.250 161.850 337.050 162.750 ;
        RECT 338.400 160.050 339.450 164.400 ;
        RECT 340.950 164.250 342.750 165.150 ;
        RECT 343.950 163.950 346.050 166.050 ;
        RECT 347.250 164.250 349.050 165.150 ;
        RECT 349.950 163.950 352.050 166.050 ;
        RECT 355.950 163.950 358.050 166.050 ;
        RECT 359.250 164.850 361.050 165.750 ;
        RECT 340.950 160.950 343.050 163.050 ;
        RECT 344.250 161.850 345.750 162.750 ;
        RECT 346.950 162.450 349.050 163.050 ;
        RECT 350.400 162.450 351.450 163.950 ;
        RECT 346.950 161.400 351.450 162.450 ;
        RECT 346.950 160.950 349.050 161.400 ;
        RECT 347.400 160.050 348.450 160.950 ;
        RECT 296.400 158.400 300.450 159.450 ;
        RECT 292.950 154.950 295.050 157.050 ;
        RECT 274.950 136.950 277.050 139.050 ;
        RECT 289.950 133.950 292.050 136.050 ;
        RECT 290.400 133.050 291.450 133.950 ;
        RECT 274.950 130.950 277.050 133.050 ;
        RECT 289.950 130.950 292.050 133.050 ;
        RECT 275.400 127.050 276.450 130.950 ;
        RECT 290.400 130.050 291.450 130.950 ;
        RECT 296.400 130.050 297.450 158.400 ;
        RECT 304.950 157.950 307.050 160.050 ;
        RECT 331.950 158.850 334.050 159.750 ;
        RECT 337.950 157.950 340.050 160.050 ;
        RECT 340.950 157.950 343.050 160.050 ;
        RECT 346.950 157.950 349.050 160.050 ;
        RECT 298.950 130.950 301.050 133.050 ;
        RECT 287.250 128.250 288.750 129.150 ;
        RECT 289.950 127.950 292.050 130.050 ;
        RECT 295.950 127.950 298.050 130.050 ;
        RECT 296.400 127.050 297.450 127.950 ;
        RECT 274.950 124.950 277.050 127.050 ;
        RECT 283.950 125.850 285.750 126.750 ;
        RECT 286.950 124.950 289.050 127.050 ;
        RECT 290.250 125.850 292.050 126.750 ;
        RECT 295.950 124.950 298.050 127.050 ;
        RECT 271.950 121.950 274.050 124.050 ;
        RECT 274.950 122.850 277.050 123.750 ;
        RECT 277.950 122.250 280.050 123.150 ;
        RECT 287.400 121.050 288.450 124.950 ;
        RECT 292.950 122.250 295.050 123.150 ;
        RECT 295.950 122.850 298.050 123.750 ;
        RECT 268.950 118.950 271.050 121.050 ;
        RECT 277.950 118.950 280.050 121.050 ;
        RECT 286.950 118.950 289.050 121.050 ;
        RECT 292.950 118.950 295.050 121.050 ;
        RECT 278.400 118.050 279.450 118.950 ;
        RECT 277.950 115.950 280.050 118.050 ;
        RECT 289.950 115.950 292.050 118.050 ;
        RECT 274.950 112.950 277.050 115.050 ;
        RECT 262.950 109.950 265.050 112.050 ;
        RECT 254.400 104.400 258.450 105.450 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 239.400 100.050 240.450 100.950 ;
        RECT 238.950 97.950 241.050 100.050 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 254.400 97.050 255.450 104.400 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 256.950 97.950 259.050 100.050 ;
        RECT 232.950 94.950 235.050 97.050 ;
        RECT 236.250 95.250 238.050 96.150 ;
        RECT 238.950 95.850 241.050 96.750 ;
        RECT 241.950 95.250 244.050 96.150 ;
        RECT 244.950 95.250 247.050 96.150 ;
        RECT 247.950 95.850 250.050 96.750 ;
        RECT 250.950 95.250 252.750 96.150 ;
        RECT 253.950 94.950 256.050 97.050 ;
        RECT 232.950 92.850 234.750 93.750 ;
        RECT 235.950 91.950 238.050 94.050 ;
        RECT 238.950 91.950 241.050 94.050 ;
        RECT 241.950 93.450 244.050 94.050 ;
        RECT 244.950 93.450 247.050 94.050 ;
        RECT 241.950 92.400 247.050 93.450 ;
        RECT 241.950 91.950 244.050 92.400 ;
        RECT 244.950 91.950 247.050 92.400 ;
        RECT 250.950 91.950 253.050 94.050 ;
        RECT 254.250 92.850 256.050 93.750 ;
        RECT 236.400 91.050 237.450 91.950 ;
        RECT 235.950 88.950 238.050 91.050 ;
        RECT 224.400 77.400 228.450 78.450 ;
        RECT 208.950 67.950 211.050 70.050 ;
        RECT 202.950 61.950 205.050 64.050 ;
        RECT 205.950 61.950 208.050 64.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 196.950 56.250 199.050 57.150 ;
        RECT 199.950 55.950 202.050 58.050 ;
        RECT 191.400 55.050 192.450 55.950 ;
        RECT 160.950 53.850 162.750 54.750 ;
        RECT 163.950 52.950 166.050 55.050 ;
        RECT 167.250 53.850 169.050 54.750 ;
        RECT 169.950 52.950 172.050 55.050 ;
        RECT 172.950 53.250 174.750 54.150 ;
        RECT 175.950 52.950 178.050 55.050 ;
        RECT 179.250 53.250 180.750 54.150 ;
        RECT 181.950 52.950 184.050 55.050 ;
        RECT 185.250 53.250 187.050 54.150 ;
        RECT 187.950 53.250 189.750 54.150 ;
        RECT 190.950 52.950 193.050 55.050 ;
        RECT 194.250 53.250 195.750 54.150 ;
        RECT 196.950 52.950 199.050 55.050 ;
        RECT 157.950 46.950 160.050 49.050 ;
        RECT 154.950 43.950 157.050 46.050 ;
        RECT 142.950 40.950 145.050 43.050 ;
        RECT 136.950 37.950 139.050 40.050 ;
        RECT 133.950 34.950 136.050 37.050 ;
        RECT 134.400 34.050 135.450 34.950 ;
        RECT 121.950 31.950 124.050 34.050 ;
        RECT 127.950 31.950 130.050 34.050 ;
        RECT 133.950 31.950 136.050 34.050 ;
        RECT 151.950 31.950 154.050 34.050 ;
        RECT 101.400 29.400 105.450 30.450 ;
        RECT 113.400 29.400 120.450 30.450 ;
        RECT 88.950 25.950 91.050 28.050 ;
        RECT 94.950 25.950 97.050 28.050 ;
        RECT 101.400 25.050 102.450 29.400 ;
        RECT 113.400 28.050 114.450 29.400 ;
        RECT 119.400 28.050 120.450 29.400 ;
        RECT 122.400 28.050 123.450 31.950 ;
        RECT 112.950 25.950 115.050 28.050 ;
        RECT 115.950 25.950 118.050 28.050 ;
        RECT 118.950 25.950 121.050 28.050 ;
        RECT 121.950 25.950 124.050 28.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 23.250 94.050 24.150 ;
        RECT 94.950 23.850 97.050 24.750 ;
        RECT 97.950 23.250 99.750 24.150 ;
        RECT 100.950 22.950 103.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 113.250 23.250 115.050 24.150 ;
        RECT 115.950 23.850 118.050 24.750 ;
        RECT 118.950 23.250 121.050 24.150 ;
        RECT 121.950 23.850 124.050 24.750 ;
        RECT 124.950 23.250 127.050 24.150 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 82.950 19.950 85.050 22.050 ;
        RECT 86.250 20.250 88.050 21.150 ;
        RECT 89.400 19.050 90.450 22.950 ;
        RECT 91.950 19.950 94.050 22.050 ;
        RECT 97.950 19.950 100.050 22.050 ;
        RECT 101.250 20.850 103.050 21.750 ;
        RECT 109.950 20.850 111.750 21.750 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 118.950 19.950 121.050 22.050 ;
        RECT 124.950 19.950 127.050 22.050 ;
        RECT 64.950 18.450 67.050 19.050 ;
        RECT 62.400 17.400 67.050 18.450 ;
        RECT 68.250 17.850 69.750 18.750 ;
        RECT 64.950 16.950 67.050 17.400 ;
        RECT 70.950 16.950 73.050 19.050 ;
        RECT 74.250 17.850 76.050 18.750 ;
        RECT 76.950 17.850 78.750 18.750 ;
        RECT 79.950 16.950 82.050 19.050 ;
        RECT 83.250 17.850 84.750 18.750 ;
        RECT 85.950 16.950 88.050 19.050 ;
        RECT 88.950 16.950 91.050 19.050 ;
        RECT 10.950 14.850 13.050 15.750 ;
        RECT 70.950 14.850 73.050 15.750 ;
        RECT 79.950 14.850 82.050 15.750 ;
        RECT 86.400 15.450 87.450 16.950 ;
        RECT 92.400 16.050 93.450 19.950 ;
        RECT 98.400 19.050 99.450 19.950 ;
        RECT 97.950 16.950 100.050 19.050 ;
        RECT 125.400 16.050 126.450 19.950 ;
        RECT 131.400 19.050 132.450 22.950 ;
        RECT 134.400 22.050 135.450 31.950 ;
        RECT 142.950 28.950 145.050 31.050 ;
        RECT 143.400 25.050 144.450 28.950 ;
        RECT 152.400 28.050 153.450 31.950 ;
        RECT 155.400 31.050 156.450 43.950 ;
        RECT 164.400 34.050 165.450 52.950 ;
        RECT 172.950 49.950 175.050 52.050 ;
        RECT 176.250 50.850 177.750 51.750 ;
        RECT 178.950 49.950 181.050 52.050 ;
        RECT 182.250 50.850 183.750 51.750 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 187.950 49.950 190.050 52.050 ;
        RECT 191.250 50.850 192.750 51.750 ;
        RECT 193.950 49.950 196.050 52.050 ;
        RECT 166.950 46.950 169.050 49.050 ;
        RECT 175.950 46.950 178.050 49.050 ;
        RECT 167.400 34.050 168.450 46.950 ;
        RECT 169.950 43.950 172.050 46.050 ;
        RECT 163.950 31.950 166.050 34.050 ;
        RECT 166.950 31.950 169.050 34.050 ;
        RECT 154.950 28.950 157.050 31.050 ;
        RECT 160.950 28.950 163.050 31.050 ;
        RECT 145.950 25.950 148.050 28.050 ;
        RECT 151.950 25.950 154.050 28.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 140.250 23.250 141.750 24.150 ;
        RECT 142.950 22.950 145.050 25.050 ;
        RECT 146.400 22.050 147.450 25.950 ;
        RECT 155.400 25.050 156.450 28.950 ;
        RECT 161.400 25.050 162.450 28.950 ;
        RECT 164.400 25.050 165.450 31.950 ;
        RECT 170.400 25.050 171.450 43.950 ;
        RECT 176.400 25.050 177.450 46.950 ;
        RECT 179.400 43.050 180.450 49.950 ;
        RECT 188.400 46.050 189.450 49.950 ;
        RECT 187.950 43.950 190.050 46.050 ;
        RECT 178.950 40.950 181.050 43.050 ;
        RECT 190.950 34.950 193.050 37.050 ;
        RECT 181.950 28.950 184.050 31.050 ;
        RECT 148.950 23.250 151.050 24.150 ;
        RECT 151.950 23.850 154.050 24.750 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 158.250 23.250 159.750 24.150 ;
        RECT 160.950 22.950 163.050 25.050 ;
        RECT 163.950 22.950 166.050 25.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 173.250 23.250 174.750 24.150 ;
        RECT 175.950 22.950 178.050 25.050 ;
        RECT 164.400 22.050 165.450 22.950 ;
        RECT 133.950 19.950 136.050 22.050 ;
        RECT 137.250 20.850 138.750 21.750 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 143.250 20.850 145.050 21.750 ;
        RECT 145.950 19.950 148.050 22.050 ;
        RECT 148.950 19.950 151.050 22.050 ;
        RECT 154.950 20.850 156.750 21.750 ;
        RECT 157.950 19.950 160.050 22.050 ;
        RECT 161.250 20.850 162.750 21.750 ;
        RECT 163.950 19.950 166.050 22.050 ;
        RECT 166.950 19.950 169.050 22.050 ;
        RECT 169.950 20.850 171.750 21.750 ;
        RECT 172.950 19.950 175.050 22.050 ;
        RECT 176.250 20.850 177.750 21.750 ;
        RECT 178.950 19.950 181.050 22.050 ;
        RECT 149.400 19.050 150.450 19.950 ;
        RECT 130.950 16.950 133.050 19.050 ;
        RECT 133.950 17.850 136.050 18.750 ;
        RECT 148.950 16.950 151.050 19.050 ;
        RECT 163.950 17.850 166.050 18.750 ;
        RECT 167.400 18.450 168.450 19.950 ;
        RECT 173.400 18.450 174.450 19.950 ;
        RECT 167.400 17.400 174.450 18.450 ;
        RECT 178.950 17.850 181.050 18.750 ;
        RECT 88.950 15.450 91.050 16.050 ;
        RECT 86.400 14.400 91.050 15.450 ;
        RECT 88.950 13.950 91.050 14.400 ;
        RECT 91.950 13.950 94.050 16.050 ;
        RECT 124.950 13.950 127.050 16.050 ;
        RECT 182.400 10.050 183.450 28.950 ;
        RECT 191.400 22.050 192.450 34.950 ;
        RECT 194.400 31.050 195.450 49.950 ;
        RECT 200.400 43.050 201.450 55.950 ;
        RECT 203.400 55.050 204.450 61.950 ;
        RECT 209.400 55.050 210.450 67.950 ;
        RECT 217.950 58.950 220.050 61.050 ;
        RECT 218.400 55.050 219.450 58.950 ;
        RECT 223.950 56.250 226.050 57.150 ;
        RECT 202.950 52.950 205.050 55.050 ;
        RECT 205.950 53.250 208.050 54.150 ;
        RECT 208.950 52.950 211.050 55.050 ;
        RECT 211.950 53.250 214.050 54.150 ;
        RECT 214.950 53.250 216.750 54.150 ;
        RECT 217.950 52.950 220.050 55.050 ;
        RECT 221.250 53.250 222.750 54.150 ;
        RECT 223.950 52.950 226.050 55.050 ;
        RECT 205.950 49.950 208.050 52.050 ;
        RECT 209.250 50.250 210.750 51.150 ;
        RECT 211.950 49.950 214.050 52.050 ;
        RECT 214.950 49.950 217.050 52.050 ;
        RECT 218.250 50.850 219.750 51.750 ;
        RECT 220.950 49.950 223.050 52.050 ;
        RECT 199.950 40.950 202.050 43.050 ;
        RECT 206.400 40.050 207.450 49.950 ;
        RECT 208.950 46.950 211.050 49.050 ;
        RECT 211.950 46.950 214.050 49.050 ;
        RECT 209.400 40.050 210.450 46.950 ;
        RECT 205.950 37.950 208.050 40.050 ;
        RECT 208.950 37.950 211.050 40.050 ;
        RECT 212.400 37.050 213.450 46.950 ;
        RECT 215.400 43.050 216.450 49.950 ;
        RECT 217.950 46.950 220.050 49.050 ;
        RECT 220.950 46.950 223.050 49.050 ;
        RECT 214.950 40.950 217.050 43.050 ;
        RECT 205.950 34.950 208.050 37.050 ;
        RECT 211.950 34.950 214.050 37.050 ;
        RECT 193.950 28.950 196.050 31.050 ;
        RECT 199.950 22.950 202.050 25.050 ;
        RECT 200.400 22.050 201.450 22.950 ;
        RECT 206.400 22.050 207.450 34.950 ;
        RECT 214.950 25.950 217.050 28.050 ;
        RECT 215.400 25.050 216.450 25.950 ;
        RECT 218.400 25.050 219.450 46.950 ;
        RECT 221.400 40.050 222.450 46.950 ;
        RECT 224.400 46.050 225.450 52.950 ;
        RECT 223.950 43.950 226.050 46.050 ;
        RECT 220.950 37.950 223.050 40.050 ;
        RECT 227.400 28.050 228.450 77.400 ;
        RECT 229.950 76.950 232.050 79.050 ;
        RECT 232.950 76.950 235.050 79.050 ;
        RECT 230.400 55.050 231.450 76.950 ;
        RECT 233.400 58.050 234.450 76.950 ;
        RECT 236.400 58.050 237.450 88.950 ;
        RECT 239.400 79.050 240.450 91.950 ;
        RECT 245.400 79.050 246.450 91.950 ;
        RECT 251.400 90.450 252.450 91.950 ;
        RECT 257.400 91.050 258.450 97.950 ;
        RECT 260.400 94.050 261.450 100.950 ;
        RECT 265.950 97.950 268.050 100.050 ;
        RECT 271.950 97.950 274.050 100.050 ;
        RECT 266.400 94.050 267.450 97.950 ;
        RECT 259.950 93.450 262.050 94.050 ;
        RECT 262.950 93.450 265.050 94.050 ;
        RECT 259.950 92.400 265.050 93.450 ;
        RECT 259.950 91.950 262.050 92.400 ;
        RECT 262.950 91.950 265.050 92.400 ;
        RECT 265.950 91.950 268.050 94.050 ;
        RECT 269.250 92.250 271.050 93.150 ;
        RECT 251.400 89.400 255.450 90.450 ;
        RECT 250.950 85.950 253.050 88.050 ;
        RECT 238.950 76.950 241.050 79.050 ;
        RECT 244.950 76.950 247.050 79.050 ;
        RECT 238.950 64.950 241.050 67.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 229.950 52.950 232.050 55.050 ;
        RECT 232.950 54.450 235.050 55.050 ;
        RECT 232.950 53.400 237.450 54.450 ;
        RECT 232.950 52.950 235.050 53.400 ;
        RECT 229.950 50.250 232.050 51.150 ;
        RECT 232.950 50.850 235.050 51.750 ;
        RECT 229.950 46.950 232.050 49.050 ;
        RECT 230.400 43.050 231.450 46.950 ;
        RECT 229.950 40.950 232.050 43.050 ;
        RECT 236.400 40.050 237.450 53.400 ;
        RECT 239.400 43.050 240.450 64.950 ;
        RECT 244.950 58.950 247.050 61.050 ;
        RECT 245.400 55.050 246.450 58.950 ;
        RECT 251.400 58.050 252.450 85.950 ;
        RECT 254.400 79.050 255.450 89.400 ;
        RECT 256.950 88.950 259.050 91.050 ;
        RECT 259.950 89.850 261.750 90.750 ;
        RECT 262.950 88.950 265.050 91.050 ;
        RECT 266.250 89.850 267.750 90.750 ;
        RECT 268.950 88.950 271.050 91.050 ;
        RECT 262.950 86.850 265.050 87.750 ;
        RECT 265.950 85.950 268.050 88.050 ;
        RECT 253.950 76.950 256.050 79.050 ;
        RECT 259.950 73.950 262.050 76.050 ;
        RECT 256.950 70.950 259.050 73.050 ;
        RECT 257.400 69.450 258.450 70.950 ;
        RECT 254.400 68.400 258.450 69.450 ;
        RECT 254.400 64.050 255.450 68.400 ;
        RECT 253.950 61.950 256.050 64.050 ;
        RECT 256.950 61.950 259.050 64.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 257.400 55.050 258.450 61.950 ;
        RECT 260.400 55.050 261.450 73.950 ;
        RECT 266.400 73.050 267.450 85.950 ;
        RECT 269.400 73.050 270.450 88.950 ;
        RECT 272.400 82.050 273.450 97.950 ;
        RECT 275.400 97.050 276.450 112.950 ;
        RECT 274.950 94.950 277.050 97.050 ;
        RECT 280.950 96.450 283.050 97.050 ;
        RECT 283.950 96.450 286.050 97.050 ;
        RECT 278.250 95.250 279.750 96.150 ;
        RECT 280.950 95.400 286.050 96.450 ;
        RECT 280.950 94.950 283.050 95.400 ;
        RECT 283.950 94.950 286.050 95.400 ;
        RECT 274.950 92.850 276.750 93.750 ;
        RECT 277.950 91.950 280.050 94.050 ;
        RECT 281.250 92.850 282.750 93.750 ;
        RECT 283.950 93.450 286.050 94.050 ;
        RECT 283.950 92.400 288.450 93.450 ;
        RECT 283.950 91.950 286.050 92.400 ;
        RECT 274.950 88.950 277.050 91.050 ;
        RECT 271.950 79.950 274.050 82.050 ;
        RECT 275.400 79.050 276.450 88.950 ;
        RECT 278.400 88.050 279.450 91.950 ;
        RECT 283.950 89.850 286.050 90.750 ;
        RECT 277.950 85.950 280.050 88.050 ;
        RECT 283.950 85.950 286.050 88.050 ;
        RECT 284.400 85.050 285.450 85.950 ;
        RECT 283.950 82.950 286.050 85.050 ;
        RECT 274.950 76.950 277.050 79.050 ;
        RECT 274.950 73.950 277.050 76.050 ;
        RECT 265.950 70.950 268.050 73.050 ;
        RECT 268.950 70.950 271.050 73.050 ;
        RECT 265.950 59.250 268.050 60.150 ;
        RECT 271.950 58.950 274.050 61.050 ;
        RECT 272.400 58.050 273.450 58.950 ;
        RECT 262.950 56.250 264.750 57.150 ;
        RECT 265.950 55.950 268.050 58.050 ;
        RECT 269.250 56.250 270.750 57.150 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 241.950 53.250 243.750 54.150 ;
        RECT 244.950 52.950 247.050 55.050 ;
        RECT 250.950 52.950 253.050 55.050 ;
        RECT 256.950 52.950 259.050 55.050 ;
        RECT 259.950 52.950 262.050 55.050 ;
        RECT 262.950 52.950 265.050 55.050 ;
        RECT 241.950 49.950 244.050 52.050 ;
        RECT 245.250 50.850 247.050 51.750 ;
        RECT 247.950 50.250 250.050 51.150 ;
        RECT 250.950 50.850 253.050 51.750 ;
        RECT 253.950 50.250 256.050 51.150 ;
        RECT 256.950 50.850 259.050 51.750 ;
        RECT 259.950 49.950 262.050 52.050 ;
        RECT 262.950 49.950 265.050 52.050 ;
        RECT 238.950 40.950 241.050 43.050 ;
        RECT 235.950 37.950 238.050 40.050 ;
        RECT 242.400 31.050 243.450 49.950 ;
        RECT 247.950 46.950 250.050 49.050 ;
        RECT 250.950 46.950 253.050 49.050 ;
        RECT 253.950 46.950 256.050 49.050 ;
        RECT 248.400 40.050 249.450 46.950 ;
        RECT 247.950 37.950 250.050 40.050 ;
        RECT 244.950 34.950 247.050 37.050 ;
        RECT 251.400 36.450 252.450 46.950 ;
        RECT 254.400 46.050 255.450 46.950 ;
        RECT 253.950 43.950 256.050 46.050 ;
        RECT 260.400 42.450 261.450 49.950 ;
        RECT 263.400 46.050 264.450 49.950 ;
        RECT 262.950 43.950 265.050 46.050 ;
        RECT 260.400 41.400 264.450 42.450 ;
        RECT 248.400 35.400 252.450 36.450 ;
        RECT 229.950 28.950 232.050 31.050 ;
        RECT 241.950 28.950 244.050 31.050 ;
        RECT 223.950 25.950 226.050 28.050 ;
        RECT 226.950 25.950 229.050 28.050 ;
        RECT 214.950 22.950 217.050 25.050 ;
        RECT 217.950 22.950 220.050 25.050 ;
        RECT 221.250 23.250 223.050 24.150 ;
        RECT 223.950 23.850 226.050 24.750 ;
        RECT 226.950 23.250 229.050 24.150 ;
        RECT 215.400 22.050 216.450 22.950 ;
        RECT 230.400 22.050 231.450 28.950 ;
        RECT 232.950 22.950 235.050 25.050 ;
        RECT 184.950 19.950 187.050 22.050 ;
        RECT 190.950 19.950 193.050 22.050 ;
        RECT 194.250 20.250 196.050 21.150 ;
        RECT 199.950 19.950 202.050 22.050 ;
        RECT 205.950 19.950 208.050 22.050 ;
        RECT 209.250 20.250 211.050 21.150 ;
        RECT 214.950 19.950 217.050 22.050 ;
        RECT 217.950 20.850 219.750 21.750 ;
        RECT 220.950 19.950 223.050 22.050 ;
        RECT 226.950 19.950 229.050 22.050 ;
        RECT 229.950 19.950 232.050 22.050 ;
        RECT 227.400 19.050 228.450 19.950 ;
        RECT 233.400 19.050 234.450 22.950 ;
        RECT 242.400 22.050 243.450 28.950 ;
        RECT 235.950 19.950 238.050 22.050 ;
        RECT 239.250 20.250 241.050 21.150 ;
        RECT 241.950 19.950 244.050 22.050 ;
        RECT 245.400 19.050 246.450 34.950 ;
        RECT 248.400 25.050 249.450 35.400 ;
        RECT 253.950 34.950 256.050 37.050 ;
        RECT 254.400 30.450 255.450 34.950 ;
        RECT 251.400 29.400 255.450 30.450 ;
        RECT 251.400 28.050 252.450 29.400 ;
        RECT 250.950 25.950 253.050 28.050 ;
        RECT 253.950 25.950 256.050 28.050 ;
        RECT 259.950 25.950 262.050 28.050 ;
        RECT 247.950 22.950 250.050 25.050 ;
        RECT 251.250 23.250 253.050 24.150 ;
        RECT 253.950 23.850 256.050 24.750 ;
        RECT 256.950 23.250 259.050 24.150 ;
        RECT 260.400 22.050 261.450 25.950 ;
        RECT 263.400 25.050 264.450 41.400 ;
        RECT 266.400 40.050 267.450 55.950 ;
        RECT 268.950 52.950 271.050 55.050 ;
        RECT 272.250 53.850 274.050 54.750 ;
        RECT 269.400 43.050 270.450 52.950 ;
        RECT 275.400 52.050 276.450 73.950 ;
        RECT 287.400 70.050 288.450 92.400 ;
        RECT 280.950 67.950 283.050 70.050 ;
        RECT 286.950 67.950 289.050 70.050 ;
        RECT 277.950 64.950 280.050 67.050 ;
        RECT 278.400 55.050 279.450 64.950 ;
        RECT 281.400 55.050 282.450 67.950 ;
        RECT 286.950 64.950 289.050 67.050 ;
        RECT 283.950 61.950 286.050 64.050 ;
        RECT 284.400 55.050 285.450 61.950 ;
        RECT 287.400 61.050 288.450 64.950 ;
        RECT 286.950 58.950 289.050 61.050 ;
        RECT 290.400 60.450 291.450 115.950 ;
        RECT 293.400 109.050 294.450 118.950 ;
        RECT 299.400 118.050 300.450 130.950 ;
        RECT 305.400 130.050 306.450 157.950 ;
        RECT 322.950 139.950 325.050 142.050 ;
        RECT 310.950 131.250 313.050 132.150 ;
        RECT 304.950 127.950 307.050 130.050 ;
        RECT 308.250 128.250 309.750 129.150 ;
        RECT 310.950 127.950 313.050 130.050 ;
        RECT 314.250 128.250 316.050 129.150 ;
        RECT 304.950 125.850 306.750 126.750 ;
        RECT 307.950 124.950 310.050 127.050 ;
        RECT 301.950 118.950 304.050 121.050 ;
        RECT 298.950 115.950 301.050 118.050 ;
        RECT 298.950 112.950 301.050 115.050 ;
        RECT 295.950 109.950 298.050 112.050 ;
        RECT 292.950 106.950 295.050 109.050 ;
        RECT 296.400 105.450 297.450 109.950 ;
        RECT 293.400 104.400 297.450 105.450 ;
        RECT 293.400 97.050 294.450 104.400 ;
        RECT 299.400 100.050 300.450 112.950 ;
        RECT 302.400 100.050 303.450 118.950 ;
        RECT 307.950 115.950 310.050 118.050 ;
        RECT 304.950 106.950 307.050 109.050 ;
        RECT 298.950 97.950 301.050 100.050 ;
        RECT 301.950 97.950 304.050 100.050 ;
        RECT 305.400 97.050 306.450 106.950 ;
        RECT 308.400 106.050 309.450 115.950 ;
        RECT 307.950 103.950 310.050 106.050 ;
        RECT 311.400 97.050 312.450 127.950 ;
        RECT 313.950 124.950 316.050 127.050 ;
        RECT 319.950 124.950 322.050 127.050 ;
        RECT 314.400 120.450 315.450 124.950 ;
        RECT 316.950 122.250 319.050 123.150 ;
        RECT 319.950 122.850 322.050 123.750 ;
        RECT 316.950 120.450 319.050 121.050 ;
        RECT 314.400 119.400 319.050 120.450 ;
        RECT 316.950 118.950 319.050 119.400 ;
        RECT 313.950 103.950 316.050 106.050 ;
        RECT 292.950 94.950 295.050 97.050 ;
        RECT 296.250 95.250 298.050 96.150 ;
        RECT 298.950 95.850 301.050 96.750 ;
        RECT 301.950 95.250 304.050 96.150 ;
        RECT 304.950 94.950 307.050 97.050 ;
        RECT 308.250 95.250 309.750 96.150 ;
        RECT 310.950 94.950 313.050 97.050 ;
        RECT 314.400 94.050 315.450 103.950 ;
        RECT 317.400 100.050 318.450 118.950 ;
        RECT 319.950 109.950 322.050 112.050 ;
        RECT 316.950 97.950 319.050 100.050 ;
        RECT 316.950 94.950 319.050 97.050 ;
        RECT 292.950 92.850 294.750 93.750 ;
        RECT 295.950 91.950 298.050 94.050 ;
        RECT 298.950 91.950 301.050 94.050 ;
        RECT 301.950 91.950 304.050 94.050 ;
        RECT 304.950 92.850 306.750 93.750 ;
        RECT 307.950 91.950 310.050 94.050 ;
        RECT 311.250 92.850 312.750 93.750 ;
        RECT 313.950 91.950 316.050 94.050 ;
        RECT 296.400 91.050 297.450 91.950 ;
        RECT 295.950 88.950 298.050 91.050 ;
        RECT 299.400 73.050 300.450 91.950 ;
        RECT 302.400 84.450 303.450 91.950 ;
        RECT 302.400 83.400 306.450 84.450 ;
        RECT 305.400 82.050 306.450 83.400 ;
        RECT 301.950 79.950 304.050 82.050 ;
        RECT 304.950 79.950 307.050 82.050 ;
        RECT 298.950 70.950 301.050 73.050 ;
        RECT 292.950 60.450 295.050 61.050 ;
        RECT 290.400 59.400 295.050 60.450 ;
        RECT 292.950 58.950 295.050 59.400 ;
        RECT 293.400 58.050 294.450 58.950 ;
        RECT 302.400 58.050 303.450 79.950 ;
        RECT 308.400 79.050 309.450 91.950 ;
        RECT 317.400 91.050 318.450 94.950 ;
        RECT 313.950 89.850 316.050 90.750 ;
        RECT 316.950 88.950 319.050 91.050 ;
        RECT 316.950 85.950 319.050 88.050 ;
        RECT 307.950 76.950 310.050 79.050 ;
        RECT 317.400 64.050 318.450 85.950 ;
        RECT 320.400 79.050 321.450 109.950 ;
        RECT 323.400 103.050 324.450 139.950 ;
        RECT 334.950 128.250 337.050 129.150 ;
        RECT 325.950 125.250 327.750 126.150 ;
        RECT 328.950 124.950 331.050 127.050 ;
        RECT 332.250 125.250 333.750 126.150 ;
        RECT 334.950 124.950 337.050 127.050 ;
        RECT 325.950 121.950 328.050 124.050 ;
        RECT 329.250 122.850 330.750 123.750 ;
        RECT 331.950 121.950 334.050 124.050 ;
        RECT 335.400 121.050 336.450 124.950 ;
        RECT 341.400 124.050 342.450 157.950 ;
        RECT 362.400 133.050 363.450 203.400 ;
        RECT 371.400 202.050 372.450 250.950 ;
        RECT 380.400 241.050 381.450 265.950 ;
        RECT 383.400 253.050 384.450 272.400 ;
        RECT 394.950 272.250 397.050 273.150 ;
        RECT 385.950 269.250 387.750 270.150 ;
        RECT 388.950 268.950 391.050 271.050 ;
        RECT 392.250 269.250 393.750 270.150 ;
        RECT 394.950 268.950 397.050 271.050 ;
        RECT 385.950 265.950 388.050 268.050 ;
        RECT 389.250 266.850 390.750 267.750 ;
        RECT 391.950 267.450 394.050 268.050 ;
        RECT 398.400 267.450 399.450 295.950 ;
        RECT 400.950 292.950 403.050 295.050 ;
        RECT 391.950 266.400 399.450 267.450 ;
        RECT 401.400 273.450 402.450 292.950 ;
        RECT 410.400 277.050 411.450 304.950 ;
        RECT 412.950 298.950 415.050 301.050 ;
        RECT 409.950 274.950 412.050 277.050 ;
        RECT 403.950 273.450 406.050 274.050 ;
        RECT 401.400 272.400 406.050 273.450 ;
        RECT 391.950 265.950 394.050 266.400 ;
        RECT 386.400 265.050 387.450 265.950 ;
        RECT 385.950 262.950 388.050 265.050 ;
        RECT 382.950 250.950 385.050 253.050 ;
        RECT 382.950 247.950 385.050 250.050 ;
        RECT 383.400 241.050 384.450 247.950 ;
        RECT 401.400 247.050 402.450 272.400 ;
        RECT 403.950 271.950 406.050 272.400 ;
        RECT 407.250 272.250 408.750 273.150 ;
        RECT 409.950 271.950 412.050 274.050 ;
        RECT 403.950 269.850 405.750 270.750 ;
        RECT 406.950 268.950 409.050 271.050 ;
        RECT 410.250 269.850 412.050 270.750 ;
        RECT 403.950 267.450 406.050 268.050 ;
        RECT 407.400 267.450 408.450 268.950 ;
        RECT 403.950 266.400 408.450 267.450 ;
        RECT 403.950 265.950 406.050 266.400 ;
        RECT 413.400 247.050 414.450 298.950 ;
        RECT 422.400 292.050 423.450 373.950 ;
        RECT 430.950 350.400 433.050 352.500 ;
        RECT 424.950 341.250 427.050 342.150 ;
        RECT 427.950 340.950 430.050 343.050 ;
        RECT 424.950 339.450 427.050 340.050 ;
        RECT 428.400 339.450 429.450 340.950 ;
        RECT 424.950 338.400 429.450 339.450 ;
        RECT 424.950 337.950 427.050 338.400 ;
        RECT 431.400 333.600 432.600 350.400 ;
        RECT 430.950 331.500 433.050 333.600 ;
        RECT 434.400 328.050 435.450 385.950 ;
        RECT 437.400 385.050 438.450 415.950 ;
        RECT 440.400 405.600 441.600 422.400 ;
        RECT 439.950 403.500 442.050 405.600 ;
        RECT 436.950 382.950 439.050 385.050 ;
        RECT 443.400 384.450 444.450 424.950 ;
        RECT 445.950 413.250 448.050 414.150 ;
        RECT 445.950 409.950 448.050 412.050 ;
        RECT 449.400 397.050 450.450 427.950 ;
        RECT 451.950 413.250 454.050 414.150 ;
        RECT 451.950 409.950 454.050 412.050 ;
        RECT 452.400 409.050 453.450 409.950 ;
        RECT 451.950 406.950 454.050 409.050 ;
        RECT 455.400 403.050 456.450 448.950 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 454.950 400.950 457.050 403.050 ;
        RECT 448.950 394.950 451.050 397.050 ;
        RECT 449.400 385.050 450.450 394.950 ;
        RECT 454.950 385.950 457.050 388.050 ;
        RECT 455.400 385.050 456.450 385.950 ;
        RECT 443.400 383.400 447.450 384.450 ;
        RECT 436.950 380.250 438.750 381.150 ;
        RECT 439.950 379.950 442.050 382.050 ;
        RECT 443.250 380.250 445.050 381.150 ;
        RECT 436.950 376.950 439.050 379.050 ;
        RECT 440.250 377.850 441.750 378.750 ;
        RECT 442.950 376.950 445.050 379.050 ;
        RECT 443.400 376.050 444.450 376.950 ;
        RECT 442.950 373.950 445.050 376.050 ;
        RECT 446.400 364.050 447.450 383.400 ;
        RECT 448.950 382.950 451.050 385.050 ;
        RECT 454.950 382.950 457.050 385.050 ;
        RECT 448.950 380.850 451.050 381.750 ;
        RECT 454.950 380.850 457.050 381.750 ;
        RECT 436.950 361.950 439.050 364.050 ;
        RECT 445.950 361.950 448.050 364.050 ;
        RECT 433.950 325.950 436.050 328.050 ;
        RECT 437.400 325.050 438.450 361.950 ;
        RECT 458.400 348.450 459.450 445.950 ;
        RECT 464.400 442.050 465.450 457.950 ;
        RECT 467.400 457.050 468.450 460.950 ;
        RECT 473.400 460.050 474.450 460.950 ;
        RECT 472.950 457.950 475.050 460.050 ;
        RECT 479.400 457.050 480.450 481.950 ;
        RECT 488.400 469.050 489.450 484.950 ;
        RECT 491.400 481.050 492.450 491.400 ;
        RECT 496.950 488.250 499.050 489.150 ;
        RECT 512.400 487.050 513.450 520.950 ;
        RECT 518.400 492.450 519.450 547.950 ;
        RECT 521.400 535.050 522.450 557.400 ;
        RECT 523.950 557.250 526.050 558.150 ;
        RECT 523.950 555.450 526.050 556.050 ;
        RECT 527.400 555.450 528.450 562.950 ;
        RECT 529.950 559.950 532.050 562.050 ;
        RECT 535.950 559.950 538.050 562.050 ;
        RECT 529.950 557.850 532.050 558.750 ;
        RECT 532.950 557.250 535.050 558.150 ;
        RECT 523.950 554.400 528.450 555.450 ;
        RECT 523.950 553.950 526.050 554.400 ;
        RECT 532.950 553.950 535.050 556.050 ;
        RECT 536.400 555.450 537.450 559.950 ;
        RECT 542.400 559.050 543.450 562.950 ;
        RECT 547.950 560.250 550.050 561.150 ;
        RECT 538.950 557.250 540.750 558.150 ;
        RECT 541.950 556.950 544.050 559.050 ;
        RECT 547.950 558.450 550.050 559.050 ;
        RECT 551.400 558.450 552.450 574.950 ;
        RECT 562.950 560.250 565.050 561.150 ;
        RECT 545.250 557.250 546.750 558.150 ;
        RECT 547.950 557.400 552.450 558.450 ;
        RECT 547.950 556.950 550.050 557.400 ;
        RECT 553.950 557.250 555.750 558.150 ;
        RECT 556.950 556.950 559.050 559.050 ;
        RECT 560.250 557.250 561.750 558.150 ;
        RECT 562.950 556.950 565.050 559.050 ;
        RECT 538.950 555.450 541.050 556.050 ;
        RECT 536.400 554.400 541.050 555.450 ;
        RECT 542.250 554.850 543.750 555.750 ;
        RECT 544.950 555.450 547.050 556.050 ;
        RECT 553.950 555.450 556.050 556.050 ;
        RECT 538.950 553.950 541.050 554.400 ;
        RECT 544.950 554.400 556.050 555.450 ;
        RECT 557.250 554.850 558.750 555.750 ;
        RECT 544.950 553.950 547.050 554.400 ;
        RECT 553.950 553.950 556.050 554.400 ;
        RECT 559.950 553.950 562.050 556.050 ;
        RECT 539.400 541.050 540.450 553.950 ;
        RECT 544.950 544.950 547.050 547.050 ;
        RECT 523.950 538.950 526.050 541.050 ;
        RECT 538.950 538.950 541.050 541.050 ;
        RECT 520.950 532.950 523.050 535.050 ;
        RECT 520.950 529.950 523.050 532.050 ;
        RECT 521.400 502.050 522.450 529.950 ;
        RECT 524.400 529.050 525.450 538.950 ;
        RECT 529.950 532.950 532.050 535.050 ;
        RECT 535.950 532.950 538.050 535.050 ;
        RECT 526.950 529.950 529.050 532.050 ;
        RECT 530.400 529.050 531.450 532.950 ;
        RECT 536.400 532.050 537.450 532.950 ;
        RECT 535.950 529.950 538.050 532.050 ;
        RECT 523.950 526.950 526.050 529.050 ;
        RECT 527.250 527.850 528.750 528.750 ;
        RECT 529.950 526.950 532.050 529.050 ;
        RECT 532.950 527.250 535.050 528.150 ;
        RECT 535.950 527.850 538.050 528.750 ;
        RECT 538.950 527.250 540.750 528.150 ;
        RECT 541.950 526.950 544.050 529.050 ;
        RECT 523.950 524.850 526.050 525.750 ;
        RECT 529.950 524.850 532.050 525.750 ;
        RECT 532.950 523.950 535.050 526.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 542.250 524.850 544.050 525.750 ;
        RECT 523.950 520.950 526.050 523.050 ;
        RECT 520.950 499.950 523.050 502.050 ;
        RECT 520.950 496.950 523.050 499.050 ;
        RECT 515.400 491.400 519.450 492.450 ;
        RECT 515.400 490.050 516.450 491.400 ;
        RECT 514.950 487.950 517.050 490.050 ;
        RECT 517.950 488.250 520.050 489.150 ;
        RECT 493.950 484.950 496.050 487.050 ;
        RECT 496.950 484.950 499.050 487.050 ;
        RECT 500.250 485.250 501.750 486.150 ;
        RECT 502.950 484.950 505.050 487.050 ;
        RECT 506.250 485.250 508.050 486.150 ;
        RECT 508.950 485.250 510.750 486.150 ;
        RECT 511.950 484.950 514.050 487.050 ;
        RECT 515.250 485.250 516.750 486.150 ;
        RECT 517.950 484.950 520.050 487.050 ;
        RECT 490.950 478.950 493.050 481.050 ;
        RECT 487.950 466.950 490.050 469.050 ;
        RECT 481.950 457.950 484.050 460.050 ;
        RECT 466.950 454.950 469.050 457.050 ;
        RECT 470.250 455.250 472.050 456.150 ;
        RECT 472.950 455.850 475.050 456.750 ;
        RECT 475.950 455.250 478.050 456.150 ;
        RECT 478.950 454.950 481.050 457.050 ;
        RECT 482.250 455.850 483.750 456.750 ;
        RECT 484.950 456.450 487.050 457.050 ;
        RECT 484.950 455.400 489.450 456.450 ;
        RECT 484.950 454.950 487.050 455.400 ;
        RECT 466.950 452.850 468.750 453.750 ;
        RECT 469.950 451.950 472.050 454.050 ;
        RECT 472.950 451.950 475.050 454.050 ;
        RECT 475.950 451.950 478.050 454.050 ;
        RECT 478.950 452.850 481.050 453.750 ;
        RECT 484.950 452.850 487.050 453.750 ;
        RECT 470.400 451.050 471.450 451.950 ;
        RECT 469.950 448.950 472.050 451.050 ;
        RECT 463.950 439.950 466.050 442.050 ;
        RECT 464.400 433.050 465.450 439.950 ;
        RECT 463.950 430.950 466.050 433.050 ;
        RECT 460.950 423.300 463.050 425.400 ;
        RECT 461.250 419.700 462.450 423.300 ;
        RECT 460.950 417.600 463.050 419.700 ;
        RECT 463.950 418.950 466.050 421.050 ;
        RECT 461.250 405.600 462.450 417.600 ;
        RECT 464.400 412.050 465.450 418.950 ;
        RECT 463.950 409.950 466.050 412.050 ;
        RECT 463.950 407.850 466.050 408.750 ;
        RECT 460.950 403.500 463.050 405.600 ;
        RECT 466.950 403.950 469.050 406.050 ;
        RECT 467.400 385.050 468.450 403.950 ;
        RECT 473.400 400.050 474.450 451.950 ;
        RECT 488.400 448.050 489.450 455.400 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 475.950 422.400 478.050 424.500 ;
        RECT 476.400 405.600 477.600 422.400 ;
        RECT 481.950 413.250 484.050 414.150 ;
        RECT 487.950 413.250 490.050 414.150 ;
        RECT 481.950 409.950 484.050 412.050 ;
        RECT 487.950 409.950 490.050 412.050 ;
        RECT 482.400 406.050 483.450 409.950 ;
        RECT 488.400 409.050 489.450 409.950 ;
        RECT 487.950 406.950 490.050 409.050 ;
        RECT 475.950 403.500 478.050 405.600 ;
        RECT 481.950 403.950 484.050 406.050 ;
        RECT 491.400 405.450 492.450 478.950 ;
        RECT 494.400 451.050 495.450 484.950 ;
        RECT 497.400 484.050 498.450 484.950 ;
        RECT 518.400 484.050 519.450 484.950 ;
        RECT 496.950 481.950 499.050 484.050 ;
        RECT 499.950 481.950 502.050 484.050 ;
        RECT 503.250 482.850 504.750 483.750 ;
        RECT 505.950 481.950 508.050 484.050 ;
        RECT 508.950 481.950 511.050 484.050 ;
        RECT 512.250 482.850 513.750 483.750 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 517.950 481.950 520.050 484.050 ;
        RECT 500.400 475.050 501.450 481.950 ;
        RECT 499.950 472.950 502.050 475.050 ;
        RECT 496.950 461.400 499.050 463.500 ;
        RECT 506.400 463.050 507.450 481.950 ;
        RECT 509.400 481.050 510.450 481.950 ;
        RECT 508.950 478.950 511.050 481.050 ;
        RECT 508.950 463.950 511.050 466.050 ;
        RECT 493.950 448.950 496.050 451.050 ;
        RECT 488.400 404.400 492.450 405.450 ;
        RECT 481.950 400.950 484.050 403.050 ;
        RECT 472.950 397.950 475.050 400.050 ;
        RECT 460.950 382.950 463.050 385.050 ;
        RECT 464.250 383.250 465.750 384.150 ;
        RECT 466.950 382.950 469.050 385.050 ;
        RECT 460.950 380.850 462.750 381.750 ;
        RECT 463.950 379.950 466.050 382.050 ;
        RECT 467.250 380.850 468.750 381.750 ;
        RECT 469.950 379.950 472.050 382.050 ;
        RECT 469.950 377.850 472.050 378.750 ;
        RECT 463.950 352.950 466.050 355.050 ;
        RECT 455.400 347.400 459.450 348.450 ;
        RECT 442.950 344.250 445.050 345.150 ;
        RECT 448.950 343.950 451.050 346.050 ;
        RECT 449.400 343.050 450.450 343.950 ;
        RECT 442.950 340.950 445.050 343.050 ;
        RECT 446.250 341.250 447.750 342.150 ;
        RECT 448.950 340.950 451.050 343.050 ;
        RECT 452.250 341.250 454.050 342.150 ;
        RECT 439.950 337.950 442.050 340.050 ;
        RECT 440.400 337.050 441.450 337.950 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 436.950 322.950 439.050 325.050 ;
        RECT 430.950 317.400 433.050 319.500 ;
        RECT 431.400 300.600 432.600 317.400 ;
        RECT 436.950 310.950 439.050 313.050 ;
        RECT 440.400 312.450 441.450 334.950 ;
        RECT 443.400 331.050 444.450 340.950 ;
        RECT 445.950 337.950 448.050 340.050 ;
        RECT 449.250 338.850 450.750 339.750 ;
        RECT 451.950 337.950 454.050 340.050 ;
        RECT 442.950 328.950 445.050 331.050 ;
        RECT 452.400 328.050 453.450 337.950 ;
        RECT 445.950 325.950 448.050 328.050 ;
        RECT 451.950 325.950 454.050 328.050 ;
        RECT 442.950 312.450 445.050 313.050 ;
        RECT 440.400 311.400 445.050 312.450 ;
        RECT 436.950 308.850 439.050 309.750 ;
        RECT 436.950 304.950 439.050 307.050 ;
        RECT 430.950 298.500 433.050 300.600 ;
        RECT 421.950 289.950 424.050 292.050 ;
        RECT 433.950 272.250 436.050 273.150 ;
        RECT 415.950 269.250 418.050 270.150 ;
        RECT 421.950 269.250 424.050 270.150 ;
        RECT 424.950 269.250 426.750 270.150 ;
        RECT 427.950 268.950 430.050 271.050 ;
        RECT 431.250 269.250 432.750 270.150 ;
        RECT 433.950 268.950 436.050 271.050 ;
        RECT 437.400 268.050 438.450 304.950 ;
        RECT 440.400 280.050 441.450 311.400 ;
        RECT 442.950 310.950 445.050 311.400 ;
        RECT 442.950 308.850 445.050 309.750 ;
        RECT 439.950 277.950 442.050 280.050 ;
        RECT 442.950 268.950 445.050 271.050 ;
        RECT 415.950 265.950 418.050 268.050 ;
        RECT 419.250 266.250 420.750 267.150 ;
        RECT 421.950 265.950 424.050 268.050 ;
        RECT 424.950 265.950 427.050 268.050 ;
        RECT 428.250 266.850 429.750 267.750 ;
        RECT 430.950 265.950 433.050 268.050 ;
        RECT 436.950 265.950 439.050 268.050 ;
        RECT 439.950 266.250 442.050 267.150 ;
        RECT 442.950 266.850 445.050 267.750 ;
        RECT 416.400 253.050 417.450 265.950 ;
        RECT 422.400 265.050 423.450 265.950 ;
        RECT 425.400 265.050 426.450 265.950 ;
        RECT 418.950 262.950 421.050 265.050 ;
        RECT 421.950 262.950 424.050 265.050 ;
        RECT 424.950 262.950 427.050 265.050 ;
        RECT 439.950 262.950 442.050 265.050 ;
        RECT 415.950 250.950 418.050 253.050 ;
        RECT 391.950 244.950 394.050 247.050 ;
        RECT 400.950 244.950 403.050 247.050 ;
        RECT 406.950 244.950 409.050 247.050 ;
        RECT 412.950 244.950 415.050 247.050 ;
        RECT 388.950 241.950 391.050 244.050 ;
        RECT 389.400 241.050 390.450 241.950 ;
        RECT 379.950 238.950 382.050 241.050 ;
        RECT 382.950 238.950 385.050 241.050 ;
        RECT 386.250 239.250 387.750 240.150 ;
        RECT 388.950 238.950 391.050 241.050 ;
        RECT 379.950 235.950 382.050 238.050 ;
        RECT 383.250 236.850 384.750 237.750 ;
        RECT 385.950 235.950 388.050 238.050 ;
        RECT 389.250 236.850 391.050 237.750 ;
        RECT 392.400 235.050 393.450 244.950 ;
        RECT 407.400 241.050 408.450 244.950 ;
        RECT 409.950 241.950 412.050 244.050 ;
        RECT 419.400 243.450 420.450 262.950 ;
        RECT 424.950 250.950 427.050 253.050 ;
        RECT 425.400 244.050 426.450 250.950 ;
        RECT 440.400 247.050 441.450 262.950 ;
        RECT 439.950 244.950 442.050 247.050 ;
        RECT 421.950 243.450 424.050 244.050 ;
        RECT 419.400 242.400 424.050 243.450 ;
        RECT 421.950 241.950 424.050 242.400 ;
        RECT 424.950 241.950 427.050 244.050 ;
        RECT 439.950 241.950 442.050 244.050 ;
        RECT 394.950 238.950 397.050 241.050 ;
        RECT 403.950 238.950 406.050 241.050 ;
        RECT 406.950 238.950 409.050 241.050 ;
        RECT 410.250 239.850 411.750 240.750 ;
        RECT 412.950 240.450 415.050 241.050 ;
        RECT 412.950 239.400 417.450 240.450 ;
        RECT 412.950 238.950 415.050 239.400 ;
        RECT 394.950 236.850 397.050 237.750 ;
        RECT 397.950 236.250 400.050 237.150 ;
        RECT 403.950 236.850 406.050 237.750 ;
        RECT 406.950 236.850 409.050 237.750 ;
        RECT 412.950 236.850 415.050 237.750 ;
        RECT 416.400 235.050 417.450 239.400 ;
        RECT 418.950 239.250 421.050 240.150 ;
        RECT 421.950 239.850 424.050 240.750 ;
        RECT 424.950 239.250 426.750 240.150 ;
        RECT 427.950 238.950 430.050 241.050 ;
        RECT 433.950 238.950 436.050 241.050 ;
        RECT 436.950 238.950 439.050 241.050 ;
        RECT 440.250 239.850 441.750 240.750 ;
        RECT 442.950 238.950 445.050 241.050 ;
        RECT 418.950 235.950 421.050 238.050 ;
        RECT 424.950 235.950 427.050 238.050 ;
        RECT 428.250 236.850 430.050 237.750 ;
        RECT 430.950 235.950 433.050 238.050 ;
        RECT 379.950 233.850 382.050 234.750 ;
        RECT 382.950 232.950 385.050 235.050 ;
        RECT 391.950 232.950 394.050 235.050 ;
        RECT 397.950 232.950 400.050 235.050 ;
        RECT 415.950 232.950 418.050 235.050 ;
        RECT 364.950 199.950 367.050 202.050 ;
        RECT 368.250 200.250 369.750 201.150 ;
        RECT 370.950 199.950 373.050 202.050 ;
        RECT 364.950 197.850 366.750 198.750 ;
        RECT 367.950 196.950 370.050 199.050 ;
        RECT 371.250 197.850 373.050 198.750 ;
        RECT 376.950 196.950 379.050 199.050 ;
        RECT 368.400 193.050 369.450 196.950 ;
        RECT 373.950 194.250 376.050 195.150 ;
        RECT 376.950 194.850 379.050 195.750 ;
        RECT 383.400 195.450 384.450 232.950 ;
        RECT 419.400 232.050 420.450 235.950 ;
        RECT 418.950 229.950 421.050 232.050 ;
        RECT 397.950 202.950 400.050 205.050 ;
        RECT 388.950 199.950 391.050 202.050 ;
        RECT 385.950 197.250 388.050 198.150 ;
        RECT 389.400 196.050 390.450 199.950 ;
        RECT 398.400 199.050 399.450 202.950 ;
        RECT 403.950 200.250 406.050 201.150 ;
        RECT 406.950 199.950 409.050 202.050 ;
        RECT 421.950 199.950 424.050 202.050 ;
        RECT 391.950 197.250 394.050 198.150 ;
        RECT 394.950 197.250 396.750 198.150 ;
        RECT 397.950 196.950 400.050 199.050 ;
        RECT 403.950 198.450 406.050 199.050 ;
        RECT 407.400 198.450 408.450 199.950 ;
        RECT 422.400 199.050 423.450 199.950 ;
        RECT 401.250 197.250 402.750 198.150 ;
        RECT 403.950 197.400 408.450 198.450 ;
        RECT 403.950 196.950 406.050 197.400 ;
        RECT 412.950 197.250 414.750 198.150 ;
        RECT 415.950 196.950 418.050 199.050 ;
        RECT 419.250 197.250 420.750 198.150 ;
        RECT 421.950 196.950 424.050 199.050 ;
        RECT 425.250 197.250 427.050 198.150 ;
        RECT 385.950 195.450 388.050 196.050 ;
        RECT 383.400 194.400 388.050 195.450 ;
        RECT 385.950 193.950 388.050 194.400 ;
        RECT 388.950 193.950 391.050 196.050 ;
        RECT 391.950 193.950 394.050 196.050 ;
        RECT 394.950 193.950 397.050 196.050 ;
        RECT 398.250 194.850 399.750 195.750 ;
        RECT 400.950 193.950 403.050 196.050 ;
        RECT 412.950 193.950 415.050 196.050 ;
        RECT 416.250 194.850 417.750 195.750 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 422.250 194.850 423.750 195.750 ;
        RECT 424.950 193.950 427.050 196.050 ;
        RECT 367.950 190.950 370.050 193.050 ;
        RECT 373.950 190.950 376.050 193.050 ;
        RECT 392.400 172.050 393.450 193.950 ;
        RECT 419.400 187.050 420.450 193.950 ;
        RECT 418.950 184.950 421.050 187.050 ;
        RECT 403.950 178.950 406.050 181.050 ;
        RECT 394.950 175.950 397.050 178.050 ;
        RECT 370.950 171.450 373.050 172.050 ;
        RECT 370.950 170.400 375.450 171.450 ;
        RECT 370.950 169.950 373.050 170.400 ;
        RECT 367.950 167.250 370.050 168.150 ;
        RECT 370.950 167.850 373.050 168.750 ;
        RECT 367.950 163.950 370.050 166.050 ;
        RECT 374.400 145.050 375.450 170.400 ;
        RECT 391.950 169.950 394.050 172.050 ;
        RECT 395.400 169.050 396.450 175.950 ;
        RECT 400.950 172.950 403.050 175.050 ;
        RECT 401.400 169.050 402.450 172.950 ;
        RECT 404.400 172.050 405.450 178.950 ;
        RECT 427.950 175.950 430.050 178.050 ;
        RECT 421.950 173.400 424.050 175.500 ;
        RECT 403.950 169.950 406.050 172.050 ;
        RECT 404.400 169.050 405.450 169.950 ;
        RECT 388.950 166.950 391.050 169.050 ;
        RECT 392.250 167.250 393.750 168.150 ;
        RECT 394.950 166.950 397.050 169.050 ;
        RECT 398.250 167.250 399.750 168.150 ;
        RECT 400.950 166.950 403.050 169.050 ;
        RECT 403.950 166.950 406.050 169.050 ;
        RECT 409.950 166.950 412.050 169.050 ;
        RECT 418.950 166.950 421.050 169.050 ;
        RECT 376.950 164.250 378.750 165.150 ;
        RECT 379.950 163.950 382.050 166.050 ;
        RECT 383.250 164.250 385.050 165.150 ;
        RECT 388.950 164.850 390.750 165.750 ;
        RECT 391.950 163.950 394.050 166.050 ;
        RECT 395.250 164.850 396.750 165.750 ;
        RECT 397.950 163.950 400.050 166.050 ;
        RECT 401.250 164.850 403.050 165.750 ;
        RECT 403.950 164.850 406.050 165.750 ;
        RECT 409.950 164.850 412.050 165.750 ;
        RECT 398.400 163.050 399.450 163.950 ;
        RECT 376.950 160.950 379.050 163.050 ;
        RECT 380.250 161.850 381.750 162.750 ;
        RECT 382.950 160.950 385.050 163.050 ;
        RECT 397.950 160.950 400.050 163.050 ;
        RECT 376.950 145.950 379.050 148.050 ;
        RECT 373.950 142.950 376.050 145.050 ;
        RECT 361.950 130.950 364.050 133.050 ;
        RECT 367.950 131.250 370.050 132.150 ;
        RECT 352.950 127.950 355.050 130.050 ;
        RECT 364.950 128.250 366.750 129.150 ;
        RECT 367.950 127.950 370.050 130.050 ;
        RECT 371.250 128.250 372.750 129.150 ;
        RECT 373.950 127.950 376.050 130.050 ;
        RECT 353.400 127.050 354.450 127.950 ;
        RECT 343.950 125.250 345.750 126.150 ;
        RECT 346.950 124.950 349.050 127.050 ;
        RECT 352.950 124.950 355.050 127.050 ;
        RECT 358.950 124.950 361.050 127.050 ;
        RECT 364.950 124.950 367.050 127.050 ;
        RECT 340.950 121.950 343.050 124.050 ;
        RECT 343.950 121.950 346.050 124.050 ;
        RECT 347.250 122.850 349.050 123.750 ;
        RECT 349.950 122.250 352.050 123.150 ;
        RECT 352.950 122.850 355.050 123.750 ;
        RECT 355.950 122.250 358.050 123.150 ;
        RECT 358.950 122.850 361.050 123.750 ;
        RECT 344.400 121.050 345.450 121.950 ;
        RECT 325.950 118.950 328.050 121.050 ;
        RECT 334.950 118.950 337.050 121.050 ;
        RECT 343.950 118.950 346.050 121.050 ;
        RECT 349.950 118.950 352.050 121.050 ;
        RECT 355.950 118.950 358.050 121.050 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 326.400 94.050 327.450 118.950 ;
        RECT 337.950 115.950 340.050 118.050 ;
        RECT 328.950 112.950 331.050 115.050 ;
        RECT 322.950 92.250 324.750 93.150 ;
        RECT 325.950 91.950 328.050 94.050 ;
        RECT 329.400 91.050 330.450 112.950 ;
        RECT 338.400 97.050 339.450 115.950 ;
        RECT 340.950 109.950 343.050 112.050 ;
        RECT 341.400 97.050 342.450 109.950 ;
        RECT 350.400 103.050 351.450 118.950 ;
        RECT 356.400 106.050 357.450 118.950 ;
        RECT 364.950 112.950 367.050 115.050 ;
        RECT 355.950 103.950 358.050 106.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 355.950 100.950 358.050 103.050 ;
        RECT 346.950 97.950 349.050 100.050 ;
        RECT 349.950 97.950 352.050 100.050 ;
        RECT 347.400 97.050 348.450 97.950 ;
        RECT 350.400 97.050 351.450 97.950 ;
        RECT 356.400 97.050 357.450 100.950 ;
        RECT 361.950 97.950 364.050 100.050 ;
        RECT 331.950 94.950 334.050 97.050 ;
        RECT 337.950 94.950 340.050 97.050 ;
        RECT 340.950 94.950 343.050 97.050 ;
        RECT 344.250 95.250 345.750 96.150 ;
        RECT 346.950 94.950 349.050 97.050 ;
        RECT 349.950 94.950 352.050 97.050 ;
        RECT 353.250 95.250 354.750 96.150 ;
        RECT 355.950 94.950 358.050 97.050 ;
        RECT 358.950 94.950 361.050 97.050 ;
        RECT 332.400 94.050 333.450 94.950 ;
        RECT 359.400 94.050 360.450 94.950 ;
        RECT 331.950 93.450 334.050 94.050 ;
        RECT 337.950 93.450 340.050 94.050 ;
        RECT 331.950 92.400 340.050 93.450 ;
        RECT 341.250 92.850 342.750 93.750 ;
        RECT 331.950 91.950 334.050 92.400 ;
        RECT 322.950 88.950 325.050 91.050 ;
        RECT 326.250 89.850 327.750 90.750 ;
        RECT 328.950 88.950 331.050 91.050 ;
        RECT 332.250 89.850 334.050 90.750 ;
        RECT 325.950 85.950 328.050 88.050 ;
        RECT 328.950 86.850 331.050 87.750 ;
        RECT 326.400 82.050 327.450 85.950 ;
        RECT 325.950 79.950 328.050 82.050 ;
        RECT 319.950 76.950 322.050 79.050 ;
        RECT 319.950 70.950 322.050 73.050 ;
        RECT 325.950 70.950 328.050 73.050 ;
        RECT 304.950 61.950 307.050 64.050 ;
        RECT 316.950 61.950 319.050 64.050 ;
        RECT 305.400 58.050 306.450 61.950 ;
        RECT 320.400 60.450 321.450 70.950 ;
        RECT 326.400 61.050 327.450 70.950 ;
        RECT 328.950 67.950 331.050 70.050 ;
        RECT 317.400 59.400 321.450 60.450 ;
        RECT 317.400 58.050 318.450 59.400 ;
        RECT 325.950 58.950 328.050 61.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 296.250 56.250 297.750 57.150 ;
        RECT 301.950 55.950 304.050 58.050 ;
        RECT 304.950 55.950 307.050 58.050 ;
        RECT 308.250 56.250 309.750 57.150 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 322.950 57.450 325.050 58.050 ;
        RECT 320.250 56.250 321.750 57.150 ;
        RECT 322.950 56.400 327.450 57.450 ;
        RECT 322.950 55.950 325.050 56.400 ;
        RECT 277.950 52.950 280.050 55.050 ;
        RECT 280.950 52.950 283.050 55.050 ;
        RECT 283.950 52.950 286.050 55.050 ;
        RECT 287.250 53.250 289.050 54.150 ;
        RECT 292.950 53.850 294.750 54.750 ;
        RECT 295.950 52.950 298.050 55.050 ;
        RECT 299.250 53.850 301.050 54.750 ;
        RECT 301.950 52.950 304.050 55.050 ;
        RECT 304.950 53.850 306.750 54.750 ;
        RECT 307.950 52.950 310.050 55.050 ;
        RECT 311.250 53.850 313.050 54.750 ;
        RECT 316.950 53.850 318.750 54.750 ;
        RECT 319.950 52.950 322.050 55.050 ;
        RECT 323.250 53.850 325.050 54.750 ;
        RECT 274.950 49.950 277.050 52.050 ;
        RECT 277.950 50.850 280.050 51.750 ;
        RECT 280.950 50.250 283.050 51.150 ;
        RECT 283.950 50.850 285.750 51.750 ;
        RECT 286.950 49.950 289.050 52.050 ;
        RECT 277.950 46.950 280.050 49.050 ;
        RECT 280.950 46.950 283.050 49.050 ;
        RECT 268.950 40.950 271.050 43.050 ;
        RECT 265.950 37.950 268.050 40.050 ;
        RECT 265.950 28.950 268.050 31.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 266.400 22.050 267.450 28.950 ;
        RECT 278.400 22.050 279.450 46.950 ;
        RECT 281.400 40.050 282.450 46.950 ;
        RECT 292.950 43.950 295.050 46.050 ;
        RECT 280.950 37.950 283.050 40.050 ;
        RECT 293.400 28.050 294.450 43.950 ;
        RECT 296.400 40.050 297.450 52.950 ;
        RECT 302.400 49.050 303.450 52.950 ;
        RECT 307.950 49.950 310.050 52.050 ;
        RECT 301.950 46.950 304.050 49.050 ;
        RECT 304.950 46.950 307.050 49.050 ;
        RECT 305.400 46.050 306.450 46.950 ;
        RECT 298.950 43.950 301.050 46.050 ;
        RECT 304.950 43.950 307.050 46.050 ;
        RECT 295.950 37.950 298.050 40.050 ;
        RECT 292.950 25.950 295.050 28.050 ;
        RECT 293.400 25.050 294.450 25.950 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 247.950 20.850 249.750 21.750 ;
        RECT 250.950 19.950 253.050 22.050 ;
        RECT 253.950 19.950 256.050 22.050 ;
        RECT 256.950 19.950 259.050 22.050 ;
        RECT 259.950 19.950 262.050 22.050 ;
        RECT 265.950 19.950 268.050 22.050 ;
        RECT 269.250 20.250 271.050 21.150 ;
        RECT 274.950 20.250 276.750 21.150 ;
        RECT 277.950 19.950 280.050 22.050 ;
        RECT 281.250 20.250 283.050 21.150 ;
        RECT 286.950 20.850 289.050 21.750 ;
        RECT 292.950 20.850 295.050 21.750 ;
        RECT 184.950 17.850 186.750 18.750 ;
        RECT 187.950 16.950 190.050 19.050 ;
        RECT 191.250 17.850 192.750 18.750 ;
        RECT 193.950 16.950 196.050 19.050 ;
        RECT 199.950 17.850 201.750 18.750 ;
        RECT 202.950 16.950 205.050 19.050 ;
        RECT 206.250 17.850 207.750 18.750 ;
        RECT 208.950 16.950 211.050 19.050 ;
        RECT 226.950 16.950 229.050 19.050 ;
        RECT 229.950 17.850 231.750 18.750 ;
        RECT 232.950 16.950 235.050 19.050 ;
        RECT 236.250 17.850 237.750 18.750 ;
        RECT 238.950 16.950 241.050 19.050 ;
        RECT 244.950 16.950 247.050 19.050 ;
        RECT 209.400 16.050 210.450 16.950 ;
        RECT 187.950 14.850 190.050 15.750 ;
        RECT 202.950 14.850 205.050 15.750 ;
        RECT 208.950 13.950 211.050 16.050 ;
        RECT 227.400 10.050 228.450 16.950 ;
        RECT 254.400 16.050 255.450 19.950 ;
        RECT 257.400 19.050 258.450 19.950 ;
        RECT 256.950 16.950 259.050 19.050 ;
        RECT 259.950 17.850 261.750 18.750 ;
        RECT 262.950 16.950 265.050 19.050 ;
        RECT 266.250 17.850 267.750 18.750 ;
        RECT 268.950 16.950 271.050 19.050 ;
        RECT 274.950 16.950 277.050 19.050 ;
        RECT 278.250 17.850 279.750 18.750 ;
        RECT 286.950 16.950 289.050 19.050 ;
        RECT 269.400 16.050 270.450 16.950 ;
        RECT 232.950 14.850 235.050 15.750 ;
        RECT 253.950 13.950 256.050 16.050 ;
        RECT 262.950 14.850 265.050 15.750 ;
        RECT 268.950 13.950 271.050 16.050 ;
        RECT 275.400 13.050 276.450 16.950 ;
        RECT 287.400 13.050 288.450 16.950 ;
        RECT 299.400 16.050 300.450 43.950 ;
        RECT 301.950 31.950 304.050 34.050 ;
        RECT 302.400 25.050 303.450 31.950 ;
        RECT 308.400 28.050 309.450 49.950 ;
        RECT 320.400 46.050 321.450 52.950 ;
        RECT 319.950 43.950 322.050 46.050 ;
        RECT 310.950 34.950 313.050 37.050 ;
        RECT 311.400 28.050 312.450 34.950 ;
        RECT 326.400 34.050 327.450 56.400 ;
        RECT 329.400 55.050 330.450 67.950 ;
        RECT 335.400 55.050 336.450 92.400 ;
        RECT 337.950 91.950 340.050 92.400 ;
        RECT 343.950 91.950 346.050 94.050 ;
        RECT 347.250 92.850 349.050 93.750 ;
        RECT 349.950 92.850 351.750 93.750 ;
        RECT 352.950 91.950 355.050 94.050 ;
        RECT 356.250 92.850 357.750 93.750 ;
        RECT 358.950 91.950 361.050 94.050 ;
        RECT 337.950 89.850 340.050 90.750 ;
        RECT 340.950 88.950 343.050 91.050 ;
        RECT 343.950 88.950 346.050 91.050 ;
        RECT 358.950 89.850 361.050 90.750 ;
        RECT 341.400 67.050 342.450 88.950 ;
        RECT 344.400 73.050 345.450 88.950 ;
        RECT 362.400 76.050 363.450 97.950 ;
        RECT 365.400 94.050 366.450 112.950 ;
        RECT 368.400 106.050 369.450 127.950 ;
        RECT 370.950 124.950 373.050 127.050 ;
        RECT 374.250 125.850 376.050 126.750 ;
        RECT 367.950 103.950 370.050 106.050 ;
        RECT 371.400 103.050 372.450 124.950 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 377.400 100.050 378.450 145.950 ;
        RECT 382.950 142.950 385.050 145.050 ;
        RECT 383.400 130.050 384.450 142.950 ;
        RECT 388.950 131.250 391.050 132.150 ;
        RECT 419.400 130.050 420.450 166.950 ;
        RECT 422.400 156.600 423.600 173.400 ;
        RECT 428.400 169.050 429.450 175.950 ;
        RECT 431.400 175.050 432.450 235.950 ;
        RECT 434.400 235.050 435.450 238.950 ;
        RECT 436.950 236.850 439.050 237.750 ;
        RECT 442.950 236.850 445.050 237.750 ;
        RECT 433.950 232.950 436.050 235.050 ;
        RECT 436.950 229.950 439.050 232.050 ;
        RECT 433.950 206.400 436.050 208.500 ;
        RECT 434.400 189.600 435.600 206.400 ;
        RECT 433.950 187.500 436.050 189.600 ;
        RECT 430.950 172.950 433.050 175.050 ;
        RECT 433.950 172.950 436.050 175.050 ;
        RECT 434.400 169.050 435.450 172.950 ;
        RECT 427.950 166.950 430.050 169.050 ;
        RECT 433.950 166.950 436.050 169.050 ;
        RECT 427.950 164.850 430.050 165.750 ;
        RECT 433.950 164.850 436.050 165.750 ;
        RECT 437.400 160.050 438.450 229.950 ;
        RECT 446.400 205.050 447.450 325.950 ;
        RECT 448.950 316.950 451.050 319.050 ;
        RECT 451.950 317.400 454.050 319.500 ;
        RECT 455.400 319.050 456.450 347.400 ;
        RECT 457.950 344.250 460.050 345.150 ;
        RECT 464.400 343.050 465.450 352.950 ;
        RECT 473.400 346.050 474.450 397.950 ;
        RECT 478.950 382.950 481.050 385.050 ;
        RECT 478.950 380.850 481.050 381.750 ;
        RECT 472.950 343.950 475.050 346.050 ;
        RECT 478.950 344.250 481.050 345.150 ;
        RECT 473.400 343.050 474.450 343.950 ;
        RECT 457.950 340.950 460.050 343.050 ;
        RECT 461.250 341.250 462.750 342.150 ;
        RECT 463.950 340.950 466.050 343.050 ;
        RECT 467.250 341.250 469.050 342.150 ;
        RECT 469.950 341.250 471.750 342.150 ;
        RECT 472.950 340.950 475.050 343.050 ;
        RECT 476.250 341.250 477.750 342.150 ;
        RECT 478.950 340.950 481.050 343.050 ;
        RECT 458.400 340.050 459.450 340.950 ;
        RECT 479.400 340.050 480.450 340.950 ;
        RECT 457.950 337.950 460.050 340.050 ;
        RECT 460.950 337.950 463.050 340.050 ;
        RECT 464.250 338.850 465.750 339.750 ;
        RECT 466.950 337.950 469.050 340.050 ;
        RECT 469.950 337.950 472.050 340.050 ;
        RECT 473.250 338.850 474.750 339.750 ;
        RECT 475.950 337.950 478.050 340.050 ;
        RECT 478.950 337.950 481.050 340.050 ;
        RECT 467.400 331.050 468.450 337.950 ;
        RECT 466.950 328.950 469.050 331.050 ;
        RECT 449.400 244.050 450.450 316.950 ;
        RECT 452.250 305.400 453.450 317.400 ;
        RECT 454.950 316.950 457.050 319.050 ;
        RECT 454.950 314.250 457.050 315.150 ;
        RECT 457.950 313.950 460.050 316.050 ;
        RECT 467.400 315.450 468.450 328.950 ;
        RECT 470.400 328.050 471.450 337.950 ;
        RECT 482.400 334.050 483.450 400.950 ;
        RECT 484.950 388.950 487.050 391.050 ;
        RECT 485.400 385.050 486.450 388.950 ;
        RECT 484.950 382.950 487.050 385.050 ;
        RECT 484.950 380.850 487.050 381.750 ;
        RECT 488.400 370.050 489.450 404.400 ;
        RECT 494.400 394.050 495.450 448.950 ;
        RECT 497.400 444.600 498.600 461.400 ;
        RECT 505.950 460.950 508.050 463.050 ;
        RECT 509.400 457.050 510.450 463.950 ;
        RECT 515.400 457.050 516.450 481.950 ;
        RECT 521.400 481.050 522.450 496.950 ;
        RECT 524.400 490.050 525.450 520.950 ;
        RECT 529.950 499.950 532.050 502.050 ;
        RECT 530.400 490.050 531.450 499.950 ;
        RECT 539.400 499.050 540.450 523.950 ;
        RECT 538.950 496.950 541.050 499.050 ;
        RECT 545.400 498.450 546.450 544.950 ;
        RECT 547.950 535.950 550.050 538.050 ;
        RECT 548.400 532.050 549.450 535.950 ;
        RECT 550.950 532.950 553.050 535.050 ;
        RECT 547.950 529.950 550.050 532.050 ;
        RECT 551.400 529.050 552.450 532.950 ;
        RECT 563.400 532.050 564.450 556.950 ;
        RECT 572.400 550.050 573.450 586.950 ;
        RECT 574.950 566.400 577.050 568.500 ;
        RECT 571.950 547.950 574.050 550.050 ;
        RECT 575.400 549.600 576.600 566.400 ;
        RECT 580.950 557.250 583.050 558.150 ;
        RECT 583.950 556.950 586.050 559.050 ;
        RECT 586.950 557.250 589.050 558.150 ;
        RECT 580.950 553.950 583.050 556.050 ;
        RECT 584.400 552.450 585.450 556.950 ;
        RECT 586.950 553.950 589.050 556.050 ;
        RECT 581.400 551.400 585.450 552.450 ;
        RECT 574.950 547.500 577.050 549.600 ;
        RECT 571.950 538.950 574.050 541.050 ;
        RECT 562.950 529.950 565.050 532.050 ;
        RECT 572.400 529.050 573.450 538.950 ;
        RECT 547.950 527.850 549.750 528.750 ;
        RECT 550.950 526.950 553.050 529.050 ;
        RECT 565.950 528.450 568.050 529.050 ;
        RECT 556.950 527.250 559.050 528.150 ;
        RECT 563.400 527.400 568.050 528.450 ;
        RECT 563.400 526.050 564.450 527.400 ;
        RECT 565.950 526.950 568.050 527.400 ;
        RECT 569.250 527.250 570.750 528.150 ;
        RECT 571.950 526.950 574.050 529.050 ;
        RECT 575.250 527.250 576.750 528.150 ;
        RECT 577.950 526.950 580.050 529.050 ;
        RECT 550.950 524.850 553.050 525.750 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 562.950 523.950 565.050 526.050 ;
        RECT 565.950 524.850 567.750 525.750 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 572.250 524.850 573.750 525.750 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 578.250 524.850 580.050 525.750 ;
        RECT 575.400 520.050 576.450 523.950 ;
        RECT 565.950 517.950 568.050 520.050 ;
        RECT 574.950 517.950 577.050 520.050 ;
        RECT 566.400 499.050 567.450 517.950 ;
        RECT 581.400 511.050 582.450 551.400 ;
        RECT 587.400 538.050 588.450 553.950 ;
        RECT 586.950 535.950 589.050 538.050 ;
        RECT 593.400 532.050 594.450 602.400 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 605.400 601.050 606.450 607.950 ;
        RECT 598.950 600.450 601.050 601.050 ;
        RECT 596.400 599.400 601.050 600.450 ;
        RECT 602.250 599.850 603.750 600.750 ;
        RECT 596.400 595.050 597.450 599.400 ;
        RECT 598.950 598.950 601.050 599.400 ;
        RECT 604.950 598.950 607.050 601.050 ;
        RECT 607.950 598.950 610.050 601.050 ;
        RECT 598.950 596.850 601.050 597.750 ;
        RECT 604.950 596.850 607.050 597.750 ;
        RECT 607.950 596.850 610.050 597.750 ;
        RECT 595.950 592.950 598.050 595.050 ;
        RECT 611.400 594.450 612.450 607.950 ;
        RECT 614.400 607.050 615.450 607.950 ;
        RECT 613.950 604.950 616.050 607.050 ;
        RECT 616.950 598.950 619.050 601.050 ;
        RECT 613.950 596.250 616.050 597.150 ;
        RECT 616.950 596.850 619.050 597.750 ;
        RECT 613.950 594.450 616.050 595.050 ;
        RECT 620.400 594.450 621.450 607.950 ;
        RECT 622.950 601.950 625.050 604.050 ;
        RECT 623.400 601.050 624.450 601.950 ;
        RECT 622.950 598.950 625.050 601.050 ;
        RECT 626.250 599.250 627.750 600.150 ;
        RECT 628.950 598.950 631.050 601.050 ;
        RECT 632.400 598.050 633.450 613.950 ;
        RECT 622.950 596.850 624.750 597.750 ;
        RECT 625.950 595.950 628.050 598.050 ;
        RECT 629.250 596.850 630.750 597.750 ;
        RECT 631.950 595.950 634.050 598.050 ;
        RECT 611.400 593.400 616.050 594.450 ;
        RECT 613.950 592.950 616.050 593.400 ;
        RECT 617.400 593.400 621.450 594.450 ;
        RECT 631.950 593.850 634.050 594.750 ;
        RECT 607.950 574.950 610.050 577.050 ;
        RECT 595.950 567.300 598.050 569.400 ;
        RECT 596.250 563.700 597.450 567.300 ;
        RECT 595.950 561.600 598.050 563.700 ;
        RECT 596.250 549.600 597.450 561.600 ;
        RECT 604.950 557.250 607.050 558.150 ;
        RECT 598.950 555.450 601.050 556.050 ;
        RECT 598.950 554.400 603.450 555.450 ;
        RECT 598.950 553.950 601.050 554.400 ;
        RECT 598.950 551.850 601.050 552.750 ;
        RECT 595.950 547.500 598.050 549.600 ;
        RECT 598.950 533.400 601.050 535.500 ;
        RECT 586.950 529.950 589.050 532.050 ;
        RECT 592.950 529.950 595.050 532.050 ;
        RECT 595.950 530.250 598.050 531.150 ;
        RECT 587.400 526.050 588.450 529.950 ;
        RECT 592.950 526.950 595.050 529.050 ;
        RECT 595.950 526.950 598.050 529.050 ;
        RECT 583.950 524.250 585.750 525.150 ;
        RECT 586.950 523.950 589.050 526.050 ;
        RECT 590.250 524.250 592.050 525.150 ;
        RECT 583.950 520.950 586.050 523.050 ;
        RECT 587.250 521.850 588.750 522.750 ;
        RECT 589.950 520.950 592.050 523.050 ;
        RECT 584.400 520.050 585.450 520.950 ;
        RECT 590.400 520.050 591.450 520.950 ;
        RECT 583.950 517.950 586.050 520.050 ;
        RECT 589.950 517.950 592.050 520.050 ;
        RECT 580.950 508.950 583.050 511.050 ;
        RECT 545.400 497.400 549.450 498.450 ;
        RECT 539.400 496.050 540.450 496.950 ;
        RECT 535.950 493.950 538.050 496.050 ;
        RECT 538.950 493.950 541.050 496.050 ;
        RECT 544.950 493.950 547.050 496.050 ;
        RECT 536.400 490.050 537.450 493.950 ;
        RECT 523.950 487.950 526.050 490.050 ;
        RECT 527.250 488.250 528.750 489.150 ;
        RECT 529.950 487.950 532.050 490.050 ;
        RECT 535.950 487.950 538.050 490.050 ;
        RECT 539.250 488.250 540.750 489.150 ;
        RECT 541.950 487.950 544.050 490.050 ;
        RECT 523.950 485.850 525.750 486.750 ;
        RECT 526.950 484.950 529.050 487.050 ;
        RECT 530.250 485.850 532.050 486.750 ;
        RECT 535.950 485.850 537.750 486.750 ;
        RECT 538.950 484.950 541.050 487.050 ;
        RECT 542.250 485.850 544.050 486.750 ;
        RECT 520.950 478.950 523.050 481.050 ;
        RECT 517.950 461.400 520.050 463.500 ;
        RECT 502.950 454.950 505.050 457.050 ;
        RECT 508.950 454.950 511.050 457.050 ;
        RECT 514.950 454.950 517.050 457.050 ;
        RECT 502.950 452.850 505.050 453.750 ;
        RECT 508.950 452.850 511.050 453.750 ;
        RECT 508.950 448.950 511.050 451.050 ;
        RECT 518.250 449.400 519.450 461.400 ;
        RECT 523.950 460.950 526.050 463.050 ;
        RECT 520.950 458.250 523.050 459.150 ;
        RECT 520.950 456.450 523.050 457.050 ;
        RECT 524.400 456.450 525.450 460.950 ;
        RECT 520.950 455.400 525.450 456.450 ;
        RECT 520.950 454.950 523.050 455.400 ;
        RECT 496.950 442.500 499.050 444.600 ;
        RECT 505.950 442.950 508.050 445.050 ;
        RECT 496.950 423.300 499.050 425.400 ;
        RECT 497.250 419.700 498.450 423.300 ;
        RECT 496.950 417.600 499.050 419.700 ;
        RECT 497.250 405.600 498.450 417.600 ;
        RECT 499.950 411.450 502.050 412.050 ;
        RECT 499.950 410.400 504.450 411.450 ;
        RECT 499.950 409.950 502.050 410.400 ;
        RECT 499.950 407.850 502.050 408.750 ;
        RECT 496.950 403.500 499.050 405.600 ;
        RECT 493.950 391.950 496.050 394.050 ;
        RECT 503.400 388.050 504.450 410.400 ;
        RECT 499.950 385.950 502.050 388.050 ;
        RECT 502.950 385.950 505.050 388.050 ;
        RECT 500.400 385.050 501.450 385.950 ;
        RECT 506.400 385.050 507.450 442.950 ;
        RECT 509.400 415.050 510.450 448.950 ;
        RECT 517.950 447.300 520.050 449.400 ;
        RECT 518.250 443.700 519.450 447.300 ;
        RECT 514.950 439.950 517.050 442.050 ;
        RECT 517.950 441.600 520.050 443.700 ;
        RECT 508.950 412.950 511.050 415.050 ;
        RECT 508.950 410.850 511.050 411.750 ;
        RECT 511.950 410.250 514.050 411.150 ;
        RECT 515.400 409.050 516.450 439.950 ;
        RECT 527.400 420.450 528.450 484.950 ;
        RECT 545.400 472.050 546.450 493.950 ;
        RECT 548.400 490.050 549.450 497.400 ;
        RECT 565.950 496.950 568.050 499.050 ;
        RECT 566.400 490.050 567.450 496.950 ;
        RECT 593.400 493.050 594.450 526.950 ;
        RECT 596.400 493.050 597.450 526.950 ;
        RECT 599.550 521.400 600.750 533.400 ;
        RECT 598.950 519.300 601.050 521.400 ;
        RECT 602.400 520.050 603.450 554.400 ;
        RECT 604.950 553.950 607.050 556.050 ;
        RECT 608.400 555.450 609.450 574.950 ;
        RECT 610.950 557.250 613.050 558.150 ;
        RECT 610.950 555.450 613.050 556.050 ;
        RECT 608.400 554.400 613.050 555.450 ;
        RECT 610.950 553.950 613.050 554.400 ;
        RECT 617.400 555.450 618.450 593.400 ;
        RECT 635.400 580.050 636.450 613.950 ;
        RECT 634.950 577.950 637.050 580.050 ;
        RECT 638.400 562.050 639.450 617.400 ;
        RECT 644.400 616.050 645.450 664.950 ;
        RECT 659.400 661.050 660.450 670.950 ;
        RECT 662.550 665.400 663.750 677.400 ;
        RECT 670.950 672.450 673.050 673.050 ;
        RECT 670.950 671.400 675.450 672.450 ;
        RECT 670.950 670.950 673.050 671.400 ;
        RECT 670.950 668.850 673.050 669.750 ;
        RECT 661.950 663.300 664.050 665.400 ;
        RECT 658.950 658.950 661.050 661.050 ;
        RECT 662.550 659.700 663.750 663.300 ;
        RECT 661.950 657.600 664.050 659.700 ;
        RECT 646.950 628.950 649.050 631.050 ;
        RECT 649.950 629.250 652.050 630.150 ;
        RECT 655.950 629.250 658.050 630.150 ;
        RECT 661.950 629.250 663.750 630.150 ;
        RECT 664.950 628.950 667.050 631.050 ;
        RECT 670.950 628.950 673.050 631.050 ;
        RECT 647.400 621.450 648.450 628.950 ;
        RECT 649.950 625.950 652.050 628.050 ;
        RECT 653.250 626.250 654.750 627.150 ;
        RECT 655.950 625.950 658.050 628.050 ;
        RECT 661.950 625.950 664.050 628.050 ;
        RECT 665.250 626.850 667.050 627.750 ;
        RECT 667.950 626.250 670.050 627.150 ;
        RECT 670.950 626.850 673.050 627.750 ;
        RECT 650.400 625.050 651.450 625.950 ;
        RECT 649.950 622.950 652.050 625.050 ;
        RECT 652.950 622.950 655.050 625.050 ;
        RECT 653.400 621.450 654.450 622.950 ;
        RECT 647.400 620.400 654.450 621.450 ;
        RECT 656.400 619.050 657.450 625.950 ;
        RECT 662.400 619.050 663.450 625.950 ;
        RECT 667.950 622.950 670.050 625.050 ;
        RECT 674.400 622.050 675.450 671.400 ;
        RECT 676.950 670.950 679.050 673.050 ;
        RECT 676.950 668.850 679.050 669.750 ;
        RECT 683.400 660.600 684.600 677.400 ;
        RECT 691.950 676.950 694.050 679.050 ;
        RECT 692.400 673.050 693.450 676.950 ;
        RECT 691.950 670.950 694.050 673.050 ;
        RECT 691.950 668.850 694.050 669.750 ;
        RECT 697.950 668.850 700.050 669.750 ;
        RECT 700.950 667.950 703.050 670.050 ;
        RECT 703.950 668.250 705.750 669.150 ;
        RECT 706.950 667.950 709.050 670.050 ;
        RECT 710.250 668.250 712.050 669.150 ;
        RECT 691.950 664.950 694.050 667.050 ;
        RECT 682.950 658.500 685.050 660.600 ;
        RECT 679.950 639.300 682.050 641.400 ;
        RECT 680.550 635.700 681.750 639.300 ;
        RECT 679.950 633.600 682.050 635.700 ;
        RECT 682.950 634.950 685.050 637.050 ;
        RECT 676.950 625.950 679.050 628.050 ;
        RECT 676.950 623.850 679.050 624.750 ;
        RECT 673.950 619.950 676.050 622.050 ;
        RECT 676.950 619.950 679.050 622.050 ;
        RECT 680.550 621.600 681.750 633.600 ;
        RECT 655.950 616.950 658.050 619.050 ;
        RECT 661.950 616.950 664.050 619.050 ;
        RECT 643.950 613.950 646.050 616.050 ;
        RECT 667.950 605.400 670.050 607.500 ;
        RECT 658.950 603.450 661.050 604.050 ;
        RECT 658.950 602.400 663.450 603.450 ;
        RECT 658.950 601.950 661.050 602.400 ;
        RECT 640.950 598.950 643.050 601.050 ;
        RECT 643.950 598.950 646.050 601.050 ;
        RECT 649.950 600.450 652.050 601.050 ;
        RECT 647.250 599.250 648.750 600.150 ;
        RECT 649.950 599.400 654.450 600.450 ;
        RECT 649.950 598.950 652.050 599.400 ;
        RECT 641.400 598.050 642.450 598.950 ;
        RECT 640.950 595.950 643.050 598.050 ;
        RECT 644.250 596.850 645.750 597.750 ;
        RECT 646.950 595.950 649.050 598.050 ;
        RECT 650.250 596.850 652.050 597.750 ;
        RECT 653.400 597.450 654.450 599.400 ;
        RECT 655.950 599.250 658.050 600.150 ;
        RECT 658.950 599.850 661.050 600.750 ;
        RECT 662.400 600.450 663.450 602.400 ;
        RECT 664.950 602.250 667.050 603.150 ;
        RECT 664.950 600.450 667.050 601.050 ;
        RECT 662.400 599.400 667.050 600.450 ;
        RECT 664.950 598.950 667.050 599.400 ;
        RECT 655.950 597.450 658.050 598.050 ;
        RECT 653.400 596.400 658.050 597.450 ;
        RECT 655.950 595.950 658.050 596.400 ;
        RECT 661.950 595.950 664.050 598.050 ;
        RECT 640.950 593.850 643.050 594.750 ;
        RECT 643.950 577.950 646.050 580.050 ;
        RECT 637.950 559.950 640.050 562.050 ;
        RECT 619.950 557.250 622.050 558.150 ;
        RECT 625.950 557.250 628.050 558.150 ;
        RECT 628.950 556.950 631.050 559.050 ;
        RECT 634.950 556.950 637.050 559.050 ;
        RECT 638.250 557.250 640.050 558.150 ;
        RECT 640.950 556.950 643.050 559.050 ;
        RECT 619.950 555.450 622.050 556.050 ;
        RECT 617.400 554.400 622.050 555.450 ;
        RECT 605.400 535.050 606.450 553.950 ;
        RECT 617.400 550.050 618.450 554.400 ;
        RECT 619.950 553.950 622.050 554.400 ;
        RECT 623.250 554.250 624.750 555.150 ;
        RECT 625.950 553.950 628.050 556.050 ;
        RECT 628.950 554.850 631.050 555.750 ;
        RECT 631.950 554.250 634.050 555.150 ;
        RECT 634.950 554.850 636.750 555.750 ;
        RECT 637.950 553.950 640.050 556.050 ;
        RECT 622.950 550.950 625.050 553.050 ;
        RECT 616.950 547.950 619.050 550.050 ;
        RECT 613.950 538.950 616.050 541.050 ;
        RECT 607.950 535.950 610.050 538.050 ;
        RECT 604.950 532.950 607.050 535.050 ;
        RECT 604.950 529.950 607.050 532.050 ;
        RECT 599.550 515.700 600.750 519.300 ;
        RECT 601.950 517.950 604.050 520.050 ;
        RECT 598.950 513.600 601.050 515.700 ;
        RECT 583.950 490.950 586.050 493.050 ;
        RECT 586.950 490.950 589.050 493.050 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 595.950 490.950 598.050 493.050 ;
        RECT 601.950 490.950 604.050 493.050 ;
        RECT 547.950 487.950 550.050 490.050 ;
        RECT 551.250 488.250 552.750 489.150 ;
        RECT 553.950 487.950 556.050 490.050 ;
        RECT 559.950 489.450 562.050 490.050 ;
        RECT 557.400 488.400 562.050 489.450 ;
        RECT 547.950 485.850 549.750 486.750 ;
        RECT 550.950 484.950 553.050 487.050 ;
        RECT 554.250 485.850 556.050 486.750 ;
        RECT 535.950 469.950 538.050 472.050 ;
        RECT 544.950 469.950 547.050 472.050 ;
        RECT 532.950 461.400 535.050 463.500 ;
        RECT 533.400 444.600 534.600 461.400 ;
        RECT 532.950 442.500 535.050 444.600 ;
        RECT 527.400 419.400 531.450 420.450 ;
        RECT 530.400 418.050 531.450 419.400 ;
        RECT 529.950 415.950 532.050 418.050 ;
        RECT 532.950 415.950 535.050 418.050 ;
        RECT 533.400 415.050 534.450 415.950 ;
        RECT 517.950 413.250 520.050 414.150 ;
        RECT 523.950 413.250 526.050 414.150 ;
        RECT 529.950 413.250 531.750 414.150 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 517.950 409.950 520.050 412.050 ;
        RECT 521.250 410.250 522.750 411.150 ;
        RECT 523.950 409.950 526.050 412.050 ;
        RECT 529.950 409.950 532.050 412.050 ;
        RECT 533.250 410.850 535.050 411.750 ;
        RECT 511.950 406.950 514.050 409.050 ;
        RECT 514.950 406.950 517.050 409.050 ;
        RECT 512.400 385.050 513.450 406.950 ;
        RECT 518.400 403.050 519.450 409.950 ;
        RECT 520.950 406.950 523.050 409.050 ;
        RECT 517.950 400.950 520.050 403.050 ;
        RECT 521.400 397.050 522.450 406.950 ;
        RECT 523.950 403.950 526.050 406.050 ;
        RECT 517.950 394.950 520.050 397.050 ;
        RECT 520.950 394.950 523.050 397.050 ;
        RECT 518.400 385.050 519.450 394.950 ;
        RECT 520.950 388.950 523.050 391.050 ;
        RECT 521.400 385.050 522.450 388.950 ;
        RECT 524.400 385.050 525.450 403.950 ;
        RECT 530.400 400.050 531.450 409.950 ;
        RECT 529.950 397.950 532.050 400.050 ;
        RECT 529.950 391.950 532.050 394.050 ;
        RECT 499.950 382.950 502.050 385.050 ;
        RECT 503.250 383.250 504.750 384.150 ;
        RECT 505.950 382.950 508.050 385.050 ;
        RECT 509.250 383.250 510.750 384.150 ;
        RECT 511.950 382.950 514.050 385.050 ;
        RECT 517.950 382.950 520.050 385.050 ;
        RECT 520.950 382.950 523.050 385.050 ;
        RECT 523.950 382.950 526.050 385.050 ;
        RECT 490.950 380.250 492.750 381.150 ;
        RECT 493.950 379.950 496.050 382.050 ;
        RECT 497.250 380.250 499.050 381.150 ;
        RECT 499.950 380.850 501.750 381.750 ;
        RECT 502.950 379.950 505.050 382.050 ;
        RECT 506.250 380.850 507.750 381.750 ;
        RECT 508.950 379.950 511.050 382.050 ;
        RECT 512.250 380.850 514.050 381.750 ;
        RECT 517.950 380.850 520.050 381.750 ;
        RECT 490.950 376.950 493.050 379.050 ;
        RECT 494.250 377.850 495.750 378.750 ;
        RECT 496.950 376.950 499.050 379.050 ;
        RECT 491.400 376.050 492.450 376.950 ;
        RECT 490.950 373.950 493.050 376.050 ;
        RECT 487.950 367.950 490.050 370.050 ;
        RECT 490.950 351.300 493.050 353.400 ;
        RECT 491.550 347.700 492.750 351.300 ;
        RECT 490.950 345.600 493.050 347.700 ;
        RECT 493.950 346.950 496.050 349.050 ;
        RECT 484.950 337.950 487.050 340.050 ;
        RECT 487.950 337.950 490.050 340.050 ;
        RECT 481.950 331.950 484.050 334.050 ;
        RECT 469.950 325.950 472.050 328.050 ;
        RECT 475.950 325.950 478.050 328.050 ;
        RECT 469.950 315.450 472.050 316.050 ;
        RECT 467.400 314.400 472.050 315.450 ;
        RECT 469.950 313.950 472.050 314.400 ;
        RECT 454.950 312.450 457.050 313.050 ;
        RECT 458.400 312.450 459.450 313.950 ;
        RECT 476.400 313.050 477.450 325.950 ;
        RECT 478.950 316.950 481.050 319.050 ;
        RECT 479.400 316.050 480.450 316.950 ;
        RECT 478.950 313.950 481.050 316.050 ;
        RECT 481.950 313.950 484.050 316.050 ;
        RECT 482.400 313.050 483.450 313.950 ;
        RECT 454.950 311.400 459.450 312.450 ;
        RECT 454.950 310.950 457.050 311.400 ;
        RECT 451.950 303.300 454.050 305.400 ;
        RECT 452.250 299.700 453.450 303.300 ;
        RECT 451.950 297.600 454.050 299.700 ;
        RECT 458.400 274.050 459.450 311.400 ;
        RECT 463.950 310.950 466.050 313.050 ;
        RECT 467.250 311.250 469.050 312.150 ;
        RECT 469.950 311.850 472.050 312.750 ;
        RECT 472.950 311.250 475.050 312.150 ;
        RECT 475.950 310.950 478.050 313.050 ;
        RECT 479.250 311.850 480.750 312.750 ;
        RECT 481.950 310.950 484.050 313.050 ;
        RECT 463.950 308.850 465.750 309.750 ;
        RECT 466.950 307.950 469.050 310.050 ;
        RECT 469.950 307.950 472.050 310.050 ;
        RECT 472.950 307.950 475.050 310.050 ;
        RECT 475.950 308.850 478.050 309.750 ;
        RECT 481.950 308.850 484.050 309.750 ;
        RECT 467.400 307.050 468.450 307.950 ;
        RECT 466.950 304.950 469.050 307.050 ;
        RECT 470.400 301.050 471.450 307.950 ;
        RECT 469.950 298.950 472.050 301.050 ;
        RECT 466.950 279.300 469.050 281.400 ;
        RECT 467.550 275.700 468.750 279.300 ;
        RECT 472.950 277.950 475.050 280.050 ;
        RECT 457.950 271.950 460.050 274.050 ;
        RECT 466.950 273.600 469.050 275.700 ;
        RECT 451.950 269.250 454.050 270.150 ;
        RECT 457.950 269.250 460.050 270.150 ;
        RECT 451.950 265.950 454.050 268.050 ;
        RECT 455.250 266.250 456.750 267.150 ;
        RECT 457.950 265.950 460.050 268.050 ;
        RECT 460.950 265.950 463.050 268.050 ;
        RECT 463.950 265.950 466.050 268.050 ;
        RECT 452.400 244.050 453.450 265.950 ;
        RECT 454.950 262.950 457.050 265.050 ;
        RECT 461.400 244.050 462.450 265.950 ;
        RECT 463.950 263.850 466.050 264.750 ;
        RECT 467.550 261.600 468.750 273.600 ;
        RECT 469.950 271.950 472.050 274.050 ;
        RECT 466.950 259.500 469.050 261.600 ;
        RECT 470.400 256.050 471.450 271.950 ;
        RECT 473.400 267.450 474.450 277.950 ;
        RECT 475.950 269.250 478.050 270.150 ;
        RECT 481.950 269.250 484.050 270.150 ;
        RECT 475.950 267.450 478.050 268.050 ;
        RECT 473.400 266.400 478.050 267.450 ;
        RECT 475.950 265.950 478.050 266.400 ;
        RECT 481.950 265.950 484.050 268.050 ;
        RECT 469.950 253.950 472.050 256.050 ;
        RECT 482.400 247.050 483.450 265.950 ;
        RECT 469.950 244.950 472.050 247.050 ;
        RECT 481.950 244.950 484.050 247.050 ;
        RECT 448.950 241.950 451.050 244.050 ;
        RECT 451.950 243.450 454.050 244.050 ;
        RECT 451.950 242.400 456.450 243.450 ;
        RECT 451.950 241.950 454.050 242.400 ;
        RECT 448.950 239.250 451.050 240.150 ;
        RECT 451.950 239.850 454.050 240.750 ;
        RECT 448.950 235.950 451.050 238.050 ;
        RECT 455.400 213.450 456.450 242.400 ;
        RECT 460.950 241.950 463.050 244.050 ;
        RECT 470.400 241.050 471.450 244.950 ;
        RECT 485.400 241.050 486.450 337.950 ;
        RECT 487.950 335.850 490.050 336.750 ;
        RECT 491.550 333.600 492.750 345.600 ;
        RECT 490.950 331.500 493.050 333.600 ;
        RECT 494.400 331.050 495.450 346.950 ;
        RECT 499.950 341.250 502.050 342.150 ;
        RECT 499.950 337.950 502.050 340.050 ;
        RECT 500.400 337.050 501.450 337.950 ;
        RECT 499.950 334.950 502.050 337.050 ;
        RECT 503.400 334.050 504.450 379.950 ;
        RECT 509.400 379.050 510.450 379.950 ;
        RECT 508.950 376.950 511.050 379.050 ;
        RECT 511.950 350.400 514.050 352.500 ;
        RECT 505.950 341.250 508.050 342.150 ;
        RECT 505.950 337.950 508.050 340.050 ;
        RECT 502.950 331.950 505.050 334.050 ;
        RECT 512.400 333.600 513.600 350.400 ;
        RECT 511.950 331.500 514.050 333.600 ;
        RECT 493.950 328.950 496.050 331.050 ;
        RECT 487.950 322.950 490.050 325.050 ;
        RECT 488.400 310.050 489.450 322.950 ;
        RECT 490.950 319.950 493.050 322.050 ;
        RECT 491.400 313.050 492.450 319.950 ;
        RECT 511.950 317.400 514.050 319.500 ;
        RECT 490.950 310.950 493.050 313.050 ;
        RECT 494.250 311.250 495.750 312.150 ;
        RECT 496.950 310.950 499.050 313.050 ;
        RECT 502.950 312.450 505.050 313.050 ;
        RECT 500.250 311.250 501.750 312.150 ;
        RECT 502.950 311.400 507.450 312.450 ;
        RECT 502.950 310.950 505.050 311.400 ;
        RECT 487.950 307.950 490.050 310.050 ;
        RECT 490.950 308.850 492.750 309.750 ;
        RECT 493.950 307.950 496.050 310.050 ;
        RECT 497.250 308.850 498.750 309.750 ;
        RECT 499.950 307.950 502.050 310.050 ;
        RECT 503.250 308.850 505.050 309.750 ;
        RECT 490.950 289.950 493.050 292.050 ;
        RECT 487.950 278.400 490.050 280.500 ;
        RECT 488.400 261.600 489.600 278.400 ;
        RECT 487.950 259.500 490.050 261.600 ;
        RECT 487.950 253.950 490.050 256.050 ;
        RECT 457.950 239.250 460.050 240.150 ;
        RECT 460.950 239.850 463.050 240.750 ;
        RECT 463.950 238.950 466.050 241.050 ;
        RECT 467.250 239.250 468.750 240.150 ;
        RECT 469.950 238.950 472.050 241.050 ;
        RECT 475.950 238.950 478.050 241.050 ;
        RECT 484.950 238.950 487.050 241.050 ;
        RECT 457.950 235.950 460.050 238.050 ;
        RECT 463.950 236.850 465.750 237.750 ;
        RECT 466.950 235.950 469.050 238.050 ;
        RECT 470.250 236.850 471.750 237.750 ;
        RECT 472.950 235.950 475.050 238.050 ;
        RECT 472.950 233.850 475.050 234.750 ;
        RECT 476.400 232.050 477.450 238.950 ;
        RECT 478.950 236.250 480.750 237.150 ;
        RECT 481.950 235.950 484.050 238.050 ;
        RECT 485.250 236.250 487.050 237.150 ;
        RECT 478.950 232.950 481.050 235.050 ;
        RECT 482.250 233.850 483.750 234.750 ;
        RECT 484.950 232.950 487.050 235.050 ;
        RECT 479.400 232.050 480.450 232.950 ;
        RECT 475.950 229.950 478.050 232.050 ;
        RECT 478.950 229.950 481.050 232.050 ;
        RECT 452.400 212.400 456.450 213.450 ;
        RECT 445.950 202.950 448.050 205.050 ;
        RECT 439.950 197.250 442.050 198.150 ;
        RECT 445.950 197.250 448.050 198.150 ;
        RECT 448.950 196.950 451.050 199.050 ;
        RECT 439.950 193.950 442.050 196.050 ;
        RECT 445.950 193.950 448.050 196.050 ;
        RECT 440.400 190.050 441.450 193.950 ;
        RECT 446.400 193.050 447.450 193.950 ;
        RECT 445.950 190.950 448.050 193.050 ;
        RECT 439.950 187.950 442.050 190.050 ;
        RECT 442.950 173.400 445.050 175.500 ;
        RECT 446.400 175.050 447.450 190.950 ;
        RECT 443.250 161.400 444.450 173.400 ;
        RECT 445.950 172.950 448.050 175.050 ;
        RECT 449.400 172.050 450.450 196.950 ;
        RECT 445.950 170.250 448.050 171.150 ;
        RECT 448.950 169.950 451.050 172.050 ;
        RECT 445.950 166.950 448.050 169.050 ;
        RECT 449.400 162.450 450.450 169.950 ;
        RECT 452.400 169.050 453.450 212.400 ;
        RECT 454.950 207.300 457.050 209.400 ;
        RECT 488.400 208.050 489.450 253.950 ;
        RECT 455.250 203.700 456.450 207.300 ;
        RECT 487.950 205.950 490.050 208.050 ;
        RECT 454.950 201.600 457.050 203.700 ;
        RECT 475.950 202.950 478.050 205.050 ;
        RECT 487.950 202.950 490.050 205.050 ;
        RECT 455.250 189.600 456.450 201.600 ;
        RECT 463.950 199.950 466.050 202.050 ;
        RECT 457.950 193.950 460.050 196.050 ;
        RECT 460.950 193.950 463.050 196.050 ;
        RECT 457.950 191.850 460.050 192.750 ;
        RECT 454.950 187.500 457.050 189.600 ;
        RECT 451.950 166.950 454.050 169.050 ;
        RECT 451.950 164.250 453.750 165.150 ;
        RECT 454.950 163.950 457.050 166.050 ;
        RECT 458.250 164.250 460.050 165.150 ;
        RECT 451.950 162.450 454.050 163.050 ;
        RECT 449.400 161.400 454.050 162.450 ;
        RECT 455.250 161.850 456.750 162.750 ;
        RECT 457.950 162.450 460.050 163.050 ;
        RECT 461.400 162.450 462.450 193.950 ;
        RECT 464.400 192.450 465.450 199.950 ;
        RECT 466.950 197.250 469.050 198.150 ;
        RECT 472.950 197.250 475.050 198.150 ;
        RECT 466.950 193.950 469.050 196.050 ;
        RECT 472.950 195.450 475.050 196.050 ;
        RECT 476.400 195.450 477.450 202.950 ;
        RECT 481.950 199.950 484.050 202.050 ;
        RECT 482.400 199.050 483.450 199.950 ;
        RECT 488.400 199.050 489.450 202.950 ;
        RECT 478.950 197.250 480.750 198.150 ;
        RECT 481.950 196.950 484.050 199.050 ;
        RECT 487.950 196.950 490.050 199.050 ;
        RECT 470.250 194.250 471.750 195.150 ;
        RECT 472.950 194.400 477.450 195.450 ;
        RECT 472.950 193.950 475.050 194.400 ;
        RECT 478.950 193.950 481.050 196.050 ;
        RECT 482.250 194.850 484.050 195.750 ;
        RECT 484.950 194.250 487.050 195.150 ;
        RECT 487.950 194.850 490.050 195.750 ;
        RECT 469.950 192.450 472.050 193.050 ;
        RECT 464.400 191.400 472.050 192.450 ;
        RECT 469.950 190.950 472.050 191.400 ;
        RECT 479.400 190.050 480.450 193.950 ;
        RECT 484.950 190.950 487.050 193.050 ;
        RECT 485.400 190.050 486.450 190.950 ;
        RECT 478.950 187.950 481.050 190.050 ;
        RECT 484.950 187.950 487.050 190.050 ;
        RECT 491.400 181.050 492.450 289.950 ;
        RECT 500.400 277.050 501.450 307.950 ;
        RECT 506.400 307.050 507.450 311.400 ;
        RECT 505.950 304.950 508.050 307.050 ;
        RECT 512.400 300.600 513.600 317.400 ;
        RECT 517.950 310.950 520.050 313.050 ;
        RECT 517.950 308.850 520.050 309.750 ;
        RECT 511.950 298.500 514.050 300.600 ;
        RECT 493.950 274.950 496.050 277.050 ;
        RECT 499.950 274.950 502.050 277.050 ;
        RECT 517.950 274.950 520.050 277.050 ;
        RECT 494.400 267.450 495.450 274.950 ;
        RECT 518.400 274.050 519.450 274.950 ;
        RECT 505.950 272.250 508.050 273.150 ;
        RECT 511.950 271.950 514.050 274.050 ;
        RECT 515.250 272.250 516.750 273.150 ;
        RECT 517.950 271.950 520.050 274.050 ;
        RECT 496.950 269.250 498.750 270.150 ;
        RECT 499.950 268.950 502.050 271.050 ;
        RECT 503.250 269.250 504.750 270.150 ;
        RECT 505.950 268.950 508.050 271.050 ;
        RECT 511.950 269.850 513.750 270.750 ;
        RECT 514.950 268.950 517.050 271.050 ;
        RECT 518.250 269.850 520.050 270.750 ;
        RECT 496.950 267.450 499.050 268.050 ;
        RECT 494.400 266.400 499.050 267.450 ;
        RECT 500.250 266.850 501.750 267.750 ;
        RECT 496.950 265.950 499.050 266.400 ;
        RECT 502.950 265.950 505.050 268.050 ;
        RECT 505.950 265.950 508.050 268.050 ;
        RECT 503.400 262.050 504.450 265.950 ;
        RECT 502.950 259.950 505.050 262.050 ;
        RECT 499.950 247.950 502.050 250.050 ;
        RECT 496.950 244.950 499.050 247.050 ;
        RECT 497.400 238.050 498.450 244.950 ;
        RECT 500.400 241.050 501.450 247.950 ;
        RECT 502.950 241.950 505.050 244.050 ;
        RECT 499.950 238.950 502.050 241.050 ;
        RECT 493.950 236.250 495.750 237.150 ;
        RECT 496.950 235.950 499.050 238.050 ;
        RECT 500.250 236.250 502.050 237.150 ;
        RECT 493.950 232.950 496.050 235.050 ;
        RECT 497.250 233.850 498.750 234.750 ;
        RECT 499.950 232.950 502.050 235.050 ;
        RECT 494.400 229.050 495.450 232.950 ;
        RECT 500.400 232.050 501.450 232.950 ;
        RECT 499.950 229.950 502.050 232.050 ;
        RECT 493.950 226.950 496.050 229.050 ;
        RECT 493.950 205.950 496.050 208.050 ;
        RECT 496.950 206.400 499.050 208.500 ;
        RECT 490.950 178.950 493.050 181.050 ;
        RECT 469.950 172.950 472.050 175.050 ;
        RECT 470.400 169.050 471.450 172.950 ;
        RECT 475.950 169.950 478.050 172.050 ;
        RECT 481.950 169.950 484.050 172.050 ;
        RECT 476.400 169.050 477.450 169.950 ;
        RECT 482.400 169.050 483.450 169.950 ;
        RECT 469.950 166.950 472.050 169.050 ;
        RECT 473.250 167.250 474.750 168.150 ;
        RECT 475.950 166.950 478.050 169.050 ;
        RECT 481.950 166.950 484.050 169.050 ;
        RECT 487.950 166.950 490.050 169.050 ;
        RECT 466.950 163.950 469.050 166.050 ;
        RECT 470.250 164.850 471.750 165.750 ;
        RECT 472.950 163.950 475.050 166.050 ;
        RECT 476.250 164.850 478.050 165.750 ;
        RECT 481.950 164.850 484.050 165.750 ;
        RECT 487.950 164.850 490.050 165.750 ;
        RECT 436.950 157.950 439.050 160.050 ;
        RECT 442.950 159.300 445.050 161.400 ;
        RECT 451.950 160.950 454.050 161.400 ;
        RECT 457.950 161.400 462.450 162.450 ;
        RECT 466.950 161.850 469.050 162.750 ;
        RECT 473.400 162.450 474.450 163.950 ;
        RECT 473.400 161.400 477.450 162.450 ;
        RECT 457.950 160.950 460.050 161.400 ;
        RECT 421.950 154.500 424.050 156.600 ;
        RECT 443.250 155.700 444.450 159.300 ;
        RECT 448.950 157.950 451.050 160.050 ;
        RECT 442.950 153.600 445.050 155.700 ;
        RECT 382.950 127.950 385.050 130.050 ;
        RECT 386.250 128.250 387.750 129.150 ;
        RECT 388.950 127.950 391.050 130.050 ;
        RECT 392.250 128.250 394.050 129.150 ;
        RECT 412.950 127.950 415.050 130.050 ;
        RECT 416.250 128.250 417.750 129.150 ;
        RECT 418.950 127.950 421.050 130.050 ;
        RECT 433.950 127.950 436.050 130.050 ;
        RECT 439.950 127.950 442.050 130.050 ;
        RECT 389.400 127.050 390.450 127.950 ;
        RECT 434.400 127.050 435.450 127.950 ;
        RECT 382.950 125.850 384.750 126.750 ;
        RECT 385.950 124.950 388.050 127.050 ;
        RECT 388.950 124.950 391.050 127.050 ;
        RECT 391.950 124.950 394.050 127.050 ;
        RECT 394.950 124.950 397.050 127.050 ;
        RECT 400.950 124.950 403.050 127.050 ;
        RECT 404.250 125.250 406.050 126.150 ;
        RECT 412.950 125.850 414.750 126.750 ;
        RECT 415.950 124.950 418.050 127.050 ;
        RECT 419.250 125.850 421.050 126.750 ;
        RECT 424.950 125.250 426.750 126.150 ;
        RECT 427.950 124.950 430.050 127.050 ;
        RECT 431.250 125.250 432.750 126.150 ;
        RECT 433.950 124.950 436.050 127.050 ;
        RECT 437.250 125.250 439.050 126.150 ;
        RECT 386.400 121.050 387.450 124.950 ;
        RECT 385.950 118.950 388.050 121.050 ;
        RECT 389.400 114.450 390.450 124.950 ;
        RECT 392.400 124.050 393.450 124.950 ;
        RECT 391.950 121.950 394.050 124.050 ;
        RECT 394.950 122.850 397.050 123.750 ;
        RECT 397.950 122.250 400.050 123.150 ;
        RECT 400.950 122.850 402.750 123.750 ;
        RECT 403.950 121.950 406.050 124.050 ;
        RECT 424.950 121.950 427.050 124.050 ;
        RECT 428.250 122.850 429.750 123.750 ;
        RECT 430.950 121.950 433.050 124.050 ;
        RECT 434.250 122.850 435.750 123.750 ;
        RECT 436.950 121.950 439.050 124.050 ;
        RECT 392.400 117.450 393.450 121.950 ;
        RECT 397.950 118.950 400.050 121.050 ;
        RECT 392.400 116.400 396.450 117.450 ;
        RECT 389.400 113.400 393.450 114.450 ;
        RECT 385.950 109.950 388.050 112.050 ;
        RECT 379.950 106.950 382.050 109.050 ;
        RECT 367.950 97.950 370.050 100.050 ;
        RECT 376.950 97.950 379.050 100.050 ;
        RECT 368.400 94.050 369.450 97.950 ;
        RECT 370.950 94.950 373.050 97.050 ;
        RECT 371.400 94.050 372.450 94.950 ;
        RECT 380.400 94.050 381.450 106.950 ;
        RECT 386.400 94.050 387.450 109.950 ;
        RECT 364.950 91.950 367.050 94.050 ;
        RECT 367.950 91.950 370.050 94.050 ;
        RECT 370.950 91.950 373.050 94.050 ;
        RECT 374.250 92.250 376.050 93.150 ;
        RECT 376.950 91.950 379.050 94.050 ;
        RECT 379.950 91.950 382.050 94.050 ;
        RECT 385.950 91.950 388.050 94.050 ;
        RECT 389.250 92.250 391.050 93.150 ;
        RECT 364.950 89.850 366.750 90.750 ;
        RECT 367.950 88.950 370.050 91.050 ;
        RECT 371.250 89.850 372.750 90.750 ;
        RECT 373.950 88.950 376.050 91.050 ;
        RECT 367.950 86.850 370.050 87.750 ;
        RECT 361.950 73.950 364.050 76.050 ;
        RECT 343.950 70.950 346.050 73.050 ;
        RECT 340.950 64.950 343.050 67.050 ;
        RECT 361.950 61.950 364.050 64.050 ;
        RECT 349.950 58.950 352.050 61.050 ;
        RECT 350.400 58.050 351.450 58.950 ;
        RECT 343.950 57.450 346.050 58.050 ;
        RECT 341.400 56.400 346.050 57.450 ;
        RECT 328.950 52.950 331.050 55.050 ;
        RECT 331.950 53.250 334.050 54.150 ;
        RECT 334.950 52.950 337.050 55.050 ;
        RECT 337.950 53.250 340.050 54.150 ;
        RECT 341.400 52.050 342.450 56.400 ;
        RECT 343.950 55.950 346.050 56.400 ;
        RECT 347.250 56.250 348.750 57.150 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 343.950 53.850 345.750 54.750 ;
        RECT 346.950 52.950 349.050 55.050 ;
        RECT 350.250 53.850 352.050 54.750 ;
        RECT 352.950 53.250 355.050 54.150 ;
        RECT 358.950 53.250 361.050 54.150 ;
        RECT 347.400 52.050 348.450 52.950 ;
        RECT 328.950 49.950 331.050 52.050 ;
        RECT 331.950 49.950 334.050 52.050 ;
        RECT 335.250 50.250 336.750 51.150 ;
        RECT 337.950 49.950 340.050 52.050 ;
        RECT 340.950 49.950 343.050 52.050 ;
        RECT 346.950 49.950 349.050 52.050 ;
        RECT 352.950 49.950 355.050 52.050 ;
        RECT 356.250 50.250 357.750 51.150 ;
        RECT 358.950 49.950 361.050 52.050 ;
        RECT 329.400 43.050 330.450 49.950 ;
        RECT 332.400 49.050 333.450 49.950 ;
        RECT 331.950 46.950 334.050 49.050 ;
        RECT 334.950 46.950 337.050 49.050 ;
        RECT 328.950 40.950 331.050 43.050 ;
        RECT 319.950 31.950 322.050 34.050 ;
        RECT 325.950 31.950 328.050 34.050 ;
        RECT 328.950 31.950 331.050 34.050 ;
        RECT 307.950 25.950 310.050 28.050 ;
        RECT 310.950 25.950 313.050 28.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 301.950 20.850 304.050 21.750 ;
        RECT 304.950 20.250 307.050 21.150 ;
        RECT 304.950 18.450 307.050 19.050 ;
        RECT 308.400 18.450 309.450 25.950 ;
        RECT 311.400 25.050 312.450 25.950 ;
        RECT 320.400 25.050 321.450 31.950 ;
        RECT 325.950 28.950 328.050 31.050 ;
        RECT 310.950 22.950 313.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 326.400 22.050 327.450 28.950 ;
        RECT 329.400 22.050 330.450 31.950 ;
        RECT 331.950 22.950 334.050 25.050 ;
        RECT 335.400 24.450 336.450 46.950 ;
        RECT 338.400 46.050 339.450 49.950 ;
        RECT 355.950 46.950 358.050 49.050 ;
        RECT 359.400 46.050 360.450 49.950 ;
        RECT 337.950 43.950 340.050 46.050 ;
        RECT 358.950 43.950 361.050 46.050 ;
        RECT 337.950 40.950 340.050 43.050 ;
        RECT 338.400 31.050 339.450 40.950 ;
        RECT 358.950 37.950 361.050 40.050 ;
        RECT 337.950 28.950 340.050 31.050 ;
        RECT 352.950 28.950 355.050 31.050 ;
        RECT 338.400 27.450 339.450 28.950 ;
        RECT 353.400 28.050 354.450 28.950 ;
        RECT 338.400 26.400 342.450 27.450 ;
        RECT 341.400 25.050 342.450 26.400 ;
        RECT 352.950 25.950 355.050 28.050 ;
        RECT 353.400 25.050 354.450 25.950 ;
        RECT 359.400 25.050 360.450 37.950 ;
        RECT 362.400 31.050 363.450 61.950 ;
        RECT 367.950 59.250 370.050 60.150 ;
        RECT 364.950 56.250 366.750 57.150 ;
        RECT 367.950 55.950 370.050 58.050 ;
        RECT 371.250 56.250 372.750 57.150 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 364.950 52.950 367.050 55.050 ;
        RECT 364.950 49.950 367.050 52.050 ;
        RECT 361.950 28.950 364.050 31.050 ;
        RECT 365.400 25.050 366.450 49.950 ;
        RECT 368.400 34.050 369.450 55.950 ;
        RECT 370.950 52.950 373.050 55.050 ;
        RECT 374.250 53.850 376.050 54.750 ;
        RECT 371.400 52.050 372.450 52.950 ;
        RECT 370.950 49.950 373.050 52.050 ;
        RECT 367.950 31.950 370.050 34.050 ;
        RECT 377.400 25.050 378.450 91.950 ;
        RECT 379.950 89.850 381.750 90.750 ;
        RECT 382.950 88.950 385.050 91.050 ;
        RECT 386.250 89.850 387.750 90.750 ;
        RECT 388.950 90.450 391.050 91.050 ;
        RECT 392.400 90.450 393.450 113.400 ;
        RECT 388.950 89.400 393.450 90.450 ;
        RECT 388.950 88.950 391.050 89.400 ;
        RECT 382.950 86.850 385.050 87.750 ;
        RECT 395.400 64.050 396.450 116.400 ;
        RECT 424.950 101.400 427.050 103.500 ;
        RECT 400.950 97.950 403.050 100.050 ;
        RECT 397.950 95.250 400.050 96.150 ;
        RECT 400.950 95.850 403.050 96.750 ;
        RECT 403.950 94.950 406.050 97.050 ;
        RECT 415.950 94.950 418.050 97.050 ;
        RECT 404.400 94.050 405.450 94.950 ;
        RECT 397.950 91.950 400.050 94.050 ;
        RECT 400.950 91.950 403.050 94.050 ;
        RECT 403.950 91.950 406.050 94.050 ;
        RECT 409.950 91.950 412.050 94.050 ;
        RECT 413.250 92.250 415.050 93.150 ;
        RECT 398.400 91.050 399.450 91.950 ;
        RECT 397.950 88.950 400.050 91.050 ;
        RECT 401.400 82.050 402.450 91.950 ;
        RECT 403.950 89.850 405.750 90.750 ;
        RECT 406.950 88.950 409.050 91.050 ;
        RECT 410.250 89.850 411.750 90.750 ;
        RECT 412.950 88.950 415.050 91.050 ;
        RECT 406.950 86.850 409.050 87.750 ;
        RECT 400.950 79.950 403.050 82.050 ;
        RECT 409.950 79.950 412.050 82.050 ;
        RECT 382.950 61.950 385.050 64.050 ;
        RECT 394.950 61.950 397.050 64.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 380.400 46.050 381.450 55.950 ;
        RECT 383.400 55.050 384.450 61.950 ;
        RECT 385.950 58.950 388.050 61.050 ;
        RECT 397.950 59.250 400.050 60.150 ;
        RECT 403.950 58.950 406.050 61.050 ;
        RECT 386.400 55.050 387.450 58.950 ;
        RECT 391.950 57.450 394.050 58.050 ;
        RECT 389.400 56.400 394.050 57.450 ;
        RECT 382.950 52.950 385.050 55.050 ;
        RECT 385.950 52.950 388.050 55.050 ;
        RECT 382.950 50.850 385.050 51.750 ;
        RECT 385.950 50.250 388.050 51.150 ;
        RECT 385.950 48.450 388.050 49.050 ;
        RECT 389.400 48.450 390.450 56.400 ;
        RECT 391.950 55.950 394.050 56.400 ;
        RECT 395.250 56.250 396.750 57.150 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 401.250 56.250 403.050 57.150 ;
        RECT 391.950 53.850 393.750 54.750 ;
        RECT 394.950 52.950 397.050 55.050 ;
        RECT 385.950 47.400 390.450 48.450 ;
        RECT 385.950 46.950 388.050 47.400 ;
        RECT 379.950 43.950 382.050 46.050 ;
        RECT 382.950 28.950 385.050 31.050 ;
        RECT 383.400 28.050 384.450 28.950 ;
        RECT 382.950 25.950 385.050 28.050 ;
        RECT 388.950 25.950 391.050 28.050 ;
        RECT 389.400 25.050 390.450 25.950 ;
        RECT 395.400 25.050 396.450 52.950 ;
        RECT 398.400 49.050 399.450 55.950 ;
        RECT 404.400 55.050 405.450 58.950 ;
        RECT 410.400 58.050 411.450 79.950 ;
        RECT 413.400 61.050 414.450 88.950 ;
        RECT 412.950 58.950 415.050 61.050 ;
        RECT 409.950 55.950 412.050 58.050 ;
        RECT 410.400 55.050 411.450 55.950 ;
        RECT 416.400 55.050 417.450 94.950 ;
        RECT 425.400 84.600 426.600 101.400 ;
        RECT 431.400 97.050 432.450 121.950 ;
        RECT 436.950 106.950 439.050 109.050 ;
        RECT 437.400 97.050 438.450 106.950 ;
        RECT 440.400 97.050 441.450 127.950 ;
        RECT 442.950 124.950 445.050 127.050 ;
        RECT 442.950 122.850 445.050 123.750 ;
        RECT 445.950 122.250 448.050 123.150 ;
        RECT 445.950 118.950 448.050 121.050 ;
        RECT 449.400 115.050 450.450 157.950 ;
        RECT 476.400 127.050 477.450 161.400 ;
        RECT 490.950 128.250 493.050 129.150 ;
        RECT 451.950 125.250 454.050 126.150 ;
        RECT 457.950 125.250 460.050 126.150 ;
        RECT 460.950 124.950 463.050 127.050 ;
        RECT 475.950 126.450 478.050 127.050 ;
        RECT 463.950 125.250 466.050 126.150 ;
        RECT 469.950 125.250 472.050 126.150 ;
        RECT 475.950 125.400 480.450 126.450 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 451.950 121.950 454.050 124.050 ;
        RECT 455.250 122.250 456.750 123.150 ;
        RECT 457.950 121.950 460.050 124.050 ;
        RECT 452.400 121.050 453.450 121.950 ;
        RECT 451.950 118.950 454.050 121.050 ;
        RECT 454.950 118.950 457.050 121.050 ;
        RECT 448.950 112.950 451.050 115.050 ;
        RECT 442.950 106.950 445.050 109.050 ;
        RECT 430.950 94.950 433.050 97.050 ;
        RECT 436.950 94.950 439.050 97.050 ;
        RECT 439.950 94.950 442.050 97.050 ;
        RECT 430.950 92.850 433.050 93.750 ;
        RECT 436.950 92.850 439.050 93.750 ;
        RECT 424.950 82.500 427.050 84.600 ;
        RECT 430.950 61.950 433.050 64.050 ;
        RECT 427.950 55.950 430.050 58.050 ;
        RECT 400.950 52.950 403.050 55.050 ;
        RECT 403.950 52.950 406.050 55.050 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 413.250 53.250 415.050 54.150 ;
        RECT 415.950 52.950 418.050 55.050 ;
        RECT 418.950 53.250 421.050 54.150 ;
        RECT 424.950 53.250 427.050 54.150 ;
        RECT 403.950 50.850 406.050 51.750 ;
        RECT 406.950 50.250 409.050 51.150 ;
        RECT 409.950 50.850 411.750 51.750 ;
        RECT 412.950 49.950 415.050 52.050 ;
        RECT 418.950 49.950 421.050 52.050 ;
        RECT 422.250 50.250 423.750 51.150 ;
        RECT 424.950 49.950 427.050 52.050 ;
        RECT 428.400 49.050 429.450 55.950 ;
        RECT 431.400 52.050 432.450 61.950 ;
        RECT 440.400 58.050 441.450 94.950 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 437.250 56.250 438.750 57.150 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 433.950 53.850 435.750 54.750 ;
        RECT 436.950 52.950 439.050 55.050 ;
        RECT 440.250 53.850 442.050 54.750 ;
        RECT 430.950 49.950 433.050 52.050 ;
        RECT 397.950 46.950 400.050 49.050 ;
        RECT 406.950 46.950 409.050 49.050 ;
        RECT 421.950 46.950 424.050 49.050 ;
        RECT 427.950 46.950 430.050 49.050 ;
        RECT 397.950 37.950 400.050 40.050 ;
        RECT 403.950 37.950 406.050 40.050 ;
        RECT 335.400 23.400 339.450 24.450 ;
        RECT 332.400 22.050 333.450 22.950 ;
        RECT 310.950 20.850 313.050 21.750 ;
        RECT 313.950 20.850 316.050 21.750 ;
        RECT 319.950 20.850 322.050 21.750 ;
        RECT 325.950 19.950 328.050 22.050 ;
        RECT 328.950 19.950 331.050 22.050 ;
        RECT 331.950 19.950 334.050 22.050 ;
        RECT 335.250 20.250 337.050 21.150 ;
        RECT 329.400 19.050 330.450 19.950 ;
        RECT 338.400 19.050 339.450 23.400 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 344.250 23.250 345.750 24.150 ;
        RECT 346.950 22.950 349.050 25.050 ;
        RECT 350.250 23.250 351.750 24.150 ;
        RECT 352.950 22.950 355.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 362.250 23.250 363.750 24.150 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 376.950 22.950 379.050 25.050 ;
        RECT 380.250 23.250 382.050 24.150 ;
        RECT 382.950 23.850 385.050 24.750 ;
        RECT 385.950 23.250 388.050 24.150 ;
        RECT 388.950 22.950 391.050 25.050 ;
        RECT 392.250 23.250 393.750 24.150 ;
        RECT 394.950 22.950 397.050 25.050 ;
        RECT 398.400 22.050 399.450 37.950 ;
        RECT 404.400 28.050 405.450 37.950 ;
        RECT 407.400 36.450 408.450 46.950 ;
        RECT 443.400 37.050 444.450 106.950 ;
        RECT 445.950 101.400 448.050 103.500 ;
        RECT 446.250 89.400 447.450 101.400 ;
        RECT 448.950 98.250 451.050 99.150 ;
        RECT 448.950 96.450 451.050 97.050 ;
        RECT 452.400 96.450 453.450 118.950 ;
        RECT 455.400 100.050 456.450 118.950 ;
        RECT 461.400 118.050 462.450 124.950 ;
        RECT 463.950 121.950 466.050 124.050 ;
        RECT 467.250 122.250 468.750 123.150 ;
        RECT 469.950 121.950 472.050 124.050 ;
        RECT 472.950 122.250 475.050 123.150 ;
        RECT 475.950 122.850 478.050 123.750 ;
        RECT 464.400 121.050 465.450 121.950 ;
        RECT 463.950 118.950 466.050 121.050 ;
        RECT 466.950 118.950 469.050 121.050 ;
        RECT 467.400 118.050 468.450 118.950 ;
        RECT 470.400 118.050 471.450 121.950 ;
        RECT 472.950 118.950 475.050 121.050 ;
        RECT 479.400 118.050 480.450 125.400 ;
        RECT 481.950 125.250 483.750 126.150 ;
        RECT 484.950 124.950 487.050 127.050 ;
        RECT 488.250 125.250 489.750 126.150 ;
        RECT 490.950 124.950 493.050 127.050 ;
        RECT 481.950 121.950 484.050 124.050 ;
        RECT 485.250 122.850 486.750 123.750 ;
        RECT 487.950 121.950 490.050 124.050 ;
        RECT 460.950 115.950 463.050 118.050 ;
        RECT 466.950 115.950 469.050 118.050 ;
        RECT 469.950 115.950 472.050 118.050 ;
        RECT 478.950 115.950 481.050 118.050 ;
        RECT 460.950 112.950 463.050 115.050 ;
        RECT 454.950 97.950 457.050 100.050 ;
        RECT 455.400 97.050 456.450 97.950 ;
        RECT 461.400 97.050 462.450 112.950 ;
        RECT 467.400 99.450 468.450 115.950 ;
        RECT 482.400 100.050 483.450 121.950 ;
        RECT 491.400 100.050 492.450 124.950 ;
        RECT 469.950 99.450 472.050 100.050 ;
        RECT 467.400 98.400 472.050 99.450 ;
        RECT 469.950 97.950 472.050 98.400 ;
        RECT 478.950 97.950 481.050 100.050 ;
        RECT 481.950 97.950 484.050 100.050 ;
        RECT 484.950 97.950 487.050 100.050 ;
        RECT 490.950 97.950 493.050 100.050 ;
        RECT 448.950 95.400 453.450 96.450 ;
        RECT 448.950 94.950 451.050 95.400 ;
        RECT 454.950 94.950 457.050 97.050 ;
        RECT 458.250 95.250 459.750 96.150 ;
        RECT 460.950 94.950 463.050 97.050 ;
        RECT 469.950 95.850 472.050 96.750 ;
        RECT 472.950 95.250 475.050 96.150 ;
        RECT 475.950 94.950 478.050 97.050 ;
        RECT 478.950 95.850 481.050 96.750 ;
        RECT 481.950 95.250 484.050 96.150 ;
        RECT 454.950 92.850 456.750 93.750 ;
        RECT 457.950 91.950 460.050 94.050 ;
        RECT 461.250 92.850 462.750 93.750 ;
        RECT 463.950 91.950 466.050 94.050 ;
        RECT 472.950 91.950 475.050 94.050 ;
        RECT 458.400 91.050 459.450 91.950 ;
        RECT 445.950 87.300 448.050 89.400 ;
        RECT 457.950 88.950 460.050 91.050 ;
        RECT 463.950 89.850 466.050 90.750 ;
        RECT 446.250 83.700 447.450 87.300 ;
        RECT 445.950 81.600 448.050 83.700 ;
        RECT 445.950 56.250 448.050 57.150 ;
        RECT 451.950 55.950 454.050 58.050 ;
        RECT 452.400 55.050 453.450 55.950 ;
        RECT 445.950 52.950 448.050 55.050 ;
        RECT 449.250 53.250 450.750 54.150 ;
        RECT 451.950 52.950 454.050 55.050 ;
        RECT 455.250 53.250 457.050 54.150 ;
        RECT 446.400 46.050 447.450 52.950 ;
        RECT 448.950 49.950 451.050 52.050 ;
        RECT 452.250 50.850 453.750 51.750 ;
        RECT 454.950 49.950 457.050 52.050 ;
        RECT 445.950 43.950 448.050 46.050 ;
        RECT 407.400 35.400 411.450 36.450 ;
        RECT 403.950 25.950 406.050 28.050 ;
        RECT 403.950 23.850 406.050 24.750 ;
        RECT 406.950 23.250 409.050 24.150 ;
        RECT 340.950 20.850 342.750 21.750 ;
        RECT 343.950 19.950 346.050 22.050 ;
        RECT 347.250 20.850 348.750 21.750 ;
        RECT 349.950 19.950 352.050 22.050 ;
        RECT 353.250 20.850 355.050 21.750 ;
        RECT 358.950 20.850 360.750 21.750 ;
        RECT 361.950 19.950 364.050 22.050 ;
        RECT 365.250 20.850 366.750 21.750 ;
        RECT 367.950 21.450 370.050 22.050 ;
        RECT 367.950 20.400 372.450 21.450 ;
        RECT 376.950 20.850 378.750 21.750 ;
        RECT 367.950 19.950 370.050 20.400 ;
        RECT 304.950 17.400 309.450 18.450 ;
        RECT 325.950 17.850 327.750 18.750 ;
        RECT 304.950 16.950 307.050 17.400 ;
        RECT 298.950 13.950 301.050 16.050 ;
        RECT 308.400 13.050 309.450 17.400 ;
        RECT 328.950 16.950 331.050 19.050 ;
        RECT 332.250 17.850 333.750 18.750 ;
        RECT 334.950 16.950 337.050 19.050 ;
        RECT 337.950 16.950 340.050 19.050 ;
        RECT 335.400 16.050 336.450 16.950 ;
        RECT 328.950 14.850 331.050 15.750 ;
        RECT 334.950 13.950 337.050 16.050 ;
        RECT 344.400 13.050 345.450 19.950 ;
        RECT 367.950 17.850 370.050 18.750 ;
        RECT 371.400 16.050 372.450 20.400 ;
        RECT 379.950 19.950 382.050 22.050 ;
        RECT 385.950 19.950 388.050 22.050 ;
        RECT 388.950 20.850 390.750 21.750 ;
        RECT 391.950 19.950 394.050 22.050 ;
        RECT 395.250 20.850 396.750 21.750 ;
        RECT 397.950 19.950 400.050 22.050 ;
        RECT 406.950 19.950 409.050 22.050 ;
        RECT 380.400 19.050 381.450 19.950 ;
        RECT 392.400 19.050 393.450 19.950 ;
        RECT 379.950 16.950 382.050 19.050 ;
        RECT 391.950 16.950 394.050 19.050 ;
        RECT 397.950 17.850 400.050 18.750 ;
        RECT 370.950 13.950 373.050 16.050 ;
        RECT 410.400 13.050 411.450 35.400 ;
        RECT 442.950 34.950 445.050 37.050 ;
        RECT 415.950 28.950 418.050 31.050 ;
        RECT 442.950 29.400 445.050 31.500 ;
        RECT 416.400 25.050 417.450 28.950 ;
        RECT 427.950 25.950 430.050 28.050 ;
        RECT 415.950 22.950 418.050 25.050 ;
        RECT 427.950 23.850 430.050 24.750 ;
        RECT 430.950 23.250 433.050 24.150 ;
        RECT 412.950 19.950 415.050 22.050 ;
        RECT 416.400 19.050 417.450 22.950 ;
        RECT 418.950 19.950 421.050 22.050 ;
        RECT 422.250 20.250 424.050 21.150 ;
        RECT 430.950 19.950 433.050 22.050 ;
        RECT 412.950 17.850 414.750 18.750 ;
        RECT 415.950 16.950 418.050 19.050 ;
        RECT 419.250 17.850 420.750 18.750 ;
        RECT 421.950 16.950 424.050 19.050 ;
        RECT 415.950 14.850 418.050 15.750 ;
        RECT 422.400 13.050 423.450 16.950 ;
        RECT 274.950 10.950 277.050 13.050 ;
        RECT 286.950 10.950 289.050 13.050 ;
        RECT 307.950 10.950 310.050 13.050 ;
        RECT 343.950 10.950 346.050 13.050 ;
        RECT 409.950 10.950 412.050 13.050 ;
        RECT 421.950 10.950 424.050 13.050 ;
        RECT 443.400 12.600 444.600 29.400 ;
        RECT 449.400 25.050 450.450 49.950 ;
        RECT 451.950 34.950 454.050 37.050 ;
        RECT 452.400 27.450 453.450 34.950 ;
        RECT 455.400 31.050 456.450 49.950 ;
        RECT 458.400 49.050 459.450 88.950 ;
        RECT 476.400 88.050 477.450 94.950 ;
        RECT 481.950 91.950 484.050 94.050 ;
        RECT 482.400 88.050 483.450 91.950 ;
        RECT 485.400 91.050 486.450 97.950 ;
        RECT 494.400 97.050 495.450 205.950 ;
        RECT 497.400 189.600 498.600 206.400 ;
        RECT 496.950 187.500 499.050 189.600 ;
        RECT 500.400 172.050 501.450 229.950 ;
        RECT 503.400 229.050 504.450 241.950 ;
        RECT 506.400 241.050 507.450 265.950 ;
        RECT 521.400 259.050 522.450 382.950 ;
        RECT 523.950 380.850 526.050 381.750 ;
        RECT 530.400 355.050 531.450 391.950 ;
        RECT 532.950 384.450 535.050 385.050 ;
        RECT 536.400 384.450 537.450 469.950 ;
        RECT 544.950 463.950 547.050 466.050 ;
        RECT 545.400 457.050 546.450 463.950 ;
        RECT 551.400 460.050 552.450 484.950 ;
        RECT 557.400 466.050 558.450 488.400 ;
        RECT 559.950 487.950 562.050 488.400 ;
        RECT 563.250 488.250 564.750 489.150 ;
        RECT 565.950 487.950 568.050 490.050 ;
        RECT 580.950 487.950 583.050 490.050 ;
        RECT 559.950 485.850 561.750 486.750 ;
        RECT 562.950 484.950 565.050 487.050 ;
        RECT 566.250 485.850 568.050 486.750 ;
        RECT 571.950 485.250 574.050 486.150 ;
        RECT 577.950 485.250 580.050 486.150 ;
        RECT 563.400 484.050 564.450 484.950 ;
        RECT 562.950 481.950 565.050 484.050 ;
        RECT 571.950 481.950 574.050 484.050 ;
        RECT 572.400 475.050 573.450 481.950 ;
        RECT 571.950 472.950 574.050 475.050 ;
        RECT 574.950 472.950 577.050 475.050 ;
        RECT 556.950 463.950 559.050 466.050 ;
        RECT 553.950 461.400 556.050 463.500 ;
        RECT 557.400 463.050 558.450 463.950 ;
        RECT 550.950 457.950 553.050 460.050 ;
        RECT 538.950 456.450 541.050 457.050 ;
        RECT 538.950 455.400 543.450 456.450 ;
        RECT 538.950 454.950 541.050 455.400 ;
        RECT 542.400 454.050 543.450 455.400 ;
        RECT 544.950 454.950 547.050 457.050 ;
        RECT 550.950 454.950 553.050 457.050 ;
        RECT 538.950 452.850 541.050 453.750 ;
        RECT 541.950 451.950 544.050 454.050 ;
        RECT 544.950 452.850 547.050 453.750 ;
        RECT 547.950 448.950 550.050 451.050 ;
        RECT 544.950 430.950 547.050 433.050 ;
        RECT 541.950 422.400 544.050 424.500 ;
        RECT 538.950 415.950 541.050 418.050 ;
        RECT 539.400 412.050 540.450 415.950 ;
        RECT 538.950 409.950 541.050 412.050 ;
        RECT 542.400 405.600 543.600 422.400 ;
        RECT 541.950 403.500 544.050 405.600 ;
        RECT 541.950 394.950 544.050 397.050 ;
        RECT 532.950 383.400 537.450 384.450 ;
        RECT 532.950 382.950 535.050 383.400 ;
        RECT 532.950 380.850 535.050 381.750 ;
        RECT 536.400 376.050 537.450 383.400 ;
        RECT 538.950 382.950 541.050 385.050 ;
        RECT 538.950 380.850 541.050 381.750 ;
        RECT 532.950 373.950 535.050 376.050 ;
        RECT 535.950 373.950 538.050 376.050 ;
        RECT 529.950 352.950 532.050 355.050 ;
        RECT 523.950 344.250 526.050 345.150 ;
        RECT 530.400 343.050 531.450 352.950 ;
        RECT 533.400 346.050 534.450 373.950 ;
        RECT 535.950 352.950 538.050 355.050 ;
        RECT 532.950 343.950 535.050 346.050 ;
        RECT 523.950 340.950 526.050 343.050 ;
        RECT 527.250 341.250 528.750 342.150 ;
        RECT 529.950 340.950 532.050 343.050 ;
        RECT 533.250 341.250 535.050 342.150 ;
        RECT 526.950 337.950 529.050 340.050 ;
        RECT 530.250 338.850 531.750 339.750 ;
        RECT 532.950 339.450 535.050 340.050 ;
        RECT 536.400 339.450 537.450 352.950 ;
        RECT 542.400 343.050 543.450 394.950 ;
        RECT 545.400 349.050 546.450 430.950 ;
        RECT 548.400 418.050 549.450 448.950 ;
        RECT 551.400 430.050 552.450 454.950 ;
        RECT 554.250 449.400 555.450 461.400 ;
        RECT 556.950 460.950 559.050 463.050 ;
        RECT 565.950 460.950 568.050 463.050 ;
        RECT 566.400 460.050 567.450 460.950 ;
        RECT 556.950 458.250 559.050 459.150 ;
        RECT 565.950 457.950 568.050 460.050 ;
        RECT 556.950 454.950 559.050 457.050 ;
        RECT 562.950 454.950 565.050 457.050 ;
        RECT 566.250 455.850 567.750 456.750 ;
        RECT 568.950 454.950 571.050 457.050 ;
        RECT 557.400 451.050 558.450 454.950 ;
        RECT 562.950 452.850 565.050 453.750 ;
        RECT 565.950 451.950 568.050 454.050 ;
        RECT 568.950 452.850 571.050 453.750 ;
        RECT 571.950 451.950 574.050 454.050 ;
        RECT 553.950 447.300 556.050 449.400 ;
        RECT 556.950 448.950 559.050 451.050 ;
        RECT 554.250 443.700 555.450 447.300 ;
        RECT 556.950 445.950 559.050 448.050 ;
        RECT 553.950 441.600 556.050 443.700 ;
        RECT 550.950 427.950 553.050 430.050 ;
        RECT 547.950 415.950 550.050 418.050 ;
        RECT 547.950 413.250 550.050 414.150 ;
        RECT 547.950 409.950 550.050 412.050 ;
        RECT 551.400 411.450 552.450 427.950 ;
        RECT 553.950 413.250 556.050 414.150 ;
        RECT 553.950 411.450 556.050 412.050 ;
        RECT 551.400 410.400 556.050 411.450 ;
        RECT 553.950 409.950 556.050 410.400 ;
        RECT 547.950 389.400 550.050 391.500 ;
        RECT 548.400 372.600 549.600 389.400 ;
        RECT 550.950 388.950 553.050 391.050 ;
        RECT 547.950 370.500 550.050 372.600 ;
        RECT 551.400 355.050 552.450 388.950 ;
        RECT 553.950 382.950 556.050 385.050 ;
        RECT 553.950 380.850 556.050 381.750 ;
        RECT 550.950 352.950 553.050 355.050 ;
        RECT 553.950 352.950 556.050 355.050 ;
        RECT 544.950 346.950 547.050 349.050 ;
        RECT 547.950 346.950 550.050 349.050 ;
        RECT 548.400 343.050 549.450 346.950 ;
        RECT 538.950 341.250 541.050 342.150 ;
        RECT 541.950 340.950 544.050 343.050 ;
        RECT 544.950 341.250 547.050 342.150 ;
        RECT 547.950 340.950 550.050 343.050 ;
        RECT 550.950 341.250 553.050 342.150 ;
        RECT 532.950 338.400 537.450 339.450 ;
        RECT 532.950 337.950 535.050 338.400 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 524.400 313.050 525.450 334.950 ;
        RECT 526.950 331.950 529.050 334.050 ;
        RECT 523.950 310.950 526.050 313.050 ;
        RECT 523.950 308.850 526.050 309.750 ;
        RECT 527.400 274.050 528.450 331.950 ;
        RECT 536.400 328.050 537.450 338.400 ;
        RECT 538.950 337.950 541.050 340.050 ;
        RECT 542.250 338.250 543.750 339.150 ;
        RECT 544.950 337.950 547.050 340.050 ;
        RECT 547.950 338.250 549.750 339.150 ;
        RECT 550.950 337.950 553.050 340.050 ;
        RECT 539.400 337.050 540.450 337.950 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 538.950 328.950 541.050 331.050 ;
        RECT 535.950 325.950 538.050 328.050 ;
        RECT 529.950 316.950 532.050 319.050 ;
        RECT 532.950 317.400 535.050 319.500 ;
        RECT 530.400 313.050 531.450 316.950 ;
        RECT 529.950 310.950 532.050 313.050 ;
        RECT 533.250 305.400 534.450 317.400 ;
        RECT 535.950 314.250 538.050 315.150 ;
        RECT 535.950 310.950 538.050 313.050 ;
        RECT 532.950 303.300 535.050 305.400 ;
        RECT 533.250 299.700 534.450 303.300 ;
        RECT 532.950 297.600 535.050 299.700 ;
        RECT 529.950 279.300 532.050 281.400 ;
        RECT 530.550 275.700 531.750 279.300 ;
        RECT 532.950 277.950 535.050 280.050 ;
        RECT 526.950 271.950 529.050 274.050 ;
        RECT 529.950 273.600 532.050 275.700 ;
        RECT 527.400 268.050 528.450 271.950 ;
        RECT 526.950 265.950 529.050 268.050 ;
        RECT 526.950 263.850 529.050 264.750 ;
        RECT 530.550 261.600 531.750 273.600 ;
        RECT 529.950 259.500 532.050 261.600 ;
        RECT 520.950 256.950 523.050 259.050 ;
        RECT 523.950 245.400 526.050 247.500 ;
        RECT 508.950 241.950 511.050 244.050 ;
        RECT 509.400 241.050 510.450 241.950 ;
        RECT 505.950 238.950 508.050 241.050 ;
        RECT 508.950 238.950 511.050 241.050 ;
        RECT 512.250 239.250 513.750 240.150 ;
        RECT 514.950 238.950 517.050 241.050 ;
        RECT 520.950 238.950 523.050 241.050 ;
        RECT 505.950 235.950 508.050 238.050 ;
        RECT 509.250 236.850 510.750 237.750 ;
        RECT 511.950 235.950 514.050 238.050 ;
        RECT 515.250 236.850 517.050 237.750 ;
        RECT 512.400 235.050 513.450 235.950 ;
        RECT 505.950 233.850 508.050 234.750 ;
        RECT 511.950 232.950 514.050 235.050 ;
        RECT 521.400 232.050 522.450 238.950 ;
        RECT 520.950 229.950 523.050 232.050 ;
        RECT 502.950 226.950 505.050 229.050 ;
        RECT 505.950 226.950 508.050 229.050 ;
        RECT 524.400 228.600 525.600 245.400 ;
        RECT 526.950 244.950 529.050 247.050 ;
        RECT 502.950 197.250 505.050 198.150 ;
        RECT 502.950 193.950 505.050 196.050 ;
        RECT 503.400 187.050 504.450 193.950 ;
        RECT 502.950 184.950 505.050 187.050 ;
        RECT 506.400 183.450 507.450 226.950 ;
        RECT 523.950 226.500 526.050 228.600 ;
        RECT 517.950 207.300 520.050 209.400 ;
        RECT 518.250 203.700 519.450 207.300 ;
        RECT 517.950 201.600 520.050 203.700 ;
        RECT 508.950 197.250 511.050 198.150 ;
        RECT 508.950 193.950 511.050 196.050 ;
        RECT 509.400 193.050 510.450 193.950 ;
        RECT 508.950 190.950 511.050 193.050 ;
        RECT 509.400 187.050 510.450 190.950 ;
        RECT 518.250 189.600 519.450 201.600 ;
        RECT 520.950 193.950 523.050 196.050 ;
        RECT 520.950 191.850 523.050 192.750 ;
        RECT 517.950 187.500 520.050 189.600 ;
        RECT 508.950 184.950 511.050 187.050 ;
        RECT 503.400 182.400 507.450 183.450 ;
        RECT 499.950 169.950 502.050 172.050 ;
        RECT 500.400 169.050 501.450 169.950 ;
        RECT 499.950 166.950 502.050 169.050 ;
        RECT 499.950 164.850 502.050 165.750 ;
        RECT 503.400 162.450 504.450 182.400 ;
        RECT 517.950 181.950 520.050 184.050 ;
        RECT 505.950 178.950 508.050 181.050 ;
        RECT 506.400 178.050 507.450 178.950 ;
        RECT 505.950 175.950 508.050 178.050 ;
        RECT 506.400 169.050 507.450 175.950 ;
        RECT 505.950 168.450 508.050 169.050 ;
        RECT 508.950 168.450 511.050 169.050 ;
        RECT 505.950 167.400 511.050 168.450 ;
        RECT 505.950 166.950 508.050 167.400 ;
        RECT 508.950 166.950 511.050 167.400 ;
        RECT 514.950 168.450 517.050 169.050 ;
        RECT 518.400 168.450 519.450 181.950 ;
        RECT 520.950 172.950 523.050 175.050 ;
        RECT 514.950 167.400 519.450 168.450 ;
        RECT 514.950 166.950 517.050 167.400 ;
        RECT 505.950 164.850 508.050 165.750 ;
        RECT 508.950 164.850 511.050 165.750 ;
        RECT 514.950 164.850 517.050 165.750 ;
        RECT 503.400 161.400 507.450 162.450 ;
        RECT 496.950 127.950 499.050 130.050 ;
        RECT 500.250 128.250 501.750 129.150 ;
        RECT 502.950 127.950 505.050 130.050 ;
        RECT 506.400 127.050 507.450 161.400 ;
        RECT 514.950 135.300 517.050 137.400 ;
        RECT 515.550 131.700 516.750 135.300 ;
        RECT 508.950 127.950 511.050 130.050 ;
        RECT 514.950 129.600 517.050 131.700 ;
        RECT 496.950 125.850 498.750 126.750 ;
        RECT 499.950 124.950 502.050 127.050 ;
        RECT 503.250 125.850 505.050 126.750 ;
        RECT 505.950 124.950 508.050 127.050 ;
        RECT 509.400 115.050 510.450 127.950 ;
        RECT 511.950 121.950 514.050 124.050 ;
        RECT 511.950 119.850 514.050 120.750 ;
        RECT 515.550 117.600 516.750 129.600 ;
        RECT 514.950 115.500 517.050 117.600 ;
        RECT 499.950 112.950 502.050 115.050 ;
        RECT 508.950 112.950 511.050 115.050 ;
        RECT 487.950 94.950 490.050 97.050 ;
        RECT 493.950 94.950 496.050 97.050 ;
        RECT 488.400 94.050 489.450 94.950 ;
        RECT 487.950 91.950 490.050 94.050 ;
        RECT 490.950 91.950 493.050 94.050 ;
        RECT 493.950 91.950 496.050 94.050 ;
        RECT 497.250 92.250 499.050 93.150 ;
        RECT 491.400 91.050 492.450 91.950 ;
        RECT 484.950 88.950 487.050 91.050 ;
        RECT 487.950 89.850 489.750 90.750 ;
        RECT 490.950 88.950 493.050 91.050 ;
        RECT 494.250 89.850 495.750 90.750 ;
        RECT 496.950 90.450 499.050 91.050 ;
        RECT 500.400 90.450 501.450 112.950 ;
        RECT 502.950 100.950 505.050 103.050 ;
        RECT 496.950 89.400 501.450 90.450 ;
        RECT 496.950 88.950 499.050 89.400 ;
        RECT 475.950 85.950 478.050 88.050 ;
        RECT 481.950 85.950 484.050 88.050 ;
        RECT 490.950 86.850 493.050 87.750 ;
        RECT 503.400 58.050 504.450 100.950 ;
        RECT 518.400 100.050 519.450 167.400 ;
        RECT 521.400 124.050 522.450 172.950 ;
        RECT 523.950 167.250 526.050 168.150 ;
        RECT 523.950 125.250 526.050 126.150 ;
        RECT 520.950 121.950 523.050 124.050 ;
        RECT 523.950 121.950 526.050 124.050 ;
        RECT 524.400 121.050 525.450 121.950 ;
        RECT 523.950 118.950 526.050 121.050 ;
        RECT 524.400 109.050 525.450 118.950 ;
        RECT 523.950 106.950 526.050 109.050 ;
        RECT 527.400 103.050 528.450 244.950 ;
        RECT 529.950 241.950 532.050 244.050 ;
        RECT 530.400 241.050 531.450 241.950 ;
        RECT 529.950 238.950 532.050 241.050 ;
        RECT 533.400 240.450 534.450 277.950 ;
        RECT 539.400 273.450 540.450 328.950 ;
        RECT 542.400 316.050 543.450 334.950 ;
        RECT 550.950 319.950 553.050 322.050 ;
        RECT 541.950 313.950 544.050 316.050 ;
        RECT 541.950 310.950 544.050 313.050 ;
        RECT 545.250 311.250 546.750 312.150 ;
        RECT 547.950 310.950 550.050 313.050 ;
        RECT 551.400 310.050 552.450 319.950 ;
        RECT 541.950 308.850 543.750 309.750 ;
        RECT 544.950 307.950 547.050 310.050 ;
        RECT 548.250 308.850 549.750 309.750 ;
        RECT 550.950 307.950 553.050 310.050 ;
        RECT 545.400 301.050 546.450 307.950 ;
        RECT 550.950 305.850 553.050 306.750 ;
        RECT 544.950 298.950 547.050 301.050 ;
        RECT 541.950 289.950 544.050 292.050 ;
        RECT 536.400 272.400 540.450 273.450 ;
        RECT 536.400 267.450 537.450 272.400 ;
        RECT 538.950 269.250 541.050 270.150 ;
        RECT 538.950 267.450 541.050 268.050 ;
        RECT 536.400 266.400 541.050 267.450 ;
        RECT 538.950 265.950 541.050 266.400 ;
        RECT 535.950 262.950 538.050 265.050 ;
        RECT 542.400 264.450 543.450 289.950 ;
        RECT 547.950 277.950 550.050 280.050 ;
        RECT 550.950 278.400 553.050 280.500 ;
        RECT 544.950 269.250 547.050 270.150 ;
        RECT 544.950 265.950 547.050 268.050 ;
        RECT 539.400 263.400 543.450 264.450 ;
        RECT 536.400 259.050 537.450 262.950 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 536.400 244.050 537.450 256.950 ;
        RECT 535.950 241.950 538.050 244.050 ;
        RECT 535.950 240.450 538.050 241.050 ;
        RECT 533.400 239.400 538.050 240.450 ;
        RECT 535.950 238.950 538.050 239.400 ;
        RECT 529.950 236.850 532.050 237.750 ;
        RECT 535.950 236.850 538.050 237.750 ;
        RECT 535.950 232.950 538.050 235.050 ;
        RECT 529.950 196.950 532.050 199.050 ;
        RECT 529.950 194.850 532.050 195.750 ;
        RECT 532.950 194.250 535.050 195.150 ;
        RECT 532.950 190.950 535.050 193.050 ;
        RECT 536.400 169.050 537.450 232.950 ;
        RECT 539.400 220.050 540.450 263.400 ;
        RECT 545.400 262.050 546.450 265.950 ;
        RECT 544.950 259.950 547.050 262.050 ;
        RECT 541.950 250.950 544.050 253.050 ;
        RECT 542.400 226.050 543.450 250.950 ;
        RECT 544.950 245.400 547.050 247.500 ;
        RECT 548.400 247.050 549.450 277.950 ;
        RECT 551.400 261.600 552.600 278.400 ;
        RECT 550.950 259.500 553.050 261.600 ;
        RECT 545.250 233.400 546.450 245.400 ;
        RECT 547.950 244.950 550.050 247.050 ;
        RECT 554.400 244.050 555.450 352.950 ;
        RECT 557.400 349.050 558.450 445.950 ;
        RECT 566.400 439.050 567.450 451.950 ;
        RECT 572.400 445.050 573.450 451.950 ;
        RECT 571.950 442.950 574.050 445.050 ;
        RECT 559.950 436.950 562.050 439.050 ;
        RECT 565.950 436.950 568.050 439.050 ;
        RECT 560.400 406.050 561.450 436.950 ;
        RECT 575.400 433.050 576.450 472.950 ;
        RECT 577.950 466.950 580.050 469.050 ;
        RECT 578.400 457.050 579.450 466.950 ;
        RECT 581.400 457.050 582.450 487.950 ;
        RECT 584.400 460.050 585.450 490.950 ;
        RECT 587.400 490.050 588.450 490.950 ;
        RECT 586.950 487.950 589.050 490.050 ;
        RECT 592.950 489.450 595.050 490.050 ;
        RECT 590.250 488.250 591.750 489.150 ;
        RECT 592.950 488.400 597.450 489.450 ;
        RECT 592.950 487.950 595.050 488.400 ;
        RECT 586.950 485.850 588.750 486.750 ;
        RECT 589.950 484.950 592.050 487.050 ;
        RECT 593.250 485.850 595.050 486.750 ;
        RECT 586.950 469.950 589.050 472.050 ;
        RECT 583.950 457.950 586.050 460.050 ;
        RECT 587.400 457.050 588.450 469.950 ;
        RECT 577.950 454.950 580.050 457.050 ;
        RECT 580.950 454.950 583.050 457.050 ;
        RECT 584.250 455.250 585.750 456.150 ;
        RECT 586.950 454.950 589.050 457.050 ;
        RECT 577.950 451.950 580.050 454.050 ;
        RECT 581.250 452.850 582.750 453.750 ;
        RECT 583.950 451.950 586.050 454.050 ;
        RECT 587.250 452.850 589.050 453.750 ;
        RECT 590.400 453.450 591.450 484.950 ;
        RECT 592.950 481.950 595.050 484.050 ;
        RECT 593.400 457.050 594.450 481.950 ;
        RECT 596.400 478.050 597.450 488.400 ;
        RECT 602.400 487.050 603.450 490.950 ;
        RECT 605.400 490.050 606.450 529.950 ;
        RECT 608.400 529.050 609.450 535.950 ;
        RECT 614.400 529.050 615.450 538.950 ;
        RECT 607.950 526.950 610.050 529.050 ;
        RECT 613.950 526.950 616.050 529.050 ;
        RECT 607.950 524.850 610.050 525.750 ;
        RECT 613.950 524.850 616.050 525.750 ;
        RECT 610.950 496.950 613.050 499.050 ;
        RECT 604.950 487.950 607.050 490.050 ;
        RECT 598.950 485.250 601.050 486.150 ;
        RECT 601.950 484.950 604.050 487.050 ;
        RECT 604.950 485.250 607.050 486.150 ;
        RECT 607.950 485.250 610.050 486.150 ;
        RECT 598.950 481.950 601.050 484.050 ;
        RECT 602.250 482.250 603.750 483.150 ;
        RECT 604.950 481.950 607.050 484.050 ;
        RECT 607.950 481.950 610.050 484.050 ;
        RECT 595.950 475.950 598.050 478.050 ;
        RECT 596.400 463.050 597.450 475.950 ;
        RECT 599.400 472.050 600.450 481.950 ;
        RECT 601.950 478.950 604.050 481.050 ;
        RECT 601.950 472.950 604.050 475.050 ;
        RECT 598.950 469.950 601.050 472.050 ;
        RECT 602.400 469.050 603.450 472.950 ;
        RECT 598.950 466.950 601.050 469.050 ;
        RECT 601.950 466.950 604.050 469.050 ;
        RECT 595.950 460.950 598.050 463.050 ;
        RECT 599.400 459.450 600.450 466.950 ;
        RECT 605.400 463.050 606.450 481.950 ;
        RECT 608.400 475.050 609.450 481.950 ;
        RECT 607.950 472.950 610.050 475.050 ;
        RECT 611.400 469.050 612.450 496.950 ;
        RECT 613.950 485.250 616.050 486.150 ;
        RECT 617.400 481.050 618.450 547.950 ;
        RECT 623.400 544.050 624.450 550.950 ;
        RECT 626.400 547.050 627.450 553.950 ;
        RECT 628.950 550.950 631.050 553.050 ;
        RECT 631.950 550.950 634.050 553.050 ;
        RECT 625.950 544.950 628.050 547.050 ;
        RECT 622.950 541.950 625.050 544.050 ;
        RECT 619.950 533.400 622.050 535.500 ;
        RECT 620.400 516.600 621.600 533.400 ;
        RECT 622.950 532.950 625.050 535.050 ;
        RECT 619.950 514.500 622.050 516.600 ;
        RECT 623.400 514.050 624.450 532.950 ;
        RECT 622.950 511.950 625.050 514.050 ;
        RECT 622.950 486.450 625.050 487.050 ;
        RECT 620.400 485.400 625.050 486.450 ;
        RECT 616.950 478.950 619.050 481.050 ;
        RECT 610.950 466.950 613.050 469.050 ;
        RECT 616.950 463.950 619.050 466.050 ;
        RECT 601.950 460.950 604.050 463.050 ;
        RECT 604.950 460.950 607.050 463.050 ;
        RECT 596.400 458.400 600.450 459.450 ;
        RECT 596.400 457.050 597.450 458.400 ;
        RECT 602.400 457.050 603.450 460.950 ;
        RECT 605.400 457.050 606.450 460.950 ;
        RECT 613.950 457.950 616.050 460.050 ;
        RECT 592.950 454.950 595.050 457.050 ;
        RECT 595.950 454.950 598.050 457.050 ;
        RECT 599.250 455.250 600.750 456.150 ;
        RECT 601.950 454.950 604.050 457.050 ;
        RECT 604.950 454.950 607.050 457.050 ;
        RECT 608.250 455.250 609.750 456.150 ;
        RECT 610.950 454.950 613.050 457.050 ;
        RECT 614.400 454.050 615.450 457.950 ;
        RECT 617.400 454.050 618.450 463.950 ;
        RECT 620.400 463.050 621.450 485.400 ;
        RECT 622.950 484.950 625.050 485.400 ;
        RECT 629.400 484.050 630.450 550.950 ;
        RECT 632.400 550.050 633.450 550.950 ;
        RECT 631.950 547.950 634.050 550.050 ;
        RECT 641.400 544.050 642.450 556.950 ;
        RECT 644.400 555.450 645.450 577.950 ;
        RECT 647.400 577.050 648.450 595.950 ;
        RECT 646.950 574.950 649.050 577.050 ;
        RECT 649.950 567.300 652.050 569.400 ;
        RECT 650.550 563.700 651.750 567.300 ;
        RECT 649.950 561.600 652.050 563.700 ;
        RECT 646.950 555.450 649.050 556.050 ;
        RECT 644.400 554.400 649.050 555.450 ;
        RECT 644.400 547.050 645.450 554.400 ;
        RECT 646.950 553.950 649.050 554.400 ;
        RECT 646.950 551.850 649.050 552.750 ;
        RECT 650.550 549.600 651.750 561.600 ;
        RECT 649.950 547.500 652.050 549.600 ;
        RECT 643.950 544.950 646.050 547.050 ;
        RECT 640.950 541.950 643.050 544.050 ;
        RECT 646.950 541.950 649.050 544.050 ;
        RECT 634.950 533.400 637.050 535.500 ;
        RECT 631.950 530.250 634.050 531.150 ;
        RECT 631.950 526.950 634.050 529.050 ;
        RECT 632.400 514.050 633.450 526.950 ;
        RECT 635.550 521.400 636.750 533.400 ;
        RECT 643.950 526.950 646.050 529.050 ;
        RECT 643.950 524.850 646.050 525.750 ;
        RECT 634.950 519.300 637.050 521.400 ;
        RECT 635.550 515.700 636.750 519.300 ;
        RECT 631.950 511.950 634.050 514.050 ;
        RECT 634.950 513.600 637.050 515.700 ;
        RECT 647.400 490.050 648.450 541.950 ;
        RECT 656.400 541.050 657.450 595.950 ;
        RECT 658.950 557.250 661.050 558.150 ;
        RECT 658.950 553.950 661.050 556.050 ;
        RECT 655.950 538.950 658.050 541.050 ;
        RECT 655.950 533.400 658.050 535.500 ;
        RECT 649.950 528.450 652.050 529.050 ;
        RECT 649.950 527.400 654.450 528.450 ;
        RECT 649.950 526.950 652.050 527.400 ;
        RECT 649.950 524.850 652.050 525.750 ;
        RECT 653.400 520.050 654.450 527.400 ;
        RECT 649.950 517.950 652.050 520.050 ;
        RECT 652.950 517.950 655.050 520.050 ;
        RECT 650.400 490.050 651.450 517.950 ;
        RECT 656.400 516.600 657.600 533.400 ;
        RECT 659.400 529.050 660.450 553.950 ;
        RECT 662.400 544.050 663.450 595.950 ;
        RECT 668.550 593.400 669.750 605.400 ;
        RECT 677.400 601.050 678.450 619.950 ;
        RECT 679.950 619.500 682.050 621.600 ;
        RECT 683.400 615.450 684.450 634.950 ;
        RECT 688.950 629.250 691.050 630.150 ;
        RECT 688.950 625.950 691.050 628.050 ;
        RECT 689.400 622.050 690.450 625.950 ;
        RECT 688.950 619.950 691.050 622.050 ;
        RECT 680.400 614.400 684.450 615.450 ;
        RECT 676.950 598.950 679.050 601.050 ;
        RECT 676.950 596.850 679.050 597.750 ;
        RECT 667.950 591.300 670.050 593.400 ;
        RECT 668.550 587.700 669.750 591.300 ;
        RECT 667.950 585.600 670.050 587.700 ;
        RECT 670.950 566.400 673.050 568.500 ;
        RECT 664.950 557.250 667.050 558.150 ;
        RECT 664.950 553.950 667.050 556.050 ;
        RECT 671.400 549.600 672.600 566.400 ;
        RECT 680.400 565.050 681.450 614.400 ;
        RECT 688.950 605.400 691.050 607.500 ;
        RECT 682.950 598.950 685.050 601.050 ;
        RECT 682.950 596.850 685.050 597.750 ;
        RECT 689.400 588.600 690.600 605.400 ;
        RECT 688.950 586.500 691.050 588.600 ;
        RECT 673.950 562.950 676.050 565.050 ;
        RECT 679.950 562.950 682.050 565.050 ;
        RECT 670.950 547.500 673.050 549.600 ;
        RECT 661.950 541.950 664.050 544.050 ;
        RECT 661.950 538.950 664.050 541.050 ;
        RECT 658.950 526.950 661.050 529.050 ;
        RECT 659.400 526.050 660.450 526.950 ;
        RECT 658.950 523.950 661.050 526.050 ;
        RECT 655.950 514.500 658.050 516.600 ;
        RECT 662.400 493.050 663.450 538.950 ;
        RECT 667.950 527.250 670.050 528.150 ;
        RECT 670.950 526.950 673.050 529.050 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 668.400 496.050 669.450 523.950 ;
        RECT 667.950 493.950 670.050 496.050 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 671.400 492.450 672.450 526.950 ;
        RECT 674.400 499.050 675.450 562.950 ;
        RECT 679.950 557.250 682.050 558.150 ;
        RECT 685.950 557.250 688.050 558.150 ;
        RECT 679.950 553.950 682.050 556.050 ;
        RECT 673.950 496.950 676.050 499.050 ;
        RECT 668.400 491.400 672.450 492.450 ;
        RECT 631.950 488.250 634.050 489.150 ;
        RECT 646.950 487.950 649.050 490.050 ;
        RECT 649.950 487.950 652.050 490.050 ;
        RECT 661.950 488.250 664.050 489.150 ;
        RECT 631.950 484.950 634.050 487.050 ;
        RECT 635.250 485.250 636.750 486.150 ;
        RECT 637.950 484.950 640.050 487.050 ;
        RECT 646.950 486.450 649.050 487.050 ;
        RECT 641.250 485.250 643.050 486.150 ;
        RECT 644.400 485.400 649.050 486.450 ;
        RECT 622.950 482.850 625.050 483.750 ;
        RECT 625.950 482.250 628.050 483.150 ;
        RECT 628.950 481.950 631.050 484.050 ;
        RECT 625.950 478.950 628.050 481.050 ;
        RECT 632.400 480.450 633.450 484.950 ;
        RECT 634.950 481.950 637.050 484.050 ;
        RECT 638.250 482.850 639.750 483.750 ;
        RECT 640.950 481.950 643.050 484.050 ;
        RECT 632.400 479.400 636.450 480.450 ;
        RECT 626.400 478.050 627.450 478.950 ;
        RECT 625.950 475.950 628.050 478.050 ;
        RECT 631.950 472.950 634.050 475.050 ;
        RECT 619.950 460.950 622.050 463.050 ;
        RECT 620.400 457.050 621.450 460.950 ;
        RECT 628.950 457.950 631.050 460.050 ;
        RECT 619.950 454.950 622.050 457.050 ;
        RECT 623.250 455.250 624.750 456.150 ;
        RECT 625.950 454.950 628.050 457.050 ;
        RECT 629.400 454.050 630.450 457.950 ;
        RECT 592.950 453.450 595.050 454.050 ;
        RECT 590.400 452.400 595.050 453.450 ;
        RECT 596.250 452.850 597.750 453.750 ;
        RECT 592.950 451.950 595.050 452.400 ;
        RECT 598.950 451.950 601.050 454.050 ;
        RECT 602.250 452.850 604.050 453.750 ;
        RECT 604.950 452.850 606.750 453.750 ;
        RECT 607.950 451.950 610.050 454.050 ;
        RECT 611.250 452.850 612.750 453.750 ;
        RECT 613.950 451.950 616.050 454.050 ;
        RECT 616.950 451.950 619.050 454.050 ;
        RECT 619.950 452.850 621.750 453.750 ;
        RECT 622.950 451.950 625.050 454.050 ;
        RECT 626.250 452.850 627.750 453.750 ;
        RECT 628.950 451.950 631.050 454.050 ;
        RECT 577.950 449.850 580.050 450.750 ;
        RECT 592.950 449.850 595.050 450.750 ;
        RECT 595.950 448.950 598.050 451.050 ;
        RECT 613.950 449.850 616.050 450.750 ;
        RECT 616.950 448.950 619.050 451.050 ;
        RECT 619.950 448.950 622.050 451.050 ;
        RECT 574.950 430.950 577.050 433.050 ;
        RECT 562.950 423.300 565.050 425.400 ;
        RECT 571.950 424.950 574.050 427.050 ;
        RECT 563.250 419.700 564.450 423.300 ;
        RECT 565.950 421.950 568.050 424.050 ;
        RECT 562.950 417.600 565.050 419.700 ;
        RECT 559.950 403.950 562.050 406.050 ;
        RECT 563.250 405.600 564.450 417.600 ;
        RECT 566.400 412.050 567.450 421.950 ;
        RECT 568.950 415.950 571.050 418.050 ;
        RECT 565.950 409.950 568.050 412.050 ;
        RECT 565.950 407.850 568.050 408.750 ;
        RECT 562.950 403.500 565.050 405.600 ;
        RECT 569.400 400.050 570.450 415.950 ;
        RECT 568.950 397.950 571.050 400.050 ;
        RECT 565.950 391.950 568.050 394.050 ;
        RECT 559.950 384.450 562.050 385.050 ;
        RECT 559.950 383.400 564.450 384.450 ;
        RECT 559.950 382.950 562.050 383.400 ;
        RECT 559.950 380.850 562.050 381.750 ;
        RECT 556.950 346.950 559.050 349.050 ;
        RECT 556.950 340.950 559.050 343.050 ;
        RECT 559.950 340.950 562.050 343.050 ;
        RECT 556.950 338.850 559.050 339.750 ;
        RECT 556.950 334.950 559.050 337.050 ;
        RECT 557.400 292.050 558.450 334.950 ;
        RECT 556.950 289.950 559.050 292.050 ;
        RECT 560.400 273.450 561.450 340.950 ;
        RECT 563.400 331.050 564.450 383.400 ;
        RECT 566.400 382.050 567.450 391.950 ;
        RECT 568.950 389.400 571.050 391.500 ;
        RECT 572.400 391.050 573.450 424.950 ;
        RECT 589.950 421.950 592.050 424.050 ;
        RECT 577.950 418.950 580.050 421.050 ;
        RECT 578.400 415.050 579.450 418.950 ;
        RECT 583.950 415.950 586.050 418.050 ;
        RECT 584.400 415.050 585.450 415.950 ;
        RECT 574.950 413.250 576.750 414.150 ;
        RECT 577.950 412.950 580.050 415.050 ;
        RECT 581.250 413.250 582.750 414.150 ;
        RECT 583.950 412.950 586.050 415.050 ;
        RECT 587.250 413.250 589.050 414.150 ;
        RECT 574.950 409.950 577.050 412.050 ;
        RECT 578.250 410.850 579.750 411.750 ;
        RECT 580.950 409.950 583.050 412.050 ;
        RECT 584.250 410.850 585.750 411.750 ;
        RECT 586.950 409.950 589.050 412.050 ;
        RECT 575.400 409.050 576.450 409.950 ;
        RECT 574.950 406.950 577.050 409.050 ;
        RECT 587.400 408.450 588.450 409.950 ;
        RECT 584.400 407.400 588.450 408.450 ;
        RECT 565.950 379.950 568.050 382.050 ;
        RECT 569.250 377.400 570.450 389.400 ;
        RECT 571.950 388.950 574.050 391.050 ;
        RECT 571.950 386.250 574.050 387.150 ;
        RECT 571.950 382.950 574.050 385.050 ;
        RECT 568.950 375.300 571.050 377.400 ;
        RECT 572.400 376.050 573.450 382.950 ;
        RECT 569.250 371.700 570.450 375.300 ;
        RECT 571.950 373.950 574.050 376.050 ;
        RECT 568.950 369.600 571.050 371.700 ;
        RECT 565.950 358.950 568.050 361.050 ;
        RECT 566.400 349.050 567.450 358.950 ;
        RECT 571.950 355.950 574.050 358.050 ;
        RECT 565.950 346.950 568.050 349.050 ;
        RECT 572.400 346.050 573.450 355.950 ;
        RECT 565.950 343.950 568.050 346.050 ;
        RECT 569.250 344.250 570.750 345.150 ;
        RECT 571.950 343.950 574.050 346.050 ;
        RECT 565.950 341.850 567.750 342.750 ;
        RECT 568.950 340.950 571.050 343.050 ;
        RECT 572.250 341.850 574.050 342.750 ;
        RECT 565.950 337.950 568.050 340.050 ;
        RECT 562.950 328.950 565.050 331.050 ;
        RECT 562.950 317.400 565.050 319.500 ;
        RECT 563.400 300.600 564.600 317.400 ;
        RECT 562.950 298.500 565.050 300.600 ;
        RECT 566.400 273.450 567.450 337.950 ;
        RECT 569.400 322.050 570.450 340.950 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 575.400 339.450 576.450 406.950 ;
        RECT 584.400 406.050 585.450 407.400 ;
        RECT 590.400 406.050 591.450 421.950 ;
        RECT 596.400 415.050 597.450 448.950 ;
        RECT 613.950 445.950 616.050 448.050 ;
        RECT 604.950 421.950 607.050 424.050 ;
        RECT 605.400 415.050 606.450 421.950 ;
        RECT 610.950 416.250 613.050 417.150 ;
        RECT 592.950 413.250 595.050 414.150 ;
        RECT 595.950 412.950 598.050 415.050 ;
        RECT 598.950 413.250 601.050 414.150 ;
        RECT 601.950 413.250 603.750 414.150 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 608.250 413.250 609.750 414.150 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 592.950 409.950 595.050 412.050 ;
        RECT 596.250 410.250 597.750 411.150 ;
        RECT 598.950 409.950 601.050 412.050 ;
        RECT 601.950 409.950 604.050 412.050 ;
        RECT 605.250 410.850 606.750 411.750 ;
        RECT 607.950 409.950 610.050 412.050 ;
        RECT 577.950 403.950 580.050 406.050 ;
        RECT 583.950 403.950 586.050 406.050 ;
        RECT 589.950 403.950 592.050 406.050 ;
        RECT 578.400 373.050 579.450 403.950 ;
        RECT 586.950 388.950 589.050 391.050 ;
        RECT 587.400 388.050 588.450 388.950 ;
        RECT 593.400 388.050 594.450 409.950 ;
        RECT 595.950 406.950 598.050 409.050 ;
        RECT 599.400 406.050 600.450 409.950 ;
        RECT 602.400 409.050 603.450 409.950 ;
        RECT 601.950 406.950 604.050 409.050 ;
        RECT 607.950 406.950 610.050 409.050 ;
        RECT 598.950 403.950 601.050 406.050 ;
        RECT 599.400 397.050 600.450 403.950 ;
        RECT 598.950 394.950 601.050 397.050 ;
        RECT 608.400 394.050 609.450 406.950 ;
        RECT 611.400 406.050 612.450 412.950 ;
        RECT 610.950 403.950 613.050 406.050 ;
        RECT 595.950 391.950 598.050 394.050 ;
        RECT 607.950 391.950 610.050 394.050 ;
        RECT 596.400 388.050 597.450 391.950 ;
        RECT 614.400 391.050 615.450 445.950 ;
        RECT 617.400 409.050 618.450 448.950 ;
        RECT 620.400 424.050 621.450 448.950 ;
        RECT 623.400 445.050 624.450 451.950 ;
        RECT 625.950 448.950 628.050 451.050 ;
        RECT 628.950 449.850 631.050 450.750 ;
        RECT 622.950 442.950 625.050 445.050 ;
        RECT 619.950 421.950 622.050 424.050 ;
        RECT 619.950 416.250 622.050 417.150 ;
        RECT 626.400 415.050 627.450 448.950 ;
        RECT 632.400 418.050 633.450 472.950 ;
        RECT 635.400 469.050 636.450 479.400 ;
        RECT 637.950 478.950 640.050 481.050 ;
        RECT 640.950 478.950 643.050 481.050 ;
        RECT 638.400 475.050 639.450 478.950 ;
        RECT 637.950 472.950 640.050 475.050 ;
        RECT 637.950 469.950 640.050 472.050 ;
        RECT 634.950 466.950 637.050 469.050 ;
        RECT 634.950 457.950 637.050 460.050 ;
        RECT 638.400 459.450 639.450 469.950 ;
        RECT 641.400 463.050 642.450 478.950 ;
        RECT 644.400 472.050 645.450 485.400 ;
        RECT 646.950 484.950 649.050 485.400 ;
        RECT 652.950 485.250 654.750 486.150 ;
        RECT 655.950 484.950 658.050 487.050 ;
        RECT 659.250 485.250 660.750 486.150 ;
        RECT 661.950 484.950 664.050 487.050 ;
        RECT 646.950 482.850 649.050 483.750 ;
        RECT 649.950 482.250 652.050 483.150 ;
        RECT 652.950 481.950 655.050 484.050 ;
        RECT 656.250 482.850 657.750 483.750 ;
        RECT 658.950 481.950 661.050 484.050 ;
        RECT 661.950 481.950 664.050 484.050 ;
        RECT 649.950 478.950 652.050 481.050 ;
        RECT 643.950 469.950 646.050 472.050 ;
        RECT 643.950 466.950 646.050 469.050 ;
        RECT 640.950 460.950 643.050 463.050 ;
        RECT 638.400 458.400 642.450 459.450 ;
        RECT 634.950 455.850 637.050 456.750 ;
        RECT 637.950 455.250 640.050 456.150 ;
        RECT 634.950 451.950 637.050 454.050 ;
        RECT 637.950 453.450 640.050 454.050 ;
        RECT 641.400 453.450 642.450 458.400 ;
        RECT 644.400 457.050 645.450 466.950 ;
        RECT 646.950 460.950 649.050 463.050 ;
        RECT 650.400 462.450 651.450 478.950 ;
        RECT 653.400 478.050 654.450 481.950 ;
        RECT 652.950 475.950 655.050 478.050 ;
        RECT 653.400 469.050 654.450 475.950 ;
        RECT 659.400 475.050 660.450 481.950 ;
        RECT 658.950 472.950 661.050 475.050 ;
        RECT 655.950 469.950 658.050 472.050 ;
        RECT 652.950 466.950 655.050 469.050 ;
        RECT 650.400 461.400 654.450 462.450 ;
        RECT 643.950 454.950 646.050 457.050 ;
        RECT 637.950 452.400 642.450 453.450 ;
        RECT 637.950 451.950 640.050 452.400 ;
        RECT 643.950 451.950 646.050 454.050 ;
        RECT 635.400 442.050 636.450 451.950 ;
        RECT 647.400 451.050 648.450 460.950 ;
        RECT 649.950 457.950 652.050 460.050 ;
        RECT 650.400 454.050 651.450 457.950 ;
        RECT 653.400 457.050 654.450 461.400 ;
        RECT 652.950 454.950 655.050 457.050 ;
        RECT 649.950 451.950 652.050 454.050 ;
        RECT 653.250 452.250 655.050 453.150 ;
        RECT 640.950 450.450 643.050 451.050 ;
        RECT 638.400 449.400 643.050 450.450 ;
        RECT 643.950 449.850 645.750 450.750 ;
        RECT 634.950 439.950 637.050 442.050 ;
        RECT 638.400 427.050 639.450 449.400 ;
        RECT 640.950 448.950 643.050 449.400 ;
        RECT 646.950 448.950 649.050 451.050 ;
        RECT 650.250 449.850 651.750 450.750 ;
        RECT 652.950 448.950 655.050 451.050 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 446.850 649.050 447.750 ;
        RECT 641.400 439.050 642.450 445.950 ;
        RECT 640.950 436.950 643.050 439.050 ;
        RECT 640.950 427.950 643.050 430.050 ;
        RECT 637.950 424.950 640.050 427.050 ;
        RECT 631.950 415.950 634.050 418.050 ;
        RECT 619.950 412.950 622.050 415.050 ;
        RECT 623.250 413.250 624.750 414.150 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 629.250 413.250 631.050 414.150 ;
        RECT 631.950 413.250 634.050 414.150 ;
        RECT 637.950 413.250 640.050 414.150 ;
        RECT 622.950 409.950 625.050 412.050 ;
        RECT 626.250 410.850 627.750 411.750 ;
        RECT 628.950 409.950 631.050 412.050 ;
        RECT 631.950 409.950 634.050 412.050 ;
        RECT 635.250 410.250 636.750 411.150 ;
        RECT 637.950 409.950 640.050 412.050 ;
        RECT 616.950 406.950 619.050 409.050 ;
        RECT 616.950 403.950 619.050 406.050 ;
        RECT 601.950 388.950 604.050 391.050 ;
        RECT 613.950 388.950 616.050 391.050 ;
        RECT 586.950 385.950 589.050 388.050 ;
        RECT 592.950 385.950 595.050 388.050 ;
        RECT 595.950 385.950 598.050 388.050 ;
        RECT 580.950 382.950 583.050 385.050 ;
        RECT 584.250 383.250 586.050 384.150 ;
        RECT 586.950 383.850 589.050 384.750 ;
        RECT 589.950 383.250 592.050 384.150 ;
        RECT 592.950 382.950 595.050 385.050 ;
        RECT 596.250 383.850 597.750 384.750 ;
        RECT 598.950 382.950 601.050 385.050 ;
        RECT 580.950 380.850 582.750 381.750 ;
        RECT 583.950 379.950 586.050 382.050 ;
        RECT 589.950 379.950 592.050 382.050 ;
        RECT 592.950 380.850 595.050 381.750 ;
        RECT 595.950 379.950 598.050 382.050 ;
        RECT 598.950 380.850 601.050 381.750 ;
        RECT 590.400 373.050 591.450 379.950 ;
        RECT 577.950 370.950 580.050 373.050 ;
        RECT 589.950 370.950 592.050 373.050 ;
        RECT 592.950 370.950 595.050 373.050 ;
        RECT 580.950 352.950 583.050 355.050 ;
        RECT 581.400 343.050 582.450 352.950 ;
        RECT 590.400 346.050 591.450 370.950 ;
        RECT 593.400 346.050 594.450 370.950 ;
        RECT 596.400 349.050 597.450 379.950 ;
        RECT 602.400 361.050 603.450 388.950 ;
        RECT 610.950 385.950 613.050 388.050 ;
        RECT 604.950 382.950 607.050 385.050 ;
        RECT 607.950 383.250 610.050 384.150 ;
        RECT 605.400 376.050 606.450 382.950 ;
        RECT 604.950 373.950 607.050 376.050 ;
        RECT 611.400 370.050 612.450 385.950 ;
        RECT 613.950 373.950 616.050 376.050 ;
        RECT 610.950 367.950 613.050 370.050 ;
        RECT 607.950 364.950 610.050 367.050 ;
        RECT 601.950 358.950 604.050 361.050 ;
        RECT 598.950 355.950 601.050 358.050 ;
        RECT 595.950 346.950 598.050 349.050 ;
        RECT 589.950 343.950 592.050 346.050 ;
        RECT 592.950 343.950 595.050 346.050 ;
        RECT 599.400 343.050 600.450 355.950 ;
        RECT 608.400 346.050 609.450 364.950 ;
        RECT 607.950 343.950 610.050 346.050 ;
        RECT 577.950 341.250 579.750 342.150 ;
        RECT 580.950 340.950 583.050 343.050 ;
        RECT 584.250 341.250 585.750 342.150 ;
        RECT 586.950 340.950 589.050 343.050 ;
        RECT 590.250 341.250 592.050 342.150 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 595.950 341.250 597.750 342.150 ;
        RECT 598.950 340.950 601.050 343.050 ;
        RECT 602.250 341.250 603.750 342.150 ;
        RECT 604.950 340.950 607.050 343.050 ;
        RECT 608.250 341.250 610.050 342.150 ;
        RECT 577.950 339.450 580.050 340.050 ;
        RECT 575.400 338.400 580.050 339.450 ;
        RECT 581.250 338.850 582.750 339.750 ;
        RECT 577.950 337.950 580.050 338.400 ;
        RECT 583.950 337.950 586.050 340.050 ;
        RECT 587.250 338.850 588.750 339.750 ;
        RECT 589.950 337.950 592.050 340.050 ;
        RECT 572.400 322.050 573.450 337.950 ;
        RECT 578.400 337.050 579.450 337.950 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 584.400 336.450 585.450 337.950 ;
        RECT 589.950 336.450 592.050 337.050 ;
        RECT 584.400 335.400 592.050 336.450 ;
        RECT 589.950 334.950 592.050 335.400 ;
        RECT 574.950 328.950 577.050 331.050 ;
        RECT 568.950 319.950 571.050 322.050 ;
        RECT 571.950 319.950 574.050 322.050 ;
        RECT 575.400 316.050 576.450 328.950 ;
        RECT 589.950 319.950 592.050 322.050 ;
        RECT 583.950 317.400 586.050 319.500 ;
        RECT 571.950 313.950 574.050 316.050 ;
        RECT 574.950 313.950 577.050 316.050 ;
        RECT 568.950 310.950 571.050 313.050 ;
        RECT 568.950 308.850 571.050 309.750 ;
        RECT 572.400 304.050 573.450 313.950 ;
        RECT 575.400 313.050 576.450 313.950 ;
        RECT 574.950 310.950 577.050 313.050 ;
        RECT 580.950 310.950 583.050 313.050 ;
        RECT 574.950 308.850 577.050 309.750 ;
        RECT 568.950 301.950 571.050 304.050 ;
        RECT 571.950 301.950 574.050 304.050 ;
        RECT 557.400 272.400 561.450 273.450 ;
        RECT 563.400 272.400 567.450 273.450 ;
        RECT 553.950 243.450 556.050 244.050 ;
        RECT 547.950 242.250 550.050 243.150 ;
        RECT 551.400 242.400 556.050 243.450 ;
        RECT 557.400 243.450 558.450 272.400 ;
        RECT 559.950 269.250 562.050 270.150 ;
        RECT 559.950 265.950 562.050 268.050 ;
        RECT 560.400 265.050 561.450 265.950 ;
        RECT 563.400 265.050 564.450 272.400 ;
        RECT 565.950 269.250 568.050 270.150 ;
        RECT 565.950 265.950 568.050 268.050 ;
        RECT 559.950 262.950 562.050 265.050 ;
        RECT 562.950 262.950 565.050 265.050 ;
        RECT 569.400 261.450 570.450 301.950 ;
        RECT 571.950 274.950 574.050 277.050 ;
        RECT 572.400 273.450 573.450 274.950 ;
        RECT 581.400 274.050 582.450 310.950 ;
        RECT 584.250 305.400 585.450 317.400 ;
        RECT 586.950 314.250 589.050 315.150 ;
        RECT 586.950 312.450 589.050 313.050 ;
        RECT 590.400 312.450 591.450 319.950 ;
        RECT 586.950 311.400 591.450 312.450 ;
        RECT 586.950 310.950 589.050 311.400 ;
        RECT 586.950 307.950 589.050 310.050 ;
        RECT 583.950 303.300 586.050 305.400 ;
        RECT 584.250 299.700 585.450 303.300 ;
        RECT 583.950 297.600 586.050 299.700 ;
        RECT 583.950 289.950 586.050 292.050 ;
        RECT 574.950 273.450 577.050 274.050 ;
        RECT 572.400 272.400 577.050 273.450 ;
        RECT 572.400 268.050 573.450 272.400 ;
        RECT 574.950 271.950 577.050 272.400 ;
        RECT 578.250 272.250 579.750 273.150 ;
        RECT 580.950 271.950 583.050 274.050 ;
        RECT 574.950 269.850 576.750 270.750 ;
        RECT 577.950 268.950 580.050 271.050 ;
        RECT 581.250 269.850 583.050 270.750 ;
        RECT 571.950 265.950 574.050 268.050 ;
        RECT 580.950 265.950 583.050 268.050 ;
        RECT 571.950 262.950 574.050 265.050 ;
        RECT 566.400 260.400 570.450 261.450 ;
        RECT 566.400 247.050 567.450 260.400 ;
        RECT 568.950 256.950 571.050 259.050 ;
        RECT 569.400 253.050 570.450 256.950 ;
        RECT 568.950 250.950 571.050 253.050 ;
        RECT 565.950 244.950 568.050 247.050 ;
        RECT 569.400 244.050 570.450 250.950 ;
        RECT 557.400 242.400 561.450 243.450 ;
        RECT 547.950 240.450 550.050 241.050 ;
        RECT 551.400 240.450 552.450 242.400 ;
        RECT 553.950 241.950 556.050 242.400 ;
        RECT 547.950 239.400 552.450 240.450 ;
        RECT 553.950 239.850 556.050 240.750 ;
        RECT 547.950 238.950 550.050 239.400 ;
        RECT 556.950 239.250 559.050 240.150 ;
        RECT 556.950 235.950 559.050 238.050 ;
        RECT 544.950 231.300 547.050 233.400 ;
        RECT 557.400 232.050 558.450 235.950 ;
        RECT 545.250 227.700 546.450 231.300 ;
        RECT 556.950 229.950 559.050 232.050 ;
        RECT 541.950 223.950 544.050 226.050 ;
        RECT 544.950 225.600 547.050 227.700 ;
        RECT 538.950 217.950 541.050 220.050 ;
        RECT 542.400 199.050 543.450 223.950 ;
        RECT 547.950 217.950 550.050 220.050 ;
        RECT 538.950 197.250 541.050 198.150 ;
        RECT 541.950 196.950 544.050 199.050 ;
        RECT 544.950 197.250 547.050 198.150 ;
        RECT 538.950 193.950 541.050 196.050 ;
        RECT 542.250 194.250 543.750 195.150 ;
        RECT 544.950 193.950 547.050 196.050 ;
        RECT 538.950 190.950 541.050 193.050 ;
        RECT 541.950 190.950 544.050 193.050 ;
        RECT 544.950 190.950 547.050 193.050 ;
        RECT 539.400 189.450 540.450 190.950 ;
        RECT 545.400 189.450 546.450 190.950 ;
        RECT 539.400 188.400 546.450 189.450 ;
        RECT 541.950 184.950 544.050 187.050 ;
        RECT 535.950 166.950 538.050 169.050 ;
        RECT 538.950 166.950 541.050 169.050 ;
        RECT 535.950 134.400 538.050 136.500 ;
        RECT 529.950 125.250 532.050 126.150 ;
        RECT 529.950 121.950 532.050 124.050 ;
        RECT 536.400 117.600 537.600 134.400 ;
        RECT 539.400 124.050 540.450 166.950 ;
        RECT 542.400 165.450 543.450 184.950 ;
        RECT 544.950 167.250 547.050 168.150 ;
        RECT 544.950 165.450 547.050 166.050 ;
        RECT 542.400 164.400 547.050 165.450 ;
        RECT 544.950 163.950 547.050 164.400 ;
        RECT 545.400 130.050 546.450 163.950 ;
        RECT 548.400 148.050 549.450 217.950 ;
        RECT 560.400 202.050 561.450 242.400 ;
        RECT 562.950 241.950 565.050 244.050 ;
        RECT 568.950 241.950 571.050 244.050 ;
        RECT 563.400 237.450 564.450 241.950 ;
        RECT 565.950 239.250 568.050 240.150 ;
        RECT 568.950 239.850 571.050 240.750 ;
        RECT 565.950 237.450 568.050 238.050 ;
        RECT 563.400 236.400 568.050 237.450 ;
        RECT 565.950 235.950 568.050 236.400 ;
        RECT 568.950 235.950 571.050 238.050 ;
        RECT 565.950 232.950 568.050 235.050 ;
        RECT 559.950 199.950 562.050 202.050 ;
        RECT 550.950 197.250 553.050 198.150 ;
        RECT 556.950 197.250 559.050 198.150 ;
        RECT 562.950 196.950 565.050 199.050 ;
        RECT 550.950 193.950 553.050 196.050 ;
        RECT 554.250 194.250 555.750 195.150 ;
        RECT 556.950 193.950 559.050 196.050 ;
        RECT 559.950 194.250 562.050 195.150 ;
        RECT 562.950 194.850 565.050 195.750 ;
        RECT 551.400 193.050 552.450 193.950 ;
        RECT 550.950 190.950 553.050 193.050 ;
        RECT 553.950 190.950 556.050 193.050 ;
        RECT 557.400 192.450 558.450 193.950 ;
        RECT 559.950 192.450 562.050 193.050 ;
        RECT 557.400 191.400 562.050 192.450 ;
        RECT 559.950 190.950 562.050 191.400 ;
        RECT 553.950 167.250 556.050 168.150 ;
        RECT 547.950 145.950 550.050 148.050 ;
        RECT 562.950 134.400 565.050 136.500 ;
        RECT 544.950 127.950 547.050 130.050 ;
        RECT 556.950 127.950 559.050 130.050 ;
        RECT 544.950 125.250 547.050 126.150 ;
        RECT 550.950 125.250 553.050 126.150 ;
        RECT 538.950 121.950 541.050 124.050 ;
        RECT 544.950 121.950 547.050 124.050 ;
        RECT 550.950 121.950 553.050 124.050 ;
        RECT 535.950 115.500 538.050 117.600 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 544.950 101.400 547.050 103.500 ;
        RECT 551.400 103.050 552.450 121.950 ;
        RECT 557.400 121.050 558.450 127.950 ;
        RECT 556.950 118.950 559.050 121.050 ;
        RECT 508.950 97.950 511.050 100.050 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 523.950 97.950 526.050 100.050 ;
        RECT 535.950 97.950 538.050 100.050 ;
        RECT 505.950 95.250 508.050 96.150 ;
        RECT 508.950 95.850 511.050 96.750 ;
        RECT 511.950 94.950 514.050 97.050 ;
        RECT 505.950 91.950 508.050 94.050 ;
        RECT 512.400 90.450 513.450 94.950 ;
        RECT 514.950 92.250 516.750 93.150 ;
        RECT 517.950 91.950 520.050 94.050 ;
        RECT 521.250 92.250 523.050 93.150 ;
        RECT 514.950 90.450 517.050 91.050 ;
        RECT 512.400 89.400 517.050 90.450 ;
        RECT 518.250 89.850 519.750 90.750 ;
        RECT 520.950 90.450 523.050 91.050 ;
        RECT 524.400 90.450 525.450 97.950 ;
        RECT 536.400 97.050 537.450 97.950 ;
        RECT 529.950 94.950 532.050 97.050 ;
        RECT 533.250 95.250 534.750 96.150 ;
        RECT 535.950 94.950 538.050 97.050 ;
        RECT 526.950 91.950 529.050 94.050 ;
        RECT 530.250 92.850 531.750 93.750 ;
        RECT 532.950 91.950 535.050 94.050 ;
        RECT 536.250 92.850 538.050 93.750 ;
        RECT 514.950 88.950 517.050 89.400 ;
        RECT 520.950 89.400 525.450 90.450 ;
        RECT 526.950 89.850 529.050 90.750 ;
        RECT 520.950 88.950 523.050 89.400 ;
        RECT 521.400 64.050 522.450 88.950 ;
        RECT 545.400 84.600 546.600 101.400 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 557.400 97.050 558.450 118.950 ;
        RECT 563.400 117.600 564.600 134.400 ;
        RECT 562.950 115.500 565.050 117.600 ;
        RECT 566.400 109.050 567.450 232.950 ;
        RECT 569.400 193.050 570.450 235.950 ;
        RECT 572.400 235.050 573.450 262.950 ;
        RECT 581.400 262.050 582.450 265.950 ;
        RECT 580.950 259.950 583.050 262.050 ;
        RECT 577.950 253.950 580.050 256.050 ;
        RECT 574.950 247.950 577.050 250.050 ;
        RECT 575.400 241.050 576.450 247.950 ;
        RECT 578.400 241.050 579.450 253.950 ;
        RECT 584.400 253.050 585.450 289.950 ;
        RECT 587.400 280.050 588.450 307.950 ;
        RECT 586.950 277.950 589.050 280.050 ;
        RECT 593.400 274.050 594.450 340.950 ;
        RECT 595.950 337.950 598.050 340.050 ;
        RECT 599.250 338.850 600.750 339.750 ;
        RECT 601.950 337.950 604.050 340.050 ;
        RECT 605.250 338.850 606.750 339.750 ;
        RECT 607.950 337.950 610.050 340.050 ;
        RECT 596.400 337.050 597.450 337.950 ;
        RECT 595.950 334.950 598.050 337.050 ;
        RECT 598.950 336.450 601.050 337.050 ;
        RECT 608.400 336.450 609.450 337.950 ;
        RECT 598.950 335.400 609.450 336.450 ;
        RECT 598.950 334.950 601.050 335.400 ;
        RECT 601.950 331.950 604.050 334.050 ;
        RECT 604.950 331.950 607.050 334.050 ;
        RECT 598.950 317.400 601.050 319.500 ;
        RECT 595.950 314.250 598.050 315.150 ;
        RECT 595.950 310.950 598.050 313.050 ;
        RECT 599.550 305.400 600.750 317.400 ;
        RECT 598.950 303.300 601.050 305.400 ;
        RECT 599.550 299.700 600.750 303.300 ;
        RECT 598.950 297.600 601.050 299.700 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 586.950 272.250 589.050 273.150 ;
        RECT 592.950 271.950 595.050 274.050 ;
        RECT 586.950 268.950 589.050 271.050 ;
        RECT 590.250 269.250 591.750 270.150 ;
        RECT 592.950 268.950 595.050 271.050 ;
        RECT 596.250 269.250 598.050 270.150 ;
        RECT 586.950 267.450 589.050 268.050 ;
        RECT 589.950 267.450 592.050 268.050 ;
        RECT 586.950 266.400 592.050 267.450 ;
        RECT 593.250 266.850 594.750 267.750 ;
        RECT 586.950 265.950 589.050 266.400 ;
        RECT 589.950 265.950 592.050 266.400 ;
        RECT 595.950 265.950 598.050 268.050 ;
        RECT 599.400 264.450 600.450 292.950 ;
        RECT 602.400 292.050 603.450 331.950 ;
        RECT 605.400 313.050 606.450 331.950 ;
        RECT 607.950 313.950 610.050 316.050 ;
        RECT 608.400 313.050 609.450 313.950 ;
        RECT 604.950 310.950 607.050 313.050 ;
        RECT 607.950 310.950 610.050 313.050 ;
        RECT 607.950 308.850 610.050 309.750 ;
        RECT 607.950 301.950 610.050 304.050 ;
        RECT 601.950 289.950 604.050 292.050 ;
        RECT 601.950 272.250 604.050 273.150 ;
        RECT 608.400 271.050 609.450 301.950 ;
        RECT 611.400 295.050 612.450 367.950 ;
        RECT 614.400 315.450 615.450 373.950 ;
        RECT 617.400 367.050 618.450 403.950 ;
        RECT 623.400 403.050 624.450 409.950 ;
        RECT 629.400 409.050 630.450 409.950 ;
        RECT 625.950 406.950 628.050 409.050 ;
        RECT 628.950 406.950 631.050 409.050 ;
        RECT 622.950 400.950 625.050 403.050 ;
        RECT 619.950 397.950 622.050 400.050 ;
        RECT 616.950 364.950 619.050 367.050 ;
        RECT 616.950 350.400 619.050 352.500 ;
        RECT 620.400 352.050 621.450 397.950 ;
        RECT 622.950 391.950 625.050 394.050 ;
        RECT 617.400 333.600 618.600 350.400 ;
        RECT 619.950 349.950 622.050 352.050 ;
        RECT 623.400 345.450 624.450 391.950 ;
        RECT 620.400 344.400 624.450 345.450 ;
        RECT 616.950 331.500 619.050 333.600 ;
        RECT 620.400 324.450 621.450 344.400 ;
        RECT 622.950 341.250 625.050 342.150 ;
        RECT 622.950 337.950 625.050 340.050 ;
        RECT 623.400 337.050 624.450 337.950 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 620.400 323.400 624.450 324.450 ;
        RECT 619.950 317.400 622.050 319.500 ;
        RECT 614.400 314.400 618.450 315.450 ;
        RECT 613.950 310.950 616.050 313.050 ;
        RECT 613.950 308.850 616.050 309.750 ;
        RECT 610.950 292.950 613.050 295.050 ;
        RECT 617.400 280.050 618.450 314.400 ;
        RECT 620.400 300.600 621.600 317.400 ;
        RECT 619.950 298.500 622.050 300.600 ;
        RECT 623.400 294.450 624.450 323.400 ;
        RECT 620.400 293.400 624.450 294.450 ;
        RECT 616.950 277.950 619.050 280.050 ;
        RECT 601.950 268.950 604.050 271.050 ;
        RECT 605.250 269.250 606.750 270.150 ;
        RECT 607.950 268.950 610.050 271.050 ;
        RECT 611.250 269.250 613.050 270.150 ;
        RECT 616.950 269.250 619.050 270.150 ;
        RECT 596.400 263.400 600.450 264.450 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 583.950 250.950 586.050 253.050 ;
        RECT 583.950 247.950 586.050 250.050 ;
        RECT 584.400 241.050 585.450 247.950 ;
        RECT 589.950 241.950 592.050 244.050 ;
        RECT 593.400 241.050 594.450 256.950 ;
        RECT 574.950 238.950 577.050 241.050 ;
        RECT 577.950 238.950 580.050 241.050 ;
        RECT 583.950 240.450 586.050 241.050 ;
        RECT 586.950 240.450 589.050 241.050 ;
        RECT 581.250 239.250 582.750 240.150 ;
        RECT 583.950 239.400 589.050 240.450 ;
        RECT 590.250 239.850 591.750 240.750 ;
        RECT 583.950 238.950 586.050 239.400 ;
        RECT 586.950 238.950 589.050 239.400 ;
        RECT 592.950 238.950 595.050 241.050 ;
        RECT 574.950 235.950 577.050 238.050 ;
        RECT 578.250 236.850 579.750 237.750 ;
        RECT 580.950 235.950 583.050 238.050 ;
        RECT 584.250 236.850 586.050 237.750 ;
        RECT 586.950 236.850 589.050 237.750 ;
        RECT 592.950 236.850 595.050 237.750 ;
        RECT 571.950 232.950 574.050 235.050 ;
        RECT 574.950 233.850 577.050 234.750 ;
        RECT 596.400 234.450 597.450 263.400 ;
        RECT 598.950 259.950 601.050 262.050 ;
        RECT 599.400 255.450 600.450 259.950 ;
        RECT 602.400 259.050 603.450 268.950 ;
        RECT 604.950 265.950 607.050 268.050 ;
        RECT 608.250 266.850 609.750 267.750 ;
        RECT 610.950 265.950 613.050 268.050 ;
        RECT 613.950 266.250 615.750 267.150 ;
        RECT 616.950 265.950 619.050 268.050 ;
        RECT 604.950 262.950 607.050 265.050 ;
        RECT 607.950 262.950 610.050 265.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 599.400 254.400 603.450 255.450 ;
        RECT 602.400 244.050 603.450 254.400 ;
        RECT 601.950 241.950 604.050 244.050 ;
        RECT 605.400 241.050 606.450 262.950 ;
        RECT 608.400 250.050 609.450 262.950 ;
        RECT 611.400 262.050 612.450 265.950 ;
        RECT 613.950 262.950 616.050 265.050 ;
        RECT 610.950 259.950 613.050 262.050 ;
        RECT 614.400 256.050 615.450 262.950 ;
        RECT 610.950 253.950 613.050 256.050 ;
        RECT 613.950 253.950 616.050 256.050 ;
        RECT 607.950 247.950 610.050 250.050 ;
        RECT 611.400 246.450 612.450 253.950 ;
        RECT 617.400 250.050 618.450 265.950 ;
        RECT 613.950 247.950 616.050 250.050 ;
        RECT 616.950 247.950 619.050 250.050 ;
        RECT 608.400 245.400 612.450 246.450 ;
        RECT 598.950 238.950 601.050 241.050 ;
        RECT 602.250 239.850 603.750 240.750 ;
        RECT 604.950 238.950 607.050 241.050 ;
        RECT 598.950 236.850 601.050 237.750 ;
        RECT 601.950 235.950 604.050 238.050 ;
        RECT 604.950 236.850 607.050 237.750 ;
        RECT 593.400 233.400 597.450 234.450 ;
        RECT 574.950 207.300 577.050 209.400 ;
        RECT 575.550 203.700 576.750 207.300 ;
        RECT 574.950 201.600 577.050 203.700 ;
        RECT 593.400 202.050 594.450 233.400 ;
        RECT 595.950 206.400 598.050 208.500 ;
        RECT 571.950 193.950 574.050 196.050 ;
        RECT 568.950 190.950 571.050 193.050 ;
        RECT 571.950 191.850 574.050 192.750 ;
        RECT 575.550 189.600 576.750 201.600 ;
        RECT 577.950 199.950 580.050 202.050 ;
        RECT 580.950 199.950 583.050 202.050 ;
        RECT 592.950 199.950 595.050 202.050 ;
        RECT 574.950 187.500 577.050 189.600 ;
        RECT 578.400 172.050 579.450 199.950 ;
        RECT 581.400 190.050 582.450 199.950 ;
        RECT 583.950 197.250 586.050 198.150 ;
        RECT 589.950 197.250 592.050 198.150 ;
        RECT 583.950 193.950 586.050 196.050 ;
        RECT 589.950 193.950 592.050 196.050 ;
        RECT 580.950 187.950 583.050 190.050 ;
        RECT 584.400 172.050 585.450 193.950 ;
        RECT 596.400 189.600 597.600 206.400 ;
        RECT 595.950 187.500 598.050 189.600 ;
        RECT 602.400 181.050 603.450 235.950 ;
        RECT 608.400 232.050 609.450 245.400 ;
        RECT 614.400 244.050 615.450 247.950 ;
        RECT 610.950 241.950 613.050 244.050 ;
        RECT 613.950 241.950 616.050 244.050 ;
        RECT 620.400 243.450 621.450 293.400 ;
        RECT 622.950 289.950 625.050 292.050 ;
        RECT 623.400 271.050 624.450 289.950 ;
        RECT 622.950 268.950 625.050 271.050 ;
        RECT 622.950 266.850 625.050 267.750 ;
        RECT 622.950 247.950 625.050 250.050 ;
        RECT 623.400 244.050 624.450 247.950 ;
        RECT 626.400 244.050 627.450 406.950 ;
        RECT 632.400 397.050 633.450 409.950 ;
        RECT 634.950 406.950 637.050 409.050 ;
        RECT 634.950 403.950 637.050 406.050 ;
        RECT 631.950 394.950 634.050 397.050 ;
        RECT 628.950 383.250 631.050 384.150 ;
        RECT 628.950 379.950 631.050 382.050 ;
        RECT 631.950 379.950 634.050 382.050 ;
        RECT 628.950 341.250 631.050 342.150 ;
        RECT 632.400 340.050 633.450 379.950 ;
        RECT 635.400 373.050 636.450 403.950 ;
        RECT 638.400 379.050 639.450 409.950 ;
        RECT 641.400 409.050 642.450 427.950 ;
        RECT 640.950 406.950 643.050 409.050 ;
        RECT 640.950 389.400 643.050 391.500 ;
        RECT 637.950 376.950 640.050 379.050 ;
        RECT 634.950 370.950 637.050 373.050 ;
        RECT 641.400 372.600 642.600 389.400 ;
        RECT 640.950 370.500 643.050 372.600 ;
        RECT 637.950 351.300 640.050 353.400 ;
        RECT 638.250 347.700 639.450 351.300 ;
        RECT 637.950 345.600 640.050 347.700 ;
        RECT 628.950 339.450 631.050 340.050 ;
        RECT 631.950 339.450 634.050 340.050 ;
        RECT 628.950 338.400 634.050 339.450 ;
        RECT 628.950 337.950 631.050 338.400 ;
        RECT 631.950 337.950 634.050 338.400 ;
        RECT 629.400 316.050 630.450 337.950 ;
        RECT 634.950 334.950 637.050 337.050 ;
        RECT 635.400 327.450 636.450 334.950 ;
        RECT 638.250 333.600 639.450 345.600 ;
        RECT 640.950 339.450 643.050 340.050 ;
        RECT 644.400 339.450 645.450 445.950 ;
        RECT 646.950 439.950 649.050 442.050 ;
        RECT 647.400 406.050 648.450 439.950 ;
        RECT 649.950 422.400 652.050 424.500 ;
        RECT 646.950 403.950 649.050 406.050 ;
        RECT 650.400 405.600 651.600 422.400 ;
        RECT 656.400 417.450 657.450 469.950 ;
        RECT 658.950 466.950 661.050 469.050 ;
        RECT 659.400 460.050 660.450 466.950 ;
        RECT 662.400 463.050 663.450 481.950 ;
        RECT 665.400 478.050 666.450 490.950 ;
        RECT 664.950 475.950 667.050 478.050 ;
        RECT 661.950 460.950 664.050 463.050 ;
        RECT 664.950 461.400 667.050 463.500 ;
        RECT 658.950 457.950 661.050 460.050 ;
        RECT 661.950 458.250 664.050 459.150 ;
        RECT 653.400 416.400 657.450 417.450 ;
        RECT 649.950 403.500 652.050 405.600 ;
        RECT 653.400 387.450 654.450 416.400 ;
        RECT 655.950 413.250 658.050 414.150 ;
        RECT 655.950 409.950 658.050 412.050 ;
        RECT 659.400 397.050 660.450 457.950 ;
        RECT 661.950 454.950 664.050 457.050 ;
        RECT 661.950 451.950 664.050 454.050 ;
        RECT 662.400 445.050 663.450 451.950 ;
        RECT 665.550 449.400 666.750 461.400 ;
        RECT 664.950 447.300 667.050 449.400 ;
        RECT 661.950 442.950 664.050 445.050 ;
        RECT 665.550 443.700 666.750 447.300 ;
        RECT 664.950 441.600 667.050 443.700 ;
        RECT 664.950 430.950 667.050 433.050 ;
        RECT 661.950 413.250 664.050 414.150 ;
        RECT 661.950 409.950 664.050 412.050 ;
        RECT 662.400 409.050 663.450 409.950 ;
        RECT 665.400 409.050 666.450 430.950 ;
        RECT 661.950 406.950 664.050 409.050 ;
        RECT 664.950 406.950 667.050 409.050 ;
        RECT 658.950 394.950 661.050 397.050 ;
        RECT 661.950 389.400 664.050 391.500 ;
        RECT 653.400 386.400 657.450 387.450 ;
        RECT 646.950 382.950 649.050 385.050 ;
        RECT 652.950 384.450 655.050 385.050 ;
        RECT 650.400 383.400 655.050 384.450 ;
        RECT 650.400 382.050 651.450 383.400 ;
        RECT 652.950 382.950 655.050 383.400 ;
        RECT 646.950 380.850 649.050 381.750 ;
        RECT 649.950 379.950 652.050 382.050 ;
        RECT 652.950 380.850 655.050 381.750 ;
        RECT 646.950 376.950 649.050 379.050 ;
        RECT 640.950 338.400 645.450 339.450 ;
        RECT 640.950 337.950 643.050 338.400 ;
        RECT 640.950 335.850 643.050 336.750 ;
        RECT 637.950 331.500 640.050 333.600 ;
        RECT 647.400 333.450 648.450 376.950 ;
        RECT 652.950 351.300 655.050 353.400 ;
        RECT 653.550 347.700 654.750 351.300 ;
        RECT 649.950 343.950 652.050 346.050 ;
        RECT 652.950 345.600 655.050 347.700 ;
        RECT 650.400 340.050 651.450 343.950 ;
        RECT 649.950 337.950 652.050 340.050 ;
        RECT 649.950 335.850 652.050 336.750 ;
        RECT 653.550 333.600 654.750 345.600 ;
        RECT 647.400 332.400 651.450 333.450 ;
        RECT 635.400 326.400 639.450 327.450 ;
        RECT 628.950 313.950 631.050 316.050 ;
        RECT 638.400 313.050 639.450 326.400 ;
        RECT 643.950 319.950 646.050 322.050 ;
        RECT 644.400 313.050 645.450 319.950 ;
        RECT 646.950 316.950 649.050 319.050 ;
        RECT 647.400 316.050 648.450 316.950 ;
        RECT 650.400 316.050 651.450 332.400 ;
        RECT 652.950 331.500 655.050 333.600 ;
        RECT 656.400 322.050 657.450 386.400 ;
        RECT 662.250 377.400 663.450 389.400 ;
        RECT 664.950 386.250 667.050 387.150 ;
        RECT 664.950 382.950 667.050 385.050 ;
        RECT 665.400 382.050 666.450 382.950 ;
        RECT 664.950 379.950 667.050 382.050 ;
        RECT 661.950 375.300 664.050 377.400 ;
        RECT 664.950 376.950 667.050 379.050 ;
        RECT 662.250 371.700 663.450 375.300 ;
        RECT 661.950 369.600 664.050 371.700 ;
        RECT 661.950 341.250 664.050 342.150 ;
        RECT 661.950 337.950 664.050 340.050 ;
        RECT 662.400 322.050 663.450 337.950 ;
        RECT 655.950 319.950 658.050 322.050 ;
        RECT 661.950 319.950 664.050 322.050 ;
        RECT 646.950 313.950 649.050 316.050 ;
        RECT 649.950 313.950 652.050 316.050 ;
        RECT 652.950 313.950 655.050 316.050 ;
        RECT 661.950 313.950 664.050 316.050 ;
        RECT 631.950 312.450 634.050 313.050 ;
        RECT 629.400 311.400 634.050 312.450 ;
        RECT 629.400 292.050 630.450 311.400 ;
        RECT 631.950 310.950 634.050 311.400 ;
        RECT 635.250 311.250 636.750 312.150 ;
        RECT 637.950 310.950 640.050 313.050 ;
        RECT 641.250 311.250 642.750 312.150 ;
        RECT 643.950 310.950 646.050 313.050 ;
        RECT 646.950 311.850 649.050 312.750 ;
        RECT 649.950 311.250 652.050 312.150 ;
        RECT 631.950 308.850 633.750 309.750 ;
        RECT 634.950 307.950 637.050 310.050 ;
        RECT 638.250 308.850 639.750 309.750 ;
        RECT 640.950 307.950 643.050 310.050 ;
        RECT 644.250 308.850 646.050 309.750 ;
        RECT 646.950 307.950 649.050 310.050 ;
        RECT 649.950 307.950 652.050 310.050 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 635.400 289.050 636.450 307.950 ;
        RECT 628.950 286.950 631.050 289.050 ;
        RECT 634.950 286.950 637.050 289.050 ;
        RECT 617.400 242.400 621.450 243.450 ;
        RECT 610.950 239.850 613.050 240.750 ;
        RECT 613.950 239.250 616.050 240.150 ;
        RECT 613.950 235.950 616.050 238.050 ;
        RECT 607.950 229.950 610.050 232.050 ;
        RECT 613.950 200.250 616.050 201.150 ;
        RECT 604.950 197.250 606.750 198.150 ;
        RECT 607.950 196.950 610.050 199.050 ;
        RECT 611.250 197.250 612.750 198.150 ;
        RECT 613.950 196.950 616.050 199.050 ;
        RECT 604.950 193.950 607.050 196.050 ;
        RECT 608.250 194.850 609.750 195.750 ;
        RECT 610.950 193.950 613.050 196.050 ;
        RECT 605.400 187.050 606.450 193.950 ;
        RECT 604.950 184.950 607.050 187.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 601.950 178.950 604.050 181.050 ;
        RECT 571.950 169.950 574.050 172.050 ;
        RECT 577.950 169.950 580.050 172.050 ;
        RECT 583.950 169.950 586.050 172.050 ;
        RECT 568.950 125.250 571.050 126.150 ;
        RECT 568.950 121.950 571.050 124.050 ;
        RECT 565.950 106.950 568.050 109.050 ;
        RECT 565.950 101.400 568.050 103.500 ;
        RECT 550.950 94.950 553.050 97.050 ;
        RECT 556.950 94.950 559.050 97.050 ;
        RECT 550.950 92.850 553.050 93.750 ;
        RECT 556.950 92.850 559.050 93.750 ;
        RECT 566.250 89.400 567.450 101.400 ;
        RECT 572.400 100.050 573.450 169.950 ;
        RECT 574.950 167.250 577.050 168.150 ;
        RECT 580.950 166.950 583.050 169.050 ;
        RECT 584.400 166.050 585.450 169.950 ;
        RECT 586.950 166.950 589.050 169.050 ;
        RECT 574.950 163.950 577.050 166.050 ;
        RECT 577.950 163.950 580.050 166.050 ;
        RECT 580.950 164.850 583.050 165.750 ;
        RECT 583.950 163.950 586.050 166.050 ;
        RECT 586.950 164.850 589.050 165.750 ;
        RECT 574.950 125.250 577.050 126.150 ;
        RECT 574.950 123.450 577.050 124.050 ;
        RECT 578.400 123.450 579.450 163.950 ;
        RECT 586.950 145.950 589.050 148.050 ;
        RECT 583.950 135.300 586.050 137.400 ;
        RECT 584.250 131.700 585.450 135.300 ;
        RECT 583.950 129.600 586.050 131.700 ;
        RECT 574.950 122.400 579.450 123.450 ;
        RECT 574.950 121.950 577.050 122.400 ;
        RECT 578.400 121.050 579.450 122.400 ;
        RECT 577.950 118.950 580.050 121.050 ;
        RECT 584.250 117.600 585.450 129.600 ;
        RECT 587.400 124.050 588.450 145.950 ;
        RECT 590.400 144.450 591.450 178.950 ;
        RECT 610.950 173.400 613.050 175.500 ;
        RECT 607.950 170.250 610.050 171.150 ;
        RECT 601.950 166.950 604.050 169.050 ;
        RECT 607.950 166.950 610.050 169.050 ;
        RECT 592.950 164.250 594.750 165.150 ;
        RECT 595.950 163.950 598.050 166.050 ;
        RECT 599.250 164.250 601.050 165.150 ;
        RECT 592.950 160.950 595.050 163.050 ;
        RECT 596.250 161.850 597.750 162.750 ;
        RECT 598.950 162.450 601.050 163.050 ;
        RECT 602.400 162.450 603.450 166.950 ;
        RECT 604.950 163.950 607.050 166.050 ;
        RECT 598.950 161.400 603.450 162.450 ;
        RECT 598.950 160.950 601.050 161.400 ;
        RECT 593.400 148.050 594.450 160.950 ;
        RECT 592.950 145.950 595.050 148.050 ;
        RECT 590.400 143.400 594.450 144.450 ;
        RECT 589.950 127.950 592.050 130.050 ;
        RECT 586.950 121.950 589.050 124.050 ;
        RECT 586.950 119.850 589.050 120.750 ;
        RECT 590.400 118.050 591.450 127.950 ;
        RECT 583.950 115.500 586.050 117.600 ;
        RECT 589.950 115.950 592.050 118.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 589.950 100.950 592.050 103.050 ;
        RECT 568.950 98.250 571.050 99.150 ;
        RECT 571.950 97.950 574.050 100.050 ;
        RECT 575.400 97.050 576.450 100.950 ;
        RECT 568.950 94.950 571.050 97.050 ;
        RECT 574.950 94.950 577.050 97.050 ;
        RECT 578.250 95.250 579.750 96.150 ;
        RECT 580.950 94.950 583.050 97.050 ;
        RECT 586.950 94.950 589.050 97.050 ;
        RECT 565.950 87.300 568.050 89.400 ;
        RECT 544.950 82.500 547.050 84.600 ;
        RECT 566.250 83.700 567.450 87.300 ;
        RECT 565.950 81.600 568.050 83.700 ;
        RECT 569.400 82.050 570.450 94.950 ;
        RECT 571.950 91.950 574.050 94.050 ;
        RECT 574.950 92.850 576.750 93.750 ;
        RECT 577.950 91.950 580.050 94.050 ;
        RECT 581.250 92.850 582.750 93.750 ;
        RECT 583.950 91.950 586.050 94.050 ;
        RECT 568.950 79.950 571.050 82.050 ;
        RECT 520.950 61.950 523.050 64.050 ;
        RECT 521.400 58.050 522.450 61.950 ;
        RECT 541.950 58.950 544.050 61.050 ;
        RECT 544.950 58.950 547.050 61.050 ;
        RECT 568.950 58.950 571.050 61.050 ;
        RECT 460.950 56.250 463.050 57.150 ;
        RECT 466.950 55.950 469.050 58.050 ;
        RECT 496.950 56.250 499.050 57.150 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 508.950 55.950 511.050 58.050 ;
        RECT 520.950 55.950 523.050 58.050 ;
        RECT 467.400 55.050 468.450 55.950 ;
        RECT 460.950 52.950 463.050 55.050 ;
        RECT 464.250 53.250 465.750 54.150 ;
        RECT 466.950 52.950 469.050 55.050 ;
        RECT 487.950 54.450 490.050 55.050 ;
        RECT 470.250 53.250 472.050 54.150 ;
        RECT 475.950 53.250 478.050 54.150 ;
        RECT 481.950 53.250 484.050 54.150 ;
        RECT 485.400 53.400 490.050 54.450 ;
        RECT 485.400 52.050 486.450 53.400 ;
        RECT 487.950 52.950 490.050 53.400 ;
        RECT 496.950 52.950 499.050 55.050 ;
        RECT 500.250 53.250 501.750 54.150 ;
        RECT 502.950 52.950 505.050 55.050 ;
        RECT 506.250 53.250 508.050 54.150 ;
        RECT 463.950 49.950 466.050 52.050 ;
        RECT 467.250 50.850 468.750 51.750 ;
        RECT 469.950 49.950 472.050 52.050 ;
        RECT 475.950 49.950 478.050 52.050 ;
        RECT 481.950 51.450 484.050 52.050 ;
        RECT 484.950 51.450 487.050 52.050 ;
        RECT 479.250 50.250 480.750 51.150 ;
        RECT 481.950 50.400 487.050 51.450 ;
        RECT 487.950 50.850 490.050 51.750 ;
        RECT 481.950 49.950 484.050 50.400 ;
        RECT 484.950 49.950 487.050 50.400 ;
        RECT 490.950 50.250 493.050 51.150 ;
        RECT 499.950 49.950 502.050 52.050 ;
        RECT 503.250 50.850 504.750 51.750 ;
        RECT 505.950 51.450 508.050 52.050 ;
        RECT 509.400 51.450 510.450 55.950 ;
        RECT 511.950 53.250 513.750 54.150 ;
        RECT 514.950 52.950 517.050 55.050 ;
        RECT 520.950 54.450 523.050 55.050 ;
        RECT 520.950 53.400 525.450 54.450 ;
        RECT 520.950 52.950 523.050 53.400 ;
        RECT 505.950 50.400 510.450 51.450 ;
        RECT 505.950 49.950 508.050 50.400 ;
        RECT 511.950 49.950 514.050 52.050 ;
        RECT 515.250 50.850 517.050 51.750 ;
        RECT 517.950 50.250 520.050 51.150 ;
        RECT 520.950 50.850 523.050 51.750 ;
        RECT 457.950 46.950 460.050 49.050 ;
        RECT 464.400 46.050 465.450 49.950 ;
        RECT 463.950 43.950 466.050 46.050 ;
        RECT 460.950 31.950 463.050 34.050 ;
        RECT 454.950 28.950 457.050 31.050 ;
        RECT 454.950 27.450 457.050 28.050 ;
        RECT 452.400 26.400 457.050 27.450 ;
        RECT 454.950 25.950 457.050 26.400 ;
        RECT 455.400 25.050 456.450 25.950 ;
        RECT 461.400 25.050 462.450 31.950 ;
        RECT 463.950 29.400 466.050 31.500 ;
        RECT 448.950 22.950 451.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 448.950 20.850 451.050 21.750 ;
        RECT 454.950 20.850 457.050 21.750 ;
        RECT 464.250 17.400 465.450 29.400 ;
        RECT 466.950 26.250 469.050 27.150 ;
        RECT 466.950 22.950 469.050 25.050 ;
        RECT 470.400 22.050 471.450 49.950 ;
        RECT 478.950 46.950 481.050 49.050 ;
        RECT 490.950 46.950 493.050 49.050 ;
        RECT 479.400 43.050 480.450 46.950 ;
        RECT 478.950 40.950 481.050 43.050 ;
        RECT 491.400 40.050 492.450 46.950 ;
        RECT 490.950 37.950 493.050 40.050 ;
        RECT 500.400 37.050 501.450 49.950 ;
        RECT 512.400 49.050 513.450 49.950 ;
        RECT 511.950 46.950 514.050 49.050 ;
        RECT 517.950 46.950 520.050 49.050 ;
        RECT 524.400 46.050 525.450 53.400 ;
        RECT 526.950 53.250 529.050 54.150 ;
        RECT 532.950 53.250 535.050 54.150 ;
        RECT 538.950 53.250 541.050 54.150 ;
        RECT 542.400 52.050 543.450 58.950 ;
        RECT 545.400 55.050 546.450 58.950 ;
        RECT 569.400 58.050 570.450 58.950 ;
        RECT 550.950 57.450 553.050 58.050 ;
        RECT 548.400 56.400 553.050 57.450 ;
        RECT 556.950 57.450 559.050 58.050 ;
        RECT 544.950 52.950 547.050 55.050 ;
        RECT 526.950 49.950 529.050 52.050 ;
        RECT 530.250 50.250 531.750 51.150 ;
        RECT 532.950 49.950 535.050 52.050 ;
        RECT 535.950 50.250 537.750 51.150 ;
        RECT 538.950 49.950 541.050 52.050 ;
        RECT 541.950 49.950 544.050 52.050 ;
        RECT 544.950 50.850 547.050 51.750 ;
        RECT 502.950 43.950 505.050 46.050 ;
        RECT 523.950 43.950 526.050 46.050 ;
        RECT 499.950 34.950 502.050 37.050 ;
        RECT 472.950 31.950 475.050 34.050 ;
        RECT 473.400 28.050 474.450 31.950 ;
        RECT 478.950 28.950 481.050 31.050 ;
        RECT 496.950 29.400 499.050 31.500 ;
        RECT 472.950 25.950 475.050 28.050 ;
        RECT 472.950 23.850 475.050 24.750 ;
        RECT 475.950 23.250 478.050 24.150 ;
        RECT 469.950 19.950 472.050 22.050 ;
        RECT 475.950 21.450 478.050 22.050 ;
        RECT 479.400 21.450 480.450 28.950 ;
        RECT 487.950 27.450 490.050 28.050 ;
        RECT 487.950 26.400 492.450 27.450 ;
        RECT 487.950 25.950 490.050 26.400 ;
        RECT 491.400 25.050 492.450 26.400 ;
        RECT 484.950 23.250 487.050 24.150 ;
        RECT 487.950 23.850 490.050 24.750 ;
        RECT 490.950 22.950 493.050 25.050 ;
        RECT 475.950 20.400 480.450 21.450 ;
        RECT 475.950 19.950 478.050 20.400 ;
        RECT 484.950 19.950 487.050 22.050 ;
        RECT 463.950 15.300 466.050 17.400 ;
        RECT 442.950 10.500 445.050 12.600 ;
        RECT 464.250 11.700 465.450 15.300 ;
        RECT 497.400 12.600 498.600 29.400 ;
        RECT 503.400 25.050 504.450 43.950 ;
        RECT 527.400 43.050 528.450 49.950 ;
        RECT 529.950 46.950 532.050 49.050 ;
        RECT 526.950 40.950 529.050 43.050 ;
        RECT 517.950 29.400 520.050 31.500 ;
        RECT 508.950 25.950 511.050 28.050 ;
        RECT 509.400 25.050 510.450 25.950 ;
        RECT 502.950 22.950 505.050 25.050 ;
        RECT 508.950 22.950 511.050 25.050 ;
        RECT 502.950 20.850 505.050 21.750 ;
        RECT 508.950 20.850 511.050 21.750 ;
        RECT 518.250 17.400 519.450 29.400 ;
        RECT 533.400 28.050 534.450 49.950 ;
        RECT 539.400 49.050 540.450 49.950 ;
        RECT 548.400 49.050 549.450 56.400 ;
        RECT 550.950 55.950 553.050 56.400 ;
        RECT 554.250 56.250 555.750 57.150 ;
        RECT 556.950 56.400 561.450 57.450 ;
        RECT 556.950 55.950 559.050 56.400 ;
        RECT 550.950 53.850 552.750 54.750 ;
        RECT 553.950 52.950 556.050 55.050 ;
        RECT 557.250 53.850 559.050 54.750 ;
        RECT 535.950 46.950 538.050 49.050 ;
        RECT 538.950 46.950 541.050 49.050 ;
        RECT 547.950 46.950 550.050 49.050 ;
        RECT 536.400 46.050 537.450 46.950 ;
        RECT 560.400 46.050 561.450 56.400 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 566.250 56.250 567.750 57.150 ;
        RECT 568.950 55.950 571.050 58.050 ;
        RECT 562.950 53.850 564.750 54.750 ;
        RECT 565.950 52.950 568.050 55.050 ;
        RECT 569.250 53.850 571.050 54.750 ;
        RECT 535.950 43.950 538.050 46.050 ;
        RECT 559.950 43.950 562.050 46.050 ;
        RECT 535.950 37.950 538.050 40.050 ;
        RECT 520.950 26.250 523.050 27.150 ;
        RECT 532.950 25.950 535.050 28.050 ;
        RECT 536.400 25.050 537.450 37.950 ;
        RECT 559.950 34.950 562.050 37.050 ;
        RECT 544.950 29.400 547.050 31.500 ;
        RECT 541.950 26.250 544.050 27.150 ;
        RECT 520.950 22.950 523.050 25.050 ;
        RECT 529.950 22.950 532.050 25.050 ;
        RECT 533.250 23.850 534.750 24.750 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 529.950 20.850 532.050 21.750 ;
        RECT 535.950 20.850 538.050 21.750 ;
        RECT 545.550 17.400 546.750 29.400 ;
        RECT 553.950 25.950 556.050 28.050 ;
        RECT 554.400 25.050 555.450 25.950 ;
        RECT 560.400 25.050 561.450 34.950 ;
        RECT 565.950 29.400 568.050 31.500 ;
        RECT 553.950 22.950 556.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 553.950 20.850 556.050 21.750 ;
        RECT 559.950 20.850 562.050 21.750 ;
        RECT 517.950 15.300 520.050 17.400 ;
        RECT 544.950 15.300 547.050 17.400 ;
        RECT 181.950 7.950 184.050 10.050 ;
        RECT 226.950 7.950 229.050 10.050 ;
        RECT 463.950 9.600 466.050 11.700 ;
        RECT 496.950 10.500 499.050 12.600 ;
        RECT 518.250 11.700 519.450 15.300 ;
        RECT 545.550 11.700 546.750 15.300 ;
        RECT 566.400 12.600 567.600 29.400 ;
        RECT 568.950 25.950 571.050 28.050 ;
        RECT 569.400 22.050 570.450 25.950 ;
        RECT 572.400 25.050 573.450 91.950 ;
        RECT 578.400 90.450 579.450 91.950 ;
        RECT 575.400 89.400 579.450 90.450 ;
        RECT 583.950 89.850 586.050 90.750 ;
        RECT 575.400 55.050 576.450 89.400 ;
        RECT 587.400 88.050 588.450 94.950 ;
        RECT 590.400 90.450 591.450 100.950 ;
        RECT 593.400 97.050 594.450 143.400 ;
        RECT 605.400 130.050 606.450 163.950 ;
        RECT 608.400 163.050 609.450 166.950 ;
        RECT 607.950 160.950 610.050 163.050 ;
        RECT 611.550 161.400 612.750 173.400 ;
        RECT 610.950 159.300 613.050 161.400 ;
        RECT 611.550 155.700 612.750 159.300 ;
        RECT 610.950 153.600 613.050 155.700 ;
        RECT 613.950 135.300 616.050 137.400 ;
        RECT 614.550 131.700 615.750 135.300 ;
        RECT 595.950 128.250 598.050 129.150 ;
        RECT 601.950 127.950 604.050 130.050 ;
        RECT 604.950 127.950 607.050 130.050 ;
        RECT 613.950 129.600 616.050 131.700 ;
        RECT 602.400 127.050 603.450 127.950 ;
        RECT 595.950 124.950 598.050 127.050 ;
        RECT 599.250 125.250 600.750 126.150 ;
        RECT 601.950 124.950 604.050 127.050 ;
        RECT 605.250 125.250 607.050 126.150 ;
        RECT 598.950 121.950 601.050 124.050 ;
        RECT 602.250 122.850 603.750 123.750 ;
        RECT 604.950 121.950 607.050 124.050 ;
        RECT 610.950 121.950 613.050 124.050 ;
        RECT 605.400 103.050 606.450 121.950 ;
        RECT 610.950 119.850 613.050 120.750 ;
        RECT 610.950 115.950 613.050 118.050 ;
        RECT 614.550 117.600 615.750 129.600 ;
        RECT 617.400 123.450 618.450 242.400 ;
        RECT 622.950 241.950 625.050 244.050 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 629.400 241.050 630.450 286.950 ;
        RECT 641.400 277.050 642.450 307.950 ;
        RECT 647.400 303.450 648.450 307.950 ;
        RECT 650.400 307.050 651.450 307.950 ;
        RECT 649.950 304.950 652.050 307.050 ;
        RECT 647.400 302.400 651.450 303.450 ;
        RECT 640.950 274.950 643.050 277.050 ;
        RECT 631.950 268.950 634.050 271.050 ;
        RECT 637.950 268.950 640.050 271.050 ;
        RECT 643.950 268.950 646.050 271.050 ;
        RECT 647.250 269.250 649.050 270.150 ;
        RECT 650.400 268.050 651.450 302.400 ;
        RECT 653.400 271.050 654.450 313.950 ;
        RECT 665.400 313.050 666.450 376.950 ;
        RECT 668.400 376.050 669.450 491.400 ;
        RECT 676.950 490.950 679.050 493.050 ;
        RECT 677.400 490.050 678.450 490.950 ;
        RECT 670.950 487.950 673.050 490.050 ;
        RECT 674.250 488.250 675.750 489.150 ;
        RECT 676.950 487.950 679.050 490.050 ;
        RECT 670.950 485.850 672.750 486.750 ;
        RECT 673.950 484.950 676.050 487.050 ;
        RECT 677.250 485.850 679.050 486.750 ;
        RECT 670.950 460.950 673.050 463.050 ;
        RECT 673.950 460.950 676.050 463.050 ;
        RECT 671.400 430.050 672.450 460.950 ;
        RECT 674.400 457.050 675.450 460.950 ;
        RECT 680.400 459.450 681.450 553.950 ;
        RECT 688.950 527.250 691.050 528.150 ;
        RECT 682.950 523.950 685.050 526.050 ;
        RECT 677.400 458.400 681.450 459.450 ;
        RECT 673.950 454.950 676.050 457.050 ;
        RECT 673.950 452.850 676.050 453.750 ;
        RECT 670.950 427.950 673.050 430.050 ;
        RECT 670.950 423.300 673.050 425.400 ;
        RECT 671.250 419.700 672.450 423.300 ;
        RECT 670.950 417.600 673.050 419.700 ;
        RECT 671.250 405.600 672.450 417.600 ;
        RECT 673.950 415.950 676.050 418.050 ;
        RECT 674.400 412.050 675.450 415.950 ;
        RECT 673.950 409.950 676.050 412.050 ;
        RECT 673.950 407.850 676.050 408.750 ;
        RECT 670.950 403.500 673.050 405.600 ;
        RECT 677.400 403.050 678.450 458.400 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 679.950 452.850 682.050 453.750 ;
        RECT 683.400 448.050 684.450 523.950 ;
        RECT 692.400 519.450 693.450 664.950 ;
        RECT 701.400 646.050 702.450 667.950 ;
        RECT 703.950 664.950 706.050 667.050 ;
        RECT 707.250 665.850 708.750 666.750 ;
        RECT 709.950 664.950 712.050 667.050 ;
        RECT 700.950 643.950 703.050 646.050 ;
        RECT 700.950 638.400 703.050 640.500 ;
        RECT 694.950 629.250 697.050 630.150 ;
        RECT 694.950 625.950 697.050 628.050 ;
        RECT 695.400 619.050 696.450 625.950 ;
        RECT 701.400 621.600 702.600 638.400 ;
        RECT 700.950 619.500 703.050 621.600 ;
        RECT 694.950 616.950 697.050 619.050 ;
        RECT 697.950 599.850 700.050 600.750 ;
        RECT 700.950 599.250 703.050 600.150 ;
        RECT 700.950 595.950 703.050 598.050 ;
        RECT 694.950 586.950 697.050 589.050 ;
        RECT 695.400 559.050 696.450 586.950 ;
        RECT 704.400 567.450 705.450 664.950 ;
        RECT 709.950 643.950 712.050 646.050 ;
        RECT 706.950 628.950 709.050 631.050 ;
        RECT 707.400 598.050 708.450 628.950 ;
        RECT 706.950 595.950 709.050 598.050 ;
        RECT 704.400 566.400 708.450 567.450 ;
        RECT 703.950 562.950 706.050 565.050 ;
        RECT 704.400 559.050 705.450 562.950 ;
        RECT 694.950 556.950 697.050 559.050 ;
        RECT 703.950 556.950 706.050 559.050 ;
        RECT 694.950 554.850 697.050 555.750 ;
        RECT 697.950 554.250 700.050 555.150 ;
        RECT 700.950 554.250 703.050 555.150 ;
        RECT 703.950 554.850 706.050 555.750 ;
        RECT 694.950 526.950 697.050 529.050 ;
        RECT 698.250 527.250 699.750 528.150 ;
        RECT 700.950 526.950 703.050 529.050 ;
        RECT 694.950 524.850 696.750 525.750 ;
        RECT 697.950 523.950 700.050 526.050 ;
        RECT 701.250 524.850 702.750 525.750 ;
        RECT 703.950 523.950 706.050 526.050 ;
        RECT 700.950 520.950 703.050 523.050 ;
        RECT 703.950 521.850 706.050 522.750 ;
        RECT 689.400 518.400 693.450 519.450 ;
        RECT 685.950 494.400 688.050 496.500 ;
        RECT 686.400 477.600 687.600 494.400 ;
        RECT 685.950 475.500 688.050 477.600 ;
        RECT 685.950 461.400 688.050 463.500 ;
        RECT 682.950 445.950 685.050 448.050 ;
        RECT 686.400 444.600 687.600 461.400 ;
        RECT 689.400 451.050 690.450 518.400 ;
        RECT 697.950 517.950 700.050 520.050 ;
        RECT 694.950 493.950 697.050 496.050 ;
        RECT 691.950 485.250 694.050 486.150 ;
        RECT 691.950 481.950 694.050 484.050 ;
        RECT 695.400 483.450 696.450 493.950 ;
        RECT 698.400 490.050 699.450 517.950 ;
        RECT 701.400 493.050 702.450 520.950 ;
        RECT 707.400 501.450 708.450 566.400 ;
        RECT 704.400 500.400 708.450 501.450 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 697.950 487.950 700.050 490.050 ;
        RECT 697.950 485.250 700.050 486.150 ;
        RECT 700.950 484.950 703.050 487.050 ;
        RECT 697.950 483.450 700.050 484.050 ;
        RECT 695.400 482.400 700.050 483.450 ;
        RECT 692.400 457.050 693.450 481.950 ;
        RECT 695.400 463.050 696.450 482.400 ;
        RECT 697.950 481.950 700.050 482.400 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 698.400 466.050 699.450 478.950 ;
        RECT 697.950 463.950 700.050 466.050 ;
        RECT 694.950 460.950 697.050 463.050 ;
        RECT 697.950 460.950 700.050 463.050 ;
        RECT 698.400 459.450 699.450 460.950 ;
        RECT 701.400 460.050 702.450 484.950 ;
        RECT 704.400 484.050 705.450 500.400 ;
        RECT 706.950 495.300 709.050 497.400 ;
        RECT 707.250 491.700 708.450 495.300 ;
        RECT 706.950 489.600 709.050 491.700 ;
        RECT 703.950 481.950 706.050 484.050 ;
        RECT 695.400 458.400 699.450 459.450 ;
        RECT 695.400 457.050 696.450 458.400 ;
        RECT 700.950 457.950 703.050 460.050 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 694.950 454.950 697.050 457.050 ;
        RECT 698.250 455.250 699.750 456.150 ;
        RECT 700.950 454.950 703.050 457.050 ;
        RECT 704.400 456.450 705.450 481.950 ;
        RECT 707.250 477.600 708.450 489.600 ;
        RECT 710.400 487.050 711.450 643.950 ;
        RECT 715.950 556.950 718.050 559.050 ;
        RECT 712.950 523.950 715.050 526.050 ;
        RECT 709.950 484.950 712.050 487.050 ;
        RECT 709.950 481.950 712.050 484.050 ;
        RECT 709.950 479.850 712.050 480.750 ;
        RECT 706.950 475.500 709.050 477.600 ;
        RECT 709.950 475.950 712.050 478.050 ;
        RECT 710.400 463.050 711.450 475.950 ;
        RECT 709.950 460.950 712.050 463.050 ;
        RECT 709.950 457.950 712.050 460.050 ;
        RECT 704.400 455.400 708.450 456.450 ;
        RECT 691.950 451.950 694.050 454.050 ;
        RECT 694.950 452.850 696.750 453.750 ;
        RECT 697.950 451.950 700.050 454.050 ;
        RECT 701.250 452.850 702.750 453.750 ;
        RECT 703.950 451.950 706.050 454.050 ;
        RECT 688.950 448.950 691.050 451.050 ;
        RECT 685.950 442.500 688.050 444.600 ;
        RECT 692.400 439.050 693.450 451.950 ;
        RECT 698.400 451.050 699.450 451.950 ;
        RECT 697.950 448.950 700.050 451.050 ;
        RECT 700.950 448.950 703.050 451.050 ;
        RECT 703.950 449.850 706.050 450.750 ;
        RECT 691.950 436.950 694.050 439.050 ;
        RECT 701.400 421.050 702.450 448.950 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 682.950 418.950 685.050 421.050 ;
        RECT 691.950 418.950 694.050 421.050 ;
        RECT 700.950 418.950 703.050 421.050 ;
        RECT 683.400 415.050 684.450 418.950 ;
        RECT 688.950 416.250 691.050 417.150 ;
        RECT 679.950 413.250 681.750 414.150 ;
        RECT 682.950 412.950 685.050 415.050 ;
        RECT 686.250 413.250 687.750 414.150 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 679.950 409.950 682.050 412.050 ;
        RECT 683.250 410.850 684.750 411.750 ;
        RECT 685.950 409.950 688.050 412.050 ;
        RECT 680.400 409.050 681.450 409.950 ;
        RECT 689.400 409.050 690.450 412.950 ;
        RECT 679.950 406.950 682.050 409.050 ;
        RECT 688.950 406.950 691.050 409.050 ;
        RECT 682.950 403.950 685.050 406.050 ;
        RECT 676.950 400.950 679.050 403.050 ;
        RECT 670.950 385.950 673.050 388.050 ;
        RECT 671.400 385.050 672.450 385.950 ;
        RECT 670.950 382.950 673.050 385.050 ;
        RECT 674.250 383.250 675.750 384.150 ;
        RECT 676.950 382.950 679.050 385.050 ;
        RECT 679.950 382.950 682.050 385.050 ;
        RECT 680.400 382.050 681.450 382.950 ;
        RECT 670.950 380.850 672.750 381.750 ;
        RECT 673.950 379.950 676.050 382.050 ;
        RECT 677.250 380.850 678.750 381.750 ;
        RECT 679.950 379.950 682.050 382.050 ;
        RECT 667.950 373.950 670.050 376.050 ;
        RECT 674.400 373.050 675.450 379.950 ;
        RECT 683.400 379.050 684.450 403.950 ;
        RECT 692.400 385.050 693.450 418.950 ;
        RECT 701.400 418.050 702.450 418.950 ;
        RECT 694.950 415.950 697.050 418.050 ;
        RECT 698.250 416.250 699.750 417.150 ;
        RECT 700.950 415.950 703.050 418.050 ;
        RECT 694.950 413.850 696.750 414.750 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 701.250 413.850 703.050 414.750 ;
        RECT 694.950 409.950 697.050 412.050 ;
        RECT 688.950 382.950 691.050 385.050 ;
        RECT 691.950 382.950 694.050 385.050 ;
        RECT 689.400 382.050 690.450 382.950 ;
        RECT 685.950 380.250 687.750 381.150 ;
        RECT 688.950 379.950 691.050 382.050 ;
        RECT 692.250 380.250 694.050 381.150 ;
        RECT 695.400 379.050 696.450 409.950 ;
        RECT 698.400 409.050 699.450 412.950 ;
        RECT 700.950 409.950 703.050 412.050 ;
        RECT 697.950 406.950 700.050 409.050 ;
        RECT 701.400 382.050 702.450 409.950 ;
        RECT 704.400 406.050 705.450 445.950 ;
        RECT 703.950 403.950 706.050 406.050 ;
        RECT 697.950 380.250 699.750 381.150 ;
        RECT 700.950 379.950 703.050 382.050 ;
        RECT 704.250 380.250 706.050 381.150 ;
        RECT 679.950 377.850 682.050 378.750 ;
        RECT 682.950 376.950 685.050 379.050 ;
        RECT 685.950 376.950 688.050 379.050 ;
        RECT 689.250 377.850 690.750 378.750 ;
        RECT 691.950 376.950 694.050 379.050 ;
        RECT 694.950 376.950 697.050 379.050 ;
        RECT 697.950 376.950 700.050 379.050 ;
        RECT 701.250 377.850 702.750 378.750 ;
        RECT 703.950 376.950 706.050 379.050 ;
        RECT 673.950 370.950 676.050 373.050 ;
        RECT 673.950 350.400 676.050 352.500 ;
        RECT 686.400 352.050 687.450 376.950 ;
        RECT 692.400 373.050 693.450 376.950 ;
        RECT 698.400 376.050 699.450 376.950 ;
        RECT 697.950 373.950 700.050 376.050 ;
        RECT 691.950 370.950 694.050 373.050 ;
        RECT 667.950 341.250 670.050 342.150 ;
        RECT 667.950 337.950 670.050 340.050 ;
        RECT 674.400 333.600 675.600 350.400 ;
        RECT 685.950 349.950 688.050 352.050 ;
        RECT 698.400 351.450 699.450 373.950 ;
        RECT 703.950 370.950 706.050 373.050 ;
        RECT 695.400 350.400 699.450 351.450 ;
        RECT 685.950 346.950 688.050 349.050 ;
        RECT 679.950 343.950 682.050 346.050 ;
        RECT 673.950 331.500 676.050 333.600 ;
        RECT 680.400 325.050 681.450 343.950 ;
        RECT 686.400 343.050 687.450 346.950 ;
        RECT 691.950 344.250 694.050 345.150 ;
        RECT 682.950 341.250 684.750 342.150 ;
        RECT 685.950 340.950 688.050 343.050 ;
        RECT 689.250 341.250 690.750 342.150 ;
        RECT 691.950 340.950 694.050 343.050 ;
        RECT 682.950 337.950 685.050 340.050 ;
        RECT 686.250 338.850 687.750 339.750 ;
        RECT 688.950 337.950 691.050 340.050 ;
        RECT 683.400 328.050 684.450 337.950 ;
        RECT 682.950 325.950 685.050 328.050 ;
        RECT 695.400 327.450 696.450 350.400 ;
        RECT 704.400 349.050 705.450 370.950 ;
        RECT 703.950 346.950 706.050 349.050 ;
        RECT 704.400 346.050 705.450 346.950 ;
        RECT 697.950 343.950 700.050 346.050 ;
        RECT 701.250 344.250 702.750 345.150 ;
        RECT 703.950 343.950 706.050 346.050 ;
        RECT 697.950 341.850 699.750 342.750 ;
        RECT 700.950 340.950 703.050 343.050 ;
        RECT 704.250 341.850 706.050 342.750 ;
        RECT 700.950 337.950 703.050 340.050 ;
        RECT 695.400 326.400 699.450 327.450 ;
        RECT 679.950 322.950 682.050 325.050 ;
        RECT 688.950 322.950 691.050 325.050 ;
        RECT 679.950 319.950 682.050 322.050 ;
        RECT 670.950 316.950 673.050 319.050 ;
        RECT 671.400 313.050 672.450 316.950 ;
        RECT 673.950 313.950 676.050 316.050 ;
        RECT 658.950 312.450 661.050 313.050 ;
        RECT 656.400 311.400 661.050 312.450 ;
        RECT 662.250 311.850 663.750 312.750 ;
        RECT 664.950 312.450 667.050 313.050 ;
        RECT 656.400 310.050 657.450 311.400 ;
        RECT 658.950 310.950 661.050 311.400 ;
        RECT 664.950 311.400 669.450 312.450 ;
        RECT 664.950 310.950 667.050 311.400 ;
        RECT 655.950 307.950 658.050 310.050 ;
        RECT 658.950 308.850 661.050 309.750 ;
        RECT 664.950 308.850 667.050 309.750 ;
        RECT 668.400 273.450 669.450 311.400 ;
        RECT 670.950 310.950 673.050 313.050 ;
        RECT 674.250 311.850 675.750 312.750 ;
        RECT 676.950 310.950 679.050 313.050 ;
        RECT 670.950 308.850 673.050 309.750 ;
        RECT 673.950 307.950 676.050 310.050 ;
        RECT 676.950 308.850 679.050 309.750 ;
        RECT 670.950 279.300 673.050 281.400 ;
        RECT 671.550 275.700 672.750 279.300 ;
        RECT 670.950 273.600 673.050 275.700 ;
        RECT 665.400 272.400 669.450 273.450 ;
        RECT 652.950 268.950 655.050 271.050 ;
        RECT 655.950 269.250 658.050 270.150 ;
        RECT 661.950 269.250 664.050 270.150 ;
        RECT 631.950 266.850 634.050 267.750 ;
        RECT 634.950 266.250 637.050 267.150 ;
        RECT 637.950 266.850 640.050 267.750 ;
        RECT 640.950 266.250 643.050 267.150 ;
        RECT 643.950 266.850 645.750 267.750 ;
        RECT 646.950 265.950 649.050 268.050 ;
        RECT 649.950 265.950 652.050 268.050 ;
        RECT 653.400 267.450 654.450 268.950 ;
        RECT 655.950 267.450 658.050 268.050 ;
        RECT 653.400 266.400 658.050 267.450 ;
        RECT 655.950 265.950 658.050 266.400 ;
        RECT 659.250 266.250 660.750 267.150 ;
        RECT 661.950 265.950 664.050 268.050 ;
        RECT 634.950 262.950 637.050 265.050 ;
        RECT 640.950 262.950 643.050 265.050 ;
        RECT 634.950 259.950 637.050 262.050 ;
        RECT 631.950 253.950 634.050 256.050 ;
        RECT 632.400 244.050 633.450 253.950 ;
        RECT 631.950 241.950 634.050 244.050 ;
        RECT 635.400 241.050 636.450 259.950 ;
        RECT 641.400 256.050 642.450 262.950 ;
        RECT 640.950 253.950 643.050 256.050 ;
        RECT 643.950 250.950 646.050 253.050 ;
        RECT 640.950 247.950 643.050 250.050 ;
        RECT 637.950 241.950 640.050 244.050 ;
        RECT 641.400 241.050 642.450 247.950 ;
        RECT 619.950 239.250 622.050 240.150 ;
        RECT 622.950 239.850 625.050 240.750 ;
        RECT 625.950 239.250 627.750 240.150 ;
        RECT 628.950 238.950 631.050 241.050 ;
        RECT 634.950 240.450 637.050 241.050 ;
        RECT 632.400 239.400 637.050 240.450 ;
        RECT 638.250 239.850 639.750 240.750 ;
        RECT 632.400 238.050 633.450 239.400 ;
        RECT 634.950 238.950 637.050 239.400 ;
        RECT 640.950 238.950 643.050 241.050 ;
        RECT 619.950 235.950 622.050 238.050 ;
        RECT 625.950 235.950 628.050 238.050 ;
        RECT 629.250 236.850 631.050 237.750 ;
        RECT 631.950 235.950 634.050 238.050 ;
        RECT 634.950 236.850 637.050 237.750 ;
        RECT 637.950 235.950 640.050 238.050 ;
        RECT 640.950 236.850 643.050 237.750 ;
        RECT 620.400 232.050 621.450 235.950 ;
        RECT 619.950 229.950 622.050 232.050 ;
        RECT 626.400 211.050 627.450 235.950 ;
        RECT 631.950 232.950 634.050 235.050 ;
        RECT 628.950 229.950 631.050 232.050 ;
        RECT 625.950 208.950 628.050 211.050 ;
        RECT 625.950 205.950 628.050 208.050 ;
        RECT 619.950 202.950 622.050 205.050 ;
        RECT 620.400 202.050 621.450 202.950 ;
        RECT 626.400 202.050 627.450 205.950 ;
        RECT 619.950 199.950 622.050 202.050 ;
        RECT 623.250 200.250 624.750 201.150 ;
        RECT 625.950 199.950 628.050 202.050 ;
        RECT 619.950 197.850 621.750 198.750 ;
        RECT 622.950 196.950 625.050 199.050 ;
        RECT 626.250 197.850 628.050 198.750 ;
        RECT 619.950 169.950 622.050 172.050 ;
        RECT 625.950 169.950 628.050 172.050 ;
        RECT 620.400 169.050 621.450 169.950 ;
        RECT 626.400 169.050 627.450 169.950 ;
        RECT 619.950 166.950 622.050 169.050 ;
        RECT 625.950 166.950 628.050 169.050 ;
        RECT 619.950 164.850 622.050 165.750 ;
        RECT 625.950 164.850 628.050 165.750 ;
        RECT 629.400 163.050 630.450 229.950 ;
        RECT 632.400 226.050 633.450 232.950 ;
        RECT 638.400 232.050 639.450 235.950 ;
        RECT 637.950 229.950 640.050 232.050 ;
        RECT 631.950 223.950 634.050 226.050 ;
        RECT 644.400 214.050 645.450 250.950 ;
        RECT 647.400 250.050 648.450 265.950 ;
        RECT 650.400 264.450 651.450 265.950 ;
        RECT 650.400 263.400 654.450 264.450 ;
        RECT 649.950 253.950 652.050 256.050 ;
        RECT 646.950 247.950 649.050 250.050 ;
        RECT 650.400 244.050 651.450 253.950 ;
        RECT 653.400 244.050 654.450 263.400 ;
        RECT 658.950 262.950 661.050 265.050 ;
        RECT 658.950 259.950 661.050 262.050 ;
        RECT 649.950 241.950 652.050 244.050 ;
        RECT 652.950 241.950 655.050 244.050 ;
        RECT 646.950 239.250 649.050 240.150 ;
        RECT 649.950 239.850 652.050 240.750 ;
        RECT 652.950 239.250 654.750 240.150 ;
        RECT 655.950 238.950 658.050 241.050 ;
        RECT 646.950 235.950 649.050 238.050 ;
        RECT 652.950 235.950 655.050 238.050 ;
        RECT 656.250 236.850 658.050 237.750 ;
        RECT 647.400 235.050 648.450 235.950 ;
        RECT 646.950 232.950 649.050 235.050 ;
        RECT 652.950 232.950 655.050 235.050 ;
        RECT 637.950 211.950 640.050 214.050 ;
        RECT 643.950 211.950 646.050 214.050 ;
        RECT 631.950 202.950 634.050 205.050 ;
        RECT 632.400 195.450 633.450 202.950 ;
        RECT 634.950 197.250 637.050 198.150 ;
        RECT 634.950 195.450 637.050 196.050 ;
        RECT 632.400 194.400 637.050 195.450 ;
        RECT 634.950 193.950 637.050 194.400 ;
        RECT 631.950 173.400 634.050 175.500 ;
        RECT 628.950 160.950 631.050 163.050 ;
        RECT 632.400 156.600 633.600 173.400 ;
        RECT 631.950 154.500 634.050 156.600 ;
        RECT 634.950 134.400 637.050 136.500 ;
        RECT 622.950 125.250 625.050 126.150 ;
        RECT 628.950 125.250 631.050 126.150 ;
        RECT 617.400 122.400 621.450 123.450 ;
        RECT 616.950 118.950 619.050 121.050 ;
        RECT 604.950 100.950 607.050 103.050 ;
        RECT 607.950 101.400 610.050 103.500 ;
        RECT 601.950 97.950 604.050 100.050 ;
        RECT 604.950 98.250 607.050 99.150 ;
        RECT 592.950 94.950 595.050 97.050 ;
        RECT 592.950 92.250 594.750 93.150 ;
        RECT 595.950 91.950 598.050 94.050 ;
        RECT 599.250 92.250 601.050 93.150 ;
        RECT 592.950 90.450 595.050 91.050 ;
        RECT 590.400 89.400 595.050 90.450 ;
        RECT 596.250 89.850 597.750 90.750 ;
        RECT 592.950 88.950 595.050 89.400 ;
        RECT 598.950 88.950 601.050 91.050 ;
        RECT 586.950 85.950 589.050 88.050 ;
        RECT 598.950 79.950 601.050 82.050 ;
        RECT 583.950 61.950 586.050 64.050 ;
        RECT 577.950 56.250 580.050 57.150 ;
        RECT 584.400 55.050 585.450 61.950 ;
        RECT 574.950 52.950 577.050 55.050 ;
        RECT 577.950 52.950 580.050 55.050 ;
        RECT 581.250 53.250 582.750 54.150 ;
        RECT 583.950 52.950 586.050 55.050 ;
        RECT 592.950 54.450 595.050 55.050 ;
        RECT 587.250 53.250 589.050 54.150 ;
        RECT 590.400 53.400 595.050 54.450 ;
        RECT 578.400 52.050 579.450 52.950 ;
        RECT 577.950 49.950 580.050 52.050 ;
        RECT 580.950 49.950 583.050 52.050 ;
        RECT 584.250 50.850 585.750 51.750 ;
        RECT 586.950 51.450 589.050 52.050 ;
        RECT 590.400 51.450 591.450 53.400 ;
        RECT 592.950 52.950 595.050 53.400 ;
        RECT 586.950 50.400 591.450 51.450 ;
        RECT 592.950 50.850 595.050 51.750 ;
        RECT 586.950 49.950 589.050 50.400 ;
        RECT 595.950 50.250 598.050 51.150 ;
        RECT 581.400 43.050 582.450 49.950 ;
        RECT 580.950 40.950 583.050 43.050 ;
        RECT 587.400 40.050 588.450 49.950 ;
        RECT 595.950 46.950 598.050 49.050 ;
        RECT 596.400 46.050 597.450 46.950 ;
        RECT 589.950 43.950 592.050 46.050 ;
        RECT 595.950 43.950 598.050 46.050 ;
        RECT 586.950 37.950 589.050 40.050 ;
        RECT 574.950 25.950 577.050 28.050 ;
        RECT 590.400 25.050 591.450 43.950 ;
        RECT 595.950 37.950 598.050 40.050 ;
        RECT 592.950 31.950 595.050 34.050 ;
        RECT 571.950 22.950 574.050 25.050 ;
        RECT 574.950 23.850 577.050 24.750 ;
        RECT 577.950 23.250 580.050 24.150 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 587.250 23.250 588.750 24.150 ;
        RECT 589.950 22.950 592.050 25.050 ;
        RECT 568.950 19.950 571.050 22.050 ;
        RECT 577.950 21.450 580.050 22.050 ;
        RECT 581.400 21.450 582.450 22.950 ;
        RECT 593.400 22.050 594.450 31.950 ;
        RECT 577.950 20.400 582.450 21.450 ;
        RECT 583.950 20.850 585.750 21.750 ;
        RECT 577.950 19.950 580.050 20.400 ;
        RECT 586.950 19.950 589.050 22.050 ;
        RECT 590.250 20.850 591.750 21.750 ;
        RECT 592.950 19.950 595.050 22.050 ;
        RECT 587.400 19.050 588.450 19.950 ;
        RECT 596.400 19.050 597.450 37.950 ;
        RECT 599.400 28.050 600.450 79.950 ;
        RECT 602.400 55.050 603.450 97.950 ;
        RECT 604.950 94.950 607.050 97.050 ;
        RECT 605.400 91.050 606.450 94.950 ;
        RECT 604.950 88.950 607.050 91.050 ;
        RECT 608.550 89.400 609.750 101.400 ;
        RECT 607.950 87.300 610.050 89.400 ;
        RECT 608.550 83.700 609.750 87.300 ;
        RECT 607.950 81.600 610.050 83.700 ;
        RECT 611.400 55.050 612.450 115.950 ;
        RECT 613.950 115.500 616.050 117.600 ;
        RECT 617.400 97.050 618.450 118.950 ;
        RECT 613.950 94.950 616.050 97.050 ;
        RECT 616.950 94.950 619.050 97.050 ;
        RECT 614.400 88.050 615.450 94.950 ;
        RECT 616.950 92.850 619.050 93.750 ;
        RECT 613.950 85.950 616.050 88.050 ;
        RECT 613.950 63.300 616.050 65.400 ;
        RECT 614.550 59.700 615.750 63.300 ;
        RECT 613.950 57.600 616.050 59.700 ;
        RECT 601.950 52.950 604.050 55.050 ;
        RECT 610.950 52.950 613.050 55.050 ;
        RECT 601.950 50.850 604.050 51.750 ;
        RECT 604.950 50.250 607.050 51.150 ;
        RECT 610.950 49.950 613.050 52.050 ;
        RECT 604.950 46.950 607.050 49.050 ;
        RECT 610.950 47.850 613.050 48.750 ;
        RECT 614.550 45.600 615.750 57.600 ;
        RECT 616.950 49.950 619.050 52.050 ;
        RECT 617.400 46.050 618.450 49.950 ;
        RECT 620.400 49.050 621.450 122.400 ;
        RECT 622.950 121.950 625.050 124.050 ;
        RECT 628.950 121.950 631.050 124.050 ;
        RECT 623.400 121.050 624.450 121.950 ;
        RECT 622.950 118.950 625.050 121.050 ;
        RECT 625.950 118.950 628.050 121.050 ;
        RECT 622.950 94.950 625.050 97.050 ;
        RECT 622.950 92.850 625.050 93.750 ;
        RECT 622.950 53.250 625.050 54.150 ;
        RECT 622.950 51.450 625.050 52.050 ;
        RECT 626.400 51.450 627.450 118.950 ;
        RECT 629.400 115.050 630.450 121.950 ;
        RECT 635.400 117.600 636.600 134.400 ;
        RECT 638.400 124.050 639.450 211.950 ;
        RECT 643.950 208.950 646.050 211.050 ;
        RECT 644.400 201.450 645.450 208.950 ;
        RECT 653.400 202.050 654.450 232.950 ;
        RECT 655.950 226.950 658.050 229.050 ;
        RECT 646.950 201.450 649.050 202.050 ;
        RECT 644.400 200.400 649.050 201.450 ;
        RECT 640.950 197.250 643.050 198.150 ;
        RECT 640.950 193.950 643.050 196.050 ;
        RECT 641.400 178.050 642.450 193.950 ;
        RECT 640.950 175.950 643.050 178.050 ;
        RECT 644.400 169.050 645.450 200.400 ;
        RECT 646.950 199.950 649.050 200.400 ;
        RECT 650.250 200.250 651.750 201.150 ;
        RECT 652.950 199.950 655.050 202.050 ;
        RECT 646.950 197.850 648.750 198.750 ;
        RECT 649.950 196.950 652.050 199.050 ;
        RECT 653.250 197.850 655.050 198.750 ;
        RECT 656.400 196.050 657.450 226.950 ;
        RECT 659.400 208.050 660.450 259.950 ;
        RECT 661.950 250.950 664.050 253.050 ;
        RECT 662.400 250.050 663.450 250.950 ;
        RECT 665.400 250.050 666.450 272.400 ;
        RECT 667.950 268.950 670.050 271.050 ;
        RECT 668.400 268.050 669.450 268.950 ;
        RECT 667.950 265.950 670.050 268.050 ;
        RECT 667.950 263.850 670.050 264.750 ;
        RECT 671.550 261.600 672.750 273.600 ;
        RECT 674.400 268.050 675.450 307.950 ;
        RECT 676.950 274.950 679.050 277.050 ;
        RECT 673.950 265.950 676.050 268.050 ;
        RECT 670.950 259.500 673.050 261.600 ;
        RECT 667.950 256.950 670.050 259.050 ;
        RECT 661.950 247.950 664.050 250.050 ;
        RECT 664.950 247.950 667.050 250.050 ;
        RECT 662.400 244.050 663.450 247.950 ;
        RECT 661.950 241.950 664.050 244.050 ;
        RECT 661.950 239.850 664.050 240.750 ;
        RECT 664.950 239.250 667.050 240.150 ;
        RECT 664.950 235.950 667.050 238.050 ;
        RECT 668.400 235.050 669.450 256.950 ;
        RECT 670.950 253.950 673.050 256.050 ;
        RECT 671.400 244.050 672.450 253.950 ;
        RECT 677.400 244.050 678.450 274.950 ;
        RECT 680.400 273.450 681.450 319.950 ;
        RECT 685.950 317.400 688.050 319.500 ;
        RECT 682.950 314.250 685.050 315.150 ;
        RECT 682.950 310.950 685.050 313.050 ;
        RECT 683.400 277.050 684.450 310.950 ;
        RECT 686.550 305.400 687.750 317.400 ;
        RECT 685.950 303.300 688.050 305.400 ;
        RECT 686.550 299.700 687.750 303.300 ;
        RECT 685.950 297.600 688.050 299.700 ;
        RECT 682.950 274.950 685.050 277.050 ;
        RECT 680.400 272.400 684.450 273.450 ;
        RECT 679.950 269.250 682.050 270.150 ;
        RECT 679.950 267.450 682.050 268.050 ;
        RECT 683.400 267.450 684.450 272.400 ;
        RECT 685.950 269.250 688.050 270.150 ;
        RECT 679.950 266.400 684.450 267.450 ;
        RECT 679.950 265.950 682.050 266.400 ;
        RECT 685.950 265.950 688.050 268.050 ;
        RECT 689.400 262.050 690.450 322.950 ;
        RECT 694.950 319.950 697.050 322.050 ;
        RECT 695.400 313.050 696.450 319.950 ;
        RECT 694.950 310.950 697.050 313.050 ;
        RECT 694.950 308.850 697.050 309.750 ;
        RECT 691.950 278.400 694.050 280.500 ;
        RECT 688.950 259.950 691.050 262.050 ;
        RECT 692.400 261.600 693.600 278.400 ;
        RECT 698.400 274.050 699.450 326.400 ;
        RECT 701.400 313.050 702.450 337.950 ;
        RECT 707.400 324.450 708.450 455.400 ;
        RECT 710.400 454.050 711.450 457.950 ;
        RECT 709.950 451.950 712.050 454.050 ;
        RECT 709.950 448.950 712.050 451.050 ;
        RECT 710.400 340.050 711.450 448.950 ;
        RECT 713.400 412.050 714.450 523.950 ;
        RECT 716.400 463.050 717.450 556.950 ;
        RECT 715.950 460.950 718.050 463.050 ;
        RECT 715.950 457.950 718.050 460.050 ;
        RECT 716.400 439.050 717.450 457.950 ;
        RECT 715.950 436.950 718.050 439.050 ;
        RECT 712.950 409.950 715.050 412.050 ;
        RECT 715.950 349.950 718.050 352.050 ;
        RECT 709.950 337.950 712.050 340.050 ;
        RECT 704.400 323.400 708.450 324.450 ;
        RECT 700.950 310.950 703.050 313.050 ;
        RECT 700.950 308.850 703.050 309.750 ;
        RECT 704.400 274.050 705.450 323.400 ;
        RECT 706.950 317.400 709.050 319.500 ;
        RECT 707.400 300.600 708.600 317.400 ;
        RECT 706.950 298.500 709.050 300.600 ;
        RECT 697.950 271.950 700.050 274.050 ;
        RECT 703.950 271.950 706.050 274.050 ;
        RECT 707.250 272.250 708.750 273.150 ;
        RECT 709.950 271.950 712.050 274.050 ;
        RECT 691.950 259.500 694.050 261.600 ;
        RECT 698.400 259.050 699.450 271.950 ;
        RECT 703.950 269.850 705.750 270.750 ;
        RECT 706.950 268.950 709.050 271.050 ;
        RECT 710.250 269.850 712.050 270.750 ;
        RECT 700.950 265.950 703.050 268.050 ;
        RECT 697.950 256.950 700.050 259.050 ;
        RECT 697.950 250.950 700.050 253.050 ;
        RECT 679.950 247.950 682.050 250.050 ;
        RECT 670.950 241.950 673.050 244.050 ;
        RECT 676.950 241.950 679.050 244.050 ;
        RECT 670.950 239.850 673.050 240.750 ;
        RECT 673.950 239.250 676.050 240.150 ;
        RECT 676.950 238.950 679.050 241.050 ;
        RECT 673.950 235.950 676.050 238.050 ;
        RECT 667.950 232.950 670.050 235.050 ;
        RECT 670.950 232.950 673.050 235.050 ;
        RECT 658.950 205.950 661.050 208.050 ;
        RECT 671.400 205.050 672.450 232.950 ;
        RECT 670.950 202.950 673.050 205.050 ;
        RECT 658.950 200.250 661.050 201.150 ;
        RECT 658.950 196.950 661.050 199.050 ;
        RECT 662.250 197.250 663.750 198.150 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 671.400 198.450 672.450 202.950 ;
        RECT 677.400 201.450 678.450 238.950 ;
        RECT 680.400 237.450 681.450 247.950 ;
        RECT 685.950 241.950 688.050 244.050 ;
        RECT 682.950 239.250 685.050 240.150 ;
        RECT 685.950 239.850 688.050 240.750 ;
        RECT 688.950 238.950 691.050 241.050 ;
        RECT 692.250 239.250 693.750 240.150 ;
        RECT 694.950 238.950 697.050 241.050 ;
        RECT 698.400 238.050 699.450 250.950 ;
        RECT 701.400 244.050 702.450 265.950 ;
        RECT 700.950 241.950 703.050 244.050 ;
        RECT 707.400 241.050 708.450 268.950 ;
        RECT 716.400 241.050 717.450 349.950 ;
        RECT 700.950 238.950 703.050 241.050 ;
        RECT 706.950 238.950 709.050 241.050 ;
        RECT 712.950 238.950 715.050 241.050 ;
        RECT 715.950 238.950 718.050 241.050 ;
        RECT 682.950 237.450 685.050 238.050 ;
        RECT 680.400 236.400 685.050 237.450 ;
        RECT 688.950 236.850 690.750 237.750 ;
        RECT 682.950 235.950 685.050 236.400 ;
        RECT 691.950 235.950 694.050 238.050 ;
        RECT 695.250 236.850 696.750 237.750 ;
        RECT 697.950 235.950 700.050 238.050 ;
        RECT 697.950 233.850 700.050 234.750 ;
        RECT 694.950 228.450 697.050 229.050 ;
        RECT 697.950 228.450 700.050 229.050 ;
        RECT 694.950 227.400 700.050 228.450 ;
        RECT 694.950 226.950 697.050 227.400 ;
        RECT 697.950 226.950 700.050 227.400 ;
        RECT 701.400 205.050 702.450 238.950 ;
        RECT 703.950 236.250 705.750 237.150 ;
        RECT 706.950 235.950 709.050 238.050 ;
        RECT 710.250 236.250 712.050 237.150 ;
        RECT 703.950 232.950 706.050 235.050 ;
        RECT 707.250 233.850 708.750 234.750 ;
        RECT 709.950 232.950 712.050 235.050 ;
        RECT 694.950 202.950 697.050 205.050 ;
        RECT 700.950 202.950 703.050 205.050 ;
        RECT 703.950 202.950 706.050 205.050 ;
        RECT 673.950 200.250 676.050 201.150 ;
        RECT 677.400 200.400 681.450 201.450 ;
        RECT 680.400 199.050 681.450 200.400 ;
        RECT 673.950 198.450 676.050 199.050 ;
        RECT 668.250 197.250 670.050 198.150 ;
        RECT 671.400 197.400 676.050 198.450 ;
        RECT 655.950 193.950 658.050 196.050 ;
        RECT 661.950 193.950 664.050 196.050 ;
        RECT 665.250 194.850 666.750 195.750 ;
        RECT 667.950 193.950 670.050 196.050 ;
        RECT 668.400 190.050 669.450 193.950 ;
        RECT 667.950 187.950 670.050 190.050 ;
        RECT 664.950 172.950 667.050 175.050 ;
        RECT 658.950 169.950 661.050 172.050 ;
        RECT 659.400 169.050 660.450 169.950 ;
        RECT 643.950 166.950 646.050 169.050 ;
        RECT 649.950 166.950 652.050 169.050 ;
        RECT 652.950 166.950 655.050 169.050 ;
        RECT 656.250 167.250 657.750 168.150 ;
        RECT 658.950 166.950 661.050 169.050 ;
        RECT 640.950 164.250 642.750 165.150 ;
        RECT 643.950 163.950 646.050 166.050 ;
        RECT 647.250 164.250 649.050 165.150 ;
        RECT 640.950 160.950 643.050 163.050 ;
        RECT 644.250 161.850 645.750 162.750 ;
        RECT 646.950 162.450 649.050 163.050 ;
        RECT 650.400 162.450 651.450 166.950 ;
        RECT 652.950 164.850 654.750 165.750 ;
        RECT 655.950 163.950 658.050 166.050 ;
        RECT 659.250 164.850 660.750 165.750 ;
        RECT 661.950 163.950 664.050 166.050 ;
        RECT 665.400 163.050 666.450 172.950 ;
        RECT 671.400 168.450 672.450 197.400 ;
        RECT 673.950 196.950 676.050 197.400 ;
        RECT 677.250 197.250 678.750 198.150 ;
        RECT 679.950 196.950 682.050 199.050 ;
        RECT 683.250 197.250 685.050 198.150 ;
        RECT 685.950 197.250 688.050 198.150 ;
        RECT 691.950 197.250 694.050 198.150 ;
        RECT 673.950 193.950 676.050 196.050 ;
        RECT 676.950 193.950 679.050 196.050 ;
        RECT 680.250 194.850 681.750 195.750 ;
        RECT 682.950 193.950 685.050 196.050 ;
        RECT 685.950 193.950 688.050 196.050 ;
        RECT 691.950 195.450 694.050 196.050 ;
        RECT 695.400 195.450 696.450 202.950 ;
        RECT 700.950 196.950 703.050 199.050 ;
        RECT 689.250 194.250 690.750 195.150 ;
        RECT 691.950 194.400 696.450 195.450 ;
        RECT 691.950 193.950 694.050 194.400 ;
        RECT 674.400 169.050 675.450 193.950 ;
        RECT 677.400 193.050 678.450 193.950 ;
        RECT 676.950 190.950 679.050 193.050 ;
        RECT 683.400 172.050 684.450 193.950 ;
        RECT 686.400 193.050 687.450 193.950 ;
        RECT 685.950 190.950 688.050 193.050 ;
        RECT 688.950 190.950 691.050 193.050 ;
        RECT 689.400 190.050 690.450 190.950 ;
        RECT 688.950 187.950 691.050 190.050 ;
        RECT 685.950 172.950 688.050 175.050 ;
        RECT 682.950 171.450 685.050 172.050 ;
        RECT 680.400 170.400 685.050 171.450 ;
        RECT 680.400 169.050 681.450 170.400 ;
        RECT 682.950 169.950 685.050 170.400 ;
        RECT 686.400 169.050 687.450 172.950 ;
        RECT 695.400 169.050 696.450 194.400 ;
        RECT 697.950 194.250 700.050 195.150 ;
        RECT 700.950 194.850 703.050 195.750 ;
        RECT 697.950 190.950 700.050 193.050 ;
        RECT 668.400 167.400 672.450 168.450 ;
        RECT 646.950 161.400 651.450 162.450 ;
        RECT 661.950 161.850 664.050 162.750 ;
        RECT 646.950 160.950 649.050 161.400 ;
        RECT 664.950 160.950 667.050 163.050 ;
        RECT 649.950 134.400 652.050 136.500 ;
        RECT 637.950 121.950 640.050 124.050 ;
        RECT 646.950 121.950 649.050 124.050 ;
        RECT 634.950 115.500 637.050 117.600 ;
        RECT 628.950 112.950 631.050 115.050 ;
        RECT 631.950 106.950 634.050 109.050 ;
        RECT 628.950 101.400 631.050 103.500 ;
        RECT 629.400 84.600 630.600 101.400 ;
        RECT 632.400 91.050 633.450 106.950 ;
        RECT 634.950 91.950 637.050 94.050 ;
        RECT 637.950 92.250 639.750 93.150 ;
        RECT 640.950 91.950 643.050 94.050 ;
        RECT 644.250 92.250 646.050 93.150 ;
        RECT 631.950 88.950 634.050 91.050 ;
        RECT 628.950 82.500 631.050 84.600 ;
        RECT 635.400 69.450 636.450 91.950 ;
        RECT 637.950 88.950 640.050 91.050 ;
        RECT 641.250 89.850 642.750 90.750 ;
        RECT 643.950 88.950 646.050 91.050 ;
        RECT 647.400 90.450 648.450 121.950 ;
        RECT 650.400 117.600 651.600 134.400 ;
        RECT 655.950 125.250 658.050 126.150 ;
        RECT 661.950 125.250 664.050 126.150 ;
        RECT 668.400 124.050 669.450 167.400 ;
        RECT 673.950 166.950 676.050 169.050 ;
        RECT 679.950 166.950 682.050 169.050 ;
        RECT 683.250 167.250 684.750 168.150 ;
        RECT 685.950 166.950 688.050 169.050 ;
        RECT 694.950 166.950 697.050 169.050 ;
        RECT 670.950 164.250 672.750 165.150 ;
        RECT 673.950 163.950 676.050 166.050 ;
        RECT 677.250 164.250 679.050 165.150 ;
        RECT 679.950 164.850 681.750 165.750 ;
        RECT 682.950 163.950 685.050 166.050 ;
        RECT 686.250 164.850 687.750 165.750 ;
        RECT 688.950 163.950 691.050 166.050 ;
        RECT 694.950 165.450 697.050 166.050 ;
        RECT 698.400 165.450 699.450 190.950 ;
        RECT 704.400 169.050 705.450 202.950 ;
        RECT 709.950 199.950 712.050 202.050 ;
        RECT 710.400 199.050 711.450 199.950 ;
        RECT 713.400 199.050 714.450 238.950 ;
        RECT 715.950 235.950 718.050 238.050 ;
        RECT 716.400 205.050 717.450 235.950 ;
        RECT 715.950 202.950 718.050 205.050 ;
        RECT 706.950 196.950 709.050 199.050 ;
        RECT 709.950 196.950 712.050 199.050 ;
        RECT 712.950 196.950 715.050 199.050 ;
        RECT 700.950 166.950 703.050 169.050 ;
        RECT 703.950 166.950 706.050 169.050 ;
        RECT 701.400 166.050 702.450 166.950 ;
        RECT 692.400 164.400 699.450 165.450 ;
        RECT 670.950 160.950 673.050 163.050 ;
        RECT 674.250 161.850 675.750 162.750 ;
        RECT 676.950 160.950 679.050 163.050 ;
        RECT 682.950 160.950 685.050 163.050 ;
        RECT 688.950 161.850 691.050 162.750 ;
        RECT 677.400 157.050 678.450 160.950 ;
        RECT 676.950 154.950 679.050 157.050 ;
        RECT 670.950 135.300 673.050 137.400 ;
        RECT 673.950 136.950 676.050 139.050 ;
        RECT 671.250 131.700 672.450 135.300 ;
        RECT 670.950 129.600 673.050 131.700 ;
        RECT 655.950 121.950 658.050 124.050 ;
        RECT 661.950 121.950 664.050 124.050 ;
        RECT 667.950 121.950 670.050 124.050 ;
        RECT 656.400 118.050 657.450 121.950 ;
        RECT 662.400 121.050 663.450 121.950 ;
        RECT 661.950 118.950 664.050 121.050 ;
        RECT 649.950 115.500 652.050 117.600 ;
        RECT 655.950 115.950 658.050 118.050 ;
        RECT 671.250 117.600 672.450 129.600 ;
        RECT 674.400 124.050 675.450 136.950 ;
        RECT 683.400 136.050 684.450 160.950 ;
        RECT 692.400 139.050 693.450 164.400 ;
        RECT 694.950 163.950 697.050 164.400 ;
        RECT 700.950 163.950 703.050 166.050 ;
        RECT 704.250 164.250 706.050 165.150 ;
        RECT 694.950 161.850 696.750 162.750 ;
        RECT 697.950 160.950 700.050 163.050 ;
        RECT 701.250 161.850 702.750 162.750 ;
        RECT 703.950 160.950 706.050 163.050 ;
        RECT 697.950 158.850 700.050 159.750 ;
        RECT 700.950 157.950 703.050 160.050 ;
        RECT 691.950 136.950 694.050 139.050 ;
        RECT 697.950 136.950 700.050 139.050 ;
        RECT 682.950 133.950 685.050 136.050 ;
        RECT 683.400 127.050 684.450 133.950 ;
        RECT 691.950 130.950 694.050 133.050 ;
        RECT 688.950 128.250 691.050 129.150 ;
        RECT 679.950 125.250 681.750 126.150 ;
        RECT 682.950 124.950 685.050 127.050 ;
        RECT 688.950 126.450 691.050 127.050 ;
        RECT 692.400 126.450 693.450 130.950 ;
        RECT 698.400 127.050 699.450 136.950 ;
        RECT 701.400 130.050 702.450 157.950 ;
        RECT 704.400 157.050 705.450 160.950 ;
        RECT 703.950 154.950 706.050 157.050 ;
        RECT 700.950 127.950 703.050 130.050 ;
        RECT 703.950 128.250 706.050 129.150 ;
        RECT 686.250 125.250 687.750 126.150 ;
        RECT 688.950 125.400 693.450 126.450 ;
        RECT 688.950 124.950 691.050 125.400 ;
        RECT 694.950 125.250 696.750 126.150 ;
        RECT 697.950 124.950 700.050 127.050 ;
        RECT 703.950 126.450 706.050 127.050 ;
        RECT 707.400 126.450 708.450 196.950 ;
        RECT 709.950 194.850 712.050 195.750 ;
        RECT 712.950 194.250 715.050 195.150 ;
        RECT 712.950 169.950 715.050 172.050 ;
        RECT 709.950 166.950 712.050 169.050 ;
        RECT 710.400 133.050 711.450 166.950 ;
        RECT 713.400 139.050 714.450 169.950 ;
        RECT 712.950 136.950 715.050 139.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 709.950 130.950 712.050 133.050 ;
        RECT 701.250 125.250 702.750 126.150 ;
        RECT 703.950 125.400 708.450 126.450 ;
        RECT 703.950 124.950 706.050 125.400 ;
        RECT 673.950 121.950 676.050 124.050 ;
        RECT 679.950 121.950 682.050 124.050 ;
        RECT 683.250 122.850 684.750 123.750 ;
        RECT 685.950 123.450 688.050 124.050 ;
        RECT 685.950 122.400 690.450 123.450 ;
        RECT 685.950 121.950 688.050 122.400 ;
        RECT 673.950 119.850 676.050 120.750 ;
        RECT 670.950 115.500 673.050 117.600 ;
        RECT 667.950 112.950 670.050 115.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 649.950 92.250 651.750 93.150 ;
        RECT 652.950 91.950 655.050 94.050 ;
        RECT 656.250 92.250 658.050 93.150 ;
        RECT 649.950 90.450 652.050 91.050 ;
        RECT 647.400 89.400 652.050 90.450 ;
        RECT 653.250 89.850 654.750 90.750 ;
        RECT 655.950 90.450 658.050 91.050 ;
        RECT 659.400 90.450 660.450 100.950 ;
        RECT 668.400 97.050 669.450 112.950 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 674.400 97.050 675.450 100.950 ;
        RECT 667.950 94.950 670.050 97.050 ;
        RECT 671.250 95.250 672.750 96.150 ;
        RECT 673.950 94.950 676.050 97.050 ;
        RECT 664.950 91.950 667.050 94.050 ;
        RECT 668.250 92.850 669.750 93.750 ;
        RECT 670.950 91.950 673.050 94.050 ;
        RECT 674.250 92.850 676.050 93.750 ;
        RECT 649.950 88.950 652.050 89.400 ;
        RECT 655.950 89.400 660.450 90.450 ;
        RECT 664.950 89.850 667.050 90.750 ;
        RECT 655.950 88.950 658.050 89.400 ;
        RECT 635.400 68.400 639.450 69.450 ;
        RECT 634.950 62.400 637.050 64.500 ;
        RECT 628.950 53.250 631.050 54.150 ;
        RECT 622.950 50.400 627.450 51.450 ;
        RECT 622.950 49.950 625.050 50.400 ;
        RECT 628.950 49.950 631.050 52.050 ;
        RECT 619.950 46.950 622.050 49.050 ;
        RECT 613.950 43.500 616.050 45.600 ;
        RECT 616.950 43.950 619.050 46.050 ;
        RECT 604.950 37.950 607.050 40.050 ;
        RECT 598.950 25.950 601.050 28.050 ;
        RECT 601.950 25.950 604.050 28.050 ;
        RECT 605.400 25.050 606.450 37.950 ;
        RECT 613.950 27.450 616.050 28.050 ;
        RECT 608.400 26.400 616.050 27.450 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 602.250 23.850 603.750 24.750 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 608.400 22.050 609.450 26.400 ;
        RECT 613.950 25.950 616.050 26.400 ;
        RECT 617.400 25.050 618.450 43.950 ;
        RECT 629.400 43.050 630.450 49.950 ;
        RECT 635.400 45.600 636.600 62.400 ;
        RECT 638.400 52.050 639.450 68.400 ;
        RECT 644.400 64.050 645.450 88.950 ;
        RECT 671.400 79.050 672.450 91.950 ;
        RECT 670.950 76.950 673.050 79.050 ;
        RECT 680.400 64.050 681.450 121.950 ;
        RECT 682.950 101.400 685.050 103.500 ;
        RECT 683.400 84.600 684.600 101.400 ;
        RECT 689.400 97.050 690.450 122.400 ;
        RECT 694.950 121.950 697.050 124.050 ;
        RECT 698.250 122.850 699.750 123.750 ;
        RECT 700.950 123.450 703.050 124.050 ;
        RECT 700.950 122.400 705.450 123.450 ;
        RECT 700.950 121.950 703.050 122.400 ;
        RECT 694.950 118.950 697.050 121.050 ;
        RECT 700.950 118.950 703.050 121.050 ;
        RECT 695.400 97.050 696.450 118.950 ;
        RECT 701.400 97.050 702.450 118.950 ;
        RECT 704.400 118.050 705.450 122.400 ;
        RECT 703.950 115.950 706.050 118.050 ;
        RECT 703.950 101.400 706.050 103.500 ;
        RECT 688.950 94.950 691.050 97.050 ;
        RECT 694.950 96.450 697.050 97.050 ;
        RECT 692.400 95.400 697.050 96.450 ;
        RECT 688.950 92.850 691.050 93.750 ;
        RECT 682.950 82.500 685.050 84.600 ;
        RECT 643.950 61.950 646.050 64.050 ;
        RECT 670.950 61.950 673.050 64.050 ;
        RECT 679.950 61.950 682.050 64.050 ;
        RECT 685.950 63.300 688.050 65.400 ;
        RECT 640.950 58.950 643.050 61.050 ;
        RECT 652.950 58.950 655.050 61.050 ;
        RECT 637.950 49.950 640.050 52.050 ;
        RECT 634.950 43.500 637.050 45.600 ;
        RECT 628.950 40.950 631.050 43.050 ;
        RECT 626.400 29.400 633.450 30.450 ;
        RECT 626.400 28.050 627.450 29.400 ;
        RECT 625.950 25.950 628.050 28.050 ;
        RECT 628.950 25.950 631.050 28.050 ;
        RECT 632.400 27.450 633.450 29.400 ;
        RECT 632.400 26.400 636.450 27.450 ;
        RECT 626.400 25.050 627.450 25.950 ;
        RECT 635.400 25.050 636.450 26.400 ;
        RECT 641.400 25.050 642.450 58.950 ;
        RECT 653.400 58.050 654.450 58.950 ;
        RECT 646.950 55.950 649.050 58.050 ;
        RECT 650.250 56.250 651.750 57.150 ;
        RECT 652.950 55.950 655.050 58.050 ;
        RECT 655.950 55.950 658.050 58.050 ;
        RECT 658.950 56.250 661.050 57.150 ;
        RECT 646.950 53.850 648.750 54.750 ;
        RECT 649.950 52.950 652.050 55.050 ;
        RECT 653.250 53.850 655.050 54.750 ;
        RECT 656.400 34.050 657.450 55.950 ;
        RECT 658.950 52.950 661.050 55.050 ;
        RECT 662.250 53.250 663.750 54.150 ;
        RECT 664.950 52.950 667.050 55.050 ;
        RECT 668.250 53.250 670.050 54.150 ;
        RECT 659.400 52.050 660.450 52.950 ;
        RECT 658.950 49.950 661.050 52.050 ;
        RECT 661.950 49.950 664.050 52.050 ;
        RECT 665.250 50.850 666.750 51.750 ;
        RECT 667.950 51.450 670.050 52.050 ;
        RECT 671.400 51.450 672.450 61.950 ;
        RECT 686.550 59.700 687.750 63.300 ;
        RECT 685.950 57.600 688.050 59.700 ;
        RECT 673.950 52.950 676.050 55.050 ;
        RECT 667.950 50.400 672.450 51.450 ;
        RECT 673.950 50.850 676.050 51.750 ;
        RECT 682.950 51.450 685.050 52.050 ;
        RECT 667.950 49.950 670.050 50.400 ;
        RECT 676.950 50.250 679.050 51.150 ;
        RECT 680.400 50.400 685.050 51.450 ;
        RECT 662.400 46.050 663.450 49.950 ;
        RECT 670.950 46.950 673.050 49.050 ;
        RECT 676.950 48.450 679.050 49.050 ;
        RECT 680.400 48.450 681.450 50.400 ;
        RECT 682.950 49.950 685.050 50.400 ;
        RECT 676.950 47.400 681.450 48.450 ;
        RECT 682.950 47.850 685.050 48.750 ;
        RECT 676.950 46.950 679.050 47.400 ;
        RECT 661.950 43.950 664.050 46.050 ;
        RECT 655.950 31.950 658.050 34.050 ;
        RECT 649.950 25.950 652.050 28.050 ;
        RECT 610.950 22.950 613.050 25.050 ;
        RECT 614.250 23.850 615.750 24.750 ;
        RECT 616.950 22.950 619.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 629.250 23.850 630.750 24.750 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 634.950 22.950 637.050 25.050 ;
        RECT 638.250 23.250 639.750 24.150 ;
        RECT 640.950 22.950 643.050 25.050 ;
        RECT 598.950 20.850 601.050 21.750 ;
        RECT 604.950 20.850 607.050 21.750 ;
        RECT 607.950 19.950 610.050 22.050 ;
        RECT 610.950 20.850 613.050 21.750 ;
        RECT 616.950 20.850 619.050 21.750 ;
        RECT 625.950 20.850 628.050 21.750 ;
        RECT 631.950 20.850 634.050 21.750 ;
        RECT 634.950 20.850 636.750 21.750 ;
        RECT 637.950 19.950 640.050 22.050 ;
        RECT 641.250 20.850 642.750 21.750 ;
        RECT 643.950 19.950 646.050 22.050 ;
        RECT 586.950 16.950 589.050 19.050 ;
        RECT 592.950 17.850 595.050 18.750 ;
        RECT 595.950 16.950 598.050 19.050 ;
        RECT 643.950 17.850 646.050 18.750 ;
        RECT 650.400 18.450 651.450 25.950 ;
        RECT 656.400 22.050 657.450 31.950 ;
        RECT 661.950 25.950 664.050 28.050 ;
        RECT 667.950 25.950 670.050 28.050 ;
        RECT 652.950 20.250 654.750 21.150 ;
        RECT 655.950 19.950 658.050 22.050 ;
        RECT 659.250 20.250 661.050 21.150 ;
        RECT 652.950 18.450 655.050 19.050 ;
        RECT 650.400 17.400 655.050 18.450 ;
        RECT 656.250 17.850 657.750 18.750 ;
        RECT 658.950 18.450 661.050 19.050 ;
        RECT 662.400 18.450 663.450 25.950 ;
        RECT 671.400 25.050 672.450 46.950 ;
        RECT 686.550 45.600 687.750 57.600 ;
        RECT 692.400 51.450 693.450 95.400 ;
        RECT 694.950 94.950 697.050 95.400 ;
        RECT 697.950 94.950 700.050 97.050 ;
        RECT 700.950 94.950 703.050 97.050 ;
        RECT 694.950 92.850 697.050 93.750 ;
        RECT 694.950 53.250 697.050 54.150 ;
        RECT 694.950 51.450 697.050 52.050 ;
        RECT 692.400 50.400 697.050 51.450 ;
        RECT 694.950 49.950 697.050 50.400 ;
        RECT 685.950 43.500 688.050 45.600 ;
        RECT 676.950 28.950 679.050 31.050 ;
        RECT 677.400 28.050 678.450 28.950 ;
        RECT 673.950 25.950 676.050 28.050 ;
        RECT 676.950 25.950 679.050 28.050 ;
        RECT 691.950 25.950 694.050 28.050 ;
        RECT 698.400 27.450 699.450 94.950 ;
        RECT 704.250 89.400 705.450 101.400 ;
        RECT 706.950 98.250 709.050 99.150 ;
        RECT 706.950 94.950 709.050 97.050 ;
        RECT 703.950 87.300 706.050 89.400 ;
        RECT 704.250 83.700 705.450 87.300 ;
        RECT 703.950 81.600 706.050 83.700 ;
        RECT 703.950 76.950 706.050 79.050 ;
        RECT 700.950 53.250 703.050 54.150 ;
        RECT 700.950 49.950 703.050 52.050 ;
        RECT 701.400 46.050 702.450 49.950 ;
        RECT 700.950 43.950 703.050 46.050 ;
        RECT 704.400 39.450 705.450 76.950 ;
        RECT 706.950 62.400 709.050 64.500 ;
        RECT 707.400 45.600 708.600 62.400 ;
        RECT 706.950 43.500 709.050 45.600 ;
        RECT 704.400 38.400 708.450 39.450 ;
        RECT 700.950 27.450 703.050 28.050 ;
        RECT 698.400 26.400 703.050 27.450 ;
        RECT 700.950 25.950 703.050 26.400 ;
        RECT 677.400 25.050 678.450 25.950 ;
        RECT 664.950 23.250 667.050 24.150 ;
        RECT 667.950 23.850 670.050 24.750 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 674.250 23.850 675.750 24.750 ;
        RECT 676.950 22.950 679.050 25.050 ;
        RECT 679.950 22.950 682.050 25.050 ;
        RECT 664.950 19.950 667.050 22.050 ;
        RECT 670.950 20.850 673.050 21.750 ;
        RECT 676.950 20.850 679.050 21.750 ;
        RECT 652.950 16.950 655.050 17.400 ;
        RECT 658.950 17.400 663.450 18.450 ;
        RECT 658.950 16.950 661.050 17.400 ;
        RECT 665.400 16.050 666.450 19.950 ;
        RECT 680.400 18.450 681.450 22.950 ;
        RECT 682.950 20.250 684.750 21.150 ;
        RECT 685.950 19.950 688.050 22.050 ;
        RECT 689.250 20.250 691.050 21.150 ;
        RECT 682.950 18.450 685.050 19.050 ;
        RECT 680.400 17.400 685.050 18.450 ;
        RECT 686.250 17.850 687.750 18.750 ;
        RECT 688.950 18.450 691.050 19.050 ;
        RECT 692.400 18.450 693.450 25.950 ;
        RECT 697.950 23.250 700.050 24.150 ;
        RECT 700.950 23.850 703.050 24.750 ;
        RECT 707.400 22.050 708.450 38.400 ;
        RECT 713.400 22.050 714.450 133.950 ;
        RECT 697.950 19.950 700.050 22.050 ;
        RECT 703.950 20.250 705.750 21.150 ;
        RECT 706.950 19.950 709.050 22.050 ;
        RECT 710.250 20.250 712.050 21.150 ;
        RECT 712.950 19.950 715.050 22.050 ;
        RECT 682.950 16.950 685.050 17.400 ;
        RECT 688.950 17.400 693.450 18.450 ;
        RECT 688.950 16.950 691.050 17.400 ;
        RECT 703.950 16.950 706.050 19.050 ;
        RECT 707.250 17.850 708.750 18.750 ;
        RECT 709.950 16.950 712.050 19.050 ;
        RECT 710.400 16.050 711.450 16.950 ;
        RECT 664.950 13.950 667.050 16.050 ;
        RECT 709.950 13.950 712.050 16.050 ;
        RECT 517.950 9.600 520.050 11.700 ;
        RECT 544.950 9.600 547.050 11.700 ;
        RECT 565.950 10.500 568.050 12.600 ;
      LAYER metal3 ;
        RECT 184.950 684.600 187.050 685.050 ;
        RECT 229.950 684.600 232.050 685.050 ;
        RECT 184.950 683.400 232.050 684.600 ;
        RECT 184.950 682.950 187.050 683.400 ;
        RECT 229.950 682.950 232.050 683.400 ;
        RECT 16.950 681.600 19.050 682.050 ;
        RECT 28.950 681.600 31.050 682.050 ;
        RECT 16.950 680.400 31.050 681.600 ;
        RECT 16.950 679.950 19.050 680.400 ;
        RECT 28.950 679.950 31.050 680.400 ;
        RECT 133.950 681.600 136.050 682.050 ;
        RECT 193.950 681.600 196.050 682.050 ;
        RECT 133.950 680.400 196.050 681.600 ;
        RECT 133.950 679.950 136.050 680.400 ;
        RECT 193.950 679.950 196.050 680.400 ;
        RECT 217.950 681.600 220.050 682.050 ;
        RECT 244.950 681.600 247.050 682.050 ;
        RECT 217.950 680.400 247.050 681.600 ;
        RECT 217.950 679.950 220.050 680.400 ;
        RECT 244.950 679.950 247.050 680.400 ;
        RECT 340.950 681.600 343.050 682.050 ;
        RECT 349.950 681.600 352.050 682.050 ;
        RECT 340.950 680.400 352.050 681.600 ;
        RECT 340.950 679.950 343.050 680.400 ;
        RECT 349.950 679.950 352.050 680.400 ;
        RECT 499.950 681.600 502.050 682.050 ;
        RECT 514.950 681.600 517.050 682.050 ;
        RECT 499.950 680.400 517.050 681.600 ;
        RECT 499.950 679.950 502.050 680.400 ;
        RECT 514.950 679.950 517.050 680.400 ;
        RECT 4.950 678.600 7.050 679.050 ;
        RECT 73.950 678.600 76.050 679.050 ;
        RECT 4.950 677.400 76.050 678.600 ;
        RECT 4.950 676.950 7.050 677.400 ;
        RECT 73.950 676.950 76.050 677.400 ;
        RECT 106.950 678.600 109.050 679.050 ;
        RECT 214.950 678.600 217.050 679.050 ;
        RECT 241.950 678.600 244.050 679.050 ;
        RECT 253.950 678.600 256.050 679.050 ;
        RECT 271.950 678.600 274.050 679.050 ;
        RECT 106.950 677.400 274.050 678.600 ;
        RECT 106.950 676.950 109.050 677.400 ;
        RECT 214.950 676.950 217.050 677.400 ;
        RECT 241.950 676.950 244.050 677.400 ;
        RECT 253.950 676.950 256.050 677.400 ;
        RECT 271.950 676.950 274.050 677.400 ;
        RECT 292.950 678.600 295.050 679.050 ;
        RECT 301.950 678.600 304.050 679.050 ;
        RECT 292.950 677.400 304.050 678.600 ;
        RECT 292.950 676.950 295.050 677.400 ;
        RECT 301.950 676.950 304.050 677.400 ;
        RECT 307.950 678.600 310.050 679.050 ;
        RECT 343.950 678.600 346.050 679.050 ;
        RECT 307.950 677.400 346.050 678.600 ;
        RECT 307.950 676.950 310.050 677.400 ;
        RECT 343.950 676.950 346.050 677.400 ;
        RECT 451.950 678.600 454.050 679.050 ;
        RECT 457.950 678.600 460.050 679.050 ;
        RECT 451.950 677.400 460.050 678.600 ;
        RECT 451.950 676.950 454.050 677.400 ;
        RECT 457.950 676.950 460.050 677.400 ;
        RECT 463.950 678.600 466.050 679.050 ;
        RECT 475.950 678.600 478.050 679.050 ;
        RECT 463.950 677.400 478.050 678.600 ;
        RECT 463.950 676.950 466.050 677.400 ;
        RECT 475.950 676.950 478.050 677.400 ;
        RECT 484.950 678.600 487.050 679.050 ;
        RECT 523.950 678.600 526.050 679.050 ;
        RECT 484.950 677.400 526.050 678.600 ;
        RECT 484.950 676.950 487.050 677.400 ;
        RECT 523.950 676.950 526.050 677.400 ;
        RECT 595.950 678.600 598.050 679.050 ;
        RECT 691.950 678.600 694.050 679.050 ;
        RECT 595.950 677.400 694.050 678.600 ;
        RECT 595.950 676.950 598.050 677.400 ;
        RECT 691.950 676.950 694.050 677.400 ;
        RECT 10.950 675.600 13.050 676.050 ;
        RECT 25.950 675.600 28.050 676.050 ;
        RECT 10.950 674.400 28.050 675.600 ;
        RECT 10.950 673.950 13.050 674.400 ;
        RECT 25.950 673.950 28.050 674.400 ;
        RECT 55.950 675.600 58.050 676.050 ;
        RECT 64.950 675.600 67.050 676.050 ;
        RECT 55.950 674.400 67.050 675.600 ;
        RECT 55.950 673.950 58.050 674.400 ;
        RECT 64.950 673.950 67.050 674.400 ;
        RECT 82.950 675.600 85.050 676.050 ;
        RECT 97.950 675.600 100.050 676.050 ;
        RECT 157.950 675.600 160.050 676.050 ;
        RECT 82.950 674.400 96.600 675.600 ;
        RECT 82.950 673.950 85.050 674.400 ;
        RECT 25.950 672.600 28.050 673.050 ;
        RECT 31.950 672.600 34.050 673.050 ;
        RECT 25.950 671.400 34.050 672.600 ;
        RECT 25.950 670.950 28.050 671.400 ;
        RECT 31.950 670.950 34.050 671.400 ;
        RECT 58.950 672.600 61.050 673.050 ;
        RECT 70.950 672.600 73.050 673.050 ;
        RECT 58.950 671.400 66.600 672.600 ;
        RECT 58.950 670.950 61.050 671.400 ;
        RECT 13.950 669.600 16.050 670.050 ;
        RECT 22.950 669.600 25.050 670.050 ;
        RECT 34.950 669.600 37.050 670.050 ;
        RECT 13.950 668.400 37.050 669.600 ;
        RECT 13.950 667.950 16.050 668.400 ;
        RECT 22.950 667.950 25.050 668.400 ;
        RECT 34.950 667.950 37.050 668.400 ;
        RECT 37.950 669.600 40.050 670.050 ;
        RECT 46.950 669.600 49.050 670.050 ;
        RECT 37.950 668.400 49.050 669.600 ;
        RECT 37.950 667.950 40.050 668.400 ;
        RECT 46.950 667.950 49.050 668.400 ;
        RECT 52.950 669.600 55.050 670.050 ;
        RECT 61.950 669.600 64.050 670.050 ;
        RECT 52.950 668.400 64.050 669.600 ;
        RECT 65.400 669.600 66.600 671.400 ;
        RECT 70.950 671.400 90.600 672.600 ;
        RECT 70.950 670.950 73.050 671.400 ;
        RECT 67.950 669.600 70.050 670.050 ;
        RECT 73.950 669.600 76.050 670.050 ;
        RECT 65.400 668.400 76.050 669.600 ;
        RECT 52.950 667.950 55.050 668.400 ;
        RECT 61.950 667.950 64.050 668.400 ;
        RECT 67.950 667.950 70.050 668.400 ;
        RECT 73.950 667.950 76.050 668.400 ;
        RECT 25.950 664.950 28.050 667.050 ;
        RECT 40.950 666.600 43.050 667.050 ;
        RECT 55.950 666.600 58.050 667.050 ;
        RECT 76.950 666.600 79.050 667.050 ;
        RECT 79.950 666.600 82.050 667.050 ;
        RECT 40.950 665.400 58.050 666.600 ;
        RECT 74.400 665.400 82.050 666.600 ;
        RECT 40.950 664.950 43.050 665.400 ;
        RECT 55.950 664.950 58.050 665.400 ;
        RECT 76.950 664.950 79.050 665.400 ;
        RECT 79.950 664.950 82.050 665.400 ;
        RECT 13.950 663.600 16.050 664.050 ;
        RECT 22.950 663.600 25.050 664.050 ;
        RECT 13.950 662.400 25.050 663.600 ;
        RECT 26.400 663.600 27.600 664.950 ;
        RECT 28.950 663.600 31.050 664.050 ;
        RECT 26.400 662.400 31.050 663.600 ;
        RECT 89.400 663.600 90.600 671.400 ;
        RECT 91.950 670.950 94.050 673.050 ;
        RECT 95.400 672.600 96.600 674.400 ;
        RECT 97.950 674.400 160.050 675.600 ;
        RECT 97.950 673.950 100.050 674.400 ;
        RECT 157.950 673.950 160.050 674.400 ;
        RECT 160.950 675.600 163.050 676.050 ;
        RECT 166.950 675.600 169.050 676.050 ;
        RECT 160.950 674.400 169.050 675.600 ;
        RECT 160.950 673.950 163.050 674.400 ;
        RECT 166.950 673.950 169.050 674.400 ;
        RECT 169.950 675.600 172.050 676.050 ;
        RECT 190.950 675.600 193.050 676.050 ;
        RECT 169.950 674.400 193.050 675.600 ;
        RECT 169.950 673.950 172.050 674.400 ;
        RECT 190.950 673.950 193.050 674.400 ;
        RECT 196.950 675.600 199.050 676.050 ;
        RECT 202.950 675.600 205.050 676.050 ;
        RECT 217.950 675.600 220.050 676.050 ;
        RECT 196.950 674.400 205.050 675.600 ;
        RECT 196.950 673.950 199.050 674.400 ;
        RECT 202.950 673.950 205.050 674.400 ;
        RECT 206.400 674.400 220.050 675.600 ;
        RECT 112.950 672.600 115.050 673.050 ;
        RECT 95.400 671.400 115.050 672.600 ;
        RECT 112.950 670.950 115.050 671.400 ;
        RECT 115.950 672.600 118.050 673.050 ;
        RECT 124.950 672.600 127.050 673.050 ;
        RECT 115.950 671.400 127.050 672.600 ;
        RECT 115.950 670.950 118.050 671.400 ;
        RECT 124.950 670.950 127.050 671.400 ;
        RECT 127.950 672.600 130.050 673.050 ;
        RECT 148.950 672.600 151.050 673.050 ;
        RECT 172.950 672.600 175.050 673.050 ;
        RECT 175.950 672.600 178.050 673.050 ;
        RECT 199.950 672.600 202.050 673.050 ;
        RECT 206.400 672.600 207.600 674.400 ;
        RECT 217.950 673.950 220.050 674.400 ;
        RECT 232.950 675.600 235.050 676.050 ;
        RECT 265.950 675.600 268.050 676.050 ;
        RECT 286.950 675.600 289.050 676.050 ;
        RECT 325.950 675.600 328.050 676.050 ;
        RECT 358.950 675.600 361.050 676.050 ;
        RECT 370.950 675.600 373.050 676.050 ;
        RECT 232.950 674.400 268.050 675.600 ;
        RECT 232.950 673.950 235.050 674.400 ;
        RECT 265.950 673.950 268.050 674.400 ;
        RECT 284.400 674.400 328.050 675.600 ;
        RECT 127.950 671.400 147.600 672.600 ;
        RECT 127.950 670.950 130.050 671.400 ;
        RECT 92.400 667.050 93.600 670.950 ;
        RECT 100.950 667.950 103.050 670.050 ;
        RECT 103.950 669.600 106.050 670.050 ;
        RECT 112.950 669.600 115.050 670.050 ;
        RECT 103.950 668.400 115.050 669.600 ;
        RECT 103.950 667.950 106.050 668.400 ;
        RECT 112.950 667.950 115.050 668.400 ;
        RECT 118.950 667.950 121.050 670.050 ;
        RECT 121.950 667.950 124.050 670.050 ;
        RECT 127.950 669.600 130.050 670.050 ;
        RECT 139.950 669.600 142.050 670.050 ;
        RECT 127.950 668.400 142.050 669.600 ;
        RECT 146.400 669.600 147.600 671.400 ;
        RECT 148.950 671.400 165.600 672.600 ;
        RECT 148.950 670.950 151.050 671.400 ;
        RECT 164.400 670.050 165.600 671.400 ;
        RECT 172.950 671.400 202.050 672.600 ;
        RECT 172.950 670.950 175.050 671.400 ;
        RECT 175.950 670.950 178.050 671.400 ;
        RECT 199.950 670.950 202.050 671.400 ;
        RECT 203.400 671.400 207.600 672.600 ;
        RECT 208.950 672.600 211.050 673.050 ;
        RECT 223.950 672.600 226.050 673.050 ;
        RECT 235.950 672.600 238.050 673.050 ;
        RECT 284.400 672.600 285.600 674.400 ;
        RECT 286.950 673.950 289.050 674.400 ;
        RECT 325.950 673.950 328.050 674.400 ;
        RECT 329.400 674.400 373.050 675.600 ;
        RECT 208.950 671.400 222.600 672.600 ;
        RECT 154.950 669.600 157.050 670.050 ;
        RECT 163.950 669.600 166.050 670.050 ;
        RECT 178.950 669.600 181.050 670.050 ;
        RECT 146.400 668.400 162.600 669.600 ;
        RECT 127.950 667.950 130.050 668.400 ;
        RECT 139.950 667.950 142.050 668.400 ;
        RECT 154.950 667.950 157.050 668.400 ;
        RECT 91.950 664.950 94.050 667.050 ;
        RECT 97.950 666.600 100.050 667.050 ;
        RECT 101.400 666.600 102.600 667.950 ;
        RECT 97.950 665.400 102.600 666.600 ;
        RECT 97.950 664.950 100.050 665.400 ;
        RECT 94.950 663.600 97.050 664.050 ;
        RECT 89.400 662.400 97.050 663.600 ;
        RECT 13.950 661.950 16.050 662.400 ;
        RECT 22.950 661.950 25.050 662.400 ;
        RECT 28.950 661.950 31.050 662.400 ;
        RECT 94.950 661.950 97.050 662.400 ;
        RECT 106.950 663.600 109.050 664.050 ;
        RECT 119.400 663.600 120.600 667.950 ;
        RECT 122.400 664.050 123.600 667.950 ;
        RECT 124.950 666.600 127.050 667.050 ;
        RECT 130.950 666.600 133.050 667.050 ;
        RECT 142.950 666.600 145.050 667.050 ;
        RECT 151.950 666.600 154.050 667.050 ;
        RECT 124.950 665.400 129.600 666.600 ;
        RECT 124.950 664.950 127.050 665.400 ;
        RECT 128.400 664.050 129.600 665.400 ;
        RECT 130.950 665.400 135.600 666.600 ;
        RECT 130.950 664.950 133.050 665.400 ;
        RECT 106.950 662.400 120.600 663.600 ;
        RECT 106.950 661.950 109.050 662.400 ;
        RECT 121.950 661.950 124.050 664.050 ;
        RECT 127.950 661.950 130.050 664.050 ;
        RECT 7.950 660.600 10.050 661.050 ;
        RECT 16.950 660.600 19.050 661.050 ;
        RECT 25.950 660.600 28.050 661.050 ;
        RECT 7.950 659.400 28.050 660.600 ;
        RECT 7.950 658.950 10.050 659.400 ;
        RECT 16.950 658.950 19.050 659.400 ;
        RECT 25.950 658.950 28.050 659.400 ;
        RECT 49.950 660.600 52.050 661.050 ;
        RECT 103.950 660.600 106.050 661.050 ;
        RECT 49.950 659.400 106.050 660.600 ;
        RECT 134.400 660.600 135.600 665.400 ;
        RECT 142.950 665.400 154.050 666.600 ;
        RECT 161.400 666.600 162.600 668.400 ;
        RECT 163.950 668.400 181.050 669.600 ;
        RECT 163.950 667.950 166.050 668.400 ;
        RECT 178.950 667.950 181.050 668.400 ;
        RECT 190.950 669.600 193.050 670.050 ;
        RECT 203.400 669.600 204.600 671.400 ;
        RECT 208.950 670.950 211.050 671.400 ;
        RECT 190.950 668.400 204.600 669.600 ;
        RECT 190.950 667.950 193.050 668.400 ;
        RECT 205.950 667.950 208.050 670.050 ;
        RECT 221.400 669.600 222.600 671.400 ;
        RECT 223.950 671.400 285.600 672.600 ;
        RECT 298.950 672.600 301.050 673.050 ;
        RECT 329.400 672.600 330.600 674.400 ;
        RECT 358.950 673.950 361.050 674.400 ;
        RECT 370.950 673.950 373.050 674.400 ;
        RECT 376.950 673.950 379.050 676.050 ;
        RECT 439.950 675.600 442.050 676.050 ;
        RECT 448.950 675.600 451.050 676.050 ;
        RECT 466.950 675.600 469.050 676.050 ;
        RECT 469.950 675.600 472.050 676.050 ;
        RECT 439.950 674.400 472.050 675.600 ;
        RECT 439.950 673.950 442.050 674.400 ;
        RECT 448.950 673.950 451.050 674.400 ;
        RECT 466.950 673.950 469.050 674.400 ;
        RECT 469.950 673.950 472.050 674.400 ;
        RECT 475.950 675.600 478.050 676.050 ;
        RECT 511.950 675.600 514.050 676.050 ;
        RECT 622.950 675.600 625.050 676.050 ;
        RECT 649.950 675.600 652.050 676.050 ;
        RECT 475.950 674.400 519.600 675.600 ;
        RECT 475.950 673.950 478.050 674.400 ;
        RECT 511.950 673.950 514.050 674.400 ;
        RECT 298.950 671.400 330.600 672.600 ;
        RECT 331.950 672.600 334.050 673.050 ;
        RECT 331.950 671.400 348.600 672.600 ;
        RECT 223.950 670.950 226.050 671.400 ;
        RECT 235.950 670.950 238.050 671.400 ;
        RECT 298.950 670.950 301.050 671.400 ;
        RECT 331.950 670.950 334.050 671.400 ;
        RECT 347.400 670.050 348.600 671.400 ;
        RECT 355.950 670.950 358.050 673.050 ;
        RECT 364.950 672.600 367.050 673.050 ;
        RECT 377.400 672.600 378.600 673.950 ;
        RECT 518.400 673.050 519.600 674.400 ;
        RECT 622.950 674.400 652.050 675.600 ;
        RECT 622.950 673.950 625.050 674.400 ;
        RECT 649.950 673.950 652.050 674.400 ;
        RECT 364.950 671.400 378.600 672.600 ;
        RECT 364.950 670.950 367.050 671.400 ;
        RECT 391.950 670.950 394.050 673.050 ;
        RECT 397.950 672.600 400.050 673.050 ;
        RECT 418.950 672.600 421.050 673.050 ;
        RECT 490.950 672.600 493.050 673.050 ;
        RECT 502.950 672.600 505.050 673.050 ;
        RECT 505.950 672.600 508.050 673.050 ;
        RECT 397.950 671.400 421.050 672.600 ;
        RECT 397.950 670.950 400.050 671.400 ;
        RECT 418.950 670.950 421.050 671.400 ;
        RECT 452.400 671.400 471.600 672.600 ;
        RECT 232.950 669.600 235.050 670.050 ;
        RECT 221.400 668.400 235.050 669.600 ;
        RECT 232.950 667.950 235.050 668.400 ;
        RECT 238.950 669.600 241.050 670.050 ;
        RECT 247.950 669.600 250.050 670.050 ;
        RECT 238.950 668.400 250.050 669.600 ;
        RECT 238.950 667.950 241.050 668.400 ;
        RECT 247.950 667.950 250.050 668.400 ;
        RECT 283.950 669.600 286.050 670.050 ;
        RECT 301.950 669.600 304.050 670.050 ;
        RECT 283.950 668.400 304.050 669.600 ;
        RECT 283.950 667.950 286.050 668.400 ;
        RECT 301.950 667.950 304.050 668.400 ;
        RECT 319.950 669.600 322.050 670.050 ;
        RECT 328.950 669.600 331.050 670.050 ;
        RECT 319.950 668.400 331.050 669.600 ;
        RECT 319.950 667.950 322.050 668.400 ;
        RECT 328.950 667.950 331.050 668.400 ;
        RECT 346.950 667.950 349.050 670.050 ;
        RECT 169.950 666.600 172.050 667.050 ;
        RECT 161.400 665.400 172.050 666.600 ;
        RECT 142.950 664.950 145.050 665.400 ;
        RECT 151.950 664.950 154.050 665.400 ;
        RECT 169.950 664.950 172.050 665.400 ;
        RECT 187.950 666.600 190.050 667.050 ;
        RECT 206.400 666.600 207.600 667.950 ;
        RECT 187.950 665.400 207.600 666.600 ;
        RECT 226.950 666.600 229.050 667.050 ;
        RECT 253.950 666.600 256.050 667.050 ;
        RECT 226.950 665.400 256.050 666.600 ;
        RECT 187.950 664.950 190.050 665.400 ;
        RECT 226.950 664.950 229.050 665.400 ;
        RECT 253.950 664.950 256.050 665.400 ;
        RECT 274.950 666.600 277.050 667.050 ;
        RECT 295.950 666.600 298.050 667.050 ;
        RECT 274.950 665.400 298.050 666.600 ;
        RECT 274.950 664.950 277.050 665.400 ;
        RECT 295.950 664.950 298.050 665.400 ;
        RECT 337.950 666.600 340.050 667.050 ;
        RECT 352.950 666.600 355.050 667.050 ;
        RECT 337.950 665.400 355.050 666.600 ;
        RECT 356.400 666.600 357.600 670.950 ;
        RECT 367.950 669.600 370.050 670.050 ;
        RECT 392.400 669.600 393.600 670.950 ;
        RECT 367.950 668.400 393.600 669.600 ;
        RECT 406.950 669.600 409.050 670.050 ;
        RECT 445.950 669.600 448.050 670.050 ;
        RECT 452.400 669.600 453.600 671.400 ;
        RECT 406.950 668.400 453.600 669.600 ;
        RECT 367.950 667.950 370.050 668.400 ;
        RECT 406.950 667.950 409.050 668.400 ;
        RECT 445.950 667.950 448.050 668.400 ;
        RECT 454.950 667.950 457.050 670.050 ;
        RECT 460.950 669.600 463.050 670.050 ;
        RECT 466.950 669.600 469.050 670.050 ;
        RECT 460.950 668.400 469.050 669.600 ;
        RECT 470.400 669.600 471.600 671.400 ;
        RECT 490.950 671.400 508.050 672.600 ;
        RECT 490.950 670.950 493.050 671.400 ;
        RECT 502.950 670.950 505.050 671.400 ;
        RECT 505.950 670.950 508.050 671.400 ;
        RECT 517.950 670.950 520.050 673.050 ;
        RECT 535.950 672.600 538.050 673.050 ;
        RECT 556.950 672.600 559.050 673.050 ;
        RECT 535.950 671.400 559.050 672.600 ;
        RECT 535.950 670.950 538.050 671.400 ;
        RECT 556.950 670.950 559.050 671.400 ;
        RECT 616.950 672.600 619.050 673.050 ;
        RECT 640.950 672.600 643.050 673.050 ;
        RECT 616.950 671.400 643.050 672.600 ;
        RECT 616.950 670.950 619.050 671.400 ;
        RECT 640.950 670.950 643.050 671.400 ;
        RECT 646.950 672.600 649.050 673.050 ;
        RECT 676.950 672.600 679.050 673.050 ;
        RECT 646.950 671.400 679.050 672.600 ;
        RECT 646.950 670.950 649.050 671.400 ;
        RECT 676.950 670.950 679.050 671.400 ;
        RECT 487.950 669.600 490.050 670.050 ;
        RECT 493.950 669.600 496.050 670.050 ;
        RECT 470.400 668.400 496.050 669.600 ;
        RECT 460.950 667.950 463.050 668.400 ;
        RECT 466.950 667.950 469.050 668.400 ;
        RECT 487.950 667.950 490.050 668.400 ;
        RECT 493.950 667.950 496.050 668.400 ;
        RECT 508.950 669.600 511.050 670.050 ;
        RECT 553.950 669.600 556.050 670.050 ;
        RECT 508.950 668.400 556.050 669.600 ;
        RECT 508.950 667.950 511.050 668.400 ;
        RECT 553.950 667.950 556.050 668.400 ;
        RECT 559.950 669.600 562.050 670.050 ;
        RECT 568.950 669.600 571.050 670.050 ;
        RECT 559.950 668.400 571.050 669.600 ;
        RECT 559.950 667.950 562.050 668.400 ;
        RECT 568.950 667.950 571.050 668.400 ;
        RECT 634.950 669.600 637.050 670.050 ;
        RECT 643.950 669.600 646.050 670.050 ;
        RECT 634.950 668.400 646.050 669.600 ;
        RECT 634.950 667.950 637.050 668.400 ;
        RECT 643.950 667.950 646.050 668.400 ;
        RECT 700.950 669.600 703.050 670.050 ;
        RECT 706.950 669.600 709.050 670.050 ;
        RECT 700.950 668.400 709.050 669.600 ;
        RECT 700.950 667.950 703.050 668.400 ;
        RECT 706.950 667.950 709.050 668.400 ;
        RECT 373.950 666.600 376.050 667.050 ;
        RECT 356.400 665.400 376.050 666.600 ;
        RECT 337.950 664.950 340.050 665.400 ;
        RECT 352.950 664.950 355.050 665.400 ;
        RECT 373.950 664.950 376.050 665.400 ;
        RECT 379.950 666.600 382.050 667.050 ;
        RECT 400.950 666.600 403.050 667.050 ;
        RECT 379.950 665.400 403.050 666.600 ;
        RECT 455.400 666.600 456.600 667.950 ;
        RECT 460.950 666.600 463.050 667.050 ;
        RECT 455.400 665.400 463.050 666.600 ;
        RECT 379.950 664.950 382.050 665.400 ;
        RECT 400.950 664.950 403.050 665.400 ;
        RECT 460.950 664.950 463.050 665.400 ;
        RECT 547.950 666.600 550.050 667.050 ;
        RECT 565.950 666.600 568.050 667.050 ;
        RECT 613.950 666.600 616.050 667.050 ;
        RECT 547.950 665.400 616.050 666.600 ;
        RECT 547.950 664.950 550.050 665.400 ;
        RECT 565.950 664.950 568.050 665.400 ;
        RECT 613.950 664.950 616.050 665.400 ;
        RECT 625.950 666.600 628.050 667.050 ;
        RECT 643.950 666.600 646.050 667.050 ;
        RECT 625.950 665.400 646.050 666.600 ;
        RECT 625.950 664.950 628.050 665.400 ;
        RECT 643.950 664.950 646.050 665.400 ;
        RECT 691.950 666.600 694.050 667.050 ;
        RECT 709.950 666.600 712.050 667.050 ;
        RECT 691.950 665.400 712.050 666.600 ;
        RECT 691.950 664.950 694.050 665.400 ;
        RECT 709.950 664.950 712.050 665.400 ;
        RECT 136.950 663.600 139.050 664.050 ;
        RECT 163.950 663.600 166.050 664.050 ;
        RECT 136.950 662.400 166.050 663.600 ;
        RECT 136.950 661.950 139.050 662.400 ;
        RECT 163.950 661.950 166.050 662.400 ;
        RECT 175.950 663.600 178.050 664.050 ;
        RECT 202.950 663.600 205.050 664.050 ;
        RECT 238.950 663.600 241.050 664.050 ;
        RECT 364.950 663.600 367.050 664.050 ;
        RECT 175.950 662.400 192.600 663.600 ;
        RECT 175.950 661.950 178.050 662.400 ;
        RECT 157.950 660.600 160.050 661.050 ;
        RECT 187.950 660.600 190.050 661.050 ;
        RECT 134.400 659.400 156.600 660.600 ;
        RECT 49.950 658.950 52.050 659.400 ;
        RECT 103.950 658.950 106.050 659.400 ;
        RECT 97.950 657.600 100.050 658.050 ;
        RECT 109.950 657.600 112.050 658.050 ;
        RECT 97.950 656.400 112.050 657.600 ;
        RECT 155.400 657.600 156.600 659.400 ;
        RECT 157.950 659.400 190.050 660.600 ;
        RECT 191.400 660.600 192.600 662.400 ;
        RECT 202.950 662.400 367.050 663.600 ;
        RECT 202.950 661.950 205.050 662.400 ;
        RECT 238.950 661.950 241.050 662.400 ;
        RECT 364.950 661.950 367.050 662.400 ;
        RECT 385.950 663.600 388.050 664.050 ;
        RECT 394.950 663.600 397.050 664.050 ;
        RECT 385.950 662.400 397.050 663.600 ;
        RECT 385.950 661.950 388.050 662.400 ;
        RECT 394.950 661.950 397.050 662.400 ;
        RECT 451.950 663.600 454.050 664.050 ;
        RECT 478.950 663.600 481.050 664.050 ;
        RECT 451.950 662.400 481.050 663.600 ;
        RECT 451.950 661.950 454.050 662.400 ;
        RECT 478.950 661.950 481.050 662.400 ;
        RECT 211.950 660.600 214.050 661.050 ;
        RECT 191.400 659.400 214.050 660.600 ;
        RECT 157.950 658.950 160.050 659.400 ;
        RECT 187.950 658.950 190.050 659.400 ;
        RECT 211.950 658.950 214.050 659.400 ;
        RECT 232.950 660.600 235.050 661.050 ;
        RECT 262.950 660.600 265.050 661.050 ;
        RECT 304.950 660.600 307.050 661.050 ;
        RECT 232.950 659.400 307.050 660.600 ;
        RECT 232.950 658.950 235.050 659.400 ;
        RECT 262.950 658.950 265.050 659.400 ;
        RECT 304.950 658.950 307.050 659.400 ;
        RECT 628.950 660.600 631.050 661.050 ;
        RECT 658.950 660.600 661.050 661.050 ;
        RECT 628.950 659.400 661.050 660.600 ;
        RECT 628.950 658.950 631.050 659.400 ;
        RECT 658.950 658.950 661.050 659.400 ;
        RECT 181.950 657.600 184.050 658.050 ;
        RECT 155.400 656.400 184.050 657.600 ;
        RECT 97.950 655.950 100.050 656.400 ;
        RECT 109.950 655.950 112.050 656.400 ;
        RECT 181.950 655.950 184.050 656.400 ;
        RECT 19.950 654.600 22.050 655.050 ;
        RECT 82.950 654.600 85.050 655.050 ;
        RECT 88.950 654.600 91.050 655.050 ;
        RECT 121.950 654.600 124.050 655.050 ;
        RECT 136.950 654.600 139.050 655.050 ;
        RECT 19.950 653.400 139.050 654.600 ;
        RECT 19.950 652.950 22.050 653.400 ;
        RECT 82.950 652.950 85.050 653.400 ;
        RECT 88.950 652.950 91.050 653.400 ;
        RECT 121.950 652.950 124.050 653.400 ;
        RECT 136.950 652.950 139.050 653.400 ;
        RECT 142.950 654.600 145.050 655.050 ;
        RECT 160.950 654.600 163.050 655.050 ;
        RECT 172.950 654.600 175.050 655.050 ;
        RECT 142.950 653.400 175.050 654.600 ;
        RECT 142.950 652.950 145.050 653.400 ;
        RECT 160.950 652.950 163.050 653.400 ;
        RECT 172.950 652.950 175.050 653.400 ;
        RECT 67.950 648.600 70.050 649.050 ;
        RECT 85.950 648.600 88.050 649.050 ;
        RECT 67.950 647.400 88.050 648.600 ;
        RECT 67.950 646.950 70.050 647.400 ;
        RECT 85.950 646.950 88.050 647.400 ;
        RECT 268.950 648.600 271.050 649.050 ;
        RECT 283.950 648.600 286.050 649.050 ;
        RECT 289.950 648.600 292.050 649.050 ;
        RECT 313.950 648.600 316.050 649.050 ;
        RECT 268.950 647.400 316.050 648.600 ;
        RECT 268.950 646.950 271.050 647.400 ;
        RECT 283.950 646.950 286.050 647.400 ;
        RECT 289.950 646.950 292.050 647.400 ;
        RECT 313.950 646.950 316.050 647.400 ;
        RECT 604.950 645.600 607.050 646.050 ;
        RECT 613.950 645.600 616.050 646.050 ;
        RECT 619.950 645.600 622.050 646.050 ;
        RECT 604.950 644.400 622.050 645.600 ;
        RECT 604.950 643.950 607.050 644.400 ;
        RECT 613.950 643.950 616.050 644.400 ;
        RECT 619.950 643.950 622.050 644.400 ;
        RECT 700.950 645.600 703.050 646.050 ;
        RECT 709.950 645.600 712.050 646.050 ;
        RECT 700.950 644.400 712.050 645.600 ;
        RECT 700.950 643.950 703.050 644.400 ;
        RECT 709.950 643.950 712.050 644.400 ;
        RECT 52.950 642.600 55.050 643.050 ;
        RECT 61.950 642.600 64.050 643.050 ;
        RECT 52.950 641.400 64.050 642.600 ;
        RECT 52.950 640.950 55.050 641.400 ;
        RECT 61.950 640.950 64.050 641.400 ;
        RECT 316.950 642.600 319.050 643.050 ;
        RECT 478.950 642.600 481.050 643.050 ;
        RECT 316.950 641.400 481.050 642.600 ;
        RECT 316.950 640.950 319.050 641.400 ;
        RECT 478.950 640.950 481.050 641.400 ;
        RECT 250.950 639.600 253.050 640.050 ;
        RECT 466.950 639.600 469.050 640.050 ;
        RECT 487.950 639.600 490.050 640.050 ;
        RECT 250.950 638.400 300.600 639.600 ;
        RECT 250.950 637.950 253.050 638.400 ;
        RECT 4.950 636.600 7.050 637.050 ;
        RECT 13.950 636.600 16.050 637.050 ;
        RECT 4.950 635.400 16.050 636.600 ;
        RECT 4.950 634.950 7.050 635.400 ;
        RECT 13.950 634.950 16.050 635.400 ;
        RECT 208.950 636.600 211.050 637.050 ;
        RECT 232.950 636.600 235.050 637.050 ;
        RECT 268.950 636.600 271.050 637.050 ;
        RECT 289.950 636.600 292.050 637.050 ;
        RECT 208.950 635.400 222.600 636.600 ;
        RECT 208.950 634.950 211.050 635.400 ;
        RECT 221.400 634.050 222.600 635.400 ;
        RECT 232.950 635.400 292.050 636.600 ;
        RECT 232.950 634.950 235.050 635.400 ;
        RECT 268.950 634.950 271.050 635.400 ;
        RECT 289.950 634.950 292.050 635.400 ;
        RECT 10.950 633.600 13.050 634.050 ;
        RECT 22.950 633.600 25.050 634.050 ;
        RECT 31.950 633.600 34.050 634.050 ;
        RECT 46.950 633.600 49.050 634.050 ;
        RECT 97.950 633.600 100.050 634.050 ;
        RECT 118.950 633.600 121.050 634.050 ;
        RECT 136.950 633.600 139.050 634.050 ;
        RECT 10.950 632.400 18.600 633.600 ;
        RECT 10.950 631.950 13.050 632.400 ;
        RECT 13.950 628.950 16.050 631.050 ;
        RECT 10.950 627.600 13.050 628.050 ;
        RECT 14.400 627.600 15.600 628.950 ;
        RECT 10.950 626.400 15.600 627.600 ;
        RECT 10.950 625.950 13.050 626.400 ;
        RECT 17.400 625.050 18.600 632.400 ;
        RECT 22.950 632.400 27.600 633.600 ;
        RECT 22.950 631.950 25.050 632.400 ;
        RECT 19.950 630.600 22.050 631.050 ;
        RECT 26.400 630.600 27.600 632.400 ;
        RECT 31.950 632.400 39.600 633.600 ;
        RECT 31.950 631.950 34.050 632.400 ;
        RECT 34.950 630.600 37.050 631.050 ;
        RECT 19.950 629.400 24.600 630.600 ;
        RECT 26.400 629.400 37.050 630.600 ;
        RECT 38.400 630.600 39.600 632.400 ;
        RECT 46.950 632.400 75.600 633.600 ;
        RECT 46.950 631.950 49.050 632.400 ;
        RECT 61.950 630.600 64.050 631.050 ;
        RECT 70.950 630.600 73.050 631.050 ;
        RECT 38.400 629.400 42.600 630.600 ;
        RECT 19.950 628.950 22.050 629.400 ;
        RECT 23.400 627.600 24.600 629.400 ;
        RECT 34.950 628.950 37.050 629.400 ;
        RECT 37.950 627.600 40.050 628.050 ;
        RECT 23.400 626.400 40.050 627.600 ;
        RECT 41.400 627.600 42.600 629.400 ;
        RECT 47.400 629.400 73.050 630.600 ;
        RECT 74.400 630.600 75.600 632.400 ;
        RECT 97.950 632.400 108.600 633.600 ;
        RECT 97.950 631.950 100.050 632.400 ;
        RECT 76.950 630.600 79.050 631.050 ;
        RECT 74.400 629.400 79.050 630.600 ;
        RECT 43.950 627.600 46.050 628.050 ;
        RECT 41.400 626.400 46.050 627.600 ;
        RECT 37.950 625.950 40.050 626.400 ;
        RECT 43.950 625.950 46.050 626.400 ;
        RECT 47.400 625.050 48.600 629.400 ;
        RECT 61.950 628.950 64.050 629.400 ;
        RECT 70.950 628.950 73.050 629.400 ;
        RECT 76.950 628.950 79.050 629.400 ;
        RECT 103.950 628.950 106.050 631.050 ;
        RECT 107.400 630.600 108.600 632.400 ;
        RECT 118.950 632.400 139.050 633.600 ;
        RECT 118.950 631.950 121.050 632.400 ;
        RECT 136.950 631.950 139.050 632.400 ;
        RECT 157.950 633.600 160.050 634.050 ;
        RECT 166.950 633.600 169.050 634.050 ;
        RECT 157.950 632.400 169.050 633.600 ;
        RECT 157.950 631.950 160.050 632.400 ;
        RECT 166.950 631.950 169.050 632.400 ;
        RECT 193.950 633.600 196.050 634.050 ;
        RECT 214.950 633.600 217.050 634.050 ;
        RECT 193.950 632.400 219.600 633.600 ;
        RECT 193.950 631.950 196.050 632.400 ;
        RECT 214.950 631.950 217.050 632.400 ;
        RECT 218.400 631.050 219.600 632.400 ;
        RECT 220.950 631.950 223.050 634.050 ;
        RECT 274.950 631.950 277.050 634.050 ;
        RECT 280.950 631.950 283.050 634.050 ;
        RECT 286.950 633.600 289.050 634.050 ;
        RECT 295.950 633.600 298.050 634.050 ;
        RECT 286.950 632.400 298.050 633.600 ;
        RECT 286.950 631.950 289.050 632.400 ;
        RECT 295.950 631.950 298.050 632.400 ;
        RECT 115.950 630.600 118.050 631.050 ;
        RECT 107.400 629.400 118.050 630.600 ;
        RECT 115.950 628.950 118.050 629.400 ;
        RECT 142.950 628.950 145.050 631.050 ;
        RECT 184.950 630.600 187.050 631.050 ;
        RECT 196.950 630.600 199.050 631.050 ;
        RECT 184.950 629.400 199.050 630.600 ;
        RECT 184.950 628.950 187.050 629.400 ;
        RECT 196.950 628.950 199.050 629.400 ;
        RECT 217.950 630.600 220.050 631.050 ;
        RECT 232.950 630.600 235.050 631.050 ;
        RECT 217.950 629.400 235.050 630.600 ;
        RECT 217.950 628.950 220.050 629.400 ;
        RECT 232.950 628.950 235.050 629.400 ;
        RECT 259.950 630.600 262.050 631.050 ;
        RECT 271.950 630.600 274.050 631.050 ;
        RECT 259.950 629.400 274.050 630.600 ;
        RECT 259.950 628.950 262.050 629.400 ;
        RECT 271.950 628.950 274.050 629.400 ;
        RECT 52.950 627.600 55.050 628.050 ;
        RECT 58.950 627.600 61.050 628.050 ;
        RECT 52.950 626.400 61.050 627.600 ;
        RECT 52.950 625.950 55.050 626.400 ;
        RECT 58.950 625.950 61.050 626.400 ;
        RECT 73.950 627.600 76.050 628.050 ;
        RECT 104.400 627.600 105.600 628.950 ;
        RECT 121.950 627.600 124.050 628.050 ;
        RECT 73.950 626.400 124.050 627.600 ;
        RECT 73.950 625.950 76.050 626.400 ;
        RECT 121.950 625.950 124.050 626.400 ;
        RECT 127.950 627.600 130.050 628.050 ;
        RECT 133.950 627.600 136.050 628.050 ;
        RECT 127.950 626.400 136.050 627.600 ;
        RECT 143.400 627.600 144.600 628.950 ;
        RECT 163.950 627.600 166.050 628.050 ;
        RECT 143.400 626.400 166.050 627.600 ;
        RECT 127.950 625.950 130.050 626.400 ;
        RECT 133.950 625.950 136.050 626.400 ;
        RECT 163.950 625.950 166.050 626.400 ;
        RECT 184.950 627.600 187.050 628.050 ;
        RECT 190.950 627.600 193.050 628.050 ;
        RECT 184.950 626.400 193.050 627.600 ;
        RECT 184.950 625.950 187.050 626.400 ;
        RECT 190.950 625.950 193.050 626.400 ;
        RECT 199.950 627.600 202.050 628.050 ;
        RECT 208.950 627.600 211.050 628.050 ;
        RECT 199.950 626.400 211.050 627.600 ;
        RECT 199.950 625.950 202.050 626.400 ;
        RECT 208.950 625.950 211.050 626.400 ;
        RECT 262.950 627.600 265.050 628.050 ;
        RECT 275.400 627.600 276.600 631.950 ;
        RECT 262.950 626.400 276.600 627.600 ;
        RECT 262.950 625.950 265.050 626.400 ;
        RECT 16.950 622.950 19.050 625.050 ;
        RECT 46.950 622.950 49.050 625.050 ;
        RECT 82.950 624.600 85.050 625.050 ;
        RECT 100.950 624.600 103.050 625.050 ;
        RECT 82.950 623.400 103.050 624.600 ;
        RECT 82.950 622.950 85.050 623.400 ;
        RECT 100.950 622.950 103.050 623.400 ;
        RECT 103.950 624.600 106.050 625.050 ;
        RECT 106.950 624.600 109.050 625.050 ;
        RECT 112.950 624.600 115.050 625.050 ;
        RECT 103.950 623.400 115.050 624.600 ;
        RECT 103.950 622.950 106.050 623.400 ;
        RECT 106.950 622.950 109.050 623.400 ;
        RECT 112.950 622.950 115.050 623.400 ;
        RECT 130.950 624.600 133.050 625.050 ;
        RECT 139.950 624.600 142.050 625.050 ;
        RECT 130.950 623.400 142.050 624.600 ;
        RECT 130.950 622.950 133.050 623.400 ;
        RECT 139.950 622.950 142.050 623.400 ;
        RECT 223.950 624.600 226.050 625.050 ;
        RECT 250.950 624.600 253.050 625.050 ;
        RECT 281.400 624.600 282.600 631.950 ;
        RECT 283.950 628.950 286.050 631.050 ;
        RECT 299.400 630.600 300.600 638.400 ;
        RECT 466.950 638.400 490.050 639.600 ;
        RECT 466.950 637.950 469.050 638.400 ;
        RECT 487.950 637.950 490.050 638.400 ;
        RECT 400.950 636.600 403.050 637.050 ;
        RECT 490.950 636.600 493.050 637.050 ;
        RECT 400.950 635.400 493.050 636.600 ;
        RECT 400.950 634.950 403.050 635.400 ;
        RECT 490.950 634.950 493.050 635.400 ;
        RECT 508.950 636.600 511.050 637.050 ;
        RECT 523.950 636.600 526.050 637.050 ;
        RECT 508.950 635.400 526.050 636.600 ;
        RECT 508.950 634.950 511.050 635.400 ;
        RECT 523.950 634.950 526.050 635.400 ;
        RECT 547.950 636.600 550.050 637.050 ;
        RECT 556.950 636.600 559.050 637.050 ;
        RECT 628.950 636.600 631.050 637.050 ;
        RECT 547.950 635.400 631.050 636.600 ;
        RECT 547.950 634.950 550.050 635.400 ;
        RECT 556.950 634.950 559.050 635.400 ;
        RECT 628.950 634.950 631.050 635.400 ;
        RECT 631.950 636.600 634.050 637.050 ;
        RECT 682.950 636.600 685.050 637.050 ;
        RECT 631.950 635.400 685.050 636.600 ;
        RECT 631.950 634.950 634.050 635.400 ;
        RECT 682.950 634.950 685.050 635.400 ;
        RECT 301.950 633.600 304.050 634.050 ;
        RECT 436.950 633.600 439.050 634.050 ;
        RECT 463.950 633.600 466.050 634.050 ;
        RECT 301.950 632.400 315.600 633.600 ;
        RECT 301.950 631.950 304.050 632.400 ;
        RECT 314.400 631.050 315.600 632.400 ;
        RECT 436.950 632.400 466.050 633.600 ;
        RECT 436.950 631.950 439.050 632.400 ;
        RECT 463.950 631.950 466.050 632.400 ;
        RECT 484.950 631.950 487.050 634.050 ;
        RECT 496.950 633.600 499.050 634.050 ;
        RECT 541.950 633.600 544.050 634.050 ;
        RECT 550.950 633.600 553.050 634.050 ;
        RECT 496.950 632.400 553.050 633.600 ;
        RECT 496.950 631.950 499.050 632.400 ;
        RECT 541.950 631.950 544.050 632.400 ;
        RECT 550.950 631.950 553.050 632.400 ;
        RECT 589.950 633.600 592.050 634.050 ;
        RECT 619.950 633.600 622.050 634.050 ;
        RECT 589.950 632.400 622.050 633.600 ;
        RECT 589.950 631.950 592.050 632.400 ;
        RECT 619.950 631.950 622.050 632.400 ;
        RECT 290.400 629.400 300.600 630.600 ;
        RECT 284.400 627.600 285.600 628.950 ;
        RECT 290.400 628.050 291.600 629.400 ;
        RECT 313.950 628.950 316.050 631.050 ;
        RECT 373.950 630.600 376.050 631.050 ;
        RECT 430.950 630.600 433.050 631.050 ;
        RECT 451.950 630.600 454.050 631.050 ;
        RECT 373.950 629.400 429.600 630.600 ;
        RECT 373.950 628.950 376.050 629.400 ;
        RECT 284.400 626.400 288.600 627.600 ;
        RECT 283.950 624.600 286.050 625.050 ;
        RECT 223.950 623.400 286.050 624.600 ;
        RECT 287.400 624.600 288.600 626.400 ;
        RECT 289.950 625.950 292.050 628.050 ;
        RECT 352.950 627.600 355.050 628.050 ;
        RECT 382.950 627.600 385.050 628.050 ;
        RECT 352.950 626.400 385.050 627.600 ;
        RECT 352.950 625.950 355.050 626.400 ;
        RECT 382.950 625.950 385.050 626.400 ;
        RECT 388.950 627.600 391.050 628.050 ;
        RECT 394.950 627.600 397.050 628.050 ;
        RECT 388.950 626.400 397.050 627.600 ;
        RECT 428.400 627.600 429.600 629.400 ;
        RECT 430.950 629.400 454.050 630.600 ;
        RECT 430.950 628.950 433.050 629.400 ;
        RECT 451.950 628.950 454.050 629.400 ;
        RECT 457.950 630.600 460.050 631.050 ;
        RECT 466.950 630.600 469.050 631.050 ;
        RECT 457.950 629.400 469.050 630.600 ;
        RECT 485.400 630.600 486.600 631.950 ;
        RECT 493.950 630.600 496.050 631.050 ;
        RECT 485.400 629.400 496.050 630.600 ;
        RECT 457.950 628.950 460.050 629.400 ;
        RECT 466.950 628.950 469.050 629.400 ;
        RECT 493.950 628.950 496.050 629.400 ;
        RECT 571.950 630.600 574.050 631.050 ;
        RECT 574.950 630.600 577.050 631.050 ;
        RECT 571.950 629.400 591.600 630.600 ;
        RECT 571.950 628.950 574.050 629.400 ;
        RECT 574.950 628.950 577.050 629.400 ;
        RECT 439.950 627.600 442.050 628.050 ;
        RECT 428.400 626.400 442.050 627.600 ;
        RECT 388.950 625.950 391.050 626.400 ;
        RECT 394.950 625.950 397.050 626.400 ;
        RECT 439.950 625.950 442.050 626.400 ;
        RECT 445.950 627.600 448.050 628.050 ;
        RECT 452.400 627.600 453.600 628.950 ;
        RECT 445.950 626.400 453.600 627.600 ;
        RECT 481.950 627.600 484.050 628.050 ;
        RECT 523.950 627.600 526.050 628.050 ;
        RECT 481.950 626.400 526.050 627.600 ;
        RECT 445.950 625.950 448.050 626.400 ;
        RECT 481.950 625.950 484.050 626.400 ;
        RECT 523.950 625.950 526.050 626.400 ;
        RECT 541.950 627.600 544.050 628.050 ;
        RECT 565.950 627.600 568.050 628.050 ;
        RECT 541.950 626.400 568.050 627.600 ;
        RECT 541.950 625.950 544.050 626.400 ;
        RECT 565.950 625.950 568.050 626.400 ;
        RECT 580.950 627.600 583.050 628.050 ;
        RECT 586.950 627.600 589.050 628.050 ;
        RECT 580.950 626.400 589.050 627.600 ;
        RECT 590.400 627.600 591.600 629.400 ;
        RECT 625.950 628.950 628.050 631.050 ;
        RECT 646.950 630.600 649.050 631.050 ;
        RECT 664.950 630.600 667.050 631.050 ;
        RECT 646.950 629.400 667.050 630.600 ;
        RECT 646.950 628.950 649.050 629.400 ;
        RECT 664.950 628.950 667.050 629.400 ;
        RECT 670.950 630.600 673.050 631.050 ;
        RECT 706.950 630.600 709.050 631.050 ;
        RECT 670.950 629.400 709.050 630.600 ;
        RECT 670.950 628.950 673.050 629.400 ;
        RECT 706.950 628.950 709.050 629.400 ;
        RECT 607.950 627.600 610.050 628.050 ;
        RECT 590.400 626.400 610.050 627.600 ;
        RECT 580.950 625.950 583.050 626.400 ;
        RECT 586.950 625.950 589.050 626.400 ;
        RECT 607.950 625.950 610.050 626.400 ;
        RECT 295.950 624.600 298.050 625.050 ;
        RECT 287.400 623.400 298.050 624.600 ;
        RECT 223.950 622.950 226.050 623.400 ;
        RECT 250.950 622.950 253.050 623.400 ;
        RECT 283.950 622.950 286.050 623.400 ;
        RECT 295.950 622.950 298.050 623.400 ;
        RECT 376.950 624.600 379.050 625.050 ;
        RECT 382.950 624.600 385.050 625.050 ;
        RECT 376.950 623.400 385.050 624.600 ;
        RECT 376.950 622.950 379.050 623.400 ;
        RECT 382.950 622.950 385.050 623.400 ;
        RECT 388.950 624.600 391.050 625.050 ;
        RECT 427.950 624.600 430.050 625.050 ;
        RECT 388.950 623.400 430.050 624.600 ;
        RECT 388.950 622.950 391.050 623.400 ;
        RECT 427.950 622.950 430.050 623.400 ;
        RECT 442.950 624.600 445.050 625.050 ;
        RECT 460.950 624.600 463.050 625.050 ;
        RECT 463.950 624.600 466.050 625.050 ;
        RECT 442.950 623.400 466.050 624.600 ;
        RECT 442.950 622.950 445.050 623.400 ;
        RECT 460.950 622.950 463.050 623.400 ;
        RECT 463.950 622.950 466.050 623.400 ;
        RECT 487.950 624.600 490.050 625.050 ;
        RECT 499.950 624.600 502.050 625.050 ;
        RECT 487.950 623.400 502.050 624.600 ;
        RECT 487.950 622.950 490.050 623.400 ;
        RECT 499.950 622.950 502.050 623.400 ;
        RECT 505.950 624.600 508.050 625.050 ;
        RECT 514.950 624.600 517.050 625.050 ;
        RECT 505.950 623.400 517.050 624.600 ;
        RECT 505.950 622.950 508.050 623.400 ;
        RECT 514.950 622.950 517.050 623.400 ;
        RECT 547.950 624.600 550.050 625.050 ;
        RECT 559.950 624.600 562.050 625.050 ;
        RECT 547.950 623.400 562.050 624.600 ;
        RECT 547.950 622.950 550.050 623.400 ;
        RECT 559.950 622.950 562.050 623.400 ;
        RECT 610.950 624.600 613.050 625.050 ;
        RECT 626.400 624.600 627.600 628.950 ;
        RECT 655.950 627.600 658.050 628.050 ;
        RECT 676.950 627.600 679.050 628.050 ;
        RECT 655.950 626.400 679.050 627.600 ;
        RECT 655.950 625.950 658.050 626.400 ;
        RECT 676.950 625.950 679.050 626.400 ;
        RECT 610.950 623.400 627.600 624.600 ;
        RECT 628.950 624.600 631.050 625.050 ;
        RECT 649.950 624.600 652.050 625.050 ;
        RECT 667.950 624.600 670.050 625.050 ;
        RECT 628.950 623.400 670.050 624.600 ;
        RECT 610.950 622.950 613.050 623.400 ;
        RECT 628.950 622.950 631.050 623.400 ;
        RECT 649.950 622.950 652.050 623.400 ;
        RECT 667.950 622.950 670.050 623.400 ;
        RECT 7.950 621.600 10.050 622.050 ;
        RECT 43.950 621.600 46.050 622.050 ;
        RECT 7.950 620.400 46.050 621.600 ;
        RECT 7.950 619.950 10.050 620.400 ;
        RECT 43.950 619.950 46.050 620.400 ;
        RECT 88.950 621.600 91.050 622.050 ;
        RECT 115.950 621.600 118.050 622.050 ;
        RECT 88.950 620.400 118.050 621.600 ;
        RECT 88.950 619.950 91.050 620.400 ;
        RECT 115.950 619.950 118.050 620.400 ;
        RECT 133.950 621.600 136.050 622.050 ;
        RECT 154.950 621.600 157.050 622.050 ;
        RECT 169.950 621.600 172.050 622.050 ;
        RECT 133.950 620.400 172.050 621.600 ;
        RECT 133.950 619.950 136.050 620.400 ;
        RECT 154.950 619.950 157.050 620.400 ;
        RECT 169.950 619.950 172.050 620.400 ;
        RECT 178.950 621.600 181.050 622.050 ;
        RECT 217.950 621.600 220.050 622.050 ;
        RECT 178.950 620.400 220.050 621.600 ;
        RECT 178.950 619.950 181.050 620.400 ;
        RECT 217.950 619.950 220.050 620.400 ;
        RECT 277.950 621.600 280.050 622.050 ;
        RECT 310.950 621.600 313.050 622.050 ;
        RECT 277.950 620.400 313.050 621.600 ;
        RECT 277.950 619.950 280.050 620.400 ;
        RECT 310.950 619.950 313.050 620.400 ;
        RECT 436.950 621.600 439.050 622.050 ;
        RECT 442.950 621.600 445.050 622.050 ;
        RECT 448.950 621.600 451.050 622.050 ;
        RECT 436.950 620.400 451.050 621.600 ;
        RECT 436.950 619.950 439.050 620.400 ;
        RECT 442.950 619.950 445.050 620.400 ;
        RECT 448.950 619.950 451.050 620.400 ;
        RECT 586.950 621.600 589.050 622.050 ;
        RECT 673.950 621.600 676.050 622.050 ;
        RECT 676.950 621.600 679.050 622.050 ;
        RECT 688.950 621.600 691.050 622.050 ;
        RECT 586.950 620.400 691.050 621.600 ;
        RECT 586.950 619.950 589.050 620.400 ;
        RECT 673.950 619.950 676.050 620.400 ;
        RECT 676.950 619.950 679.050 620.400 ;
        RECT 688.950 619.950 691.050 620.400 ;
        RECT 25.950 618.600 28.050 619.050 ;
        RECT 55.950 618.600 58.050 619.050 ;
        RECT 25.950 617.400 58.050 618.600 ;
        RECT 25.950 616.950 28.050 617.400 ;
        RECT 55.950 616.950 58.050 617.400 ;
        RECT 76.950 618.600 79.050 619.050 ;
        RECT 88.950 618.600 91.050 619.050 ;
        RECT 76.950 617.400 91.050 618.600 ;
        RECT 76.950 616.950 79.050 617.400 ;
        RECT 88.950 616.950 91.050 617.400 ;
        RECT 160.950 618.600 163.050 619.050 ;
        RECT 199.950 618.600 202.050 619.050 ;
        RECT 160.950 617.400 202.050 618.600 ;
        RECT 160.950 616.950 163.050 617.400 ;
        RECT 199.950 616.950 202.050 617.400 ;
        RECT 211.950 618.600 214.050 619.050 ;
        RECT 256.950 618.600 259.050 619.050 ;
        RECT 319.950 618.600 322.050 619.050 ;
        RECT 325.950 618.600 328.050 619.050 ;
        RECT 211.950 617.400 328.050 618.600 ;
        RECT 211.950 616.950 214.050 617.400 ;
        RECT 256.950 616.950 259.050 617.400 ;
        RECT 319.950 616.950 322.050 617.400 ;
        RECT 325.950 616.950 328.050 617.400 ;
        RECT 412.950 618.600 415.050 619.050 ;
        RECT 454.950 618.600 457.050 619.050 ;
        RECT 412.950 617.400 457.050 618.600 ;
        RECT 412.950 616.950 415.050 617.400 ;
        RECT 454.950 616.950 457.050 617.400 ;
        RECT 472.950 618.600 475.050 619.050 ;
        RECT 655.950 618.600 658.050 619.050 ;
        RECT 472.950 617.400 658.050 618.600 ;
        RECT 472.950 616.950 475.050 617.400 ;
        RECT 655.950 616.950 658.050 617.400 ;
        RECT 661.950 618.600 664.050 619.050 ;
        RECT 694.950 618.600 697.050 619.050 ;
        RECT 661.950 617.400 697.050 618.600 ;
        RECT 661.950 616.950 664.050 617.400 ;
        RECT 694.950 616.950 697.050 617.400 ;
        RECT 22.950 615.600 25.050 616.050 ;
        RECT 64.950 615.600 67.050 616.050 ;
        RECT 22.950 614.400 67.050 615.600 ;
        RECT 22.950 613.950 25.050 614.400 ;
        RECT 64.950 613.950 67.050 614.400 ;
        RECT 202.950 615.600 205.050 616.050 ;
        RECT 211.950 615.600 214.050 616.050 ;
        RECT 202.950 614.400 214.050 615.600 ;
        RECT 202.950 613.950 205.050 614.400 ;
        RECT 211.950 613.950 214.050 614.400 ;
        RECT 241.950 615.600 244.050 616.050 ;
        RECT 247.950 615.600 250.050 616.050 ;
        RECT 256.950 615.600 259.050 616.050 ;
        RECT 241.950 614.400 259.050 615.600 ;
        RECT 241.950 613.950 244.050 614.400 ;
        RECT 247.950 613.950 250.050 614.400 ;
        RECT 256.950 613.950 259.050 614.400 ;
        RECT 298.950 615.600 301.050 616.050 ;
        RECT 310.950 615.600 313.050 616.050 ;
        RECT 346.950 615.600 349.050 616.050 ;
        RECT 298.950 614.400 349.050 615.600 ;
        RECT 298.950 613.950 301.050 614.400 ;
        RECT 310.950 613.950 313.050 614.400 ;
        RECT 346.950 613.950 349.050 614.400 ;
        RECT 532.950 615.600 535.050 616.050 ;
        RECT 553.950 615.600 556.050 616.050 ;
        RECT 532.950 614.400 556.050 615.600 ;
        RECT 532.950 613.950 535.050 614.400 ;
        RECT 553.950 613.950 556.050 614.400 ;
        RECT 604.950 615.600 607.050 616.050 ;
        RECT 631.950 615.600 634.050 616.050 ;
        RECT 604.950 614.400 634.050 615.600 ;
        RECT 604.950 613.950 607.050 614.400 ;
        RECT 631.950 613.950 634.050 614.400 ;
        RECT 634.950 615.600 637.050 616.050 ;
        RECT 643.950 615.600 646.050 616.050 ;
        RECT 634.950 614.400 646.050 615.600 ;
        RECT 634.950 613.950 637.050 614.400 ;
        RECT 643.950 613.950 646.050 614.400 ;
        RECT 22.950 612.600 25.050 613.050 ;
        RECT 40.950 612.600 43.050 613.050 ;
        RECT 49.950 612.600 52.050 613.050 ;
        RECT 22.950 611.400 52.050 612.600 ;
        RECT 22.950 610.950 25.050 611.400 ;
        RECT 40.950 610.950 43.050 611.400 ;
        RECT 49.950 610.950 52.050 611.400 ;
        RECT 229.950 612.600 232.050 613.050 ;
        RECT 280.950 612.600 283.050 613.050 ;
        RECT 229.950 611.400 283.050 612.600 ;
        RECT 229.950 610.950 232.050 611.400 ;
        RECT 280.950 610.950 283.050 611.400 ;
        RECT 340.950 612.600 343.050 613.050 ;
        RECT 406.950 612.600 409.050 613.050 ;
        RECT 421.950 612.600 424.050 613.050 ;
        RECT 529.950 612.600 532.050 613.050 ;
        RECT 547.950 612.600 550.050 613.050 ;
        RECT 580.950 612.600 583.050 613.050 ;
        RECT 340.950 611.400 583.050 612.600 ;
        RECT 340.950 610.950 343.050 611.400 ;
        RECT 406.950 610.950 409.050 611.400 ;
        RECT 421.950 610.950 424.050 611.400 ;
        RECT 529.950 610.950 532.050 611.400 ;
        RECT 547.950 610.950 550.050 611.400 ;
        RECT 580.950 610.950 583.050 611.400 ;
        RECT 28.950 609.600 31.050 610.050 ;
        RECT 43.950 609.600 46.050 610.050 ;
        RECT 28.950 608.400 46.050 609.600 ;
        RECT 28.950 607.950 31.050 608.400 ;
        RECT 43.950 607.950 46.050 608.400 ;
        RECT 97.950 609.600 100.050 610.050 ;
        RECT 118.950 609.600 121.050 610.050 ;
        RECT 160.950 609.600 163.050 610.050 ;
        RECT 97.950 608.400 163.050 609.600 ;
        RECT 97.950 607.950 100.050 608.400 ;
        RECT 118.950 607.950 121.050 608.400 ;
        RECT 160.950 607.950 163.050 608.400 ;
        RECT 271.950 609.600 274.050 610.050 ;
        RECT 337.950 609.600 340.050 610.050 ;
        RECT 271.950 608.400 340.050 609.600 ;
        RECT 271.950 607.950 274.050 608.400 ;
        RECT 337.950 607.950 340.050 608.400 ;
        RECT 502.950 609.600 505.050 610.050 ;
        RECT 604.950 609.600 607.050 610.050 ;
        RECT 610.950 609.600 613.050 610.050 ;
        RECT 502.950 608.400 613.050 609.600 ;
        RECT 502.950 607.950 505.050 608.400 ;
        RECT 604.950 607.950 607.050 608.400 ;
        RECT 610.950 607.950 613.050 608.400 ;
        RECT 613.950 609.600 616.050 610.050 ;
        RECT 619.950 609.600 622.050 610.050 ;
        RECT 628.950 609.600 631.050 610.050 ;
        RECT 613.950 608.400 631.050 609.600 ;
        RECT 613.950 607.950 616.050 608.400 ;
        RECT 619.950 607.950 622.050 608.400 ;
        RECT 628.950 607.950 631.050 608.400 ;
        RECT 7.950 606.600 10.050 607.050 ;
        RECT 55.950 606.600 58.050 607.050 ;
        RECT 7.950 605.400 58.050 606.600 ;
        RECT 7.950 604.950 10.050 605.400 ;
        RECT 55.950 604.950 58.050 605.400 ;
        RECT 61.950 606.600 64.050 607.050 ;
        RECT 127.950 606.600 130.050 607.050 ;
        RECT 139.950 606.600 142.050 607.050 ;
        RECT 61.950 605.400 142.050 606.600 ;
        RECT 61.950 604.950 64.050 605.400 ;
        RECT 127.950 604.950 130.050 605.400 ;
        RECT 139.950 604.950 142.050 605.400 ;
        RECT 142.950 606.600 145.050 607.050 ;
        RECT 181.950 606.600 184.050 607.050 ;
        RECT 205.950 606.600 208.050 607.050 ;
        RECT 142.950 605.400 208.050 606.600 ;
        RECT 142.950 604.950 145.050 605.400 ;
        RECT 181.950 604.950 184.050 605.400 ;
        RECT 205.950 604.950 208.050 605.400 ;
        RECT 268.950 606.600 271.050 607.050 ;
        RECT 289.950 606.600 292.050 607.050 ;
        RECT 268.950 605.400 292.050 606.600 ;
        RECT 268.950 604.950 271.050 605.400 ;
        RECT 289.950 604.950 292.050 605.400 ;
        RECT 307.950 606.600 310.050 607.050 ;
        RECT 340.950 606.600 343.050 607.050 ;
        RECT 355.950 606.600 358.050 607.050 ;
        RECT 307.950 605.400 358.050 606.600 ;
        RECT 307.950 604.950 310.050 605.400 ;
        RECT 340.950 604.950 343.050 605.400 ;
        RECT 355.950 604.950 358.050 605.400 ;
        RECT 409.950 606.600 412.050 607.050 ;
        RECT 448.950 606.600 451.050 607.050 ;
        RECT 409.950 605.400 451.050 606.600 ;
        RECT 409.950 604.950 412.050 605.400 ;
        RECT 448.950 604.950 451.050 605.400 ;
        RECT 484.950 606.600 487.050 607.050 ;
        RECT 550.950 606.600 553.050 607.050 ;
        RECT 484.950 605.400 553.050 606.600 ;
        RECT 484.950 604.950 487.050 605.400 ;
        RECT 550.950 604.950 553.050 605.400 ;
        RECT 577.950 606.600 580.050 607.050 ;
        RECT 589.950 606.600 592.050 607.050 ;
        RECT 613.950 606.600 616.050 607.050 ;
        RECT 577.950 605.400 616.050 606.600 ;
        RECT 577.950 604.950 580.050 605.400 ;
        RECT 589.950 604.950 592.050 605.400 ;
        RECT 613.950 604.950 616.050 605.400 ;
        RECT 10.950 603.600 13.050 604.050 ;
        RECT 31.950 603.600 34.050 604.050 ;
        RECT 10.950 602.400 34.050 603.600 ;
        RECT 10.950 601.950 13.050 602.400 ;
        RECT 31.950 601.950 34.050 602.400 ;
        RECT 49.950 603.600 52.050 604.050 ;
        RECT 73.950 603.600 76.050 604.050 ;
        RECT 106.950 603.600 109.050 604.050 ;
        RECT 184.950 603.600 187.050 604.050 ;
        RECT 202.950 603.600 205.050 604.050 ;
        RECT 214.950 603.600 217.050 604.050 ;
        RECT 49.950 602.400 96.600 603.600 ;
        RECT 49.950 601.950 52.050 602.400 ;
        RECT 73.950 601.950 76.050 602.400 ;
        RECT 64.950 600.600 67.050 601.050 ;
        RECT 76.950 600.600 79.050 601.050 ;
        RECT 91.950 600.600 94.050 601.050 ;
        RECT 64.950 599.400 79.050 600.600 ;
        RECT 64.950 598.950 67.050 599.400 ;
        RECT 76.950 598.950 79.050 599.400 ;
        RECT 80.400 599.400 94.050 600.600 ;
        RECT 37.950 597.600 40.050 598.050 ;
        RECT 40.950 597.600 43.050 598.050 ;
        RECT 80.400 597.600 81.600 599.400 ;
        RECT 91.950 598.950 94.050 599.400 ;
        RECT 95.400 598.050 96.600 602.400 ;
        RECT 106.950 602.400 217.050 603.600 ;
        RECT 106.950 601.950 109.050 602.400 ;
        RECT 184.950 601.950 187.050 602.400 ;
        RECT 202.950 601.950 205.050 602.400 ;
        RECT 214.950 601.950 217.050 602.400 ;
        RECT 220.950 603.600 223.050 604.050 ;
        RECT 247.950 603.600 250.050 604.050 ;
        RECT 271.950 603.600 274.050 604.050 ;
        RECT 220.950 602.400 231.600 603.600 ;
        RECT 220.950 601.950 223.050 602.400 ;
        RECT 115.950 600.600 118.050 601.050 ;
        RECT 110.400 599.400 118.050 600.600 ;
        RECT 37.950 596.400 81.600 597.600 ;
        RECT 82.950 597.600 85.050 598.050 ;
        RECT 82.950 596.400 93.600 597.600 ;
        RECT 37.950 595.950 40.050 596.400 ;
        RECT 40.950 595.950 43.050 596.400 ;
        RECT 82.950 595.950 85.050 596.400 ;
        RECT 4.950 594.600 7.050 595.050 ;
        RECT 28.950 594.600 31.050 595.050 ;
        RECT 4.950 593.400 31.050 594.600 ;
        RECT 41.400 594.600 42.600 595.950 ;
        RECT 52.950 594.600 55.050 595.050 ;
        RECT 41.400 593.400 55.050 594.600 ;
        RECT 92.400 594.600 93.600 596.400 ;
        RECT 94.950 595.950 97.050 598.050 ;
        RECT 100.950 595.950 103.050 598.050 ;
        RECT 101.400 594.600 102.600 595.950 ;
        RECT 92.400 593.400 102.600 594.600 ;
        RECT 4.950 592.950 7.050 593.400 ;
        RECT 28.950 592.950 31.050 593.400 ;
        RECT 52.950 592.950 55.050 593.400 ;
        RECT 19.950 591.600 22.050 592.050 ;
        RECT 67.950 591.600 70.050 592.050 ;
        RECT 85.950 591.600 88.050 592.050 ;
        RECT 19.950 590.400 88.050 591.600 ;
        RECT 19.950 589.950 22.050 590.400 ;
        RECT 67.950 589.950 70.050 590.400 ;
        RECT 85.950 589.950 88.050 590.400 ;
        RECT 97.950 591.600 100.050 592.050 ;
        RECT 110.400 591.600 111.600 599.400 ;
        RECT 115.950 598.950 118.050 599.400 ;
        RECT 148.950 600.600 151.050 601.050 ;
        RECT 151.950 600.600 154.050 601.050 ;
        RECT 148.950 599.400 154.050 600.600 ;
        RECT 148.950 598.950 151.050 599.400 ;
        RECT 151.950 598.950 154.050 599.400 ;
        RECT 208.950 600.600 211.050 601.050 ;
        RECT 226.950 600.600 229.050 601.050 ;
        RECT 208.950 599.400 229.050 600.600 ;
        RECT 208.950 598.950 211.050 599.400 ;
        RECT 226.950 598.950 229.050 599.400 ;
        RECT 112.950 597.600 115.050 598.050 ;
        RECT 121.950 597.600 124.050 598.050 ;
        RECT 145.950 597.600 148.050 598.050 ;
        RECT 112.950 596.400 124.050 597.600 ;
        RECT 112.950 595.950 115.050 596.400 ;
        RECT 121.950 595.950 124.050 596.400 ;
        RECT 143.400 596.400 148.050 597.600 ;
        RECT 113.400 592.050 114.600 595.950 ;
        RECT 115.950 594.600 118.050 595.050 ;
        RECT 124.950 594.600 127.050 595.050 ;
        RECT 115.950 593.400 127.050 594.600 ;
        RECT 115.950 592.950 118.050 593.400 ;
        RECT 124.950 592.950 127.050 593.400 ;
        RECT 97.950 590.400 111.600 591.600 ;
        RECT 97.950 589.950 100.050 590.400 ;
        RECT 112.950 589.950 115.050 592.050 ;
        RECT 125.400 591.600 126.600 592.950 ;
        RECT 130.950 591.600 133.050 592.050 ;
        RECT 125.400 590.400 133.050 591.600 ;
        RECT 143.400 591.600 144.600 596.400 ;
        RECT 145.950 595.950 148.050 596.400 ;
        RECT 145.950 594.600 148.050 595.050 ;
        RECT 149.400 594.600 150.600 598.950 ;
        RECT 154.950 597.600 157.050 598.050 ;
        RECT 169.950 597.600 172.050 598.050 ;
        RECT 154.950 596.400 172.050 597.600 ;
        RECT 154.950 595.950 157.050 596.400 ;
        RECT 169.950 595.950 172.050 596.400 ;
        RECT 193.950 597.600 196.050 598.050 ;
        RECT 199.950 597.600 202.050 598.050 ;
        RECT 193.950 596.400 202.050 597.600 ;
        RECT 193.950 595.950 196.050 596.400 ;
        RECT 199.950 595.950 202.050 596.400 ;
        RECT 145.950 593.400 150.600 594.600 ;
        RECT 163.950 594.600 166.050 595.050 ;
        RECT 178.950 594.600 181.050 595.050 ;
        RECT 163.950 593.400 181.050 594.600 ;
        RECT 145.950 592.950 148.050 593.400 ;
        RECT 163.950 592.950 166.050 593.400 ;
        RECT 178.950 592.950 181.050 593.400 ;
        RECT 208.950 594.600 211.050 595.050 ;
        RECT 217.950 594.600 220.050 595.050 ;
        RECT 208.950 593.400 220.050 594.600 ;
        RECT 208.950 592.950 211.050 593.400 ;
        RECT 217.950 592.950 220.050 593.400 ;
        RECT 223.950 594.600 226.050 595.050 ;
        RECT 230.400 594.600 231.600 602.400 ;
        RECT 247.950 602.400 274.050 603.600 ;
        RECT 247.950 601.950 250.050 602.400 ;
        RECT 271.950 601.950 274.050 602.400 ;
        RECT 286.950 603.600 289.050 604.050 ;
        RECT 292.950 603.600 295.050 604.050 ;
        RECT 286.950 602.400 295.050 603.600 ;
        RECT 286.950 601.950 289.050 602.400 ;
        RECT 292.950 601.950 295.050 602.400 ;
        RECT 358.950 603.600 361.050 604.050 ;
        RECT 364.950 603.600 367.050 604.050 ;
        RECT 358.950 602.400 367.050 603.600 ;
        RECT 358.950 601.950 361.050 602.400 ;
        RECT 364.950 601.950 367.050 602.400 ;
        RECT 385.950 603.600 388.050 604.050 ;
        RECT 457.950 603.600 460.050 604.050 ;
        RECT 385.950 602.400 460.050 603.600 ;
        RECT 385.950 601.950 388.050 602.400 ;
        RECT 457.950 601.950 460.050 602.400 ;
        RECT 460.950 603.600 463.050 604.050 ;
        RECT 481.950 603.600 484.050 604.050 ;
        RECT 490.950 603.600 493.050 604.050 ;
        RECT 496.950 603.600 499.050 604.050 ;
        RECT 460.950 602.400 499.050 603.600 ;
        RECT 460.950 601.950 463.050 602.400 ;
        RECT 481.950 601.950 484.050 602.400 ;
        RECT 490.950 601.950 493.050 602.400 ;
        RECT 496.950 601.950 499.050 602.400 ;
        RECT 499.950 603.600 502.050 604.050 ;
        RECT 517.950 603.600 520.050 604.050 ;
        RECT 499.950 602.400 520.050 603.600 ;
        RECT 499.950 601.950 502.050 602.400 ;
        RECT 517.950 601.950 520.050 602.400 ;
        RECT 520.950 603.600 523.050 604.050 ;
        RECT 562.950 603.600 565.050 604.050 ;
        RECT 586.950 603.600 589.050 604.050 ;
        RECT 520.950 602.400 565.050 603.600 ;
        RECT 520.950 601.950 523.050 602.400 ;
        RECT 562.950 601.950 565.050 602.400 ;
        RECT 575.400 602.400 589.050 603.600 ;
        RECT 238.950 600.600 241.050 601.050 ;
        RECT 244.950 600.600 247.050 601.050 ;
        RECT 238.950 599.400 247.050 600.600 ;
        RECT 238.950 598.950 241.050 599.400 ;
        RECT 244.950 598.950 247.050 599.400 ;
        RECT 250.950 600.600 253.050 601.050 ;
        RECT 253.950 600.600 256.050 601.050 ;
        RECT 262.950 600.600 265.050 601.050 ;
        RECT 250.950 599.400 265.050 600.600 ;
        RECT 250.950 598.950 253.050 599.400 ;
        RECT 253.950 598.950 256.050 599.400 ;
        RECT 262.950 598.950 265.050 599.400 ;
        RECT 265.950 598.950 268.050 601.050 ;
        RECT 274.950 598.950 277.050 601.050 ;
        RECT 340.950 600.600 343.050 601.050 ;
        RECT 352.950 600.600 355.050 601.050 ;
        RECT 340.950 599.400 355.050 600.600 ;
        RECT 340.950 598.950 343.050 599.400 ;
        RECT 352.950 598.950 355.050 599.400 ;
        RECT 415.950 598.950 418.050 601.050 ;
        RECT 463.950 600.600 466.050 601.050 ;
        RECT 463.950 599.400 486.600 600.600 ;
        RECT 463.950 598.950 466.050 599.400 ;
        RECT 223.950 593.400 231.600 594.600 ;
        RECT 223.950 592.950 226.050 593.400 ;
        RECT 154.950 591.600 157.050 592.050 ;
        RECT 143.400 590.400 157.050 591.600 ;
        RECT 130.950 589.950 133.050 590.400 ;
        RECT 154.950 589.950 157.050 590.400 ;
        RECT 211.950 591.600 214.050 592.050 ;
        RECT 220.950 591.600 223.050 592.050 ;
        RECT 229.950 591.600 232.050 592.050 ;
        RECT 211.950 590.400 232.050 591.600 ;
        RECT 266.400 591.600 267.600 598.950 ;
        RECT 275.400 595.050 276.600 598.950 ;
        RECT 286.950 597.600 289.050 598.050 ;
        RECT 295.950 597.600 298.050 598.050 ;
        RECT 286.950 596.400 298.050 597.600 ;
        RECT 286.950 595.950 289.050 596.400 ;
        RECT 295.950 595.950 298.050 596.400 ;
        RECT 313.950 597.600 316.050 598.050 ;
        RECT 322.950 597.600 325.050 598.050 ;
        RECT 313.950 596.400 325.050 597.600 ;
        RECT 313.950 595.950 316.050 596.400 ;
        RECT 322.950 595.950 325.050 596.400 ;
        RECT 331.950 597.600 334.050 598.050 ;
        RECT 343.950 597.600 346.050 598.050 ;
        RECT 331.950 596.400 346.050 597.600 ;
        RECT 331.950 595.950 334.050 596.400 ;
        RECT 343.950 595.950 346.050 596.400 ;
        RECT 391.950 597.600 394.050 598.050 ;
        RECT 416.400 597.600 417.600 598.950 ;
        RECT 391.950 596.400 417.600 597.600 ;
        RECT 436.950 597.600 439.050 598.050 ;
        RECT 445.950 597.600 448.050 598.050 ;
        RECT 436.950 596.400 448.050 597.600 ;
        RECT 391.950 595.950 394.050 596.400 ;
        RECT 436.950 595.950 439.050 596.400 ;
        RECT 445.950 595.950 448.050 596.400 ;
        RECT 451.950 597.600 454.050 598.050 ;
        RECT 472.950 597.600 475.050 598.050 ;
        RECT 451.950 596.400 475.050 597.600 ;
        RECT 485.400 597.600 486.600 599.400 ;
        RECT 502.950 598.950 505.050 601.050 ;
        RECT 505.950 600.600 508.050 601.050 ;
        RECT 511.950 600.600 514.050 601.050 ;
        RECT 505.950 599.400 514.050 600.600 ;
        RECT 505.950 598.950 508.050 599.400 ;
        RECT 511.950 598.950 514.050 599.400 ;
        RECT 514.950 598.950 517.050 601.050 ;
        RECT 553.950 600.600 556.050 601.050 ;
        RECT 571.950 600.600 574.050 601.050 ;
        RECT 553.950 599.400 574.050 600.600 ;
        RECT 553.950 598.950 556.050 599.400 ;
        RECT 571.950 598.950 574.050 599.400 ;
        RECT 487.950 597.600 490.050 598.050 ;
        RECT 485.400 596.400 490.050 597.600 ;
        RECT 451.950 595.950 454.050 596.400 ;
        RECT 472.950 595.950 475.050 596.400 ;
        RECT 487.950 595.950 490.050 596.400 ;
        RECT 503.400 595.050 504.600 598.950 ;
        RECT 515.400 597.600 516.600 598.950 ;
        RECT 575.400 598.050 576.600 602.400 ;
        RECT 586.950 601.950 589.050 602.400 ;
        RECT 601.950 603.600 604.050 604.050 ;
        RECT 622.950 603.600 625.050 604.050 ;
        RECT 601.950 602.400 625.050 603.600 ;
        RECT 601.950 601.950 604.050 602.400 ;
        RECT 622.950 601.950 625.050 602.400 ;
        RECT 583.950 600.600 586.050 601.050 ;
        RECT 578.400 599.400 586.050 600.600 ;
        RECT 578.400 598.050 579.600 599.400 ;
        RECT 583.950 598.950 586.050 599.400 ;
        RECT 598.950 600.600 601.050 601.050 ;
        RECT 607.950 600.600 610.050 601.050 ;
        RECT 598.950 599.400 610.050 600.600 ;
        RECT 598.950 598.950 601.050 599.400 ;
        RECT 607.950 598.950 610.050 599.400 ;
        RECT 616.950 600.600 619.050 601.050 ;
        RECT 628.950 600.600 631.050 601.050 ;
        RECT 640.950 600.600 643.050 601.050 ;
        RECT 616.950 599.400 627.600 600.600 ;
        RECT 616.950 598.950 619.050 599.400 ;
        RECT 626.400 598.050 627.600 599.400 ;
        RECT 628.950 599.400 643.050 600.600 ;
        RECT 628.950 598.950 631.050 599.400 ;
        RECT 640.950 598.950 643.050 599.400 ;
        RECT 643.950 600.600 646.050 601.050 ;
        RECT 682.950 600.600 685.050 601.050 ;
        RECT 643.950 599.400 685.050 600.600 ;
        RECT 643.950 598.950 646.050 599.400 ;
        RECT 682.950 598.950 685.050 599.400 ;
        RECT 526.950 597.600 529.050 598.050 ;
        RECT 506.400 596.400 529.050 597.600 ;
        RECT 506.400 595.050 507.600 596.400 ;
        RECT 526.950 595.950 529.050 596.400 ;
        RECT 574.950 595.950 577.050 598.050 ;
        RECT 577.950 595.950 580.050 598.050 ;
        RECT 625.950 595.950 628.050 598.050 ;
        RECT 631.950 597.600 634.050 598.050 ;
        RECT 646.950 597.600 649.050 598.050 ;
        RECT 631.950 596.400 649.050 597.600 ;
        RECT 631.950 595.950 634.050 596.400 ;
        RECT 646.950 595.950 649.050 596.400 ;
        RECT 661.950 597.600 664.050 598.050 ;
        RECT 700.950 597.600 703.050 598.050 ;
        RECT 706.950 597.600 709.050 598.050 ;
        RECT 661.950 596.400 709.050 597.600 ;
        RECT 661.950 595.950 664.050 596.400 ;
        RECT 700.950 595.950 703.050 596.400 ;
        RECT 706.950 595.950 709.050 596.400 ;
        RECT 274.950 592.950 277.050 595.050 ;
        RECT 277.950 594.600 280.050 595.050 ;
        RECT 298.950 594.600 301.050 595.050 ;
        RECT 277.950 593.400 301.050 594.600 ;
        RECT 277.950 592.950 280.050 593.400 ;
        RECT 298.950 592.950 301.050 593.400 ;
        RECT 400.950 594.600 403.050 595.050 ;
        RECT 415.950 594.600 418.050 595.050 ;
        RECT 400.950 593.400 418.050 594.600 ;
        RECT 400.950 592.950 403.050 593.400 ;
        RECT 415.950 592.950 418.050 593.400 ;
        RECT 439.950 594.600 442.050 595.050 ;
        RECT 469.950 594.600 472.050 595.050 ;
        RECT 439.950 593.400 472.050 594.600 ;
        RECT 439.950 592.950 442.050 593.400 ;
        RECT 469.950 592.950 472.050 593.400 ;
        RECT 502.950 592.950 505.050 595.050 ;
        RECT 505.950 592.950 508.050 595.050 ;
        RECT 550.950 594.600 553.050 595.050 ;
        RECT 595.950 594.600 598.050 595.050 ;
        RECT 550.950 593.400 598.050 594.600 ;
        RECT 550.950 592.950 553.050 593.400 ;
        RECT 595.950 592.950 598.050 593.400 ;
        RECT 271.950 591.600 274.050 592.050 ;
        RECT 266.400 590.400 274.050 591.600 ;
        RECT 211.950 589.950 214.050 590.400 ;
        RECT 220.950 589.950 223.050 590.400 ;
        RECT 229.950 589.950 232.050 590.400 ;
        RECT 271.950 589.950 274.050 590.400 ;
        RECT 475.950 591.600 478.050 592.050 ;
        RECT 535.950 591.600 538.050 592.050 ;
        RECT 577.950 591.600 580.050 592.050 ;
        RECT 475.950 590.400 580.050 591.600 ;
        RECT 475.950 589.950 478.050 590.400 ;
        RECT 535.950 589.950 538.050 590.400 ;
        RECT 577.950 589.950 580.050 590.400 ;
        RECT 37.950 588.600 40.050 589.050 ;
        RECT 64.950 588.600 67.050 589.050 ;
        RECT 79.950 588.600 82.050 589.050 ;
        RECT 37.950 587.400 82.050 588.600 ;
        RECT 37.950 586.950 40.050 587.400 ;
        RECT 64.950 586.950 67.050 587.400 ;
        RECT 79.950 586.950 82.050 587.400 ;
        RECT 103.950 588.600 106.050 589.050 ;
        RECT 127.950 588.600 130.050 589.050 ;
        RECT 103.950 587.400 130.050 588.600 ;
        RECT 103.950 586.950 106.050 587.400 ;
        RECT 127.950 586.950 130.050 587.400 ;
        RECT 571.950 588.600 574.050 589.050 ;
        RECT 580.950 588.600 583.050 589.050 ;
        RECT 694.950 588.600 697.050 589.050 ;
        RECT 571.950 587.400 697.050 588.600 ;
        RECT 571.950 586.950 574.050 587.400 ;
        RECT 580.950 586.950 583.050 587.400 ;
        RECT 694.950 586.950 697.050 587.400 ;
        RECT 7.950 585.600 10.050 586.050 ;
        RECT 46.950 585.600 49.050 586.050 ;
        RECT 58.950 585.600 61.050 586.050 ;
        RECT 7.950 584.400 61.050 585.600 ;
        RECT 7.950 583.950 10.050 584.400 ;
        RECT 46.950 583.950 49.050 584.400 ;
        RECT 58.950 583.950 61.050 584.400 ;
        RECT 79.950 585.600 82.050 586.050 ;
        RECT 88.950 585.600 91.050 586.050 ;
        RECT 79.950 584.400 91.050 585.600 ;
        RECT 79.950 583.950 82.050 584.400 ;
        RECT 88.950 583.950 91.050 584.400 ;
        RECT 166.950 585.600 169.050 586.050 ;
        RECT 184.950 585.600 187.050 586.050 ;
        RECT 190.950 585.600 193.050 586.050 ;
        RECT 166.950 584.400 193.050 585.600 ;
        RECT 166.950 583.950 169.050 584.400 ;
        RECT 184.950 583.950 187.050 584.400 ;
        RECT 190.950 583.950 193.050 584.400 ;
        RECT 22.950 582.600 25.050 583.050 ;
        RECT 25.950 582.600 28.050 583.050 ;
        RECT 55.950 582.600 58.050 583.050 ;
        RECT 22.950 581.400 58.050 582.600 ;
        RECT 22.950 580.950 25.050 581.400 ;
        RECT 25.950 580.950 28.050 581.400 ;
        RECT 55.950 580.950 58.050 581.400 ;
        RECT 199.950 579.600 202.050 580.050 ;
        RECT 226.950 579.600 229.050 580.050 ;
        RECT 235.950 579.600 238.050 580.050 ;
        RECT 199.950 578.400 238.050 579.600 ;
        RECT 199.950 577.950 202.050 578.400 ;
        RECT 226.950 577.950 229.050 578.400 ;
        RECT 235.950 577.950 238.050 578.400 ;
        RECT 634.950 579.600 637.050 580.050 ;
        RECT 643.950 579.600 646.050 580.050 ;
        RECT 634.950 578.400 646.050 579.600 ;
        RECT 634.950 577.950 637.050 578.400 ;
        RECT 643.950 577.950 646.050 578.400 ;
        RECT 550.950 576.600 553.050 577.050 ;
        RECT 607.950 576.600 610.050 577.050 ;
        RECT 646.950 576.600 649.050 577.050 ;
        RECT 550.950 575.400 649.050 576.600 ;
        RECT 550.950 574.950 553.050 575.400 ;
        RECT 607.950 574.950 610.050 575.400 ;
        RECT 646.950 574.950 649.050 575.400 ;
        RECT 130.950 570.600 133.050 571.050 ;
        RECT 154.950 570.600 157.050 571.050 ;
        RECT 175.950 570.600 178.050 571.050 ;
        RECT 130.950 569.400 178.050 570.600 ;
        RECT 130.950 568.950 133.050 569.400 ;
        RECT 154.950 568.950 157.050 569.400 ;
        RECT 175.950 568.950 178.050 569.400 ;
        RECT 124.950 567.600 127.050 568.050 ;
        RECT 142.950 567.600 145.050 568.050 ;
        RECT 124.950 566.400 145.050 567.600 ;
        RECT 124.950 565.950 127.050 566.400 ;
        RECT 142.950 565.950 145.050 566.400 ;
        RECT 61.950 564.600 64.050 565.050 ;
        RECT 88.950 564.600 91.050 565.050 ;
        RECT 61.950 563.400 91.050 564.600 ;
        RECT 61.950 562.950 64.050 563.400 ;
        RECT 88.950 562.950 91.050 563.400 ;
        RECT 94.950 564.600 97.050 565.050 ;
        RECT 148.950 564.600 151.050 565.050 ;
        RECT 94.950 563.400 151.050 564.600 ;
        RECT 94.950 562.950 97.050 563.400 ;
        RECT 137.400 562.050 138.600 563.400 ;
        RECT 148.950 562.950 151.050 563.400 ;
        RECT 211.950 564.600 214.050 565.050 ;
        RECT 244.950 564.600 247.050 565.050 ;
        RECT 211.950 563.400 247.050 564.600 ;
        RECT 211.950 562.950 214.050 563.400 ;
        RECT 244.950 562.950 247.050 563.400 ;
        RECT 283.950 564.600 286.050 565.050 ;
        RECT 292.950 564.600 295.050 565.050 ;
        RECT 283.950 563.400 295.050 564.600 ;
        RECT 283.950 562.950 286.050 563.400 ;
        RECT 292.950 562.950 295.050 563.400 ;
        RECT 472.950 564.600 475.050 565.050 ;
        RECT 526.950 564.600 529.050 565.050 ;
        RECT 541.950 564.600 544.050 565.050 ;
        RECT 472.950 563.400 544.050 564.600 ;
        RECT 472.950 562.950 475.050 563.400 ;
        RECT 526.950 562.950 529.050 563.400 ;
        RECT 541.950 562.950 544.050 563.400 ;
        RECT 673.950 564.600 676.050 565.050 ;
        RECT 679.950 564.600 682.050 565.050 ;
        RECT 703.950 564.600 706.050 565.050 ;
        RECT 673.950 563.400 706.050 564.600 ;
        RECT 673.950 562.950 676.050 563.400 ;
        RECT 679.950 562.950 682.050 563.400 ;
        RECT 703.950 562.950 706.050 563.400 ;
        RECT 10.950 559.950 13.050 562.050 ;
        RECT 19.950 559.950 22.050 562.050 ;
        RECT 58.950 561.600 61.050 562.050 ;
        RECT 76.950 561.600 79.050 562.050 ;
        RECT 58.950 560.400 79.050 561.600 ;
        RECT 58.950 559.950 61.050 560.400 ;
        RECT 76.950 559.950 79.050 560.400 ;
        RECT 101.400 560.400 126.600 561.600 ;
        RECT 7.950 556.950 10.050 559.050 ;
        RECT 8.400 553.050 9.600 556.950 ;
        RECT 11.400 556.050 12.600 559.950 ;
        RECT 16.950 556.950 19.050 559.050 ;
        RECT 10.950 553.950 13.050 556.050 ;
        RECT 17.400 553.050 18.600 556.950 ;
        RECT 20.400 555.600 21.600 559.950 ;
        RECT 22.950 558.600 25.050 559.050 ;
        RECT 31.950 558.600 34.050 559.050 ;
        RECT 22.950 557.400 34.050 558.600 ;
        RECT 22.950 556.950 25.050 557.400 ;
        RECT 31.950 556.950 34.050 557.400 ;
        RECT 43.950 556.950 46.050 559.050 ;
        RECT 49.950 556.950 52.050 559.050 ;
        RECT 52.950 558.600 55.050 559.050 ;
        RECT 73.950 558.600 76.050 559.050 ;
        RECT 52.950 557.400 76.050 558.600 ;
        RECT 52.950 556.950 55.050 557.400 ;
        RECT 73.950 556.950 76.050 557.400 ;
        RECT 22.950 555.600 25.050 556.050 ;
        RECT 44.400 555.600 45.600 556.950 ;
        RECT 20.400 554.400 25.050 555.600 ;
        RECT 22.950 553.950 25.050 554.400 ;
        RECT 35.400 554.400 45.600 555.600 ;
        RECT 50.400 555.600 51.600 556.950 ;
        RECT 77.400 556.050 78.600 559.950 ;
        RECT 85.950 558.600 88.050 559.050 ;
        RECT 101.400 558.600 102.600 560.400 ;
        RECT 85.950 557.400 102.600 558.600 ;
        RECT 85.950 556.950 88.050 557.400 ;
        RECT 103.950 556.950 106.050 559.050 ;
        RECT 109.950 558.600 112.050 559.050 ;
        RECT 118.950 558.600 121.050 559.050 ;
        RECT 109.950 557.400 121.050 558.600 ;
        RECT 125.400 558.600 126.600 560.400 ;
        RECT 136.950 559.950 139.050 562.050 ;
        RECT 154.950 561.600 157.050 562.050 ;
        RECT 160.950 561.600 163.050 562.050 ;
        RECT 143.400 560.400 153.600 561.600 ;
        RECT 143.400 558.600 144.600 560.400 ;
        RECT 125.400 557.400 144.600 558.600 ;
        RECT 109.950 556.950 112.050 557.400 ;
        RECT 118.950 556.950 121.050 557.400 ;
        RECT 145.950 556.950 148.050 559.050 ;
        RECT 152.400 558.600 153.600 560.400 ;
        RECT 154.950 560.400 163.050 561.600 ;
        RECT 154.950 559.950 157.050 560.400 ;
        RECT 160.950 559.950 163.050 560.400 ;
        RECT 166.950 561.600 169.050 562.050 ;
        RECT 205.950 561.600 208.050 562.050 ;
        RECT 235.950 561.600 238.050 562.050 ;
        RECT 166.950 560.400 238.050 561.600 ;
        RECT 166.950 559.950 169.050 560.400 ;
        RECT 205.950 559.950 208.050 560.400 ;
        RECT 235.950 559.950 238.050 560.400 ;
        RECT 289.950 559.950 292.050 562.050 ;
        RECT 295.950 561.600 298.050 562.050 ;
        RECT 322.950 561.600 325.050 562.050 ;
        RECT 295.950 560.400 325.050 561.600 ;
        RECT 295.950 559.950 298.050 560.400 ;
        RECT 322.950 559.950 325.050 560.400 ;
        RECT 490.950 561.600 493.050 562.050 ;
        RECT 508.950 561.600 511.050 562.050 ;
        RECT 490.950 560.400 511.050 561.600 ;
        RECT 490.950 559.950 493.050 560.400 ;
        RECT 508.950 559.950 511.050 560.400 ;
        RECT 529.950 561.600 532.050 562.050 ;
        RECT 535.950 561.600 538.050 562.050 ;
        RECT 637.950 561.600 640.050 562.050 ;
        RECT 529.950 560.400 538.050 561.600 ;
        RECT 529.950 559.950 532.050 560.400 ;
        RECT 535.950 559.950 538.050 560.400 ;
        RECT 632.400 560.400 640.050 561.600 ;
        RECT 157.950 558.600 160.050 559.050 ;
        RECT 152.400 557.400 160.050 558.600 ;
        RECT 157.950 556.950 160.050 557.400 ;
        RECT 163.950 558.600 166.050 559.050 ;
        RECT 178.950 558.600 181.050 559.050 ;
        RECT 163.950 557.400 181.050 558.600 ;
        RECT 163.950 556.950 166.050 557.400 ;
        RECT 178.950 556.950 181.050 557.400 ;
        RECT 190.950 558.600 193.050 559.050 ;
        RECT 202.950 558.600 205.050 559.050 ;
        RECT 190.950 557.400 205.050 558.600 ;
        RECT 190.950 556.950 193.050 557.400 ;
        RECT 202.950 556.950 205.050 557.400 ;
        RECT 214.950 558.600 217.050 559.050 ;
        RECT 223.950 558.600 226.050 559.050 ;
        RECT 214.950 557.400 226.050 558.600 ;
        RECT 214.950 556.950 217.050 557.400 ;
        RECT 223.950 556.950 226.050 557.400 ;
        RECT 229.950 558.600 232.050 559.050 ;
        RECT 238.950 558.600 241.050 559.050 ;
        RECT 229.950 557.400 241.050 558.600 ;
        RECT 229.950 556.950 232.050 557.400 ;
        RECT 238.950 556.950 241.050 557.400 ;
        RECT 250.950 556.950 253.050 559.050 ;
        RECT 262.950 556.950 265.050 559.050 ;
        RECT 290.400 558.600 291.600 559.950 ;
        RECT 307.950 558.600 310.050 559.050 ;
        RECT 290.400 557.400 310.050 558.600 ;
        RECT 307.950 556.950 310.050 557.400 ;
        RECT 346.950 558.600 349.050 559.050 ;
        RECT 394.950 558.600 397.050 559.050 ;
        RECT 346.950 557.400 397.050 558.600 ;
        RECT 346.950 556.950 349.050 557.400 ;
        RECT 394.950 556.950 397.050 557.400 ;
        RECT 400.950 556.950 403.050 559.050 ;
        RECT 445.950 556.950 448.050 559.050 ;
        RECT 472.950 556.950 475.050 559.050 ;
        RECT 481.950 558.600 484.050 559.050 ;
        RECT 490.950 558.600 493.050 559.050 ;
        RECT 481.950 557.400 493.050 558.600 ;
        RECT 481.950 556.950 484.050 557.400 ;
        RECT 490.950 556.950 493.050 557.400 ;
        RECT 493.950 558.600 496.050 559.050 ;
        RECT 496.950 558.600 499.050 559.050 ;
        RECT 493.950 557.400 499.050 558.600 ;
        RECT 493.950 556.950 496.050 557.400 ;
        RECT 496.950 556.950 499.050 557.400 ;
        RECT 499.950 558.600 502.050 559.050 ;
        RECT 499.950 557.400 516.600 558.600 ;
        RECT 499.950 556.950 502.050 557.400 ;
        RECT 52.950 555.600 55.050 556.050 ;
        RECT 50.400 554.400 55.050 555.600 ;
        RECT 35.400 553.050 36.600 554.400 ;
        RECT 52.950 553.950 55.050 554.400 ;
        RECT 76.950 553.950 79.050 556.050 ;
        RECT 79.950 555.600 82.050 556.050 ;
        RECT 85.950 555.600 88.050 556.050 ;
        RECT 79.950 554.400 88.050 555.600 ;
        RECT 79.950 553.950 82.050 554.400 ;
        RECT 85.950 553.950 88.050 554.400 ;
        RECT 100.950 553.950 103.050 556.050 ;
        RECT 7.950 550.950 10.050 553.050 ;
        RECT 16.950 550.950 19.050 553.050 ;
        RECT 34.950 550.950 37.050 553.050 ;
        RECT 37.950 552.600 40.050 553.050 ;
        RECT 46.950 552.600 49.050 553.050 ;
        RECT 61.950 552.600 64.050 553.050 ;
        RECT 101.400 552.600 102.600 553.950 ;
        RECT 104.400 553.050 105.600 556.950 ;
        RECT 112.950 555.600 115.050 556.050 ;
        RECT 139.950 555.600 142.050 556.050 ;
        RECT 112.950 554.400 142.050 555.600 ;
        RECT 146.400 555.600 147.600 556.950 ;
        RECT 151.950 555.600 154.050 556.050 ;
        RECT 146.400 554.400 154.050 555.600 ;
        RECT 112.950 553.950 115.050 554.400 ;
        RECT 139.950 553.950 142.050 554.400 ;
        RECT 151.950 553.950 154.050 554.400 ;
        RECT 157.950 555.600 160.050 556.050 ;
        RECT 169.950 555.600 172.050 556.050 ;
        RECT 157.950 554.400 172.050 555.600 ;
        RECT 157.950 553.950 160.050 554.400 ;
        RECT 169.950 553.950 172.050 554.400 ;
        RECT 220.950 555.600 223.050 556.050 ;
        RECT 226.950 555.600 229.050 556.050 ;
        RECT 220.950 554.400 229.050 555.600 ;
        RECT 220.950 553.950 223.050 554.400 ;
        RECT 226.950 553.950 229.050 554.400 ;
        RECT 232.950 555.600 235.050 556.050 ;
        RECT 251.400 555.600 252.600 556.950 ;
        RECT 232.950 554.400 252.600 555.600 ;
        RECT 253.950 555.600 256.050 556.050 ;
        RECT 256.950 555.600 259.050 556.050 ;
        RECT 259.950 555.600 262.050 556.050 ;
        RECT 253.950 554.400 262.050 555.600 ;
        RECT 232.950 553.950 235.050 554.400 ;
        RECT 253.950 553.950 256.050 554.400 ;
        RECT 256.950 553.950 259.050 554.400 ;
        RECT 259.950 553.950 262.050 554.400 ;
        RECT 263.400 553.050 264.600 556.950 ;
        RECT 265.950 555.600 268.050 556.050 ;
        RECT 271.950 555.600 274.050 556.050 ;
        RECT 292.950 555.600 295.050 556.050 ;
        RECT 265.950 554.400 295.050 555.600 ;
        RECT 265.950 553.950 268.050 554.400 ;
        RECT 271.950 553.950 274.050 554.400 ;
        RECT 292.950 553.950 295.050 554.400 ;
        RECT 373.950 555.600 376.050 556.050 ;
        RECT 379.950 555.600 382.050 556.050 ;
        RECT 391.950 555.600 394.050 556.050 ;
        RECT 373.950 554.400 394.050 555.600 ;
        RECT 373.950 553.950 376.050 554.400 ;
        RECT 379.950 553.950 382.050 554.400 ;
        RECT 391.950 553.950 394.050 554.400 ;
        RECT 401.400 553.050 402.600 556.950 ;
        RECT 406.950 555.600 409.050 556.050 ;
        RECT 430.950 555.600 433.050 556.050 ;
        RECT 406.950 554.400 433.050 555.600 ;
        RECT 406.950 553.950 409.050 554.400 ;
        RECT 430.950 553.950 433.050 554.400 ;
        RECT 436.950 555.600 439.050 556.050 ;
        RECT 446.400 555.600 447.600 556.950 ;
        RECT 436.950 554.400 447.600 555.600 ;
        RECT 473.400 555.600 474.600 556.950 ;
        RECT 487.950 555.600 490.050 556.050 ;
        RECT 473.400 554.400 490.050 555.600 ;
        RECT 497.400 555.600 498.600 556.950 ;
        RECT 497.400 554.400 501.600 555.600 ;
        RECT 436.950 553.950 439.050 554.400 ;
        RECT 487.950 553.950 490.050 554.400 ;
        RECT 37.950 551.400 102.600 552.600 ;
        RECT 37.950 550.950 40.050 551.400 ;
        RECT 46.950 550.950 49.050 551.400 ;
        RECT 61.950 550.950 64.050 551.400 ;
        RECT 103.950 550.950 106.050 553.050 ;
        RECT 124.950 552.600 127.050 553.050 ;
        RECT 136.950 552.600 139.050 553.050 ;
        RECT 124.950 551.400 139.050 552.600 ;
        RECT 124.950 550.950 127.050 551.400 ;
        RECT 136.950 550.950 139.050 551.400 ;
        RECT 139.950 552.600 142.050 553.050 ;
        RECT 145.950 552.600 148.050 553.050 ;
        RECT 139.950 551.400 148.050 552.600 ;
        RECT 139.950 550.950 142.050 551.400 ;
        RECT 145.950 550.950 148.050 551.400 ;
        RECT 160.950 552.600 163.050 553.050 ;
        RECT 175.950 552.600 178.050 553.050 ;
        RECT 160.950 551.400 178.050 552.600 ;
        RECT 160.950 550.950 163.050 551.400 ;
        RECT 175.950 550.950 178.050 551.400 ;
        RECT 181.950 552.600 184.050 553.050 ;
        RECT 187.950 552.600 190.050 553.050 ;
        RECT 181.950 551.400 190.050 552.600 ;
        RECT 181.950 550.950 184.050 551.400 ;
        RECT 187.950 550.950 190.050 551.400 ;
        RECT 208.950 552.600 211.050 553.050 ;
        RECT 211.950 552.600 214.050 553.050 ;
        RECT 217.950 552.600 220.050 553.050 ;
        RECT 208.950 551.400 220.050 552.600 ;
        RECT 208.950 550.950 211.050 551.400 ;
        RECT 211.950 550.950 214.050 551.400 ;
        RECT 217.950 550.950 220.050 551.400 ;
        RECT 235.950 552.600 238.050 553.050 ;
        RECT 241.950 552.600 244.050 553.050 ;
        RECT 247.950 552.600 250.050 553.050 ;
        RECT 235.950 551.400 250.050 552.600 ;
        RECT 235.950 550.950 238.050 551.400 ;
        RECT 241.950 550.950 244.050 551.400 ;
        RECT 247.950 550.950 250.050 551.400 ;
        RECT 262.950 550.950 265.050 553.050 ;
        RECT 280.950 552.600 283.050 553.050 ;
        RECT 286.950 552.600 289.050 553.050 ;
        RECT 280.950 551.400 289.050 552.600 ;
        RECT 280.950 550.950 283.050 551.400 ;
        RECT 286.950 550.950 289.050 551.400 ;
        RECT 292.950 552.600 295.050 553.050 ;
        RECT 298.950 552.600 301.050 553.050 ;
        RECT 292.950 551.400 301.050 552.600 ;
        RECT 292.950 550.950 295.050 551.400 ;
        RECT 298.950 550.950 301.050 551.400 ;
        RECT 367.950 552.600 370.050 553.050 ;
        RECT 397.950 552.600 400.050 553.050 ;
        RECT 367.950 551.400 400.050 552.600 ;
        RECT 367.950 550.950 370.050 551.400 ;
        RECT 397.950 550.950 400.050 551.400 ;
        RECT 400.950 550.950 403.050 553.050 ;
        RECT 412.950 552.600 415.050 553.050 ;
        RECT 418.950 552.600 421.050 553.050 ;
        RECT 412.950 551.400 421.050 552.600 ;
        RECT 412.950 550.950 415.050 551.400 ;
        RECT 418.950 550.950 421.050 551.400 ;
        RECT 433.950 552.600 436.050 553.050 ;
        RECT 442.950 552.600 445.050 553.050 ;
        RECT 433.950 551.400 445.050 552.600 ;
        RECT 433.950 550.950 436.050 551.400 ;
        RECT 442.950 550.950 445.050 551.400 ;
        RECT 460.950 552.600 463.050 553.050 ;
        RECT 478.950 552.600 481.050 553.050 ;
        RECT 460.950 551.400 481.050 552.600 ;
        RECT 500.400 552.600 501.600 554.400 ;
        RECT 515.400 553.050 516.600 557.400 ;
        RECT 556.950 556.950 559.050 559.050 ;
        RECT 583.950 558.600 586.050 559.050 ;
        RECT 628.950 558.600 631.050 559.050 ;
        RECT 583.950 557.400 631.050 558.600 ;
        RECT 583.950 556.950 586.050 557.400 ;
        RECT 628.950 556.950 631.050 557.400 ;
        RECT 532.950 555.600 535.050 556.050 ;
        RECT 557.400 555.600 558.600 556.950 ;
        RECT 532.950 554.400 558.600 555.600 ;
        RECT 559.950 555.600 562.050 556.050 ;
        RECT 580.950 555.600 583.050 556.050 ;
        RECT 632.400 555.600 633.600 560.400 ;
        RECT 637.950 559.950 640.050 560.400 ;
        RECT 634.950 558.600 637.050 559.050 ;
        RECT 640.950 558.600 643.050 559.050 ;
        RECT 634.950 557.400 643.050 558.600 ;
        RECT 634.950 556.950 637.050 557.400 ;
        RECT 640.950 556.950 643.050 557.400 ;
        RECT 694.950 558.600 697.050 559.050 ;
        RECT 715.950 558.600 718.050 559.050 ;
        RECT 694.950 557.400 718.050 558.600 ;
        RECT 694.950 556.950 697.050 557.400 ;
        RECT 715.950 556.950 718.050 557.400 ;
        RECT 559.950 554.400 583.050 555.600 ;
        RECT 532.950 553.950 535.050 554.400 ;
        RECT 559.950 553.950 562.050 554.400 ;
        RECT 580.950 553.950 583.050 554.400 ;
        RECT 629.400 554.400 633.600 555.600 ;
        RECT 637.950 555.600 640.050 556.050 ;
        RECT 664.950 555.600 667.050 556.050 ;
        RECT 637.950 554.400 667.050 555.600 ;
        RECT 629.400 553.050 630.600 554.400 ;
        RECT 637.950 553.950 640.050 554.400 ;
        RECT 664.950 553.950 667.050 554.400 ;
        RECT 505.950 552.600 508.050 553.050 ;
        RECT 500.400 551.400 508.050 552.600 ;
        RECT 460.950 550.950 463.050 551.400 ;
        RECT 478.950 550.950 481.050 551.400 ;
        RECT 505.950 550.950 508.050 551.400 ;
        RECT 514.950 550.950 517.050 553.050 ;
        RECT 628.950 550.950 631.050 553.050 ;
        RECT 10.950 549.600 13.050 550.050 ;
        RECT 19.950 549.600 22.050 550.050 ;
        RECT 10.950 548.400 22.050 549.600 ;
        RECT 10.950 547.950 13.050 548.400 ;
        RECT 19.950 547.950 22.050 548.400 ;
        RECT 25.950 549.600 28.050 550.050 ;
        RECT 55.950 549.600 58.050 550.050 ;
        RECT 25.950 548.400 58.050 549.600 ;
        RECT 25.950 547.950 28.050 548.400 ;
        RECT 55.950 547.950 58.050 548.400 ;
        RECT 76.950 549.600 79.050 550.050 ;
        RECT 139.950 549.600 142.050 550.050 ;
        RECT 76.950 548.400 142.050 549.600 ;
        RECT 76.950 547.950 79.050 548.400 ;
        RECT 139.950 547.950 142.050 548.400 ;
        RECT 187.950 549.600 190.050 550.050 ;
        RECT 232.950 549.600 235.050 550.050 ;
        RECT 187.950 548.400 235.050 549.600 ;
        RECT 187.950 547.950 190.050 548.400 ;
        RECT 232.950 547.950 235.050 548.400 ;
        RECT 274.950 549.600 277.050 550.050 ;
        RECT 358.950 549.600 361.050 550.050 ;
        RECT 274.950 548.400 361.050 549.600 ;
        RECT 274.950 547.950 277.050 548.400 ;
        RECT 358.950 547.950 361.050 548.400 ;
        RECT 388.950 549.600 391.050 550.050 ;
        RECT 412.950 549.600 415.050 550.050 ;
        RECT 388.950 548.400 415.050 549.600 ;
        RECT 388.950 547.950 391.050 548.400 ;
        RECT 412.950 547.950 415.050 548.400 ;
        RECT 442.950 549.600 445.050 550.050 ;
        RECT 466.950 549.600 469.050 550.050 ;
        RECT 502.950 549.600 505.050 550.050 ;
        RECT 442.950 548.400 505.050 549.600 ;
        RECT 442.950 547.950 445.050 548.400 ;
        RECT 466.950 547.950 469.050 548.400 ;
        RECT 502.950 547.950 505.050 548.400 ;
        RECT 517.950 549.600 520.050 550.050 ;
        RECT 571.950 549.600 574.050 550.050 ;
        RECT 517.950 548.400 574.050 549.600 ;
        RECT 517.950 547.950 520.050 548.400 ;
        RECT 571.950 547.950 574.050 548.400 ;
        RECT 616.950 549.600 619.050 550.050 ;
        RECT 631.950 549.600 634.050 550.050 ;
        RECT 616.950 548.400 634.050 549.600 ;
        RECT 616.950 547.950 619.050 548.400 ;
        RECT 631.950 547.950 634.050 548.400 ;
        RECT 7.950 546.600 10.050 547.050 ;
        RECT 13.950 546.600 16.050 547.050 ;
        RECT 7.950 545.400 16.050 546.600 ;
        RECT 7.950 544.950 10.050 545.400 ;
        RECT 13.950 544.950 16.050 545.400 ;
        RECT 34.950 546.600 37.050 547.050 ;
        RECT 46.950 546.600 49.050 547.050 ;
        RECT 34.950 545.400 49.050 546.600 ;
        RECT 34.950 544.950 37.050 545.400 ;
        RECT 46.950 544.950 49.050 545.400 ;
        RECT 64.950 546.600 67.050 547.050 ;
        RECT 67.950 546.600 70.050 547.050 ;
        RECT 118.950 546.600 121.050 547.050 ;
        RECT 64.950 545.400 121.050 546.600 ;
        RECT 64.950 544.950 67.050 545.400 ;
        RECT 67.950 544.950 70.050 545.400 ;
        RECT 118.950 544.950 121.050 545.400 ;
        RECT 160.950 546.600 163.050 547.050 ;
        RECT 205.950 546.600 208.050 547.050 ;
        RECT 244.950 546.600 247.050 547.050 ;
        RECT 286.950 546.600 289.050 547.050 ;
        RECT 160.950 545.400 289.050 546.600 ;
        RECT 160.950 544.950 163.050 545.400 ;
        RECT 205.950 544.950 208.050 545.400 ;
        RECT 244.950 544.950 247.050 545.400 ;
        RECT 286.950 544.950 289.050 545.400 ;
        RECT 421.950 546.600 424.050 547.050 ;
        RECT 448.950 546.600 451.050 547.050 ;
        RECT 469.950 546.600 472.050 547.050 ;
        RECT 421.950 545.400 472.050 546.600 ;
        RECT 421.950 544.950 424.050 545.400 ;
        RECT 448.950 544.950 451.050 545.400 ;
        RECT 469.950 544.950 472.050 545.400 ;
        RECT 508.950 546.600 511.050 547.050 ;
        RECT 544.950 546.600 547.050 547.050 ;
        RECT 508.950 545.400 547.050 546.600 ;
        RECT 508.950 544.950 511.050 545.400 ;
        RECT 544.950 544.950 547.050 545.400 ;
        RECT 625.950 546.600 628.050 547.050 ;
        RECT 643.950 546.600 646.050 547.050 ;
        RECT 625.950 545.400 646.050 546.600 ;
        RECT 625.950 544.950 628.050 545.400 ;
        RECT 643.950 544.950 646.050 545.400 ;
        RECT 4.950 543.600 7.050 544.050 ;
        RECT 13.950 543.600 16.050 544.050 ;
        RECT 4.950 542.400 16.050 543.600 ;
        RECT 4.950 541.950 7.050 542.400 ;
        RECT 13.950 541.950 16.050 542.400 ;
        RECT 16.950 543.600 19.050 544.050 ;
        RECT 55.950 543.600 58.050 544.050 ;
        RECT 103.950 543.600 106.050 544.050 ;
        RECT 16.950 542.400 106.050 543.600 ;
        RECT 16.950 541.950 19.050 542.400 ;
        RECT 55.950 541.950 58.050 542.400 ;
        RECT 103.950 541.950 106.050 542.400 ;
        RECT 112.950 543.600 115.050 544.050 ;
        RECT 169.950 543.600 172.050 544.050 ;
        RECT 235.950 543.600 238.050 544.050 ;
        RECT 112.950 542.400 238.050 543.600 ;
        RECT 112.950 541.950 115.050 542.400 ;
        RECT 169.950 541.950 172.050 542.400 ;
        RECT 235.950 541.950 238.050 542.400 ;
        RECT 289.950 543.600 292.050 544.050 ;
        RECT 355.950 543.600 358.050 544.050 ;
        RECT 289.950 542.400 358.050 543.600 ;
        RECT 289.950 541.950 292.050 542.400 ;
        RECT 355.950 541.950 358.050 542.400 ;
        RECT 415.950 543.600 418.050 544.050 ;
        RECT 436.950 543.600 439.050 544.050 ;
        RECT 415.950 542.400 439.050 543.600 ;
        RECT 415.950 541.950 418.050 542.400 ;
        RECT 436.950 541.950 439.050 542.400 ;
        RECT 493.950 543.600 496.050 544.050 ;
        RECT 511.950 543.600 514.050 544.050 ;
        RECT 514.950 543.600 517.050 544.050 ;
        RECT 493.950 542.400 517.050 543.600 ;
        RECT 493.950 541.950 496.050 542.400 ;
        RECT 511.950 541.950 514.050 542.400 ;
        RECT 514.950 541.950 517.050 542.400 ;
        RECT 622.950 543.600 625.050 544.050 ;
        RECT 640.950 543.600 643.050 544.050 ;
        RECT 622.950 542.400 643.050 543.600 ;
        RECT 622.950 541.950 625.050 542.400 ;
        RECT 640.950 541.950 643.050 542.400 ;
        RECT 646.950 543.600 649.050 544.050 ;
        RECT 661.950 543.600 664.050 544.050 ;
        RECT 646.950 542.400 664.050 543.600 ;
        RECT 646.950 541.950 649.050 542.400 ;
        RECT 661.950 541.950 664.050 542.400 ;
        RECT 16.950 540.600 19.050 541.050 ;
        RECT 97.950 540.600 100.050 541.050 ;
        RECT 160.950 540.600 163.050 541.050 ;
        RECT 16.950 539.400 96.600 540.600 ;
        RECT 16.950 538.950 19.050 539.400 ;
        RECT 49.950 537.600 52.050 538.050 ;
        RECT 52.950 537.600 55.050 538.050 ;
        RECT 79.950 537.600 82.050 538.050 ;
        RECT 88.950 537.600 91.050 538.050 ;
        RECT 49.950 536.400 91.050 537.600 ;
        RECT 95.400 537.600 96.600 539.400 ;
        RECT 97.950 539.400 163.050 540.600 ;
        RECT 97.950 538.950 100.050 539.400 ;
        RECT 160.950 538.950 163.050 539.400 ;
        RECT 163.950 540.600 166.050 541.050 ;
        RECT 229.950 540.600 232.050 541.050 ;
        RECT 163.950 539.400 232.050 540.600 ;
        RECT 163.950 538.950 166.050 539.400 ;
        RECT 229.950 538.950 232.050 539.400 ;
        RECT 298.950 540.600 301.050 541.050 ;
        RECT 322.950 540.600 325.050 541.050 ;
        RECT 346.950 540.600 349.050 541.050 ;
        RECT 298.950 539.400 349.050 540.600 ;
        RECT 298.950 538.950 301.050 539.400 ;
        RECT 322.950 538.950 325.050 539.400 ;
        RECT 346.950 538.950 349.050 539.400 ;
        RECT 457.950 540.600 460.050 541.050 ;
        RECT 523.950 540.600 526.050 541.050 ;
        RECT 538.950 540.600 541.050 541.050 ;
        RECT 457.950 539.400 541.050 540.600 ;
        RECT 457.950 538.950 460.050 539.400 ;
        RECT 523.950 538.950 526.050 539.400 ;
        RECT 538.950 538.950 541.050 539.400 ;
        RECT 571.950 540.600 574.050 541.050 ;
        RECT 613.950 540.600 616.050 541.050 ;
        RECT 571.950 539.400 616.050 540.600 ;
        RECT 571.950 538.950 574.050 539.400 ;
        RECT 613.950 538.950 616.050 539.400 ;
        RECT 655.950 540.600 658.050 541.050 ;
        RECT 661.950 540.600 664.050 541.050 ;
        RECT 655.950 539.400 664.050 540.600 ;
        RECT 655.950 538.950 658.050 539.400 ;
        RECT 661.950 538.950 664.050 539.400 ;
        RECT 148.950 537.600 151.050 538.050 ;
        RECT 95.400 536.400 151.050 537.600 ;
        RECT 49.950 535.950 52.050 536.400 ;
        RECT 52.950 535.950 55.050 536.400 ;
        RECT 79.950 535.950 82.050 536.400 ;
        RECT 88.950 535.950 91.050 536.400 ;
        RECT 148.950 535.950 151.050 536.400 ;
        RECT 166.950 537.600 169.050 538.050 ;
        RECT 172.950 537.600 175.050 538.050 ;
        RECT 166.950 536.400 175.050 537.600 ;
        RECT 166.950 535.950 169.050 536.400 ;
        RECT 172.950 535.950 175.050 536.400 ;
        RECT 325.950 537.600 328.050 538.050 ;
        RECT 373.950 537.600 376.050 538.050 ;
        RECT 325.950 536.400 376.050 537.600 ;
        RECT 325.950 535.950 328.050 536.400 ;
        RECT 373.950 535.950 376.050 536.400 ;
        RECT 475.950 537.600 478.050 538.050 ;
        RECT 547.950 537.600 550.050 538.050 ;
        RECT 475.950 536.400 550.050 537.600 ;
        RECT 475.950 535.950 478.050 536.400 ;
        RECT 547.950 535.950 550.050 536.400 ;
        RECT 586.950 537.600 589.050 538.050 ;
        RECT 607.950 537.600 610.050 538.050 ;
        RECT 586.950 536.400 610.050 537.600 ;
        RECT 586.950 535.950 589.050 536.400 ;
        RECT 607.950 535.950 610.050 536.400 ;
        RECT 100.950 534.600 103.050 535.050 ;
        RECT 109.950 534.600 112.050 535.050 ;
        RECT 100.950 533.400 112.050 534.600 ;
        RECT 100.950 532.950 103.050 533.400 ;
        RECT 109.950 532.950 112.050 533.400 ;
        RECT 145.950 534.600 148.050 535.050 ;
        RECT 190.950 534.600 193.050 535.050 ;
        RECT 145.950 533.400 193.050 534.600 ;
        RECT 145.950 532.950 148.050 533.400 ;
        RECT 190.950 532.950 193.050 533.400 ;
        RECT 238.950 534.600 241.050 535.050 ;
        RECT 325.950 534.600 328.050 535.050 ;
        RECT 238.950 533.400 328.050 534.600 ;
        RECT 238.950 532.950 241.050 533.400 ;
        RECT 325.950 532.950 328.050 533.400 ;
        RECT 343.950 534.600 346.050 535.050 ;
        RECT 364.950 534.600 367.050 535.050 ;
        RECT 343.950 533.400 367.050 534.600 ;
        RECT 343.950 532.950 346.050 533.400 ;
        RECT 364.950 532.950 367.050 533.400 ;
        RECT 385.950 534.600 388.050 535.050 ;
        RECT 406.950 534.600 409.050 535.050 ;
        RECT 385.950 533.400 409.050 534.600 ;
        RECT 385.950 532.950 388.050 533.400 ;
        RECT 406.950 532.950 409.050 533.400 ;
        RECT 481.950 534.600 484.050 535.050 ;
        RECT 490.950 534.600 493.050 535.050 ;
        RECT 481.950 533.400 493.050 534.600 ;
        RECT 481.950 532.950 484.050 533.400 ;
        RECT 490.950 532.950 493.050 533.400 ;
        RECT 502.950 534.600 505.050 535.050 ;
        RECT 508.950 534.600 511.050 535.050 ;
        RECT 502.950 533.400 511.050 534.600 ;
        RECT 502.950 532.950 505.050 533.400 ;
        RECT 508.950 532.950 511.050 533.400 ;
        RECT 520.950 534.600 523.050 535.050 ;
        RECT 529.950 534.600 532.050 535.050 ;
        RECT 535.950 534.600 538.050 535.050 ;
        RECT 550.950 534.600 553.050 535.050 ;
        RECT 520.950 533.400 553.050 534.600 ;
        RECT 520.950 532.950 523.050 533.400 ;
        RECT 529.950 532.950 532.050 533.400 ;
        RECT 535.950 532.950 538.050 533.400 ;
        RECT 550.950 532.950 553.050 533.400 ;
        RECT 604.950 534.600 607.050 535.050 ;
        RECT 622.950 534.600 625.050 535.050 ;
        RECT 604.950 533.400 625.050 534.600 ;
        RECT 604.950 532.950 607.050 533.400 ;
        RECT 622.950 532.950 625.050 533.400 ;
        RECT 25.950 531.600 28.050 532.050 ;
        RECT 76.950 531.600 79.050 532.050 ;
        RECT 112.950 531.600 115.050 532.050 ;
        RECT 25.950 530.400 79.050 531.600 ;
        RECT 25.950 529.950 28.050 530.400 ;
        RECT 76.950 529.950 79.050 530.400 ;
        RECT 86.400 530.400 115.050 531.600 ;
        RECT 70.950 528.600 73.050 529.050 ;
        RECT 82.950 528.600 85.050 529.050 ;
        RECT 70.950 527.400 85.050 528.600 ;
        RECT 70.950 526.950 73.050 527.400 ;
        RECT 82.950 526.950 85.050 527.400 ;
        RECT 64.950 525.600 67.050 526.050 ;
        RECT 73.950 525.600 76.050 526.050 ;
        RECT 64.950 524.400 76.050 525.600 ;
        RECT 64.950 523.950 67.050 524.400 ;
        RECT 73.950 523.950 76.050 524.400 ;
        RECT 79.950 525.600 82.050 526.050 ;
        RECT 86.400 525.600 87.600 530.400 ;
        RECT 112.950 529.950 115.050 530.400 ;
        RECT 124.950 531.600 127.050 532.050 ;
        RECT 130.950 531.600 133.050 532.050 ;
        RECT 124.950 530.400 133.050 531.600 ;
        RECT 124.950 529.950 127.050 530.400 ;
        RECT 130.950 529.950 133.050 530.400 ;
        RECT 151.950 531.600 154.050 532.050 ;
        RECT 157.950 531.600 160.050 532.050 ;
        RECT 151.950 530.400 160.050 531.600 ;
        RECT 151.950 529.950 154.050 530.400 ;
        RECT 157.950 529.950 160.050 530.400 ;
        RECT 163.950 531.600 166.050 532.050 ;
        RECT 184.950 531.600 187.050 532.050 ;
        RECT 253.950 531.600 256.050 532.050 ;
        RECT 268.950 531.600 271.050 532.050 ;
        RECT 163.950 530.400 187.050 531.600 ;
        RECT 163.950 529.950 166.050 530.400 ;
        RECT 184.950 529.950 187.050 530.400 ;
        RECT 209.400 530.400 252.600 531.600 ;
        RECT 97.950 526.950 100.050 529.050 ;
        RECT 124.950 526.950 127.050 529.050 ;
        RECT 148.950 528.600 151.050 529.050 ;
        RECT 209.400 528.600 210.600 530.400 ;
        RECT 251.400 529.050 252.600 530.400 ;
        RECT 253.950 530.400 271.050 531.600 ;
        RECT 253.950 529.950 256.050 530.400 ;
        RECT 268.950 529.950 271.050 530.400 ;
        RECT 274.950 531.600 277.050 532.050 ;
        RECT 316.950 531.600 319.050 532.050 ;
        RECT 274.950 530.400 319.050 531.600 ;
        RECT 274.950 529.950 277.050 530.400 ;
        RECT 316.950 529.950 319.050 530.400 ;
        RECT 355.950 531.600 358.050 532.050 ;
        RECT 364.950 531.600 367.050 532.050 ;
        RECT 355.950 530.400 367.050 531.600 ;
        RECT 355.950 529.950 358.050 530.400 ;
        RECT 364.950 529.950 367.050 530.400 ;
        RECT 379.950 531.600 382.050 532.050 ;
        RECT 454.950 531.600 457.050 532.050 ;
        RECT 379.950 530.400 457.050 531.600 ;
        RECT 379.950 529.950 382.050 530.400 ;
        RECT 454.950 529.950 457.050 530.400 ;
        RECT 472.950 531.600 475.050 532.050 ;
        RECT 481.950 531.600 484.050 532.050 ;
        RECT 472.950 530.400 484.050 531.600 ;
        RECT 472.950 529.950 475.050 530.400 ;
        RECT 481.950 529.950 484.050 530.400 ;
        RECT 484.950 531.600 487.050 532.050 ;
        RECT 496.950 531.600 499.050 532.050 ;
        RECT 499.950 531.600 502.050 532.050 ;
        RECT 511.950 531.600 514.050 532.050 ;
        RECT 484.950 530.400 502.050 531.600 ;
        RECT 484.950 529.950 487.050 530.400 ;
        RECT 496.950 529.950 499.050 530.400 ;
        RECT 499.950 529.950 502.050 530.400 ;
        RECT 503.400 530.400 514.050 531.600 ;
        RECT 148.950 527.400 210.600 528.600 ;
        RECT 211.950 528.600 214.050 529.050 ;
        RECT 232.950 528.600 235.050 529.050 ;
        RECT 211.950 527.400 235.050 528.600 ;
        RECT 148.950 526.950 151.050 527.400 ;
        RECT 211.950 526.950 214.050 527.400 ;
        RECT 232.950 526.950 235.050 527.400 ;
        RECT 250.950 526.950 253.050 529.050 ;
        RECT 256.950 528.600 259.050 529.050 ;
        RECT 268.950 528.600 271.050 529.050 ;
        RECT 256.950 527.400 271.050 528.600 ;
        RECT 256.950 526.950 259.050 527.400 ;
        RECT 268.950 526.950 271.050 527.400 ;
        RECT 316.950 528.600 319.050 529.050 ;
        RECT 322.950 528.600 325.050 529.050 ;
        RECT 334.950 528.600 337.050 529.050 ;
        RECT 316.950 527.400 337.050 528.600 ;
        RECT 316.950 526.950 319.050 527.400 ;
        RECT 322.950 526.950 325.050 527.400 ;
        RECT 334.950 526.950 337.050 527.400 ;
        RECT 400.950 528.600 403.050 529.050 ;
        RECT 421.950 528.600 424.050 529.050 ;
        RECT 424.950 528.600 427.050 529.050 ;
        RECT 439.950 528.600 442.050 529.050 ;
        RECT 460.950 528.600 463.050 529.050 ;
        RECT 469.950 528.600 472.050 529.050 ;
        RECT 400.950 527.400 459.600 528.600 ;
        RECT 400.950 526.950 403.050 527.400 ;
        RECT 421.950 526.950 424.050 527.400 ;
        RECT 424.950 526.950 427.050 527.400 ;
        RECT 439.950 526.950 442.050 527.400 ;
        RECT 79.950 524.400 87.600 525.600 ;
        RECT 79.950 523.950 82.050 524.400 ;
        RECT 10.950 522.600 13.050 523.050 ;
        RECT 16.950 522.600 19.050 523.050 ;
        RECT 10.950 521.400 19.050 522.600 ;
        RECT 10.950 520.950 13.050 521.400 ;
        RECT 16.950 520.950 19.050 521.400 ;
        RECT 82.950 522.600 85.050 523.050 ;
        RECT 98.400 522.600 99.600 526.950 ;
        RECT 103.950 523.950 106.050 526.050 ;
        RECT 125.400 525.600 126.600 526.950 ;
        RECT 130.950 525.600 133.050 526.050 ;
        RECT 125.400 524.400 133.050 525.600 ;
        RECT 130.950 523.950 133.050 524.400 ;
        RECT 133.950 525.600 136.050 526.050 ;
        RECT 151.950 525.600 154.050 526.050 ;
        RECT 133.950 524.400 154.050 525.600 ;
        RECT 133.950 523.950 136.050 524.400 ;
        RECT 151.950 523.950 154.050 524.400 ;
        RECT 154.950 525.600 157.050 526.050 ;
        RECT 166.950 525.600 169.050 526.050 ;
        RECT 154.950 524.400 169.050 525.600 ;
        RECT 154.950 523.950 157.050 524.400 ;
        RECT 166.950 523.950 169.050 524.400 ;
        RECT 172.950 525.600 175.050 526.050 ;
        RECT 184.950 525.600 187.050 526.050 ;
        RECT 172.950 524.400 187.050 525.600 ;
        RECT 172.950 523.950 175.050 524.400 ;
        RECT 184.950 523.950 187.050 524.400 ;
        RECT 196.950 525.600 199.050 526.050 ;
        RECT 214.950 525.600 217.050 526.050 ;
        RECT 196.950 524.400 217.050 525.600 ;
        RECT 196.950 523.950 199.050 524.400 ;
        RECT 214.950 523.950 217.050 524.400 ;
        RECT 262.950 525.600 265.050 526.050 ;
        RECT 277.950 525.600 280.050 526.050 ;
        RECT 262.950 524.400 280.050 525.600 ;
        RECT 262.950 523.950 265.050 524.400 ;
        RECT 277.950 523.950 280.050 524.400 ;
        RECT 298.950 525.600 301.050 526.050 ;
        RECT 337.950 525.600 340.050 526.050 ;
        RECT 349.950 525.600 352.050 526.050 ;
        RECT 298.950 524.400 318.600 525.600 ;
        RECT 298.950 523.950 301.050 524.400 ;
        RECT 82.950 521.400 99.600 522.600 ;
        RECT 82.950 520.950 85.050 521.400 ;
        RECT 104.400 520.050 105.600 523.950 ;
        RECT 317.400 523.050 318.600 524.400 ;
        RECT 337.950 524.400 352.050 525.600 ;
        RECT 337.950 523.950 340.050 524.400 ;
        RECT 349.950 523.950 352.050 524.400 ;
        RECT 358.950 525.600 361.050 526.050 ;
        RECT 403.950 525.600 406.050 526.050 ;
        RECT 358.950 524.400 406.050 525.600 ;
        RECT 358.950 523.950 361.050 524.400 ;
        RECT 403.950 523.950 406.050 524.400 ;
        RECT 409.950 525.600 412.050 526.050 ;
        RECT 430.950 525.600 433.050 526.050 ;
        RECT 409.950 524.400 433.050 525.600 ;
        RECT 458.400 525.600 459.600 527.400 ;
        RECT 460.950 527.400 472.050 528.600 ;
        RECT 460.950 526.950 463.050 527.400 ;
        RECT 469.950 526.950 472.050 527.400 ;
        RECT 475.950 528.600 478.050 529.050 ;
        RECT 487.950 528.600 490.050 529.050 ;
        RECT 503.400 528.600 504.600 530.400 ;
        RECT 511.950 529.950 514.050 530.400 ;
        RECT 514.950 531.600 517.050 532.050 ;
        RECT 520.950 531.600 523.050 532.050 ;
        RECT 526.950 531.600 529.050 532.050 ;
        RECT 547.950 531.600 550.050 532.050 ;
        RECT 514.950 530.400 519.600 531.600 ;
        RECT 514.950 529.950 517.050 530.400 ;
        RECT 475.950 527.400 490.050 528.600 ;
        RECT 475.950 526.950 478.050 527.400 ;
        RECT 487.950 526.950 490.050 527.400 ;
        RECT 500.400 527.400 504.600 528.600 ;
        RECT 518.400 528.600 519.600 530.400 ;
        RECT 520.950 530.400 529.050 531.600 ;
        RECT 520.950 529.950 523.050 530.400 ;
        RECT 526.950 529.950 529.050 530.400 ;
        RECT 533.400 530.400 550.050 531.600 ;
        RECT 518.400 527.400 525.600 528.600 ;
        RECT 478.950 525.600 481.050 526.050 ;
        RECT 458.400 524.400 481.050 525.600 ;
        RECT 409.950 523.950 412.050 524.400 ;
        RECT 430.950 523.950 433.050 524.400 ;
        RECT 478.950 523.950 481.050 524.400 ;
        RECT 484.950 525.600 487.050 526.050 ;
        RECT 500.400 525.600 501.600 527.400 ;
        RECT 484.950 524.400 501.600 525.600 ;
        RECT 508.950 525.600 511.050 526.050 ;
        RECT 514.950 525.600 517.050 526.050 ;
        RECT 508.950 524.400 517.050 525.600 ;
        RECT 484.950 523.950 487.050 524.400 ;
        RECT 508.950 523.950 511.050 524.400 ;
        RECT 514.950 523.950 517.050 524.400 ;
        RECT 524.400 523.050 525.600 527.400 ;
        RECT 533.400 526.050 534.600 530.400 ;
        RECT 547.950 529.950 550.050 530.400 ;
        RECT 562.950 531.600 565.050 532.050 ;
        RECT 586.950 531.600 589.050 532.050 ;
        RECT 562.950 530.400 589.050 531.600 ;
        RECT 562.950 529.950 565.050 530.400 ;
        RECT 586.950 529.950 589.050 530.400 ;
        RECT 592.950 531.600 595.050 532.050 ;
        RECT 604.950 531.600 607.050 532.050 ;
        RECT 592.950 530.400 607.050 531.600 ;
        RECT 592.950 529.950 595.050 530.400 ;
        RECT 604.950 529.950 607.050 530.400 ;
        RECT 541.950 528.600 544.050 529.050 ;
        RECT 577.950 528.600 580.050 529.050 ;
        RECT 592.950 528.600 595.050 529.050 ;
        RECT 541.950 527.400 570.600 528.600 ;
        RECT 541.950 526.950 544.050 527.400 ;
        RECT 569.400 526.050 570.600 527.400 ;
        RECT 577.950 527.400 595.050 528.600 ;
        RECT 577.950 526.950 580.050 527.400 ;
        RECT 592.950 526.950 595.050 527.400 ;
        RECT 607.950 528.600 610.050 529.050 ;
        RECT 643.950 528.600 646.050 529.050 ;
        RECT 658.950 528.600 661.050 529.050 ;
        RECT 607.950 527.400 661.050 528.600 ;
        RECT 607.950 526.950 610.050 527.400 ;
        RECT 643.950 526.950 646.050 527.400 ;
        RECT 658.950 526.950 661.050 527.400 ;
        RECT 670.950 528.600 673.050 529.050 ;
        RECT 694.950 528.600 697.050 529.050 ;
        RECT 670.950 527.400 697.050 528.600 ;
        RECT 670.950 526.950 673.050 527.400 ;
        RECT 694.950 526.950 697.050 527.400 ;
        RECT 700.950 526.950 703.050 529.050 ;
        RECT 532.950 523.950 535.050 526.050 ;
        RECT 556.950 525.600 559.050 526.050 ;
        RECT 562.950 525.600 565.050 526.050 ;
        RECT 556.950 524.400 565.050 525.600 ;
        RECT 556.950 523.950 559.050 524.400 ;
        RECT 562.950 523.950 565.050 524.400 ;
        RECT 568.950 523.950 571.050 526.050 ;
        RECT 658.950 525.600 661.050 526.050 ;
        RECT 667.950 525.600 670.050 526.050 ;
        RECT 658.950 524.400 670.050 525.600 ;
        RECT 658.950 523.950 661.050 524.400 ;
        RECT 667.950 523.950 670.050 524.400 ;
        RECT 682.950 525.600 685.050 526.050 ;
        RECT 697.950 525.600 700.050 526.050 ;
        RECT 682.950 524.400 700.050 525.600 ;
        RECT 682.950 523.950 685.050 524.400 ;
        RECT 697.950 523.950 700.050 524.400 ;
        RECT 701.400 523.050 702.600 526.950 ;
        RECT 703.950 525.600 706.050 526.050 ;
        RECT 712.950 525.600 715.050 526.050 ;
        RECT 703.950 524.400 715.050 525.600 ;
        RECT 703.950 523.950 706.050 524.400 ;
        RECT 712.950 523.950 715.050 524.400 ;
        RECT 148.950 522.600 151.050 523.050 ;
        RECT 154.950 522.600 157.050 523.050 ;
        RECT 148.950 521.400 157.050 522.600 ;
        RECT 148.950 520.950 151.050 521.400 ;
        RECT 154.950 520.950 157.050 521.400 ;
        RECT 163.950 522.600 166.050 523.050 ;
        RECT 178.950 522.600 181.050 523.050 ;
        RECT 163.950 521.400 181.050 522.600 ;
        RECT 163.950 520.950 166.050 521.400 ;
        RECT 178.950 520.950 181.050 521.400 ;
        RECT 199.950 522.600 202.050 523.050 ;
        RECT 205.950 522.600 208.050 523.050 ;
        RECT 199.950 521.400 208.050 522.600 ;
        RECT 199.950 520.950 202.050 521.400 ;
        RECT 205.950 520.950 208.050 521.400 ;
        RECT 238.950 522.600 241.050 523.050 ;
        RECT 250.950 522.600 253.050 523.050 ;
        RECT 283.950 522.600 286.050 523.050 ;
        RECT 238.950 521.400 286.050 522.600 ;
        RECT 238.950 520.950 241.050 521.400 ;
        RECT 250.950 520.950 253.050 521.400 ;
        RECT 283.950 520.950 286.050 521.400 ;
        RECT 286.950 522.600 289.050 523.050 ;
        RECT 292.950 522.600 295.050 523.050 ;
        RECT 295.950 522.600 298.050 523.050 ;
        RECT 286.950 521.400 298.050 522.600 ;
        RECT 286.950 520.950 289.050 521.400 ;
        RECT 292.950 520.950 295.050 521.400 ;
        RECT 295.950 520.950 298.050 521.400 ;
        RECT 316.950 520.950 319.050 523.050 ;
        RECT 433.950 522.600 436.050 523.050 ;
        RECT 442.950 522.600 445.050 523.050 ;
        RECT 433.950 521.400 445.050 522.600 ;
        RECT 433.950 520.950 436.050 521.400 ;
        RECT 442.950 520.950 445.050 521.400 ;
        RECT 475.950 522.600 478.050 523.050 ;
        RECT 493.950 522.600 496.050 523.050 ;
        RECT 475.950 521.400 496.050 522.600 ;
        RECT 475.950 520.950 478.050 521.400 ;
        RECT 493.950 520.950 496.050 521.400 ;
        RECT 523.950 520.950 526.050 523.050 ;
        RECT 700.950 520.950 703.050 523.050 ;
        RECT 103.950 517.950 106.050 520.050 ;
        RECT 259.950 519.600 262.050 520.050 ;
        RECT 119.400 518.400 262.050 519.600 ;
        RECT 43.950 516.600 46.050 517.050 ;
        RECT 119.400 516.600 120.600 518.400 ;
        RECT 259.950 517.950 262.050 518.400 ;
        RECT 262.950 519.600 265.050 520.050 ;
        RECT 271.950 519.600 274.050 520.050 ;
        RECT 262.950 518.400 274.050 519.600 ;
        RECT 262.950 517.950 265.050 518.400 ;
        RECT 271.950 517.950 274.050 518.400 ;
        RECT 301.950 519.600 304.050 520.050 ;
        RECT 313.950 519.600 316.050 520.050 ;
        RECT 301.950 518.400 316.050 519.600 ;
        RECT 301.950 517.950 304.050 518.400 ;
        RECT 313.950 517.950 316.050 518.400 ;
        RECT 448.950 519.600 451.050 520.050 ;
        RECT 484.950 519.600 487.050 520.050 ;
        RECT 448.950 518.400 487.050 519.600 ;
        RECT 448.950 517.950 451.050 518.400 ;
        RECT 484.950 517.950 487.050 518.400 ;
        RECT 565.950 519.600 568.050 520.050 ;
        RECT 574.950 519.600 577.050 520.050 ;
        RECT 583.950 519.600 586.050 520.050 ;
        RECT 565.950 518.400 586.050 519.600 ;
        RECT 565.950 517.950 568.050 518.400 ;
        RECT 574.950 517.950 577.050 518.400 ;
        RECT 583.950 517.950 586.050 518.400 ;
        RECT 589.950 519.600 592.050 520.050 ;
        RECT 601.950 519.600 604.050 520.050 ;
        RECT 649.950 519.600 652.050 520.050 ;
        RECT 589.950 518.400 652.050 519.600 ;
        RECT 589.950 517.950 592.050 518.400 ;
        RECT 601.950 517.950 604.050 518.400 ;
        RECT 649.950 517.950 652.050 518.400 ;
        RECT 652.950 519.600 655.050 520.050 ;
        RECT 697.950 519.600 700.050 520.050 ;
        RECT 652.950 518.400 700.050 519.600 ;
        RECT 652.950 517.950 655.050 518.400 ;
        RECT 697.950 517.950 700.050 518.400 ;
        RECT 43.950 515.400 120.600 516.600 ;
        RECT 121.950 516.600 124.050 517.050 ;
        RECT 160.950 516.600 163.050 517.050 ;
        RECT 121.950 515.400 163.050 516.600 ;
        RECT 43.950 514.950 46.050 515.400 ;
        RECT 121.950 514.950 124.050 515.400 ;
        RECT 160.950 514.950 163.050 515.400 ;
        RECT 277.950 516.600 280.050 517.050 ;
        RECT 283.950 516.600 286.050 517.050 ;
        RECT 277.950 515.400 286.050 516.600 ;
        RECT 277.950 514.950 280.050 515.400 ;
        RECT 283.950 514.950 286.050 515.400 ;
        RECT 250.950 513.600 253.050 514.050 ;
        RECT 313.950 513.600 316.050 514.050 ;
        RECT 250.950 512.400 316.050 513.600 ;
        RECT 250.950 511.950 253.050 512.400 ;
        RECT 313.950 511.950 316.050 512.400 ;
        RECT 412.950 513.600 415.050 514.050 ;
        RECT 622.950 513.600 625.050 514.050 ;
        RECT 631.950 513.600 634.050 514.050 ;
        RECT 412.950 512.400 634.050 513.600 ;
        RECT 412.950 511.950 415.050 512.400 ;
        RECT 622.950 511.950 625.050 512.400 ;
        RECT 631.950 511.950 634.050 512.400 ;
        RECT 1.950 510.600 4.050 511.050 ;
        RECT 43.950 510.600 46.050 511.050 ;
        RECT 1.950 509.400 46.050 510.600 ;
        RECT 1.950 508.950 4.050 509.400 ;
        RECT 43.950 508.950 46.050 509.400 ;
        RECT 91.950 510.600 94.050 511.050 ;
        RECT 127.950 510.600 130.050 511.050 ;
        RECT 91.950 509.400 130.050 510.600 ;
        RECT 91.950 508.950 94.050 509.400 ;
        RECT 127.950 508.950 130.050 509.400 ;
        RECT 139.950 510.600 142.050 511.050 ;
        RECT 151.950 510.600 154.050 511.050 ;
        RECT 139.950 509.400 154.050 510.600 ;
        RECT 139.950 508.950 142.050 509.400 ;
        RECT 151.950 508.950 154.050 509.400 ;
        RECT 181.950 510.600 184.050 511.050 ;
        RECT 220.950 510.600 223.050 511.050 ;
        RECT 256.950 510.600 259.050 511.050 ;
        RECT 265.950 510.600 268.050 511.050 ;
        RECT 181.950 509.400 268.050 510.600 ;
        RECT 181.950 508.950 184.050 509.400 ;
        RECT 220.950 508.950 223.050 509.400 ;
        RECT 256.950 508.950 259.050 509.400 ;
        RECT 265.950 508.950 268.050 509.400 ;
        RECT 493.950 510.600 496.050 511.050 ;
        RECT 580.950 510.600 583.050 511.050 ;
        RECT 493.950 509.400 583.050 510.600 ;
        RECT 493.950 508.950 496.050 509.400 ;
        RECT 580.950 508.950 583.050 509.400 ;
        RECT 106.950 507.600 109.050 508.050 ;
        RECT 112.950 507.600 115.050 508.050 ;
        RECT 163.950 507.600 166.050 508.050 ;
        RECT 250.950 507.600 253.050 508.050 ;
        RECT 106.950 506.400 150.600 507.600 ;
        RECT 106.950 505.950 109.050 506.400 ;
        RECT 112.950 505.950 115.050 506.400 ;
        RECT 37.950 504.600 40.050 505.050 ;
        RECT 79.950 504.600 82.050 505.050 ;
        RECT 37.950 503.400 82.050 504.600 ;
        RECT 37.950 502.950 40.050 503.400 ;
        RECT 79.950 502.950 82.050 503.400 ;
        RECT 100.950 504.600 103.050 505.050 ;
        RECT 109.950 504.600 112.050 505.050 ;
        RECT 100.950 503.400 112.050 504.600 ;
        RECT 100.950 502.950 103.050 503.400 ;
        RECT 109.950 502.950 112.050 503.400 ;
        RECT 136.950 504.600 139.050 505.050 ;
        RECT 145.950 504.600 148.050 505.050 ;
        RECT 136.950 503.400 148.050 504.600 ;
        RECT 149.400 504.600 150.600 506.400 ;
        RECT 163.950 506.400 253.050 507.600 ;
        RECT 163.950 505.950 166.050 506.400 ;
        RECT 250.950 505.950 253.050 506.400 ;
        RECT 205.950 504.600 208.050 505.050 ;
        RECT 149.400 503.400 208.050 504.600 ;
        RECT 136.950 502.950 139.050 503.400 ;
        RECT 145.950 502.950 148.050 503.400 ;
        RECT 205.950 502.950 208.050 503.400 ;
        RECT 259.950 504.600 262.050 505.050 ;
        RECT 289.950 504.600 292.050 505.050 ;
        RECT 259.950 503.400 292.050 504.600 ;
        RECT 259.950 502.950 262.050 503.400 ;
        RECT 289.950 502.950 292.050 503.400 ;
        RECT 352.950 504.600 355.050 505.050 ;
        RECT 376.950 504.600 379.050 505.050 ;
        RECT 352.950 503.400 379.050 504.600 ;
        RECT 352.950 502.950 355.050 503.400 ;
        RECT 376.950 502.950 379.050 503.400 ;
        RECT 37.950 501.600 40.050 502.050 ;
        RECT 94.950 501.600 97.050 502.050 ;
        RECT 37.950 500.400 97.050 501.600 ;
        RECT 37.950 499.950 40.050 500.400 ;
        RECT 94.950 499.950 97.050 500.400 ;
        RECT 115.950 501.600 118.050 502.050 ;
        RECT 163.950 501.600 166.050 502.050 ;
        RECT 115.950 500.400 166.050 501.600 ;
        RECT 115.950 499.950 118.050 500.400 ;
        RECT 163.950 499.950 166.050 500.400 ;
        RECT 214.950 501.600 217.050 502.050 ;
        RECT 322.950 501.600 325.050 502.050 ;
        RECT 214.950 500.400 325.050 501.600 ;
        RECT 214.950 499.950 217.050 500.400 ;
        RECT 322.950 499.950 325.050 500.400 ;
        RECT 520.950 501.600 523.050 502.050 ;
        RECT 529.950 501.600 532.050 502.050 ;
        RECT 520.950 500.400 532.050 501.600 ;
        RECT 520.950 499.950 523.050 500.400 ;
        RECT 529.950 499.950 532.050 500.400 ;
        RECT 46.950 498.600 49.050 499.050 ;
        RECT 58.950 498.600 61.050 499.050 ;
        RECT 46.950 497.400 61.050 498.600 ;
        RECT 46.950 496.950 49.050 497.400 ;
        RECT 58.950 496.950 61.050 497.400 ;
        RECT 67.950 498.600 70.050 499.050 ;
        RECT 76.950 498.600 79.050 499.050 ;
        RECT 181.950 498.600 184.050 499.050 ;
        RECT 67.950 497.400 184.050 498.600 ;
        RECT 67.950 496.950 70.050 497.400 ;
        RECT 76.950 496.950 79.050 497.400 ;
        RECT 181.950 496.950 184.050 497.400 ;
        RECT 244.950 498.600 247.050 499.050 ;
        RECT 319.950 498.600 322.050 499.050 ;
        RECT 244.950 497.400 322.050 498.600 ;
        RECT 244.950 496.950 247.050 497.400 ;
        RECT 319.950 496.950 322.050 497.400 ;
        RECT 472.950 498.600 475.050 499.050 ;
        RECT 520.950 498.600 523.050 499.050 ;
        RECT 472.950 497.400 523.050 498.600 ;
        RECT 472.950 496.950 475.050 497.400 ;
        RECT 520.950 496.950 523.050 497.400 ;
        RECT 538.950 498.600 541.050 499.050 ;
        RECT 565.950 498.600 568.050 499.050 ;
        RECT 538.950 497.400 568.050 498.600 ;
        RECT 538.950 496.950 541.050 497.400 ;
        RECT 565.950 496.950 568.050 497.400 ;
        RECT 610.950 498.600 613.050 499.050 ;
        RECT 673.950 498.600 676.050 499.050 ;
        RECT 610.950 497.400 676.050 498.600 ;
        RECT 610.950 496.950 613.050 497.400 ;
        RECT 673.950 496.950 676.050 497.400 ;
        RECT 67.950 495.600 70.050 496.050 ;
        RECT 82.950 495.600 85.050 496.050 ;
        RECT 67.950 494.400 85.050 495.600 ;
        RECT 67.950 493.950 70.050 494.400 ;
        RECT 82.950 493.950 85.050 494.400 ;
        RECT 88.950 495.600 91.050 496.050 ;
        RECT 340.950 495.600 343.050 496.050 ;
        RECT 349.950 495.600 352.050 496.050 ;
        RECT 358.950 495.600 361.050 496.050 ;
        RECT 88.950 494.400 123.600 495.600 ;
        RECT 88.950 493.950 91.050 494.400 ;
        RECT 4.950 492.600 7.050 493.050 ;
        RECT 43.950 492.600 46.050 493.050 ;
        RECT 4.950 491.400 46.050 492.600 ;
        RECT 122.400 492.600 123.600 494.400 ;
        RECT 340.950 494.400 361.050 495.600 ;
        RECT 340.950 493.950 343.050 494.400 ;
        RECT 349.950 493.950 352.050 494.400 ;
        RECT 358.950 493.950 361.050 494.400 ;
        RECT 490.950 495.600 493.050 496.050 ;
        RECT 535.950 495.600 538.050 496.050 ;
        RECT 490.950 494.400 538.050 495.600 ;
        RECT 490.950 493.950 493.050 494.400 ;
        RECT 535.950 493.950 538.050 494.400 ;
        RECT 538.950 495.600 541.050 496.050 ;
        RECT 544.950 495.600 547.050 496.050 ;
        RECT 538.950 494.400 547.050 495.600 ;
        RECT 538.950 493.950 541.050 494.400 ;
        RECT 544.950 493.950 547.050 494.400 ;
        RECT 667.950 495.600 670.050 496.050 ;
        RECT 694.950 495.600 697.050 496.050 ;
        RECT 667.950 494.400 697.050 495.600 ;
        RECT 667.950 493.950 670.050 494.400 ;
        RECT 694.950 493.950 697.050 494.400 ;
        RECT 136.950 492.600 139.050 493.050 ;
        RECT 122.400 491.400 139.050 492.600 ;
        RECT 4.950 490.950 7.050 491.400 ;
        RECT 43.950 490.950 46.050 491.400 ;
        RECT 136.950 490.950 139.050 491.400 ;
        RECT 148.950 492.600 151.050 493.050 ;
        RECT 271.950 492.600 274.050 493.050 ;
        RECT 292.950 492.600 295.050 493.050 ;
        RECT 304.950 492.600 307.050 493.050 ;
        RECT 148.950 491.400 307.050 492.600 ;
        RECT 148.950 490.950 151.050 491.400 ;
        RECT 271.950 490.950 274.050 491.400 ;
        RECT 292.950 490.950 295.050 491.400 ;
        RECT 304.950 490.950 307.050 491.400 ;
        RECT 340.950 492.600 343.050 493.050 ;
        RECT 352.950 492.600 355.050 493.050 ;
        RECT 340.950 491.400 355.050 492.600 ;
        RECT 340.950 490.950 343.050 491.400 ;
        RECT 352.950 490.950 355.050 491.400 ;
        RECT 463.950 492.600 466.050 493.050 ;
        RECT 481.950 492.600 484.050 493.050 ;
        RECT 463.950 491.400 484.050 492.600 ;
        RECT 463.950 490.950 466.050 491.400 ;
        RECT 481.950 490.950 484.050 491.400 ;
        RECT 583.950 492.600 586.050 493.050 ;
        RECT 586.950 492.600 589.050 493.050 ;
        RECT 592.950 492.600 595.050 493.050 ;
        RECT 583.950 491.400 595.050 492.600 ;
        RECT 583.950 490.950 586.050 491.400 ;
        RECT 586.950 490.950 589.050 491.400 ;
        RECT 592.950 490.950 595.050 491.400 ;
        RECT 595.950 492.600 598.050 493.050 ;
        RECT 601.950 492.600 604.050 493.050 ;
        RECT 595.950 491.400 604.050 492.600 ;
        RECT 595.950 490.950 598.050 491.400 ;
        RECT 601.950 490.950 604.050 491.400 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 664.950 492.600 667.050 493.050 ;
        RECT 676.950 492.600 679.050 493.050 ;
        RECT 700.950 492.600 703.050 493.050 ;
        RECT 664.950 491.400 679.050 492.600 ;
        RECT 664.950 490.950 667.050 491.400 ;
        RECT 676.950 490.950 679.050 491.400 ;
        RECT 695.400 491.400 703.050 492.600 ;
        RECT 16.950 489.600 19.050 490.050 ;
        RECT 64.950 489.600 67.050 490.050 ;
        RECT 70.950 489.600 73.050 490.050 ;
        RECT 88.950 489.600 91.050 490.050 ;
        RECT 16.950 488.400 54.600 489.600 ;
        RECT 16.950 487.950 19.050 488.400 ;
        RECT 25.950 486.600 28.050 487.050 ;
        RECT 23.400 485.400 28.050 486.600 ;
        RECT 23.400 483.600 24.600 485.400 ;
        RECT 25.950 484.950 28.050 485.400 ;
        RECT 53.400 484.050 54.600 488.400 ;
        RECT 64.950 488.400 91.050 489.600 ;
        RECT 64.950 487.950 67.050 488.400 ;
        RECT 70.950 487.950 73.050 488.400 ;
        RECT 88.950 487.950 91.050 488.400 ;
        RECT 97.950 489.600 100.050 490.050 ;
        RECT 121.950 489.600 124.050 490.050 ;
        RECT 130.950 489.600 133.050 490.050 ;
        RECT 97.950 488.400 124.050 489.600 ;
        RECT 97.950 487.950 100.050 488.400 ;
        RECT 121.950 487.950 124.050 488.400 ;
        RECT 128.400 488.400 133.050 489.600 ;
        RECT 55.950 486.600 58.050 487.050 ;
        RECT 61.950 486.600 64.050 487.050 ;
        RECT 55.950 485.400 64.050 486.600 ;
        RECT 55.950 484.950 58.050 485.400 ;
        RECT 61.950 484.950 64.050 485.400 ;
        RECT 128.400 484.050 129.600 488.400 ;
        RECT 130.950 487.950 133.050 488.400 ;
        RECT 187.950 489.600 190.050 490.050 ;
        RECT 190.950 489.600 193.050 490.050 ;
        RECT 187.950 488.400 204.600 489.600 ;
        RECT 187.950 487.950 190.050 488.400 ;
        RECT 190.950 487.950 193.050 488.400 ;
        RECT 203.400 487.050 204.600 488.400 ;
        RECT 208.950 487.950 211.050 490.050 ;
        RECT 223.950 489.600 226.050 490.050 ;
        RECT 226.950 489.600 229.050 490.050 ;
        RECT 238.950 489.600 241.050 490.050 ;
        RECT 223.950 488.400 241.050 489.600 ;
        RECT 223.950 487.950 226.050 488.400 ;
        RECT 226.950 487.950 229.050 488.400 ;
        RECT 238.950 487.950 241.050 488.400 ;
        RECT 244.950 487.950 247.050 490.050 ;
        RECT 253.950 489.600 256.050 490.050 ;
        RECT 253.950 488.400 273.600 489.600 ;
        RECT 253.950 487.950 256.050 488.400 ;
        RECT 139.950 486.600 142.050 487.050 ;
        RECT 148.950 486.600 151.050 487.050 ;
        RECT 160.950 486.600 163.050 487.050 ;
        RECT 139.950 485.400 151.050 486.600 ;
        RECT 139.950 484.950 142.050 485.400 ;
        RECT 148.950 484.950 151.050 485.400 ;
        RECT 158.400 485.400 163.050 486.600 ;
        RECT 17.400 482.400 24.600 483.600 ;
        RECT 25.950 483.600 28.050 484.050 ;
        RECT 31.950 483.600 34.050 484.050 ;
        RECT 25.950 482.400 34.050 483.600 ;
        RECT 1.950 480.600 4.050 481.050 ;
        RECT 13.950 480.600 16.050 481.050 ;
        RECT 1.950 479.400 16.050 480.600 ;
        RECT 1.950 478.950 4.050 479.400 ;
        RECT 13.950 478.950 16.050 479.400 ;
        RECT 17.400 477.600 18.600 482.400 ;
        RECT 25.950 481.950 28.050 482.400 ;
        RECT 31.950 481.950 34.050 482.400 ;
        RECT 52.950 481.950 55.050 484.050 ;
        RECT 64.950 483.600 67.050 484.050 ;
        RECT 70.950 483.600 73.050 484.050 ;
        RECT 64.950 482.400 73.050 483.600 ;
        RECT 64.950 481.950 67.050 482.400 ;
        RECT 70.950 481.950 73.050 482.400 ;
        RECT 88.950 483.600 91.050 484.050 ;
        RECT 109.950 483.600 112.050 484.050 ;
        RECT 88.950 482.400 112.050 483.600 ;
        RECT 88.950 481.950 91.050 482.400 ;
        RECT 109.950 481.950 112.050 482.400 ;
        RECT 127.950 481.950 130.050 484.050 ;
        RECT 133.950 483.600 136.050 484.050 ;
        RECT 158.400 483.600 159.600 485.400 ;
        RECT 160.950 484.950 163.050 485.400 ;
        RECT 190.950 486.600 193.050 487.050 ;
        RECT 196.950 486.600 199.050 487.050 ;
        RECT 190.950 485.400 199.050 486.600 ;
        RECT 190.950 484.950 193.050 485.400 ;
        RECT 196.950 484.950 199.050 485.400 ;
        RECT 202.950 484.950 205.050 487.050 ;
        RECT 133.950 482.400 159.600 483.600 ;
        RECT 160.950 483.600 163.050 484.050 ;
        RECT 166.950 483.600 169.050 484.050 ;
        RECT 209.400 483.600 210.600 487.950 ;
        RECT 232.950 486.600 235.050 487.050 ;
        RECT 241.950 486.600 244.050 487.050 ;
        RECT 232.950 485.400 244.050 486.600 ;
        RECT 232.950 484.950 235.050 485.400 ;
        RECT 241.950 484.950 244.050 485.400 ;
        RECT 160.950 482.400 210.600 483.600 ;
        RECT 214.950 483.600 217.050 484.050 ;
        RECT 229.950 483.600 232.050 484.050 ;
        RECT 214.950 482.400 232.050 483.600 ;
        RECT 245.400 483.600 246.600 487.950 ;
        RECT 253.950 483.600 256.050 484.050 ;
        RECT 245.400 482.400 256.050 483.600 ;
        RECT 133.950 481.950 136.050 482.400 ;
        RECT 160.950 481.950 163.050 482.400 ;
        RECT 166.950 481.950 169.050 482.400 ;
        RECT 214.950 481.950 217.050 482.400 ;
        RECT 229.950 481.950 232.050 482.400 ;
        RECT 253.950 481.950 256.050 482.400 ;
        RECT 256.950 483.600 259.050 484.050 ;
        RECT 268.950 483.600 271.050 484.050 ;
        RECT 256.950 482.400 271.050 483.600 ;
        RECT 256.950 481.950 259.050 482.400 ;
        RECT 268.950 481.950 271.050 482.400 ;
        RECT 19.950 480.600 22.050 481.050 ;
        RECT 34.950 480.600 37.050 481.050 ;
        RECT 52.950 480.600 55.050 481.050 ;
        RECT 82.950 480.600 85.050 481.050 ;
        RECT 19.950 479.400 85.050 480.600 ;
        RECT 19.950 478.950 22.050 479.400 ;
        RECT 34.950 478.950 37.050 479.400 ;
        RECT 52.950 478.950 55.050 479.400 ;
        RECT 82.950 478.950 85.050 479.400 ;
        RECT 121.950 480.600 124.050 481.050 ;
        RECT 124.950 480.600 127.050 481.050 ;
        RECT 175.950 480.600 178.050 481.050 ;
        RECT 121.950 479.400 178.050 480.600 ;
        RECT 121.950 478.950 124.050 479.400 ;
        RECT 124.950 478.950 127.050 479.400 ;
        RECT 175.950 478.950 178.050 479.400 ;
        RECT 199.950 480.600 202.050 481.050 ;
        RECT 217.950 480.600 220.050 481.050 ;
        RECT 199.950 479.400 220.050 480.600 ;
        RECT 199.950 478.950 202.050 479.400 ;
        RECT 217.950 478.950 220.050 479.400 ;
        RECT 232.950 480.600 235.050 481.050 ;
        RECT 256.950 480.600 259.050 481.050 ;
        RECT 232.950 479.400 259.050 480.600 ;
        RECT 272.400 480.600 273.600 488.400 ;
        RECT 310.950 487.950 313.050 490.050 ;
        RECT 316.950 489.600 319.050 490.050 ;
        RECT 343.950 489.600 346.050 490.050 ;
        RECT 316.950 488.400 339.600 489.600 ;
        RECT 316.950 487.950 319.050 488.400 ;
        RECT 311.400 484.050 312.600 487.950 ;
        RECT 338.400 487.050 339.600 488.400 ;
        RECT 343.950 488.400 360.600 489.600 ;
        RECT 343.950 487.950 346.050 488.400 ;
        RECT 319.950 486.600 322.050 487.050 ;
        RECT 317.400 485.400 322.050 486.600 ;
        RECT 317.400 484.050 318.600 485.400 ;
        RECT 319.950 484.950 322.050 485.400 ;
        RECT 322.950 486.600 325.050 487.050 ;
        RECT 322.950 485.400 330.600 486.600 ;
        RECT 322.950 484.950 325.050 485.400 ;
        RECT 329.400 484.050 330.600 485.400 ;
        RECT 331.950 484.950 334.050 487.050 ;
        RECT 337.950 484.950 340.050 487.050 ;
        RECT 349.950 484.950 352.050 487.050 ;
        RECT 274.950 483.600 277.050 484.050 ;
        RECT 280.950 483.600 283.050 484.050 ;
        RECT 274.950 482.400 283.050 483.600 ;
        RECT 274.950 481.950 277.050 482.400 ;
        RECT 280.950 481.950 283.050 482.400 ;
        RECT 289.950 481.950 292.050 484.050 ;
        RECT 310.950 481.950 313.050 484.050 ;
        RECT 316.950 481.950 319.050 484.050 ;
        RECT 328.950 481.950 331.050 484.050 ;
        RECT 274.950 480.600 277.050 481.050 ;
        RECT 272.400 479.400 277.050 480.600 ;
        RECT 232.950 478.950 235.050 479.400 ;
        RECT 256.950 478.950 259.050 479.400 ;
        RECT 274.950 478.950 277.050 479.400 ;
        RECT 280.950 480.600 283.050 481.050 ;
        RECT 290.400 480.600 291.600 481.950 ;
        RECT 280.950 479.400 291.600 480.600 ;
        RECT 310.950 480.600 313.050 481.050 ;
        RECT 332.400 480.600 333.600 484.950 ;
        RECT 334.950 483.600 337.050 484.050 ;
        RECT 340.950 483.600 343.050 484.050 ;
        RECT 334.950 482.400 343.050 483.600 ;
        RECT 334.950 481.950 337.050 482.400 ;
        RECT 340.950 481.950 343.050 482.400 ;
        RECT 350.400 481.050 351.600 484.950 ;
        RECT 359.400 484.050 360.600 488.400 ;
        RECT 469.950 487.950 472.050 490.050 ;
        RECT 514.950 489.600 517.050 490.050 ;
        RECT 506.400 488.400 517.050 489.600 ;
        RECT 442.950 486.600 445.050 487.050 ;
        RECT 451.950 486.600 454.050 487.050 ;
        RECT 442.950 485.400 454.050 486.600 ;
        RECT 442.950 484.950 445.050 485.400 ;
        RECT 451.950 484.950 454.050 485.400 ;
        RECT 457.950 486.600 460.050 487.050 ;
        RECT 463.950 486.600 466.050 487.050 ;
        RECT 457.950 485.400 466.050 486.600 ;
        RECT 457.950 484.950 460.050 485.400 ;
        RECT 463.950 484.950 466.050 485.400 ;
        RECT 470.400 484.050 471.600 487.950 ;
        RECT 472.950 486.600 475.050 487.050 ;
        RECT 493.950 486.600 496.050 487.050 ;
        RECT 502.950 486.600 505.050 487.050 ;
        RECT 472.950 485.400 505.050 486.600 ;
        RECT 472.950 484.950 475.050 485.400 ;
        RECT 493.950 484.950 496.050 485.400 ;
        RECT 502.950 484.950 505.050 485.400 ;
        RECT 506.400 484.050 507.600 488.400 ;
        RECT 514.950 487.950 517.050 488.400 ;
        RECT 529.950 489.600 532.050 490.050 ;
        RECT 541.950 489.600 544.050 490.050 ;
        RECT 529.950 488.400 544.050 489.600 ;
        RECT 529.950 487.950 532.050 488.400 ;
        RECT 541.950 487.950 544.050 488.400 ;
        RECT 553.950 487.950 556.050 490.050 ;
        RECT 580.950 489.600 583.050 490.050 ;
        RECT 604.950 489.600 607.050 490.050 ;
        RECT 646.950 489.600 649.050 490.050 ;
        RECT 580.950 488.400 607.050 489.600 ;
        RECT 580.950 487.950 583.050 488.400 ;
        RECT 604.950 487.950 607.050 488.400 ;
        RECT 623.400 488.400 642.600 489.600 ;
        RECT 538.950 486.600 541.050 487.050 ;
        RECT 554.400 486.600 555.600 487.950 ;
        RECT 601.950 486.600 604.050 487.050 ;
        RECT 623.400 486.600 624.600 488.400 ;
        RECT 538.950 485.400 555.600 486.600 ;
        RECT 593.400 485.400 604.050 486.600 ;
        RECT 538.950 484.950 541.050 485.400 ;
        RECT 593.400 484.050 594.600 485.400 ;
        RECT 601.950 484.950 604.050 485.400 ;
        RECT 611.400 485.400 624.600 486.600 ;
        RECT 358.950 481.950 361.050 484.050 ;
        RECT 367.950 481.950 370.050 484.050 ;
        RECT 415.950 483.600 418.050 484.050 ;
        RECT 424.950 483.600 427.050 484.050 ;
        RECT 445.950 483.600 448.050 484.050 ;
        RECT 415.950 482.400 448.050 483.600 ;
        RECT 415.950 481.950 418.050 482.400 ;
        RECT 424.950 481.950 427.050 482.400 ;
        RECT 445.950 481.950 448.050 482.400 ;
        RECT 454.950 483.600 457.050 484.050 ;
        RECT 466.950 483.600 469.050 484.050 ;
        RECT 454.950 482.400 469.050 483.600 ;
        RECT 454.950 481.950 457.050 482.400 ;
        RECT 466.950 481.950 469.050 482.400 ;
        RECT 469.950 481.950 472.050 484.050 ;
        RECT 484.950 483.600 487.050 484.050 ;
        RECT 496.950 483.600 499.050 484.050 ;
        RECT 484.950 482.400 499.050 483.600 ;
        RECT 484.950 481.950 487.050 482.400 ;
        RECT 496.950 481.950 499.050 482.400 ;
        RECT 505.950 481.950 508.050 484.050 ;
        RECT 517.950 483.600 520.050 484.050 ;
        RECT 562.950 483.600 565.050 484.050 ;
        RECT 517.950 482.400 565.050 483.600 ;
        RECT 517.950 481.950 520.050 482.400 ;
        RECT 562.950 481.950 565.050 482.400 ;
        RECT 592.950 481.950 595.050 484.050 ;
        RECT 598.950 483.600 601.050 484.050 ;
        RECT 611.400 483.600 612.600 485.400 ;
        RECT 637.950 484.950 640.050 487.050 ;
        RECT 598.950 482.400 612.600 483.600 ;
        RECT 628.950 483.600 631.050 484.050 ;
        RECT 634.950 483.600 637.050 484.050 ;
        RECT 628.950 482.400 637.050 483.600 ;
        RECT 598.950 481.950 601.050 482.400 ;
        RECT 628.950 481.950 631.050 482.400 ;
        RECT 634.950 481.950 637.050 482.400 ;
        RECT 310.950 479.400 333.600 480.600 ;
        RECT 280.950 478.950 283.050 479.400 ;
        RECT 310.950 478.950 313.050 479.400 ;
        RECT 349.950 478.950 352.050 481.050 ;
        RECT 368.400 478.050 369.600 481.950 ;
        RECT 638.400 481.050 639.600 484.950 ;
        RECT 641.400 484.050 642.600 488.400 ;
        RECT 644.400 488.400 649.050 489.600 ;
        RECT 640.950 481.950 643.050 484.050 ;
        RECT 382.950 480.600 385.050 481.050 ;
        RECT 427.950 480.600 430.050 481.050 ;
        RECT 382.950 479.400 430.050 480.600 ;
        RECT 382.950 478.950 385.050 479.400 ;
        RECT 427.950 478.950 430.050 479.400 ;
        RECT 454.950 480.600 457.050 481.050 ;
        RECT 463.950 480.600 466.050 481.050 ;
        RECT 454.950 479.400 466.050 480.600 ;
        RECT 454.950 478.950 457.050 479.400 ;
        RECT 463.950 478.950 466.050 479.400 ;
        RECT 475.950 480.600 478.050 481.050 ;
        RECT 490.950 480.600 493.050 481.050 ;
        RECT 475.950 479.400 493.050 480.600 ;
        RECT 475.950 478.950 478.050 479.400 ;
        RECT 490.950 478.950 493.050 479.400 ;
        RECT 508.950 480.600 511.050 481.050 ;
        RECT 520.950 480.600 523.050 481.050 ;
        RECT 508.950 479.400 523.050 480.600 ;
        RECT 508.950 478.950 511.050 479.400 ;
        RECT 520.950 478.950 523.050 479.400 ;
        RECT 601.950 480.600 604.050 481.050 ;
        RECT 616.950 480.600 619.050 481.050 ;
        RECT 601.950 479.400 619.050 480.600 ;
        RECT 601.950 478.950 604.050 479.400 ;
        RECT 616.950 478.950 619.050 479.400 ;
        RECT 637.950 478.950 640.050 481.050 ;
        RECT 640.950 480.600 643.050 481.050 ;
        RECT 644.400 480.600 645.600 488.400 ;
        RECT 646.950 487.950 649.050 488.400 ;
        RECT 649.950 489.600 652.050 490.050 ;
        RECT 662.400 489.600 663.600 490.950 ;
        RECT 670.950 489.600 673.050 490.050 ;
        RECT 649.950 488.400 660.600 489.600 ;
        RECT 662.400 488.400 673.050 489.600 ;
        RECT 649.950 487.950 652.050 488.400 ;
        RECT 655.950 484.950 658.050 487.050 ;
        RECT 640.950 479.400 645.600 480.600 ;
        RECT 649.950 480.600 652.050 481.050 ;
        RECT 656.400 480.600 657.600 484.950 ;
        RECT 659.400 483.600 660.600 488.400 ;
        RECT 670.950 487.950 673.050 488.400 ;
        RECT 661.950 486.600 664.050 487.050 ;
        RECT 673.950 486.600 676.050 487.050 ;
        RECT 661.950 485.400 676.050 486.600 ;
        RECT 661.950 484.950 664.050 485.400 ;
        RECT 673.950 484.950 676.050 485.400 ;
        RECT 661.950 483.600 664.050 484.050 ;
        RECT 659.400 482.400 664.050 483.600 ;
        RECT 661.950 481.950 664.050 482.400 ;
        RECT 649.950 479.400 657.600 480.600 ;
        RECT 640.950 478.950 643.050 479.400 ;
        RECT 649.950 478.950 652.050 479.400 ;
        RECT 19.950 477.600 22.050 478.050 ;
        RECT 17.400 476.400 22.050 477.600 ;
        RECT 19.950 475.950 22.050 476.400 ;
        RECT 22.950 477.600 25.050 478.050 ;
        RECT 46.950 477.600 49.050 478.050 ;
        RECT 22.950 476.400 49.050 477.600 ;
        RECT 22.950 475.950 25.050 476.400 ;
        RECT 46.950 475.950 49.050 476.400 ;
        RECT 49.950 477.600 52.050 478.050 ;
        RECT 55.950 477.600 58.050 478.050 ;
        RECT 49.950 476.400 58.050 477.600 ;
        RECT 49.950 475.950 52.050 476.400 ;
        RECT 55.950 475.950 58.050 476.400 ;
        RECT 67.950 477.600 70.050 478.050 ;
        RECT 88.950 477.600 91.050 478.050 ;
        RECT 67.950 476.400 91.050 477.600 ;
        RECT 67.950 475.950 70.050 476.400 ;
        RECT 88.950 475.950 91.050 476.400 ;
        RECT 97.950 477.600 100.050 478.050 ;
        RECT 115.950 477.600 118.050 478.050 ;
        RECT 97.950 476.400 118.050 477.600 ;
        RECT 97.950 475.950 100.050 476.400 ;
        RECT 115.950 475.950 118.050 476.400 ;
        RECT 130.950 477.600 133.050 478.050 ;
        RECT 223.950 477.600 226.050 478.050 ;
        RECT 130.950 476.400 226.050 477.600 ;
        RECT 130.950 475.950 133.050 476.400 ;
        RECT 223.950 475.950 226.050 476.400 ;
        RECT 226.950 477.600 229.050 478.050 ;
        RECT 298.950 477.600 301.050 478.050 ;
        RECT 226.950 476.400 301.050 477.600 ;
        RECT 226.950 475.950 229.050 476.400 ;
        RECT 298.950 475.950 301.050 476.400 ;
        RECT 367.950 475.950 370.050 478.050 ;
        RECT 406.950 477.600 409.050 478.050 ;
        RECT 460.950 477.600 463.050 478.050 ;
        RECT 406.950 476.400 463.050 477.600 ;
        RECT 406.950 475.950 409.050 476.400 ;
        RECT 460.950 475.950 463.050 476.400 ;
        RECT 595.950 477.600 598.050 478.050 ;
        RECT 625.950 477.600 628.050 478.050 ;
        RECT 652.950 477.600 655.050 478.050 ;
        RECT 664.950 477.600 667.050 478.050 ;
        RECT 595.950 476.400 667.050 477.600 ;
        RECT 695.400 477.600 696.600 491.400 ;
        RECT 700.950 490.950 703.050 491.400 ;
        RECT 697.950 487.950 700.050 490.050 ;
        RECT 698.400 481.050 699.600 487.950 ;
        RECT 700.950 486.600 703.050 487.050 ;
        RECT 709.950 486.600 712.050 487.050 ;
        RECT 700.950 485.400 712.050 486.600 ;
        RECT 700.950 484.950 703.050 485.400 ;
        RECT 709.950 484.950 712.050 485.400 ;
        RECT 703.950 483.600 706.050 484.050 ;
        RECT 709.950 483.600 712.050 484.050 ;
        RECT 703.950 482.400 712.050 483.600 ;
        RECT 703.950 481.950 706.050 482.400 ;
        RECT 709.950 481.950 712.050 482.400 ;
        RECT 697.950 478.950 700.050 481.050 ;
        RECT 709.950 477.600 712.050 478.050 ;
        RECT 695.400 476.400 712.050 477.600 ;
        RECT 595.950 475.950 598.050 476.400 ;
        RECT 625.950 475.950 628.050 476.400 ;
        RECT 652.950 475.950 655.050 476.400 ;
        RECT 664.950 475.950 667.050 476.400 ;
        RECT 709.950 475.950 712.050 476.400 ;
        RECT 13.950 474.600 16.050 475.050 ;
        RECT 58.950 474.600 61.050 475.050 ;
        RECT 13.950 473.400 61.050 474.600 ;
        RECT 13.950 472.950 16.050 473.400 ;
        RECT 58.950 472.950 61.050 473.400 ;
        RECT 67.950 474.600 70.050 475.050 ;
        RECT 85.950 474.600 88.050 475.050 ;
        RECT 67.950 473.400 88.050 474.600 ;
        RECT 67.950 472.950 70.050 473.400 ;
        RECT 85.950 472.950 88.050 473.400 ;
        RECT 91.950 474.600 94.050 475.050 ;
        RECT 97.950 474.600 100.050 475.050 ;
        RECT 91.950 473.400 100.050 474.600 ;
        RECT 91.950 472.950 94.050 473.400 ;
        RECT 97.950 472.950 100.050 473.400 ;
        RECT 112.950 474.600 115.050 475.050 ;
        RECT 130.950 474.600 133.050 475.050 ;
        RECT 112.950 473.400 133.050 474.600 ;
        RECT 112.950 472.950 115.050 473.400 ;
        RECT 130.950 472.950 133.050 473.400 ;
        RECT 139.950 474.600 142.050 475.050 ;
        RECT 145.950 474.600 148.050 475.050 ;
        RECT 139.950 473.400 148.050 474.600 ;
        RECT 139.950 472.950 142.050 473.400 ;
        RECT 145.950 472.950 148.050 473.400 ;
        RECT 169.950 474.600 172.050 475.050 ;
        RECT 181.950 474.600 184.050 475.050 ;
        RECT 169.950 473.400 184.050 474.600 ;
        RECT 169.950 472.950 172.050 473.400 ;
        RECT 181.950 472.950 184.050 473.400 ;
        RECT 184.950 474.600 187.050 475.050 ;
        RECT 211.950 474.600 214.050 475.050 ;
        RECT 184.950 473.400 214.050 474.600 ;
        RECT 184.950 472.950 187.050 473.400 ;
        RECT 211.950 472.950 214.050 473.400 ;
        RECT 220.950 474.600 223.050 475.050 ;
        RECT 241.950 474.600 244.050 475.050 ;
        RECT 220.950 473.400 244.050 474.600 ;
        RECT 220.950 472.950 223.050 473.400 ;
        RECT 241.950 472.950 244.050 473.400 ;
        RECT 253.950 474.600 256.050 475.050 ;
        RECT 265.950 474.600 268.050 475.050 ;
        RECT 253.950 473.400 268.050 474.600 ;
        RECT 253.950 472.950 256.050 473.400 ;
        RECT 265.950 472.950 268.050 473.400 ;
        RECT 268.950 474.600 271.050 475.050 ;
        RECT 400.950 474.600 403.050 475.050 ;
        RECT 415.950 474.600 418.050 475.050 ;
        RECT 268.950 473.400 399.600 474.600 ;
        RECT 268.950 472.950 271.050 473.400 ;
        RECT 19.950 471.600 22.050 472.050 ;
        RECT 43.950 471.600 46.050 472.050 ;
        RECT 19.950 470.400 46.050 471.600 ;
        RECT 19.950 469.950 22.050 470.400 ;
        RECT 43.950 469.950 46.050 470.400 ;
        RECT 94.950 471.600 97.050 472.050 ;
        RECT 100.950 471.600 103.050 472.050 ;
        RECT 94.950 470.400 103.050 471.600 ;
        RECT 94.950 469.950 97.050 470.400 ;
        RECT 100.950 469.950 103.050 470.400 ;
        RECT 166.950 471.600 169.050 472.050 ;
        RECT 208.950 471.600 211.050 472.050 ;
        RECT 166.950 470.400 211.050 471.600 ;
        RECT 166.950 469.950 169.050 470.400 ;
        RECT 208.950 469.950 211.050 470.400 ;
        RECT 259.950 471.600 262.050 472.050 ;
        RECT 271.950 471.600 274.050 472.050 ;
        RECT 259.950 470.400 274.050 471.600 ;
        RECT 259.950 469.950 262.050 470.400 ;
        RECT 271.950 469.950 274.050 470.400 ;
        RECT 286.950 471.600 289.050 472.050 ;
        RECT 295.950 471.600 298.050 472.050 ;
        RECT 286.950 470.400 298.050 471.600 ;
        RECT 286.950 469.950 289.050 470.400 ;
        RECT 295.950 469.950 298.050 470.400 ;
        RECT 355.950 471.600 358.050 472.050 ;
        RECT 394.950 471.600 397.050 472.050 ;
        RECT 355.950 470.400 397.050 471.600 ;
        RECT 398.400 471.600 399.600 473.400 ;
        RECT 400.950 473.400 418.050 474.600 ;
        RECT 400.950 472.950 403.050 473.400 ;
        RECT 415.950 472.950 418.050 473.400 ;
        RECT 433.950 474.600 436.050 475.050 ;
        RECT 499.950 474.600 502.050 475.050 ;
        RECT 571.950 474.600 574.050 475.050 ;
        RECT 433.950 473.400 502.050 474.600 ;
        RECT 433.950 472.950 436.050 473.400 ;
        RECT 499.950 472.950 502.050 473.400 ;
        RECT 503.400 473.400 574.050 474.600 ;
        RECT 503.400 471.600 504.600 473.400 ;
        RECT 571.950 472.950 574.050 473.400 ;
        RECT 574.950 474.600 577.050 475.050 ;
        RECT 601.950 474.600 604.050 475.050 ;
        RECT 574.950 473.400 604.050 474.600 ;
        RECT 574.950 472.950 577.050 473.400 ;
        RECT 601.950 472.950 604.050 473.400 ;
        RECT 607.950 474.600 610.050 475.050 ;
        RECT 631.950 474.600 634.050 475.050 ;
        RECT 607.950 473.400 634.050 474.600 ;
        RECT 607.950 472.950 610.050 473.400 ;
        RECT 631.950 472.950 634.050 473.400 ;
        RECT 637.950 474.600 640.050 475.050 ;
        RECT 658.950 474.600 661.050 475.050 ;
        RECT 637.950 473.400 661.050 474.600 ;
        RECT 637.950 472.950 640.050 473.400 ;
        RECT 658.950 472.950 661.050 473.400 ;
        RECT 398.400 470.400 504.600 471.600 ;
        RECT 535.950 471.600 538.050 472.050 ;
        RECT 544.950 471.600 547.050 472.050 ;
        RECT 535.950 470.400 547.050 471.600 ;
        RECT 355.950 469.950 358.050 470.400 ;
        RECT 394.950 469.950 397.050 470.400 ;
        RECT 535.950 469.950 538.050 470.400 ;
        RECT 544.950 469.950 547.050 470.400 ;
        RECT 586.950 471.600 589.050 472.050 ;
        RECT 598.950 471.600 601.050 472.050 ;
        RECT 637.950 471.600 640.050 472.050 ;
        RECT 586.950 470.400 640.050 471.600 ;
        RECT 586.950 469.950 589.050 470.400 ;
        RECT 598.950 469.950 601.050 470.400 ;
        RECT 637.950 469.950 640.050 470.400 ;
        RECT 643.950 471.600 646.050 472.050 ;
        RECT 655.950 471.600 658.050 472.050 ;
        RECT 643.950 470.400 658.050 471.600 ;
        RECT 643.950 469.950 646.050 470.400 ;
        RECT 655.950 469.950 658.050 470.400 ;
        RECT 34.950 468.600 37.050 469.050 ;
        RECT 40.950 468.600 43.050 469.050 ;
        RECT 64.950 468.600 67.050 469.050 ;
        RECT 34.950 467.400 67.050 468.600 ;
        RECT 34.950 466.950 37.050 467.400 ;
        RECT 40.950 466.950 43.050 467.400 ;
        RECT 64.950 466.950 67.050 467.400 ;
        RECT 136.950 468.600 139.050 469.050 ;
        RECT 181.950 468.600 184.050 469.050 ;
        RECT 136.950 467.400 184.050 468.600 ;
        RECT 136.950 466.950 139.050 467.400 ;
        RECT 181.950 466.950 184.050 467.400 ;
        RECT 259.950 468.600 262.050 469.050 ;
        RECT 292.950 468.600 295.050 469.050 ;
        RECT 259.950 467.400 295.050 468.600 ;
        RECT 259.950 466.950 262.050 467.400 ;
        RECT 292.950 466.950 295.050 467.400 ;
        RECT 322.950 468.600 325.050 469.050 ;
        RECT 376.950 468.600 379.050 469.050 ;
        RECT 322.950 467.400 379.050 468.600 ;
        RECT 322.950 466.950 325.050 467.400 ;
        RECT 376.950 466.950 379.050 467.400 ;
        RECT 445.950 468.600 448.050 469.050 ;
        RECT 487.950 468.600 490.050 469.050 ;
        RECT 445.950 467.400 490.050 468.600 ;
        RECT 445.950 466.950 448.050 467.400 ;
        RECT 487.950 466.950 490.050 467.400 ;
        RECT 577.950 468.600 580.050 469.050 ;
        RECT 598.950 468.600 601.050 469.050 ;
        RECT 577.950 467.400 601.050 468.600 ;
        RECT 577.950 466.950 580.050 467.400 ;
        RECT 598.950 466.950 601.050 467.400 ;
        RECT 601.950 468.600 604.050 469.050 ;
        RECT 610.950 468.600 613.050 469.050 ;
        RECT 601.950 467.400 613.050 468.600 ;
        RECT 601.950 466.950 604.050 467.400 ;
        RECT 610.950 466.950 613.050 467.400 ;
        RECT 634.950 468.600 637.050 469.050 ;
        RECT 643.950 468.600 646.050 469.050 ;
        RECT 634.950 467.400 646.050 468.600 ;
        RECT 634.950 466.950 637.050 467.400 ;
        RECT 643.950 466.950 646.050 467.400 ;
        RECT 652.950 468.600 655.050 469.050 ;
        RECT 658.950 468.600 661.050 469.050 ;
        RECT 652.950 467.400 661.050 468.600 ;
        RECT 652.950 466.950 655.050 467.400 ;
        RECT 658.950 466.950 661.050 467.400 ;
        RECT 70.950 465.600 73.050 466.050 ;
        RECT 82.950 465.600 85.050 466.050 ;
        RECT 70.950 464.400 85.050 465.600 ;
        RECT 70.950 463.950 73.050 464.400 ;
        RECT 82.950 463.950 85.050 464.400 ;
        RECT 85.950 465.600 88.050 466.050 ;
        RECT 88.950 465.600 91.050 466.050 ;
        RECT 118.950 465.600 121.050 466.050 ;
        RECT 148.950 465.600 151.050 466.050 ;
        RECT 160.950 465.600 163.050 466.050 ;
        RECT 85.950 464.400 117.600 465.600 ;
        RECT 85.950 463.950 88.050 464.400 ;
        RECT 88.950 463.950 91.050 464.400 ;
        RECT 37.950 462.600 40.050 463.050 ;
        RECT 11.400 461.400 40.050 462.600 ;
        RECT 4.950 454.950 7.050 457.050 ;
        RECT 5.400 451.050 6.600 454.950 ;
        RECT 11.400 451.050 12.600 461.400 ;
        RECT 37.950 460.950 40.050 461.400 ;
        RECT 76.950 462.600 79.050 463.050 ;
        RECT 88.950 462.600 91.050 463.050 ;
        RECT 76.950 461.400 91.050 462.600 ;
        RECT 116.400 462.600 117.600 464.400 ;
        RECT 118.950 464.400 151.050 465.600 ;
        RECT 118.950 463.950 121.050 464.400 ;
        RECT 148.950 463.950 151.050 464.400 ;
        RECT 152.400 464.400 163.050 465.600 ;
        RECT 152.400 462.600 153.600 464.400 ;
        RECT 160.950 463.950 163.050 464.400 ;
        RECT 175.950 465.600 178.050 466.050 ;
        RECT 223.950 465.600 226.050 466.050 ;
        RECT 247.950 465.600 250.050 466.050 ;
        RECT 262.950 465.600 265.050 466.050 ;
        RECT 277.950 465.600 280.050 466.050 ;
        RECT 175.950 464.400 198.600 465.600 ;
        RECT 175.950 463.950 178.050 464.400 ;
        RECT 116.400 461.400 153.600 462.600 ;
        RECT 154.950 462.600 157.050 463.050 ;
        RECT 178.950 462.600 181.050 463.050 ;
        RECT 154.950 461.400 181.050 462.600 ;
        RECT 76.950 460.950 79.050 461.400 ;
        RECT 88.950 460.950 91.050 461.400 ;
        RECT 154.950 460.950 157.050 461.400 ;
        RECT 178.950 460.950 181.050 461.400 ;
        RECT 187.950 462.600 190.050 463.050 ;
        RECT 193.950 462.600 196.050 463.050 ;
        RECT 187.950 461.400 196.050 462.600 ;
        RECT 197.400 462.600 198.600 464.400 ;
        RECT 223.950 464.400 280.050 465.600 ;
        RECT 223.950 463.950 226.050 464.400 ;
        RECT 247.950 463.950 250.050 464.400 ;
        RECT 262.950 463.950 265.050 464.400 ;
        RECT 277.950 463.950 280.050 464.400 ;
        RECT 280.950 465.600 283.050 466.050 ;
        RECT 304.950 465.600 307.050 466.050 ;
        RECT 325.950 465.600 328.050 466.050 ;
        RECT 280.950 464.400 328.050 465.600 ;
        RECT 280.950 463.950 283.050 464.400 ;
        RECT 304.950 463.950 307.050 464.400 ;
        RECT 325.950 463.950 328.050 464.400 ;
        RECT 352.950 465.600 355.050 466.050 ;
        RECT 406.950 465.600 409.050 466.050 ;
        RECT 352.950 464.400 409.050 465.600 ;
        RECT 352.950 463.950 355.050 464.400 ;
        RECT 406.950 463.950 409.050 464.400 ;
        RECT 427.950 465.600 430.050 466.050 ;
        RECT 430.950 465.600 433.050 466.050 ;
        RECT 433.950 465.600 436.050 466.050 ;
        RECT 427.950 464.400 436.050 465.600 ;
        RECT 427.950 463.950 430.050 464.400 ;
        RECT 430.950 463.950 433.050 464.400 ;
        RECT 433.950 463.950 436.050 464.400 ;
        RECT 508.950 465.600 511.050 466.050 ;
        RECT 544.950 465.600 547.050 466.050 ;
        RECT 508.950 464.400 547.050 465.600 ;
        RECT 508.950 463.950 511.050 464.400 ;
        RECT 544.950 463.950 547.050 464.400 ;
        RECT 556.950 465.600 559.050 466.050 ;
        RECT 616.950 465.600 619.050 466.050 ;
        RECT 556.950 464.400 619.050 465.600 ;
        RECT 556.950 463.950 559.050 464.400 ;
        RECT 616.950 463.950 619.050 464.400 ;
        RECT 697.950 465.600 700.050 466.050 ;
        RECT 697.950 464.400 720.600 465.600 ;
        RECT 697.950 463.950 700.050 464.400 ;
        RECT 220.950 462.600 223.050 463.050 ;
        RECT 197.400 461.400 223.050 462.600 ;
        RECT 187.950 460.950 190.050 461.400 ;
        RECT 193.950 460.950 196.050 461.400 ;
        RECT 220.950 460.950 223.050 461.400 ;
        RECT 226.950 462.600 229.050 463.050 ;
        RECT 256.950 462.600 259.050 463.050 ;
        RECT 313.950 462.600 316.050 463.050 ;
        RECT 319.950 462.600 322.050 463.050 ;
        RECT 226.950 461.400 322.050 462.600 ;
        RECT 226.950 460.950 229.050 461.400 ;
        RECT 256.950 460.950 259.050 461.400 ;
        RECT 313.950 460.950 316.050 461.400 ;
        RECT 319.950 460.950 322.050 461.400 ;
        RECT 340.950 462.600 343.050 463.050 ;
        RECT 367.950 462.600 370.050 463.050 ;
        RECT 340.950 461.400 370.050 462.600 ;
        RECT 340.950 460.950 343.050 461.400 ;
        RECT 367.950 460.950 370.050 461.400 ;
        RECT 427.950 462.600 430.050 463.050 ;
        RECT 466.950 462.600 469.050 463.050 ;
        RECT 427.950 461.400 469.050 462.600 ;
        RECT 427.950 460.950 430.050 461.400 ;
        RECT 466.950 460.950 469.050 461.400 ;
        RECT 472.950 462.600 475.050 463.050 ;
        RECT 505.950 462.600 508.050 463.050 ;
        RECT 472.950 461.400 508.050 462.600 ;
        RECT 472.950 460.950 475.050 461.400 ;
        RECT 505.950 460.950 508.050 461.400 ;
        RECT 523.950 462.600 526.050 463.050 ;
        RECT 556.950 462.600 559.050 463.050 ;
        RECT 523.950 461.400 559.050 462.600 ;
        RECT 523.950 460.950 526.050 461.400 ;
        RECT 556.950 460.950 559.050 461.400 ;
        RECT 565.950 462.600 568.050 463.050 ;
        RECT 595.950 462.600 598.050 463.050 ;
        RECT 601.950 462.600 604.050 463.050 ;
        RECT 565.950 461.400 588.600 462.600 ;
        RECT 565.950 460.950 568.050 461.400 ;
        RECT 22.950 459.600 25.050 460.050 ;
        RECT 79.950 459.600 82.050 460.050 ;
        RECT 14.400 458.400 25.050 459.600 ;
        RECT 14.400 454.050 15.600 458.400 ;
        RECT 22.950 457.950 25.050 458.400 ;
        RECT 53.400 458.400 82.050 459.600 ;
        RECT 16.950 454.950 19.050 457.050 ;
        RECT 13.950 451.950 16.050 454.050 ;
        RECT 4.950 448.950 7.050 451.050 ;
        RECT 10.950 448.950 13.050 451.050 ;
        RECT 17.400 450.600 18.600 454.950 ;
        RECT 43.950 453.600 46.050 454.050 ;
        RECT 41.400 452.400 46.050 453.600 ;
        RECT 31.950 450.600 34.050 451.050 ;
        RECT 17.400 449.400 34.050 450.600 ;
        RECT 31.950 448.950 34.050 449.400 ;
        RECT 7.950 447.600 10.050 448.050 ;
        RECT 13.950 447.600 16.050 448.050 ;
        RECT 7.950 446.400 16.050 447.600 ;
        RECT 41.400 447.600 42.600 452.400 ;
        RECT 43.950 451.950 46.050 452.400 ;
        RECT 43.950 450.600 46.050 451.050 ;
        RECT 53.400 450.600 54.600 458.400 ;
        RECT 79.950 457.950 82.050 458.400 ;
        RECT 124.950 459.600 127.050 460.050 ;
        RECT 151.950 459.600 154.050 460.050 ;
        RECT 124.950 458.400 154.050 459.600 ;
        RECT 124.950 457.950 127.050 458.400 ;
        RECT 151.950 457.950 154.050 458.400 ;
        RECT 172.950 457.950 175.050 460.050 ;
        RECT 175.950 459.600 178.050 460.050 ;
        RECT 175.950 458.400 267.600 459.600 ;
        RECT 175.950 457.950 178.050 458.400 ;
        RECT 55.950 456.600 58.050 457.050 ;
        RECT 76.950 456.600 79.050 457.050 ;
        RECT 55.950 455.400 79.050 456.600 ;
        RECT 55.950 454.950 58.050 455.400 ;
        RECT 76.950 454.950 79.050 455.400 ;
        RECT 88.950 456.600 91.050 457.050 ;
        RECT 112.950 456.600 115.050 457.050 ;
        RECT 124.950 456.600 127.050 457.050 ;
        RECT 88.950 455.400 108.600 456.600 ;
        RECT 88.950 454.950 91.050 455.400 ;
        RECT 79.950 453.600 82.050 454.050 ;
        RECT 88.950 453.600 91.050 454.050 ;
        RECT 79.950 452.400 91.050 453.600 ;
        RECT 79.950 451.950 82.050 452.400 ;
        RECT 88.950 451.950 91.050 452.400 ;
        RECT 103.950 451.950 106.050 454.050 ;
        RECT 43.950 449.400 54.600 450.600 ;
        RECT 43.950 448.950 46.050 449.400 ;
        RECT 70.950 447.600 73.050 448.050 ;
        RECT 41.400 446.400 73.050 447.600 ;
        RECT 7.950 445.950 10.050 446.400 ;
        RECT 13.950 445.950 16.050 446.400 ;
        RECT 70.950 445.950 73.050 446.400 ;
        RECT 100.950 447.600 103.050 448.050 ;
        RECT 104.400 447.600 105.600 451.950 ;
        RECT 107.400 451.050 108.600 455.400 ;
        RECT 112.950 455.400 127.050 456.600 ;
        RECT 112.950 454.950 115.050 455.400 ;
        RECT 124.950 454.950 127.050 455.400 ;
        RECT 127.950 454.950 130.050 457.050 ;
        RECT 145.950 454.950 148.050 457.050 ;
        RECT 173.400 456.600 174.600 457.950 ;
        RECT 173.400 455.400 183.600 456.600 ;
        RECT 128.400 453.600 129.600 454.950 ;
        RECT 122.400 452.400 129.600 453.600 ;
        RECT 146.400 453.600 147.600 454.950 ;
        RECT 175.950 453.600 178.050 454.050 ;
        RECT 146.400 452.400 178.050 453.600 ;
        RECT 122.400 451.050 123.600 452.400 ;
        RECT 175.950 451.950 178.050 452.400 ;
        RECT 106.950 448.950 109.050 451.050 ;
        RECT 121.950 448.950 124.050 451.050 ;
        RECT 139.950 450.600 142.050 451.050 ;
        RECT 148.950 450.600 151.050 451.050 ;
        RECT 139.950 449.400 151.050 450.600 ;
        RECT 182.400 450.600 183.600 455.400 ;
        RECT 190.950 454.950 193.050 457.050 ;
        RECT 235.950 456.600 238.050 457.050 ;
        RECT 230.400 455.400 238.050 456.600 ;
        RECT 184.950 453.600 187.050 454.050 ;
        RECT 191.400 453.600 192.600 454.950 ;
        RECT 226.950 453.600 229.050 454.050 ;
        RECT 184.950 452.400 229.050 453.600 ;
        RECT 184.950 451.950 187.050 452.400 ;
        RECT 226.950 451.950 229.050 452.400 ;
        RECT 187.950 450.600 190.050 451.050 ;
        RECT 182.400 449.400 190.050 450.600 ;
        RECT 139.950 448.950 142.050 449.400 ;
        RECT 148.950 448.950 151.050 449.400 ;
        RECT 187.950 448.950 190.050 449.400 ;
        RECT 190.950 450.600 193.050 451.050 ;
        RECT 211.950 450.600 214.050 451.050 ;
        RECT 220.950 450.600 223.050 451.050 ;
        RECT 190.950 449.400 223.050 450.600 ;
        RECT 230.400 450.600 231.600 455.400 ;
        RECT 235.950 454.950 238.050 455.400 ;
        RECT 241.950 456.600 244.050 457.050 ;
        RECT 262.950 456.600 265.050 457.050 ;
        RECT 241.950 455.400 265.050 456.600 ;
        RECT 241.950 454.950 244.050 455.400 ;
        RECT 262.950 454.950 265.050 455.400 ;
        RECT 266.400 454.050 267.600 458.400 ;
        RECT 289.950 457.950 292.050 460.050 ;
        RECT 316.950 459.600 319.050 460.050 ;
        RECT 316.950 458.400 357.600 459.600 ;
        RECT 316.950 457.950 319.050 458.400 ;
        RECT 283.950 456.600 286.050 457.050 ;
        RECT 269.400 455.400 286.050 456.600 ;
        RECT 232.950 453.600 235.050 454.050 ;
        RECT 232.950 452.400 255.600 453.600 ;
        RECT 232.950 451.950 235.050 452.400 ;
        RECT 254.400 451.050 255.600 452.400 ;
        RECT 265.950 451.950 268.050 454.050 ;
        RECT 269.400 451.050 270.600 455.400 ;
        RECT 283.950 454.950 286.050 455.400 ;
        RECT 271.950 451.950 274.050 454.050 ;
        RECT 280.950 453.600 283.050 454.050 ;
        RECT 290.400 453.600 291.600 457.950 ;
        RECT 319.950 456.600 322.050 457.050 ;
        RECT 328.950 456.600 331.050 457.050 ;
        RECT 319.950 455.400 331.050 456.600 ;
        RECT 319.950 454.950 322.050 455.400 ;
        RECT 328.950 454.950 331.050 455.400 ;
        RECT 334.950 456.600 337.050 457.050 ;
        RECT 343.950 456.600 346.050 457.050 ;
        RECT 352.950 456.600 355.050 457.050 ;
        RECT 334.950 455.400 346.050 456.600 ;
        RECT 334.950 454.950 337.050 455.400 ;
        RECT 343.950 454.950 346.050 455.400 ;
        RECT 350.400 455.400 355.050 456.600 ;
        RECT 280.950 452.400 291.600 453.600 ;
        RECT 307.950 453.600 310.050 454.050 ;
        RECT 310.950 453.600 313.050 454.050 ;
        RECT 316.950 453.600 319.050 454.050 ;
        RECT 307.950 452.400 319.050 453.600 ;
        RECT 280.950 451.950 283.050 452.400 ;
        RECT 307.950 451.950 310.050 452.400 ;
        RECT 310.950 451.950 313.050 452.400 ;
        RECT 316.950 451.950 319.050 452.400 ;
        RECT 322.950 453.600 325.050 454.050 ;
        RECT 331.950 453.600 334.050 454.050 ;
        RECT 322.950 452.400 334.050 453.600 ;
        RECT 322.950 451.950 325.050 452.400 ;
        RECT 331.950 451.950 334.050 452.400 ;
        RECT 346.950 451.950 349.050 454.050 ;
        RECT 232.950 450.600 235.050 451.050 ;
        RECT 230.400 449.400 235.050 450.600 ;
        RECT 190.950 448.950 193.050 449.400 ;
        RECT 211.950 448.950 214.050 449.400 ;
        RECT 220.950 448.950 223.050 449.400 ;
        RECT 232.950 448.950 235.050 449.400 ;
        RECT 253.950 448.950 256.050 451.050 ;
        RECT 268.950 448.950 271.050 451.050 ;
        RECT 100.950 446.400 105.600 447.600 ;
        RECT 115.950 447.600 118.050 448.050 ;
        RECT 133.950 447.600 136.050 448.050 ;
        RECT 184.950 447.600 187.050 448.050 ;
        RECT 115.950 446.400 187.050 447.600 ;
        RECT 100.950 445.950 103.050 446.400 ;
        RECT 115.950 445.950 118.050 446.400 ;
        RECT 133.950 445.950 136.050 446.400 ;
        RECT 184.950 445.950 187.050 446.400 ;
        RECT 247.950 447.600 250.050 448.050 ;
        RECT 272.400 447.600 273.600 451.950 ;
        RECT 274.950 450.600 277.050 451.050 ;
        RECT 295.950 450.600 298.050 451.050 ;
        RECT 274.950 449.400 298.050 450.600 ;
        RECT 274.950 448.950 277.050 449.400 ;
        RECT 295.950 448.950 298.050 449.400 ;
        RECT 310.950 450.600 313.050 451.050 ;
        RECT 343.950 450.600 346.050 451.050 ;
        RECT 310.950 449.400 346.050 450.600 ;
        RECT 310.950 448.950 313.050 449.400 ;
        RECT 343.950 448.950 346.050 449.400 ;
        RECT 247.950 446.400 273.600 447.600 ;
        RECT 347.400 447.600 348.600 451.950 ;
        RECT 350.400 451.050 351.600 455.400 ;
        RECT 352.950 454.950 355.050 455.400 ;
        RECT 356.400 454.050 357.600 458.400 ;
        RECT 364.950 457.950 367.050 460.050 ;
        RECT 391.950 459.600 394.050 460.050 ;
        RECT 412.950 459.600 415.050 460.050 ;
        RECT 418.950 459.600 421.050 460.050 ;
        RECT 391.950 458.400 421.050 459.600 ;
        RECT 391.950 457.950 394.050 458.400 ;
        RECT 412.950 457.950 415.050 458.400 ;
        RECT 418.950 457.950 421.050 458.400 ;
        RECT 457.950 459.600 460.050 460.050 ;
        RECT 463.950 459.600 466.050 460.050 ;
        RECT 457.950 458.400 466.050 459.600 ;
        RECT 457.950 457.950 460.050 458.400 ;
        RECT 463.950 457.950 466.050 458.400 ;
        RECT 481.950 457.950 484.050 460.050 ;
        RECT 550.950 459.600 553.050 460.050 ;
        RECT 539.400 458.400 553.050 459.600 ;
        RECT 365.400 456.600 366.600 457.950 ;
        RECT 359.400 455.400 366.600 456.600 ;
        RECT 376.950 456.600 379.050 457.050 ;
        RECT 397.950 456.600 400.050 457.050 ;
        RECT 400.950 456.600 403.050 457.050 ;
        RECT 376.950 455.400 403.050 456.600 ;
        RECT 355.950 451.950 358.050 454.050 ;
        RECT 359.400 451.050 360.600 455.400 ;
        RECT 376.950 454.950 379.050 455.400 ;
        RECT 397.950 454.950 400.050 455.400 ;
        RECT 400.950 454.950 403.050 455.400 ;
        RECT 403.950 454.950 406.050 457.050 ;
        RECT 454.950 454.950 457.050 457.050 ;
        RECT 460.950 456.600 463.050 457.050 ;
        RECT 478.950 456.600 481.050 457.050 ;
        RECT 460.950 455.400 481.050 456.600 ;
        RECT 460.950 454.950 463.050 455.400 ;
        RECT 361.950 453.600 364.050 454.050 ;
        RECT 367.950 453.600 370.050 454.050 ;
        RECT 361.950 452.400 370.050 453.600 ;
        RECT 361.950 451.950 364.050 452.400 ;
        RECT 367.950 451.950 370.050 452.400 ;
        RECT 370.950 453.600 373.050 454.050 ;
        RECT 379.950 453.600 382.050 454.050 ;
        RECT 370.950 452.400 382.050 453.600 ;
        RECT 370.950 451.950 373.050 452.400 ;
        RECT 379.950 451.950 382.050 452.400 ;
        RECT 349.950 448.950 352.050 451.050 ;
        RECT 358.950 448.950 361.050 451.050 ;
        RECT 379.950 450.600 382.050 451.050 ;
        RECT 404.400 450.600 405.600 454.950 ;
        RECT 406.950 451.950 409.050 454.050 ;
        RECT 455.400 453.600 456.600 454.950 ;
        RECT 476.400 454.050 477.600 455.400 ;
        RECT 478.950 454.950 481.050 455.400 ;
        RECT 472.950 453.600 475.050 454.050 ;
        RECT 455.400 452.400 475.050 453.600 ;
        RECT 472.950 451.950 475.050 452.400 ;
        RECT 475.950 451.950 478.050 454.050 ;
        RECT 482.400 453.600 483.600 457.950 ;
        RECT 502.950 456.600 505.050 457.050 ;
        RECT 514.950 456.600 517.050 457.050 ;
        RECT 502.950 455.400 517.050 456.600 ;
        RECT 502.950 454.950 505.050 455.400 ;
        RECT 514.950 454.950 517.050 455.400 ;
        RECT 479.400 452.400 483.600 453.600 ;
        RECT 379.950 449.400 405.600 450.600 ;
        RECT 379.950 448.950 382.050 449.400 ;
        RECT 367.950 447.600 370.050 448.050 ;
        RECT 347.400 446.400 370.050 447.600 ;
        RECT 247.950 445.950 250.050 446.400 ;
        RECT 367.950 445.950 370.050 446.400 ;
        RECT 388.950 447.600 391.050 448.050 ;
        RECT 407.400 447.600 408.600 451.950 ;
        RECT 409.950 450.600 412.050 451.050 ;
        RECT 424.950 450.600 427.050 451.050 ;
        RECT 409.950 449.400 427.050 450.600 ;
        RECT 409.950 448.950 412.050 449.400 ;
        RECT 424.950 448.950 427.050 449.400 ;
        RECT 448.950 450.600 451.050 451.050 ;
        RECT 454.950 450.600 457.050 451.050 ;
        RECT 448.950 449.400 457.050 450.600 ;
        RECT 448.950 448.950 451.050 449.400 ;
        RECT 454.950 448.950 457.050 449.400 ;
        RECT 469.950 450.600 472.050 451.050 ;
        RECT 479.400 450.600 480.600 452.400 ;
        RECT 469.950 449.400 480.600 450.600 ;
        RECT 493.950 450.600 496.050 451.050 ;
        RECT 508.950 450.600 511.050 451.050 ;
        RECT 493.950 449.400 511.050 450.600 ;
        RECT 469.950 448.950 472.050 449.400 ;
        RECT 493.950 448.950 496.050 449.400 ;
        RECT 508.950 448.950 511.050 449.400 ;
        RECT 388.950 446.400 408.600 447.600 ;
        RECT 445.950 447.600 448.050 448.050 ;
        RECT 457.950 447.600 460.050 448.050 ;
        RECT 487.950 447.600 490.050 448.050 ;
        RECT 445.950 446.400 490.050 447.600 ;
        RECT 539.400 447.600 540.600 458.400 ;
        RECT 550.950 457.950 553.050 458.400 ;
        RECT 583.950 457.950 586.050 460.050 ;
        RECT 587.400 459.600 588.600 461.400 ;
        RECT 595.950 461.400 604.050 462.600 ;
        RECT 595.950 460.950 598.050 461.400 ;
        RECT 601.950 460.950 604.050 461.400 ;
        RECT 604.950 462.600 607.050 463.050 ;
        RECT 619.950 462.600 622.050 463.050 ;
        RECT 646.950 462.600 649.050 463.050 ;
        RECT 661.950 462.600 664.050 463.050 ;
        RECT 604.950 461.400 649.050 462.600 ;
        RECT 604.950 460.950 607.050 461.400 ;
        RECT 619.950 460.950 622.050 461.400 ;
        RECT 646.950 460.950 649.050 461.400 ;
        RECT 656.400 461.400 664.050 462.600 ;
        RECT 613.950 459.600 616.050 460.050 ;
        RECT 628.950 459.600 631.050 460.050 ;
        RECT 634.950 459.600 637.050 460.050 ;
        RECT 649.950 459.600 652.050 460.050 ;
        RECT 587.400 458.400 652.050 459.600 ;
        RECT 613.950 457.950 616.050 458.400 ;
        RECT 628.950 457.950 631.050 458.400 ;
        RECT 634.950 457.950 637.050 458.400 ;
        RECT 649.950 457.950 652.050 458.400 ;
        RECT 544.950 456.600 547.050 457.050 ;
        RECT 550.950 456.600 553.050 457.050 ;
        RECT 544.950 455.400 553.050 456.600 ;
        RECT 544.950 454.950 547.050 455.400 ;
        RECT 550.950 454.950 553.050 455.400 ;
        RECT 556.950 456.600 559.050 457.050 ;
        RECT 562.950 456.600 565.050 457.050 ;
        RECT 556.950 455.400 565.050 456.600 ;
        RECT 556.950 454.950 559.050 455.400 ;
        RECT 562.950 454.950 565.050 455.400 ;
        RECT 568.950 454.950 571.050 457.050 ;
        RECT 577.950 456.600 580.050 457.050 ;
        RECT 584.400 456.600 585.600 457.950 ;
        RECT 592.950 456.600 595.050 457.050 ;
        RECT 610.950 456.600 613.050 457.050 ;
        RECT 577.950 455.400 582.600 456.600 ;
        RECT 584.400 455.400 591.600 456.600 ;
        RECT 577.950 454.950 580.050 455.400 ;
        RECT 541.950 453.600 544.050 454.050 ;
        RECT 565.950 453.600 568.050 454.050 ;
        RECT 569.400 453.600 570.600 454.950 ;
        RECT 541.950 452.400 570.600 453.600 ;
        RECT 571.950 453.600 574.050 454.050 ;
        RECT 577.950 453.600 580.050 454.050 ;
        RECT 571.950 452.400 580.050 453.600 ;
        RECT 581.400 453.600 582.600 455.400 ;
        RECT 583.950 453.600 586.050 454.050 ;
        RECT 581.400 452.400 586.050 453.600 ;
        RECT 590.400 453.600 591.600 455.400 ;
        RECT 592.950 455.400 597.600 456.600 ;
        RECT 592.950 454.950 595.050 455.400 ;
        RECT 590.400 452.400 594.600 453.600 ;
        RECT 541.950 451.950 544.050 452.400 ;
        RECT 565.950 451.950 568.050 452.400 ;
        RECT 571.950 451.950 574.050 452.400 ;
        RECT 577.950 451.950 580.050 452.400 ;
        RECT 583.950 451.950 586.050 452.400 ;
        RECT 547.950 450.600 550.050 451.050 ;
        RECT 556.950 450.600 559.050 451.050 ;
        RECT 547.950 449.400 559.050 450.600 ;
        RECT 547.950 448.950 550.050 449.400 ;
        RECT 556.950 448.950 559.050 449.400 ;
        RECT 556.950 447.600 559.050 448.050 ;
        RECT 539.400 446.400 559.050 447.600 ;
        RECT 593.400 447.600 594.600 452.400 ;
        RECT 596.400 451.050 597.600 455.400 ;
        RECT 610.950 455.400 621.600 456.600 ;
        RECT 610.950 454.950 613.050 455.400 ;
        RECT 598.950 453.600 601.050 454.050 ;
        RECT 607.950 453.600 610.050 454.050 ;
        RECT 616.950 453.600 619.050 454.050 ;
        RECT 598.950 452.400 603.600 453.600 ;
        RECT 598.950 451.950 601.050 452.400 ;
        RECT 595.950 448.950 598.050 451.050 ;
        RECT 602.400 450.600 603.600 452.400 ;
        RECT 607.950 452.400 619.050 453.600 ;
        RECT 607.950 451.950 610.050 452.400 ;
        RECT 616.950 451.950 619.050 452.400 ;
        RECT 620.400 451.050 621.600 455.400 ;
        RECT 625.950 454.950 628.050 457.050 ;
        RECT 643.950 456.600 646.050 457.050 ;
        RECT 652.950 456.600 655.050 457.050 ;
        RECT 638.400 455.400 646.050 456.600 ;
        RECT 626.400 451.050 627.600 454.950 ;
        RECT 634.950 453.600 637.050 454.050 ;
        RECT 638.400 453.600 639.600 455.400 ;
        RECT 643.950 454.950 646.050 455.400 ;
        RECT 647.400 455.400 655.050 456.600 ;
        RECT 656.400 456.600 657.600 461.400 ;
        RECT 661.950 460.950 664.050 461.400 ;
        RECT 670.950 462.600 673.050 463.050 ;
        RECT 673.950 462.600 676.050 463.050 ;
        RECT 694.950 462.600 697.050 463.050 ;
        RECT 670.950 461.400 697.050 462.600 ;
        RECT 670.950 460.950 673.050 461.400 ;
        RECT 673.950 460.950 676.050 461.400 ;
        RECT 694.950 460.950 697.050 461.400 ;
        RECT 697.950 462.600 700.050 463.050 ;
        RECT 715.950 462.600 718.050 463.050 ;
        RECT 697.950 461.400 718.050 462.600 ;
        RECT 697.950 460.950 700.050 461.400 ;
        RECT 715.950 460.950 718.050 461.400 ;
        RECT 658.950 459.600 661.050 460.050 ;
        RECT 700.950 459.600 703.050 460.050 ;
        RECT 709.950 459.600 712.050 460.050 ;
        RECT 658.950 458.400 681.600 459.600 ;
        RECT 658.950 457.950 661.050 458.400 ;
        RECT 680.400 457.050 681.600 458.400 ;
        RECT 700.950 458.400 712.050 459.600 ;
        RECT 700.950 457.950 703.050 458.400 ;
        RECT 709.950 457.950 712.050 458.400 ;
        RECT 715.950 459.600 718.050 460.050 ;
        RECT 719.400 459.600 720.600 464.400 ;
        RECT 715.950 458.400 720.600 459.600 ;
        RECT 715.950 457.950 718.050 458.400 ;
        RECT 661.950 456.600 664.050 457.050 ;
        RECT 656.400 455.400 660.600 456.600 ;
        RECT 643.950 453.600 646.050 454.050 ;
        RECT 634.950 452.400 639.600 453.600 ;
        RECT 641.400 452.400 646.050 453.600 ;
        RECT 634.950 451.950 637.050 452.400 ;
        RECT 616.950 450.600 619.050 451.050 ;
        RECT 602.400 449.400 619.050 450.600 ;
        RECT 616.950 448.950 619.050 449.400 ;
        RECT 619.950 448.950 622.050 451.050 ;
        RECT 625.950 448.950 628.050 451.050 ;
        RECT 641.400 448.050 642.600 452.400 ;
        RECT 643.950 451.950 646.050 452.400 ;
        RECT 647.400 450.600 648.600 455.400 ;
        RECT 652.950 454.950 655.050 455.400 ;
        RECT 659.400 453.600 660.600 455.400 ;
        RECT 661.950 455.400 666.600 456.600 ;
        RECT 661.950 454.950 664.050 455.400 ;
        RECT 661.950 453.600 664.050 454.050 ;
        RECT 659.400 452.400 664.050 453.600 ;
        RECT 665.400 453.600 666.600 455.400 ;
        RECT 679.950 454.950 682.050 457.050 ;
        RECT 691.950 456.600 694.050 457.050 ;
        RECT 700.950 456.600 703.050 457.050 ;
        RECT 691.950 455.400 703.050 456.600 ;
        RECT 691.950 454.950 694.050 455.400 ;
        RECT 700.950 454.950 703.050 455.400 ;
        RECT 691.950 453.600 694.050 454.050 ;
        RECT 665.400 452.400 694.050 453.600 ;
        RECT 661.950 451.950 664.050 452.400 ;
        RECT 691.950 451.950 694.050 452.400 ;
        RECT 703.950 453.600 706.050 454.050 ;
        RECT 709.950 453.600 712.050 454.050 ;
        RECT 703.950 452.400 712.050 453.600 ;
        RECT 703.950 451.950 706.050 452.400 ;
        RECT 709.950 451.950 712.050 452.400 ;
        RECT 644.400 449.400 648.600 450.600 ;
        RECT 652.950 450.600 655.050 451.050 ;
        RECT 688.950 450.600 691.050 451.050 ;
        RECT 697.950 450.600 700.050 451.050 ;
        RECT 700.950 450.600 703.050 451.050 ;
        RECT 652.950 449.400 703.050 450.600 ;
        RECT 644.400 448.050 645.600 449.400 ;
        RECT 652.950 448.950 655.050 449.400 ;
        RECT 688.950 448.950 691.050 449.400 ;
        RECT 697.950 448.950 700.050 449.400 ;
        RECT 700.950 448.950 703.050 449.400 ;
        RECT 613.950 447.600 616.050 448.050 ;
        RECT 593.400 446.400 616.050 447.600 ;
        RECT 388.950 445.950 391.050 446.400 ;
        RECT 445.950 445.950 448.050 446.400 ;
        RECT 457.950 445.950 460.050 446.400 ;
        RECT 487.950 445.950 490.050 446.400 ;
        RECT 556.950 445.950 559.050 446.400 ;
        RECT 613.950 445.950 616.050 446.400 ;
        RECT 640.950 445.950 643.050 448.050 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 682.950 447.600 685.050 448.050 ;
        RECT 703.950 447.600 706.050 448.050 ;
        RECT 682.950 446.400 706.050 447.600 ;
        RECT 682.950 445.950 685.050 446.400 ;
        RECT 703.950 445.950 706.050 446.400 ;
        RECT 64.950 444.600 67.050 445.050 ;
        RECT 103.950 444.600 106.050 445.050 ;
        RECT 64.950 443.400 106.050 444.600 ;
        RECT 64.950 442.950 67.050 443.400 ;
        RECT 103.950 442.950 106.050 443.400 ;
        RECT 106.950 444.600 109.050 445.050 ;
        RECT 130.950 444.600 133.050 445.050 ;
        RECT 106.950 443.400 133.050 444.600 ;
        RECT 106.950 442.950 109.050 443.400 ;
        RECT 130.950 442.950 133.050 443.400 ;
        RECT 151.950 444.600 154.050 445.050 ;
        RECT 157.950 444.600 160.050 445.050 ;
        RECT 151.950 443.400 160.050 444.600 ;
        RECT 151.950 442.950 154.050 443.400 ;
        RECT 157.950 442.950 160.050 443.400 ;
        RECT 193.950 444.600 196.050 445.050 ;
        RECT 238.950 444.600 241.050 445.050 ;
        RECT 193.950 443.400 241.050 444.600 ;
        RECT 193.950 442.950 196.050 443.400 ;
        RECT 238.950 442.950 241.050 443.400 ;
        RECT 505.950 444.600 508.050 445.050 ;
        RECT 571.950 444.600 574.050 445.050 ;
        RECT 505.950 443.400 574.050 444.600 ;
        RECT 505.950 442.950 508.050 443.400 ;
        RECT 571.950 442.950 574.050 443.400 ;
        RECT 622.950 444.600 625.050 445.050 ;
        RECT 661.950 444.600 664.050 445.050 ;
        RECT 622.950 443.400 664.050 444.600 ;
        RECT 622.950 442.950 625.050 443.400 ;
        RECT 661.950 442.950 664.050 443.400 ;
        RECT 1.950 441.600 4.050 442.050 ;
        RECT 25.950 441.600 28.050 442.050 ;
        RECT 1.950 440.400 28.050 441.600 ;
        RECT 1.950 439.950 4.050 440.400 ;
        RECT 25.950 439.950 28.050 440.400 ;
        RECT 73.950 441.600 76.050 442.050 ;
        RECT 91.950 441.600 94.050 442.050 ;
        RECT 112.950 441.600 115.050 442.050 ;
        RECT 73.950 440.400 115.050 441.600 ;
        RECT 73.950 439.950 76.050 440.400 ;
        RECT 91.950 439.950 94.050 440.400 ;
        RECT 112.950 439.950 115.050 440.400 ;
        RECT 142.950 441.600 145.050 442.050 ;
        RECT 163.950 441.600 166.050 442.050 ;
        RECT 268.950 441.600 271.050 442.050 ;
        RECT 142.950 440.400 271.050 441.600 ;
        RECT 142.950 439.950 145.050 440.400 ;
        RECT 163.950 439.950 166.050 440.400 ;
        RECT 268.950 439.950 271.050 440.400 ;
        RECT 463.950 441.600 466.050 442.050 ;
        RECT 514.950 441.600 517.050 442.050 ;
        RECT 463.950 440.400 517.050 441.600 ;
        RECT 463.950 439.950 466.050 440.400 ;
        RECT 514.950 439.950 517.050 440.400 ;
        RECT 634.950 441.600 637.050 442.050 ;
        RECT 646.950 441.600 649.050 442.050 ;
        RECT 634.950 440.400 649.050 441.600 ;
        RECT 634.950 439.950 637.050 440.400 ;
        RECT 646.950 439.950 649.050 440.400 ;
        RECT 7.950 438.600 10.050 439.050 ;
        RECT 46.950 438.600 49.050 439.050 ;
        RECT 7.950 437.400 49.050 438.600 ;
        RECT 7.950 436.950 10.050 437.400 ;
        RECT 46.950 436.950 49.050 437.400 ;
        RECT 82.950 438.600 85.050 439.050 ;
        RECT 217.950 438.600 220.050 439.050 ;
        RECT 82.950 437.400 220.050 438.600 ;
        RECT 82.950 436.950 85.050 437.400 ;
        RECT 217.950 436.950 220.050 437.400 ;
        RECT 223.950 438.600 226.050 439.050 ;
        RECT 253.950 438.600 256.050 439.050 ;
        RECT 223.950 437.400 256.050 438.600 ;
        RECT 223.950 436.950 226.050 437.400 ;
        RECT 253.950 436.950 256.050 437.400 ;
        RECT 559.950 438.600 562.050 439.050 ;
        RECT 565.950 438.600 568.050 439.050 ;
        RECT 559.950 437.400 568.050 438.600 ;
        RECT 559.950 436.950 562.050 437.400 ;
        RECT 565.950 436.950 568.050 437.400 ;
        RECT 640.950 438.600 643.050 439.050 ;
        RECT 691.950 438.600 694.050 439.050 ;
        RECT 715.950 438.600 718.050 439.050 ;
        RECT 640.950 437.400 718.050 438.600 ;
        RECT 640.950 436.950 643.050 437.400 ;
        RECT 691.950 436.950 694.050 437.400 ;
        RECT 715.950 436.950 718.050 437.400 ;
        RECT 37.950 435.600 40.050 436.050 ;
        RECT 85.950 435.600 88.050 436.050 ;
        RECT 37.950 434.400 88.050 435.600 ;
        RECT 37.950 433.950 40.050 434.400 ;
        RECT 85.950 433.950 88.050 434.400 ;
        RECT 97.950 435.600 100.050 436.050 ;
        RECT 130.950 435.600 133.050 436.050 ;
        RECT 253.950 435.600 256.050 436.050 ;
        RECT 97.950 434.400 133.050 435.600 ;
        RECT 97.950 433.950 100.050 434.400 ;
        RECT 130.950 433.950 133.050 434.400 ;
        RECT 134.400 434.400 256.050 435.600 ;
        RECT 52.950 432.600 55.050 433.050 ;
        RECT 134.400 432.600 135.600 434.400 ;
        RECT 253.950 433.950 256.050 434.400 ;
        RECT 52.950 431.400 135.600 432.600 ;
        RECT 166.950 432.600 169.050 433.050 ;
        RECT 175.950 432.600 178.050 433.050 ;
        RECT 166.950 431.400 178.050 432.600 ;
        RECT 52.950 430.950 55.050 431.400 ;
        RECT 166.950 430.950 169.050 431.400 ;
        RECT 175.950 430.950 178.050 431.400 ;
        RECT 202.950 432.600 205.050 433.050 ;
        RECT 250.950 432.600 253.050 433.050 ;
        RECT 202.950 431.400 253.050 432.600 ;
        RECT 202.950 430.950 205.050 431.400 ;
        RECT 250.950 430.950 253.050 431.400 ;
        RECT 262.950 432.600 265.050 433.050 ;
        RECT 463.950 432.600 466.050 433.050 ;
        RECT 262.950 431.400 466.050 432.600 ;
        RECT 262.950 430.950 265.050 431.400 ;
        RECT 463.950 430.950 466.050 431.400 ;
        RECT 544.950 432.600 547.050 433.050 ;
        RECT 574.950 432.600 577.050 433.050 ;
        RECT 664.950 432.600 667.050 433.050 ;
        RECT 544.950 431.400 667.050 432.600 ;
        RECT 544.950 430.950 547.050 431.400 ;
        RECT 574.950 430.950 577.050 431.400 ;
        RECT 664.950 430.950 667.050 431.400 ;
        RECT 28.950 429.600 31.050 430.050 ;
        RECT 232.950 429.600 235.050 430.050 ;
        RECT 415.950 429.600 418.050 430.050 ;
        RECT 448.950 429.600 451.050 430.050 ;
        RECT 28.950 428.400 451.050 429.600 ;
        RECT 28.950 427.950 31.050 428.400 ;
        RECT 232.950 427.950 235.050 428.400 ;
        RECT 415.950 427.950 418.050 428.400 ;
        RECT 448.950 427.950 451.050 428.400 ;
        RECT 550.950 429.600 553.050 430.050 ;
        RECT 640.950 429.600 643.050 430.050 ;
        RECT 670.950 429.600 673.050 430.050 ;
        RECT 550.950 428.400 673.050 429.600 ;
        RECT 550.950 427.950 553.050 428.400 ;
        RECT 640.950 427.950 643.050 428.400 ;
        RECT 670.950 427.950 673.050 428.400 ;
        RECT 10.950 426.600 13.050 427.050 ;
        RECT 82.950 426.600 85.050 427.050 ;
        RECT 10.950 425.400 85.050 426.600 ;
        RECT 10.950 424.950 13.050 425.400 ;
        RECT 82.950 424.950 85.050 425.400 ;
        RECT 337.950 426.600 340.050 427.050 ;
        RECT 442.950 426.600 445.050 427.050 ;
        RECT 337.950 425.400 445.050 426.600 ;
        RECT 337.950 424.950 340.050 425.400 ;
        RECT 442.950 424.950 445.050 425.400 ;
        RECT 571.950 426.600 574.050 427.050 ;
        RECT 637.950 426.600 640.050 427.050 ;
        RECT 571.950 425.400 640.050 426.600 ;
        RECT 571.950 424.950 574.050 425.400 ;
        RECT 637.950 424.950 640.050 425.400 ;
        RECT 34.950 423.600 37.050 424.050 ;
        RECT 40.950 423.600 43.050 424.050 ;
        RECT 34.950 422.400 43.050 423.600 ;
        RECT 34.950 421.950 37.050 422.400 ;
        RECT 40.950 421.950 43.050 422.400 ;
        RECT 82.950 423.600 85.050 424.050 ;
        RECT 100.950 423.600 103.050 424.050 ;
        RECT 124.950 423.600 127.050 424.050 ;
        RECT 82.950 422.400 93.600 423.600 ;
        RECT 82.950 421.950 85.050 422.400 ;
        RECT 49.950 420.600 52.050 421.050 ;
        RECT 49.950 419.400 66.600 420.600 ;
        RECT 49.950 418.950 52.050 419.400 ;
        RECT 1.950 417.600 4.050 418.050 ;
        RECT 19.950 417.600 22.050 418.050 ;
        RECT 1.950 416.400 22.050 417.600 ;
        RECT 1.950 415.950 4.050 416.400 ;
        RECT 19.950 415.950 22.050 416.400 ;
        RECT 22.950 415.950 25.050 418.050 ;
        RECT 31.950 415.950 34.050 418.050 ;
        RECT 43.950 417.600 46.050 418.050 ;
        RECT 52.950 417.600 55.050 418.050 ;
        RECT 43.950 416.400 55.050 417.600 ;
        RECT 43.950 415.950 46.050 416.400 ;
        RECT 52.950 415.950 55.050 416.400 ;
        RECT 55.950 417.600 58.050 418.050 ;
        RECT 55.950 416.400 63.600 417.600 ;
        RECT 55.950 415.950 58.050 416.400 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 7.950 412.950 10.050 415.050 ;
        RECT 5.400 409.050 6.600 412.950 ;
        RECT 8.400 411.600 9.600 412.950 ;
        RECT 16.950 411.600 19.050 412.050 ;
        RECT 8.400 410.400 19.050 411.600 ;
        RECT 23.400 411.600 24.600 415.950 ;
        RECT 28.950 412.950 31.050 415.050 ;
        RECT 25.950 411.600 28.050 412.050 ;
        RECT 23.400 410.400 28.050 411.600 ;
        RECT 16.950 409.950 19.050 410.400 ;
        RECT 25.950 409.950 28.050 410.400 ;
        RECT 29.400 409.050 30.600 412.950 ;
        RECT 4.950 406.950 7.050 409.050 ;
        RECT 28.950 406.950 31.050 409.050 ;
        RECT 32.400 408.600 33.600 415.950 ;
        RECT 34.950 414.600 37.050 415.050 ;
        RECT 58.950 414.600 61.050 415.050 ;
        RECT 34.950 413.400 61.050 414.600 ;
        RECT 34.950 412.950 37.050 413.400 ;
        RECT 58.950 412.950 61.050 413.400 ;
        RECT 62.400 412.050 63.600 416.400 ;
        RECT 65.400 414.600 66.600 419.400 ;
        RECT 79.950 418.950 82.050 421.050 ;
        RECT 92.400 420.600 93.600 422.400 ;
        RECT 100.950 422.400 127.050 423.600 ;
        RECT 100.950 421.950 103.050 422.400 ;
        RECT 124.950 421.950 127.050 422.400 ;
        RECT 253.950 423.600 256.050 424.050 ;
        RECT 373.950 423.600 376.050 424.050 ;
        RECT 253.950 422.400 376.050 423.600 ;
        RECT 253.950 421.950 256.050 422.400 ;
        RECT 373.950 421.950 376.050 422.400 ;
        RECT 565.950 423.600 568.050 424.050 ;
        RECT 589.950 423.600 592.050 424.050 ;
        RECT 565.950 422.400 592.050 423.600 ;
        RECT 565.950 421.950 568.050 422.400 ;
        RECT 589.950 421.950 592.050 422.400 ;
        RECT 604.950 423.600 607.050 424.050 ;
        RECT 619.950 423.600 622.050 424.050 ;
        RECT 604.950 422.400 622.050 423.600 ;
        RECT 604.950 421.950 607.050 422.400 ;
        RECT 619.950 421.950 622.050 422.400 ;
        RECT 92.400 419.400 99.600 420.600 ;
        RECT 73.950 414.600 76.050 415.050 ;
        RECT 65.400 413.400 76.050 414.600 ;
        RECT 73.950 412.950 76.050 413.400 ;
        RECT 37.950 411.600 40.050 412.050 ;
        RECT 40.950 411.600 43.050 412.050 ;
        RECT 55.950 411.600 58.050 412.050 ;
        RECT 37.950 410.400 58.050 411.600 ;
        RECT 37.950 409.950 40.050 410.400 ;
        RECT 40.950 409.950 43.050 410.400 ;
        RECT 55.950 409.950 58.050 410.400 ;
        RECT 61.950 409.950 64.050 412.050 ;
        RECT 64.950 411.600 67.050 412.050 ;
        RECT 73.950 411.600 76.050 412.050 ;
        RECT 64.950 410.400 76.050 411.600 ;
        RECT 80.400 411.600 81.600 418.950 ;
        RECT 85.950 415.950 88.050 418.050 ;
        RECT 86.400 412.050 87.600 415.950 ;
        RECT 98.400 414.600 99.600 419.400 ;
        RECT 106.950 418.950 109.050 421.050 ;
        RECT 112.950 420.600 115.050 421.050 ;
        RECT 178.950 420.600 181.050 421.050 ;
        RECT 205.950 420.600 208.050 421.050 ;
        RECT 262.950 420.600 265.050 421.050 ;
        RECT 112.950 419.400 265.050 420.600 ;
        RECT 112.950 418.950 115.050 419.400 ;
        RECT 178.950 418.950 181.050 419.400 ;
        RECT 205.950 418.950 208.050 419.400 ;
        RECT 262.950 418.950 265.050 419.400 ;
        RECT 265.950 420.600 268.050 421.050 ;
        RECT 283.950 420.600 286.050 421.050 ;
        RECT 265.950 419.400 286.050 420.600 ;
        RECT 265.950 418.950 268.050 419.400 ;
        RECT 283.950 418.950 286.050 419.400 ;
        RECT 301.950 420.600 304.050 421.050 ;
        RECT 307.950 420.600 310.050 421.050 ;
        RECT 301.950 419.400 310.050 420.600 ;
        RECT 301.950 418.950 304.050 419.400 ;
        RECT 307.950 418.950 310.050 419.400 ;
        RECT 334.950 420.600 337.050 421.050 ;
        RECT 370.950 420.600 373.050 421.050 ;
        RECT 334.950 419.400 373.050 420.600 ;
        RECT 334.950 418.950 337.050 419.400 ;
        RECT 370.950 418.950 373.050 419.400 ;
        RECT 373.950 420.600 376.050 421.050 ;
        RECT 394.950 420.600 397.050 421.050 ;
        RECT 373.950 419.400 397.050 420.600 ;
        RECT 373.950 418.950 376.050 419.400 ;
        RECT 394.950 418.950 397.050 419.400 ;
        RECT 421.950 420.600 424.050 421.050 ;
        RECT 463.950 420.600 466.050 421.050 ;
        RECT 577.950 420.600 580.050 421.050 ;
        RECT 421.950 419.400 580.050 420.600 ;
        RECT 421.950 418.950 424.050 419.400 ;
        RECT 463.950 418.950 466.050 419.400 ;
        RECT 577.950 418.950 580.050 419.400 ;
        RECT 682.950 420.600 685.050 421.050 ;
        RECT 691.950 420.600 694.050 421.050 ;
        RECT 700.950 420.600 703.050 421.050 ;
        RECT 682.950 419.400 703.050 420.600 ;
        RECT 682.950 418.950 685.050 419.400 ;
        RECT 691.950 418.950 694.050 419.400 ;
        RECT 700.950 418.950 703.050 419.400 ;
        RECT 95.400 413.400 99.600 414.600 ;
        RECT 82.950 411.600 85.050 412.050 ;
        RECT 80.400 410.400 85.050 411.600 ;
        RECT 64.950 409.950 67.050 410.400 ;
        RECT 73.950 409.950 76.050 410.400 ;
        RECT 82.950 409.950 85.050 410.400 ;
        RECT 85.950 409.950 88.050 412.050 ;
        RECT 91.950 411.600 94.050 412.050 ;
        RECT 95.400 411.600 96.600 413.400 ;
        RECT 91.950 410.400 96.600 411.600 ;
        RECT 100.950 411.600 103.050 412.050 ;
        RECT 107.400 411.600 108.600 418.950 ;
        RECT 163.950 417.600 166.050 418.050 ;
        RECT 178.950 417.600 181.050 418.050 ;
        RECT 163.950 416.400 181.050 417.600 ;
        RECT 163.950 415.950 166.050 416.400 ;
        RECT 178.950 415.950 181.050 416.400 ;
        RECT 187.950 417.600 190.050 418.050 ;
        RECT 187.950 416.400 210.600 417.600 ;
        RECT 187.950 415.950 190.050 416.400 ;
        RECT 124.950 414.600 127.050 415.050 ;
        RECT 151.950 414.600 154.050 415.050 ;
        RECT 202.950 414.600 205.050 415.050 ;
        RECT 124.950 413.400 150.600 414.600 ;
        RECT 124.950 412.950 127.050 413.400 ;
        RECT 100.950 410.400 108.600 411.600 ;
        RECT 109.950 411.600 112.050 412.050 ;
        RECT 121.950 411.600 124.050 412.050 ;
        RECT 127.950 411.600 130.050 412.050 ;
        RECT 109.950 410.400 114.600 411.600 ;
        RECT 91.950 409.950 94.050 410.400 ;
        RECT 100.950 409.950 103.050 410.400 ;
        RECT 109.950 409.950 112.050 410.400 ;
        RECT 43.950 408.600 46.050 409.050 ;
        RECT 32.400 407.400 46.050 408.600 ;
        RECT 43.950 406.950 46.050 407.400 ;
        RECT 52.950 408.600 55.050 409.050 ;
        RECT 79.950 408.600 82.050 409.050 ;
        RECT 52.950 407.400 82.050 408.600 ;
        RECT 113.400 408.600 114.600 410.400 ;
        RECT 121.950 410.400 130.050 411.600 ;
        RECT 121.950 409.950 124.050 410.400 ;
        RECT 127.950 409.950 130.050 410.400 ;
        RECT 133.950 411.600 136.050 412.050 ;
        RECT 136.950 411.600 139.050 412.050 ;
        RECT 145.950 411.600 148.050 412.050 ;
        RECT 133.950 410.400 148.050 411.600 ;
        RECT 149.400 411.600 150.600 413.400 ;
        RECT 151.950 413.400 205.050 414.600 ;
        RECT 151.950 412.950 154.050 413.400 ;
        RECT 202.950 412.950 205.050 413.400 ;
        RECT 157.950 411.600 160.050 412.050 ;
        RECT 149.400 410.400 160.050 411.600 ;
        RECT 133.950 409.950 136.050 410.400 ;
        RECT 136.950 409.950 139.050 410.400 ;
        RECT 145.950 409.950 148.050 410.400 ;
        RECT 157.950 409.950 160.050 410.400 ;
        RECT 160.950 411.600 163.050 412.050 ;
        RECT 172.950 411.600 175.050 412.050 ;
        RECT 160.950 410.400 175.050 411.600 ;
        RECT 160.950 409.950 163.050 410.400 ;
        RECT 172.950 409.950 175.050 410.400 ;
        RECT 175.950 411.600 178.050 412.050 ;
        RECT 205.950 411.600 208.050 412.050 ;
        RECT 175.950 410.400 208.050 411.600 ;
        RECT 175.950 409.950 178.050 410.400 ;
        RECT 205.950 409.950 208.050 410.400 ;
        RECT 151.950 408.600 154.050 409.050 ;
        RECT 193.950 408.600 196.050 409.050 ;
        RECT 209.400 408.600 210.600 416.400 ;
        RECT 244.950 415.950 247.050 418.050 ;
        RECT 274.950 415.950 277.050 418.050 ;
        RECT 295.950 417.600 298.050 418.050 ;
        RECT 331.950 417.600 334.050 418.050 ;
        RECT 295.950 416.400 334.050 417.600 ;
        RECT 295.950 415.950 298.050 416.400 ;
        RECT 331.950 415.950 334.050 416.400 ;
        RECT 352.950 417.600 355.050 418.050 ;
        RECT 364.950 417.600 367.050 418.050 ;
        RECT 352.950 416.400 367.050 417.600 ;
        RECT 352.950 415.950 355.050 416.400 ;
        RECT 364.950 415.950 367.050 416.400 ;
        RECT 370.950 417.600 373.050 418.050 ;
        RECT 382.950 417.600 385.050 418.050 ;
        RECT 388.950 417.600 391.050 418.050 ;
        RECT 370.950 416.400 391.050 417.600 ;
        RECT 370.950 415.950 373.050 416.400 ;
        RECT 382.950 415.950 385.050 416.400 ;
        RECT 388.950 415.950 391.050 416.400 ;
        RECT 427.950 417.600 430.050 418.050 ;
        RECT 436.950 417.600 439.050 418.050 ;
        RECT 529.950 417.600 532.050 418.050 ;
        RECT 427.950 416.400 439.050 417.600 ;
        RECT 427.950 415.950 430.050 416.400 ;
        RECT 436.950 415.950 439.050 416.400 ;
        RECT 524.400 416.400 532.050 417.600 ;
        RECT 217.950 414.600 220.050 415.050 ;
        RECT 245.400 414.600 246.600 415.950 ;
        RECT 271.950 414.600 274.050 415.050 ;
        RECT 217.950 413.400 274.050 414.600 ;
        RECT 217.950 412.950 220.050 413.400 ;
        RECT 271.950 412.950 274.050 413.400 ;
        RECT 275.400 412.050 276.600 415.950 ;
        RECT 277.950 414.600 280.050 415.050 ;
        RECT 283.950 414.600 286.050 415.050 ;
        RECT 277.950 413.400 286.050 414.600 ;
        RECT 277.950 412.950 280.050 413.400 ;
        RECT 283.950 412.950 286.050 413.400 ;
        RECT 289.950 414.600 292.050 415.050 ;
        RECT 322.950 414.600 325.050 415.050 ;
        RECT 340.950 414.600 343.050 415.050 ;
        RECT 289.950 413.400 325.050 414.600 ;
        RECT 289.950 412.950 292.050 413.400 ;
        RECT 322.950 412.950 325.050 413.400 ;
        RECT 332.400 413.400 343.050 414.600 ;
        RECT 262.950 409.950 265.050 412.050 ;
        RECT 274.950 409.950 277.050 412.050 ;
        RECT 277.950 411.600 280.050 412.050 ;
        RECT 298.950 411.600 301.050 412.050 ;
        RECT 277.950 410.400 301.050 411.600 ;
        RECT 277.950 409.950 280.050 410.400 ;
        RECT 298.950 409.950 301.050 410.400 ;
        RECT 319.950 411.600 322.050 412.050 ;
        RECT 332.400 411.600 333.600 413.400 ;
        RECT 340.950 412.950 343.050 413.400 ;
        RECT 349.950 414.600 352.050 415.050 ;
        RECT 355.950 414.600 358.050 415.050 ;
        RECT 349.950 413.400 358.050 414.600 ;
        RECT 349.950 412.950 352.050 413.400 ;
        RECT 355.950 412.950 358.050 413.400 ;
        RECT 361.950 412.950 364.050 415.050 ;
        RECT 394.950 414.600 397.050 415.050 ;
        RECT 383.400 413.400 397.050 414.600 ;
        RECT 319.950 410.400 333.600 411.600 ;
        RECT 362.400 411.600 363.600 412.950 ;
        RECT 383.400 412.050 384.600 413.400 ;
        RECT 394.950 412.950 397.050 413.400 ;
        RECT 409.950 412.950 412.050 415.050 ;
        RECT 415.950 414.600 418.050 415.050 ;
        RECT 424.950 414.600 427.050 415.050 ;
        RECT 415.950 413.400 427.050 414.600 ;
        RECT 415.950 412.950 418.050 413.400 ;
        RECT 424.950 412.950 427.050 413.400 ;
        RECT 364.950 411.600 367.050 412.050 ;
        RECT 362.400 410.400 367.050 411.600 ;
        RECT 319.950 409.950 322.050 410.400 ;
        RECT 364.950 409.950 367.050 410.400 ;
        RECT 376.950 411.600 379.050 412.050 ;
        RECT 382.950 411.600 385.050 412.050 ;
        RECT 376.950 410.400 385.050 411.600 ;
        RECT 376.950 409.950 379.050 410.400 ;
        RECT 382.950 409.950 385.050 410.400 ;
        RECT 385.950 411.600 388.050 412.050 ;
        RECT 410.400 411.600 411.600 412.950 ;
        RECT 524.400 412.050 525.600 416.400 ;
        RECT 529.950 415.950 532.050 416.400 ;
        RECT 532.950 417.600 535.050 418.050 ;
        RECT 538.950 417.600 541.050 418.050 ;
        RECT 547.950 417.600 550.050 418.050 ;
        RECT 532.950 416.400 550.050 417.600 ;
        RECT 532.950 415.950 535.050 416.400 ;
        RECT 538.950 415.950 541.050 416.400 ;
        RECT 547.950 415.950 550.050 416.400 ;
        RECT 568.950 417.600 571.050 418.050 ;
        RECT 583.950 417.600 586.050 418.050 ;
        RECT 631.950 417.600 634.050 418.050 ;
        RECT 568.950 416.400 586.050 417.600 ;
        RECT 568.950 415.950 571.050 416.400 ;
        RECT 583.950 415.950 586.050 416.400 ;
        RECT 593.400 416.400 621.600 417.600 ;
        RECT 385.950 410.400 411.600 411.600 ;
        RECT 412.950 411.600 415.050 412.050 ;
        RECT 445.950 411.600 448.050 412.050 ;
        RECT 412.950 410.400 448.050 411.600 ;
        RECT 385.950 409.950 388.050 410.400 ;
        RECT 412.950 409.950 415.050 410.400 ;
        RECT 445.950 409.950 448.050 410.400 ;
        RECT 523.950 409.950 526.050 412.050 ;
        RECT 538.950 411.600 541.050 412.050 ;
        RECT 547.950 411.600 550.050 412.050 ;
        RECT 538.950 410.400 550.050 411.600 ;
        RECT 538.950 409.950 541.050 410.400 ;
        RECT 547.950 409.950 550.050 410.400 ;
        RECT 580.950 411.600 583.050 412.050 ;
        RECT 593.400 411.600 594.600 416.400 ;
        RECT 620.400 415.050 621.600 416.400 ;
        RECT 629.400 416.400 634.050 417.600 ;
        RECT 595.950 414.600 598.050 415.050 ;
        RECT 595.950 413.400 603.600 414.600 ;
        RECT 595.950 412.950 598.050 413.400 ;
        RECT 580.950 410.400 594.600 411.600 ;
        RECT 602.400 411.600 603.600 413.400 ;
        RECT 619.950 412.950 622.050 415.050 ;
        RECT 629.400 414.600 630.600 416.400 ;
        RECT 631.950 415.950 634.050 416.400 ;
        RECT 673.950 417.600 676.050 418.050 ;
        RECT 694.950 417.600 697.050 418.050 ;
        RECT 673.950 416.400 697.050 417.600 ;
        RECT 673.950 415.950 676.050 416.400 ;
        RECT 694.950 415.950 697.050 416.400 ;
        RECT 626.400 413.400 630.600 414.600 ;
        RECT 607.950 411.600 610.050 412.050 ;
        RECT 626.400 411.600 627.600 413.400 ;
        RECT 695.400 412.050 696.600 415.950 ;
        RECT 602.400 410.400 606.600 411.600 ;
        RECT 580.950 409.950 583.050 410.400 ;
        RECT 113.400 407.400 120.600 408.600 ;
        RECT 52.950 406.950 55.050 407.400 ;
        RECT 79.950 406.950 82.050 407.400 ;
        RECT 1.950 405.600 4.050 406.050 ;
        RECT 7.950 405.600 10.050 406.050 ;
        RECT 31.950 405.600 34.050 406.050 ;
        RECT 1.950 404.400 34.050 405.600 ;
        RECT 1.950 403.950 4.050 404.400 ;
        RECT 7.950 403.950 10.050 404.400 ;
        RECT 31.950 403.950 34.050 404.400 ;
        RECT 49.950 405.600 52.050 406.050 ;
        RECT 91.950 405.600 94.050 406.050 ;
        RECT 49.950 404.400 94.050 405.600 ;
        RECT 49.950 403.950 52.050 404.400 ;
        RECT 91.950 403.950 94.050 404.400 ;
        RECT 97.950 405.600 100.050 406.050 ;
        RECT 115.950 405.600 118.050 406.050 ;
        RECT 97.950 404.400 118.050 405.600 ;
        RECT 119.400 405.600 120.600 407.400 ;
        RECT 151.950 407.400 196.050 408.600 ;
        RECT 151.950 406.950 154.050 407.400 ;
        RECT 193.950 406.950 196.050 407.400 ;
        RECT 197.400 407.400 210.600 408.600 ;
        RECT 263.400 408.600 264.600 409.950 ;
        RECT 283.950 408.600 286.050 409.050 ;
        RECT 313.950 408.600 316.050 409.050 ;
        RECT 263.400 407.400 316.050 408.600 ;
        RECT 154.950 405.600 157.050 406.050 ;
        RECT 166.950 405.600 169.050 406.050 ;
        RECT 181.950 405.600 184.050 406.050 ;
        RECT 119.400 404.400 184.050 405.600 ;
        RECT 97.950 403.950 100.050 404.400 ;
        RECT 115.950 403.950 118.050 404.400 ;
        RECT 154.950 403.950 157.050 404.400 ;
        RECT 166.950 403.950 169.050 404.400 ;
        RECT 181.950 403.950 184.050 404.400 ;
        RECT 187.950 405.600 190.050 406.050 ;
        RECT 197.400 405.600 198.600 407.400 ;
        RECT 283.950 406.950 286.050 407.400 ;
        RECT 313.950 406.950 316.050 407.400 ;
        RECT 328.950 408.600 331.050 409.050 ;
        RECT 337.950 408.600 340.050 409.050 ;
        RECT 346.950 408.600 349.050 409.050 ;
        RECT 328.950 407.400 349.050 408.600 ;
        RECT 328.950 406.950 331.050 407.400 ;
        RECT 337.950 406.950 340.050 407.400 ;
        RECT 346.950 406.950 349.050 407.400 ;
        RECT 397.950 408.600 400.050 409.050 ;
        RECT 406.950 408.600 409.050 409.050 ;
        RECT 397.950 407.400 409.050 408.600 ;
        RECT 397.950 406.950 400.050 407.400 ;
        RECT 406.950 406.950 409.050 407.400 ;
        RECT 430.950 408.600 433.050 409.050 ;
        RECT 451.950 408.600 454.050 409.050 ;
        RECT 487.950 408.600 490.050 409.050 ;
        RECT 430.950 407.400 490.050 408.600 ;
        RECT 430.950 406.950 433.050 407.400 ;
        RECT 451.950 406.950 454.050 407.400 ;
        RECT 487.950 406.950 490.050 407.400 ;
        RECT 511.950 408.600 514.050 409.050 ;
        RECT 514.950 408.600 517.050 409.050 ;
        RECT 574.950 408.600 577.050 409.050 ;
        RECT 511.950 407.400 577.050 408.600 ;
        RECT 511.950 406.950 514.050 407.400 ;
        RECT 514.950 406.950 517.050 407.400 ;
        RECT 574.950 406.950 577.050 407.400 ;
        RECT 595.950 408.600 598.050 409.050 ;
        RECT 601.950 408.600 604.050 409.050 ;
        RECT 595.950 407.400 604.050 408.600 ;
        RECT 605.400 408.600 606.600 410.400 ;
        RECT 607.950 410.400 627.600 411.600 ;
        RECT 655.950 411.600 658.050 412.050 ;
        RECT 685.950 411.600 688.050 412.050 ;
        RECT 655.950 410.400 688.050 411.600 ;
        RECT 607.950 409.950 610.050 410.400 ;
        RECT 655.950 409.950 658.050 410.400 ;
        RECT 685.950 409.950 688.050 410.400 ;
        RECT 694.950 409.950 697.050 412.050 ;
        RECT 700.950 411.600 703.050 412.050 ;
        RECT 712.950 411.600 715.050 412.050 ;
        RECT 700.950 410.400 715.050 411.600 ;
        RECT 700.950 409.950 703.050 410.400 ;
        RECT 712.950 409.950 715.050 410.400 ;
        RECT 607.950 408.600 610.050 409.050 ;
        RECT 605.400 407.400 610.050 408.600 ;
        RECT 595.950 406.950 598.050 407.400 ;
        RECT 601.950 406.950 604.050 407.400 ;
        RECT 607.950 406.950 610.050 407.400 ;
        RECT 616.950 408.600 619.050 409.050 ;
        RECT 625.950 408.600 628.050 409.050 ;
        RECT 616.950 407.400 628.050 408.600 ;
        RECT 616.950 406.950 619.050 407.400 ;
        RECT 625.950 406.950 628.050 407.400 ;
        RECT 628.950 408.600 631.050 409.050 ;
        RECT 634.950 408.600 637.050 409.050 ;
        RECT 628.950 407.400 637.050 408.600 ;
        RECT 628.950 406.950 631.050 407.400 ;
        RECT 634.950 406.950 637.050 407.400 ;
        RECT 640.950 408.600 643.050 409.050 ;
        RECT 661.950 408.600 664.050 409.050 ;
        RECT 640.950 407.400 664.050 408.600 ;
        RECT 640.950 406.950 643.050 407.400 ;
        RECT 661.950 406.950 664.050 407.400 ;
        RECT 664.950 408.600 667.050 409.050 ;
        RECT 679.950 408.600 682.050 409.050 ;
        RECT 664.950 407.400 682.050 408.600 ;
        RECT 664.950 406.950 667.050 407.400 ;
        RECT 679.950 406.950 682.050 407.400 ;
        RECT 688.950 408.600 691.050 409.050 ;
        RECT 697.950 408.600 700.050 409.050 ;
        RECT 688.950 407.400 700.050 408.600 ;
        RECT 688.950 406.950 691.050 407.400 ;
        RECT 697.950 406.950 700.050 407.400 ;
        RECT 187.950 404.400 198.600 405.600 ;
        RECT 244.950 405.600 247.050 406.050 ;
        RECT 277.950 405.600 280.050 406.050 ;
        RECT 244.950 404.400 280.050 405.600 ;
        RECT 187.950 403.950 190.050 404.400 ;
        RECT 244.950 403.950 247.050 404.400 ;
        RECT 277.950 403.950 280.050 404.400 ;
        RECT 292.950 405.600 295.050 406.050 ;
        RECT 307.950 405.600 310.050 406.050 ;
        RECT 292.950 404.400 310.050 405.600 ;
        RECT 292.950 403.950 295.050 404.400 ;
        RECT 307.950 403.950 310.050 404.400 ;
        RECT 340.950 405.600 343.050 406.050 ;
        RECT 367.950 405.600 370.050 406.050 ;
        RECT 379.950 405.600 382.050 406.050 ;
        RECT 340.950 404.400 382.050 405.600 ;
        RECT 340.950 403.950 343.050 404.400 ;
        RECT 367.950 403.950 370.050 404.400 ;
        RECT 379.950 403.950 382.050 404.400 ;
        RECT 406.950 405.600 409.050 406.050 ;
        RECT 418.950 405.600 421.050 406.050 ;
        RECT 406.950 404.400 421.050 405.600 ;
        RECT 406.950 403.950 409.050 404.400 ;
        RECT 418.950 403.950 421.050 404.400 ;
        RECT 466.950 405.600 469.050 406.050 ;
        RECT 481.950 405.600 484.050 406.050 ;
        RECT 466.950 404.400 484.050 405.600 ;
        RECT 466.950 403.950 469.050 404.400 ;
        RECT 481.950 403.950 484.050 404.400 ;
        RECT 523.950 405.600 526.050 406.050 ;
        RECT 559.950 405.600 562.050 406.050 ;
        RECT 577.950 405.600 580.050 406.050 ;
        RECT 583.950 405.600 586.050 406.050 ;
        RECT 523.950 404.400 586.050 405.600 ;
        RECT 523.950 403.950 526.050 404.400 ;
        RECT 559.950 403.950 562.050 404.400 ;
        RECT 577.950 403.950 580.050 404.400 ;
        RECT 583.950 403.950 586.050 404.400 ;
        RECT 589.950 405.600 592.050 406.050 ;
        RECT 598.950 405.600 601.050 406.050 ;
        RECT 589.950 404.400 601.050 405.600 ;
        RECT 589.950 403.950 592.050 404.400 ;
        RECT 598.950 403.950 601.050 404.400 ;
        RECT 610.950 405.600 613.050 406.050 ;
        RECT 616.950 405.600 619.050 406.050 ;
        RECT 610.950 404.400 619.050 405.600 ;
        RECT 610.950 403.950 613.050 404.400 ;
        RECT 616.950 403.950 619.050 404.400 ;
        RECT 634.950 405.600 637.050 406.050 ;
        RECT 646.950 405.600 649.050 406.050 ;
        RECT 634.950 404.400 649.050 405.600 ;
        RECT 634.950 403.950 637.050 404.400 ;
        RECT 646.950 403.950 649.050 404.400 ;
        RECT 682.950 405.600 685.050 406.050 ;
        RECT 703.950 405.600 706.050 406.050 ;
        RECT 682.950 404.400 706.050 405.600 ;
        RECT 682.950 403.950 685.050 404.400 ;
        RECT 703.950 403.950 706.050 404.400 ;
        RECT 253.950 402.600 256.050 403.050 ;
        RECT 224.400 401.400 256.050 402.600 ;
        RECT 7.950 399.600 10.050 400.050 ;
        RECT 13.950 399.600 16.050 400.050 ;
        RECT 46.950 399.600 49.050 400.050 ;
        RECT 7.950 398.400 49.050 399.600 ;
        RECT 7.950 397.950 10.050 398.400 ;
        RECT 13.950 397.950 16.050 398.400 ;
        RECT 46.950 397.950 49.050 398.400 ;
        RECT 61.950 399.600 64.050 400.050 ;
        RECT 121.950 399.600 124.050 400.050 ;
        RECT 61.950 398.400 124.050 399.600 ;
        RECT 61.950 397.950 64.050 398.400 ;
        RECT 121.950 397.950 124.050 398.400 ;
        RECT 124.950 399.600 127.050 400.050 ;
        RECT 145.950 399.600 148.050 400.050 ;
        RECT 124.950 398.400 148.050 399.600 ;
        RECT 124.950 397.950 127.050 398.400 ;
        RECT 145.950 397.950 148.050 398.400 ;
        RECT 199.950 399.600 202.050 400.050 ;
        RECT 224.400 399.600 225.600 401.400 ;
        RECT 253.950 400.950 256.050 401.400 ;
        RECT 265.950 402.600 268.050 403.050 ;
        RECT 286.950 402.600 289.050 403.050 ;
        RECT 265.950 401.400 289.050 402.600 ;
        RECT 265.950 400.950 268.050 401.400 ;
        RECT 286.950 400.950 289.050 401.400 ;
        RECT 304.950 402.600 307.050 403.050 ;
        RECT 313.950 402.600 316.050 403.050 ;
        RECT 304.950 401.400 316.050 402.600 ;
        RECT 304.950 400.950 307.050 401.400 ;
        RECT 313.950 400.950 316.050 401.400 ;
        RECT 316.950 402.600 319.050 403.050 ;
        RECT 343.950 402.600 346.050 403.050 ;
        RECT 394.950 402.600 397.050 403.050 ;
        RECT 316.950 401.400 397.050 402.600 ;
        RECT 316.950 400.950 319.050 401.400 ;
        RECT 343.950 400.950 346.050 401.400 ;
        RECT 394.950 400.950 397.050 401.400 ;
        RECT 454.950 402.600 457.050 403.050 ;
        RECT 481.950 402.600 484.050 403.050 ;
        RECT 517.950 402.600 520.050 403.050 ;
        RECT 454.950 401.400 520.050 402.600 ;
        RECT 454.950 400.950 457.050 401.400 ;
        RECT 481.950 400.950 484.050 401.400 ;
        RECT 517.950 400.950 520.050 401.400 ;
        RECT 622.950 402.600 625.050 403.050 ;
        RECT 676.950 402.600 679.050 403.050 ;
        RECT 622.950 401.400 679.050 402.600 ;
        RECT 622.950 400.950 625.050 401.400 ;
        RECT 676.950 400.950 679.050 401.400 ;
        RECT 199.950 398.400 225.600 399.600 ;
        RECT 247.950 399.600 250.050 400.050 ;
        RECT 274.950 399.600 277.050 400.050 ;
        RECT 247.950 398.400 277.050 399.600 ;
        RECT 199.950 397.950 202.050 398.400 ;
        RECT 247.950 397.950 250.050 398.400 ;
        RECT 274.950 397.950 277.050 398.400 ;
        RECT 340.950 399.600 343.050 400.050 ;
        RECT 376.950 399.600 379.050 400.050 ;
        RECT 340.950 398.400 379.050 399.600 ;
        RECT 340.950 397.950 343.050 398.400 ;
        RECT 376.950 397.950 379.050 398.400 ;
        RECT 472.950 399.600 475.050 400.050 ;
        RECT 529.950 399.600 532.050 400.050 ;
        RECT 472.950 398.400 532.050 399.600 ;
        RECT 472.950 397.950 475.050 398.400 ;
        RECT 529.950 397.950 532.050 398.400 ;
        RECT 568.950 399.600 571.050 400.050 ;
        RECT 619.950 399.600 622.050 400.050 ;
        RECT 568.950 398.400 622.050 399.600 ;
        RECT 568.950 397.950 571.050 398.400 ;
        RECT 619.950 397.950 622.050 398.400 ;
        RECT 118.950 396.600 121.050 397.050 ;
        RECT 139.950 396.600 142.050 397.050 ;
        RECT 118.950 395.400 142.050 396.600 ;
        RECT 118.950 394.950 121.050 395.400 ;
        RECT 139.950 394.950 142.050 395.400 ;
        RECT 148.950 396.600 151.050 397.050 ;
        RECT 169.950 396.600 172.050 397.050 ;
        RECT 148.950 395.400 172.050 396.600 ;
        RECT 148.950 394.950 151.050 395.400 ;
        RECT 169.950 394.950 172.050 395.400 ;
        RECT 172.950 396.600 175.050 397.050 ;
        RECT 184.950 396.600 187.050 397.050 ;
        RECT 172.950 395.400 187.050 396.600 ;
        RECT 172.950 394.950 175.050 395.400 ;
        RECT 184.950 394.950 187.050 395.400 ;
        RECT 250.950 396.600 253.050 397.050 ;
        RECT 310.950 396.600 313.050 397.050 ;
        RECT 250.950 395.400 313.050 396.600 ;
        RECT 250.950 394.950 253.050 395.400 ;
        RECT 310.950 394.950 313.050 395.400 ;
        RECT 328.950 396.600 331.050 397.050 ;
        RECT 343.950 396.600 346.050 397.050 ;
        RECT 358.950 396.600 361.050 397.050 ;
        RECT 328.950 395.400 361.050 396.600 ;
        RECT 328.950 394.950 331.050 395.400 ;
        RECT 343.950 394.950 346.050 395.400 ;
        RECT 358.950 394.950 361.050 395.400 ;
        RECT 448.950 396.600 451.050 397.050 ;
        RECT 517.950 396.600 520.050 397.050 ;
        RECT 448.950 395.400 520.050 396.600 ;
        RECT 448.950 394.950 451.050 395.400 ;
        RECT 517.950 394.950 520.050 395.400 ;
        RECT 520.950 396.600 523.050 397.050 ;
        RECT 541.950 396.600 544.050 397.050 ;
        RECT 520.950 395.400 544.050 396.600 ;
        RECT 520.950 394.950 523.050 395.400 ;
        RECT 541.950 394.950 544.050 395.400 ;
        RECT 598.950 396.600 601.050 397.050 ;
        RECT 631.950 396.600 634.050 397.050 ;
        RECT 658.950 396.600 661.050 397.050 ;
        RECT 598.950 395.400 661.050 396.600 ;
        RECT 598.950 394.950 601.050 395.400 ;
        RECT 631.950 394.950 634.050 395.400 ;
        RECT 658.950 394.950 661.050 395.400 ;
        RECT 13.950 393.600 16.050 394.050 ;
        RECT 25.950 393.600 28.050 394.050 ;
        RECT 52.950 393.600 55.050 394.050 ;
        RECT 13.950 392.400 55.050 393.600 ;
        RECT 13.950 391.950 16.050 392.400 ;
        RECT 25.950 391.950 28.050 392.400 ;
        RECT 52.950 391.950 55.050 392.400 ;
        RECT 64.950 393.600 67.050 394.050 ;
        RECT 91.950 393.600 94.050 394.050 ;
        RECT 64.950 392.400 94.050 393.600 ;
        RECT 64.950 391.950 67.050 392.400 ;
        RECT 91.950 391.950 94.050 392.400 ;
        RECT 118.950 393.600 121.050 394.050 ;
        RECT 127.950 393.600 130.050 394.050 ;
        RECT 154.950 393.600 157.050 394.050 ;
        RECT 118.950 392.400 157.050 393.600 ;
        RECT 118.950 391.950 121.050 392.400 ;
        RECT 127.950 391.950 130.050 392.400 ;
        RECT 154.950 391.950 157.050 392.400 ;
        RECT 193.950 393.600 196.050 394.050 ;
        RECT 247.950 393.600 250.050 394.050 ;
        RECT 193.950 392.400 250.050 393.600 ;
        RECT 193.950 391.950 196.050 392.400 ;
        RECT 247.950 391.950 250.050 392.400 ;
        RECT 493.950 393.600 496.050 394.050 ;
        RECT 529.950 393.600 532.050 394.050 ;
        RECT 493.950 392.400 532.050 393.600 ;
        RECT 493.950 391.950 496.050 392.400 ;
        RECT 529.950 391.950 532.050 392.400 ;
        RECT 565.950 393.600 568.050 394.050 ;
        RECT 595.950 393.600 598.050 394.050 ;
        RECT 565.950 392.400 598.050 393.600 ;
        RECT 565.950 391.950 568.050 392.400 ;
        RECT 595.950 391.950 598.050 392.400 ;
        RECT 607.950 393.600 610.050 394.050 ;
        RECT 622.950 393.600 625.050 394.050 ;
        RECT 607.950 392.400 625.050 393.600 ;
        RECT 607.950 391.950 610.050 392.400 ;
        RECT 622.950 391.950 625.050 392.400 ;
        RECT 22.950 390.600 25.050 391.050 ;
        RECT 37.950 390.600 40.050 391.050 ;
        RECT 82.950 390.600 85.050 391.050 ;
        RECT 88.950 390.600 91.050 391.050 ;
        RECT 22.950 389.400 91.050 390.600 ;
        RECT 22.950 388.950 25.050 389.400 ;
        RECT 37.950 388.950 40.050 389.400 ;
        RECT 4.950 387.600 7.050 388.050 ;
        RECT 19.950 387.600 22.050 388.050 ;
        RECT 4.950 386.400 22.050 387.600 ;
        RECT 4.950 385.950 7.050 386.400 ;
        RECT 19.950 385.950 22.050 386.400 ;
        RECT 1.950 384.600 4.050 385.050 ;
        RECT 10.950 384.600 13.050 385.050 ;
        RECT 58.950 384.600 61.050 385.050 ;
        RECT 1.950 383.400 21.600 384.600 ;
        RECT 1.950 382.950 4.050 383.400 ;
        RECT 10.950 382.950 13.050 383.400 ;
        RECT 7.950 381.600 10.050 382.050 ;
        RECT 16.950 381.600 19.050 382.050 ;
        RECT 7.950 380.400 19.050 381.600 ;
        RECT 20.400 381.600 21.600 383.400 ;
        RECT 38.400 383.400 61.050 384.600 ;
        RECT 38.400 382.050 39.600 383.400 ;
        RECT 58.950 382.950 61.050 383.400 ;
        RECT 62.400 382.050 63.600 389.400 ;
        RECT 82.950 388.950 85.050 389.400 ;
        RECT 88.950 388.950 91.050 389.400 ;
        RECT 175.950 390.600 178.050 391.050 ;
        RECT 184.950 390.600 187.050 391.050 ;
        RECT 175.950 389.400 187.050 390.600 ;
        RECT 175.950 388.950 178.050 389.400 ;
        RECT 184.950 388.950 187.050 389.400 ;
        RECT 199.950 390.600 202.050 391.050 ;
        RECT 223.950 390.600 226.050 391.050 ;
        RECT 238.950 390.600 241.050 391.050 ;
        RECT 268.950 390.600 271.050 391.050 ;
        RECT 199.950 389.400 271.050 390.600 ;
        RECT 199.950 388.950 202.050 389.400 ;
        RECT 223.950 388.950 226.050 389.400 ;
        RECT 238.950 388.950 241.050 389.400 ;
        RECT 268.950 388.950 271.050 389.400 ;
        RECT 355.950 390.600 358.050 391.050 ;
        RECT 403.950 390.600 406.050 391.050 ;
        RECT 355.950 389.400 406.050 390.600 ;
        RECT 355.950 388.950 358.050 389.400 ;
        RECT 403.950 388.950 406.050 389.400 ;
        RECT 484.950 390.600 487.050 391.050 ;
        RECT 520.950 390.600 523.050 391.050 ;
        RECT 484.950 389.400 523.050 390.600 ;
        RECT 484.950 388.950 487.050 389.400 ;
        RECT 520.950 388.950 523.050 389.400 ;
        RECT 550.950 390.600 553.050 391.050 ;
        RECT 571.950 390.600 574.050 391.050 ;
        RECT 586.950 390.600 589.050 391.050 ;
        RECT 550.950 389.400 589.050 390.600 ;
        RECT 550.950 388.950 553.050 389.400 ;
        RECT 571.950 388.950 574.050 389.400 ;
        RECT 586.950 388.950 589.050 389.400 ;
        RECT 601.950 390.600 604.050 391.050 ;
        RECT 613.950 390.600 616.050 391.050 ;
        RECT 601.950 389.400 616.050 390.600 ;
        RECT 601.950 388.950 604.050 389.400 ;
        RECT 613.950 388.950 616.050 389.400 ;
        RECT 67.950 385.950 70.050 388.050 ;
        RECT 76.950 387.600 79.050 388.050 ;
        RECT 91.950 387.600 94.050 388.050 ;
        RECT 76.950 386.400 94.050 387.600 ;
        RECT 76.950 385.950 79.050 386.400 ;
        RECT 91.950 385.950 94.050 386.400 ;
        RECT 136.950 387.600 139.050 388.050 ;
        RECT 142.950 387.600 145.050 388.050 ;
        RECT 136.950 386.400 145.050 387.600 ;
        RECT 136.950 385.950 139.050 386.400 ;
        RECT 142.950 385.950 145.050 386.400 ;
        RECT 145.950 387.600 148.050 388.050 ;
        RECT 178.950 387.600 181.050 388.050 ;
        RECT 145.950 386.400 181.050 387.600 ;
        RECT 145.950 385.950 148.050 386.400 ;
        RECT 178.950 385.950 181.050 386.400 ;
        RECT 184.950 387.600 187.050 388.050 ;
        RECT 205.950 387.600 208.050 388.050 ;
        RECT 184.950 386.400 208.050 387.600 ;
        RECT 184.950 385.950 187.050 386.400 ;
        RECT 205.950 385.950 208.050 386.400 ;
        RECT 214.950 385.950 217.050 388.050 ;
        RECT 217.950 387.600 220.050 388.050 ;
        RECT 223.950 387.600 226.050 388.050 ;
        RECT 217.950 386.400 226.050 387.600 ;
        RECT 217.950 385.950 220.050 386.400 ;
        RECT 223.950 385.950 226.050 386.400 ;
        RECT 295.950 387.600 298.050 388.050 ;
        RECT 310.950 387.600 313.050 388.050 ;
        RECT 319.950 387.600 322.050 388.050 ;
        RECT 295.950 386.400 322.050 387.600 ;
        RECT 295.950 385.950 298.050 386.400 ;
        RECT 310.950 385.950 313.050 386.400 ;
        RECT 319.950 385.950 322.050 386.400 ;
        RECT 337.950 387.600 340.050 388.050 ;
        RECT 349.950 387.600 352.050 388.050 ;
        RECT 370.950 387.600 373.050 388.050 ;
        RECT 424.950 387.600 427.050 388.050 ;
        RECT 427.950 387.600 430.050 388.050 ;
        RECT 337.950 386.400 369.600 387.600 ;
        RECT 337.950 385.950 340.050 386.400 ;
        RECT 349.950 385.950 352.050 386.400 ;
        RECT 68.400 384.600 69.600 385.950 ;
        RECT 124.950 384.600 127.050 385.050 ;
        RECT 133.950 384.600 136.050 385.050 ;
        RECT 148.950 384.600 151.050 385.050 ;
        RECT 151.950 384.600 154.050 385.050 ;
        RECT 68.400 383.400 84.600 384.600 ;
        RECT 22.950 381.600 25.050 382.050 ;
        RECT 34.950 381.600 37.050 382.050 ;
        RECT 20.400 380.400 37.050 381.600 ;
        RECT 7.950 379.950 10.050 380.400 ;
        RECT 16.950 379.950 19.050 380.400 ;
        RECT 22.950 379.950 25.050 380.400 ;
        RECT 34.950 379.950 37.050 380.400 ;
        RECT 37.950 379.950 40.050 382.050 ;
        RECT 61.950 379.950 64.050 382.050 ;
        RECT 64.950 381.600 67.050 382.050 ;
        RECT 79.950 381.600 82.050 382.050 ;
        RECT 64.950 380.400 82.050 381.600 ;
        RECT 64.950 379.950 67.050 380.400 ;
        RECT 79.950 379.950 82.050 380.400 ;
        RECT 46.950 378.600 49.050 379.050 ;
        RECT 52.950 378.600 55.050 379.050 ;
        RECT 55.950 378.600 58.050 379.050 ;
        RECT 46.950 377.400 58.050 378.600 ;
        RECT 46.950 376.950 49.050 377.400 ;
        RECT 52.950 376.950 55.050 377.400 ;
        RECT 55.950 376.950 58.050 377.400 ;
        RECT 67.950 378.600 70.050 379.050 ;
        RECT 79.950 378.600 82.050 379.050 ;
        RECT 67.950 377.400 82.050 378.600 ;
        RECT 83.400 378.600 84.600 383.400 ;
        RECT 124.950 383.400 129.600 384.600 ;
        RECT 124.950 382.950 127.050 383.400 ;
        RECT 91.950 378.600 94.050 379.050 ;
        RECT 83.400 377.400 94.050 378.600 ;
        RECT 67.950 376.950 70.050 377.400 ;
        RECT 79.950 376.950 82.050 377.400 ;
        RECT 91.950 376.950 94.050 377.400 ;
        RECT 112.950 378.600 115.050 379.050 ;
        RECT 124.950 378.600 127.050 379.050 ;
        RECT 112.950 377.400 127.050 378.600 ;
        RECT 128.400 378.600 129.600 383.400 ;
        RECT 133.950 383.400 144.600 384.600 ;
        RECT 133.950 382.950 136.050 383.400 ;
        RECT 130.950 381.600 133.050 382.050 ;
        RECT 130.950 380.400 135.600 381.600 ;
        RECT 130.950 379.950 133.050 380.400 ;
        RECT 130.950 378.600 133.050 379.050 ;
        RECT 128.400 377.400 133.050 378.600 ;
        RECT 112.950 376.950 115.050 377.400 ;
        RECT 124.950 376.950 127.050 377.400 ;
        RECT 130.950 376.950 133.050 377.400 ;
        RECT 1.950 375.600 4.050 376.050 ;
        RECT 85.950 375.600 88.050 376.050 ;
        RECT 1.950 374.400 88.050 375.600 ;
        RECT 134.400 375.600 135.600 380.400 ;
        RECT 143.400 379.050 144.600 383.400 ;
        RECT 148.950 383.400 154.050 384.600 ;
        RECT 148.950 382.950 151.050 383.400 ;
        RECT 151.950 382.950 154.050 383.400 ;
        RECT 157.950 384.600 160.050 385.050 ;
        RECT 190.950 384.600 193.050 385.050 ;
        RECT 157.950 383.400 193.050 384.600 ;
        RECT 157.950 382.950 160.050 383.400 ;
        RECT 190.950 382.950 193.050 383.400 ;
        RECT 202.950 382.950 205.050 385.050 ;
        RECT 149.400 379.050 150.600 382.950 ;
        RECT 172.950 381.600 175.050 382.050 ;
        RECT 172.950 380.400 177.600 381.600 ;
        RECT 172.950 379.950 175.050 380.400 ;
        RECT 142.950 376.950 145.050 379.050 ;
        RECT 148.950 376.950 151.050 379.050 ;
        RECT 160.950 378.600 163.050 379.050 ;
        RECT 172.950 378.600 175.050 379.050 ;
        RECT 160.950 377.400 175.050 378.600 ;
        RECT 176.400 378.600 177.600 380.400 ;
        RECT 178.950 378.600 181.050 379.050 ;
        RECT 176.400 377.400 181.050 378.600 ;
        RECT 160.950 376.950 163.050 377.400 ;
        RECT 172.950 376.950 175.050 377.400 ;
        RECT 178.950 376.950 181.050 377.400 ;
        RECT 139.950 375.600 142.050 376.050 ;
        RECT 134.400 374.400 142.050 375.600 ;
        RECT 1.950 373.950 4.050 374.400 ;
        RECT 85.950 373.950 88.050 374.400 ;
        RECT 139.950 373.950 142.050 374.400 ;
        RECT 145.950 375.600 148.050 376.050 ;
        RECT 169.950 375.600 172.050 376.050 ;
        RECT 145.950 374.400 172.050 375.600 ;
        RECT 145.950 373.950 148.050 374.400 ;
        RECT 169.950 373.950 172.050 374.400 ;
        RECT 190.950 375.600 193.050 376.050 ;
        RECT 203.400 375.600 204.600 382.950 ;
        RECT 215.400 382.050 216.600 385.950 ;
        RECT 253.950 384.600 256.050 385.050 ;
        RECT 259.950 384.600 262.050 385.050 ;
        RECT 253.950 383.400 262.050 384.600 ;
        RECT 253.950 382.950 256.050 383.400 ;
        RECT 259.950 382.950 262.050 383.400 ;
        RECT 289.950 382.950 292.050 385.050 ;
        RECT 316.950 382.950 319.050 385.050 ;
        RECT 358.950 382.950 361.050 385.050 ;
        RECT 368.400 384.600 369.600 386.400 ;
        RECT 370.950 386.400 430.050 387.600 ;
        RECT 370.950 385.950 373.050 386.400 ;
        RECT 424.950 385.950 427.050 386.400 ;
        RECT 427.950 385.950 430.050 386.400 ;
        RECT 433.950 387.600 436.050 388.050 ;
        RECT 454.950 387.600 457.050 388.050 ;
        RECT 499.950 387.600 502.050 388.050 ;
        RECT 433.950 386.400 502.050 387.600 ;
        RECT 433.950 385.950 436.050 386.400 ;
        RECT 454.950 385.950 457.050 386.400 ;
        RECT 499.950 385.950 502.050 386.400 ;
        RECT 502.950 385.950 505.050 388.050 ;
        RECT 592.950 387.600 595.050 388.050 ;
        RECT 610.950 387.600 613.050 388.050 ;
        RECT 670.950 387.600 673.050 388.050 ;
        RECT 592.950 386.400 597.600 387.600 ;
        RECT 592.950 385.950 595.050 386.400 ;
        RECT 373.950 384.600 376.050 385.050 ;
        RECT 368.400 383.400 376.050 384.600 ;
        RECT 373.950 382.950 376.050 383.400 ;
        RECT 400.950 384.600 403.050 385.050 ;
        RECT 409.950 384.600 412.050 385.050 ;
        RECT 418.950 384.600 421.050 385.050 ;
        RECT 400.950 383.400 421.050 384.600 ;
        RECT 400.950 382.950 403.050 383.400 ;
        RECT 409.950 382.950 412.050 383.400 ;
        RECT 418.950 382.950 421.050 383.400 ;
        RECT 436.950 384.600 439.050 385.050 ;
        RECT 460.950 384.600 463.050 385.050 ;
        RECT 478.950 384.600 481.050 385.050 ;
        RECT 436.950 383.400 481.050 384.600 ;
        RECT 436.950 382.950 439.050 383.400 ;
        RECT 460.950 382.950 463.050 383.400 ;
        RECT 478.950 382.950 481.050 383.400 ;
        RECT 214.950 379.950 217.050 382.050 ;
        RECT 229.950 381.600 232.050 382.050 ;
        RECT 244.950 381.600 247.050 382.050 ;
        RECT 229.950 380.400 247.050 381.600 ;
        RECT 229.950 379.950 232.050 380.400 ;
        RECT 244.950 379.950 247.050 380.400 ;
        RECT 232.950 378.600 235.050 379.050 ;
        RECT 238.950 378.600 241.050 379.050 ;
        RECT 247.950 378.600 250.050 379.050 ;
        RECT 271.950 378.600 274.050 379.050 ;
        RECT 232.950 377.400 274.050 378.600 ;
        RECT 232.950 376.950 235.050 377.400 ;
        RECT 238.950 376.950 241.050 377.400 ;
        RECT 247.950 376.950 250.050 377.400 ;
        RECT 271.950 376.950 274.050 377.400 ;
        RECT 190.950 374.400 204.600 375.600 ;
        RECT 271.950 375.600 274.050 376.050 ;
        RECT 283.950 375.600 286.050 376.050 ;
        RECT 271.950 374.400 286.050 375.600 ;
        RECT 290.400 375.600 291.600 382.950 ;
        RECT 301.950 381.600 304.050 382.050 ;
        RECT 313.950 381.600 316.050 382.050 ;
        RECT 317.400 381.600 318.600 382.950 ;
        RECT 301.950 380.400 318.600 381.600 ;
        RECT 325.950 381.600 328.050 382.050 ;
        RECT 328.950 381.600 331.050 382.050 ;
        RECT 331.950 381.600 334.050 382.050 ;
        RECT 325.950 380.400 334.050 381.600 ;
        RECT 301.950 379.950 304.050 380.400 ;
        RECT 313.950 379.950 316.050 380.400 ;
        RECT 325.950 379.950 328.050 380.400 ;
        RECT 328.950 379.950 331.050 380.400 ;
        RECT 331.950 379.950 334.050 380.400 ;
        RECT 346.950 381.600 349.050 382.050 ;
        RECT 355.950 381.600 358.050 382.050 ;
        RECT 346.950 380.400 358.050 381.600 ;
        RECT 346.950 379.950 349.050 380.400 ;
        RECT 355.950 379.950 358.050 380.400 ;
        RECT 298.950 378.600 301.050 379.050 ;
        RECT 307.950 378.600 310.050 379.050 ;
        RECT 298.950 377.400 310.050 378.600 ;
        RECT 298.950 376.950 301.050 377.400 ;
        RECT 307.950 376.950 310.050 377.400 ;
        RECT 349.950 378.600 352.050 379.050 ;
        RECT 359.400 378.600 360.600 382.950 ;
        RECT 361.950 381.600 364.050 382.050 ;
        RECT 403.950 381.600 406.050 382.050 ;
        RECT 361.950 380.400 406.050 381.600 ;
        RECT 361.950 379.950 364.050 380.400 ;
        RECT 403.950 379.950 406.050 380.400 ;
        RECT 415.950 381.600 418.050 382.050 ;
        RECT 439.950 381.600 442.050 382.050 ;
        RECT 463.950 381.600 466.050 382.050 ;
        RECT 415.950 380.400 438.600 381.600 ;
        RECT 415.950 379.950 418.050 380.400 ;
        RECT 437.400 379.050 438.600 380.400 ;
        RECT 439.950 380.400 466.050 381.600 ;
        RECT 439.950 379.950 442.050 380.400 ;
        RECT 463.950 379.950 466.050 380.400 ;
        RECT 469.950 381.600 472.050 382.050 ;
        RECT 493.950 381.600 496.050 382.050 ;
        RECT 469.950 380.400 496.050 381.600 ;
        RECT 503.400 381.600 504.600 385.950 ;
        RECT 520.950 384.600 523.050 385.050 ;
        RECT 538.950 384.600 541.050 385.050 ;
        RECT 520.950 383.400 541.050 384.600 ;
        RECT 520.950 382.950 523.050 383.400 ;
        RECT 538.950 382.950 541.050 383.400 ;
        RECT 553.950 384.600 556.050 385.050 ;
        RECT 580.950 384.600 583.050 385.050 ;
        RECT 553.950 383.400 583.050 384.600 ;
        RECT 553.950 382.950 556.050 383.400 ;
        RECT 580.950 382.950 583.050 383.400 ;
        RECT 592.950 382.950 595.050 385.050 ;
        RECT 508.950 381.600 511.050 382.050 ;
        RECT 503.400 380.400 511.050 381.600 ;
        RECT 469.950 379.950 472.050 380.400 ;
        RECT 493.950 379.950 496.050 380.400 ;
        RECT 508.950 379.950 511.050 380.400 ;
        RECT 565.950 381.600 568.050 382.050 ;
        RECT 583.950 381.600 586.050 382.050 ;
        RECT 565.950 380.400 586.050 381.600 ;
        RECT 565.950 379.950 568.050 380.400 ;
        RECT 583.950 379.950 586.050 380.400 ;
        RECT 589.950 381.600 592.050 382.050 ;
        RECT 593.400 381.600 594.600 382.950 ;
        RECT 596.400 382.050 597.600 386.400 ;
        RECT 610.950 386.400 673.050 387.600 ;
        RECT 610.950 385.950 613.050 386.400 ;
        RECT 670.950 385.950 673.050 386.400 ;
        RECT 598.950 384.600 601.050 385.050 ;
        RECT 604.950 384.600 607.050 385.050 ;
        RECT 598.950 383.400 607.050 384.600 ;
        RECT 598.950 382.950 601.050 383.400 ;
        RECT 604.950 382.950 607.050 383.400 ;
        RECT 646.950 384.600 649.050 385.050 ;
        RECT 676.950 384.600 679.050 385.050 ;
        RECT 646.950 383.400 679.050 384.600 ;
        RECT 646.950 382.950 649.050 383.400 ;
        RECT 676.950 382.950 679.050 383.400 ;
        RECT 679.950 384.600 682.050 385.050 ;
        RECT 688.950 384.600 691.050 385.050 ;
        RECT 679.950 383.400 691.050 384.600 ;
        RECT 679.950 382.950 682.050 383.400 ;
        RECT 688.950 382.950 691.050 383.400 ;
        RECT 691.950 382.950 694.050 385.050 ;
        RECT 589.950 380.400 594.600 381.600 ;
        RECT 589.950 379.950 592.050 380.400 ;
        RECT 595.950 379.950 598.050 382.050 ;
        RECT 628.950 381.600 631.050 382.050 ;
        RECT 631.950 381.600 634.050 382.050 ;
        RECT 649.950 381.600 652.050 382.050 ;
        RECT 628.950 380.400 652.050 381.600 ;
        RECT 628.950 379.950 631.050 380.400 ;
        RECT 631.950 379.950 634.050 380.400 ;
        RECT 649.950 379.950 652.050 380.400 ;
        RECT 664.950 381.600 667.050 382.050 ;
        RECT 664.950 380.400 687.600 381.600 ;
        RECT 664.950 379.950 667.050 380.400 ;
        RECT 686.400 379.050 687.600 380.400 ;
        RECT 692.400 379.050 693.600 382.950 ;
        RECT 349.950 377.400 360.600 378.600 ;
        RECT 385.950 378.600 388.050 379.050 ;
        RECT 418.950 378.600 421.050 379.050 ;
        RECT 427.950 378.600 430.050 379.050 ;
        RECT 385.950 377.400 430.050 378.600 ;
        RECT 349.950 376.950 352.050 377.400 ;
        RECT 385.950 376.950 388.050 377.400 ;
        RECT 418.950 376.950 421.050 377.400 ;
        RECT 427.950 376.950 430.050 377.400 ;
        RECT 436.950 376.950 439.050 379.050 ;
        RECT 496.950 378.600 499.050 379.050 ;
        RECT 508.950 378.600 511.050 379.050 ;
        RECT 496.950 377.400 511.050 378.600 ;
        RECT 496.950 376.950 499.050 377.400 ;
        RECT 508.950 376.950 511.050 377.400 ;
        RECT 637.950 378.600 640.050 379.050 ;
        RECT 646.950 378.600 649.050 379.050 ;
        RECT 637.950 377.400 649.050 378.600 ;
        RECT 637.950 376.950 640.050 377.400 ;
        RECT 646.950 376.950 649.050 377.400 ;
        RECT 664.950 378.600 667.050 379.050 ;
        RECT 682.950 378.600 685.050 379.050 ;
        RECT 664.950 377.400 685.050 378.600 ;
        RECT 664.950 376.950 667.050 377.400 ;
        RECT 682.950 376.950 685.050 377.400 ;
        RECT 685.950 376.950 688.050 379.050 ;
        RECT 691.950 376.950 694.050 379.050 ;
        RECT 694.950 378.600 697.050 379.050 ;
        RECT 703.950 378.600 706.050 379.050 ;
        RECT 694.950 377.400 706.050 378.600 ;
        RECT 694.950 376.950 697.050 377.400 ;
        RECT 703.950 376.950 706.050 377.400 ;
        RECT 304.950 375.600 307.050 376.050 ;
        RECT 290.400 374.400 307.050 375.600 ;
        RECT 190.950 373.950 193.050 374.400 ;
        RECT 271.950 373.950 274.050 374.400 ;
        RECT 283.950 373.950 286.050 374.400 ;
        RECT 304.950 373.950 307.050 374.400 ;
        RECT 382.950 375.600 385.050 376.050 ;
        RECT 385.950 375.600 388.050 376.050 ;
        RECT 397.950 375.600 400.050 376.050 ;
        RECT 382.950 374.400 400.050 375.600 ;
        RECT 382.950 373.950 385.050 374.400 ;
        RECT 385.950 373.950 388.050 374.400 ;
        RECT 397.950 373.950 400.050 374.400 ;
        RECT 406.950 375.600 409.050 376.050 ;
        RECT 421.950 375.600 424.050 376.050 ;
        RECT 406.950 374.400 424.050 375.600 ;
        RECT 406.950 373.950 409.050 374.400 ;
        RECT 421.950 373.950 424.050 374.400 ;
        RECT 430.950 375.600 433.050 376.050 ;
        RECT 442.950 375.600 445.050 376.050 ;
        RECT 430.950 374.400 445.050 375.600 ;
        RECT 430.950 373.950 433.050 374.400 ;
        RECT 442.950 373.950 445.050 374.400 ;
        RECT 490.950 375.600 493.050 376.050 ;
        RECT 532.950 375.600 535.050 376.050 ;
        RECT 535.950 375.600 538.050 376.050 ;
        RECT 490.950 374.400 538.050 375.600 ;
        RECT 490.950 373.950 493.050 374.400 ;
        RECT 532.950 373.950 535.050 374.400 ;
        RECT 535.950 373.950 538.050 374.400 ;
        RECT 571.950 375.600 574.050 376.050 ;
        RECT 604.950 375.600 607.050 376.050 ;
        RECT 613.950 375.600 616.050 376.050 ;
        RECT 571.950 374.400 616.050 375.600 ;
        RECT 571.950 373.950 574.050 374.400 ;
        RECT 604.950 373.950 607.050 374.400 ;
        RECT 613.950 373.950 616.050 374.400 ;
        RECT 667.950 375.600 670.050 376.050 ;
        RECT 697.950 375.600 700.050 376.050 ;
        RECT 667.950 374.400 700.050 375.600 ;
        RECT 667.950 373.950 670.050 374.400 ;
        RECT 697.950 373.950 700.050 374.400 ;
        RECT 70.950 372.600 73.050 373.050 ;
        RECT 88.950 372.600 91.050 373.050 ;
        RECT 70.950 371.400 91.050 372.600 ;
        RECT 70.950 370.950 73.050 371.400 ;
        RECT 88.950 370.950 91.050 371.400 ;
        RECT 106.950 372.600 109.050 373.050 ;
        RECT 121.950 372.600 124.050 373.050 ;
        RECT 124.950 372.600 127.050 373.050 ;
        RECT 106.950 371.400 127.050 372.600 ;
        RECT 106.950 370.950 109.050 371.400 ;
        RECT 121.950 370.950 124.050 371.400 ;
        RECT 124.950 370.950 127.050 371.400 ;
        RECT 142.950 372.600 145.050 373.050 ;
        RECT 151.950 372.600 154.050 373.050 ;
        RECT 142.950 371.400 154.050 372.600 ;
        RECT 142.950 370.950 145.050 371.400 ;
        RECT 151.950 370.950 154.050 371.400 ;
        RECT 202.950 372.600 205.050 373.050 ;
        RECT 211.950 372.600 214.050 373.050 ;
        RECT 250.950 372.600 253.050 373.050 ;
        RECT 202.950 371.400 253.050 372.600 ;
        RECT 202.950 370.950 205.050 371.400 ;
        RECT 211.950 370.950 214.050 371.400 ;
        RECT 250.950 370.950 253.050 371.400 ;
        RECT 268.950 372.600 271.050 373.050 ;
        RECT 277.950 372.600 280.050 373.050 ;
        RECT 268.950 371.400 280.050 372.600 ;
        RECT 268.950 370.950 271.050 371.400 ;
        RECT 277.950 370.950 280.050 371.400 ;
        RECT 292.950 372.600 295.050 373.050 ;
        RECT 304.950 372.600 307.050 373.050 ;
        RECT 292.950 371.400 307.050 372.600 ;
        RECT 292.950 370.950 295.050 371.400 ;
        RECT 304.950 370.950 307.050 371.400 ;
        RECT 577.950 372.600 580.050 373.050 ;
        RECT 589.950 372.600 592.050 373.050 ;
        RECT 577.950 371.400 592.050 372.600 ;
        RECT 577.950 370.950 580.050 371.400 ;
        RECT 589.950 370.950 592.050 371.400 ;
        RECT 592.950 372.600 595.050 373.050 ;
        RECT 634.950 372.600 637.050 373.050 ;
        RECT 592.950 371.400 637.050 372.600 ;
        RECT 592.950 370.950 595.050 371.400 ;
        RECT 634.950 370.950 637.050 371.400 ;
        RECT 673.950 372.600 676.050 373.050 ;
        RECT 691.950 372.600 694.050 373.050 ;
        RECT 703.950 372.600 706.050 373.050 ;
        RECT 673.950 371.400 706.050 372.600 ;
        RECT 673.950 370.950 676.050 371.400 ;
        RECT 691.950 370.950 694.050 371.400 ;
        RECT 703.950 370.950 706.050 371.400 ;
        RECT 49.950 369.600 52.050 370.050 ;
        RECT 115.950 369.600 118.050 370.050 ;
        RECT 49.950 368.400 118.050 369.600 ;
        RECT 49.950 367.950 52.050 368.400 ;
        RECT 115.950 367.950 118.050 368.400 ;
        RECT 136.950 369.600 139.050 370.050 ;
        RECT 166.950 369.600 169.050 370.050 ;
        RECT 136.950 368.400 169.050 369.600 ;
        RECT 136.950 367.950 139.050 368.400 ;
        RECT 166.950 367.950 169.050 368.400 ;
        RECT 271.950 369.600 274.050 370.050 ;
        RECT 313.950 369.600 316.050 370.050 ;
        RECT 271.950 368.400 316.050 369.600 ;
        RECT 271.950 367.950 274.050 368.400 ;
        RECT 313.950 367.950 316.050 368.400 ;
        RECT 487.950 369.600 490.050 370.050 ;
        RECT 610.950 369.600 613.050 370.050 ;
        RECT 487.950 368.400 613.050 369.600 ;
        RECT 487.950 367.950 490.050 368.400 ;
        RECT 610.950 367.950 613.050 368.400 ;
        RECT 145.950 366.600 148.050 367.050 ;
        RECT 160.950 366.600 163.050 367.050 ;
        RECT 145.950 365.400 163.050 366.600 ;
        RECT 145.950 364.950 148.050 365.400 ;
        RECT 160.950 364.950 163.050 365.400 ;
        RECT 607.950 366.600 610.050 367.050 ;
        RECT 616.950 366.600 619.050 367.050 ;
        RECT 607.950 365.400 619.050 366.600 ;
        RECT 607.950 364.950 610.050 365.400 ;
        RECT 616.950 364.950 619.050 365.400 ;
        RECT 61.950 363.600 64.050 364.050 ;
        RECT 73.950 363.600 76.050 364.050 ;
        RECT 61.950 362.400 76.050 363.600 ;
        RECT 61.950 361.950 64.050 362.400 ;
        RECT 73.950 361.950 76.050 362.400 ;
        RECT 85.950 363.600 88.050 364.050 ;
        RECT 214.950 363.600 217.050 364.050 ;
        RECT 85.950 362.400 217.050 363.600 ;
        RECT 85.950 361.950 88.050 362.400 ;
        RECT 214.950 361.950 217.050 362.400 ;
        RECT 265.950 363.600 268.050 364.050 ;
        RECT 289.950 363.600 292.050 364.050 ;
        RECT 322.950 363.600 325.050 364.050 ;
        RECT 265.950 362.400 325.050 363.600 ;
        RECT 265.950 361.950 268.050 362.400 ;
        RECT 289.950 361.950 292.050 362.400 ;
        RECT 322.950 361.950 325.050 362.400 ;
        RECT 436.950 363.600 439.050 364.050 ;
        RECT 445.950 363.600 448.050 364.050 ;
        RECT 436.950 362.400 448.050 363.600 ;
        RECT 436.950 361.950 439.050 362.400 ;
        RECT 445.950 361.950 448.050 362.400 ;
        RECT 4.950 360.600 7.050 361.050 ;
        RECT 31.950 360.600 34.050 361.050 ;
        RECT 4.950 359.400 34.050 360.600 ;
        RECT 4.950 358.950 7.050 359.400 ;
        RECT 31.950 358.950 34.050 359.400 ;
        RECT 112.950 360.600 115.050 361.050 ;
        RECT 121.950 360.600 124.050 361.050 ;
        RECT 130.950 360.600 133.050 361.050 ;
        RECT 112.950 359.400 133.050 360.600 ;
        RECT 112.950 358.950 115.050 359.400 ;
        RECT 121.950 358.950 124.050 359.400 ;
        RECT 130.950 358.950 133.050 359.400 ;
        RECT 154.950 360.600 157.050 361.050 ;
        RECT 187.950 360.600 190.050 361.050 ;
        RECT 154.950 359.400 190.050 360.600 ;
        RECT 154.950 358.950 157.050 359.400 ;
        RECT 187.950 358.950 190.050 359.400 ;
        RECT 565.950 360.600 568.050 361.050 ;
        RECT 601.950 360.600 604.050 361.050 ;
        RECT 565.950 359.400 604.050 360.600 ;
        RECT 565.950 358.950 568.050 359.400 ;
        RECT 601.950 358.950 604.050 359.400 ;
        RECT 100.950 357.600 103.050 358.050 ;
        RECT 148.950 357.600 151.050 358.050 ;
        RECT 172.950 357.600 175.050 358.050 ;
        RECT 100.950 356.400 175.050 357.600 ;
        RECT 100.950 355.950 103.050 356.400 ;
        RECT 148.950 355.950 151.050 356.400 ;
        RECT 172.950 355.950 175.050 356.400 ;
        RECT 223.950 357.600 226.050 358.050 ;
        RECT 244.950 357.600 247.050 358.050 ;
        RECT 223.950 356.400 247.050 357.600 ;
        RECT 223.950 355.950 226.050 356.400 ;
        RECT 244.950 355.950 247.050 356.400 ;
        RECT 571.950 357.600 574.050 358.050 ;
        RECT 598.950 357.600 601.050 358.050 ;
        RECT 571.950 356.400 601.050 357.600 ;
        RECT 571.950 355.950 574.050 356.400 ;
        RECT 598.950 355.950 601.050 356.400 ;
        RECT 19.950 354.600 22.050 355.050 ;
        RECT 40.950 354.600 43.050 355.050 ;
        RECT 19.950 353.400 43.050 354.600 ;
        RECT 19.950 352.950 22.050 353.400 ;
        RECT 40.950 352.950 43.050 353.400 ;
        RECT 46.950 354.600 49.050 355.050 ;
        RECT 67.950 354.600 70.050 355.050 ;
        RECT 46.950 353.400 70.050 354.600 ;
        RECT 46.950 352.950 49.050 353.400 ;
        RECT 67.950 352.950 70.050 353.400 ;
        RECT 112.950 354.600 115.050 355.050 ;
        RECT 220.950 354.600 223.050 355.050 ;
        RECT 112.950 353.400 223.050 354.600 ;
        RECT 112.950 352.950 115.050 353.400 ;
        RECT 220.950 352.950 223.050 353.400 ;
        RECT 337.950 354.600 340.050 355.050 ;
        RECT 394.950 354.600 397.050 355.050 ;
        RECT 337.950 353.400 397.050 354.600 ;
        RECT 337.950 352.950 340.050 353.400 ;
        RECT 394.950 352.950 397.050 353.400 ;
        RECT 463.950 354.600 466.050 355.050 ;
        RECT 529.950 354.600 532.050 355.050 ;
        RECT 463.950 353.400 532.050 354.600 ;
        RECT 463.950 352.950 466.050 353.400 ;
        RECT 529.950 352.950 532.050 353.400 ;
        RECT 535.950 354.600 538.050 355.050 ;
        RECT 550.950 354.600 553.050 355.050 ;
        RECT 535.950 353.400 553.050 354.600 ;
        RECT 535.950 352.950 538.050 353.400 ;
        RECT 550.950 352.950 553.050 353.400 ;
        RECT 553.950 354.600 556.050 355.050 ;
        RECT 580.950 354.600 583.050 355.050 ;
        RECT 553.950 353.400 583.050 354.600 ;
        RECT 553.950 352.950 556.050 353.400 ;
        RECT 580.950 352.950 583.050 353.400 ;
        RECT 61.950 351.600 64.050 352.050 ;
        RECT 11.400 350.400 64.050 351.600 ;
        RECT 1.950 346.950 4.050 349.050 ;
        RECT 4.950 346.950 7.050 349.050 ;
        RECT 2.400 333.600 3.600 346.950 ;
        RECT 5.400 340.050 6.600 346.950 ;
        RECT 7.950 342.600 10.050 343.050 ;
        RECT 11.400 342.600 12.600 350.400 ;
        RECT 13.950 346.950 16.050 349.050 ;
        RECT 46.950 346.950 49.050 349.050 ;
        RECT 14.400 343.050 15.600 346.950 ;
        RECT 28.950 345.600 31.050 346.050 ;
        RECT 43.950 345.600 46.050 346.050 ;
        RECT 28.950 344.400 46.050 345.600 ;
        RECT 28.950 343.950 31.050 344.400 ;
        RECT 43.950 343.950 46.050 344.400 ;
        RECT 47.400 343.050 48.600 346.950 ;
        RECT 7.950 341.400 12.600 342.600 ;
        RECT 13.950 342.600 16.050 343.050 ;
        RECT 25.950 342.600 28.050 343.050 ;
        RECT 34.950 342.600 37.050 343.050 ;
        RECT 13.950 341.400 24.600 342.600 ;
        RECT 7.950 340.950 10.050 341.400 ;
        RECT 13.950 340.950 16.050 341.400 ;
        RECT 4.950 337.950 7.050 340.050 ;
        RECT 10.950 339.600 13.050 340.050 ;
        RECT 19.950 339.600 22.050 340.050 ;
        RECT 10.950 338.400 22.050 339.600 ;
        RECT 23.400 339.600 24.600 341.400 ;
        RECT 25.950 341.400 37.050 342.600 ;
        RECT 25.950 340.950 28.050 341.400 ;
        RECT 34.950 340.950 37.050 341.400 ;
        RECT 40.950 342.600 43.050 343.050 ;
        RECT 46.950 342.600 49.050 343.050 ;
        RECT 40.950 341.400 49.050 342.600 ;
        RECT 50.400 342.600 51.600 350.400 ;
        RECT 61.950 349.950 64.050 350.400 ;
        RECT 142.950 351.600 145.050 352.050 ;
        RECT 178.950 351.600 181.050 352.050 ;
        RECT 142.950 350.400 181.050 351.600 ;
        RECT 142.950 349.950 145.050 350.400 ;
        RECT 178.950 349.950 181.050 350.400 ;
        RECT 196.950 351.600 199.050 352.050 ;
        RECT 202.950 351.600 205.050 352.050 ;
        RECT 196.950 350.400 205.050 351.600 ;
        RECT 196.950 349.950 199.050 350.400 ;
        RECT 202.950 349.950 205.050 350.400 ;
        RECT 376.950 351.600 379.050 352.050 ;
        RECT 400.950 351.600 403.050 352.050 ;
        RECT 619.950 351.600 622.050 352.050 ;
        RECT 376.950 350.400 403.050 351.600 ;
        RECT 376.950 349.950 379.050 350.400 ;
        RECT 400.950 349.950 403.050 350.400 ;
        RECT 593.400 350.400 622.050 351.600 ;
        RECT 52.950 346.950 55.050 349.050 ;
        RECT 76.950 348.600 79.050 349.050 ;
        RECT 94.950 348.600 97.050 349.050 ;
        RECT 76.950 347.400 97.050 348.600 ;
        RECT 76.950 346.950 79.050 347.400 ;
        RECT 94.950 346.950 97.050 347.400 ;
        RECT 166.950 348.600 169.050 349.050 ;
        RECT 169.950 348.600 172.050 349.050 ;
        RECT 196.950 348.600 199.050 349.050 ;
        RECT 166.950 347.400 199.050 348.600 ;
        RECT 166.950 346.950 169.050 347.400 ;
        RECT 169.950 346.950 172.050 347.400 ;
        RECT 196.950 346.950 199.050 347.400 ;
        RECT 340.950 348.600 343.050 349.050 ;
        RECT 391.950 348.600 394.050 349.050 ;
        RECT 340.950 347.400 394.050 348.600 ;
        RECT 340.950 346.950 343.050 347.400 ;
        RECT 53.400 345.600 54.600 346.950 ;
        RECT 97.950 345.600 100.050 346.050 ;
        RECT 109.950 345.600 112.050 346.050 ;
        RECT 136.950 345.600 139.050 346.050 ;
        RECT 53.400 344.400 57.600 345.600 ;
        RECT 52.950 342.600 55.050 343.050 ;
        RECT 50.400 341.400 55.050 342.600 ;
        RECT 40.950 340.950 43.050 341.400 ;
        RECT 46.950 340.950 49.050 341.400 ;
        RECT 52.950 340.950 55.050 341.400 ;
        RECT 56.400 340.050 57.600 344.400 ;
        RECT 97.950 344.400 112.050 345.600 ;
        RECT 97.950 343.950 100.050 344.400 ;
        RECT 109.950 343.950 112.050 344.400 ;
        RECT 128.400 344.400 139.050 345.600 ;
        RECT 64.950 340.950 67.050 343.050 ;
        RECT 79.950 340.950 82.050 343.050 ;
        RECT 103.950 340.950 106.050 343.050 ;
        RECT 49.950 339.600 52.050 340.050 ;
        RECT 23.400 338.400 52.050 339.600 ;
        RECT 10.950 337.950 13.050 338.400 ;
        RECT 19.950 337.950 22.050 338.400 ;
        RECT 49.950 337.950 52.050 338.400 ;
        RECT 55.950 337.950 58.050 340.050 ;
        RECT 65.400 339.600 66.600 340.950 ;
        RECT 70.950 339.600 73.050 340.050 ;
        RECT 80.400 339.600 81.600 340.950 ;
        RECT 65.400 338.400 69.600 339.600 ;
        RECT 28.950 336.600 31.050 337.050 ;
        RECT 31.950 336.600 34.050 337.050 ;
        RECT 43.950 336.600 46.050 337.050 ;
        RECT 28.950 335.400 46.050 336.600 ;
        RECT 28.950 334.950 31.050 335.400 ;
        RECT 31.950 334.950 34.050 335.400 ;
        RECT 43.950 334.950 46.050 335.400 ;
        RECT 49.950 336.600 52.050 337.050 ;
        RECT 64.950 336.600 67.050 337.050 ;
        RECT 49.950 335.400 67.050 336.600 ;
        RECT 68.400 336.600 69.600 338.400 ;
        RECT 70.950 338.400 81.600 339.600 ;
        RECT 82.950 339.600 85.050 340.050 ;
        RECT 88.950 339.600 91.050 340.050 ;
        RECT 82.950 338.400 91.050 339.600 ;
        RECT 104.400 339.600 105.600 340.950 ;
        RECT 128.400 340.050 129.600 344.400 ;
        RECT 136.950 343.950 139.050 344.400 ;
        RECT 142.950 343.950 145.050 346.050 ;
        RECT 295.950 345.600 298.050 346.050 ;
        RECT 310.950 345.600 313.050 346.050 ;
        RECT 295.950 344.400 313.050 345.600 ;
        RECT 295.950 343.950 298.050 344.400 ;
        RECT 310.950 343.950 313.050 344.400 ;
        RECT 352.950 345.600 355.050 346.050 ;
        RECT 358.950 345.600 361.050 346.050 ;
        RECT 352.950 344.400 361.050 345.600 ;
        RECT 352.950 343.950 355.050 344.400 ;
        RECT 358.950 343.950 361.050 344.400 ;
        RECT 376.950 345.600 379.050 346.050 ;
        RECT 380.400 345.600 381.600 347.400 ;
        RECT 391.950 346.950 394.050 347.400 ;
        RECT 493.950 348.600 496.050 349.050 ;
        RECT 544.950 348.600 547.050 349.050 ;
        RECT 493.950 347.400 547.050 348.600 ;
        RECT 493.950 346.950 496.050 347.400 ;
        RECT 544.950 346.950 547.050 347.400 ;
        RECT 547.950 348.600 550.050 349.050 ;
        RECT 556.950 348.600 559.050 349.050 ;
        RECT 547.950 347.400 559.050 348.600 ;
        RECT 547.950 346.950 550.050 347.400 ;
        RECT 556.950 346.950 559.050 347.400 ;
        RECT 376.950 344.400 381.600 345.600 ;
        RECT 382.950 345.600 385.050 346.050 ;
        RECT 391.950 345.600 394.050 346.050 ;
        RECT 382.950 344.400 394.050 345.600 ;
        RECT 376.950 343.950 379.050 344.400 ;
        RECT 382.950 343.950 385.050 344.400 ;
        RECT 391.950 343.950 394.050 344.400 ;
        RECT 448.950 345.600 451.050 346.050 ;
        RECT 472.950 345.600 475.050 346.050 ;
        RECT 448.950 344.400 475.050 345.600 ;
        RECT 448.950 343.950 451.050 344.400 ;
        RECT 472.950 343.950 475.050 344.400 ;
        RECT 532.950 345.600 535.050 346.050 ;
        RECT 565.950 345.600 568.050 346.050 ;
        RECT 532.950 344.400 568.050 345.600 ;
        RECT 532.950 343.950 535.050 344.400 ;
        RECT 565.950 343.950 568.050 344.400 ;
        RECT 571.950 343.950 574.050 346.050 ;
        RECT 589.950 343.950 592.050 346.050 ;
        RECT 143.400 340.050 144.600 343.950 ;
        RECT 154.950 342.600 157.050 343.050 ;
        RECT 175.950 342.600 178.050 343.050 ;
        RECT 154.950 341.400 178.050 342.600 ;
        RECT 154.950 340.950 157.050 341.400 ;
        RECT 175.950 340.950 178.050 341.400 ;
        RECT 181.950 340.950 184.050 343.050 ;
        RECT 232.950 342.600 235.050 343.050 ;
        RECT 241.950 342.600 244.050 343.050 ;
        RECT 232.950 341.400 244.050 342.600 ;
        RECT 232.950 340.950 235.050 341.400 ;
        RECT 241.950 340.950 244.050 341.400 ;
        RECT 286.950 342.600 289.050 343.050 ;
        RECT 295.950 342.600 298.050 343.050 ;
        RECT 286.950 341.400 298.050 342.600 ;
        RECT 286.950 340.950 289.050 341.400 ;
        RECT 295.950 340.950 298.050 341.400 ;
        RECT 301.950 342.600 304.050 343.050 ;
        RECT 331.950 342.600 334.050 343.050 ;
        RECT 301.950 341.400 334.050 342.600 ;
        RECT 301.950 340.950 304.050 341.400 ;
        RECT 331.950 340.950 334.050 341.400 ;
        RECT 337.950 342.600 340.050 343.050 ;
        RECT 355.950 342.600 358.050 343.050 ;
        RECT 364.950 342.600 367.050 343.050 ;
        RECT 337.950 341.400 348.600 342.600 ;
        RECT 337.950 340.950 340.050 341.400 ;
        RECT 118.950 339.600 121.050 340.050 ;
        RECT 104.400 338.400 121.050 339.600 ;
        RECT 70.950 337.950 73.050 338.400 ;
        RECT 82.950 337.950 85.050 338.400 ;
        RECT 88.950 337.950 91.050 338.400 ;
        RECT 118.950 337.950 121.050 338.400 ;
        RECT 127.950 337.950 130.050 340.050 ;
        RECT 136.950 339.600 139.050 340.050 ;
        RECT 142.950 339.600 145.050 340.050 ;
        RECT 136.950 338.400 145.050 339.600 ;
        RECT 136.950 337.950 139.050 338.400 ;
        RECT 142.950 337.950 145.050 338.400 ;
        RECT 151.950 339.600 154.050 340.050 ;
        RECT 157.950 339.600 160.050 340.050 ;
        RECT 160.950 339.600 163.050 340.050 ;
        RECT 151.950 338.400 163.050 339.600 ;
        RECT 151.950 337.950 154.050 338.400 ;
        RECT 157.950 337.950 160.050 338.400 ;
        RECT 160.950 337.950 163.050 338.400 ;
        RECT 175.950 339.600 178.050 340.050 ;
        RECT 182.400 339.600 183.600 340.950 ;
        RECT 347.400 340.050 348.600 341.400 ;
        RECT 355.950 341.400 367.050 342.600 ;
        RECT 355.950 340.950 358.050 341.400 ;
        RECT 364.950 340.950 367.050 341.400 ;
        RECT 370.950 342.600 373.050 343.050 ;
        RECT 379.950 342.600 382.050 343.050 ;
        RECT 370.950 341.400 382.050 342.600 ;
        RECT 370.950 340.950 373.050 341.400 ;
        RECT 379.950 340.950 382.050 341.400 ;
        RECT 427.950 342.600 430.050 343.050 ;
        RECT 523.950 342.600 526.050 343.050 ;
        RECT 541.950 342.600 544.050 343.050 ;
        RECT 427.950 341.400 462.600 342.600 ;
        RECT 427.950 340.950 430.050 341.400 ;
        RECT 175.950 338.400 183.600 339.600 ;
        RECT 184.950 339.600 187.050 340.050 ;
        RECT 211.950 339.600 214.050 340.050 ;
        RECT 217.950 339.600 220.050 340.050 ;
        RECT 184.950 338.400 207.600 339.600 ;
        RECT 175.950 337.950 178.050 338.400 ;
        RECT 184.950 337.950 187.050 338.400 ;
        RECT 70.950 336.600 73.050 337.050 ;
        RECT 68.400 335.400 73.050 336.600 ;
        RECT 49.950 334.950 52.050 335.400 ;
        RECT 64.950 334.950 67.050 335.400 ;
        RECT 70.950 334.950 73.050 335.400 ;
        RECT 124.950 336.600 127.050 337.050 ;
        RECT 142.950 336.600 145.050 337.050 ;
        RECT 124.950 335.400 145.050 336.600 ;
        RECT 124.950 334.950 127.050 335.400 ;
        RECT 142.950 334.950 145.050 335.400 ;
        RECT 145.950 336.600 148.050 337.050 ;
        RECT 163.950 336.600 166.050 337.050 ;
        RECT 145.950 335.400 166.050 336.600 ;
        RECT 145.950 334.950 148.050 335.400 ;
        RECT 163.950 334.950 166.050 335.400 ;
        RECT 178.950 336.600 181.050 337.050 ;
        RECT 199.950 336.600 202.050 337.050 ;
        RECT 178.950 335.400 202.050 336.600 ;
        RECT 206.400 336.600 207.600 338.400 ;
        RECT 211.950 338.400 220.050 339.600 ;
        RECT 211.950 337.950 214.050 338.400 ;
        RECT 217.950 337.950 220.050 338.400 ;
        RECT 235.950 339.600 238.050 340.050 ;
        RECT 247.950 339.600 250.050 340.050 ;
        RECT 235.950 338.400 250.050 339.600 ;
        RECT 235.950 337.950 238.050 338.400 ;
        RECT 247.950 337.950 250.050 338.400 ;
        RECT 268.950 339.600 271.050 340.050 ;
        RECT 337.950 339.600 340.050 340.050 ;
        RECT 343.950 339.600 346.050 340.050 ;
        RECT 268.950 338.400 336.600 339.600 ;
        RECT 268.950 337.950 271.050 338.400 ;
        RECT 235.950 336.600 238.050 337.050 ;
        RECT 206.400 335.400 238.050 336.600 ;
        RECT 178.950 334.950 181.050 335.400 ;
        RECT 199.950 334.950 202.050 335.400 ;
        RECT 235.950 334.950 238.050 335.400 ;
        RECT 274.950 336.600 277.050 337.050 ;
        RECT 286.950 336.600 289.050 337.050 ;
        RECT 274.950 335.400 289.050 336.600 ;
        RECT 335.400 336.600 336.600 338.400 ;
        RECT 337.950 338.400 346.050 339.600 ;
        RECT 337.950 337.950 340.050 338.400 ;
        RECT 343.950 337.950 346.050 338.400 ;
        RECT 346.950 337.950 349.050 340.050 ;
        RECT 356.400 337.050 357.600 340.950 ;
        RECT 461.400 340.050 462.600 341.400 ;
        RECT 476.400 341.400 526.050 342.600 ;
        RECT 476.400 340.050 477.600 341.400 ;
        RECT 523.950 340.950 526.050 341.400 ;
        RECT 539.400 341.400 544.050 342.600 ;
        RECT 539.400 340.050 540.600 341.400 ;
        RECT 541.950 340.950 544.050 341.400 ;
        RECT 547.950 342.600 550.050 343.050 ;
        RECT 556.950 342.600 559.050 343.050 ;
        RECT 547.950 341.400 552.600 342.600 ;
        RECT 547.950 340.950 550.050 341.400 ;
        RECT 551.400 340.050 552.600 341.400 ;
        RECT 556.950 341.400 567.600 342.600 ;
        RECT 556.950 340.950 559.050 341.400 ;
        RECT 566.400 340.050 567.600 341.400 ;
        RECT 572.400 340.050 573.600 343.950 ;
        RECT 586.950 340.950 589.050 343.050 ;
        RECT 361.950 339.600 364.050 340.050 ;
        RECT 385.950 339.600 388.050 340.050 ;
        RECT 361.950 338.400 388.050 339.600 ;
        RECT 361.950 337.950 364.050 338.400 ;
        RECT 385.950 337.950 388.050 338.400 ;
        RECT 418.950 339.600 421.050 340.050 ;
        RECT 439.950 339.600 442.050 340.050 ;
        RECT 418.950 338.400 442.050 339.600 ;
        RECT 418.950 337.950 421.050 338.400 ;
        RECT 439.950 337.950 442.050 338.400 ;
        RECT 445.950 339.600 448.050 340.050 ;
        RECT 457.950 339.600 460.050 340.050 ;
        RECT 445.950 338.400 460.050 339.600 ;
        RECT 445.950 337.950 448.050 338.400 ;
        RECT 457.950 337.950 460.050 338.400 ;
        RECT 460.950 337.950 463.050 340.050 ;
        RECT 475.950 337.950 478.050 340.050 ;
        RECT 478.950 339.600 481.050 340.050 ;
        RECT 484.950 339.600 487.050 340.050 ;
        RECT 487.950 339.600 490.050 340.050 ;
        RECT 478.950 338.400 490.050 339.600 ;
        RECT 478.950 337.950 481.050 338.400 ;
        RECT 484.950 337.950 487.050 338.400 ;
        RECT 487.950 337.950 490.050 338.400 ;
        RECT 505.950 339.600 508.050 340.050 ;
        RECT 526.950 339.600 529.050 340.050 ;
        RECT 505.950 338.400 529.050 339.600 ;
        RECT 505.950 337.950 508.050 338.400 ;
        RECT 526.950 337.950 529.050 338.400 ;
        RECT 538.950 337.950 541.050 340.050 ;
        RECT 544.950 339.600 547.050 340.050 ;
        RECT 550.950 339.600 553.050 340.050 ;
        RECT 544.950 338.400 553.050 339.600 ;
        RECT 544.950 337.950 547.050 338.400 ;
        RECT 550.950 337.950 553.050 338.400 ;
        RECT 565.950 337.950 568.050 340.050 ;
        RECT 571.950 337.950 574.050 340.050 ;
        RECT 587.400 339.600 588.600 340.950 ;
        RECT 590.400 340.050 591.600 343.950 ;
        RECT 593.400 343.050 594.600 350.400 ;
        RECT 619.950 349.950 622.050 350.400 ;
        RECT 685.950 351.600 688.050 352.050 ;
        RECT 715.950 351.600 718.050 352.050 ;
        RECT 685.950 350.400 718.050 351.600 ;
        RECT 685.950 349.950 688.050 350.400 ;
        RECT 715.950 349.950 718.050 350.400 ;
        RECT 595.950 348.600 598.050 349.050 ;
        RECT 685.950 348.600 688.050 349.050 ;
        RECT 703.950 348.600 706.050 349.050 ;
        RECT 595.950 347.400 612.600 348.600 ;
        RECT 595.950 346.950 598.050 347.400 ;
        RECT 607.950 345.600 610.050 346.050 ;
        RECT 602.400 344.400 610.050 345.600 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 602.400 340.050 603.600 344.400 ;
        RECT 607.950 343.950 610.050 344.400 ;
        RECT 604.950 340.950 607.050 343.050 ;
        RECT 575.400 338.400 588.600 339.600 ;
        RECT 589.950 339.600 592.050 340.050 ;
        RECT 589.950 338.400 600.600 339.600 ;
        RECT 340.950 336.600 343.050 337.050 ;
        RECT 352.950 336.600 355.050 337.050 ;
        RECT 335.400 335.400 339.600 336.600 ;
        RECT 274.950 334.950 277.050 335.400 ;
        RECT 286.950 334.950 289.050 335.400 ;
        RECT 338.400 334.050 339.600 335.400 ;
        RECT 340.950 335.400 355.050 336.600 ;
        RECT 340.950 334.950 343.050 335.400 ;
        RECT 352.950 334.950 355.050 335.400 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 379.950 336.600 382.050 337.050 ;
        RECT 391.950 336.600 394.050 337.050 ;
        RECT 379.950 335.400 394.050 336.600 ;
        RECT 379.950 334.950 382.050 335.400 ;
        RECT 391.950 334.950 394.050 335.400 ;
        RECT 439.950 336.600 442.050 337.050 ;
        RECT 499.950 336.600 502.050 337.050 ;
        RECT 523.950 336.600 526.050 337.050 ;
        RECT 439.950 335.400 526.050 336.600 ;
        RECT 439.950 334.950 442.050 335.400 ;
        RECT 499.950 334.950 502.050 335.400 ;
        RECT 523.950 334.950 526.050 335.400 ;
        RECT 538.950 336.600 541.050 337.050 ;
        RECT 547.950 336.600 550.050 337.050 ;
        RECT 538.950 335.400 550.050 336.600 ;
        RECT 538.950 334.950 541.050 335.400 ;
        RECT 547.950 334.950 550.050 335.400 ;
        RECT 556.950 336.600 559.050 337.050 ;
        RECT 575.400 336.600 576.600 338.400 ;
        RECT 589.950 337.950 592.050 338.400 ;
        RECT 599.400 337.050 600.600 338.400 ;
        RECT 601.950 337.950 604.050 340.050 ;
        RECT 556.950 335.400 576.600 336.600 ;
        RECT 577.950 336.600 580.050 337.050 ;
        RECT 595.950 336.600 598.050 337.050 ;
        RECT 577.950 335.400 598.050 336.600 ;
        RECT 556.950 334.950 559.050 335.400 ;
        RECT 577.950 334.950 580.050 335.400 ;
        RECT 595.950 334.950 598.050 335.400 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 605.400 336.600 606.600 340.950 ;
        RECT 602.400 335.400 606.600 336.600 ;
        RECT 602.400 334.050 603.600 335.400 ;
        RECT 31.950 333.600 34.050 334.050 ;
        RECT 2.400 332.400 34.050 333.600 ;
        RECT 31.950 331.950 34.050 332.400 ;
        RECT 34.950 333.600 37.050 334.050 ;
        RECT 40.950 333.600 43.050 334.050 ;
        RECT 34.950 332.400 43.050 333.600 ;
        RECT 34.950 331.950 37.050 332.400 ;
        RECT 40.950 331.950 43.050 332.400 ;
        RECT 58.950 333.600 61.050 334.050 ;
        RECT 76.950 333.600 79.050 334.050 ;
        RECT 85.950 333.600 88.050 334.050 ;
        RECT 58.950 332.400 88.050 333.600 ;
        RECT 58.950 331.950 61.050 332.400 ;
        RECT 76.950 331.950 79.050 332.400 ;
        RECT 85.950 331.950 88.050 332.400 ;
        RECT 124.950 333.600 127.050 334.050 ;
        RECT 139.950 333.600 142.050 334.050 ;
        RECT 124.950 332.400 142.050 333.600 ;
        RECT 124.950 331.950 127.050 332.400 ;
        RECT 139.950 331.950 142.050 332.400 ;
        RECT 145.950 333.600 148.050 334.050 ;
        RECT 169.950 333.600 172.050 334.050 ;
        RECT 145.950 332.400 172.050 333.600 ;
        RECT 145.950 331.950 148.050 332.400 ;
        RECT 169.950 331.950 172.050 332.400 ;
        RECT 229.950 333.600 232.050 334.050 ;
        RECT 250.950 333.600 253.050 334.050 ;
        RECT 229.950 332.400 253.050 333.600 ;
        RECT 229.950 331.950 232.050 332.400 ;
        RECT 250.950 331.950 253.050 332.400 ;
        RECT 280.950 333.600 283.050 334.050 ;
        RECT 292.950 333.600 295.050 334.050 ;
        RECT 316.950 333.600 319.050 334.050 ;
        RECT 328.950 333.600 331.050 334.050 ;
        RECT 280.950 332.400 319.050 333.600 ;
        RECT 280.950 331.950 283.050 332.400 ;
        RECT 292.950 331.950 295.050 332.400 ;
        RECT 316.950 331.950 319.050 332.400 ;
        RECT 326.400 332.400 331.050 333.600 ;
        RECT 22.950 330.600 25.050 331.050 ;
        RECT 52.950 330.600 55.050 331.050 ;
        RECT 82.950 330.600 85.050 331.050 ;
        RECT 97.950 330.600 100.050 331.050 ;
        RECT 22.950 329.400 100.050 330.600 ;
        RECT 22.950 328.950 25.050 329.400 ;
        RECT 52.950 328.950 55.050 329.400 ;
        RECT 82.950 328.950 85.050 329.400 ;
        RECT 97.950 328.950 100.050 329.400 ;
        RECT 121.950 330.600 124.050 331.050 ;
        RECT 136.950 330.600 139.050 331.050 ;
        RECT 121.950 329.400 139.050 330.600 ;
        RECT 121.950 328.950 124.050 329.400 ;
        RECT 136.950 328.950 139.050 329.400 ;
        RECT 205.950 330.600 208.050 331.050 ;
        RECT 256.950 330.600 259.050 331.050 ;
        RECT 205.950 329.400 259.050 330.600 ;
        RECT 205.950 328.950 208.050 329.400 ;
        RECT 256.950 328.950 259.050 329.400 ;
        RECT 271.950 330.600 274.050 331.050 ;
        RECT 289.950 330.600 292.050 331.050 ;
        RECT 271.950 329.400 292.050 330.600 ;
        RECT 271.950 328.950 274.050 329.400 ;
        RECT 289.950 328.950 292.050 329.400 ;
        RECT 326.400 328.050 327.600 332.400 ;
        RECT 328.950 331.950 331.050 332.400 ;
        RECT 337.950 331.950 340.050 334.050 ;
        RECT 397.950 333.600 400.050 334.050 ;
        RECT 481.950 333.600 484.050 334.050 ;
        RECT 397.950 332.400 484.050 333.600 ;
        RECT 397.950 331.950 400.050 332.400 ;
        RECT 481.950 331.950 484.050 332.400 ;
        RECT 502.950 333.600 505.050 334.050 ;
        RECT 526.950 333.600 529.050 334.050 ;
        RECT 502.950 332.400 529.050 333.600 ;
        RECT 502.950 331.950 505.050 332.400 ;
        RECT 526.950 331.950 529.050 332.400 ;
        RECT 601.950 331.950 604.050 334.050 ;
        RECT 604.950 333.600 607.050 334.050 ;
        RECT 611.400 333.600 612.600 347.400 ;
        RECT 685.950 347.400 706.050 348.600 ;
        RECT 685.950 346.950 688.050 347.400 ;
        RECT 703.950 346.950 706.050 347.400 ;
        RECT 649.950 345.600 652.050 346.050 ;
        RECT 679.950 345.600 682.050 346.050 ;
        RECT 697.950 345.600 700.050 346.050 ;
        RECT 649.950 344.400 700.050 345.600 ;
        RECT 649.950 343.950 652.050 344.400 ;
        RECT 679.950 343.950 682.050 344.400 ;
        RECT 697.950 343.950 700.050 344.400 ;
        RECT 691.950 342.600 694.050 343.050 ;
        RECT 700.950 342.600 703.050 343.050 ;
        RECT 691.950 341.400 703.050 342.600 ;
        RECT 691.950 340.950 694.050 341.400 ;
        RECT 700.950 340.950 703.050 341.400 ;
        RECT 631.950 339.600 634.050 340.050 ;
        RECT 661.950 339.600 664.050 340.050 ;
        RECT 631.950 338.400 664.050 339.600 ;
        RECT 631.950 337.950 634.050 338.400 ;
        RECT 661.950 337.950 664.050 338.400 ;
        RECT 667.950 339.600 670.050 340.050 ;
        RECT 688.950 339.600 691.050 340.050 ;
        RECT 667.950 338.400 691.050 339.600 ;
        RECT 667.950 337.950 670.050 338.400 ;
        RECT 688.950 337.950 691.050 338.400 ;
        RECT 700.950 339.600 703.050 340.050 ;
        RECT 709.950 339.600 712.050 340.050 ;
        RECT 700.950 338.400 712.050 339.600 ;
        RECT 700.950 337.950 703.050 338.400 ;
        RECT 709.950 337.950 712.050 338.400 ;
        RECT 622.950 336.600 625.050 337.050 ;
        RECT 634.950 336.600 637.050 337.050 ;
        RECT 622.950 335.400 637.050 336.600 ;
        RECT 622.950 334.950 625.050 335.400 ;
        RECT 634.950 334.950 637.050 335.400 ;
        RECT 604.950 332.400 612.600 333.600 ;
        RECT 604.950 331.950 607.050 332.400 ;
        RECT 367.950 330.600 370.050 331.050 ;
        RECT 403.950 330.600 406.050 331.050 ;
        RECT 442.950 330.600 445.050 331.050 ;
        RECT 367.950 329.400 445.050 330.600 ;
        RECT 367.950 328.950 370.050 329.400 ;
        RECT 403.950 328.950 406.050 329.400 ;
        RECT 442.950 328.950 445.050 329.400 ;
        RECT 466.950 330.600 469.050 331.050 ;
        RECT 493.950 330.600 496.050 331.050 ;
        RECT 466.950 329.400 496.050 330.600 ;
        RECT 466.950 328.950 469.050 329.400 ;
        RECT 493.950 328.950 496.050 329.400 ;
        RECT 538.950 330.600 541.050 331.050 ;
        RECT 562.950 330.600 565.050 331.050 ;
        RECT 574.950 330.600 577.050 331.050 ;
        RECT 538.950 329.400 577.050 330.600 ;
        RECT 538.950 328.950 541.050 329.400 ;
        RECT 562.950 328.950 565.050 329.400 ;
        RECT 574.950 328.950 577.050 329.400 ;
        RECT 1.950 327.600 4.050 328.050 ;
        RECT 46.950 327.600 49.050 328.050 ;
        RECT 1.950 326.400 49.050 327.600 ;
        RECT 1.950 325.950 4.050 326.400 ;
        RECT 46.950 325.950 49.050 326.400 ;
        RECT 85.950 327.600 88.050 328.050 ;
        RECT 106.950 327.600 109.050 328.050 ;
        RECT 85.950 326.400 109.050 327.600 ;
        RECT 85.950 325.950 88.050 326.400 ;
        RECT 106.950 325.950 109.050 326.400 ;
        RECT 244.950 327.600 247.050 328.050 ;
        RECT 253.950 327.600 256.050 328.050 ;
        RECT 244.950 326.400 256.050 327.600 ;
        RECT 244.950 325.950 247.050 326.400 ;
        RECT 253.950 325.950 256.050 326.400 ;
        RECT 265.950 327.600 268.050 328.050 ;
        RECT 298.950 327.600 301.050 328.050 ;
        RECT 265.950 326.400 301.050 327.600 ;
        RECT 265.950 325.950 268.050 326.400 ;
        RECT 298.950 325.950 301.050 326.400 ;
        RECT 325.950 325.950 328.050 328.050 ;
        RECT 433.950 327.600 436.050 328.050 ;
        RECT 445.950 327.600 448.050 328.050 ;
        RECT 451.950 327.600 454.050 328.050 ;
        RECT 469.950 327.600 472.050 328.050 ;
        RECT 475.950 327.600 478.050 328.050 ;
        RECT 433.950 326.400 478.050 327.600 ;
        RECT 433.950 325.950 436.050 326.400 ;
        RECT 445.950 325.950 448.050 326.400 ;
        RECT 451.950 325.950 454.050 326.400 ;
        RECT 469.950 325.950 472.050 326.400 ;
        RECT 475.950 325.950 478.050 326.400 ;
        RECT 535.950 327.600 538.050 328.050 ;
        RECT 682.950 327.600 685.050 328.050 ;
        RECT 535.950 326.400 685.050 327.600 ;
        RECT 535.950 325.950 538.050 326.400 ;
        RECT 682.950 325.950 685.050 326.400 ;
        RECT 40.950 324.600 43.050 325.050 ;
        RECT 79.950 324.600 82.050 325.050 ;
        RECT 133.950 324.600 136.050 325.050 ;
        RECT 40.950 323.400 136.050 324.600 ;
        RECT 40.950 322.950 43.050 323.400 ;
        RECT 79.950 322.950 82.050 323.400 ;
        RECT 133.950 322.950 136.050 323.400 ;
        RECT 253.950 324.600 256.050 325.050 ;
        RECT 271.950 324.600 274.050 325.050 ;
        RECT 253.950 323.400 274.050 324.600 ;
        RECT 253.950 322.950 256.050 323.400 ;
        RECT 271.950 322.950 274.050 323.400 ;
        RECT 274.950 324.600 277.050 325.050 ;
        RECT 280.950 324.600 283.050 325.050 ;
        RECT 274.950 323.400 283.050 324.600 ;
        RECT 274.950 322.950 277.050 323.400 ;
        RECT 280.950 322.950 283.050 323.400 ;
        RECT 289.950 324.600 292.050 325.050 ;
        RECT 334.950 324.600 337.050 325.050 ;
        RECT 289.950 323.400 337.050 324.600 ;
        RECT 289.950 322.950 292.050 323.400 ;
        RECT 334.950 322.950 337.050 323.400 ;
        RECT 379.950 324.600 382.050 325.050 ;
        RECT 388.950 324.600 391.050 325.050 ;
        RECT 400.950 324.600 403.050 325.050 ;
        RECT 379.950 323.400 403.050 324.600 ;
        RECT 379.950 322.950 382.050 323.400 ;
        RECT 388.950 322.950 391.050 323.400 ;
        RECT 400.950 322.950 403.050 323.400 ;
        RECT 436.950 324.600 439.050 325.050 ;
        RECT 487.950 324.600 490.050 325.050 ;
        RECT 436.950 323.400 490.050 324.600 ;
        RECT 436.950 322.950 439.050 323.400 ;
        RECT 487.950 322.950 490.050 323.400 ;
        RECT 679.950 324.600 682.050 325.050 ;
        RECT 688.950 324.600 691.050 325.050 ;
        RECT 679.950 323.400 691.050 324.600 ;
        RECT 679.950 322.950 682.050 323.400 ;
        RECT 688.950 322.950 691.050 323.400 ;
        RECT 25.950 321.600 28.050 322.050 ;
        RECT 112.950 321.600 115.050 322.050 ;
        RECT 25.950 320.400 115.050 321.600 ;
        RECT 25.950 319.950 28.050 320.400 ;
        RECT 112.950 319.950 115.050 320.400 ;
        RECT 196.950 321.600 199.050 322.050 ;
        RECT 262.950 321.600 265.050 322.050 ;
        RECT 307.950 321.600 310.050 322.050 ;
        RECT 196.950 320.400 310.050 321.600 ;
        RECT 196.950 319.950 199.050 320.400 ;
        RECT 262.950 319.950 265.050 320.400 ;
        RECT 307.950 319.950 310.050 320.400 ;
        RECT 322.950 321.600 325.050 322.050 ;
        RECT 343.950 321.600 346.050 322.050 ;
        RECT 322.950 320.400 346.050 321.600 ;
        RECT 322.950 319.950 325.050 320.400 ;
        RECT 343.950 319.950 346.050 320.400 ;
        RECT 397.950 321.600 400.050 322.050 ;
        RECT 490.950 321.600 493.050 322.050 ;
        RECT 397.950 320.400 493.050 321.600 ;
        RECT 397.950 319.950 400.050 320.400 ;
        RECT 490.950 319.950 493.050 320.400 ;
        RECT 550.950 321.600 553.050 322.050 ;
        RECT 568.950 321.600 571.050 322.050 ;
        RECT 550.950 320.400 571.050 321.600 ;
        RECT 550.950 319.950 553.050 320.400 ;
        RECT 568.950 319.950 571.050 320.400 ;
        RECT 571.950 321.600 574.050 322.050 ;
        RECT 589.950 321.600 592.050 322.050 ;
        RECT 571.950 320.400 592.050 321.600 ;
        RECT 571.950 319.950 574.050 320.400 ;
        RECT 589.950 319.950 592.050 320.400 ;
        RECT 643.950 321.600 646.050 322.050 ;
        RECT 655.950 321.600 658.050 322.050 ;
        RECT 643.950 320.400 658.050 321.600 ;
        RECT 643.950 319.950 646.050 320.400 ;
        RECT 655.950 319.950 658.050 320.400 ;
        RECT 661.950 321.600 664.050 322.050 ;
        RECT 679.950 321.600 682.050 322.050 ;
        RECT 694.950 321.600 697.050 322.050 ;
        RECT 661.950 320.400 697.050 321.600 ;
        RECT 661.950 319.950 664.050 320.400 ;
        RECT 679.950 319.950 682.050 320.400 ;
        RECT 694.950 319.950 697.050 320.400 ;
        RECT 67.950 318.600 70.050 319.050 ;
        RECT 85.950 318.600 88.050 319.050 ;
        RECT 67.950 317.400 88.050 318.600 ;
        RECT 67.950 316.950 70.050 317.400 ;
        RECT 85.950 316.950 88.050 317.400 ;
        RECT 94.950 318.600 97.050 319.050 ;
        RECT 106.950 318.600 109.050 319.050 ;
        RECT 118.950 318.600 121.050 319.050 ;
        RECT 94.950 317.400 109.050 318.600 ;
        RECT 94.950 316.950 97.050 317.400 ;
        RECT 106.950 316.950 109.050 317.400 ;
        RECT 110.400 317.400 121.050 318.600 ;
        RECT 7.950 315.600 10.050 316.050 ;
        RECT 5.400 314.400 10.050 315.600 ;
        RECT 5.400 306.600 6.600 314.400 ;
        RECT 7.950 313.950 10.050 314.400 ;
        RECT 52.950 315.600 55.050 316.050 ;
        RECT 70.950 315.600 73.050 316.050 ;
        RECT 110.400 315.600 111.600 317.400 ;
        RECT 118.950 316.950 121.050 317.400 ;
        RECT 139.950 318.600 142.050 319.050 ;
        RECT 154.950 318.600 157.050 319.050 ;
        RECT 139.950 317.400 157.050 318.600 ;
        RECT 139.950 316.950 142.050 317.400 ;
        RECT 154.950 316.950 157.050 317.400 ;
        RECT 247.950 318.600 250.050 319.050 ;
        RECT 283.950 318.600 286.050 319.050 ;
        RECT 247.950 317.400 286.050 318.600 ;
        RECT 247.950 316.950 250.050 317.400 ;
        RECT 283.950 316.950 286.050 317.400 ;
        RECT 286.950 318.600 289.050 319.050 ;
        RECT 295.950 318.600 298.050 319.050 ;
        RECT 286.950 317.400 298.050 318.600 ;
        RECT 286.950 316.950 289.050 317.400 ;
        RECT 295.950 316.950 298.050 317.400 ;
        RECT 307.950 318.600 310.050 319.050 ;
        RECT 331.950 318.600 334.050 319.050 ;
        RECT 307.950 317.400 334.050 318.600 ;
        RECT 307.950 316.950 310.050 317.400 ;
        RECT 331.950 316.950 334.050 317.400 ;
        RECT 448.950 318.600 451.050 319.050 ;
        RECT 454.950 318.600 457.050 319.050 ;
        RECT 448.950 317.400 457.050 318.600 ;
        RECT 448.950 316.950 451.050 317.400 ;
        RECT 454.950 316.950 457.050 317.400 ;
        RECT 478.950 318.600 481.050 319.050 ;
        RECT 529.950 318.600 532.050 319.050 ;
        RECT 646.950 318.600 649.050 319.050 ;
        RECT 670.950 318.600 673.050 319.050 ;
        RECT 478.950 317.400 486.600 318.600 ;
        RECT 478.950 316.950 481.050 317.400 ;
        RECT 52.950 314.400 60.600 315.600 ;
        RECT 52.950 313.950 55.050 314.400 ;
        RECT 7.950 312.600 10.050 313.050 ;
        RECT 19.950 312.600 22.050 313.050 ;
        RECT 25.950 312.600 28.050 313.050 ;
        RECT 7.950 311.400 22.050 312.600 ;
        RECT 7.950 310.950 10.050 311.400 ;
        RECT 19.950 310.950 22.050 311.400 ;
        RECT 23.400 311.400 28.050 312.600 ;
        RECT 23.400 309.600 24.600 311.400 ;
        RECT 25.950 310.950 28.050 311.400 ;
        RECT 31.950 310.950 34.050 313.050 ;
        RECT 34.950 310.950 37.050 313.050 ;
        RECT 37.950 312.600 40.050 313.050 ;
        RECT 52.950 312.600 55.050 313.050 ;
        RECT 37.950 311.400 45.600 312.600 ;
        RECT 37.950 310.950 40.050 311.400 ;
        RECT 14.400 308.400 24.600 309.600 ;
        RECT 14.400 307.050 15.600 308.400 ;
        RECT 10.950 306.600 13.050 307.050 ;
        RECT 5.400 305.400 13.050 306.600 ;
        RECT 10.950 304.950 13.050 305.400 ;
        RECT 13.950 304.950 16.050 307.050 ;
        RECT 25.950 306.600 28.050 307.050 ;
        RECT 32.400 306.600 33.600 310.950 ;
        RECT 25.950 305.400 33.600 306.600 ;
        RECT 25.950 304.950 28.050 305.400 ;
        RECT 35.400 304.050 36.600 310.950 ;
        RECT 44.400 310.050 45.600 311.400 ;
        RECT 52.950 311.400 57.600 312.600 ;
        RECT 52.950 310.950 55.050 311.400 ;
        RECT 40.950 307.950 43.050 310.050 ;
        RECT 43.950 307.950 46.050 310.050 ;
        RECT 37.950 304.950 40.050 307.050 ;
        RECT 41.400 306.600 42.600 307.950 ;
        RECT 49.950 306.600 52.050 307.050 ;
        RECT 41.400 305.400 52.050 306.600 ;
        RECT 56.400 306.600 57.600 311.400 ;
        RECT 59.400 310.050 60.600 314.400 ;
        RECT 62.400 314.400 73.050 315.600 ;
        RECT 62.400 310.050 63.600 314.400 ;
        RECT 70.950 313.950 73.050 314.400 ;
        RECT 74.400 314.400 111.600 315.600 ;
        RECT 74.400 312.600 75.600 314.400 ;
        RECT 115.950 313.950 118.050 316.050 ;
        RECT 118.950 315.600 121.050 316.050 ;
        RECT 133.950 315.600 136.050 316.050 ;
        RECT 151.950 315.600 154.050 316.050 ;
        RECT 118.950 314.400 132.600 315.600 ;
        RECT 118.950 313.950 121.050 314.400 ;
        RECT 65.400 311.400 75.600 312.600 ;
        RECT 65.400 310.050 66.600 311.400 ;
        RECT 97.950 310.950 100.050 313.050 ;
        RECT 116.400 312.600 117.600 313.950 ;
        RECT 121.950 312.600 124.050 313.050 ;
        RECT 113.400 311.400 117.600 312.600 ;
        RECT 119.400 311.400 124.050 312.600 ;
        RECT 131.400 312.600 132.600 314.400 ;
        RECT 133.950 314.400 154.050 315.600 ;
        RECT 133.950 313.950 136.050 314.400 ;
        RECT 151.950 313.950 154.050 314.400 ;
        RECT 166.950 315.600 169.050 316.050 ;
        RECT 181.950 315.600 184.050 316.050 ;
        RECT 211.950 315.600 214.050 316.050 ;
        RECT 166.950 314.400 184.050 315.600 ;
        RECT 166.950 313.950 169.050 314.400 ;
        RECT 181.950 313.950 184.050 314.400 ;
        RECT 185.400 314.400 214.050 315.600 ;
        RECT 139.950 312.600 142.050 313.050 ;
        RECT 131.400 311.400 142.050 312.600 ;
        RECT 58.950 307.950 61.050 310.050 ;
        RECT 61.950 307.950 64.050 310.050 ;
        RECT 64.950 307.950 67.050 310.050 ;
        RECT 88.950 309.600 91.050 310.050 ;
        RECT 80.400 308.400 91.050 309.600 ;
        RECT 58.950 306.600 61.050 307.050 ;
        RECT 56.400 305.400 61.050 306.600 ;
        RECT 49.950 304.950 52.050 305.400 ;
        RECT 58.950 304.950 61.050 305.400 ;
        RECT 64.950 306.600 67.050 307.050 ;
        RECT 76.950 306.600 79.050 307.050 ;
        RECT 64.950 305.400 79.050 306.600 ;
        RECT 64.950 304.950 67.050 305.400 ;
        RECT 76.950 304.950 79.050 305.400 ;
        RECT 34.950 301.950 37.050 304.050 ;
        RECT 1.950 300.600 4.050 301.050 ;
        RECT 38.400 300.600 39.600 304.950 ;
        RECT 80.400 303.600 81.600 308.400 ;
        RECT 88.950 307.950 91.050 308.400 ;
        RECT 94.950 307.950 97.050 310.050 ;
        RECT 98.400 309.600 99.600 310.950 ;
        RECT 103.950 309.600 106.050 310.050 ;
        RECT 98.400 308.400 106.050 309.600 ;
        RECT 103.950 307.950 106.050 308.400 ;
        RECT 82.950 306.600 85.050 307.050 ;
        RECT 95.400 306.600 96.600 307.950 ;
        RECT 113.400 307.050 114.600 311.400 ;
        RECT 106.950 306.600 109.050 307.050 ;
        RECT 82.950 305.400 109.050 306.600 ;
        RECT 82.950 304.950 85.050 305.400 ;
        RECT 106.950 304.950 109.050 305.400 ;
        RECT 112.950 304.950 115.050 307.050 ;
        RECT 119.400 306.600 120.600 311.400 ;
        RECT 121.950 310.950 124.050 311.400 ;
        RECT 139.950 310.950 142.050 311.400 ;
        RECT 142.950 310.950 145.050 313.050 ;
        RECT 148.950 312.600 151.050 313.050 ;
        RECT 148.950 311.400 159.600 312.600 ;
        RECT 148.950 310.950 151.050 311.400 ;
        RECT 121.950 309.600 124.050 310.050 ;
        RECT 136.950 309.600 139.050 310.050 ;
        RECT 121.950 308.400 139.050 309.600 ;
        RECT 121.950 307.950 124.050 308.400 ;
        RECT 136.950 307.950 139.050 308.400 ;
        RECT 130.950 306.600 133.050 307.050 ;
        RECT 119.400 305.400 133.050 306.600 ;
        RECT 130.950 304.950 133.050 305.400 ;
        RECT 136.950 304.950 139.050 307.050 ;
        RECT 143.400 306.600 144.600 310.950 ;
        RECT 151.950 309.600 154.050 310.050 ;
        RECT 151.950 308.400 156.600 309.600 ;
        RECT 151.950 307.950 154.050 308.400 ;
        RECT 140.400 305.400 144.600 306.600 ;
        RECT 94.950 303.600 97.050 304.050 ;
        RECT 118.950 303.600 121.050 304.050 ;
        RECT 80.400 302.400 84.600 303.600 ;
        RECT 76.950 300.600 79.050 301.050 ;
        RECT 1.950 299.400 39.600 300.600 ;
        RECT 41.400 299.400 79.050 300.600 ;
        RECT 83.400 300.600 84.600 302.400 ;
        RECT 94.950 302.400 121.050 303.600 ;
        RECT 94.950 301.950 97.050 302.400 ;
        RECT 118.950 301.950 121.050 302.400 ;
        RECT 133.950 303.600 136.050 304.050 ;
        RECT 137.400 303.600 138.600 304.950 ;
        RECT 140.400 304.050 141.600 305.400 ;
        RECT 151.950 304.950 154.050 307.050 ;
        RECT 133.950 302.400 138.600 303.600 ;
        RECT 133.950 301.950 136.050 302.400 ;
        RECT 139.950 301.950 142.050 304.050 ;
        RECT 148.950 303.600 151.050 304.050 ;
        RECT 152.400 303.600 153.600 304.950 ;
        RECT 155.400 304.050 156.600 308.400 ;
        RECT 158.400 304.050 159.600 311.400 ;
        RECT 163.950 307.950 166.050 310.050 ;
        RECT 169.950 309.600 172.050 310.050 ;
        RECT 178.950 309.600 181.050 310.050 ;
        RECT 169.950 308.400 181.050 309.600 ;
        RECT 169.950 307.950 172.050 308.400 ;
        RECT 178.950 307.950 181.050 308.400 ;
        RECT 181.950 309.600 184.050 310.050 ;
        RECT 185.400 309.600 186.600 314.400 ;
        RECT 211.950 313.950 214.050 314.400 ;
        RECT 259.950 313.950 262.050 316.050 ;
        RECT 262.950 313.950 265.050 316.050 ;
        RECT 277.950 315.600 280.050 316.050 ;
        RECT 289.950 315.600 292.050 316.050 ;
        RECT 277.950 314.400 292.050 315.600 ;
        RECT 277.950 313.950 280.050 314.400 ;
        RECT 289.950 313.950 292.050 314.400 ;
        RECT 292.950 313.950 295.050 316.050 ;
        RECT 340.950 315.600 343.050 316.050 ;
        RECT 358.950 315.600 361.050 316.050 ;
        RECT 385.950 315.600 388.050 316.050 ;
        RECT 340.950 314.400 388.050 315.600 ;
        RECT 340.950 313.950 343.050 314.400 ;
        RECT 358.950 313.950 361.050 314.400 ;
        RECT 385.950 313.950 388.050 314.400 ;
        RECT 457.950 315.600 460.050 316.050 ;
        RECT 481.950 315.600 484.050 316.050 ;
        RECT 457.950 314.400 484.050 315.600 ;
        RECT 457.950 313.950 460.050 314.400 ;
        RECT 481.950 313.950 484.050 314.400 ;
        RECT 187.950 312.600 190.050 313.050 ;
        RECT 193.950 312.600 196.050 313.050 ;
        RECT 187.950 311.400 196.050 312.600 ;
        RECT 187.950 310.950 190.050 311.400 ;
        RECT 193.950 310.950 196.050 311.400 ;
        RECT 199.950 312.600 202.050 313.050 ;
        RECT 205.950 312.600 208.050 313.050 ;
        RECT 199.950 311.400 208.050 312.600 ;
        RECT 199.950 310.950 202.050 311.400 ;
        RECT 205.950 310.950 208.050 311.400 ;
        RECT 232.950 312.600 235.050 313.050 ;
        RECT 253.950 312.600 256.050 313.050 ;
        RECT 232.950 311.400 256.050 312.600 ;
        RECT 232.950 310.950 235.050 311.400 ;
        RECT 253.950 310.950 256.050 311.400 ;
        RECT 260.400 310.050 261.600 313.950 ;
        RECT 263.400 310.050 264.600 313.950 ;
        RECT 286.950 310.950 289.050 313.050 ;
        RECT 293.400 312.600 294.600 313.950 ;
        RECT 290.400 311.400 294.600 312.600 ;
        RECT 304.950 312.600 307.050 313.050 ;
        RECT 316.950 312.600 319.050 313.050 ;
        RECT 304.950 311.400 319.050 312.600 ;
        RECT 181.950 308.400 186.600 309.600 ;
        RECT 190.950 309.600 193.050 310.050 ;
        RECT 196.950 309.600 199.050 310.050 ;
        RECT 190.950 308.400 199.050 309.600 ;
        RECT 181.950 307.950 184.050 308.400 ;
        RECT 190.950 307.950 193.050 308.400 ;
        RECT 196.950 307.950 199.050 308.400 ;
        RECT 223.950 309.600 226.050 310.050 ;
        RECT 244.950 309.600 247.050 310.050 ;
        RECT 223.950 308.400 247.050 309.600 ;
        RECT 223.950 307.950 226.050 308.400 ;
        RECT 244.950 307.950 247.050 308.400 ;
        RECT 250.950 309.600 253.050 310.050 ;
        RECT 256.950 309.600 259.050 310.050 ;
        RECT 250.950 308.400 259.050 309.600 ;
        RECT 250.950 307.950 253.050 308.400 ;
        RECT 256.950 307.950 259.050 308.400 ;
        RECT 259.950 307.950 262.050 310.050 ;
        RECT 262.950 307.950 265.050 310.050 ;
        RECT 164.400 304.050 165.600 307.950 ;
        RECT 172.950 306.600 175.050 307.050 ;
        RECT 214.950 306.600 217.050 307.050 ;
        RECT 229.950 306.600 232.050 307.050 ;
        RECT 172.950 305.400 232.050 306.600 ;
        RECT 172.950 304.950 175.050 305.400 ;
        RECT 214.950 304.950 217.050 305.400 ;
        RECT 229.950 304.950 232.050 305.400 ;
        RECT 148.950 302.400 153.600 303.600 ;
        RECT 148.950 301.950 151.050 302.400 ;
        RECT 154.950 301.950 157.050 304.050 ;
        RECT 157.950 301.950 160.050 304.050 ;
        RECT 163.950 301.950 166.050 304.050 ;
        RECT 208.950 303.600 211.050 304.050 ;
        RECT 259.950 303.600 262.050 304.050 ;
        RECT 283.950 303.600 286.050 304.050 ;
        RECT 208.950 302.400 286.050 303.600 ;
        RECT 287.400 303.600 288.600 310.950 ;
        RECT 290.400 307.050 291.600 311.400 ;
        RECT 304.950 310.950 307.050 311.400 ;
        RECT 316.950 310.950 319.050 311.400 ;
        RECT 382.950 312.600 385.050 313.050 ;
        RECT 400.950 312.600 403.050 313.050 ;
        RECT 382.950 311.400 403.050 312.600 ;
        RECT 382.950 310.950 385.050 311.400 ;
        RECT 400.950 310.950 403.050 311.400 ;
        RECT 436.950 312.600 439.050 313.050 ;
        RECT 463.950 312.600 466.050 313.050 ;
        RECT 475.950 312.600 478.050 313.050 ;
        RECT 485.400 312.600 486.600 317.400 ;
        RECT 529.950 317.400 673.050 318.600 ;
        RECT 529.950 316.950 532.050 317.400 ;
        RECT 646.950 316.950 649.050 317.400 ;
        RECT 670.950 316.950 673.050 317.400 ;
        RECT 541.950 315.600 544.050 316.050 ;
        RECT 571.950 315.600 574.050 316.050 ;
        RECT 541.950 314.400 574.050 315.600 ;
        RECT 541.950 313.950 544.050 314.400 ;
        RECT 571.950 313.950 574.050 314.400 ;
        RECT 574.950 315.600 577.050 316.050 ;
        RECT 607.950 315.600 610.050 316.050 ;
        RECT 628.950 315.600 631.050 316.050 ;
        RECT 574.950 314.400 631.050 315.600 ;
        RECT 574.950 313.950 577.050 314.400 ;
        RECT 607.950 313.950 610.050 314.400 ;
        RECT 628.950 313.950 631.050 314.400 ;
        RECT 649.950 313.950 652.050 316.050 ;
        RECT 652.950 315.600 655.050 316.050 ;
        RECT 661.950 315.600 664.050 316.050 ;
        RECT 652.950 314.400 664.050 315.600 ;
        RECT 652.950 313.950 655.050 314.400 ;
        RECT 661.950 313.950 664.050 314.400 ;
        RECT 673.950 313.950 676.050 316.050 ;
        RECT 436.950 311.400 466.050 312.600 ;
        RECT 436.950 310.950 439.050 311.400 ;
        RECT 463.950 310.950 466.050 311.400 ;
        RECT 473.400 311.400 478.050 312.600 ;
        RECT 473.400 310.050 474.600 311.400 ;
        RECT 475.950 310.950 478.050 311.400 ;
        RECT 479.400 311.400 486.600 312.600 ;
        RECT 496.950 312.600 499.050 313.050 ;
        RECT 517.950 312.600 520.050 313.050 ;
        RECT 496.950 311.400 520.050 312.600 ;
        RECT 292.950 309.600 295.050 310.050 ;
        RECT 313.950 309.600 316.050 310.050 ;
        RECT 292.950 308.400 316.050 309.600 ;
        RECT 292.950 307.950 295.050 308.400 ;
        RECT 313.950 307.950 316.050 308.400 ;
        RECT 349.950 309.600 352.050 310.050 ;
        RECT 361.950 309.600 364.050 310.050 ;
        RECT 349.950 308.400 364.050 309.600 ;
        RECT 349.950 307.950 352.050 308.400 ;
        RECT 361.950 307.950 364.050 308.400 ;
        RECT 406.950 309.600 409.050 310.050 ;
        RECT 415.950 309.600 418.050 310.050 ;
        RECT 469.950 309.600 472.050 310.050 ;
        RECT 406.950 308.400 414.600 309.600 ;
        RECT 406.950 307.950 409.050 308.400 ;
        RECT 413.400 307.050 414.600 308.400 ;
        RECT 415.950 308.400 472.050 309.600 ;
        RECT 415.950 307.950 418.050 308.400 ;
        RECT 469.950 307.950 472.050 308.400 ;
        RECT 472.950 307.950 475.050 310.050 ;
        RECT 479.400 309.600 480.600 311.400 ;
        RECT 496.950 310.950 499.050 311.400 ;
        RECT 517.950 310.950 520.050 311.400 ;
        RECT 529.950 312.600 532.050 313.050 ;
        RECT 535.950 312.600 538.050 313.050 ;
        RECT 529.950 311.400 538.050 312.600 ;
        RECT 529.950 310.950 532.050 311.400 ;
        RECT 535.950 310.950 538.050 311.400 ;
        RECT 541.950 310.950 544.050 313.050 ;
        RECT 547.950 312.600 550.050 313.050 ;
        RECT 568.950 312.600 571.050 313.050 ;
        RECT 547.950 311.400 571.050 312.600 ;
        RECT 547.950 310.950 550.050 311.400 ;
        RECT 568.950 310.950 571.050 311.400 ;
        RECT 580.950 312.600 583.050 313.050 ;
        RECT 595.950 312.600 598.050 313.050 ;
        RECT 604.950 312.600 607.050 313.050 ;
        RECT 580.950 311.400 607.050 312.600 ;
        RECT 580.950 310.950 583.050 311.400 ;
        RECT 595.950 310.950 598.050 311.400 ;
        RECT 604.950 310.950 607.050 311.400 ;
        RECT 613.950 310.950 616.050 313.050 ;
        RECT 650.400 312.600 651.600 313.950 ;
        RECT 647.400 311.400 651.600 312.600 ;
        RECT 476.400 308.400 480.600 309.600 ;
        RECT 487.950 309.600 490.050 310.050 ;
        RECT 493.950 309.600 496.050 310.050 ;
        RECT 487.950 308.400 496.050 309.600 ;
        RECT 289.950 304.950 292.050 307.050 ;
        RECT 400.950 306.600 403.050 307.050 ;
        RECT 409.950 306.600 412.050 307.050 ;
        RECT 400.950 305.400 412.050 306.600 ;
        RECT 400.950 304.950 403.050 305.400 ;
        RECT 409.950 304.950 412.050 305.400 ;
        RECT 412.950 304.950 415.050 307.050 ;
        RECT 418.950 306.600 421.050 307.050 ;
        RECT 436.950 306.600 439.050 307.050 ;
        RECT 418.950 305.400 439.050 306.600 ;
        RECT 418.950 304.950 421.050 305.400 ;
        RECT 436.950 304.950 439.050 305.400 ;
        RECT 466.950 306.600 469.050 307.050 ;
        RECT 476.400 306.600 477.600 308.400 ;
        RECT 487.950 307.950 490.050 308.400 ;
        RECT 493.950 307.950 496.050 308.400 ;
        RECT 499.950 309.600 502.050 310.050 ;
        RECT 542.400 309.600 543.600 310.950 ;
        RECT 499.950 308.400 543.600 309.600 ;
        RECT 586.950 309.600 589.050 310.050 ;
        RECT 614.400 309.600 615.600 310.950 ;
        RECT 647.400 310.050 648.600 311.400 ;
        RECT 674.400 310.050 675.600 313.950 ;
        RECT 676.950 312.600 679.050 313.050 ;
        RECT 682.950 312.600 685.050 313.050 ;
        RECT 676.950 311.400 685.050 312.600 ;
        RECT 676.950 310.950 679.050 311.400 ;
        RECT 682.950 310.950 685.050 311.400 ;
        RECT 586.950 308.400 615.600 309.600 ;
        RECT 499.950 307.950 502.050 308.400 ;
        RECT 586.950 307.950 589.050 308.400 ;
        RECT 646.950 307.950 649.050 310.050 ;
        RECT 649.950 309.600 652.050 310.050 ;
        RECT 655.950 309.600 658.050 310.050 ;
        RECT 649.950 308.400 658.050 309.600 ;
        RECT 649.950 307.950 652.050 308.400 ;
        RECT 655.950 307.950 658.050 308.400 ;
        RECT 673.950 307.950 676.050 310.050 ;
        RECT 466.950 305.400 477.600 306.600 ;
        RECT 505.950 306.600 508.050 307.050 ;
        RECT 649.950 306.600 652.050 307.050 ;
        RECT 505.950 305.400 652.050 306.600 ;
        RECT 466.950 304.950 469.050 305.400 ;
        RECT 505.950 304.950 508.050 305.400 ;
        RECT 649.950 304.950 652.050 305.400 ;
        RECT 298.950 303.600 301.050 304.050 ;
        RECT 287.400 302.400 301.050 303.600 ;
        RECT 208.950 301.950 211.050 302.400 ;
        RECT 259.950 301.950 262.050 302.400 ;
        RECT 283.950 301.950 286.050 302.400 ;
        RECT 298.950 301.950 301.050 302.400 ;
        RECT 568.950 303.600 571.050 304.050 ;
        RECT 571.950 303.600 574.050 304.050 ;
        RECT 607.950 303.600 610.050 304.050 ;
        RECT 568.950 302.400 610.050 303.600 ;
        RECT 568.950 301.950 571.050 302.400 ;
        RECT 571.950 301.950 574.050 302.400 ;
        RECT 607.950 301.950 610.050 302.400 ;
        RECT 109.950 300.600 112.050 301.050 ;
        RECT 83.400 299.400 112.050 300.600 ;
        RECT 1.950 298.950 4.050 299.400 ;
        RECT 25.950 297.600 28.050 298.050 ;
        RECT 41.400 297.600 42.600 299.400 ;
        RECT 76.950 298.950 79.050 299.400 ;
        RECT 109.950 298.950 112.050 299.400 ;
        RECT 115.950 300.600 118.050 301.050 ;
        RECT 127.950 300.600 130.050 301.050 ;
        RECT 115.950 299.400 130.050 300.600 ;
        RECT 115.950 298.950 118.050 299.400 ;
        RECT 127.950 298.950 130.050 299.400 ;
        RECT 145.950 300.600 148.050 301.050 ;
        RECT 160.950 300.600 163.050 301.050 ;
        RECT 145.950 299.400 163.050 300.600 ;
        RECT 145.950 298.950 148.050 299.400 ;
        RECT 160.950 298.950 163.050 299.400 ;
        RECT 166.950 300.600 169.050 301.050 ;
        RECT 175.950 300.600 178.050 301.050 ;
        RECT 166.950 299.400 178.050 300.600 ;
        RECT 166.950 298.950 169.050 299.400 ;
        RECT 175.950 298.950 178.050 299.400 ;
        RECT 226.950 300.600 229.050 301.050 ;
        RECT 235.950 300.600 238.050 301.050 ;
        RECT 226.950 299.400 238.050 300.600 ;
        RECT 226.950 298.950 229.050 299.400 ;
        RECT 235.950 298.950 238.050 299.400 ;
        RECT 280.950 300.600 283.050 301.050 ;
        RECT 301.950 300.600 304.050 301.050 ;
        RECT 280.950 299.400 304.050 300.600 ;
        RECT 280.950 298.950 283.050 299.400 ;
        RECT 301.950 298.950 304.050 299.400 ;
        RECT 391.950 300.600 394.050 301.050 ;
        RECT 403.950 300.600 406.050 301.050 ;
        RECT 412.950 300.600 415.050 301.050 ;
        RECT 391.950 299.400 415.050 300.600 ;
        RECT 391.950 298.950 394.050 299.400 ;
        RECT 403.950 298.950 406.050 299.400 ;
        RECT 412.950 298.950 415.050 299.400 ;
        RECT 469.950 300.600 472.050 301.050 ;
        RECT 544.950 300.600 547.050 301.050 ;
        RECT 469.950 299.400 547.050 300.600 ;
        RECT 469.950 298.950 472.050 299.400 ;
        RECT 544.950 298.950 547.050 299.400 ;
        RECT 25.950 296.400 42.600 297.600 ;
        RECT 97.950 297.600 100.050 298.050 ;
        RECT 133.950 297.600 136.050 298.050 ;
        RECT 148.950 297.600 151.050 298.050 ;
        RECT 97.950 296.400 151.050 297.600 ;
        RECT 25.950 295.950 28.050 296.400 ;
        RECT 97.950 295.950 100.050 296.400 ;
        RECT 133.950 295.950 136.050 296.400 ;
        RECT 148.950 295.950 151.050 296.400 ;
        RECT 202.950 297.600 205.050 298.050 ;
        RECT 247.950 297.600 250.050 298.050 ;
        RECT 202.950 296.400 250.050 297.600 ;
        RECT 202.950 295.950 205.050 296.400 ;
        RECT 247.950 295.950 250.050 296.400 ;
        RECT 286.950 297.600 289.050 298.050 ;
        RECT 334.950 297.600 337.050 298.050 ;
        RECT 286.950 296.400 337.050 297.600 ;
        RECT 286.950 295.950 289.050 296.400 ;
        RECT 334.950 295.950 337.050 296.400 ;
        RECT 355.950 297.600 358.050 298.050 ;
        RECT 397.950 297.600 400.050 298.050 ;
        RECT 355.950 296.400 400.050 297.600 ;
        RECT 355.950 295.950 358.050 296.400 ;
        RECT 397.950 295.950 400.050 296.400 ;
        RECT 31.950 294.600 34.050 295.050 ;
        RECT 103.950 294.600 106.050 295.050 ;
        RECT 127.950 294.600 130.050 295.050 ;
        RECT 31.950 293.400 130.050 294.600 ;
        RECT 31.950 292.950 34.050 293.400 ;
        RECT 103.950 292.950 106.050 293.400 ;
        RECT 127.950 292.950 130.050 293.400 ;
        RECT 376.950 294.600 379.050 295.050 ;
        RECT 400.950 294.600 403.050 295.050 ;
        RECT 376.950 293.400 403.050 294.600 ;
        RECT 376.950 292.950 379.050 293.400 ;
        RECT 400.950 292.950 403.050 293.400 ;
        RECT 598.950 294.600 601.050 295.050 ;
        RECT 610.950 294.600 613.050 295.050 ;
        RECT 598.950 293.400 613.050 294.600 ;
        RECT 598.950 292.950 601.050 293.400 ;
        RECT 610.950 292.950 613.050 293.400 ;
        RECT 34.950 291.600 37.050 292.050 ;
        RECT 43.950 291.600 46.050 292.050 ;
        RECT 34.950 290.400 46.050 291.600 ;
        RECT 34.950 289.950 37.050 290.400 ;
        RECT 43.950 289.950 46.050 290.400 ;
        RECT 310.950 291.600 313.050 292.050 ;
        RECT 313.950 291.600 316.050 292.050 ;
        RECT 322.950 291.600 325.050 292.050 ;
        RECT 358.950 291.600 361.050 292.050 ;
        RECT 310.950 290.400 361.050 291.600 ;
        RECT 310.950 289.950 313.050 290.400 ;
        RECT 313.950 289.950 316.050 290.400 ;
        RECT 322.950 289.950 325.050 290.400 ;
        RECT 358.950 289.950 361.050 290.400 ;
        RECT 421.950 291.600 424.050 292.050 ;
        RECT 490.950 291.600 493.050 292.050 ;
        RECT 421.950 290.400 493.050 291.600 ;
        RECT 421.950 289.950 424.050 290.400 ;
        RECT 490.950 289.950 493.050 290.400 ;
        RECT 541.950 291.600 544.050 292.050 ;
        RECT 556.950 291.600 559.050 292.050 ;
        RECT 541.950 290.400 559.050 291.600 ;
        RECT 541.950 289.950 544.050 290.400 ;
        RECT 556.950 289.950 559.050 290.400 ;
        RECT 583.950 291.600 586.050 292.050 ;
        RECT 601.950 291.600 604.050 292.050 ;
        RECT 583.950 290.400 604.050 291.600 ;
        RECT 583.950 289.950 586.050 290.400 ;
        RECT 601.950 289.950 604.050 290.400 ;
        RECT 622.950 291.600 625.050 292.050 ;
        RECT 628.950 291.600 631.050 292.050 ;
        RECT 622.950 290.400 631.050 291.600 ;
        RECT 622.950 289.950 625.050 290.400 ;
        RECT 628.950 289.950 631.050 290.400 ;
        RECT 34.950 288.600 37.050 289.050 ;
        RECT 82.950 288.600 85.050 289.050 ;
        RECT 34.950 287.400 85.050 288.600 ;
        RECT 34.950 286.950 37.050 287.400 ;
        RECT 82.950 286.950 85.050 287.400 ;
        RECT 628.950 288.600 631.050 289.050 ;
        RECT 634.950 288.600 637.050 289.050 ;
        RECT 628.950 287.400 637.050 288.600 ;
        RECT 628.950 286.950 631.050 287.400 ;
        RECT 634.950 286.950 637.050 287.400 ;
        RECT 106.950 285.600 109.050 286.050 ;
        RECT 151.950 285.600 154.050 286.050 ;
        RECT 106.950 284.400 154.050 285.600 ;
        RECT 106.950 283.950 109.050 284.400 ;
        RECT 151.950 283.950 154.050 284.400 ;
        RECT 256.950 285.600 259.050 286.050 ;
        RECT 262.950 285.600 265.050 286.050 ;
        RECT 256.950 284.400 265.050 285.600 ;
        RECT 256.950 283.950 259.050 284.400 ;
        RECT 262.950 283.950 265.050 284.400 ;
        RECT 1.950 282.600 4.050 283.050 ;
        RECT 13.950 282.600 16.050 283.050 ;
        RECT 1.950 281.400 16.050 282.600 ;
        RECT 1.950 280.950 4.050 281.400 ;
        RECT 13.950 280.950 16.050 281.400 ;
        RECT 58.950 282.600 61.050 283.050 ;
        RECT 124.950 282.600 127.050 283.050 ;
        RECT 133.950 282.600 136.050 283.050 ;
        RECT 58.950 281.400 136.050 282.600 ;
        RECT 58.950 280.950 61.050 281.400 ;
        RECT 124.950 280.950 127.050 281.400 ;
        RECT 133.950 280.950 136.050 281.400 ;
        RECT 142.950 282.600 145.050 283.050 ;
        RECT 214.950 282.600 217.050 283.050 ;
        RECT 142.950 281.400 217.050 282.600 ;
        RECT 142.950 280.950 145.050 281.400 ;
        RECT 214.950 280.950 217.050 281.400 ;
        RECT 4.950 279.600 7.050 280.050 ;
        RECT 31.950 279.600 34.050 280.050 ;
        RECT 4.950 278.400 34.050 279.600 ;
        RECT 4.950 277.950 7.050 278.400 ;
        RECT 31.950 277.950 34.050 278.400 ;
        RECT 43.950 279.600 46.050 280.050 ;
        RECT 55.950 279.600 58.050 280.050 ;
        RECT 67.950 279.600 70.050 280.050 ;
        RECT 43.950 278.400 70.050 279.600 ;
        RECT 43.950 277.950 46.050 278.400 ;
        RECT 55.950 277.950 58.050 278.400 ;
        RECT 67.950 277.950 70.050 278.400 ;
        RECT 85.950 279.600 88.050 280.050 ;
        RECT 121.950 279.600 124.050 280.050 ;
        RECT 85.950 278.400 124.050 279.600 ;
        RECT 85.950 277.950 88.050 278.400 ;
        RECT 121.950 277.950 124.050 278.400 ;
        RECT 130.950 279.600 133.050 280.050 ;
        RECT 142.950 279.600 145.050 280.050 ;
        RECT 130.950 278.400 145.050 279.600 ;
        RECT 130.950 277.950 133.050 278.400 ;
        RECT 142.950 277.950 145.050 278.400 ;
        RECT 154.950 279.600 157.050 280.050 ;
        RECT 172.950 279.600 175.050 280.050 ;
        RECT 154.950 278.400 175.050 279.600 ;
        RECT 154.950 277.950 157.050 278.400 ;
        RECT 172.950 277.950 175.050 278.400 ;
        RECT 328.950 279.600 331.050 280.050 ;
        RECT 358.950 279.600 361.050 280.050 ;
        RECT 439.950 279.600 442.050 280.050 ;
        RECT 472.950 279.600 475.050 280.050 ;
        RECT 532.950 279.600 535.050 280.050 ;
        RECT 328.950 278.400 535.050 279.600 ;
        RECT 328.950 277.950 331.050 278.400 ;
        RECT 358.950 277.950 361.050 278.400 ;
        RECT 439.950 277.950 442.050 278.400 ;
        RECT 472.950 277.950 475.050 278.400 ;
        RECT 532.950 277.950 535.050 278.400 ;
        RECT 547.950 279.600 550.050 280.050 ;
        RECT 616.950 279.600 619.050 280.050 ;
        RECT 547.950 278.400 619.050 279.600 ;
        RECT 547.950 277.950 550.050 278.400 ;
        RECT 616.950 277.950 619.050 278.400 ;
        RECT 7.950 274.950 10.050 277.050 ;
        RECT 16.950 276.600 19.050 277.050 ;
        RECT 34.950 276.600 37.050 277.050 ;
        RECT 61.950 276.600 64.050 277.050 ;
        RECT 16.950 275.400 37.050 276.600 ;
        RECT 16.950 274.950 19.050 275.400 ;
        RECT 34.950 274.950 37.050 275.400 ;
        RECT 47.400 275.400 64.050 276.600 ;
        RECT 8.400 264.600 9.600 274.950 ;
        RECT 10.950 271.950 13.050 274.050 ;
        RECT 13.950 273.600 16.050 274.050 ;
        RECT 31.950 273.600 34.050 274.050 ;
        RECT 47.400 273.600 48.600 275.400 ;
        RECT 61.950 274.950 64.050 275.400 ;
        RECT 70.950 276.600 73.050 277.050 ;
        RECT 106.950 276.600 109.050 277.050 ;
        RECT 70.950 275.400 109.050 276.600 ;
        RECT 70.950 274.950 73.050 275.400 ;
        RECT 106.950 274.950 109.050 275.400 ;
        RECT 127.950 276.600 130.050 277.050 ;
        RECT 151.950 276.600 154.050 277.050 ;
        RECT 127.950 275.400 147.600 276.600 ;
        RECT 127.950 274.950 130.050 275.400 ;
        RECT 13.950 272.400 48.600 273.600 ;
        RECT 13.950 271.950 16.050 272.400 ;
        RECT 31.950 271.950 34.050 272.400 ;
        RECT 49.950 271.950 52.050 274.050 ;
        RECT 55.950 273.600 58.050 274.050 ;
        RECT 64.950 273.600 67.050 274.050 ;
        RECT 85.950 273.600 88.050 274.050 ;
        RECT 100.950 273.600 103.050 274.050 ;
        RECT 55.950 272.400 103.050 273.600 ;
        RECT 55.950 271.950 58.050 272.400 ;
        RECT 64.950 271.950 67.050 272.400 ;
        RECT 85.950 271.950 88.050 272.400 ;
        RECT 100.950 271.950 103.050 272.400 ;
        RECT 109.950 273.600 112.050 274.050 ;
        RECT 121.950 273.600 124.050 274.050 ;
        RECT 109.950 272.400 120.600 273.600 ;
        RECT 109.950 271.950 112.050 272.400 ;
        RECT 11.400 268.050 12.600 271.950 ;
        RECT 22.950 270.600 25.050 271.050 ;
        RECT 28.950 270.600 31.050 271.050 ;
        RECT 37.950 270.600 40.050 271.050 ;
        RECT 22.950 269.400 27.600 270.600 ;
        RECT 22.950 268.950 25.050 269.400 ;
        RECT 10.950 265.950 13.050 268.050 ;
        RECT 26.400 267.600 27.600 269.400 ;
        RECT 28.950 269.400 40.050 270.600 ;
        RECT 28.950 268.950 31.050 269.400 ;
        RECT 37.950 268.950 40.050 269.400 ;
        RECT 50.400 268.050 51.600 271.950 ;
        RECT 119.400 271.050 120.600 272.400 ;
        RECT 121.950 272.400 129.600 273.600 ;
        RECT 121.950 271.950 124.050 272.400 ;
        RECT 100.950 270.600 103.050 271.050 ;
        RECT 100.950 269.400 108.600 270.600 ;
        RECT 100.950 268.950 103.050 269.400 ;
        RECT 40.950 267.600 43.050 268.050 ;
        RECT 26.400 266.400 43.050 267.600 ;
        RECT 40.950 265.950 43.050 266.400 ;
        RECT 49.950 265.950 52.050 268.050 ;
        RECT 55.950 267.600 58.050 268.050 ;
        RECT 67.950 267.600 70.050 268.050 ;
        RECT 55.950 266.400 70.050 267.600 ;
        RECT 55.950 265.950 58.050 266.400 ;
        RECT 67.950 265.950 70.050 266.400 ;
        RECT 73.950 267.600 76.050 268.050 ;
        RECT 79.950 267.600 82.050 268.050 ;
        RECT 73.950 266.400 82.050 267.600 ;
        RECT 107.400 267.600 108.600 269.400 ;
        RECT 118.950 268.950 121.050 271.050 ;
        RECT 109.950 267.600 112.050 268.050 ;
        RECT 107.400 266.400 112.050 267.600 ;
        RECT 73.950 265.950 76.050 266.400 ;
        RECT 79.950 265.950 82.050 266.400 ;
        RECT 109.950 265.950 112.050 266.400 ;
        RECT 13.950 264.600 16.050 265.050 ;
        RECT 8.400 263.400 16.050 264.600 ;
        RECT 13.950 262.950 16.050 263.400 ;
        RECT 37.950 264.600 40.050 265.050 ;
        RECT 52.950 264.600 55.050 265.050 ;
        RECT 79.950 264.600 82.050 265.050 ;
        RECT 88.950 264.600 91.050 265.050 ;
        RECT 37.950 263.400 55.050 264.600 ;
        RECT 37.950 262.950 40.050 263.400 ;
        RECT 52.950 262.950 55.050 263.400 ;
        RECT 56.400 263.400 91.050 264.600 ;
        RECT 4.950 261.600 7.050 262.050 ;
        RECT 25.950 261.600 28.050 262.050 ;
        RECT 4.950 260.400 28.050 261.600 ;
        RECT 4.950 259.950 7.050 260.400 ;
        RECT 25.950 259.950 28.050 260.400 ;
        RECT 31.950 261.600 34.050 262.050 ;
        RECT 56.400 261.600 57.600 263.400 ;
        RECT 79.950 262.950 82.050 263.400 ;
        RECT 88.950 262.950 91.050 263.400 ;
        RECT 94.950 264.600 97.050 265.050 ;
        RECT 119.400 264.600 120.600 268.950 ;
        RECT 128.400 268.050 129.600 272.400 ;
        RECT 136.950 271.950 139.050 274.050 ;
        RECT 121.950 267.600 124.050 268.050 ;
        RECT 127.950 267.600 130.050 268.050 ;
        RECT 130.950 267.600 133.050 268.050 ;
        RECT 121.950 266.400 126.600 267.600 ;
        RECT 121.950 265.950 124.050 266.400 ;
        RECT 121.950 264.600 124.050 265.050 ;
        RECT 94.950 263.400 117.600 264.600 ;
        RECT 119.400 263.400 124.050 264.600 ;
        RECT 125.400 264.600 126.600 266.400 ;
        RECT 127.950 266.400 133.050 267.600 ;
        RECT 127.950 265.950 130.050 266.400 ;
        RECT 130.950 265.950 133.050 266.400 ;
        RECT 127.950 264.600 130.050 265.050 ;
        RECT 125.400 263.400 130.050 264.600 ;
        RECT 94.950 262.950 97.050 263.400 ;
        RECT 31.950 260.400 57.600 261.600 ;
        RECT 61.950 261.600 64.050 262.050 ;
        RECT 76.950 261.600 79.050 262.050 ;
        RECT 97.950 261.600 100.050 262.050 ;
        RECT 112.950 261.600 115.050 262.050 ;
        RECT 61.950 260.400 79.050 261.600 ;
        RECT 31.950 259.950 34.050 260.400 ;
        RECT 61.950 259.950 64.050 260.400 ;
        RECT 76.950 259.950 79.050 260.400 ;
        RECT 89.400 260.400 115.050 261.600 ;
        RECT 116.400 261.600 117.600 263.400 ;
        RECT 121.950 262.950 124.050 263.400 ;
        RECT 127.950 262.950 130.050 263.400 ;
        RECT 130.950 264.600 133.050 265.050 ;
        RECT 137.400 264.600 138.600 271.950 ;
        RECT 146.400 271.050 147.600 275.400 ;
        RECT 149.400 275.400 154.050 276.600 ;
        RECT 149.400 274.050 150.600 275.400 ;
        RECT 151.950 274.950 154.050 275.400 ;
        RECT 154.950 276.600 157.050 277.050 ;
        RECT 163.950 276.600 166.050 277.050 ;
        RECT 184.950 276.600 187.050 277.050 ;
        RECT 154.950 275.400 162.600 276.600 ;
        RECT 154.950 274.950 157.050 275.400 ;
        RECT 148.950 271.950 151.050 274.050 ;
        RECT 154.950 271.950 157.050 274.050 ;
        RECT 157.950 271.950 160.050 274.050 ;
        RECT 161.400 273.600 162.600 275.400 ;
        RECT 163.950 275.400 187.050 276.600 ;
        RECT 163.950 274.950 166.050 275.400 ;
        RECT 163.950 273.600 166.050 274.050 ;
        RECT 161.400 272.400 166.050 273.600 ;
        RECT 163.950 271.950 166.050 272.400 ;
        RECT 145.950 268.950 148.050 271.050 ;
        RECT 155.400 268.050 156.600 271.950 ;
        RECT 139.950 267.600 142.050 268.050 ;
        RECT 151.950 267.600 154.050 268.050 ;
        RECT 139.950 266.400 154.050 267.600 ;
        RECT 139.950 265.950 142.050 266.400 ;
        RECT 151.950 265.950 154.050 266.400 ;
        RECT 154.950 265.950 157.050 268.050 ;
        RECT 130.950 263.400 138.600 264.600 ;
        RECT 158.400 264.600 159.600 271.950 ;
        RECT 170.400 268.050 171.600 275.400 ;
        RECT 184.950 274.950 187.050 275.400 ;
        RECT 190.950 274.950 193.050 277.050 ;
        RECT 322.950 276.600 325.050 277.050 ;
        RECT 340.950 276.600 343.050 277.050 ;
        RECT 409.950 276.600 412.050 277.050 ;
        RECT 322.950 275.400 343.050 276.600 ;
        RECT 322.950 274.950 325.050 275.400 ;
        RECT 340.950 274.950 343.050 275.400 ;
        RECT 407.400 275.400 412.050 276.600 ;
        RECT 172.950 273.600 175.050 274.050 ;
        RECT 187.950 273.600 190.050 274.050 ;
        RECT 172.950 272.400 190.050 273.600 ;
        RECT 172.950 271.950 175.050 272.400 ;
        RECT 187.950 271.950 190.050 272.400 ;
        RECT 169.950 265.950 172.050 268.050 ;
        RECT 191.400 267.600 192.600 274.950 ;
        RECT 193.950 273.600 196.050 274.050 ;
        RECT 214.950 273.600 217.050 274.050 ;
        RECT 229.950 273.600 232.050 274.050 ;
        RECT 193.950 272.400 210.600 273.600 ;
        RECT 193.950 271.950 196.050 272.400 ;
        RECT 209.400 270.600 210.600 272.400 ;
        RECT 214.950 272.400 232.050 273.600 ;
        RECT 214.950 271.950 217.050 272.400 ;
        RECT 229.950 271.950 232.050 272.400 ;
        RECT 241.950 273.600 244.050 274.050 ;
        RECT 250.950 273.600 253.050 274.050 ;
        RECT 241.950 272.400 253.050 273.600 ;
        RECT 241.950 271.950 244.050 272.400 ;
        RECT 250.950 271.950 253.050 272.400 ;
        RECT 268.950 273.600 271.050 274.050 ;
        RECT 289.950 273.600 292.050 274.050 ;
        RECT 268.950 272.400 292.050 273.600 ;
        RECT 268.950 271.950 271.050 272.400 ;
        RECT 289.950 271.950 292.050 272.400 ;
        RECT 310.950 273.600 313.050 274.050 ;
        RECT 328.950 273.600 331.050 274.050 ;
        RECT 310.950 272.400 331.050 273.600 ;
        RECT 310.950 271.950 313.050 272.400 ;
        RECT 328.950 271.950 331.050 272.400 ;
        RECT 349.950 273.600 352.050 274.050 ;
        RECT 349.950 272.400 357.600 273.600 ;
        RECT 349.950 271.950 352.050 272.400 ;
        RECT 356.400 271.050 357.600 272.400 ;
        RECT 220.950 270.600 223.050 271.050 ;
        RECT 229.950 270.600 232.050 271.050 ;
        RECT 209.400 269.400 213.600 270.600 ;
        RECT 212.400 268.050 213.600 269.400 ;
        RECT 220.950 269.400 232.050 270.600 ;
        RECT 220.950 268.950 223.050 269.400 ;
        RECT 229.950 268.950 232.050 269.400 ;
        RECT 232.950 270.600 235.050 271.050 ;
        RECT 244.950 270.600 247.050 271.050 ;
        RECT 232.950 269.400 247.050 270.600 ;
        RECT 232.950 268.950 235.050 269.400 ;
        RECT 244.950 268.950 247.050 269.400 ;
        RECT 325.950 270.600 328.050 271.050 ;
        RECT 337.950 270.600 340.050 271.050 ;
        RECT 325.950 269.400 340.050 270.600 ;
        RECT 325.950 268.950 328.050 269.400 ;
        RECT 337.950 268.950 340.050 269.400 ;
        RECT 340.950 270.600 343.050 271.050 ;
        RECT 349.950 270.600 352.050 271.050 ;
        RECT 340.950 269.400 352.050 270.600 ;
        RECT 340.950 268.950 343.050 269.400 ;
        RECT 349.950 268.950 352.050 269.400 ;
        RECT 355.950 268.950 358.050 271.050 ;
        RECT 388.950 268.950 391.050 271.050 ;
        RECT 394.950 268.950 397.050 271.050 ;
        RECT 193.950 267.600 196.050 268.050 ;
        RECT 191.400 266.400 196.050 267.600 ;
        RECT 193.950 265.950 196.050 266.400 ;
        RECT 211.950 267.600 214.050 268.050 ;
        RECT 226.950 267.600 229.050 268.050 ;
        RECT 211.950 266.400 229.050 267.600 ;
        RECT 211.950 265.950 214.050 266.400 ;
        RECT 226.950 265.950 229.050 266.400 ;
        RECT 259.950 267.600 262.050 268.050 ;
        RECT 271.950 267.600 274.050 268.050 ;
        RECT 277.950 267.600 280.050 268.050 ;
        RECT 259.950 266.400 280.050 267.600 ;
        RECT 259.950 265.950 262.050 266.400 ;
        RECT 271.950 265.950 274.050 266.400 ;
        RECT 277.950 265.950 280.050 266.400 ;
        RECT 319.950 267.600 322.050 268.050 ;
        RECT 328.950 267.600 331.050 268.050 ;
        RECT 319.950 266.400 331.050 267.600 ;
        RECT 350.400 267.600 351.600 268.950 ;
        RECT 373.950 267.600 376.050 268.050 ;
        RECT 350.400 266.400 376.050 267.600 ;
        RECT 319.950 265.950 322.050 266.400 ;
        RECT 328.950 265.950 331.050 266.400 ;
        RECT 373.950 265.950 376.050 266.400 ;
        RECT 379.950 267.600 382.050 268.050 ;
        RECT 389.400 267.600 390.600 268.950 ;
        RECT 379.950 266.400 390.600 267.600 ;
        RECT 395.400 267.600 396.600 268.950 ;
        RECT 403.950 267.600 406.050 268.050 ;
        RECT 395.400 266.400 406.050 267.600 ;
        RECT 379.950 265.950 382.050 266.400 ;
        RECT 403.950 265.950 406.050 266.400 ;
        RECT 160.950 264.600 163.050 265.050 ;
        RECT 184.950 264.600 187.050 265.050 ;
        RECT 158.400 263.400 187.050 264.600 ;
        RECT 130.950 262.950 133.050 263.400 ;
        RECT 160.950 262.950 163.050 263.400 ;
        RECT 184.950 262.950 187.050 263.400 ;
        RECT 223.950 264.600 226.050 265.050 ;
        RECT 244.950 264.600 247.050 265.050 ;
        RECT 223.950 263.400 247.050 264.600 ;
        RECT 223.950 262.950 226.050 263.400 ;
        RECT 244.950 262.950 247.050 263.400 ;
        RECT 265.950 264.600 268.050 265.050 ;
        RECT 274.950 264.600 277.050 265.050 ;
        RECT 265.950 263.400 277.050 264.600 ;
        RECT 265.950 262.950 268.050 263.400 ;
        RECT 274.950 262.950 277.050 263.400 ;
        RECT 331.950 264.600 334.050 265.050 ;
        RECT 361.950 264.600 364.050 265.050 ;
        RECT 331.950 263.400 364.050 264.600 ;
        RECT 331.950 262.950 334.050 263.400 ;
        RECT 361.950 262.950 364.050 263.400 ;
        RECT 373.950 264.600 376.050 265.050 ;
        RECT 385.950 264.600 388.050 265.050 ;
        RECT 373.950 263.400 388.050 264.600 ;
        RECT 407.400 264.600 408.600 275.400 ;
        RECT 409.950 274.950 412.050 275.400 ;
        RECT 493.950 276.600 496.050 277.050 ;
        RECT 499.950 276.600 502.050 277.050 ;
        RECT 517.950 276.600 520.050 277.050 ;
        RECT 571.950 276.600 574.050 277.050 ;
        RECT 640.950 276.600 643.050 277.050 ;
        RECT 493.950 275.400 643.050 276.600 ;
        RECT 493.950 274.950 496.050 275.400 ;
        RECT 499.950 274.950 502.050 275.400 ;
        RECT 517.950 274.950 520.050 275.400 ;
        RECT 571.950 274.950 574.050 275.400 ;
        RECT 640.950 274.950 643.050 275.400 ;
        RECT 676.950 276.600 679.050 277.050 ;
        RECT 682.950 276.600 685.050 277.050 ;
        RECT 676.950 275.400 685.050 276.600 ;
        RECT 676.950 274.950 679.050 275.400 ;
        RECT 682.950 274.950 685.050 275.400 ;
        RECT 409.950 273.600 412.050 274.050 ;
        RECT 457.950 273.600 460.050 274.050 ;
        RECT 469.950 273.600 472.050 274.050 ;
        RECT 409.950 272.400 420.600 273.600 ;
        RECT 409.950 271.950 412.050 272.400 ;
        RECT 419.400 270.600 420.600 272.400 ;
        RECT 457.950 272.400 472.050 273.600 ;
        RECT 457.950 271.950 460.050 272.400 ;
        RECT 469.950 271.950 472.050 272.400 ;
        RECT 511.950 273.600 514.050 274.050 ;
        RECT 526.950 273.600 529.050 274.050 ;
        RECT 511.950 272.400 529.050 273.600 ;
        RECT 511.950 271.950 514.050 272.400 ;
        RECT 526.950 271.950 529.050 272.400 ;
        RECT 592.950 273.600 595.050 274.050 ;
        RECT 697.950 273.600 700.050 274.050 ;
        RECT 709.950 273.600 712.050 274.050 ;
        RECT 592.950 272.400 597.600 273.600 ;
        RECT 592.950 271.950 595.050 272.400 ;
        RECT 427.950 270.600 430.050 271.050 ;
        RECT 419.400 269.400 430.050 270.600 ;
        RECT 415.950 267.600 418.050 268.050 ;
        RECT 419.400 267.600 420.600 269.400 ;
        RECT 427.950 268.950 430.050 269.400 ;
        RECT 433.950 270.600 436.050 271.050 ;
        RECT 442.950 270.600 445.050 271.050 ;
        RECT 433.950 269.400 445.050 270.600 ;
        RECT 433.950 268.950 436.050 269.400 ;
        RECT 442.950 268.950 445.050 269.400 ;
        RECT 499.950 268.950 502.050 271.050 ;
        RECT 505.950 270.600 508.050 271.050 ;
        RECT 514.950 270.600 517.050 271.050 ;
        RECT 505.950 269.400 517.050 270.600 ;
        RECT 505.950 268.950 508.050 269.400 ;
        RECT 514.950 268.950 517.050 269.400 ;
        RECT 577.950 270.600 580.050 271.050 ;
        RECT 586.950 270.600 589.050 271.050 ;
        RECT 577.950 269.400 589.050 270.600 ;
        RECT 577.950 268.950 580.050 269.400 ;
        RECT 586.950 268.950 589.050 269.400 ;
        RECT 592.950 268.950 595.050 271.050 ;
        RECT 596.400 270.600 597.600 272.400 ;
        RECT 697.950 272.400 712.050 273.600 ;
        RECT 697.950 271.950 700.050 272.400 ;
        RECT 709.950 271.950 712.050 272.400 ;
        RECT 631.950 270.600 634.050 271.050 ;
        RECT 596.400 269.400 609.600 270.600 ;
        RECT 415.950 266.400 420.600 267.600 ;
        RECT 430.950 267.600 433.050 268.050 ;
        RECT 436.950 267.600 439.050 268.050 ;
        RECT 430.950 266.400 439.050 267.600 ;
        RECT 415.950 265.950 418.050 266.400 ;
        RECT 430.950 265.950 433.050 266.400 ;
        RECT 436.950 265.950 439.050 266.400 ;
        RECT 457.950 267.600 460.050 268.050 ;
        RECT 460.950 267.600 463.050 268.050 ;
        RECT 463.950 267.600 466.050 268.050 ;
        RECT 457.950 266.400 466.050 267.600 ;
        RECT 500.400 267.600 501.600 268.950 ;
        RECT 505.950 267.600 508.050 268.050 ;
        RECT 500.400 266.400 508.050 267.600 ;
        RECT 457.950 265.950 460.050 266.400 ;
        RECT 460.950 265.950 463.050 266.400 ;
        RECT 463.950 265.950 466.050 266.400 ;
        RECT 505.950 265.950 508.050 266.400 ;
        RECT 565.950 267.600 568.050 268.050 ;
        RECT 571.950 267.600 574.050 268.050 ;
        RECT 565.950 266.400 574.050 267.600 ;
        RECT 565.950 265.950 568.050 266.400 ;
        RECT 571.950 265.950 574.050 266.400 ;
        RECT 580.950 267.600 583.050 268.050 ;
        RECT 593.400 267.600 594.600 268.950 ;
        RECT 580.950 266.400 594.600 267.600 ;
        RECT 595.950 267.600 598.050 268.050 ;
        RECT 604.950 267.600 607.050 268.050 ;
        RECT 595.950 266.400 607.050 267.600 ;
        RECT 580.950 265.950 583.050 266.400 ;
        RECT 595.950 265.950 598.050 266.400 ;
        RECT 604.950 265.950 607.050 266.400 ;
        RECT 608.400 265.050 609.600 269.400 ;
        RECT 617.400 269.400 634.050 270.600 ;
        RECT 617.400 268.050 618.600 269.400 ;
        RECT 631.950 268.950 634.050 269.400 ;
        RECT 637.950 268.950 640.050 271.050 ;
        RECT 643.950 270.600 646.050 271.050 ;
        RECT 652.950 270.600 655.050 271.050 ;
        RECT 667.950 270.600 670.050 271.050 ;
        RECT 643.950 269.400 655.050 270.600 ;
        RECT 643.950 268.950 646.050 269.400 ;
        RECT 652.950 268.950 655.050 269.400 ;
        RECT 659.400 269.400 670.050 270.600 ;
        RECT 616.950 265.950 619.050 268.050 ;
        RECT 418.950 264.600 421.050 265.050 ;
        RECT 407.400 263.400 421.050 264.600 ;
        RECT 373.950 262.950 376.050 263.400 ;
        RECT 385.950 262.950 388.050 263.400 ;
        RECT 418.950 262.950 421.050 263.400 ;
        RECT 421.950 264.600 424.050 265.050 ;
        RECT 424.950 264.600 427.050 265.050 ;
        RECT 454.950 264.600 457.050 265.050 ;
        RECT 421.950 263.400 457.050 264.600 ;
        RECT 421.950 262.950 424.050 263.400 ;
        RECT 424.950 262.950 427.050 263.400 ;
        RECT 454.950 262.950 457.050 263.400 ;
        RECT 535.950 264.600 538.050 265.050 ;
        RECT 559.950 264.600 562.050 265.050 ;
        RECT 535.950 263.400 562.050 264.600 ;
        RECT 535.950 262.950 538.050 263.400 ;
        RECT 559.950 262.950 562.050 263.400 ;
        RECT 562.950 264.600 565.050 265.050 ;
        RECT 571.950 264.600 574.050 265.050 ;
        RECT 604.950 264.600 607.050 265.050 ;
        RECT 562.950 263.400 607.050 264.600 ;
        RECT 562.950 262.950 565.050 263.400 ;
        RECT 571.950 262.950 574.050 263.400 ;
        RECT 604.950 262.950 607.050 263.400 ;
        RECT 607.950 262.950 610.050 265.050 ;
        RECT 634.950 264.600 637.050 265.050 ;
        RECT 638.400 264.600 639.600 268.950 ;
        RECT 649.950 267.600 652.050 268.050 ;
        RECT 659.400 267.600 660.600 269.400 ;
        RECT 667.950 268.950 670.050 269.400 ;
        RECT 649.950 266.400 660.600 267.600 ;
        RECT 661.950 267.600 664.050 268.050 ;
        RECT 673.950 267.600 676.050 268.050 ;
        RECT 661.950 266.400 676.050 267.600 ;
        RECT 649.950 265.950 652.050 266.400 ;
        RECT 661.950 265.950 664.050 266.400 ;
        RECT 673.950 265.950 676.050 266.400 ;
        RECT 685.950 267.600 688.050 268.050 ;
        RECT 700.950 267.600 703.050 268.050 ;
        RECT 685.950 266.400 703.050 267.600 ;
        RECT 685.950 265.950 688.050 266.400 ;
        RECT 700.950 265.950 703.050 266.400 ;
        RECT 658.950 264.600 661.050 265.050 ;
        RECT 634.950 263.400 661.050 264.600 ;
        RECT 634.950 262.950 637.050 263.400 ;
        RECT 658.950 262.950 661.050 263.400 ;
        RECT 136.950 261.600 139.050 262.050 ;
        RECT 116.400 260.400 139.050 261.600 ;
        RECT 1.950 258.600 4.050 259.050 ;
        RECT 19.950 258.600 22.050 259.050 ;
        RECT 1.950 257.400 22.050 258.600 ;
        RECT 1.950 256.950 4.050 257.400 ;
        RECT 19.950 256.950 22.050 257.400 ;
        RECT 46.950 258.600 49.050 259.050 ;
        RECT 58.950 258.600 61.050 259.050 ;
        RECT 89.400 258.600 90.600 260.400 ;
        RECT 97.950 259.950 100.050 260.400 ;
        RECT 112.950 259.950 115.050 260.400 ;
        RECT 136.950 259.950 139.050 260.400 ;
        RECT 142.950 261.600 145.050 262.050 ;
        RECT 151.950 261.600 154.050 262.050 ;
        RECT 142.950 260.400 154.050 261.600 ;
        RECT 142.950 259.950 145.050 260.400 ;
        RECT 151.950 259.950 154.050 260.400 ;
        RECT 154.950 261.600 157.050 262.050 ;
        RECT 175.950 261.600 178.050 262.050 ;
        RECT 190.950 261.600 193.050 262.050 ;
        RECT 154.950 260.400 193.050 261.600 ;
        RECT 154.950 259.950 157.050 260.400 ;
        RECT 175.950 259.950 178.050 260.400 ;
        RECT 190.950 259.950 193.050 260.400 ;
        RECT 217.950 261.600 220.050 262.050 ;
        RECT 247.950 261.600 250.050 262.050 ;
        RECT 217.950 260.400 250.050 261.600 ;
        RECT 217.950 259.950 220.050 260.400 ;
        RECT 247.950 259.950 250.050 260.400 ;
        RECT 352.950 261.600 355.050 262.050 ;
        RECT 361.950 261.600 364.050 262.050 ;
        RECT 352.950 260.400 364.050 261.600 ;
        RECT 352.950 259.950 355.050 260.400 ;
        RECT 361.950 259.950 364.050 260.400 ;
        RECT 367.950 261.600 370.050 262.050 ;
        RECT 376.950 261.600 379.050 262.050 ;
        RECT 367.950 260.400 379.050 261.600 ;
        RECT 367.950 259.950 370.050 260.400 ;
        RECT 376.950 259.950 379.050 260.400 ;
        RECT 502.950 261.600 505.050 262.050 ;
        RECT 544.950 261.600 547.050 262.050 ;
        RECT 502.950 260.400 547.050 261.600 ;
        RECT 502.950 259.950 505.050 260.400 ;
        RECT 544.950 259.950 547.050 260.400 ;
        RECT 580.950 261.600 583.050 262.050 ;
        RECT 598.950 261.600 601.050 262.050 ;
        RECT 580.950 260.400 601.050 261.600 ;
        RECT 580.950 259.950 583.050 260.400 ;
        RECT 598.950 259.950 601.050 260.400 ;
        RECT 610.950 261.600 613.050 262.050 ;
        RECT 634.950 261.600 637.050 262.050 ;
        RECT 610.950 260.400 637.050 261.600 ;
        RECT 610.950 259.950 613.050 260.400 ;
        RECT 634.950 259.950 637.050 260.400 ;
        RECT 658.950 261.600 661.050 262.050 ;
        RECT 688.950 261.600 691.050 262.050 ;
        RECT 658.950 260.400 691.050 261.600 ;
        RECT 658.950 259.950 661.050 260.400 ;
        RECT 688.950 259.950 691.050 260.400 ;
        RECT 46.950 257.400 61.050 258.600 ;
        RECT 46.950 256.950 49.050 257.400 ;
        RECT 58.950 256.950 61.050 257.400 ;
        RECT 71.400 257.400 90.600 258.600 ;
        RECT 97.950 258.600 100.050 259.050 ;
        RECT 121.950 258.600 124.050 259.050 ;
        RECT 97.950 257.400 124.050 258.600 ;
        RECT 16.950 255.600 19.050 256.050 ;
        RECT 37.950 255.600 40.050 256.050 ;
        RECT 16.950 254.400 40.050 255.600 ;
        RECT 16.950 253.950 19.050 254.400 ;
        RECT 37.950 253.950 40.050 254.400 ;
        RECT 40.950 255.600 43.050 256.050 ;
        RECT 67.950 255.600 70.050 256.050 ;
        RECT 71.400 255.600 72.600 257.400 ;
        RECT 97.950 256.950 100.050 257.400 ;
        RECT 121.950 256.950 124.050 257.400 ;
        RECT 127.950 258.600 130.050 259.050 ;
        RECT 187.950 258.600 190.050 259.050 ;
        RECT 127.950 257.400 190.050 258.600 ;
        RECT 127.950 256.950 130.050 257.400 ;
        RECT 187.950 256.950 190.050 257.400 ;
        RECT 205.950 258.600 208.050 259.050 ;
        RECT 274.950 258.600 277.050 259.050 ;
        RECT 343.950 258.600 346.050 259.050 ;
        RECT 205.950 257.400 346.050 258.600 ;
        RECT 205.950 256.950 208.050 257.400 ;
        RECT 274.950 256.950 277.050 257.400 ;
        RECT 343.950 256.950 346.050 257.400 ;
        RECT 520.950 258.600 523.050 259.050 ;
        RECT 535.950 258.600 538.050 259.050 ;
        RECT 520.950 257.400 538.050 258.600 ;
        RECT 520.950 256.950 523.050 257.400 ;
        RECT 535.950 256.950 538.050 257.400 ;
        RECT 568.950 258.600 571.050 259.050 ;
        RECT 592.950 258.600 595.050 259.050 ;
        RECT 568.950 257.400 595.050 258.600 ;
        RECT 568.950 256.950 571.050 257.400 ;
        RECT 592.950 256.950 595.050 257.400 ;
        RECT 601.950 258.600 604.050 259.050 ;
        RECT 667.950 258.600 670.050 259.050 ;
        RECT 697.950 258.600 700.050 259.050 ;
        RECT 601.950 257.400 700.050 258.600 ;
        RECT 601.950 256.950 604.050 257.400 ;
        RECT 667.950 256.950 670.050 257.400 ;
        RECT 697.950 256.950 700.050 257.400 ;
        RECT 40.950 254.400 72.600 255.600 ;
        RECT 112.950 255.600 115.050 256.050 ;
        RECT 139.950 255.600 142.050 256.050 ;
        RECT 112.950 254.400 142.050 255.600 ;
        RECT 40.950 253.950 43.050 254.400 ;
        RECT 67.950 253.950 70.050 254.400 ;
        RECT 112.950 253.950 115.050 254.400 ;
        RECT 139.950 253.950 142.050 254.400 ;
        RECT 190.950 255.600 193.050 256.050 ;
        RECT 196.950 255.600 199.050 256.050 ;
        RECT 253.950 255.600 256.050 256.050 ;
        RECT 190.950 254.400 256.050 255.600 ;
        RECT 190.950 253.950 193.050 254.400 ;
        RECT 196.950 253.950 199.050 254.400 ;
        RECT 253.950 253.950 256.050 254.400 ;
        RECT 469.950 255.600 472.050 256.050 ;
        RECT 487.950 255.600 490.050 256.050 ;
        RECT 469.950 254.400 490.050 255.600 ;
        RECT 469.950 253.950 472.050 254.400 ;
        RECT 487.950 253.950 490.050 254.400 ;
        RECT 577.950 255.600 580.050 256.050 ;
        RECT 610.950 255.600 613.050 256.050 ;
        RECT 613.950 255.600 616.050 256.050 ;
        RECT 577.950 254.400 616.050 255.600 ;
        RECT 577.950 253.950 580.050 254.400 ;
        RECT 610.950 253.950 613.050 254.400 ;
        RECT 613.950 253.950 616.050 254.400 ;
        RECT 631.950 255.600 634.050 256.050 ;
        RECT 640.950 255.600 643.050 256.050 ;
        RECT 631.950 254.400 643.050 255.600 ;
        RECT 631.950 253.950 634.050 254.400 ;
        RECT 640.950 253.950 643.050 254.400 ;
        RECT 649.950 255.600 652.050 256.050 ;
        RECT 670.950 255.600 673.050 256.050 ;
        RECT 649.950 254.400 673.050 255.600 ;
        RECT 649.950 253.950 652.050 254.400 ;
        RECT 670.950 253.950 673.050 254.400 ;
        RECT 19.950 252.600 22.050 253.050 ;
        RECT 145.950 252.600 148.050 253.050 ;
        RECT 19.950 251.400 148.050 252.600 ;
        RECT 19.950 250.950 22.050 251.400 ;
        RECT 145.950 250.950 148.050 251.400 ;
        RECT 187.950 252.600 190.050 253.050 ;
        RECT 193.950 252.600 196.050 253.050 ;
        RECT 241.950 252.600 244.050 253.050 ;
        RECT 187.950 251.400 196.050 252.600 ;
        RECT 187.950 250.950 190.050 251.400 ;
        RECT 193.950 250.950 196.050 251.400 ;
        RECT 200.400 251.400 244.050 252.600 ;
        RECT 52.950 249.600 55.050 250.050 ;
        RECT 94.950 249.600 97.050 250.050 ;
        RECT 52.950 248.400 97.050 249.600 ;
        RECT 52.950 247.950 55.050 248.400 ;
        RECT 94.950 247.950 97.050 248.400 ;
        RECT 169.950 249.600 172.050 250.050 ;
        RECT 200.400 249.600 201.600 251.400 ;
        RECT 241.950 250.950 244.050 251.400 ;
        RECT 370.950 252.600 373.050 253.050 ;
        RECT 382.950 252.600 385.050 253.050 ;
        RECT 370.950 251.400 385.050 252.600 ;
        RECT 370.950 250.950 373.050 251.400 ;
        RECT 382.950 250.950 385.050 251.400 ;
        RECT 415.950 252.600 418.050 253.050 ;
        RECT 424.950 252.600 427.050 253.050 ;
        RECT 415.950 251.400 427.050 252.600 ;
        RECT 415.950 250.950 418.050 251.400 ;
        RECT 424.950 250.950 427.050 251.400 ;
        RECT 541.950 252.600 544.050 253.050 ;
        RECT 568.950 252.600 571.050 253.050 ;
        RECT 541.950 251.400 571.050 252.600 ;
        RECT 541.950 250.950 544.050 251.400 ;
        RECT 568.950 250.950 571.050 251.400 ;
        RECT 583.950 252.600 586.050 253.050 ;
        RECT 643.950 252.600 646.050 253.050 ;
        RECT 583.950 251.400 646.050 252.600 ;
        RECT 583.950 250.950 586.050 251.400 ;
        RECT 643.950 250.950 646.050 251.400 ;
        RECT 661.950 252.600 664.050 253.050 ;
        RECT 697.950 252.600 700.050 253.050 ;
        RECT 661.950 251.400 700.050 252.600 ;
        RECT 661.950 250.950 664.050 251.400 ;
        RECT 697.950 250.950 700.050 251.400 ;
        RECT 169.950 248.400 201.600 249.600 ;
        RECT 202.950 249.600 205.050 250.050 ;
        RECT 277.950 249.600 280.050 250.050 ;
        RECT 202.950 248.400 280.050 249.600 ;
        RECT 169.950 247.950 172.050 248.400 ;
        RECT 202.950 247.950 205.050 248.400 ;
        RECT 277.950 247.950 280.050 248.400 ;
        RECT 382.950 249.600 385.050 250.050 ;
        RECT 499.950 249.600 502.050 250.050 ;
        RECT 382.950 248.400 502.050 249.600 ;
        RECT 382.950 247.950 385.050 248.400 ;
        RECT 499.950 247.950 502.050 248.400 ;
        RECT 574.950 249.600 577.050 250.050 ;
        RECT 583.950 249.600 586.050 250.050 ;
        RECT 574.950 248.400 586.050 249.600 ;
        RECT 574.950 247.950 577.050 248.400 ;
        RECT 583.950 247.950 586.050 248.400 ;
        RECT 607.950 249.600 610.050 250.050 ;
        RECT 613.950 249.600 616.050 250.050 ;
        RECT 607.950 248.400 616.050 249.600 ;
        RECT 607.950 247.950 610.050 248.400 ;
        RECT 613.950 247.950 616.050 248.400 ;
        RECT 616.950 249.600 619.050 250.050 ;
        RECT 622.950 249.600 625.050 250.050 ;
        RECT 640.950 249.600 643.050 250.050 ;
        RECT 616.950 248.400 643.050 249.600 ;
        RECT 616.950 247.950 619.050 248.400 ;
        RECT 622.950 247.950 625.050 248.400 ;
        RECT 640.950 247.950 643.050 248.400 ;
        RECT 646.950 249.600 649.050 250.050 ;
        RECT 661.950 249.600 664.050 250.050 ;
        RECT 646.950 248.400 664.050 249.600 ;
        RECT 646.950 247.950 649.050 248.400 ;
        RECT 661.950 247.950 664.050 248.400 ;
        RECT 664.950 249.600 667.050 250.050 ;
        RECT 679.950 249.600 682.050 250.050 ;
        RECT 664.950 248.400 682.050 249.600 ;
        RECT 664.950 247.950 667.050 248.400 ;
        RECT 679.950 247.950 682.050 248.400 ;
        RECT 40.950 246.600 43.050 247.050 ;
        RECT 61.950 246.600 64.050 247.050 ;
        RECT 40.950 245.400 64.050 246.600 ;
        RECT 40.950 244.950 43.050 245.400 ;
        RECT 61.950 244.950 64.050 245.400 ;
        RECT 73.950 246.600 76.050 247.050 ;
        RECT 85.950 246.600 88.050 247.050 ;
        RECT 88.950 246.600 91.050 247.050 ;
        RECT 73.950 245.400 91.050 246.600 ;
        RECT 73.950 244.950 76.050 245.400 ;
        RECT 85.950 244.950 88.050 245.400 ;
        RECT 88.950 244.950 91.050 245.400 ;
        RECT 106.950 246.600 109.050 247.050 ;
        RECT 115.950 246.600 118.050 247.050 ;
        RECT 106.950 245.400 118.050 246.600 ;
        RECT 106.950 244.950 109.050 245.400 ;
        RECT 115.950 244.950 118.050 245.400 ;
        RECT 136.950 246.600 139.050 247.050 ;
        RECT 148.950 246.600 151.050 247.050 ;
        RECT 136.950 245.400 151.050 246.600 ;
        RECT 136.950 244.950 139.050 245.400 ;
        RECT 148.950 244.950 151.050 245.400 ;
        RECT 166.950 246.600 169.050 247.050 ;
        RECT 220.950 246.600 223.050 247.050 ;
        RECT 229.950 246.600 232.050 247.050 ;
        RECT 235.950 246.600 238.050 247.050 ;
        RECT 166.950 245.400 238.050 246.600 ;
        RECT 166.950 244.950 169.050 245.400 ;
        RECT 220.950 244.950 223.050 245.400 ;
        RECT 229.950 244.950 232.050 245.400 ;
        RECT 235.950 244.950 238.050 245.400 ;
        RECT 292.950 246.600 295.050 247.050 ;
        RECT 304.950 246.600 307.050 247.050 ;
        RECT 292.950 245.400 307.050 246.600 ;
        RECT 292.950 244.950 295.050 245.400 ;
        RECT 304.950 244.950 307.050 245.400 ;
        RECT 322.950 246.600 325.050 247.050 ;
        RECT 352.950 246.600 355.050 247.050 ;
        RECT 322.950 245.400 355.050 246.600 ;
        RECT 322.950 244.950 325.050 245.400 ;
        RECT 352.950 244.950 355.050 245.400 ;
        RECT 364.950 246.600 367.050 247.050 ;
        RECT 391.950 246.600 394.050 247.050 ;
        RECT 400.950 246.600 403.050 247.050 ;
        RECT 406.950 246.600 409.050 247.050 ;
        RECT 364.950 245.400 409.050 246.600 ;
        RECT 364.950 244.950 367.050 245.400 ;
        RECT 391.950 244.950 394.050 245.400 ;
        RECT 400.950 244.950 403.050 245.400 ;
        RECT 406.950 244.950 409.050 245.400 ;
        RECT 412.950 246.600 415.050 247.050 ;
        RECT 439.950 246.600 442.050 247.050 ;
        RECT 412.950 245.400 442.050 246.600 ;
        RECT 412.950 244.950 415.050 245.400 ;
        RECT 13.950 243.600 16.050 244.050 ;
        RECT 19.950 243.600 22.050 244.050 ;
        RECT 25.950 243.600 28.050 244.050 ;
        RECT 13.950 242.400 18.600 243.600 ;
        RECT 13.950 241.950 16.050 242.400 ;
        RECT 1.950 240.600 4.050 241.050 ;
        RECT 13.950 240.600 16.050 241.050 ;
        RECT 1.950 239.400 16.050 240.600 ;
        RECT 17.400 240.600 18.600 242.400 ;
        RECT 19.950 242.400 28.050 243.600 ;
        RECT 19.950 241.950 22.050 242.400 ;
        RECT 25.950 241.950 28.050 242.400 ;
        RECT 43.950 243.600 46.050 244.050 ;
        RECT 70.950 243.600 73.050 244.050 ;
        RECT 79.950 243.600 82.050 244.050 ;
        RECT 43.950 242.400 73.050 243.600 ;
        RECT 43.950 241.950 46.050 242.400 ;
        RECT 70.950 241.950 73.050 242.400 ;
        RECT 74.400 242.400 82.050 243.600 ;
        RECT 55.950 240.600 58.050 241.050 ;
        RECT 17.400 239.400 21.600 240.600 ;
        RECT 1.950 238.950 4.050 239.400 ;
        RECT 13.950 238.950 16.050 239.400 ;
        RECT 20.400 238.050 21.600 239.400 ;
        RECT 55.950 239.400 63.600 240.600 ;
        RECT 55.950 238.950 58.050 239.400 ;
        RECT 62.400 238.050 63.600 239.400 ;
        RECT 64.950 238.950 67.050 241.050 ;
        RECT 74.400 240.600 75.600 242.400 ;
        RECT 79.950 241.950 82.050 242.400 ;
        RECT 94.950 243.600 97.050 244.050 ;
        RECT 106.950 243.600 109.050 244.050 ;
        RECT 94.950 242.400 109.050 243.600 ;
        RECT 94.950 241.950 97.050 242.400 ;
        RECT 106.950 241.950 109.050 242.400 ;
        RECT 121.950 243.600 124.050 244.050 ;
        RECT 136.950 243.600 139.050 244.050 ;
        RECT 121.950 242.400 139.050 243.600 ;
        RECT 121.950 241.950 124.050 242.400 ;
        RECT 136.950 241.950 139.050 242.400 ;
        RECT 142.950 243.600 145.050 244.050 ;
        RECT 142.950 242.400 174.600 243.600 ;
        RECT 142.950 241.950 145.050 242.400 ;
        RECT 97.950 240.600 100.050 241.050 ;
        RECT 71.400 239.400 75.600 240.600 ;
        RECT 89.400 239.400 100.050 240.600 ;
        RECT 4.950 237.600 7.050 238.050 ;
        RECT 16.950 237.600 19.050 238.050 ;
        RECT 4.950 236.400 19.050 237.600 ;
        RECT 4.950 235.950 7.050 236.400 ;
        RECT 16.950 235.950 19.050 236.400 ;
        RECT 19.950 235.950 22.050 238.050 ;
        RECT 22.950 237.600 25.050 238.050 ;
        RECT 31.950 237.600 34.050 238.050 ;
        RECT 43.950 237.600 46.050 238.050 ;
        RECT 55.950 237.600 58.050 238.050 ;
        RECT 22.950 236.400 58.050 237.600 ;
        RECT 22.950 235.950 25.050 236.400 ;
        RECT 31.950 235.950 34.050 236.400 ;
        RECT 43.950 235.950 46.050 236.400 ;
        RECT 55.950 235.950 58.050 236.400 ;
        RECT 61.950 235.950 64.050 238.050 ;
        RECT 65.400 235.050 66.600 238.950 ;
        RECT 71.400 237.600 72.600 239.400 ;
        RECT 68.400 236.400 72.600 237.600 ;
        RECT 85.950 237.600 88.050 238.050 ;
        RECT 89.400 237.600 90.600 239.400 ;
        RECT 97.950 238.950 100.050 239.400 ;
        RECT 130.950 240.600 133.050 241.050 ;
        RECT 151.950 240.600 154.050 241.050 ;
        RECT 130.950 239.400 135.600 240.600 ;
        RECT 130.950 238.950 133.050 239.400 ;
        RECT 85.950 236.400 90.600 237.600 ;
        RECT 91.950 237.600 94.050 238.050 ;
        RECT 103.950 237.600 106.050 238.050 ;
        RECT 91.950 236.400 106.050 237.600 ;
        RECT 16.950 234.600 19.050 235.050 ;
        RECT 28.950 234.600 31.050 235.050 ;
        RECT 16.950 233.400 31.050 234.600 ;
        RECT 16.950 232.950 19.050 233.400 ;
        RECT 28.950 232.950 31.050 233.400 ;
        RECT 64.950 232.950 67.050 235.050 ;
        RECT 46.950 231.600 49.050 232.050 ;
        RECT 68.400 231.600 69.600 236.400 ;
        RECT 85.950 235.950 88.050 236.400 ;
        RECT 91.950 235.950 94.050 236.400 ;
        RECT 103.950 235.950 106.050 236.400 ;
        RECT 118.950 237.600 121.050 238.050 ;
        RECT 121.950 237.600 124.050 238.050 ;
        RECT 118.950 236.400 124.050 237.600 ;
        RECT 118.950 235.950 121.050 236.400 ;
        RECT 121.950 235.950 124.050 236.400 ;
        RECT 124.950 237.600 127.050 238.050 ;
        RECT 130.950 237.600 133.050 238.050 ;
        RECT 124.950 236.400 133.050 237.600 ;
        RECT 134.400 237.600 135.600 239.400 ;
        RECT 151.950 239.400 156.600 240.600 ;
        RECT 151.950 238.950 154.050 239.400 ;
        RECT 136.950 237.600 139.050 238.050 ;
        RECT 134.400 236.400 139.050 237.600 ;
        RECT 124.950 235.950 127.050 236.400 ;
        RECT 130.950 235.950 133.050 236.400 ;
        RECT 136.950 235.950 139.050 236.400 ;
        RECT 139.950 237.600 142.050 238.050 ;
        RECT 151.950 237.600 154.050 238.050 ;
        RECT 139.950 236.400 154.050 237.600 ;
        RECT 139.950 235.950 142.050 236.400 ;
        RECT 151.950 235.950 154.050 236.400 ;
        RECT 91.950 232.950 94.050 235.050 ;
        RECT 103.950 234.600 106.050 235.050 ;
        RECT 119.400 234.600 120.600 235.950 ;
        RECT 103.950 233.400 120.600 234.600 ;
        RECT 103.950 232.950 106.050 233.400 ;
        RECT 121.950 232.950 124.050 235.050 ;
        RECT 127.950 234.600 130.050 235.050 ;
        RECT 133.950 234.600 136.050 235.050 ;
        RECT 151.950 234.600 154.050 235.050 ;
        RECT 127.950 233.400 132.600 234.600 ;
        RECT 127.950 232.950 130.050 233.400 ;
        RECT 46.950 230.400 69.600 231.600 ;
        RECT 79.950 231.600 82.050 232.050 ;
        RECT 92.400 231.600 93.600 232.950 ;
        RECT 79.950 230.400 93.600 231.600 ;
        RECT 97.950 231.600 100.050 232.050 ;
        RECT 122.400 231.600 123.600 232.950 ;
        RECT 131.400 231.600 132.600 233.400 ;
        RECT 133.950 233.400 154.050 234.600 ;
        RECT 133.950 232.950 136.050 233.400 ;
        RECT 151.950 232.950 154.050 233.400 ;
        RECT 155.400 232.050 156.600 239.400 ;
        RECT 173.400 238.050 174.600 242.400 ;
        RECT 196.950 241.950 199.050 244.050 ;
        RECT 199.950 243.600 202.050 244.050 ;
        RECT 205.950 243.600 208.050 244.050 ;
        RECT 199.950 242.400 208.050 243.600 ;
        RECT 199.950 241.950 202.050 242.400 ;
        RECT 205.950 241.950 208.050 242.400 ;
        RECT 250.950 243.600 253.050 244.050 ;
        RECT 274.950 243.600 277.050 244.050 ;
        RECT 250.950 242.400 267.600 243.600 ;
        RECT 250.950 241.950 253.050 242.400 ;
        RECT 175.950 240.600 178.050 241.050 ;
        RECT 178.950 240.600 181.050 241.050 ;
        RECT 197.400 240.600 198.600 241.950 ;
        RECT 241.950 240.600 244.050 241.050 ;
        RECT 262.950 240.600 265.050 241.050 ;
        RECT 175.950 239.400 189.600 240.600 ;
        RECT 197.400 239.400 216.600 240.600 ;
        RECT 175.950 238.950 178.050 239.400 ;
        RECT 178.950 238.950 181.050 239.400 ;
        RECT 166.950 237.600 169.050 238.050 ;
        RECT 161.400 236.400 169.050 237.600 ;
        RECT 157.950 234.600 160.050 235.050 ;
        RECT 161.400 234.600 162.600 236.400 ;
        RECT 166.950 235.950 169.050 236.400 ;
        RECT 172.950 235.950 175.050 238.050 ;
        RECT 181.950 237.600 184.050 238.050 ;
        RECT 179.400 236.400 184.050 237.600 ;
        RECT 157.950 233.400 162.600 234.600 ;
        RECT 163.950 234.600 166.050 235.050 ;
        RECT 172.950 234.600 175.050 235.050 ;
        RECT 163.950 233.400 175.050 234.600 ;
        RECT 157.950 232.950 160.050 233.400 ;
        RECT 163.950 232.950 166.050 233.400 ;
        RECT 172.950 232.950 175.050 233.400 ;
        RECT 175.950 234.600 178.050 235.050 ;
        RECT 179.400 234.600 180.600 236.400 ;
        RECT 181.950 235.950 184.050 236.400 ;
        RECT 184.950 235.950 187.050 238.050 ;
        RECT 188.400 237.600 189.600 239.400 ;
        RECT 199.950 237.600 202.050 238.050 ;
        RECT 211.950 237.600 214.050 238.050 ;
        RECT 188.400 236.400 214.050 237.600 ;
        RECT 199.950 235.950 202.050 236.400 ;
        RECT 211.950 235.950 214.050 236.400 ;
        RECT 175.950 233.400 180.600 234.600 ;
        RECT 175.950 232.950 178.050 233.400 ;
        RECT 181.950 232.950 184.050 235.050 ;
        RECT 148.950 231.600 151.050 232.050 ;
        RECT 97.950 230.400 129.600 231.600 ;
        RECT 131.400 230.400 151.050 231.600 ;
        RECT 46.950 229.950 49.050 230.400 ;
        RECT 79.950 229.950 82.050 230.400 ;
        RECT 97.950 229.950 100.050 230.400 ;
        RECT 82.950 228.600 85.050 229.050 ;
        RECT 109.950 228.600 112.050 229.050 ;
        RECT 82.950 227.400 112.050 228.600 ;
        RECT 128.400 228.600 129.600 230.400 ;
        RECT 148.950 229.950 151.050 230.400 ;
        RECT 154.950 229.950 157.050 232.050 ;
        RECT 178.950 231.600 181.050 232.050 ;
        RECT 182.400 231.600 183.600 232.950 ;
        RECT 185.400 232.050 186.600 235.950 ;
        RECT 190.950 234.600 193.050 235.050 ;
        RECT 199.950 234.600 202.050 235.050 ;
        RECT 190.950 233.400 202.050 234.600 ;
        RECT 190.950 232.950 193.050 233.400 ;
        RECT 199.950 232.950 202.050 233.400 ;
        RECT 211.950 234.600 214.050 235.050 ;
        RECT 215.400 234.600 216.600 239.400 ;
        RECT 241.950 239.400 265.050 240.600 ;
        RECT 241.950 238.950 244.050 239.400 ;
        RECT 262.950 238.950 265.050 239.400 ;
        RECT 223.950 237.600 226.050 238.050 ;
        RECT 232.950 237.600 235.050 238.050 ;
        RECT 223.950 236.400 235.050 237.600 ;
        RECT 223.950 235.950 226.050 236.400 ;
        RECT 232.950 235.950 235.050 236.400 ;
        RECT 235.950 237.600 238.050 238.050 ;
        RECT 250.950 237.600 253.050 238.050 ;
        RECT 235.950 236.400 253.050 237.600 ;
        RECT 235.950 235.950 238.050 236.400 ;
        RECT 250.950 235.950 253.050 236.400 ;
        RECT 253.950 235.950 256.050 238.050 ;
        RECT 266.400 237.600 267.600 242.400 ;
        RECT 263.400 236.400 267.600 237.600 ;
        RECT 269.400 242.400 277.050 243.600 ;
        RECT 211.950 233.400 216.600 234.600 ;
        RECT 226.950 234.600 229.050 235.050 ;
        RECT 244.950 234.600 247.050 235.050 ;
        RECT 226.950 233.400 247.050 234.600 ;
        RECT 211.950 232.950 214.050 233.400 ;
        RECT 226.950 232.950 229.050 233.400 ;
        RECT 244.950 232.950 247.050 233.400 ;
        RECT 178.950 230.400 183.600 231.600 ;
        RECT 178.950 229.950 181.050 230.400 ;
        RECT 184.950 229.950 187.050 232.050 ;
        RECT 187.950 231.600 190.050 232.050 ;
        RECT 254.400 231.600 255.600 235.950 ;
        RECT 263.400 235.050 264.600 236.400 ;
        RECT 269.400 235.050 270.600 242.400 ;
        RECT 274.950 241.950 277.050 242.400 ;
        RECT 286.950 241.950 289.050 244.050 ;
        RECT 289.950 241.950 292.050 244.050 ;
        RECT 301.950 243.600 304.050 244.050 ;
        RECT 322.950 243.600 325.050 244.050 ;
        RECT 301.950 242.400 325.050 243.600 ;
        RECT 301.950 241.950 304.050 242.400 ;
        RECT 322.950 241.950 325.050 242.400 ;
        RECT 325.950 243.600 328.050 244.050 ;
        RECT 364.950 243.600 367.050 244.050 ;
        RECT 325.950 242.400 367.050 243.600 ;
        RECT 325.950 241.950 328.050 242.400 ;
        RECT 364.950 241.950 367.050 242.400 ;
        RECT 388.950 243.600 391.050 244.050 ;
        RECT 409.950 243.600 412.050 244.050 ;
        RECT 388.950 242.400 412.050 243.600 ;
        RECT 388.950 241.950 391.050 242.400 ;
        RECT 409.950 241.950 412.050 242.400 ;
        RECT 274.950 240.600 277.050 241.050 ;
        RECT 280.950 240.600 283.050 241.050 ;
        RECT 274.950 239.400 283.050 240.600 ;
        RECT 274.950 238.950 277.050 239.400 ;
        RECT 280.950 238.950 283.050 239.400 ;
        RECT 287.400 238.050 288.600 241.950 ;
        RECT 286.950 235.950 289.050 238.050 ;
        RECT 290.400 237.600 291.600 241.950 ;
        RECT 301.950 240.600 304.050 241.050 ;
        RECT 313.950 240.600 316.050 241.050 ;
        RECT 301.950 239.400 316.050 240.600 ;
        RECT 301.950 238.950 304.050 239.400 ;
        RECT 313.950 238.950 316.050 239.400 ;
        RECT 328.950 240.600 331.050 241.050 ;
        RECT 379.950 240.600 382.050 241.050 ;
        RECT 394.950 240.600 397.050 241.050 ;
        RECT 328.950 239.400 382.050 240.600 ;
        RECT 328.950 238.950 331.050 239.400 ;
        RECT 335.400 238.050 336.600 239.400 ;
        RECT 379.950 238.950 382.050 239.400 ;
        RECT 386.400 239.400 397.050 240.600 ;
        RECT 386.400 238.050 387.600 239.400 ;
        RECT 394.950 238.950 397.050 239.400 ;
        RECT 403.950 240.600 406.050 241.050 ;
        RECT 412.950 240.600 415.050 241.050 ;
        RECT 403.950 239.400 415.050 240.600 ;
        RECT 403.950 238.950 406.050 239.400 ;
        RECT 412.950 238.950 415.050 239.400 ;
        RECT 292.950 237.600 295.050 238.050 ;
        RECT 290.400 236.400 295.050 237.600 ;
        RECT 292.950 235.950 295.050 236.400 ;
        RECT 307.950 237.600 310.050 238.050 ;
        RECT 316.950 237.600 319.050 238.050 ;
        RECT 307.950 236.400 319.050 237.600 ;
        RECT 307.950 235.950 310.050 236.400 ;
        RECT 316.950 235.950 319.050 236.400 ;
        RECT 334.950 235.950 337.050 238.050 ;
        RECT 379.950 235.950 382.050 238.050 ;
        RECT 385.950 235.950 388.050 238.050 ;
        RECT 418.950 237.600 421.050 238.050 ;
        RECT 422.400 237.600 423.600 245.400 ;
        RECT 439.950 244.950 442.050 245.400 ;
        RECT 469.950 246.600 472.050 247.050 ;
        RECT 481.950 246.600 484.050 247.050 ;
        RECT 469.950 245.400 484.050 246.600 ;
        RECT 469.950 244.950 472.050 245.400 ;
        RECT 481.950 244.950 484.050 245.400 ;
        RECT 496.950 246.600 499.050 247.050 ;
        RECT 526.950 246.600 529.050 247.050 ;
        RECT 496.950 245.400 529.050 246.600 ;
        RECT 496.950 244.950 499.050 245.400 ;
        RECT 526.950 244.950 529.050 245.400 ;
        RECT 547.950 246.600 550.050 247.050 ;
        RECT 565.950 246.600 568.050 247.050 ;
        RECT 547.950 245.400 561.600 246.600 ;
        RECT 547.950 244.950 550.050 245.400 ;
        RECT 424.950 243.600 427.050 244.050 ;
        RECT 439.950 243.600 442.050 244.050 ;
        RECT 424.950 242.400 442.050 243.600 ;
        RECT 424.950 241.950 427.050 242.400 ;
        RECT 439.950 241.950 442.050 242.400 ;
        RECT 448.950 243.600 451.050 244.050 ;
        RECT 502.950 243.600 505.050 244.050 ;
        RECT 448.950 242.400 505.050 243.600 ;
        RECT 448.950 241.950 451.050 242.400 ;
        RECT 502.950 241.950 505.050 242.400 ;
        RECT 508.950 243.600 511.050 244.050 ;
        RECT 529.950 243.600 532.050 244.050 ;
        RECT 508.950 242.400 532.050 243.600 ;
        RECT 508.950 241.950 511.050 242.400 ;
        RECT 529.950 241.950 532.050 242.400 ;
        RECT 535.950 241.950 538.050 244.050 ;
        RECT 425.400 238.050 426.600 241.950 ;
        RECT 427.950 240.600 430.050 241.050 ;
        RECT 433.950 240.600 436.050 241.050 ;
        RECT 427.950 239.400 436.050 240.600 ;
        RECT 427.950 238.950 430.050 239.400 ;
        RECT 433.950 238.950 436.050 239.400 ;
        RECT 436.950 240.600 439.050 241.050 ;
        RECT 442.950 240.600 445.050 241.050 ;
        RECT 463.950 240.600 466.050 241.050 ;
        RECT 475.950 240.600 478.050 241.050 ;
        RECT 436.950 239.400 441.600 240.600 ;
        RECT 436.950 238.950 439.050 239.400 ;
        RECT 418.950 236.400 423.600 237.600 ;
        RECT 418.950 235.950 421.050 236.400 ;
        RECT 424.950 235.950 427.050 238.050 ;
        RECT 430.950 237.600 433.050 238.050 ;
        RECT 440.400 237.600 441.600 239.400 ;
        RECT 442.950 239.400 459.600 240.600 ;
        RECT 442.950 238.950 445.050 239.400 ;
        RECT 458.400 238.050 459.600 239.400 ;
        RECT 463.950 239.400 478.050 240.600 ;
        RECT 463.950 238.950 466.050 239.400 ;
        RECT 475.950 238.950 478.050 239.400 ;
        RECT 484.950 238.950 487.050 241.050 ;
        RECT 499.950 240.600 502.050 241.050 ;
        RECT 514.950 240.600 517.050 241.050 ;
        RECT 520.950 240.600 523.050 241.050 ;
        RECT 499.950 239.400 507.600 240.600 ;
        RECT 499.950 238.950 502.050 239.400 ;
        RECT 448.950 237.600 451.050 238.050 ;
        RECT 430.950 236.400 451.050 237.600 ;
        RECT 430.950 235.950 433.050 236.400 ;
        RECT 448.950 235.950 451.050 236.400 ;
        RECT 457.950 237.600 460.050 238.050 ;
        RECT 466.950 237.600 469.050 238.050 ;
        RECT 457.950 236.400 469.050 237.600 ;
        RECT 457.950 235.950 460.050 236.400 ;
        RECT 466.950 235.950 469.050 236.400 ;
        RECT 472.950 237.600 475.050 238.050 ;
        RECT 481.950 237.600 484.050 238.050 ;
        RECT 472.950 236.400 484.050 237.600 ;
        RECT 472.950 235.950 475.050 236.400 ;
        RECT 481.950 235.950 484.050 236.400 ;
        RECT 262.950 232.950 265.050 235.050 ;
        RECT 268.950 232.950 271.050 235.050 ;
        RECT 283.950 234.600 286.050 235.050 ;
        RECT 295.950 234.600 298.050 235.050 ;
        RECT 283.950 233.400 298.050 234.600 ;
        RECT 283.950 232.950 286.050 233.400 ;
        RECT 295.950 232.950 298.050 233.400 ;
        RECT 298.950 234.600 301.050 235.050 ;
        RECT 304.950 234.600 307.050 235.050 ;
        RECT 298.950 233.400 307.050 234.600 ;
        RECT 298.950 232.950 301.050 233.400 ;
        RECT 304.950 232.950 307.050 233.400 ;
        RECT 313.950 234.600 316.050 235.050 ;
        RECT 325.950 234.600 328.050 235.050 ;
        RECT 349.950 234.600 352.050 235.050 ;
        RECT 380.400 234.600 381.600 235.950 ;
        RECT 485.400 235.050 486.600 238.950 ;
        RECT 506.400 238.050 507.600 239.400 ;
        RECT 514.950 239.400 523.050 240.600 ;
        RECT 514.950 238.950 517.050 239.400 ;
        RECT 520.950 238.950 523.050 239.400 ;
        RECT 505.950 235.950 508.050 238.050 ;
        RECT 536.400 235.050 537.600 241.950 ;
        RECT 560.400 240.600 561.600 245.400 ;
        RECT 565.950 245.400 693.600 246.600 ;
        RECT 565.950 244.950 568.050 245.400 ;
        RECT 562.950 243.600 565.050 244.050 ;
        RECT 562.950 242.400 579.600 243.600 ;
        RECT 562.950 241.950 565.050 242.400 ;
        RECT 574.950 240.600 577.050 241.050 ;
        RECT 560.400 239.400 567.600 240.600 ;
        RECT 566.400 235.050 567.600 239.400 ;
        RECT 572.400 239.400 577.050 240.600 ;
        RECT 568.950 237.600 571.050 238.050 ;
        RECT 572.400 237.600 573.600 239.400 ;
        RECT 574.950 238.950 577.050 239.400 ;
        RECT 568.950 236.400 573.600 237.600 ;
        RECT 574.950 237.600 577.050 238.050 ;
        RECT 578.400 237.600 579.600 242.400 ;
        RECT 581.400 238.050 582.600 245.400 ;
        RECT 589.950 243.600 592.050 244.050 ;
        RECT 610.950 243.600 613.050 244.050 ;
        RECT 589.950 242.400 613.050 243.600 ;
        RECT 589.950 241.950 592.050 242.400 ;
        RECT 599.400 241.050 600.600 242.400 ;
        RECT 610.950 241.950 613.050 242.400 ;
        RECT 613.950 241.950 616.050 244.050 ;
        RECT 625.950 241.950 628.050 244.050 ;
        RECT 637.950 243.600 640.050 244.050 ;
        RECT 649.950 243.600 652.050 244.050 ;
        RECT 637.950 242.400 652.050 243.600 ;
        RECT 637.950 241.950 640.050 242.400 ;
        RECT 649.950 241.950 652.050 242.400 ;
        RECT 652.950 241.950 655.050 244.050 ;
        RECT 676.950 243.600 679.050 244.050 ;
        RECT 685.950 243.600 688.050 244.050 ;
        RECT 676.950 242.400 688.050 243.600 ;
        RECT 676.950 241.950 679.050 242.400 ;
        RECT 685.950 241.950 688.050 242.400 ;
        RECT 598.950 238.950 601.050 241.050 ;
        RECT 614.400 240.600 615.600 241.950 ;
        RECT 611.400 239.400 615.600 240.600 ;
        RECT 626.400 240.600 627.600 241.950 ;
        RECT 653.400 240.600 654.600 241.950 ;
        RECT 626.400 239.400 636.600 240.600 ;
        RECT 574.950 236.400 579.600 237.600 ;
        RECT 568.950 235.950 571.050 236.400 ;
        RECT 574.950 235.950 577.050 236.400 ;
        RECT 580.950 235.950 583.050 238.050 ;
        RECT 601.950 237.600 604.050 238.050 ;
        RECT 611.400 237.600 612.600 239.400 ;
        RECT 601.950 236.400 612.600 237.600 ;
        RECT 613.950 237.600 616.050 238.050 ;
        RECT 631.950 237.600 634.050 238.050 ;
        RECT 613.950 236.400 634.050 237.600 ;
        RECT 635.400 237.600 636.600 239.400 ;
        RECT 650.400 239.400 654.600 240.600 ;
        RECT 655.950 240.600 658.050 241.050 ;
        RECT 676.950 240.600 679.050 241.050 ;
        RECT 655.950 239.400 679.050 240.600 ;
        RECT 637.950 237.600 640.050 238.050 ;
        RECT 635.400 236.400 640.050 237.600 ;
        RECT 601.950 235.950 604.050 236.400 ;
        RECT 613.950 235.950 616.050 236.400 ;
        RECT 631.950 235.950 634.050 236.400 ;
        RECT 637.950 235.950 640.050 236.400 ;
        RECT 382.950 234.600 385.050 235.050 ;
        RECT 313.950 233.400 385.050 234.600 ;
        RECT 313.950 232.950 316.050 233.400 ;
        RECT 325.950 232.950 328.050 233.400 ;
        RECT 349.950 232.950 352.050 233.400 ;
        RECT 382.950 232.950 385.050 233.400 ;
        RECT 391.950 234.600 394.050 235.050 ;
        RECT 397.950 234.600 400.050 235.050 ;
        RECT 391.950 233.400 400.050 234.600 ;
        RECT 391.950 232.950 394.050 233.400 ;
        RECT 397.950 232.950 400.050 233.400 ;
        RECT 415.950 234.600 418.050 235.050 ;
        RECT 433.950 234.600 436.050 235.050 ;
        RECT 415.950 233.400 436.050 234.600 ;
        RECT 415.950 232.950 418.050 233.400 ;
        RECT 433.950 232.950 436.050 233.400 ;
        RECT 484.950 232.950 487.050 235.050 ;
        RECT 499.950 234.600 502.050 235.050 ;
        RECT 511.950 234.600 514.050 235.050 ;
        RECT 499.950 233.400 514.050 234.600 ;
        RECT 499.950 232.950 502.050 233.400 ;
        RECT 511.950 232.950 514.050 233.400 ;
        RECT 535.950 232.950 538.050 235.050 ;
        RECT 565.950 232.950 568.050 235.050 ;
        RECT 571.950 234.600 574.050 235.050 ;
        RECT 646.950 234.600 649.050 235.050 ;
        RECT 571.950 233.400 649.050 234.600 ;
        RECT 650.400 234.600 651.600 239.400 ;
        RECT 655.950 238.950 658.050 239.400 ;
        RECT 676.950 238.950 679.050 239.400 ;
        RECT 688.950 238.950 691.050 241.050 ;
        RECT 652.950 237.600 655.050 238.050 ;
        RECT 664.950 237.600 667.050 238.050 ;
        RECT 652.950 236.400 667.050 237.600 ;
        RECT 652.950 235.950 655.050 236.400 ;
        RECT 664.950 235.950 667.050 236.400 ;
        RECT 673.950 237.600 676.050 238.050 ;
        RECT 689.400 237.600 690.600 238.950 ;
        RECT 692.400 238.050 693.600 245.400 ;
        RECT 694.950 240.600 697.050 241.050 ;
        RECT 700.950 240.600 703.050 241.050 ;
        RECT 694.950 239.400 703.050 240.600 ;
        RECT 694.950 238.950 697.050 239.400 ;
        RECT 700.950 238.950 703.050 239.400 ;
        RECT 706.950 240.600 709.050 241.050 ;
        RECT 712.950 240.600 715.050 241.050 ;
        RECT 706.950 239.400 715.050 240.600 ;
        RECT 706.950 238.950 709.050 239.400 ;
        RECT 712.950 238.950 715.050 239.400 ;
        RECT 715.950 240.600 718.050 241.050 ;
        RECT 715.950 239.400 720.600 240.600 ;
        RECT 715.950 238.950 718.050 239.400 ;
        RECT 673.950 236.400 690.600 237.600 ;
        RECT 673.950 235.950 676.050 236.400 ;
        RECT 691.950 235.950 694.050 238.050 ;
        RECT 706.950 237.600 709.050 238.050 ;
        RECT 715.950 237.600 718.050 238.050 ;
        RECT 706.950 236.400 718.050 237.600 ;
        RECT 706.950 235.950 709.050 236.400 ;
        RECT 715.950 235.950 718.050 236.400 ;
        RECT 652.950 234.600 655.050 235.050 ;
        RECT 650.400 233.400 655.050 234.600 ;
        RECT 571.950 232.950 574.050 233.400 ;
        RECT 646.950 232.950 649.050 233.400 ;
        RECT 652.950 232.950 655.050 233.400 ;
        RECT 667.950 234.600 670.050 235.050 ;
        RECT 670.950 234.600 673.050 235.050 ;
        RECT 703.950 234.600 706.050 235.050 ;
        RECT 667.950 233.400 706.050 234.600 ;
        RECT 667.950 232.950 670.050 233.400 ;
        RECT 670.950 232.950 673.050 233.400 ;
        RECT 703.950 232.950 706.050 233.400 ;
        RECT 709.950 234.600 712.050 235.050 ;
        RECT 719.400 234.600 720.600 239.400 ;
        RECT 709.950 233.400 720.600 234.600 ;
        RECT 709.950 232.950 712.050 233.400 ;
        RECT 187.950 230.400 255.600 231.600 ;
        RECT 265.950 231.600 268.050 232.050 ;
        RECT 277.950 231.600 280.050 232.050 ;
        RECT 265.950 230.400 280.050 231.600 ;
        RECT 187.950 229.950 190.050 230.400 ;
        RECT 265.950 229.950 268.050 230.400 ;
        RECT 277.950 229.950 280.050 230.400 ;
        RECT 316.950 231.600 319.050 232.050 ;
        RECT 355.950 231.600 358.050 232.050 ;
        RECT 316.950 230.400 358.050 231.600 ;
        RECT 316.950 229.950 319.050 230.400 ;
        RECT 355.950 229.950 358.050 230.400 ;
        RECT 418.950 231.600 421.050 232.050 ;
        RECT 436.950 231.600 439.050 232.050 ;
        RECT 418.950 230.400 439.050 231.600 ;
        RECT 418.950 229.950 421.050 230.400 ;
        RECT 436.950 229.950 439.050 230.400 ;
        RECT 475.950 231.600 478.050 232.050 ;
        RECT 478.950 231.600 481.050 232.050 ;
        RECT 499.950 231.600 502.050 232.050 ;
        RECT 475.950 230.400 502.050 231.600 ;
        RECT 475.950 229.950 478.050 230.400 ;
        RECT 478.950 229.950 481.050 230.400 ;
        RECT 499.950 229.950 502.050 230.400 ;
        RECT 520.950 231.600 523.050 232.050 ;
        RECT 556.950 231.600 559.050 232.050 ;
        RECT 520.950 230.400 559.050 231.600 ;
        RECT 520.950 229.950 523.050 230.400 ;
        RECT 556.950 229.950 559.050 230.400 ;
        RECT 607.950 231.600 610.050 232.050 ;
        RECT 619.950 231.600 622.050 232.050 ;
        RECT 607.950 230.400 622.050 231.600 ;
        RECT 607.950 229.950 610.050 230.400 ;
        RECT 619.950 229.950 622.050 230.400 ;
        RECT 628.950 231.600 631.050 232.050 ;
        RECT 637.950 231.600 640.050 232.050 ;
        RECT 628.950 230.400 640.050 231.600 ;
        RECT 628.950 229.950 631.050 230.400 ;
        RECT 637.950 229.950 640.050 230.400 ;
        RECT 133.950 228.600 136.050 229.050 ;
        RECT 128.400 227.400 136.050 228.600 ;
        RECT 82.950 226.950 85.050 227.400 ;
        RECT 109.950 226.950 112.050 227.400 ;
        RECT 133.950 226.950 136.050 227.400 ;
        RECT 193.950 228.600 196.050 229.050 ;
        RECT 241.950 228.600 244.050 229.050 ;
        RECT 193.950 227.400 244.050 228.600 ;
        RECT 193.950 226.950 196.050 227.400 ;
        RECT 241.950 226.950 244.050 227.400 ;
        RECT 493.950 228.600 496.050 229.050 ;
        RECT 502.950 228.600 505.050 229.050 ;
        RECT 493.950 227.400 505.050 228.600 ;
        RECT 493.950 226.950 496.050 227.400 ;
        RECT 502.950 226.950 505.050 227.400 ;
        RECT 655.950 228.600 658.050 229.050 ;
        RECT 694.950 228.600 697.050 229.050 ;
        RECT 655.950 227.400 697.050 228.600 ;
        RECT 655.950 226.950 658.050 227.400 ;
        RECT 694.950 226.950 697.050 227.400 ;
        RECT 70.950 225.600 73.050 226.050 ;
        RECT 103.950 225.600 106.050 226.050 ;
        RECT 70.950 224.400 106.050 225.600 ;
        RECT 70.950 223.950 73.050 224.400 ;
        RECT 103.950 223.950 106.050 224.400 ;
        RECT 118.950 225.600 121.050 226.050 ;
        RECT 136.950 225.600 139.050 226.050 ;
        RECT 118.950 224.400 139.050 225.600 ;
        RECT 118.950 223.950 121.050 224.400 ;
        RECT 136.950 223.950 139.050 224.400 ;
        RECT 148.950 225.600 151.050 226.050 ;
        RECT 184.950 225.600 187.050 226.050 ;
        RECT 196.950 225.600 199.050 226.050 ;
        RECT 148.950 224.400 199.050 225.600 ;
        RECT 148.950 223.950 151.050 224.400 ;
        RECT 184.950 223.950 187.050 224.400 ;
        RECT 196.950 223.950 199.050 224.400 ;
        RECT 214.950 225.600 217.050 226.050 ;
        RECT 217.950 225.600 220.050 226.050 ;
        RECT 238.950 225.600 241.050 226.050 ;
        RECT 214.950 224.400 241.050 225.600 ;
        RECT 214.950 223.950 217.050 224.400 ;
        RECT 217.950 223.950 220.050 224.400 ;
        RECT 238.950 223.950 241.050 224.400 ;
        RECT 541.950 225.600 544.050 226.050 ;
        RECT 631.950 225.600 634.050 226.050 ;
        RECT 541.950 224.400 634.050 225.600 ;
        RECT 541.950 223.950 544.050 224.400 ;
        RECT 631.950 223.950 634.050 224.400 ;
        RECT 124.950 222.600 127.050 223.050 ;
        RECT 178.950 222.600 181.050 223.050 ;
        RECT 211.950 222.600 214.050 223.050 ;
        RECT 124.950 221.400 214.050 222.600 ;
        RECT 124.950 220.950 127.050 221.400 ;
        RECT 178.950 220.950 181.050 221.400 ;
        RECT 211.950 220.950 214.050 221.400 ;
        RECT 223.950 222.600 226.050 223.050 ;
        RECT 253.950 222.600 256.050 223.050 ;
        RECT 268.950 222.600 271.050 223.050 ;
        RECT 223.950 221.400 271.050 222.600 ;
        RECT 223.950 220.950 226.050 221.400 ;
        RECT 253.950 220.950 256.050 221.400 ;
        RECT 268.950 220.950 271.050 221.400 ;
        RECT 28.950 219.600 31.050 220.050 ;
        RECT 67.950 219.600 70.050 220.050 ;
        RECT 28.950 218.400 70.050 219.600 ;
        RECT 28.950 217.950 31.050 218.400 ;
        RECT 67.950 217.950 70.050 218.400 ;
        RECT 109.950 219.600 112.050 220.050 ;
        RECT 127.950 219.600 130.050 220.050 ;
        RECT 109.950 218.400 130.050 219.600 ;
        RECT 109.950 217.950 112.050 218.400 ;
        RECT 127.950 217.950 130.050 218.400 ;
        RECT 130.950 219.600 133.050 220.050 ;
        RECT 232.950 219.600 235.050 220.050 ;
        RECT 130.950 218.400 235.050 219.600 ;
        RECT 130.950 217.950 133.050 218.400 ;
        RECT 232.950 217.950 235.050 218.400 ;
        RECT 538.950 219.600 541.050 220.050 ;
        RECT 547.950 219.600 550.050 220.050 ;
        RECT 538.950 218.400 550.050 219.600 ;
        RECT 538.950 217.950 541.050 218.400 ;
        RECT 547.950 217.950 550.050 218.400 ;
        RECT 43.950 216.600 46.050 217.050 ;
        RECT 55.950 216.600 58.050 217.050 ;
        RECT 154.950 216.600 157.050 217.050 ;
        RECT 43.950 215.400 157.050 216.600 ;
        RECT 43.950 214.950 46.050 215.400 ;
        RECT 55.950 214.950 58.050 215.400 ;
        RECT 154.950 214.950 157.050 215.400 ;
        RECT 175.950 216.600 178.050 217.050 ;
        RECT 226.950 216.600 229.050 217.050 ;
        RECT 175.950 215.400 229.050 216.600 ;
        RECT 175.950 214.950 178.050 215.400 ;
        RECT 226.950 214.950 229.050 215.400 ;
        RECT 52.950 213.600 55.050 214.050 ;
        RECT 61.950 213.600 64.050 214.050 ;
        RECT 52.950 212.400 64.050 213.600 ;
        RECT 52.950 211.950 55.050 212.400 ;
        RECT 61.950 211.950 64.050 212.400 ;
        RECT 121.950 213.600 124.050 214.050 ;
        RECT 139.950 213.600 142.050 214.050 ;
        RECT 121.950 212.400 142.050 213.600 ;
        RECT 121.950 211.950 124.050 212.400 ;
        RECT 139.950 211.950 142.050 212.400 ;
        RECT 637.950 213.600 640.050 214.050 ;
        RECT 643.950 213.600 646.050 214.050 ;
        RECT 637.950 212.400 646.050 213.600 ;
        RECT 637.950 211.950 640.050 212.400 ;
        RECT 643.950 211.950 646.050 212.400 ;
        RECT 7.950 210.600 10.050 211.050 ;
        RECT 10.950 210.600 13.050 211.050 ;
        RECT 52.950 210.600 55.050 211.050 ;
        RECT 64.950 210.600 67.050 211.050 ;
        RECT 7.950 209.400 67.050 210.600 ;
        RECT 7.950 208.950 10.050 209.400 ;
        RECT 10.950 208.950 13.050 209.400 ;
        RECT 52.950 208.950 55.050 209.400 ;
        RECT 64.950 208.950 67.050 209.400 ;
        RECT 625.950 210.600 628.050 211.050 ;
        RECT 643.950 210.600 646.050 211.050 ;
        RECT 625.950 209.400 646.050 210.600 ;
        RECT 625.950 208.950 628.050 209.400 ;
        RECT 643.950 208.950 646.050 209.400 ;
        RECT 13.950 207.600 16.050 208.050 ;
        RECT 19.950 207.600 22.050 208.050 ;
        RECT 13.950 206.400 22.050 207.600 ;
        RECT 13.950 205.950 16.050 206.400 ;
        RECT 19.950 205.950 22.050 206.400 ;
        RECT 34.950 205.950 37.050 208.050 ;
        RECT 142.950 207.600 145.050 208.050 ;
        RECT 178.950 207.600 181.050 208.050 ;
        RECT 142.950 206.400 181.050 207.600 ;
        RECT 142.950 205.950 145.050 206.400 ;
        RECT 178.950 205.950 181.050 206.400 ;
        RECT 220.950 207.600 223.050 208.050 ;
        RECT 289.950 207.600 292.050 208.050 ;
        RECT 307.950 207.600 310.050 208.050 ;
        RECT 313.950 207.600 316.050 208.050 ;
        RECT 220.950 206.400 228.600 207.600 ;
        RECT 220.950 205.950 223.050 206.400 ;
        RECT 35.400 202.050 36.600 205.950 ;
        RECT 37.950 202.950 40.050 205.050 ;
        RECT 40.950 204.600 43.050 205.050 ;
        RECT 40.950 203.400 48.600 204.600 ;
        RECT 40.950 202.950 43.050 203.400 ;
        RECT 7.950 201.600 10.050 202.050 ;
        RECT 25.950 201.600 28.050 202.050 ;
        RECT 7.950 200.400 18.600 201.600 ;
        RECT 7.950 199.950 10.050 200.400 ;
        RECT 17.400 199.050 18.600 200.400 ;
        RECT 25.950 200.400 33.600 201.600 ;
        RECT 25.950 199.950 28.050 200.400 ;
        RECT 13.950 196.950 16.050 199.050 ;
        RECT 16.950 196.950 19.050 199.050 ;
        RECT 32.400 198.600 33.600 200.400 ;
        RECT 34.950 199.950 37.050 202.050 ;
        RECT 38.400 201.600 39.600 202.950 ;
        RECT 38.400 200.400 42.600 201.600 ;
        RECT 37.950 198.600 40.050 199.050 ;
        RECT 32.400 197.400 40.050 198.600 ;
        RECT 37.950 196.950 40.050 197.400 ;
        RECT 14.400 195.600 15.600 196.950 ;
        RECT 22.950 195.600 25.050 196.050 ;
        RECT 14.400 194.400 25.050 195.600 ;
        RECT 22.950 193.950 25.050 194.400 ;
        RECT 25.950 195.600 28.050 196.050 ;
        RECT 41.400 195.600 42.600 200.400 ;
        RECT 47.400 198.600 48.600 203.400 ;
        RECT 52.950 202.950 55.050 205.050 ;
        RECT 124.950 204.600 127.050 205.050 ;
        RECT 116.400 203.400 127.050 204.600 ;
        RECT 53.400 199.050 54.600 202.950 ;
        RECT 61.950 201.600 64.050 202.050 ;
        RECT 109.950 201.600 112.050 202.050 ;
        RECT 61.950 200.400 75.600 201.600 ;
        RECT 61.950 199.950 64.050 200.400 ;
        RECT 74.400 199.050 75.600 200.400 ;
        RECT 104.400 200.400 112.050 201.600 ;
        RECT 47.400 197.400 51.600 198.600 ;
        RECT 50.400 196.050 51.600 197.400 ;
        RECT 52.950 196.950 55.050 199.050 ;
        RECT 61.950 196.950 64.050 199.050 ;
        RECT 73.950 196.950 76.050 199.050 ;
        RECT 79.950 196.950 82.050 199.050 ;
        RECT 91.950 198.600 94.050 199.050 ;
        RECT 97.950 198.600 100.050 199.050 ;
        RECT 104.400 198.600 105.600 200.400 ;
        RECT 109.950 199.950 112.050 200.400 ;
        RECT 91.950 197.400 96.600 198.600 ;
        RECT 91.950 196.950 94.050 197.400 ;
        RECT 25.950 194.400 42.600 195.600 ;
        RECT 25.950 193.950 28.050 194.400 ;
        RECT 49.950 193.950 52.050 196.050 ;
        RECT 10.950 192.600 13.050 193.050 ;
        RECT 19.950 192.600 22.050 193.050 ;
        RECT 46.950 192.600 49.050 193.050 ;
        RECT 10.950 191.400 49.050 192.600 ;
        RECT 10.950 190.950 13.050 191.400 ;
        RECT 19.950 190.950 22.050 191.400 ;
        RECT 46.950 190.950 49.050 191.400 ;
        RECT 52.950 192.600 55.050 193.050 ;
        RECT 62.400 192.600 63.600 196.950 ;
        RECT 74.400 195.600 75.600 196.950 ;
        RECT 52.950 191.400 63.600 192.600 ;
        RECT 71.400 194.400 75.600 195.600 ;
        RECT 80.400 195.600 81.600 196.950 ;
        RECT 95.400 195.600 96.600 197.400 ;
        RECT 97.950 197.400 105.600 198.600 ;
        RECT 97.950 196.950 100.050 197.400 ;
        RECT 106.950 196.950 109.050 199.050 ;
        RECT 107.400 195.600 108.600 196.950 ;
        RECT 80.400 194.400 93.600 195.600 ;
        RECT 95.400 194.400 108.600 195.600 ;
        RECT 52.950 190.950 55.050 191.400 ;
        RECT 7.950 189.600 10.050 190.050 ;
        RECT 71.400 189.600 72.600 194.400 ;
        RECT 92.400 193.050 93.600 194.400 ;
        RECT 107.400 193.050 108.600 194.400 ;
        RECT 109.950 195.600 112.050 196.050 ;
        RECT 116.400 195.600 117.600 203.400 ;
        RECT 124.950 202.950 127.050 203.400 ;
        RECT 133.950 204.600 136.050 205.050 ;
        RECT 145.950 204.600 148.050 205.050 ;
        RECT 133.950 203.400 148.050 204.600 ;
        RECT 133.950 202.950 136.050 203.400 ;
        RECT 145.950 202.950 148.050 203.400 ;
        RECT 163.950 204.600 166.050 205.050 ;
        RECT 181.950 204.600 184.050 205.050 ;
        RECT 205.950 204.600 208.050 205.050 ;
        RECT 163.950 203.400 180.600 204.600 ;
        RECT 163.950 202.950 166.050 203.400 ;
        RECT 118.950 199.950 121.050 202.050 ;
        RECT 136.950 199.950 139.050 202.050 ;
        RECT 145.950 199.950 148.050 202.050 ;
        RECT 151.950 201.600 154.050 202.050 ;
        RECT 154.950 201.600 157.050 202.050 ;
        RECT 160.950 201.600 163.050 202.050 ;
        RECT 151.950 200.400 163.050 201.600 ;
        RECT 151.950 199.950 154.050 200.400 ;
        RECT 154.950 199.950 157.050 200.400 ;
        RECT 160.950 199.950 163.050 200.400 ;
        RECT 166.950 201.600 169.050 202.050 ;
        RECT 175.950 201.600 178.050 202.050 ;
        RECT 166.950 200.400 178.050 201.600 ;
        RECT 179.400 201.600 180.600 203.400 ;
        RECT 181.950 203.400 208.050 204.600 ;
        RECT 181.950 202.950 184.050 203.400 ;
        RECT 205.950 202.950 208.050 203.400 ;
        RECT 208.950 204.600 211.050 205.050 ;
        RECT 223.950 204.600 226.050 205.050 ;
        RECT 208.950 203.400 226.050 204.600 ;
        RECT 227.400 204.600 228.600 206.400 ;
        RECT 289.950 206.400 316.050 207.600 ;
        RECT 289.950 205.950 292.050 206.400 ;
        RECT 307.950 205.950 310.050 206.400 ;
        RECT 313.950 205.950 316.050 206.400 ;
        RECT 487.950 207.600 490.050 208.050 ;
        RECT 493.950 207.600 496.050 208.050 ;
        RECT 487.950 206.400 496.050 207.600 ;
        RECT 487.950 205.950 490.050 206.400 ;
        RECT 493.950 205.950 496.050 206.400 ;
        RECT 625.950 207.600 628.050 208.050 ;
        RECT 658.950 207.600 661.050 208.050 ;
        RECT 625.950 206.400 661.050 207.600 ;
        RECT 625.950 205.950 628.050 206.400 ;
        RECT 658.950 205.950 661.050 206.400 ;
        RECT 250.950 204.600 253.050 205.050 ;
        RECT 286.950 204.600 289.050 205.050 ;
        RECT 397.950 204.600 400.050 205.050 ;
        RECT 227.400 203.400 231.600 204.600 ;
        RECT 208.950 202.950 211.050 203.400 ;
        RECT 223.950 202.950 226.050 203.400 ;
        RECT 190.950 201.600 193.050 202.050 ;
        RECT 179.400 200.400 183.600 201.600 ;
        RECT 166.950 199.950 169.050 200.400 ;
        RECT 175.950 199.950 178.050 200.400 ;
        RECT 119.400 196.050 120.600 199.950 ;
        RECT 137.400 196.050 138.600 199.950 ;
        RECT 139.950 198.600 142.050 199.050 ;
        RECT 146.400 198.600 147.600 199.950 ;
        RECT 163.950 198.600 166.050 199.050 ;
        RECT 139.950 197.400 166.050 198.600 ;
        RECT 139.950 196.950 142.050 197.400 ;
        RECT 163.950 196.950 166.050 197.400 ;
        RECT 166.950 198.600 169.050 199.050 ;
        RECT 178.950 198.600 181.050 199.050 ;
        RECT 166.950 197.400 181.050 198.600 ;
        RECT 166.950 196.950 169.050 197.400 ;
        RECT 178.950 196.950 181.050 197.400 ;
        RECT 109.950 194.400 117.600 195.600 ;
        RECT 109.950 193.950 112.050 194.400 ;
        RECT 118.950 193.950 121.050 196.050 ;
        RECT 136.950 193.950 139.050 196.050 ;
        RECT 163.950 195.600 166.050 196.050 ;
        RECT 172.950 195.600 175.050 196.050 ;
        RECT 163.950 194.400 175.050 195.600 ;
        RECT 163.950 193.950 166.050 194.400 ;
        RECT 172.950 193.950 175.050 194.400 ;
        RECT 82.950 192.600 85.050 193.050 ;
        RECT 88.950 192.600 91.050 193.050 ;
        RECT 82.950 191.400 91.050 192.600 ;
        RECT 82.950 190.950 85.050 191.400 ;
        RECT 88.950 190.950 91.050 191.400 ;
        RECT 91.950 190.950 94.050 193.050 ;
        RECT 106.950 190.950 109.050 193.050 ;
        RECT 112.950 192.600 115.050 193.050 ;
        RECT 121.950 192.600 124.050 193.050 ;
        RECT 112.950 191.400 124.050 192.600 ;
        RECT 112.950 190.950 115.050 191.400 ;
        RECT 121.950 190.950 124.050 191.400 ;
        RECT 127.950 192.600 130.050 193.050 ;
        RECT 136.950 192.600 139.050 193.050 ;
        RECT 127.950 191.400 139.050 192.600 ;
        RECT 127.950 190.950 130.050 191.400 ;
        RECT 136.950 190.950 139.050 191.400 ;
        RECT 148.950 192.600 151.050 193.050 ;
        RECT 182.400 192.600 183.600 200.400 ;
        RECT 190.950 200.400 204.600 201.600 ;
        RECT 190.950 199.950 193.050 200.400 ;
        RECT 199.950 198.600 202.050 199.050 ;
        RECT 191.400 197.400 202.050 198.600 ;
        RECT 203.400 198.600 204.600 200.400 ;
        RECT 217.950 199.950 220.050 202.050 ;
        RECT 226.950 201.600 229.050 202.050 ;
        RECT 221.400 200.400 229.050 201.600 ;
        RECT 214.950 198.600 217.050 199.050 ;
        RECT 203.400 197.400 217.050 198.600 ;
        RECT 187.950 195.600 190.050 196.050 ;
        RECT 191.400 195.600 192.600 197.400 ;
        RECT 199.950 196.950 202.050 197.400 ;
        RECT 214.950 196.950 217.050 197.400 ;
        RECT 218.400 196.050 219.600 199.950 ;
        RECT 187.950 194.400 192.600 195.600 ;
        RECT 193.950 195.600 196.050 196.050 ;
        RECT 193.950 194.400 201.600 195.600 ;
        RECT 187.950 193.950 190.050 194.400 ;
        RECT 193.950 193.950 196.050 194.400 ;
        RECT 196.950 192.600 199.050 193.050 ;
        RECT 148.950 191.400 183.600 192.600 ;
        RECT 185.400 191.400 199.050 192.600 ;
        RECT 200.400 192.600 201.600 194.400 ;
        RECT 217.950 193.950 220.050 196.050 ;
        RECT 221.400 192.600 222.600 200.400 ;
        RECT 226.950 199.950 229.050 200.400 ;
        RECT 230.400 199.050 231.600 203.400 ;
        RECT 250.950 203.400 327.600 204.600 ;
        RECT 250.950 202.950 253.050 203.400 ;
        RECT 286.950 202.950 289.050 203.400 ;
        RECT 262.950 201.600 265.050 202.050 ;
        RECT 239.400 200.400 265.050 201.600 ;
        RECT 229.950 196.950 232.050 199.050 ;
        RECT 239.400 196.050 240.600 200.400 ;
        RECT 262.950 199.950 265.050 200.400 ;
        RECT 289.950 201.600 292.050 202.050 ;
        RECT 298.950 201.600 301.050 202.050 ;
        RECT 289.950 200.400 303.600 201.600 ;
        RECT 289.950 199.950 292.050 200.400 ;
        RECT 298.950 199.950 301.050 200.400 ;
        RECT 241.950 196.950 244.050 199.050 ;
        RECT 265.950 198.600 268.050 199.050 ;
        RECT 271.950 198.600 274.050 199.050 ;
        RECT 286.950 198.600 289.050 199.050 ;
        RECT 265.950 197.400 270.600 198.600 ;
        RECT 265.950 196.950 268.050 197.400 ;
        RECT 238.950 193.950 241.050 196.050 ;
        RECT 242.400 195.600 243.600 196.950 ;
        RECT 253.950 195.600 256.050 196.050 ;
        RECT 242.400 194.400 256.050 195.600 ;
        RECT 269.400 195.600 270.600 197.400 ;
        RECT 271.950 197.400 289.050 198.600 ;
        RECT 271.950 196.950 274.050 197.400 ;
        RECT 286.950 196.950 289.050 197.400 ;
        RECT 298.950 196.950 301.050 199.050 ;
        RECT 302.400 198.600 303.600 200.400 ;
        RECT 326.400 199.050 327.600 203.400 ;
        RECT 368.400 203.400 400.050 204.600 ;
        RECT 328.950 201.600 331.050 202.050 ;
        RECT 340.950 201.600 343.050 202.050 ;
        RECT 328.950 200.400 343.050 201.600 ;
        RECT 328.950 199.950 331.050 200.400 ;
        RECT 340.950 199.950 343.050 200.400 ;
        RECT 352.950 201.600 355.050 202.050 ;
        RECT 364.950 201.600 367.050 202.050 ;
        RECT 368.400 201.600 369.600 203.400 ;
        RECT 397.950 202.950 400.050 203.400 ;
        RECT 445.950 204.600 448.050 205.050 ;
        RECT 475.950 204.600 478.050 205.050 ;
        RECT 487.950 204.600 490.050 205.050 ;
        RECT 445.950 203.400 490.050 204.600 ;
        RECT 445.950 202.950 448.050 203.400 ;
        RECT 475.950 202.950 478.050 203.400 ;
        RECT 487.950 202.950 490.050 203.400 ;
        RECT 619.950 204.600 622.050 205.050 ;
        RECT 631.950 204.600 634.050 205.050 ;
        RECT 670.950 204.600 673.050 205.050 ;
        RECT 619.950 203.400 673.050 204.600 ;
        RECT 619.950 202.950 622.050 203.400 ;
        RECT 631.950 202.950 634.050 203.400 ;
        RECT 670.950 202.950 673.050 203.400 ;
        RECT 694.950 204.600 697.050 205.050 ;
        RECT 700.950 204.600 703.050 205.050 ;
        RECT 694.950 203.400 703.050 204.600 ;
        RECT 694.950 202.950 697.050 203.400 ;
        RECT 700.950 202.950 703.050 203.400 ;
        RECT 703.950 204.600 706.050 205.050 ;
        RECT 715.950 204.600 718.050 205.050 ;
        RECT 703.950 203.400 718.050 204.600 ;
        RECT 703.950 202.950 706.050 203.400 ;
        RECT 715.950 202.950 718.050 203.400 ;
        RECT 352.950 200.400 369.600 201.600 ;
        RECT 370.950 201.600 373.050 202.050 ;
        RECT 388.950 201.600 391.050 202.050 ;
        RECT 370.950 200.400 391.050 201.600 ;
        RECT 352.950 199.950 355.050 200.400 ;
        RECT 364.950 199.950 367.050 200.400 ;
        RECT 370.950 199.950 373.050 200.400 ;
        RECT 388.950 199.950 391.050 200.400 ;
        RECT 406.950 201.600 409.050 202.050 ;
        RECT 421.950 201.600 424.050 202.050 ;
        RECT 406.950 200.400 424.050 201.600 ;
        RECT 406.950 199.950 409.050 200.400 ;
        RECT 421.950 199.950 424.050 200.400 ;
        RECT 463.950 201.600 466.050 202.050 ;
        RECT 481.950 201.600 484.050 202.050 ;
        RECT 463.950 200.400 484.050 201.600 ;
        RECT 463.950 199.950 466.050 200.400 ;
        RECT 481.950 199.950 484.050 200.400 ;
        RECT 559.950 201.600 562.050 202.050 ;
        RECT 577.950 201.600 580.050 202.050 ;
        RECT 559.950 200.400 580.050 201.600 ;
        RECT 559.950 199.950 562.050 200.400 ;
        RECT 577.950 199.950 580.050 200.400 ;
        RECT 580.950 201.600 583.050 202.050 ;
        RECT 592.950 201.600 595.050 202.050 ;
        RECT 709.950 201.600 712.050 202.050 ;
        RECT 580.950 200.400 712.050 201.600 ;
        RECT 580.950 199.950 583.050 200.400 ;
        RECT 592.950 199.950 595.050 200.400 ;
        RECT 709.950 199.950 712.050 200.400 ;
        RECT 304.950 198.600 307.050 199.050 ;
        RECT 322.950 198.600 325.050 199.050 ;
        RECT 302.400 197.400 325.050 198.600 ;
        RECT 304.950 196.950 307.050 197.400 ;
        RECT 322.950 196.950 325.050 197.400 ;
        RECT 325.950 196.950 328.050 199.050 ;
        RECT 280.950 195.600 283.050 196.050 ;
        RECT 269.400 194.400 283.050 195.600 ;
        RECT 253.950 193.950 256.050 194.400 ;
        RECT 280.950 193.950 283.050 194.400 ;
        RECT 289.950 195.600 292.050 196.050 ;
        RECT 299.400 195.600 300.600 196.950 ;
        RECT 289.950 194.400 300.600 195.600 ;
        RECT 322.950 195.600 325.050 196.050 ;
        RECT 329.400 195.600 330.600 199.950 ;
        RECT 376.950 198.600 379.050 199.050 ;
        RECT 415.950 198.600 418.050 199.050 ;
        RECT 376.950 197.400 418.050 198.600 ;
        RECT 376.950 196.950 379.050 197.400 ;
        RECT 415.950 196.950 418.050 197.400 ;
        RECT 421.950 198.600 424.050 199.050 ;
        RECT 448.950 198.600 451.050 199.050 ;
        RECT 529.950 198.600 532.050 199.050 ;
        RECT 421.950 197.400 451.050 198.600 ;
        RECT 421.950 196.950 424.050 197.400 ;
        RECT 448.950 196.950 451.050 197.400 ;
        RECT 452.400 197.400 540.600 198.600 ;
        RECT 322.950 194.400 330.600 195.600 ;
        RECT 337.950 195.600 340.050 196.050 ;
        RECT 349.950 195.600 352.050 196.050 ;
        RECT 337.950 194.400 352.050 195.600 ;
        RECT 289.950 193.950 292.050 194.400 ;
        RECT 322.950 193.950 325.050 194.400 ;
        RECT 337.950 193.950 340.050 194.400 ;
        RECT 349.950 193.950 352.050 194.400 ;
        RECT 388.950 195.600 391.050 196.050 ;
        RECT 394.950 195.600 397.050 196.050 ;
        RECT 388.950 194.400 397.050 195.600 ;
        RECT 388.950 193.950 391.050 194.400 ;
        RECT 394.950 193.950 397.050 194.400 ;
        RECT 400.950 195.600 403.050 196.050 ;
        RECT 412.950 195.600 415.050 196.050 ;
        RECT 400.950 194.400 415.050 195.600 ;
        RECT 400.950 193.950 403.050 194.400 ;
        RECT 412.950 193.950 415.050 194.400 ;
        RECT 424.950 195.600 427.050 196.050 ;
        RECT 452.400 195.600 453.600 197.400 ;
        RECT 529.950 196.950 532.050 197.400 ;
        RECT 539.400 196.050 540.600 197.400 ;
        RECT 541.950 196.950 544.050 199.050 ;
        RECT 562.950 198.600 565.050 199.050 ;
        RECT 607.950 198.600 610.050 199.050 ;
        RECT 554.400 197.400 610.050 198.600 ;
        RECT 424.950 194.400 453.600 195.600 ;
        RECT 457.950 195.600 460.050 196.050 ;
        RECT 460.950 195.600 463.050 196.050 ;
        RECT 466.950 195.600 469.050 196.050 ;
        RECT 457.950 194.400 469.050 195.600 ;
        RECT 424.950 193.950 427.050 194.400 ;
        RECT 457.950 193.950 460.050 194.400 ;
        RECT 460.950 193.950 463.050 194.400 ;
        RECT 466.950 193.950 469.050 194.400 ;
        RECT 520.950 193.950 523.050 196.050 ;
        RECT 538.950 193.950 541.050 196.050 ;
        RECT 200.400 191.400 222.600 192.600 ;
        RECT 223.950 192.600 226.050 193.050 ;
        RECT 247.950 192.600 250.050 193.050 ;
        RECT 256.950 192.600 259.050 193.050 ;
        RECT 223.950 191.400 259.050 192.600 ;
        RECT 148.950 190.950 151.050 191.400 ;
        RECT 7.950 188.400 72.600 189.600 ;
        RECT 88.950 189.600 91.050 190.050 ;
        RECT 103.950 189.600 106.050 190.050 ;
        RECT 88.950 188.400 106.050 189.600 ;
        RECT 7.950 187.950 10.050 188.400 ;
        RECT 88.950 187.950 91.050 188.400 ;
        RECT 103.950 187.950 106.050 188.400 ;
        RECT 148.950 189.600 151.050 190.050 ;
        RECT 157.950 189.600 160.050 190.050 ;
        RECT 185.400 189.600 186.600 191.400 ;
        RECT 196.950 190.950 199.050 191.400 ;
        RECT 223.950 190.950 226.050 191.400 ;
        RECT 247.950 190.950 250.050 191.400 ;
        RECT 256.950 190.950 259.050 191.400 ;
        RECT 268.950 192.600 271.050 193.050 ;
        RECT 283.950 192.600 286.050 193.050 ;
        RECT 268.950 191.400 286.050 192.600 ;
        RECT 268.950 190.950 271.050 191.400 ;
        RECT 283.950 190.950 286.050 191.400 ;
        RECT 295.950 192.600 298.050 193.050 ;
        RECT 310.950 192.600 313.050 193.050 ;
        RECT 319.950 192.600 322.050 193.050 ;
        RECT 295.950 191.400 322.050 192.600 ;
        RECT 295.950 190.950 298.050 191.400 ;
        RECT 310.950 190.950 313.050 191.400 ;
        RECT 319.950 190.950 322.050 191.400 ;
        RECT 367.950 192.600 370.050 193.050 ;
        RECT 373.950 192.600 376.050 193.050 ;
        RECT 367.950 191.400 376.050 192.600 ;
        RECT 367.950 190.950 370.050 191.400 ;
        RECT 373.950 190.950 376.050 191.400 ;
        RECT 445.950 192.600 448.050 193.050 ;
        RECT 508.950 192.600 511.050 193.050 ;
        RECT 445.950 191.400 511.050 192.600 ;
        RECT 521.400 192.600 522.600 193.950 ;
        RECT 542.400 193.050 543.600 196.950 ;
        RECT 544.950 195.600 547.050 196.050 ;
        RECT 554.400 195.600 555.600 197.400 ;
        RECT 562.950 196.950 565.050 197.400 ;
        RECT 607.950 196.950 610.050 197.400 ;
        RECT 613.950 198.600 616.050 199.050 ;
        RECT 622.950 198.600 625.050 199.050 ;
        RECT 613.950 197.400 625.050 198.600 ;
        RECT 613.950 196.950 616.050 197.400 ;
        RECT 622.950 196.950 625.050 197.400 ;
        RECT 649.950 198.600 652.050 199.050 ;
        RECT 658.950 198.600 661.050 199.050 ;
        RECT 649.950 197.400 661.050 198.600 ;
        RECT 649.950 196.950 652.050 197.400 ;
        RECT 658.950 196.950 661.050 197.400 ;
        RECT 664.950 196.950 667.050 199.050 ;
        RECT 679.950 198.600 682.050 199.050 ;
        RECT 674.400 197.400 682.050 198.600 ;
        RECT 544.950 194.400 555.600 195.600 ;
        RECT 556.950 195.600 559.050 196.050 ;
        RECT 571.950 195.600 574.050 196.050 ;
        RECT 556.950 194.400 574.050 195.600 ;
        RECT 544.950 193.950 547.050 194.400 ;
        RECT 556.950 193.950 559.050 194.400 ;
        RECT 571.950 193.950 574.050 194.400 ;
        RECT 589.950 195.600 592.050 196.050 ;
        RECT 610.950 195.600 613.050 196.050 ;
        RECT 589.950 194.400 613.050 195.600 ;
        RECT 589.950 193.950 592.050 194.400 ;
        RECT 610.950 193.950 613.050 194.400 ;
        RECT 655.950 195.600 658.050 196.050 ;
        RECT 661.950 195.600 664.050 196.050 ;
        RECT 655.950 194.400 664.050 195.600 ;
        RECT 655.950 193.950 658.050 194.400 ;
        RECT 661.950 193.950 664.050 194.400 ;
        RECT 532.950 192.600 535.050 193.050 ;
        RECT 538.950 192.600 541.050 193.050 ;
        RECT 521.400 191.400 541.050 192.600 ;
        RECT 445.950 190.950 448.050 191.400 ;
        RECT 508.950 190.950 511.050 191.400 ;
        RECT 532.950 190.950 535.050 191.400 ;
        RECT 538.950 190.950 541.050 191.400 ;
        RECT 541.950 190.950 544.050 193.050 ;
        RECT 544.950 192.600 547.050 193.050 ;
        RECT 550.950 192.600 553.050 193.050 ;
        RECT 544.950 191.400 553.050 192.600 ;
        RECT 544.950 190.950 547.050 191.400 ;
        RECT 550.950 190.950 553.050 191.400 ;
        RECT 553.950 192.600 556.050 193.050 ;
        RECT 568.950 192.600 571.050 193.050 ;
        RECT 553.950 191.400 571.050 192.600 ;
        RECT 665.400 192.600 666.600 196.950 ;
        RECT 674.400 196.050 675.600 197.400 ;
        RECT 679.950 196.950 682.050 197.400 ;
        RECT 700.950 196.950 703.050 199.050 ;
        RECT 706.950 198.600 709.050 199.050 ;
        RECT 712.950 198.600 715.050 199.050 ;
        RECT 706.950 197.400 715.050 198.600 ;
        RECT 706.950 196.950 709.050 197.400 ;
        RECT 712.950 196.950 715.050 197.400 ;
        RECT 673.950 193.950 676.050 196.050 ;
        RECT 682.950 195.600 685.050 196.050 ;
        RECT 701.400 195.600 702.600 196.950 ;
        RECT 682.950 194.400 702.600 195.600 ;
        RECT 682.950 193.950 685.050 194.400 ;
        RECT 676.950 192.600 679.050 193.050 ;
        RECT 665.400 191.400 679.050 192.600 ;
        RECT 553.950 190.950 556.050 191.400 ;
        RECT 568.950 190.950 571.050 191.400 ;
        RECT 676.950 190.950 679.050 191.400 ;
        RECT 685.950 192.600 688.050 193.050 ;
        RECT 697.950 192.600 700.050 193.050 ;
        RECT 685.950 191.400 700.050 192.600 ;
        RECT 685.950 190.950 688.050 191.400 ;
        RECT 697.950 190.950 700.050 191.400 ;
        RECT 148.950 188.400 186.600 189.600 ;
        RECT 187.950 189.600 190.050 190.050 ;
        RECT 199.950 189.600 202.050 190.050 ;
        RECT 187.950 188.400 202.050 189.600 ;
        RECT 148.950 187.950 151.050 188.400 ;
        RECT 157.950 187.950 160.050 188.400 ;
        RECT 187.950 187.950 190.050 188.400 ;
        RECT 199.950 187.950 202.050 188.400 ;
        RECT 205.950 189.600 208.050 190.050 ;
        RECT 229.950 189.600 232.050 190.050 ;
        RECT 205.950 188.400 232.050 189.600 ;
        RECT 205.950 187.950 208.050 188.400 ;
        RECT 229.950 187.950 232.050 188.400 ;
        RECT 232.950 189.600 235.050 190.050 ;
        RECT 253.950 189.600 256.050 190.050 ;
        RECT 232.950 188.400 256.050 189.600 ;
        RECT 232.950 187.950 235.050 188.400 ;
        RECT 253.950 187.950 256.050 188.400 ;
        RECT 274.950 189.600 277.050 190.050 ;
        RECT 289.950 189.600 292.050 190.050 ;
        RECT 274.950 188.400 292.050 189.600 ;
        RECT 274.950 187.950 277.050 188.400 ;
        RECT 289.950 187.950 292.050 188.400 ;
        RECT 292.950 189.600 295.050 190.050 ;
        RECT 313.950 189.600 316.050 190.050 ;
        RECT 292.950 188.400 316.050 189.600 ;
        RECT 292.950 187.950 295.050 188.400 ;
        RECT 313.950 187.950 316.050 188.400 ;
        RECT 439.950 189.600 442.050 190.050 ;
        RECT 478.950 189.600 481.050 190.050 ;
        RECT 439.950 188.400 481.050 189.600 ;
        RECT 439.950 187.950 442.050 188.400 ;
        RECT 478.950 187.950 481.050 188.400 ;
        RECT 484.950 189.600 487.050 190.050 ;
        RECT 580.950 189.600 583.050 190.050 ;
        RECT 484.950 188.400 583.050 189.600 ;
        RECT 484.950 187.950 487.050 188.400 ;
        RECT 580.950 187.950 583.050 188.400 ;
        RECT 667.950 189.600 670.050 190.050 ;
        RECT 688.950 189.600 691.050 190.050 ;
        RECT 667.950 188.400 691.050 189.600 ;
        RECT 667.950 187.950 670.050 188.400 ;
        RECT 688.950 187.950 691.050 188.400 ;
        RECT 64.950 186.600 67.050 187.050 ;
        RECT 85.950 186.600 88.050 187.050 ;
        RECT 64.950 185.400 88.050 186.600 ;
        RECT 64.950 184.950 67.050 185.400 ;
        RECT 85.950 184.950 88.050 185.400 ;
        RECT 94.950 186.600 97.050 187.050 ;
        RECT 127.950 186.600 130.050 187.050 ;
        RECT 94.950 185.400 130.050 186.600 ;
        RECT 94.950 184.950 97.050 185.400 ;
        RECT 127.950 184.950 130.050 185.400 ;
        RECT 130.950 186.600 133.050 187.050 ;
        RECT 178.950 186.600 181.050 187.050 ;
        RECT 130.950 185.400 181.050 186.600 ;
        RECT 130.950 184.950 133.050 185.400 ;
        RECT 178.950 184.950 181.050 185.400 ;
        RECT 235.950 186.600 238.050 187.050 ;
        RECT 301.950 186.600 304.050 187.050 ;
        RECT 235.950 185.400 304.050 186.600 ;
        RECT 235.950 184.950 238.050 185.400 ;
        RECT 301.950 184.950 304.050 185.400 ;
        RECT 319.950 186.600 322.050 187.050 ;
        RECT 331.950 186.600 334.050 187.050 ;
        RECT 319.950 185.400 334.050 186.600 ;
        RECT 319.950 184.950 322.050 185.400 ;
        RECT 331.950 184.950 334.050 185.400 ;
        RECT 418.950 186.600 421.050 187.050 ;
        RECT 502.950 186.600 505.050 187.050 ;
        RECT 418.950 185.400 505.050 186.600 ;
        RECT 418.950 184.950 421.050 185.400 ;
        RECT 502.950 184.950 505.050 185.400 ;
        RECT 508.950 186.600 511.050 187.050 ;
        RECT 541.950 186.600 544.050 187.050 ;
        RECT 604.950 186.600 607.050 187.050 ;
        RECT 508.950 185.400 544.050 186.600 ;
        RECT 508.950 184.950 511.050 185.400 ;
        RECT 541.950 184.950 544.050 185.400 ;
        RECT 593.400 185.400 607.050 186.600 ;
        RECT 40.950 183.600 43.050 184.050 ;
        RECT 67.950 183.600 70.050 184.050 ;
        RECT 76.950 183.600 79.050 184.050 ;
        RECT 40.950 182.400 79.050 183.600 ;
        RECT 40.950 181.950 43.050 182.400 ;
        RECT 67.950 181.950 70.050 182.400 ;
        RECT 76.950 181.950 79.050 182.400 ;
        RECT 85.950 183.600 88.050 184.050 ;
        RECT 106.950 183.600 109.050 184.050 ;
        RECT 85.950 182.400 109.050 183.600 ;
        RECT 85.950 181.950 88.050 182.400 ;
        RECT 106.950 181.950 109.050 182.400 ;
        RECT 118.950 183.600 121.050 184.050 ;
        RECT 127.950 183.600 130.050 184.050 ;
        RECT 118.950 182.400 130.050 183.600 ;
        RECT 118.950 181.950 121.050 182.400 ;
        RECT 127.950 181.950 130.050 182.400 ;
        RECT 133.950 183.600 136.050 184.050 ;
        RECT 178.950 183.600 181.050 184.050 ;
        RECT 208.950 183.600 211.050 184.050 ;
        RECT 133.950 182.400 153.600 183.600 ;
        RECT 133.950 181.950 136.050 182.400 ;
        RECT 43.950 180.600 46.050 181.050 ;
        RECT 82.950 180.600 85.050 181.050 ;
        RECT 43.950 179.400 85.050 180.600 ;
        RECT 43.950 178.950 46.050 179.400 ;
        RECT 82.950 178.950 85.050 179.400 ;
        RECT 91.950 180.600 94.050 181.050 ;
        RECT 106.950 180.600 109.050 181.050 ;
        RECT 91.950 179.400 109.050 180.600 ;
        RECT 91.950 178.950 94.050 179.400 ;
        RECT 106.950 178.950 109.050 179.400 ;
        RECT 118.950 180.600 121.050 181.050 ;
        RECT 148.950 180.600 151.050 181.050 ;
        RECT 118.950 179.400 151.050 180.600 ;
        RECT 152.400 180.600 153.600 182.400 ;
        RECT 178.950 182.400 211.050 183.600 ;
        RECT 178.950 181.950 181.050 182.400 ;
        RECT 208.950 181.950 211.050 182.400 ;
        RECT 517.950 183.600 520.050 184.050 ;
        RECT 593.400 183.600 594.600 185.400 ;
        RECT 604.950 184.950 607.050 185.400 ;
        RECT 517.950 182.400 594.600 183.600 ;
        RECT 517.950 181.950 520.050 182.400 ;
        RECT 157.950 180.600 160.050 181.050 ;
        RECT 152.400 179.400 160.050 180.600 ;
        RECT 118.950 178.950 121.050 179.400 ;
        RECT 148.950 178.950 151.050 179.400 ;
        RECT 157.950 178.950 160.050 179.400 ;
        RECT 169.950 180.600 172.050 181.050 ;
        RECT 202.950 180.600 205.050 181.050 ;
        RECT 169.950 179.400 205.050 180.600 ;
        RECT 169.950 178.950 172.050 179.400 ;
        RECT 202.950 178.950 205.050 179.400 ;
        RECT 241.950 180.600 244.050 181.050 ;
        RECT 265.950 180.600 268.050 181.050 ;
        RECT 241.950 179.400 268.050 180.600 ;
        RECT 241.950 178.950 244.050 179.400 ;
        RECT 265.950 178.950 268.050 179.400 ;
        RECT 403.950 180.600 406.050 181.050 ;
        RECT 490.950 180.600 493.050 181.050 ;
        RECT 505.950 180.600 508.050 181.050 ;
        RECT 403.950 179.400 508.050 180.600 ;
        RECT 403.950 178.950 406.050 179.400 ;
        RECT 490.950 178.950 493.050 179.400 ;
        RECT 505.950 178.950 508.050 179.400 ;
        RECT 589.950 180.600 592.050 181.050 ;
        RECT 601.950 180.600 604.050 181.050 ;
        RECT 589.950 179.400 604.050 180.600 ;
        RECT 589.950 178.950 592.050 179.400 ;
        RECT 601.950 178.950 604.050 179.400 ;
        RECT 31.950 177.600 34.050 178.050 ;
        RECT -0.600 176.400 34.050 177.600 ;
        RECT -0.600 168.600 0.600 176.400 ;
        RECT 31.950 175.950 34.050 176.400 ;
        RECT 43.950 177.600 46.050 178.050 ;
        RECT 49.950 177.600 52.050 178.050 ;
        RECT 43.950 176.400 52.050 177.600 ;
        RECT 43.950 175.950 46.050 176.400 ;
        RECT 49.950 175.950 52.050 176.400 ;
        RECT 91.950 177.600 94.050 178.050 ;
        RECT 97.950 177.600 100.050 178.050 ;
        RECT 91.950 176.400 100.050 177.600 ;
        RECT 91.950 175.950 94.050 176.400 ;
        RECT 97.950 175.950 100.050 176.400 ;
        RECT 109.950 177.600 112.050 178.050 ;
        RECT 154.950 177.600 157.050 178.050 ;
        RECT 109.950 176.400 157.050 177.600 ;
        RECT 109.950 175.950 112.050 176.400 ;
        RECT 154.950 175.950 157.050 176.400 ;
        RECT 175.950 177.600 178.050 178.050 ;
        RECT 181.950 177.600 184.050 178.050 ;
        RECT 175.950 176.400 184.050 177.600 ;
        RECT 175.950 175.950 178.050 176.400 ;
        RECT 181.950 175.950 184.050 176.400 ;
        RECT 235.950 177.600 238.050 178.050 ;
        RECT 244.950 177.600 247.050 178.050 ;
        RECT 235.950 176.400 247.050 177.600 ;
        RECT 235.950 175.950 238.050 176.400 ;
        RECT 244.950 175.950 247.050 176.400 ;
        RECT 394.950 177.600 397.050 178.050 ;
        RECT 427.950 177.600 430.050 178.050 ;
        RECT 394.950 176.400 430.050 177.600 ;
        RECT 394.950 175.950 397.050 176.400 ;
        RECT 427.950 175.950 430.050 176.400 ;
        RECT 505.950 177.600 508.050 178.050 ;
        RECT 640.950 177.600 643.050 178.050 ;
        RECT 505.950 176.400 643.050 177.600 ;
        RECT 505.950 175.950 508.050 176.400 ;
        RECT 640.950 175.950 643.050 176.400 ;
        RECT 22.950 174.600 25.050 175.050 ;
        RECT 55.950 174.600 58.050 175.050 ;
        RECT 22.950 173.400 58.050 174.600 ;
        RECT 22.950 172.950 25.050 173.400 ;
        RECT 55.950 172.950 58.050 173.400 ;
        RECT 58.950 174.600 61.050 175.050 ;
        RECT 61.950 174.600 64.050 175.050 ;
        RECT 97.950 174.600 100.050 175.050 ;
        RECT 58.950 173.400 100.050 174.600 ;
        RECT 58.950 172.950 61.050 173.400 ;
        RECT 61.950 172.950 64.050 173.400 ;
        RECT 97.950 172.950 100.050 173.400 ;
        RECT 145.950 174.600 148.050 175.050 ;
        RECT 163.950 174.600 166.050 175.050 ;
        RECT 145.950 173.400 166.050 174.600 ;
        RECT 145.950 172.950 148.050 173.400 ;
        RECT 163.950 172.950 166.050 173.400 ;
        RECT 169.950 174.600 172.050 175.050 ;
        RECT 178.950 174.600 181.050 175.050 ;
        RECT 169.950 173.400 181.050 174.600 ;
        RECT 169.950 172.950 172.050 173.400 ;
        RECT 178.950 172.950 181.050 173.400 ;
        RECT 226.950 174.600 229.050 175.050 ;
        RECT 253.950 174.600 256.050 175.050 ;
        RECT 226.950 173.400 256.050 174.600 ;
        RECT 226.950 172.950 229.050 173.400 ;
        RECT 253.950 172.950 256.050 173.400 ;
        RECT 400.950 174.600 403.050 175.050 ;
        RECT 430.950 174.600 433.050 175.050 ;
        RECT 400.950 173.400 433.050 174.600 ;
        RECT 400.950 172.950 403.050 173.400 ;
        RECT 430.950 172.950 433.050 173.400 ;
        RECT 433.950 174.600 436.050 175.050 ;
        RECT 445.950 174.600 448.050 175.050 ;
        RECT 433.950 173.400 448.050 174.600 ;
        RECT 433.950 172.950 436.050 173.400 ;
        RECT 445.950 172.950 448.050 173.400 ;
        RECT 469.950 174.600 472.050 175.050 ;
        RECT 520.950 174.600 523.050 175.050 ;
        RECT 469.950 173.400 523.050 174.600 ;
        RECT 469.950 172.950 472.050 173.400 ;
        RECT 520.950 172.950 523.050 173.400 ;
        RECT 664.950 174.600 667.050 175.050 ;
        RECT 685.950 174.600 688.050 175.050 ;
        RECT 664.950 173.400 688.050 174.600 ;
        RECT 664.950 172.950 667.050 173.400 ;
        RECT 685.950 172.950 688.050 173.400 ;
        RECT 1.950 171.600 4.050 172.050 ;
        RECT 13.950 171.600 16.050 172.050 ;
        RECT 16.950 171.600 19.050 172.050 ;
        RECT 34.950 171.600 37.050 172.050 ;
        RECT 49.950 171.600 52.050 172.050 ;
        RECT 1.950 170.400 19.050 171.600 ;
        RECT 1.950 169.950 4.050 170.400 ;
        RECT 13.950 169.950 16.050 170.400 ;
        RECT 16.950 169.950 19.050 170.400 ;
        RECT 23.400 170.400 30.600 171.600 ;
        RECT 1.950 168.600 4.050 169.050 ;
        RECT -0.600 167.400 4.050 168.600 ;
        RECT 1.950 166.950 4.050 167.400 ;
        RECT 4.950 168.600 7.050 169.050 ;
        RECT 4.950 167.400 12.600 168.600 ;
        RECT 4.950 166.950 7.050 167.400 ;
        RECT 11.400 166.050 12.600 167.400 ;
        RECT 4.950 163.950 7.050 166.050 ;
        RECT 10.950 165.600 13.050 166.050 ;
        RECT 19.950 165.600 22.050 166.050 ;
        RECT 10.950 164.400 22.050 165.600 ;
        RECT 10.950 163.950 13.050 164.400 ;
        RECT 19.950 163.950 22.050 164.400 ;
        RECT 5.400 162.600 6.600 163.950 ;
        RECT 13.950 162.600 16.050 163.050 ;
        RECT 23.400 162.600 24.600 170.400 ;
        RECT 25.950 166.950 28.050 169.050 ;
        RECT 5.400 161.400 24.600 162.600 ;
        RECT 13.950 160.950 16.050 161.400 ;
        RECT 26.400 160.050 27.600 166.950 ;
        RECT 29.400 165.600 30.600 170.400 ;
        RECT 34.950 170.400 52.050 171.600 ;
        RECT 34.950 169.950 37.050 170.400 ;
        RECT 49.950 169.950 52.050 170.400 ;
        RECT 52.950 169.950 55.050 172.050 ;
        RECT 64.950 171.600 67.050 172.050 ;
        RECT 79.950 171.600 82.050 172.050 ;
        RECT 64.950 170.400 82.050 171.600 ;
        RECT 64.950 169.950 67.050 170.400 ;
        RECT 79.950 169.950 82.050 170.400 ;
        RECT 82.950 171.600 85.050 172.050 ;
        RECT 124.950 171.600 127.050 172.050 ;
        RECT 154.950 171.600 157.050 172.050 ;
        RECT 166.950 171.600 169.050 172.050 ;
        RECT 184.950 171.600 187.050 172.050 ;
        RECT 82.950 170.400 87.600 171.600 ;
        RECT 82.950 169.950 85.050 170.400 ;
        RECT 31.950 168.600 34.050 169.050 ;
        RECT 37.950 168.600 40.050 169.050 ;
        RECT 43.950 168.600 46.050 169.050 ;
        RECT 31.950 167.400 46.050 168.600 ;
        RECT 53.400 168.600 54.600 169.950 ;
        RECT 55.950 168.600 58.050 169.050 ;
        RECT 53.400 167.400 58.050 168.600 ;
        RECT 31.950 166.950 34.050 167.400 ;
        RECT 37.950 166.950 40.050 167.400 ;
        RECT 43.950 166.950 46.050 167.400 ;
        RECT 55.950 166.950 58.050 167.400 ;
        RECT 61.950 168.600 64.050 169.050 ;
        RECT 61.950 167.400 84.600 168.600 ;
        RECT 61.950 166.950 64.050 167.400 ;
        RECT 83.400 166.050 84.600 167.400 ;
        RECT 37.950 165.600 40.050 166.050 ;
        RECT 64.950 165.600 67.050 166.050 ;
        RECT 29.400 164.400 40.050 165.600 ;
        RECT 37.950 163.950 40.050 164.400 ;
        RECT 56.400 164.400 67.050 165.600 ;
        RECT 40.950 162.600 43.050 163.050 ;
        RECT 56.400 162.600 57.600 164.400 ;
        RECT 64.950 163.950 67.050 164.400 ;
        RECT 67.950 165.600 70.050 166.050 ;
        RECT 76.950 165.600 79.050 166.050 ;
        RECT 67.950 164.400 79.050 165.600 ;
        RECT 67.950 163.950 70.050 164.400 ;
        RECT 76.950 163.950 79.050 164.400 ;
        RECT 82.950 163.950 85.050 166.050 ;
        RECT 40.950 161.400 57.600 162.600 ;
        RECT 58.950 162.600 61.050 163.050 ;
        RECT 68.400 162.600 69.600 163.950 ;
        RECT 86.400 163.050 87.600 170.400 ;
        RECT 124.950 170.400 157.050 171.600 ;
        RECT 124.950 169.950 127.050 170.400 ;
        RECT 154.950 169.950 157.050 170.400 ;
        RECT 158.400 170.400 187.050 171.600 ;
        RECT 109.950 166.950 112.050 169.050 ;
        RECT 115.950 166.950 118.050 169.050 ;
        RECT 121.950 166.950 124.050 169.050 ;
        RECT 139.950 168.600 142.050 169.050 ;
        RECT 128.400 167.400 142.050 168.600 ;
        RECT 110.400 163.050 111.600 166.950 ;
        RECT 116.400 163.050 117.600 166.950 ;
        RECT 58.950 161.400 69.600 162.600 ;
        RECT 70.950 162.600 73.050 163.050 ;
        RECT 79.950 162.600 82.050 163.050 ;
        RECT 70.950 161.400 82.050 162.600 ;
        RECT 40.950 160.950 43.050 161.400 ;
        RECT 58.950 160.950 61.050 161.400 ;
        RECT 70.950 160.950 73.050 161.400 ;
        RECT 79.950 160.950 82.050 161.400 ;
        RECT 85.950 160.950 88.050 163.050 ;
        RECT 100.950 162.600 103.050 163.050 ;
        RECT 109.950 162.600 112.050 163.050 ;
        RECT 100.950 161.400 112.050 162.600 ;
        RECT 100.950 160.950 103.050 161.400 ;
        RECT 109.950 160.950 112.050 161.400 ;
        RECT 115.950 160.950 118.050 163.050 ;
        RECT 25.950 157.950 28.050 160.050 ;
        RECT 28.950 159.600 31.050 160.050 ;
        RECT 37.950 159.600 40.050 160.050 ;
        RECT 52.950 159.600 55.050 160.050 ;
        RECT 28.950 158.400 55.050 159.600 ;
        RECT 122.400 159.600 123.600 166.950 ;
        RECT 128.400 166.050 129.600 167.400 ;
        RECT 139.950 166.950 142.050 167.400 ;
        RECT 158.400 166.050 159.600 170.400 ;
        RECT 166.950 169.950 169.050 170.400 ;
        RECT 184.950 169.950 187.050 170.400 ;
        RECT 193.950 171.600 196.050 172.050 ;
        RECT 202.950 171.600 205.050 172.050 ;
        RECT 241.950 171.600 244.050 172.050 ;
        RECT 193.950 170.400 244.050 171.600 ;
        RECT 193.950 169.950 196.050 170.400 ;
        RECT 202.950 169.950 205.050 170.400 ;
        RECT 241.950 169.950 244.050 170.400 ;
        RECT 244.950 171.600 247.050 172.050 ;
        RECT 250.950 171.600 253.050 172.050 ;
        RECT 244.950 170.400 253.050 171.600 ;
        RECT 244.950 169.950 247.050 170.400 ;
        RECT 250.950 169.950 253.050 170.400 ;
        RECT 253.950 171.600 256.050 172.050 ;
        RECT 268.950 171.600 271.050 172.050 ;
        RECT 253.950 170.400 271.050 171.600 ;
        RECT 253.950 169.950 256.050 170.400 ;
        RECT 268.950 169.950 271.050 170.400 ;
        RECT 277.950 171.600 280.050 172.050 ;
        RECT 307.950 171.600 310.050 172.050 ;
        RECT 277.950 170.400 310.050 171.600 ;
        RECT 277.950 169.950 280.050 170.400 ;
        RECT 307.950 169.950 310.050 170.400 ;
        RECT 331.950 171.600 334.050 172.050 ;
        RECT 352.950 171.600 355.050 172.050 ;
        RECT 331.950 170.400 355.050 171.600 ;
        RECT 331.950 169.950 334.050 170.400 ;
        RECT 352.950 169.950 355.050 170.400 ;
        RECT 391.950 171.600 394.050 172.050 ;
        RECT 403.950 171.600 406.050 172.050 ;
        RECT 391.950 170.400 406.050 171.600 ;
        RECT 391.950 169.950 394.050 170.400 ;
        RECT 403.950 169.950 406.050 170.400 ;
        RECT 448.950 171.600 451.050 172.050 ;
        RECT 475.950 171.600 478.050 172.050 ;
        RECT 481.950 171.600 484.050 172.050 ;
        RECT 499.950 171.600 502.050 172.050 ;
        RECT 448.950 170.400 502.050 171.600 ;
        RECT 448.950 169.950 451.050 170.400 ;
        RECT 475.950 169.950 478.050 170.400 ;
        RECT 481.950 169.950 484.050 170.400 ;
        RECT 499.950 169.950 502.050 170.400 ;
        RECT 571.950 171.600 574.050 172.050 ;
        RECT 577.950 171.600 580.050 172.050 ;
        RECT 571.950 170.400 580.050 171.600 ;
        RECT 571.950 169.950 574.050 170.400 ;
        RECT 577.950 169.950 580.050 170.400 ;
        RECT 583.950 171.600 586.050 172.050 ;
        RECT 619.950 171.600 622.050 172.050 ;
        RECT 583.950 170.400 622.050 171.600 ;
        RECT 583.950 169.950 586.050 170.400 ;
        RECT 619.950 169.950 622.050 170.400 ;
        RECT 625.950 171.600 628.050 172.050 ;
        RECT 658.950 171.600 661.050 172.050 ;
        RECT 625.950 170.400 661.050 171.600 ;
        RECT 625.950 169.950 628.050 170.400 ;
        RECT 658.950 169.950 661.050 170.400 ;
        RECT 682.950 171.600 685.050 172.050 ;
        RECT 712.950 171.600 715.050 172.050 ;
        RECT 682.950 170.400 715.050 171.600 ;
        RECT 682.950 169.950 685.050 170.400 ;
        RECT 712.950 169.950 715.050 170.400 ;
        RECT 166.950 168.600 169.050 169.050 ;
        RECT 193.950 168.600 196.050 169.050 ;
        RECT 166.950 167.400 196.050 168.600 ;
        RECT 166.950 166.950 169.050 167.400 ;
        RECT 127.950 163.950 130.050 166.050 ;
        RECT 157.950 163.950 160.050 166.050 ;
        RECT 182.400 163.050 183.600 167.400 ;
        RECT 193.950 166.950 196.050 167.400 ;
        RECT 205.950 166.950 208.050 169.050 ;
        RECT 214.950 168.600 217.050 169.050 ;
        RECT 220.950 168.600 223.050 169.050 ;
        RECT 232.950 168.600 235.050 169.050 ;
        RECT 214.950 167.400 235.050 168.600 ;
        RECT 214.950 166.950 217.050 167.400 ;
        RECT 220.950 166.950 223.050 167.400 ;
        RECT 232.950 166.950 235.050 167.400 ;
        RECT 250.950 168.600 253.050 169.050 ;
        RECT 262.950 168.600 265.050 169.050 ;
        RECT 280.950 168.600 283.050 169.050 ;
        RECT 319.950 168.600 322.050 169.050 ;
        RECT 250.950 167.400 283.050 168.600 ;
        RECT 250.950 166.950 253.050 167.400 ;
        RECT 262.950 166.950 265.050 167.400 ;
        RECT 280.950 166.950 283.050 167.400 ;
        RECT 290.400 167.400 322.050 168.600 ;
        RECT 184.950 165.600 187.050 166.050 ;
        RECT 184.950 164.400 204.600 165.600 ;
        RECT 184.950 163.950 187.050 164.400 ;
        RECT 203.400 163.050 204.600 164.400 ;
        RECT 206.400 163.050 207.600 166.950 ;
        RECT 232.950 165.600 235.050 166.050 ;
        RECT 232.950 164.400 243.600 165.600 ;
        RECT 232.950 163.950 235.050 164.400 ;
        RECT 242.400 163.050 243.600 164.400 ;
        RECT 256.950 163.950 259.050 166.050 ;
        RECT 271.950 165.600 274.050 166.050 ;
        RECT 283.950 165.600 286.050 166.050 ;
        RECT 290.400 165.600 291.600 167.400 ;
        RECT 319.950 166.950 322.050 167.400 ;
        RECT 358.950 168.600 361.050 169.050 ;
        RECT 388.950 168.600 391.050 169.050 ;
        RECT 409.950 168.600 412.050 169.050 ;
        RECT 418.950 168.600 421.050 169.050 ;
        RECT 358.950 167.400 391.050 168.600 ;
        RECT 358.950 166.950 361.050 167.400 ;
        RECT 388.950 166.950 391.050 167.400 ;
        RECT 398.400 167.400 421.050 168.600 ;
        RECT 398.400 166.050 399.600 167.400 ;
        RECT 409.950 166.950 412.050 167.400 ;
        RECT 418.950 166.950 421.050 167.400 ;
        RECT 445.950 168.600 448.050 169.050 ;
        RECT 451.950 168.600 454.050 169.050 ;
        RECT 445.950 167.400 454.050 168.600 ;
        RECT 445.950 166.950 448.050 167.400 ;
        RECT 451.950 166.950 454.050 167.400 ;
        RECT 487.950 168.600 490.050 169.050 ;
        RECT 535.950 168.600 538.050 169.050 ;
        RECT 538.950 168.600 541.050 169.050 ;
        RECT 580.950 168.600 583.050 169.050 ;
        RECT 487.950 167.400 583.050 168.600 ;
        RECT 487.950 166.950 490.050 167.400 ;
        RECT 535.950 166.950 538.050 167.400 ;
        RECT 538.950 166.950 541.050 167.400 ;
        RECT 580.950 166.950 583.050 167.400 ;
        RECT 586.950 168.600 589.050 169.050 ;
        RECT 601.950 168.600 604.050 169.050 ;
        RECT 643.950 168.600 646.050 169.050 ;
        RECT 649.950 168.600 652.050 169.050 ;
        RECT 652.950 168.600 655.050 169.050 ;
        RECT 673.950 168.600 676.050 169.050 ;
        RECT 694.950 168.600 697.050 169.050 ;
        RECT 700.950 168.600 703.050 169.050 ;
        RECT 586.950 167.400 655.050 168.600 ;
        RECT 586.950 166.950 589.050 167.400 ;
        RECT 601.950 166.950 604.050 167.400 ;
        RECT 643.950 166.950 646.050 167.400 ;
        RECT 649.950 166.950 652.050 167.400 ;
        RECT 652.950 166.950 655.050 167.400 ;
        RECT 656.400 167.400 666.600 168.600 ;
        RECT 656.400 166.050 657.600 167.400 ;
        RECT 271.950 164.400 286.050 165.600 ;
        RECT 271.950 163.950 274.050 164.400 ;
        RECT 283.950 163.950 286.050 164.400 ;
        RECT 287.400 164.400 291.600 165.600 ;
        RECT 316.950 165.600 319.050 166.050 ;
        RECT 322.950 165.600 325.050 166.050 ;
        RECT 316.950 164.400 325.050 165.600 ;
        RECT 142.950 162.600 145.050 163.050 ;
        RECT 172.950 162.600 175.050 163.050 ;
        RECT 142.950 161.400 175.050 162.600 ;
        RECT 142.950 160.950 145.050 161.400 ;
        RECT 172.950 160.950 175.050 161.400 ;
        RECT 181.950 160.950 184.050 163.050 ;
        RECT 202.950 160.950 205.050 163.050 ;
        RECT 205.950 160.950 208.050 163.050 ;
        RECT 241.950 160.950 244.050 163.050 ;
        RECT 247.950 162.600 250.050 163.050 ;
        RECT 257.400 162.600 258.600 163.950 ;
        RECT 287.400 163.050 288.600 164.400 ;
        RECT 316.950 163.950 319.050 164.400 ;
        RECT 322.950 163.950 325.050 164.400 ;
        RECT 328.950 165.600 331.050 166.050 ;
        RECT 355.950 165.600 358.050 166.050 ;
        RECT 367.950 165.600 370.050 166.050 ;
        RECT 328.950 164.400 370.050 165.600 ;
        RECT 328.950 163.950 331.050 164.400 ;
        RECT 355.950 163.950 358.050 164.400 ;
        RECT 367.950 163.950 370.050 164.400 ;
        RECT 379.950 165.600 382.050 166.050 ;
        RECT 391.950 165.600 394.050 166.050 ;
        RECT 379.950 164.400 394.050 165.600 ;
        RECT 379.950 163.950 382.050 164.400 ;
        RECT 391.950 163.950 394.050 164.400 ;
        RECT 397.950 163.950 400.050 166.050 ;
        RECT 454.950 165.600 457.050 166.050 ;
        RECT 466.950 165.600 469.050 166.050 ;
        RECT 454.950 164.400 469.050 165.600 ;
        RECT 454.950 163.950 457.050 164.400 ;
        RECT 466.950 163.950 469.050 164.400 ;
        RECT 574.950 165.600 577.050 166.050 ;
        RECT 577.950 165.600 580.050 166.050 ;
        RECT 583.950 165.600 586.050 166.050 ;
        RECT 574.950 164.400 586.050 165.600 ;
        RECT 574.950 163.950 577.050 164.400 ;
        RECT 577.950 163.950 580.050 164.400 ;
        RECT 583.950 163.950 586.050 164.400 ;
        RECT 595.950 165.600 598.050 166.050 ;
        RECT 604.950 165.600 607.050 166.050 ;
        RECT 595.950 164.400 607.050 165.600 ;
        RECT 595.950 163.950 598.050 164.400 ;
        RECT 604.950 163.950 607.050 164.400 ;
        RECT 643.950 165.600 646.050 166.050 ;
        RECT 643.950 164.400 654.600 165.600 ;
        RECT 643.950 163.950 646.050 164.400 ;
        RECT 247.950 161.400 258.600 162.600 ;
        RECT 259.950 162.600 262.050 163.050 ;
        RECT 280.950 162.600 283.050 163.050 ;
        RECT 259.950 161.400 283.050 162.600 ;
        RECT 247.950 160.950 250.050 161.400 ;
        RECT 259.950 160.950 262.050 161.400 ;
        RECT 280.950 160.950 283.050 161.400 ;
        RECT 286.950 160.950 289.050 163.050 ;
        RECT 310.950 162.600 313.050 163.050 ;
        RECT 325.950 162.600 328.050 163.050 ;
        RECT 340.950 162.600 343.050 163.050 ;
        RECT 376.950 162.600 379.050 163.050 ;
        RECT 310.950 161.400 379.050 162.600 ;
        RECT 310.950 160.950 313.050 161.400 ;
        RECT 325.950 160.950 328.050 161.400 ;
        RECT 340.950 160.950 343.050 161.400 ;
        RECT 376.950 160.950 379.050 161.400 ;
        RECT 382.950 162.600 385.050 163.050 ;
        RECT 397.950 162.600 400.050 163.050 ;
        RECT 382.950 161.400 400.050 162.600 ;
        RECT 382.950 160.950 385.050 161.400 ;
        RECT 397.950 160.950 400.050 161.400 ;
        RECT 607.950 162.600 610.050 163.050 ;
        RECT 628.950 162.600 631.050 163.050 ;
        RECT 640.950 162.600 643.050 163.050 ;
        RECT 607.950 161.400 643.050 162.600 ;
        RECT 653.400 162.600 654.600 164.400 ;
        RECT 655.950 163.950 658.050 166.050 ;
        RECT 661.950 163.950 664.050 166.050 ;
        RECT 665.400 165.600 666.600 167.400 ;
        RECT 673.950 167.400 684.600 168.600 ;
        RECT 673.950 166.950 676.050 167.400 ;
        RECT 683.400 166.050 684.600 167.400 ;
        RECT 694.950 167.400 703.050 168.600 ;
        RECT 694.950 166.950 697.050 167.400 ;
        RECT 700.950 166.950 703.050 167.400 ;
        RECT 703.950 168.600 706.050 169.050 ;
        RECT 709.950 168.600 712.050 169.050 ;
        RECT 703.950 167.400 712.050 168.600 ;
        RECT 703.950 166.950 706.050 167.400 ;
        RECT 709.950 166.950 712.050 167.400 ;
        RECT 673.950 165.600 676.050 166.050 ;
        RECT 665.400 164.400 676.050 165.600 ;
        RECT 673.950 163.950 676.050 164.400 ;
        RECT 682.950 163.950 685.050 166.050 ;
        RECT 688.950 165.600 691.050 166.050 ;
        RECT 686.400 164.400 691.050 165.600 ;
        RECT 662.400 162.600 663.600 163.950 ;
        RECT 653.400 161.400 663.600 162.600 ;
        RECT 664.950 162.600 667.050 163.050 ;
        RECT 670.950 162.600 673.050 163.050 ;
        RECT 664.950 161.400 673.050 162.600 ;
        RECT 607.950 160.950 610.050 161.400 ;
        RECT 628.950 160.950 631.050 161.400 ;
        RECT 640.950 160.950 643.050 161.400 ;
        RECT 664.950 160.950 667.050 161.400 ;
        RECT 670.950 160.950 673.050 161.400 ;
        RECT 682.950 162.600 685.050 163.050 ;
        RECT 686.400 162.600 687.600 164.400 ;
        RECT 688.950 163.950 691.050 164.400 ;
        RECT 682.950 161.400 687.600 162.600 ;
        RECT 697.950 162.600 700.050 163.050 ;
        RECT 697.950 161.400 702.600 162.600 ;
        RECT 682.950 160.950 685.050 161.400 ;
        RECT 697.950 160.950 700.050 161.400 ;
        RECT 701.400 160.050 702.600 161.400 ;
        RECT 130.950 159.600 133.050 160.050 ;
        RECT 122.400 158.400 133.050 159.600 ;
        RECT 28.950 157.950 31.050 158.400 ;
        RECT 37.950 157.950 40.050 158.400 ;
        RECT 52.950 157.950 55.050 158.400 ;
        RECT 130.950 157.950 133.050 158.400 ;
        RECT 241.950 159.600 244.050 160.050 ;
        RECT 268.950 159.600 271.050 160.050 ;
        RECT 241.950 158.400 271.050 159.600 ;
        RECT 241.950 157.950 244.050 158.400 ;
        RECT 268.950 157.950 271.050 158.400 ;
        RECT 274.950 159.600 277.050 160.050 ;
        RECT 289.950 159.600 292.050 160.050 ;
        RECT 274.950 158.400 292.050 159.600 ;
        RECT 274.950 157.950 277.050 158.400 ;
        RECT 289.950 157.950 292.050 158.400 ;
        RECT 304.950 159.600 307.050 160.050 ;
        RECT 337.950 159.600 340.050 160.050 ;
        RECT 346.950 159.600 349.050 160.050 ;
        RECT 304.950 158.400 349.050 159.600 ;
        RECT 304.950 157.950 307.050 158.400 ;
        RECT 337.950 157.950 340.050 158.400 ;
        RECT 346.950 157.950 349.050 158.400 ;
        RECT 436.950 159.600 439.050 160.050 ;
        RECT 448.950 159.600 451.050 160.050 ;
        RECT 436.950 158.400 451.050 159.600 ;
        RECT 436.950 157.950 439.050 158.400 ;
        RECT 448.950 157.950 451.050 158.400 ;
        RECT 700.950 157.950 703.050 160.050 ;
        RECT 82.950 156.600 85.050 157.050 ;
        RECT 235.950 156.600 238.050 157.050 ;
        RECT 262.950 156.600 265.050 157.050 ;
        RECT 82.950 155.400 265.050 156.600 ;
        RECT 82.950 154.950 85.050 155.400 ;
        RECT 235.950 154.950 238.050 155.400 ;
        RECT 262.950 154.950 265.050 155.400 ;
        RECT 271.950 156.600 274.050 157.050 ;
        RECT 292.950 156.600 295.050 157.050 ;
        RECT 271.950 155.400 295.050 156.600 ;
        RECT 271.950 154.950 274.050 155.400 ;
        RECT 292.950 154.950 295.050 155.400 ;
        RECT 676.950 156.600 679.050 157.050 ;
        RECT 703.950 156.600 706.050 157.050 ;
        RECT 676.950 155.400 706.050 156.600 ;
        RECT 676.950 154.950 679.050 155.400 ;
        RECT 703.950 154.950 706.050 155.400 ;
        RECT 94.950 153.600 97.050 154.050 ;
        RECT 115.950 153.600 118.050 154.050 ;
        RECT 121.950 153.600 124.050 154.050 ;
        RECT 94.950 152.400 124.050 153.600 ;
        RECT 94.950 151.950 97.050 152.400 ;
        RECT 115.950 151.950 118.050 152.400 ;
        RECT 121.950 151.950 124.050 152.400 ;
        RECT 193.950 153.600 196.050 154.050 ;
        RECT 193.950 152.400 243.600 153.600 ;
        RECT 193.950 151.950 196.050 152.400 ;
        RECT 115.950 150.600 118.050 151.050 ;
        RECT 229.950 150.600 232.050 151.050 ;
        RECT 115.950 149.400 232.050 150.600 ;
        RECT 242.400 150.600 243.600 152.400 ;
        RECT 247.950 150.600 250.050 151.050 ;
        RECT 242.400 149.400 250.050 150.600 ;
        RECT 115.950 148.950 118.050 149.400 ;
        RECT 229.950 148.950 232.050 149.400 ;
        RECT 247.950 148.950 250.050 149.400 ;
        RECT 124.950 147.600 127.050 148.050 ;
        RECT 133.950 147.600 136.050 148.050 ;
        RECT 124.950 146.400 136.050 147.600 ;
        RECT 124.950 145.950 127.050 146.400 ;
        RECT 133.950 145.950 136.050 146.400 ;
        RECT 172.950 147.600 175.050 148.050 ;
        RECT 214.950 147.600 217.050 148.050 ;
        RECT 172.950 146.400 217.050 147.600 ;
        RECT 172.950 145.950 175.050 146.400 ;
        RECT 214.950 145.950 217.050 146.400 ;
        RECT 268.950 147.600 271.050 148.050 ;
        RECT 376.950 147.600 379.050 148.050 ;
        RECT 268.950 146.400 379.050 147.600 ;
        RECT 268.950 145.950 271.050 146.400 ;
        RECT 376.950 145.950 379.050 146.400 ;
        RECT 547.950 147.600 550.050 148.050 ;
        RECT 586.950 147.600 589.050 148.050 ;
        RECT 592.950 147.600 595.050 148.050 ;
        RECT 547.950 146.400 595.050 147.600 ;
        RECT 547.950 145.950 550.050 146.400 ;
        RECT 586.950 145.950 589.050 146.400 ;
        RECT 592.950 145.950 595.050 146.400 ;
        RECT 148.950 144.600 151.050 145.050 ;
        RECT 160.950 144.600 163.050 145.050 ;
        RECT 148.950 143.400 163.050 144.600 ;
        RECT 148.950 142.950 151.050 143.400 ;
        RECT 160.950 142.950 163.050 143.400 ;
        RECT 175.950 144.600 178.050 145.050 ;
        RECT 187.950 144.600 190.050 145.050 ;
        RECT 271.950 144.600 274.050 145.050 ;
        RECT 175.950 143.400 274.050 144.600 ;
        RECT 175.950 142.950 178.050 143.400 ;
        RECT 187.950 142.950 190.050 143.400 ;
        RECT 271.950 142.950 274.050 143.400 ;
        RECT 373.950 144.600 376.050 145.050 ;
        RECT 382.950 144.600 385.050 145.050 ;
        RECT 373.950 143.400 385.050 144.600 ;
        RECT 373.950 142.950 376.050 143.400 ;
        RECT 382.950 142.950 385.050 143.400 ;
        RECT 1.950 141.600 4.050 142.050 ;
        RECT 133.950 141.600 136.050 142.050 ;
        RECT 1.950 140.400 136.050 141.600 ;
        RECT 1.950 139.950 4.050 140.400 ;
        RECT 133.950 139.950 136.050 140.400 ;
        RECT 160.950 141.600 163.050 142.050 ;
        RECT 178.950 141.600 181.050 142.050 ;
        RECT 160.950 140.400 181.050 141.600 ;
        RECT 160.950 139.950 163.050 140.400 ;
        RECT 178.950 139.950 181.050 140.400 ;
        RECT 229.950 141.600 232.050 142.050 ;
        RECT 247.950 141.600 250.050 142.050 ;
        RECT 229.950 140.400 250.050 141.600 ;
        RECT 229.950 139.950 232.050 140.400 ;
        RECT 247.950 139.950 250.050 140.400 ;
        RECT 265.950 141.600 268.050 142.050 ;
        RECT 322.950 141.600 325.050 142.050 ;
        RECT 265.950 140.400 325.050 141.600 ;
        RECT 265.950 139.950 268.050 140.400 ;
        RECT 322.950 139.950 325.050 140.400 ;
        RECT 76.950 138.600 79.050 139.050 ;
        RECT 112.950 138.600 115.050 139.050 ;
        RECT 121.950 138.600 124.050 139.050 ;
        RECT 76.950 137.400 124.050 138.600 ;
        RECT 76.950 136.950 79.050 137.400 ;
        RECT 112.950 136.950 115.050 137.400 ;
        RECT 121.950 136.950 124.050 137.400 ;
        RECT 151.950 138.600 154.050 139.050 ;
        RECT 166.950 138.600 169.050 139.050 ;
        RECT 151.950 137.400 169.050 138.600 ;
        RECT 151.950 136.950 154.050 137.400 ;
        RECT 166.950 136.950 169.050 137.400 ;
        RECT 178.950 138.600 181.050 139.050 ;
        RECT 196.950 138.600 199.050 139.050 ;
        RECT 178.950 137.400 199.050 138.600 ;
        RECT 178.950 136.950 181.050 137.400 ;
        RECT 196.950 136.950 199.050 137.400 ;
        RECT 202.950 138.600 205.050 139.050 ;
        RECT 214.950 138.600 217.050 139.050 ;
        RECT 202.950 137.400 217.050 138.600 ;
        RECT 202.950 136.950 205.050 137.400 ;
        RECT 214.950 136.950 217.050 137.400 ;
        RECT 241.950 138.600 244.050 139.050 ;
        RECT 274.950 138.600 277.050 139.050 ;
        RECT 241.950 137.400 277.050 138.600 ;
        RECT 241.950 136.950 244.050 137.400 ;
        RECT 274.950 136.950 277.050 137.400 ;
        RECT 673.950 138.600 676.050 139.050 ;
        RECT 691.950 138.600 694.050 139.050 ;
        RECT 673.950 137.400 694.050 138.600 ;
        RECT 673.950 136.950 676.050 137.400 ;
        RECT 691.950 136.950 694.050 137.400 ;
        RECT 697.950 138.600 700.050 139.050 ;
        RECT 712.950 138.600 715.050 139.050 ;
        RECT 697.950 137.400 715.050 138.600 ;
        RECT 697.950 136.950 700.050 137.400 ;
        RECT 712.950 136.950 715.050 137.400 ;
        RECT 73.950 135.600 76.050 136.050 ;
        RECT 85.950 135.600 88.050 136.050 ;
        RECT 73.950 134.400 88.050 135.600 ;
        RECT 73.950 133.950 76.050 134.400 ;
        RECT 85.950 133.950 88.050 134.400 ;
        RECT 127.950 135.600 130.050 136.050 ;
        RECT 136.950 135.600 139.050 136.050 ;
        RECT 181.950 135.600 184.050 136.050 ;
        RECT 127.950 134.400 184.050 135.600 ;
        RECT 127.950 133.950 130.050 134.400 ;
        RECT 136.950 133.950 139.050 134.400 ;
        RECT 181.950 133.950 184.050 134.400 ;
        RECT 247.950 135.600 250.050 136.050 ;
        RECT 289.950 135.600 292.050 136.050 ;
        RECT 247.950 134.400 292.050 135.600 ;
        RECT 247.950 133.950 250.050 134.400 ;
        RECT 289.950 133.950 292.050 134.400 ;
        RECT 682.950 135.600 685.050 136.050 ;
        RECT 712.950 135.600 715.050 136.050 ;
        RECT 682.950 134.400 715.050 135.600 ;
        RECT 682.950 133.950 685.050 134.400 ;
        RECT 712.950 133.950 715.050 134.400 ;
        RECT 10.950 132.600 13.050 133.050 ;
        RECT 43.950 132.600 46.050 133.050 ;
        RECT 160.950 132.600 163.050 133.050 ;
        RECT 10.950 131.400 46.050 132.600 ;
        RECT 10.950 130.950 13.050 131.400 ;
        RECT 43.950 130.950 46.050 131.400 ;
        RECT 158.400 131.400 163.050 132.600 ;
        RECT 158.400 130.050 159.600 131.400 ;
        RECT 160.950 130.950 163.050 131.400 ;
        RECT 181.950 132.600 184.050 133.050 ;
        RECT 190.950 132.600 193.050 133.050 ;
        RECT 181.950 131.400 193.050 132.600 ;
        RECT 181.950 130.950 184.050 131.400 ;
        RECT 190.950 130.950 193.050 131.400 ;
        RECT 205.950 132.600 208.050 133.050 ;
        RECT 232.950 132.600 235.050 133.050 ;
        RECT 205.950 131.400 235.050 132.600 ;
        RECT 205.950 130.950 208.050 131.400 ;
        RECT 230.400 130.050 231.600 131.400 ;
        RECT 232.950 130.950 235.050 131.400 ;
        RECT 238.950 132.600 241.050 133.050 ;
        RECT 259.950 132.600 262.050 133.050 ;
        RECT 274.950 132.600 277.050 133.050 ;
        RECT 238.950 131.400 277.050 132.600 ;
        RECT 238.950 130.950 241.050 131.400 ;
        RECT 259.950 130.950 262.050 131.400 ;
        RECT 274.950 130.950 277.050 131.400 ;
        RECT 289.950 132.600 292.050 133.050 ;
        RECT 298.950 132.600 301.050 133.050 ;
        RECT 361.950 132.600 364.050 133.050 ;
        RECT 289.950 131.400 364.050 132.600 ;
        RECT 289.950 130.950 292.050 131.400 ;
        RECT 298.950 130.950 301.050 131.400 ;
        RECT 361.950 130.950 364.050 131.400 ;
        RECT 691.950 132.600 694.050 133.050 ;
        RECT 709.950 132.600 712.050 133.050 ;
        RECT 691.950 131.400 712.050 132.600 ;
        RECT 691.950 130.950 694.050 131.400 ;
        RECT 709.950 130.950 712.050 131.400 ;
        RECT 37.950 129.600 40.050 130.050 ;
        RECT 55.950 129.600 58.050 130.050 ;
        RECT 67.950 129.600 70.050 130.050 ;
        RECT 35.400 128.400 40.050 129.600 ;
        RECT 35.400 124.050 36.600 128.400 ;
        RECT 37.950 127.950 40.050 128.400 ;
        RECT 41.400 128.400 54.600 129.600 ;
        RECT 37.950 126.600 40.050 127.050 ;
        RECT 41.400 126.600 42.600 128.400 ;
        RECT 37.950 125.400 42.600 126.600 ;
        RECT 37.950 124.950 40.050 125.400 ;
        RECT 49.950 124.950 52.050 127.050 ;
        RECT 16.950 123.600 19.050 124.050 ;
        RECT 19.950 123.600 22.050 124.050 ;
        RECT 28.950 123.600 31.050 124.050 ;
        RECT 16.950 122.400 31.050 123.600 ;
        RECT 16.950 121.950 19.050 122.400 ;
        RECT 19.950 121.950 22.050 122.400 ;
        RECT 28.950 121.950 31.050 122.400 ;
        RECT 34.950 121.950 37.050 124.050 ;
        RECT 1.950 120.600 4.050 121.050 ;
        RECT 22.950 120.600 25.050 121.050 ;
        RECT 50.400 120.600 51.600 124.950 ;
        RECT 53.400 124.050 54.600 128.400 ;
        RECT 55.950 128.400 70.050 129.600 ;
        RECT 55.950 127.950 58.050 128.400 ;
        RECT 67.950 127.950 70.050 128.400 ;
        RECT 85.950 129.600 88.050 130.050 ;
        RECT 97.950 129.600 100.050 130.050 ;
        RECT 85.950 128.400 100.050 129.600 ;
        RECT 85.950 127.950 88.050 128.400 ;
        RECT 97.950 127.950 100.050 128.400 ;
        RECT 103.950 129.600 106.050 130.050 ;
        RECT 109.950 129.600 112.050 130.050 ;
        RECT 103.950 128.400 112.050 129.600 ;
        RECT 103.950 127.950 106.050 128.400 ;
        RECT 109.950 127.950 112.050 128.400 ;
        RECT 124.950 129.600 127.050 130.050 ;
        RECT 133.950 129.600 136.050 130.050 ;
        RECT 142.950 129.600 145.050 130.050 ;
        RECT 145.950 129.600 148.050 130.050 ;
        RECT 151.950 129.600 154.050 130.050 ;
        RECT 124.950 128.400 129.600 129.600 ;
        RECT 124.950 127.950 127.050 128.400 ;
        RECT 73.950 126.600 76.050 127.050 ;
        RECT 59.400 125.400 76.050 126.600 ;
        RECT 59.400 124.050 60.600 125.400 ;
        RECT 73.950 124.950 76.050 125.400 ;
        RECT 103.950 126.600 106.050 127.050 ;
        RECT 103.950 125.400 126.600 126.600 ;
        RECT 103.950 124.950 106.050 125.400 ;
        RECT 125.400 124.050 126.600 125.400 ;
        RECT 128.400 124.050 129.600 128.400 ;
        RECT 133.950 128.400 141.600 129.600 ;
        RECT 133.950 127.950 136.050 128.400 ;
        RECT 140.400 126.600 141.600 128.400 ;
        RECT 142.950 128.400 154.050 129.600 ;
        RECT 142.950 127.950 145.050 128.400 ;
        RECT 145.950 127.950 148.050 128.400 ;
        RECT 151.950 127.950 154.050 128.400 ;
        RECT 157.950 127.950 160.050 130.050 ;
        RECT 163.950 127.950 166.050 130.050 ;
        RECT 166.950 129.600 169.050 130.050 ;
        RECT 199.950 129.600 202.050 130.050 ;
        RECT 205.950 129.600 208.050 130.050 ;
        RECT 166.950 128.400 208.050 129.600 ;
        RECT 166.950 127.950 169.050 128.400 ;
        RECT 199.950 127.950 202.050 128.400 ;
        RECT 205.950 127.950 208.050 128.400 ;
        RECT 229.950 127.950 232.050 130.050 ;
        RECT 295.950 129.600 298.050 130.050 ;
        RECT 352.950 129.600 355.050 130.050 ;
        RECT 373.950 129.600 376.050 130.050 ;
        RECT 382.950 129.600 385.050 130.050 ;
        RECT 412.950 129.600 415.050 130.050 ;
        RECT 295.950 128.400 366.600 129.600 ;
        RECT 295.950 127.950 298.050 128.400 ;
        RECT 352.950 127.950 355.050 128.400 ;
        RECT 157.950 126.600 160.050 127.050 ;
        RECT 140.400 125.400 160.050 126.600 ;
        RECT 157.950 124.950 160.050 125.400 ;
        RECT 164.400 124.050 165.600 127.950 ;
        RECT 365.400 127.050 366.600 128.400 ;
        RECT 373.950 128.400 381.600 129.600 ;
        RECT 373.950 127.950 376.050 128.400 ;
        RECT 178.950 126.600 181.050 127.050 ;
        RECT 187.950 126.600 190.050 127.050 ;
        RECT 178.950 125.400 190.050 126.600 ;
        RECT 178.950 124.950 181.050 125.400 ;
        RECT 187.950 124.950 190.050 125.400 ;
        RECT 193.950 124.950 196.050 127.050 ;
        RECT 211.950 126.600 214.050 127.050 ;
        RECT 232.950 126.600 235.050 127.050 ;
        RECT 250.950 126.600 253.050 127.050 ;
        RECT 307.950 126.600 310.050 127.050 ;
        RECT 211.950 125.400 253.050 126.600 ;
        RECT 211.950 124.950 214.050 125.400 ;
        RECT 232.950 124.950 235.050 125.400 ;
        RECT 250.950 124.950 253.050 125.400 ;
        RECT 263.400 125.400 310.050 126.600 ;
        RECT 52.950 121.950 55.050 124.050 ;
        RECT 58.950 121.950 61.050 124.050 ;
        RECT 112.950 123.600 115.050 124.050 ;
        RECT 104.400 122.400 115.050 123.600 ;
        RECT 64.950 120.600 67.050 121.050 ;
        RECT 73.950 120.600 76.050 121.050 ;
        RECT 1.950 119.400 76.050 120.600 ;
        RECT 1.950 118.950 4.050 119.400 ;
        RECT 22.950 118.950 25.050 119.400 ;
        RECT 64.950 118.950 67.050 119.400 ;
        RECT 73.950 118.950 76.050 119.400 ;
        RECT 100.950 120.600 103.050 121.050 ;
        RECT 104.400 120.600 105.600 122.400 ;
        RECT 112.950 121.950 115.050 122.400 ;
        RECT 124.950 121.950 127.050 124.050 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 133.950 123.600 136.050 124.050 ;
        RECT 145.950 123.600 148.050 124.050 ;
        RECT 133.950 122.400 148.050 123.600 ;
        RECT 133.950 121.950 136.050 122.400 ;
        RECT 145.950 121.950 148.050 122.400 ;
        RECT 163.950 121.950 166.050 124.050 ;
        RECT 194.400 123.600 195.600 124.950 ;
        RECT 263.400 124.050 264.600 125.400 ;
        RECT 307.950 124.950 310.050 125.400 ;
        RECT 319.950 126.600 322.050 127.050 ;
        RECT 328.950 126.600 331.050 127.050 ;
        RECT 319.950 125.400 331.050 126.600 ;
        RECT 319.950 124.950 322.050 125.400 ;
        RECT 328.950 124.950 331.050 125.400 ;
        RECT 346.950 126.600 349.050 127.050 ;
        RECT 358.950 126.600 361.050 127.050 ;
        RECT 346.950 125.400 361.050 126.600 ;
        RECT 346.950 124.950 349.050 125.400 ;
        RECT 358.950 124.950 361.050 125.400 ;
        RECT 364.950 124.950 367.050 127.050 ;
        RECT 380.400 126.600 381.600 128.400 ;
        RECT 382.950 128.400 415.050 129.600 ;
        RECT 382.950 127.950 385.050 128.400 ;
        RECT 412.950 127.950 415.050 128.400 ;
        RECT 418.950 129.600 421.050 130.050 ;
        RECT 433.950 129.600 436.050 130.050 ;
        RECT 439.950 129.600 442.050 130.050 ;
        RECT 418.950 128.400 442.050 129.600 ;
        RECT 418.950 127.950 421.050 128.400 ;
        RECT 433.950 127.950 436.050 128.400 ;
        RECT 439.950 127.950 442.050 128.400 ;
        RECT 496.950 127.950 499.050 130.050 ;
        RECT 502.950 129.600 505.050 130.050 ;
        RECT 508.950 129.600 511.050 130.050 ;
        RECT 502.950 128.400 511.050 129.600 ;
        RECT 502.950 127.950 505.050 128.400 ;
        RECT 508.950 127.950 511.050 128.400 ;
        RECT 544.950 129.600 547.050 130.050 ;
        RECT 556.950 129.600 559.050 130.050 ;
        RECT 544.950 128.400 559.050 129.600 ;
        RECT 544.950 127.950 547.050 128.400 ;
        RECT 556.950 127.950 559.050 128.400 ;
        RECT 589.950 129.600 592.050 130.050 ;
        RECT 601.950 129.600 604.050 130.050 ;
        RECT 589.950 128.400 604.050 129.600 ;
        RECT 589.950 127.950 592.050 128.400 ;
        RECT 601.950 127.950 604.050 128.400 ;
        RECT 604.950 127.950 607.050 130.050 ;
        RECT 700.950 127.950 703.050 130.050 ;
        RECT 385.950 126.600 388.050 127.050 ;
        RECT 380.400 125.400 388.050 126.600 ;
        RECT 385.950 124.950 388.050 125.400 ;
        RECT 388.950 126.600 391.050 127.050 ;
        RECT 394.950 126.600 397.050 127.050 ;
        RECT 388.950 125.400 397.050 126.600 ;
        RECT 388.950 124.950 391.050 125.400 ;
        RECT 394.950 124.950 397.050 125.400 ;
        RECT 400.950 124.950 403.050 127.050 ;
        RECT 415.950 126.600 418.050 127.050 ;
        RECT 427.950 126.600 430.050 127.050 ;
        RECT 415.950 125.400 430.050 126.600 ;
        RECT 415.950 124.950 418.050 125.400 ;
        RECT 427.950 124.950 430.050 125.400 ;
        RECT 442.950 124.950 445.050 127.050 ;
        RECT 460.950 126.600 463.050 127.050 ;
        RECT 484.950 126.600 487.050 127.050 ;
        RECT 460.950 125.400 487.050 126.600 ;
        RECT 460.950 124.950 463.050 125.400 ;
        RECT 484.950 124.950 487.050 125.400 ;
        RECT 232.950 123.600 235.050 124.050 ;
        RECT 194.400 122.400 235.050 123.600 ;
        RECT 232.950 121.950 235.050 122.400 ;
        RECT 238.950 123.600 241.050 124.050 ;
        RECT 256.950 123.600 259.050 124.050 ;
        RECT 238.950 122.400 259.050 123.600 ;
        RECT 238.950 121.950 241.050 122.400 ;
        RECT 256.950 121.950 259.050 122.400 ;
        RECT 262.950 121.950 265.050 124.050 ;
        RECT 265.950 123.600 268.050 124.050 ;
        RECT 271.950 123.600 274.050 124.050 ;
        RECT 325.950 123.600 328.050 124.050 ;
        RECT 265.950 122.400 274.050 123.600 ;
        RECT 265.950 121.950 268.050 122.400 ;
        RECT 271.950 121.950 274.050 122.400 ;
        RECT 284.400 122.400 328.050 123.600 ;
        RECT 100.950 119.400 105.600 120.600 ;
        RECT 106.950 120.600 109.050 121.050 ;
        RECT 139.950 120.600 142.050 121.050 ;
        RECT 106.950 119.400 142.050 120.600 ;
        RECT 100.950 118.950 103.050 119.400 ;
        RECT 106.950 118.950 109.050 119.400 ;
        RECT 139.950 118.950 142.050 119.400 ;
        RECT 163.950 120.600 166.050 121.050 ;
        RECT 202.950 120.600 205.050 121.050 ;
        RECT 163.950 119.400 205.050 120.600 ;
        RECT 163.950 118.950 166.050 119.400 ;
        RECT 202.950 118.950 205.050 119.400 ;
        RECT 256.950 120.600 259.050 121.050 ;
        RECT 268.950 120.600 271.050 121.050 ;
        RECT 284.400 120.600 285.600 122.400 ;
        RECT 325.950 121.950 328.050 122.400 ;
        RECT 331.950 123.600 334.050 124.050 ;
        RECT 340.950 123.600 343.050 124.050 ;
        RECT 331.950 122.400 343.050 123.600 ;
        RECT 331.950 121.950 334.050 122.400 ;
        RECT 340.950 121.950 343.050 122.400 ;
        RECT 391.950 123.600 394.050 124.050 ;
        RECT 401.400 123.600 402.600 124.950 ;
        RECT 391.950 122.400 402.600 123.600 ;
        RECT 403.950 123.600 406.050 124.050 ;
        RECT 424.950 123.600 427.050 124.050 ;
        RECT 403.950 122.400 427.050 123.600 ;
        RECT 391.950 121.950 394.050 122.400 ;
        RECT 403.950 121.950 406.050 122.400 ;
        RECT 424.950 121.950 427.050 122.400 ;
        RECT 436.950 123.600 439.050 124.050 ;
        RECT 443.400 123.600 444.600 124.950 ;
        RECT 457.950 123.600 460.050 124.050 ;
        RECT 487.950 123.600 490.050 124.050 ;
        RECT 497.400 123.600 498.600 127.950 ;
        RECT 499.950 126.600 502.050 127.050 ;
        RECT 505.950 126.600 508.050 127.050 ;
        RECT 499.950 125.400 508.050 126.600 ;
        RECT 499.950 124.950 502.050 125.400 ;
        RECT 505.950 124.950 508.050 125.400 ;
        RECT 595.950 126.600 598.050 127.050 ;
        RECT 605.400 126.600 606.600 127.950 ;
        RECT 595.950 125.400 606.600 126.600 ;
        RECT 595.950 124.950 598.050 125.400 ;
        RECT 436.950 122.400 456.600 123.600 ;
        RECT 436.950 121.950 439.050 122.400 ;
        RECT 256.950 119.400 271.050 120.600 ;
        RECT 256.950 118.950 259.050 119.400 ;
        RECT 268.950 118.950 271.050 119.400 ;
        RECT 275.400 119.400 285.600 120.600 ;
        RECT 286.950 120.600 289.050 121.050 ;
        RECT 292.950 120.600 295.050 121.050 ;
        RECT 286.950 119.400 295.050 120.600 ;
        RECT 25.950 117.600 28.050 118.050 ;
        RECT 43.950 117.600 46.050 118.050 ;
        RECT 25.950 116.400 46.050 117.600 ;
        RECT 25.950 115.950 28.050 116.400 ;
        RECT 43.950 115.950 46.050 116.400 ;
        RECT 103.950 117.600 106.050 118.050 ;
        RECT 130.950 117.600 133.050 118.050 ;
        RECT 103.950 116.400 133.050 117.600 ;
        RECT 103.950 115.950 106.050 116.400 ;
        RECT 130.950 115.950 133.050 116.400 ;
        RECT 160.950 117.600 163.050 118.050 ;
        RECT 193.950 117.600 196.050 118.050 ;
        RECT 223.950 117.600 226.050 118.050 ;
        RECT 160.950 116.400 226.050 117.600 ;
        RECT 160.950 115.950 163.050 116.400 ;
        RECT 193.950 115.950 196.050 116.400 ;
        RECT 223.950 115.950 226.050 116.400 ;
        RECT 256.950 117.600 259.050 118.050 ;
        RECT 275.400 117.600 276.600 119.400 ;
        RECT 286.950 118.950 289.050 119.400 ;
        RECT 292.950 118.950 295.050 119.400 ;
        RECT 301.950 120.600 304.050 121.050 ;
        RECT 325.950 120.600 328.050 121.050 ;
        RECT 301.950 119.400 328.050 120.600 ;
        RECT 301.950 118.950 304.050 119.400 ;
        RECT 325.950 118.950 328.050 119.400 ;
        RECT 334.950 120.600 337.050 121.050 ;
        RECT 343.950 120.600 346.050 121.050 ;
        RECT 334.950 119.400 346.050 120.600 ;
        RECT 334.950 118.950 337.050 119.400 ;
        RECT 343.950 118.950 346.050 119.400 ;
        RECT 385.950 120.600 388.050 121.050 ;
        RECT 397.950 120.600 400.050 121.050 ;
        RECT 385.950 119.400 400.050 120.600 ;
        RECT 385.950 118.950 388.050 119.400 ;
        RECT 397.950 118.950 400.050 119.400 ;
        RECT 445.950 120.600 448.050 121.050 ;
        RECT 451.950 120.600 454.050 121.050 ;
        RECT 445.950 119.400 454.050 120.600 ;
        RECT 455.400 120.600 456.600 122.400 ;
        RECT 457.950 122.400 474.600 123.600 ;
        RECT 457.950 121.950 460.050 122.400 ;
        RECT 473.400 121.050 474.600 122.400 ;
        RECT 487.950 122.400 498.600 123.600 ;
        RECT 487.950 121.950 490.050 122.400 ;
        RECT 511.950 121.950 514.050 124.050 ;
        RECT 520.950 123.600 523.050 124.050 ;
        RECT 529.950 123.600 532.050 124.050 ;
        RECT 520.950 122.400 532.050 123.600 ;
        RECT 520.950 121.950 523.050 122.400 ;
        RECT 529.950 121.950 532.050 122.400 ;
        RECT 538.950 123.600 541.050 124.050 ;
        RECT 544.950 123.600 547.050 124.050 ;
        RECT 538.950 122.400 547.050 123.600 ;
        RECT 538.950 121.950 541.050 122.400 ;
        RECT 544.950 121.950 547.050 122.400 ;
        RECT 568.950 123.600 571.050 124.050 ;
        RECT 598.950 123.600 601.050 124.050 ;
        RECT 568.950 122.400 601.050 123.600 ;
        RECT 568.950 121.950 571.050 122.400 ;
        RECT 598.950 121.950 601.050 122.400 ;
        RECT 610.950 123.600 613.050 124.050 ;
        RECT 637.950 123.600 640.050 124.050 ;
        RECT 646.950 123.600 649.050 124.050 ;
        RECT 610.950 122.400 649.050 123.600 ;
        RECT 610.950 121.950 613.050 122.400 ;
        RECT 637.950 121.950 640.050 122.400 ;
        RECT 646.950 121.950 649.050 122.400 ;
        RECT 667.950 123.600 670.050 124.050 ;
        RECT 694.950 123.600 697.050 124.050 ;
        RECT 667.950 122.400 697.050 123.600 ;
        RECT 667.950 121.950 670.050 122.400 ;
        RECT 694.950 121.950 697.050 122.400 ;
        RECT 463.950 120.600 466.050 121.050 ;
        RECT 455.400 119.400 466.050 120.600 ;
        RECT 445.950 118.950 448.050 119.400 ;
        RECT 451.950 118.950 454.050 119.400 ;
        RECT 463.950 118.950 466.050 119.400 ;
        RECT 472.950 120.600 475.050 121.050 ;
        RECT 512.400 120.600 513.600 121.950 ;
        RECT 701.400 121.050 702.600 127.950 ;
        RECT 472.950 119.400 513.600 120.600 ;
        RECT 523.950 120.600 526.050 121.050 ;
        RECT 556.950 120.600 559.050 121.050 ;
        RECT 523.950 119.400 559.050 120.600 ;
        RECT 472.950 118.950 475.050 119.400 ;
        RECT 523.950 118.950 526.050 119.400 ;
        RECT 556.950 118.950 559.050 119.400 ;
        RECT 577.950 120.600 580.050 121.050 ;
        RECT 616.950 120.600 619.050 121.050 ;
        RECT 622.950 120.600 625.050 121.050 ;
        RECT 625.950 120.600 628.050 121.050 ;
        RECT 661.950 120.600 664.050 121.050 ;
        RECT 694.950 120.600 697.050 121.050 ;
        RECT 577.950 119.400 697.050 120.600 ;
        RECT 577.950 118.950 580.050 119.400 ;
        RECT 616.950 118.950 619.050 119.400 ;
        RECT 622.950 118.950 625.050 119.400 ;
        RECT 625.950 118.950 628.050 119.400 ;
        RECT 661.950 118.950 664.050 119.400 ;
        RECT 694.950 118.950 697.050 119.400 ;
        RECT 700.950 118.950 703.050 121.050 ;
        RECT 256.950 116.400 276.600 117.600 ;
        RECT 277.950 117.600 280.050 118.050 ;
        RECT 289.950 117.600 292.050 118.050 ;
        RECT 298.950 117.600 301.050 118.050 ;
        RECT 277.950 116.400 301.050 117.600 ;
        RECT 256.950 115.950 259.050 116.400 ;
        RECT 277.950 115.950 280.050 116.400 ;
        RECT 289.950 115.950 292.050 116.400 ;
        RECT 298.950 115.950 301.050 116.400 ;
        RECT 307.950 117.600 310.050 118.050 ;
        RECT 337.950 117.600 340.050 118.050 ;
        RECT 307.950 116.400 340.050 117.600 ;
        RECT 307.950 115.950 310.050 116.400 ;
        RECT 337.950 115.950 340.050 116.400 ;
        RECT 460.950 117.600 463.050 118.050 ;
        RECT 466.950 117.600 469.050 118.050 ;
        RECT 460.950 116.400 469.050 117.600 ;
        RECT 460.950 115.950 463.050 116.400 ;
        RECT 466.950 115.950 469.050 116.400 ;
        RECT 469.950 117.600 472.050 118.050 ;
        RECT 478.950 117.600 481.050 118.050 ;
        RECT 469.950 116.400 481.050 117.600 ;
        RECT 469.950 115.950 472.050 116.400 ;
        RECT 478.950 115.950 481.050 116.400 ;
        RECT 589.950 117.600 592.050 118.050 ;
        RECT 610.950 117.600 613.050 118.050 ;
        RECT 589.950 116.400 613.050 117.600 ;
        RECT 589.950 115.950 592.050 116.400 ;
        RECT 610.950 115.950 613.050 116.400 ;
        RECT 655.950 117.600 658.050 118.050 ;
        RECT 703.950 117.600 706.050 118.050 ;
        RECT 655.950 116.400 706.050 117.600 ;
        RECT 655.950 115.950 658.050 116.400 ;
        RECT 703.950 115.950 706.050 116.400 ;
        RECT 88.950 114.600 91.050 115.050 ;
        RECT 97.950 114.600 100.050 115.050 ;
        RECT 109.950 114.600 112.050 115.050 ;
        RECT 88.950 113.400 112.050 114.600 ;
        RECT 88.950 112.950 91.050 113.400 ;
        RECT 97.950 112.950 100.050 113.400 ;
        RECT 109.950 112.950 112.050 113.400 ;
        RECT 154.950 114.600 157.050 115.050 ;
        RECT 169.950 114.600 172.050 115.050 ;
        RECT 154.950 113.400 172.050 114.600 ;
        RECT 154.950 112.950 157.050 113.400 ;
        RECT 169.950 112.950 172.050 113.400 ;
        RECT 190.950 114.600 193.050 115.050 ;
        RECT 208.950 114.600 211.050 115.050 ;
        RECT 190.950 113.400 211.050 114.600 ;
        RECT 190.950 112.950 193.050 113.400 ;
        RECT 208.950 112.950 211.050 113.400 ;
        RECT 211.950 114.600 214.050 115.050 ;
        RECT 241.950 114.600 244.050 115.050 ;
        RECT 211.950 113.400 244.050 114.600 ;
        RECT 211.950 112.950 214.050 113.400 ;
        RECT 241.950 112.950 244.050 113.400 ;
        RECT 259.950 114.600 262.050 115.050 ;
        RECT 274.950 114.600 277.050 115.050 ;
        RECT 259.950 113.400 277.050 114.600 ;
        RECT 259.950 112.950 262.050 113.400 ;
        RECT 274.950 112.950 277.050 113.400 ;
        RECT 298.950 114.600 301.050 115.050 ;
        RECT 328.950 114.600 331.050 115.050 ;
        RECT 364.950 114.600 367.050 115.050 ;
        RECT 298.950 113.400 367.050 114.600 ;
        RECT 298.950 112.950 301.050 113.400 ;
        RECT 328.950 112.950 331.050 113.400 ;
        RECT 364.950 112.950 367.050 113.400 ;
        RECT 448.950 114.600 451.050 115.050 ;
        RECT 460.950 114.600 463.050 115.050 ;
        RECT 448.950 113.400 463.050 114.600 ;
        RECT 448.950 112.950 451.050 113.400 ;
        RECT 460.950 112.950 463.050 113.400 ;
        RECT 499.950 114.600 502.050 115.050 ;
        RECT 508.950 114.600 511.050 115.050 ;
        RECT 499.950 113.400 511.050 114.600 ;
        RECT 499.950 112.950 502.050 113.400 ;
        RECT 508.950 112.950 511.050 113.400 ;
        RECT 628.950 114.600 631.050 115.050 ;
        RECT 667.950 114.600 670.050 115.050 ;
        RECT 628.950 113.400 670.050 114.600 ;
        RECT 628.950 112.950 631.050 113.400 ;
        RECT 667.950 112.950 670.050 113.400 ;
        RECT 184.950 111.600 187.050 112.050 ;
        RECT 214.950 111.600 217.050 112.050 ;
        RECT 184.950 110.400 217.050 111.600 ;
        RECT 184.950 109.950 187.050 110.400 ;
        RECT 214.950 109.950 217.050 110.400 ;
        RECT 220.950 111.600 223.050 112.050 ;
        RECT 262.950 111.600 265.050 112.050 ;
        RECT 220.950 110.400 265.050 111.600 ;
        RECT 220.950 109.950 223.050 110.400 ;
        RECT 262.950 109.950 265.050 110.400 ;
        RECT 295.950 111.600 298.050 112.050 ;
        RECT 319.950 111.600 322.050 112.050 ;
        RECT 295.950 110.400 322.050 111.600 ;
        RECT 295.950 109.950 298.050 110.400 ;
        RECT 319.950 109.950 322.050 110.400 ;
        RECT 340.950 111.600 343.050 112.050 ;
        RECT 385.950 111.600 388.050 112.050 ;
        RECT 340.950 110.400 388.050 111.600 ;
        RECT 340.950 109.950 343.050 110.400 ;
        RECT 385.950 109.950 388.050 110.400 ;
        RECT 79.950 108.600 82.050 109.050 ;
        RECT 148.950 108.600 151.050 109.050 ;
        RECT 79.950 107.400 151.050 108.600 ;
        RECT 79.950 106.950 82.050 107.400 ;
        RECT 148.950 106.950 151.050 107.400 ;
        RECT 184.950 108.600 187.050 109.050 ;
        RECT 253.950 108.600 256.050 109.050 ;
        RECT 292.950 108.600 295.050 109.050 ;
        RECT 304.950 108.600 307.050 109.050 ;
        RECT 379.950 108.600 382.050 109.050 ;
        RECT 184.950 107.400 252.600 108.600 ;
        RECT 184.950 106.950 187.050 107.400 ;
        RECT 31.950 105.600 34.050 106.050 ;
        RECT 37.950 105.600 40.050 106.050 ;
        RECT 58.950 105.600 61.050 106.050 ;
        RECT 31.950 104.400 61.050 105.600 ;
        RECT 31.950 103.950 34.050 104.400 ;
        RECT 37.950 103.950 40.050 104.400 ;
        RECT 58.950 103.950 61.050 104.400 ;
        RECT 121.950 105.600 124.050 106.050 ;
        RECT 133.950 105.600 136.050 106.050 ;
        RECT 121.950 104.400 136.050 105.600 ;
        RECT 121.950 103.950 124.050 104.400 ;
        RECT 133.950 103.950 136.050 104.400 ;
        RECT 142.950 105.600 145.050 106.050 ;
        RECT 178.950 105.600 181.050 106.050 ;
        RECT 142.950 104.400 181.050 105.600 ;
        RECT 142.950 103.950 145.050 104.400 ;
        RECT 178.950 103.950 181.050 104.400 ;
        RECT 196.950 105.600 199.050 106.050 ;
        RECT 199.950 105.600 202.050 106.050 ;
        RECT 223.950 105.600 226.050 106.050 ;
        RECT 247.950 105.600 250.050 106.050 ;
        RECT 196.950 104.400 250.050 105.600 ;
        RECT 251.400 105.600 252.600 107.400 ;
        RECT 253.950 107.400 382.050 108.600 ;
        RECT 253.950 106.950 256.050 107.400 ;
        RECT 292.950 106.950 295.050 107.400 ;
        RECT 304.950 106.950 307.050 107.400 ;
        RECT 379.950 106.950 382.050 107.400 ;
        RECT 436.950 108.600 439.050 109.050 ;
        RECT 442.950 108.600 445.050 109.050 ;
        RECT 523.950 108.600 526.050 109.050 ;
        RECT 436.950 107.400 526.050 108.600 ;
        RECT 436.950 106.950 439.050 107.400 ;
        RECT 442.950 106.950 445.050 107.400 ;
        RECT 523.950 106.950 526.050 107.400 ;
        RECT 565.950 108.600 568.050 109.050 ;
        RECT 631.950 108.600 634.050 109.050 ;
        RECT 565.950 107.400 634.050 108.600 ;
        RECT 565.950 106.950 568.050 107.400 ;
        RECT 631.950 106.950 634.050 107.400 ;
        RECT 307.950 105.600 310.050 106.050 ;
        RECT 251.400 104.400 310.050 105.600 ;
        RECT 196.950 103.950 199.050 104.400 ;
        RECT 199.950 103.950 202.050 104.400 ;
        RECT 223.950 103.950 226.050 104.400 ;
        RECT 247.950 103.950 250.050 104.400 ;
        RECT 307.950 103.950 310.050 104.400 ;
        RECT 313.950 105.600 316.050 106.050 ;
        RECT 355.950 105.600 358.050 106.050 ;
        RECT 367.950 105.600 370.050 106.050 ;
        RECT 313.950 104.400 370.050 105.600 ;
        RECT 313.950 103.950 316.050 104.400 ;
        RECT 355.950 103.950 358.050 104.400 ;
        RECT 367.950 103.950 370.050 104.400 ;
        RECT 22.950 102.600 25.050 103.050 ;
        RECT 46.950 102.600 49.050 103.050 ;
        RECT 52.950 102.600 55.050 103.050 ;
        RECT 22.950 101.400 55.050 102.600 ;
        RECT 22.950 100.950 25.050 101.400 ;
        RECT 46.950 100.950 49.050 101.400 ;
        RECT 52.950 100.950 55.050 101.400 ;
        RECT 64.950 102.600 67.050 103.050 ;
        RECT 100.950 102.600 103.050 103.050 ;
        RECT 64.950 101.400 103.050 102.600 ;
        RECT 64.950 100.950 67.050 101.400 ;
        RECT 100.950 100.950 103.050 101.400 ;
        RECT 118.950 102.600 121.050 103.050 ;
        RECT 136.950 102.600 139.050 103.050 ;
        RECT 118.950 101.400 139.050 102.600 ;
        RECT 118.950 100.950 121.050 101.400 ;
        RECT 136.950 100.950 139.050 101.400 ;
        RECT 151.950 102.600 154.050 103.050 ;
        RECT 166.950 102.600 169.050 103.050 ;
        RECT 151.950 101.400 169.050 102.600 ;
        RECT 151.950 100.950 154.050 101.400 ;
        RECT 166.950 100.950 169.050 101.400 ;
        RECT 214.950 102.600 217.050 103.050 ;
        RECT 229.950 102.600 232.050 103.050 ;
        RECT 214.950 101.400 232.050 102.600 ;
        RECT 214.950 100.950 217.050 101.400 ;
        RECT 229.950 100.950 232.050 101.400 ;
        RECT 238.950 102.600 241.050 103.050 ;
        RECT 259.950 102.600 262.050 103.050 ;
        RECT 238.950 101.400 262.050 102.600 ;
        RECT 238.950 100.950 241.050 101.400 ;
        RECT 259.950 100.950 262.050 101.400 ;
        RECT 349.950 102.600 352.050 103.050 ;
        RECT 355.950 102.600 358.050 103.050 ;
        RECT 370.950 102.600 373.050 103.050 ;
        RECT 349.950 101.400 373.050 102.600 ;
        RECT 349.950 100.950 352.050 101.400 ;
        RECT 355.950 100.950 358.050 101.400 ;
        RECT 370.950 100.950 373.050 101.400 ;
        RECT 502.950 102.600 505.050 103.050 ;
        RECT 526.950 102.600 529.050 103.050 ;
        RECT 502.950 101.400 529.050 102.600 ;
        RECT 502.950 100.950 505.050 101.400 ;
        RECT 526.950 100.950 529.050 101.400 ;
        RECT 550.950 102.600 553.050 103.050 ;
        RECT 574.950 102.600 577.050 103.050 ;
        RECT 589.950 102.600 592.050 103.050 ;
        RECT 604.950 102.600 607.050 103.050 ;
        RECT 658.950 102.600 661.050 103.050 ;
        RECT 673.950 102.600 676.050 103.050 ;
        RECT 550.950 101.400 676.050 102.600 ;
        RECT 550.950 100.950 553.050 101.400 ;
        RECT 574.950 100.950 577.050 101.400 ;
        RECT 589.950 100.950 592.050 101.400 ;
        RECT 604.950 100.950 607.050 101.400 ;
        RECT 658.950 100.950 661.050 101.400 ;
        RECT 673.950 100.950 676.050 101.400 ;
        RECT 7.950 99.600 10.050 100.050 ;
        RECT 19.950 99.600 22.050 100.050 ;
        RECT 28.950 99.600 31.050 100.050 ;
        RECT 40.950 99.600 43.050 100.050 ;
        RECT 55.950 99.600 58.050 100.050 ;
        RECT 7.950 98.400 15.600 99.600 ;
        RECT 7.950 97.950 10.050 98.400 ;
        RECT 14.400 93.600 15.600 98.400 ;
        RECT 19.950 98.400 24.600 99.600 ;
        RECT 19.950 97.950 22.050 98.400 ;
        RECT 23.400 94.050 24.600 98.400 ;
        RECT 28.950 98.400 43.050 99.600 ;
        RECT 28.950 97.950 31.050 98.400 ;
        RECT 40.950 97.950 43.050 98.400 ;
        RECT 47.400 98.400 58.050 99.600 ;
        RECT 29.400 94.050 30.600 97.950 ;
        RECT 34.950 96.600 37.050 97.050 ;
        RECT 40.950 96.600 43.050 97.050 ;
        RECT 34.950 95.400 43.050 96.600 ;
        RECT 34.950 94.950 37.050 95.400 ;
        RECT 40.950 94.950 43.050 95.400 ;
        RECT 47.400 94.050 48.600 98.400 ;
        RECT 55.950 97.950 58.050 98.400 ;
        RECT 67.950 99.600 70.050 100.050 ;
        RECT 130.950 99.600 133.050 100.050 ;
        RECT 148.950 99.600 151.050 100.050 ;
        RECT 154.950 99.600 157.050 100.050 ;
        RECT 67.950 98.400 78.600 99.600 ;
        RECT 67.950 97.950 70.050 98.400 ;
        RECT 52.950 96.600 55.050 97.050 ;
        RECT 73.950 96.600 76.050 97.050 ;
        RECT 52.950 95.400 76.050 96.600 ;
        RECT 77.400 96.600 78.600 98.400 ;
        RECT 130.950 98.400 157.050 99.600 ;
        RECT 130.950 97.950 133.050 98.400 ;
        RECT 148.950 97.950 151.050 98.400 ;
        RECT 154.950 97.950 157.050 98.400 ;
        RECT 157.950 99.600 160.050 100.050 ;
        RECT 238.950 99.600 241.050 100.050 ;
        RECT 157.950 98.400 162.600 99.600 ;
        RECT 157.950 97.950 160.050 98.400 ;
        RECT 85.950 96.600 88.050 97.050 ;
        RECT 106.950 96.600 109.050 97.050 ;
        RECT 77.400 95.400 88.050 96.600 ;
        RECT 52.950 94.950 55.050 95.400 ;
        RECT 73.950 94.950 76.050 95.400 ;
        RECT 85.950 94.950 88.050 95.400 ;
        RECT 98.400 95.400 109.050 96.600 ;
        RECT 19.950 93.600 22.050 94.050 ;
        RECT 14.400 92.400 22.050 93.600 ;
        RECT 19.950 91.950 22.050 92.400 ;
        RECT 22.950 91.950 25.050 94.050 ;
        RECT 28.950 91.950 31.050 94.050 ;
        RECT 46.950 91.950 49.050 94.050 ;
        RECT 49.950 93.600 52.050 94.050 ;
        RECT 58.950 93.600 61.050 94.050 ;
        RECT 49.950 92.400 61.050 93.600 ;
        RECT 49.950 91.950 52.050 92.400 ;
        RECT 58.950 91.950 61.050 92.400 ;
        RECT 70.950 93.600 73.050 94.050 ;
        RECT 94.950 93.600 97.050 94.050 ;
        RECT 98.400 93.600 99.600 95.400 ;
        RECT 106.950 94.950 109.050 95.400 ;
        RECT 121.950 96.600 124.050 97.050 ;
        RECT 127.950 96.600 130.050 97.050 ;
        RECT 151.950 96.600 154.050 97.050 ;
        RECT 157.950 96.600 160.050 97.050 ;
        RECT 121.950 95.400 132.600 96.600 ;
        RECT 121.950 94.950 124.050 95.400 ;
        RECT 127.950 94.950 130.050 95.400 ;
        RECT 70.950 92.400 75.600 93.600 ;
        RECT 70.950 91.950 73.050 92.400 ;
        RECT 74.400 91.050 75.600 92.400 ;
        RECT 94.950 92.400 99.600 93.600 ;
        RECT 94.950 91.950 97.050 92.400 ;
        RECT 131.400 91.050 132.600 95.400 ;
        RECT 151.950 95.400 160.050 96.600 ;
        RECT 151.950 94.950 154.050 95.400 ;
        RECT 157.950 94.950 160.050 95.400 ;
        RECT 161.400 94.050 162.600 98.400 ;
        RECT 236.400 98.400 241.050 99.600 ;
        RECT 163.950 96.600 166.050 97.050 ;
        RECT 169.950 96.600 172.050 97.050 ;
        RECT 163.950 95.400 172.050 96.600 ;
        RECT 163.950 94.950 166.050 95.400 ;
        RECT 169.950 94.950 172.050 95.400 ;
        RECT 205.950 96.600 208.050 97.050 ;
        RECT 211.950 96.600 214.050 97.050 ;
        RECT 236.400 96.600 237.600 98.400 ;
        RECT 238.950 97.950 241.050 98.400 ;
        RECT 247.950 99.600 250.050 100.050 ;
        RECT 256.950 99.600 259.050 100.050 ;
        RECT 247.950 98.400 259.050 99.600 ;
        RECT 247.950 97.950 250.050 98.400 ;
        RECT 256.950 97.950 259.050 98.400 ;
        RECT 265.950 99.600 268.050 100.050 ;
        RECT 271.950 99.600 274.050 100.050 ;
        RECT 265.950 98.400 274.050 99.600 ;
        RECT 265.950 97.950 268.050 98.400 ;
        RECT 271.950 97.950 274.050 98.400 ;
        RECT 301.950 97.950 304.050 100.050 ;
        RECT 316.950 99.600 319.050 100.050 ;
        RECT 314.400 98.400 319.050 99.600 ;
        RECT 302.400 96.600 303.600 97.950 ;
        RECT 314.400 96.600 315.600 98.400 ;
        RECT 316.950 97.950 319.050 98.400 ;
        RECT 346.950 99.600 349.050 100.050 ;
        RECT 349.950 99.600 352.050 100.050 ;
        RECT 361.950 99.600 364.050 100.050 ;
        RECT 346.950 98.400 364.050 99.600 ;
        RECT 346.950 97.950 349.050 98.400 ;
        RECT 349.950 97.950 352.050 98.400 ;
        RECT 361.950 97.950 364.050 98.400 ;
        RECT 367.950 99.600 370.050 100.050 ;
        RECT 376.950 99.600 379.050 100.050 ;
        RECT 367.950 98.400 379.050 99.600 ;
        RECT 367.950 97.950 370.050 98.400 ;
        RECT 376.950 97.950 379.050 98.400 ;
        RECT 400.950 97.950 403.050 100.050 ;
        RECT 454.950 99.600 457.050 100.050 ;
        RECT 478.950 99.600 481.050 100.050 ;
        RECT 481.950 99.600 484.050 100.050 ;
        RECT 454.950 98.400 484.050 99.600 ;
        RECT 454.950 97.950 457.050 98.400 ;
        RECT 478.950 97.950 481.050 98.400 ;
        RECT 481.950 97.950 484.050 98.400 ;
        RECT 484.950 99.600 487.050 100.050 ;
        RECT 490.950 99.600 493.050 100.050 ;
        RECT 508.950 99.600 511.050 100.050 ;
        RECT 484.950 98.400 511.050 99.600 ;
        RECT 484.950 97.950 487.050 98.400 ;
        RECT 490.950 97.950 493.050 98.400 ;
        RECT 508.950 97.950 511.050 98.400 ;
        RECT 517.950 99.600 520.050 100.050 ;
        RECT 523.950 99.600 526.050 100.050 ;
        RECT 535.950 99.600 538.050 100.050 ;
        RECT 517.950 98.400 538.050 99.600 ;
        RECT 517.950 97.950 520.050 98.400 ;
        RECT 523.950 97.950 526.050 98.400 ;
        RECT 535.950 97.950 538.050 98.400 ;
        RECT 571.950 99.600 574.050 100.050 ;
        RECT 601.950 99.600 604.050 100.050 ;
        RECT 571.950 98.400 604.050 99.600 ;
        RECT 571.950 97.950 574.050 98.400 ;
        RECT 601.950 97.950 604.050 98.400 ;
        RECT 205.950 95.400 214.050 96.600 ;
        RECT 205.950 94.950 208.050 95.400 ;
        RECT 211.950 94.950 214.050 95.400 ;
        RECT 221.400 95.400 237.600 96.600 ;
        RECT 260.400 95.400 303.600 96.600 ;
        RECT 311.400 95.400 315.600 96.600 ;
        RECT 316.950 96.600 319.050 97.050 ;
        RECT 331.950 96.600 334.050 97.050 ;
        RECT 316.950 95.400 334.050 96.600 ;
        RECT 133.950 93.600 136.050 94.050 ;
        RECT 139.950 93.600 142.050 94.050 ;
        RECT 133.950 92.400 142.050 93.600 ;
        RECT 133.950 91.950 136.050 92.400 ;
        RECT 139.950 91.950 142.050 92.400 ;
        RECT 145.950 93.600 148.050 94.050 ;
        RECT 151.950 93.600 154.050 94.050 ;
        RECT 145.950 92.400 154.050 93.600 ;
        RECT 145.950 91.950 148.050 92.400 ;
        RECT 151.950 91.950 154.050 92.400 ;
        RECT 160.950 91.950 163.050 94.050 ;
        RECT 166.950 93.600 169.050 94.050 ;
        RECT 175.950 93.600 178.050 94.050 ;
        RECT 166.950 92.400 178.050 93.600 ;
        RECT 166.950 91.950 169.050 92.400 ;
        RECT 175.950 91.950 178.050 92.400 ;
        RECT 181.950 93.600 184.050 94.050 ;
        RECT 187.950 93.600 190.050 94.050 ;
        RECT 181.950 92.400 190.050 93.600 ;
        RECT 181.950 91.950 184.050 92.400 ;
        RECT 187.950 91.950 190.050 92.400 ;
        RECT 193.950 93.600 196.050 94.050 ;
        RECT 221.400 93.600 222.600 95.400 ;
        RECT 193.950 92.400 222.600 93.600 ;
        RECT 238.950 93.600 241.050 94.050 ;
        RECT 260.400 93.600 261.600 95.400 ;
        RECT 238.950 92.400 261.600 93.600 ;
        RECT 262.950 93.600 265.050 94.050 ;
        RECT 298.950 93.600 301.050 94.050 ;
        RECT 311.400 93.600 312.600 95.400 ;
        RECT 316.950 94.950 319.050 95.400 ;
        RECT 331.950 94.950 334.050 95.400 ;
        RECT 337.950 96.600 340.050 97.050 ;
        RECT 358.950 96.600 361.050 97.050 ;
        RECT 370.950 96.600 373.050 97.050 ;
        RECT 337.950 95.400 345.600 96.600 ;
        RECT 337.950 94.950 340.050 95.400 ;
        RECT 344.400 94.050 345.600 95.400 ;
        RECT 358.950 95.400 373.050 96.600 ;
        RECT 358.950 94.950 361.050 95.400 ;
        RECT 370.950 94.950 373.050 95.400 ;
        RECT 401.400 94.050 402.600 97.950 ;
        RECT 403.950 96.600 406.050 97.050 ;
        RECT 415.950 96.600 418.050 97.050 ;
        RECT 439.950 96.600 442.050 97.050 ;
        RECT 403.950 95.400 442.050 96.600 ;
        RECT 403.950 94.950 406.050 95.400 ;
        RECT 415.950 94.950 418.050 95.400 ;
        RECT 439.950 94.950 442.050 95.400 ;
        RECT 475.950 96.600 478.050 97.050 ;
        RECT 487.950 96.600 490.050 97.050 ;
        RECT 475.950 95.400 490.050 96.600 ;
        RECT 475.950 94.950 478.050 95.400 ;
        RECT 487.950 94.950 490.050 95.400 ;
        RECT 493.950 96.600 496.050 97.050 ;
        RECT 511.950 96.600 514.050 97.050 ;
        RECT 493.950 95.400 514.050 96.600 ;
        RECT 493.950 94.950 496.050 95.400 ;
        RECT 511.950 94.950 514.050 95.400 ;
        RECT 529.950 96.600 532.050 97.050 ;
        RECT 550.950 96.600 553.050 97.050 ;
        RECT 529.950 95.400 553.050 96.600 ;
        RECT 529.950 94.950 532.050 95.400 ;
        RECT 550.950 94.950 553.050 95.400 ;
        RECT 580.950 96.600 583.050 97.050 ;
        RECT 586.950 96.600 589.050 97.050 ;
        RECT 580.950 95.400 589.050 96.600 ;
        RECT 580.950 94.950 583.050 95.400 ;
        RECT 586.950 94.950 589.050 95.400 ;
        RECT 592.950 96.600 595.050 97.050 ;
        RECT 604.950 96.600 607.050 97.050 ;
        RECT 592.950 95.400 607.050 96.600 ;
        RECT 592.950 94.950 595.050 95.400 ;
        RECT 604.950 94.950 607.050 95.400 ;
        RECT 613.950 96.600 616.050 97.050 ;
        RECT 622.950 96.600 625.050 97.050 ;
        RECT 613.950 95.400 625.050 96.600 ;
        RECT 613.950 94.950 616.050 95.400 ;
        RECT 622.950 94.950 625.050 95.400 ;
        RECT 697.950 96.600 700.050 97.050 ;
        RECT 700.950 96.600 703.050 97.050 ;
        RECT 706.950 96.600 709.050 97.050 ;
        RECT 697.950 95.400 709.050 96.600 ;
        RECT 697.950 94.950 700.050 95.400 ;
        RECT 700.950 94.950 703.050 95.400 ;
        RECT 706.950 94.950 709.050 95.400 ;
        RECT 262.950 92.400 276.600 93.600 ;
        RECT 193.950 91.950 196.050 92.400 ;
        RECT 238.950 91.950 241.050 92.400 ;
        RECT 262.950 91.950 265.050 92.400 ;
        RECT 275.400 91.050 276.600 92.400 ;
        RECT 298.950 92.400 312.600 93.600 ;
        RECT 313.950 93.600 316.050 94.050 ;
        RECT 313.950 92.400 321.600 93.600 ;
        RECT 298.950 91.950 301.050 92.400 ;
        RECT 313.950 91.950 316.050 92.400 ;
        RECT 25.950 90.600 28.050 91.050 ;
        RECT 31.950 90.600 34.050 91.050 ;
        RECT 43.950 90.600 46.050 91.050 ;
        RECT 55.950 90.600 58.050 91.050 ;
        RECT 25.950 89.400 58.050 90.600 ;
        RECT 25.950 88.950 28.050 89.400 ;
        RECT 31.950 88.950 34.050 89.400 ;
        RECT 43.950 88.950 46.050 89.400 ;
        RECT 55.950 88.950 58.050 89.400 ;
        RECT 73.950 88.950 76.050 91.050 ;
        RECT 115.950 90.600 118.050 91.050 ;
        RECT 127.950 90.600 130.050 91.050 ;
        RECT 115.950 89.400 130.050 90.600 ;
        RECT 115.950 88.950 118.050 89.400 ;
        RECT 127.950 88.950 130.050 89.400 ;
        RECT 130.950 88.950 133.050 91.050 ;
        RECT 160.950 90.600 163.050 91.050 ;
        RECT 205.950 90.600 208.050 91.050 ;
        RECT 160.950 89.400 208.050 90.600 ;
        RECT 160.950 88.950 163.050 89.400 ;
        RECT 205.950 88.950 208.050 89.400 ;
        RECT 217.950 90.600 220.050 91.050 ;
        RECT 235.950 90.600 238.050 91.050 ;
        RECT 217.950 89.400 238.050 90.600 ;
        RECT 217.950 88.950 220.050 89.400 ;
        RECT 235.950 88.950 238.050 89.400 ;
        RECT 256.950 90.600 259.050 91.050 ;
        RECT 262.950 90.600 265.050 91.050 ;
        RECT 256.950 89.400 265.050 90.600 ;
        RECT 256.950 88.950 259.050 89.400 ;
        RECT 262.950 88.950 265.050 89.400 ;
        RECT 274.950 88.950 277.050 91.050 ;
        RECT 295.950 90.600 298.050 91.050 ;
        RECT 316.950 90.600 319.050 91.050 ;
        RECT 295.950 89.400 319.050 90.600 ;
        RECT 320.400 90.600 321.600 92.400 ;
        RECT 325.950 91.950 328.050 94.050 ;
        RECT 343.950 93.600 346.050 94.050 ;
        RECT 352.950 93.600 355.050 94.050 ;
        RECT 367.950 93.600 370.050 94.050 ;
        RECT 343.950 92.400 355.050 93.600 ;
        RECT 343.950 91.950 346.050 92.400 ;
        RECT 352.950 91.950 355.050 92.400 ;
        RECT 356.400 92.400 370.050 93.600 ;
        RECT 322.950 90.600 325.050 91.050 ;
        RECT 320.400 89.400 325.050 90.600 ;
        RECT 295.950 88.950 298.050 89.400 ;
        RECT 316.950 88.950 319.050 89.400 ;
        RECT 322.950 88.950 325.050 89.400 ;
        RECT 79.950 87.600 82.050 88.050 ;
        RECT 133.950 87.600 136.050 88.050 ;
        RECT 79.950 86.400 136.050 87.600 ;
        RECT 79.950 85.950 82.050 86.400 ;
        RECT 133.950 85.950 136.050 86.400 ;
        RECT 211.950 87.600 214.050 88.050 ;
        RECT 250.950 87.600 253.050 88.050 ;
        RECT 263.400 87.600 264.600 88.950 ;
        RECT 326.400 88.050 327.600 91.950 ;
        RECT 328.950 90.600 331.050 91.050 ;
        RECT 340.950 90.600 343.050 91.050 ;
        RECT 328.950 89.400 343.050 90.600 ;
        RECT 328.950 88.950 331.050 89.400 ;
        RECT 340.950 88.950 343.050 89.400 ;
        RECT 343.950 90.600 346.050 91.050 ;
        RECT 356.400 90.600 357.600 92.400 ;
        RECT 367.950 91.950 370.050 92.400 ;
        RECT 370.950 93.600 373.050 94.050 ;
        RECT 376.950 93.600 379.050 94.050 ;
        RECT 370.950 92.400 379.050 93.600 ;
        RECT 370.950 91.950 373.050 92.400 ;
        RECT 376.950 91.950 379.050 92.400 ;
        RECT 400.950 91.950 403.050 94.050 ;
        RECT 409.950 93.600 412.050 94.050 ;
        RECT 404.400 92.400 412.050 93.600 ;
        RECT 343.950 89.400 357.600 90.600 ;
        RECT 343.950 88.950 346.050 89.400 ;
        RECT 367.950 88.950 370.050 91.050 ;
        RECT 373.950 90.600 376.050 91.050 ;
        RECT 382.950 90.600 385.050 91.050 ;
        RECT 373.950 89.400 385.050 90.600 ;
        RECT 373.950 88.950 376.050 89.400 ;
        RECT 382.950 88.950 385.050 89.400 ;
        RECT 397.950 90.600 400.050 91.050 ;
        RECT 404.400 90.600 405.600 92.400 ;
        RECT 409.950 91.950 412.050 92.400 ;
        RECT 463.950 93.600 466.050 94.050 ;
        RECT 472.950 93.600 475.050 94.050 ;
        RECT 490.950 93.600 493.050 94.050 ;
        RECT 463.950 92.400 493.050 93.600 ;
        RECT 463.950 91.950 466.050 92.400 ;
        RECT 472.950 91.950 475.050 92.400 ;
        RECT 490.950 91.950 493.050 92.400 ;
        RECT 493.950 93.600 496.050 94.050 ;
        RECT 505.950 93.600 508.050 94.050 ;
        RECT 493.950 92.400 508.050 93.600 ;
        RECT 493.950 91.950 496.050 92.400 ;
        RECT 505.950 91.950 508.050 92.400 ;
        RECT 517.950 93.600 520.050 94.050 ;
        RECT 526.950 93.600 529.050 94.050 ;
        RECT 517.950 92.400 529.050 93.600 ;
        RECT 517.950 91.950 520.050 92.400 ;
        RECT 526.950 91.950 529.050 92.400 ;
        RECT 532.950 93.600 535.050 94.050 ;
        RECT 571.950 93.600 574.050 94.050 ;
        RECT 532.950 92.400 574.050 93.600 ;
        RECT 532.950 91.950 535.050 92.400 ;
        RECT 571.950 91.950 574.050 92.400 ;
        RECT 583.950 93.600 586.050 94.050 ;
        RECT 595.950 93.600 598.050 94.050 ;
        RECT 583.950 92.400 598.050 93.600 ;
        RECT 583.950 91.950 586.050 92.400 ;
        RECT 595.950 91.950 598.050 92.400 ;
        RECT 634.950 93.600 637.050 94.050 ;
        RECT 640.950 93.600 643.050 94.050 ;
        RECT 634.950 92.400 643.050 93.600 ;
        RECT 634.950 91.950 637.050 92.400 ;
        RECT 640.950 91.950 643.050 92.400 ;
        RECT 652.950 93.600 655.050 94.050 ;
        RECT 664.950 93.600 667.050 94.050 ;
        RECT 652.950 92.400 667.050 93.600 ;
        RECT 652.950 91.950 655.050 92.400 ;
        RECT 664.950 91.950 667.050 92.400 ;
        RECT 397.950 89.400 405.600 90.600 ;
        RECT 397.950 88.950 400.050 89.400 ;
        RECT 406.950 88.950 409.050 91.050 ;
        RECT 457.950 90.600 460.050 91.050 ;
        RECT 484.950 90.600 487.050 91.050 ;
        RECT 457.950 89.400 487.050 90.600 ;
        RECT 457.950 88.950 460.050 89.400 ;
        RECT 484.950 88.950 487.050 89.400 ;
        RECT 598.950 90.600 601.050 91.050 ;
        RECT 604.950 90.600 607.050 91.050 ;
        RECT 598.950 89.400 607.050 90.600 ;
        RECT 598.950 88.950 601.050 89.400 ;
        RECT 604.950 88.950 607.050 89.400 ;
        RECT 631.950 90.600 634.050 91.050 ;
        RECT 637.950 90.600 640.050 91.050 ;
        RECT 631.950 89.400 640.050 90.600 ;
        RECT 631.950 88.950 634.050 89.400 ;
        RECT 637.950 88.950 640.050 89.400 ;
        RECT 211.950 86.400 264.600 87.600 ;
        RECT 265.950 87.600 268.050 88.050 ;
        RECT 277.950 87.600 280.050 88.050 ;
        RECT 265.950 86.400 280.050 87.600 ;
        RECT 211.950 85.950 214.050 86.400 ;
        RECT 250.950 85.950 253.050 86.400 ;
        RECT 265.950 85.950 268.050 86.400 ;
        RECT 277.950 85.950 280.050 86.400 ;
        RECT 283.950 87.600 286.050 88.050 ;
        RECT 325.950 87.600 328.050 88.050 ;
        RECT 368.400 87.600 369.600 88.950 ;
        RECT 283.950 86.400 324.600 87.600 ;
        RECT 283.950 85.950 286.050 86.400 ;
        RECT 323.400 84.600 324.600 86.400 ;
        RECT 325.950 86.400 369.600 87.600 ;
        RECT 325.950 85.950 328.050 86.400 ;
        RECT 407.400 84.600 408.600 88.950 ;
        RECT 475.950 87.600 478.050 88.050 ;
        RECT 481.950 87.600 484.050 88.050 ;
        RECT 475.950 86.400 484.050 87.600 ;
        RECT 475.950 85.950 478.050 86.400 ;
        RECT 481.950 85.950 484.050 86.400 ;
        RECT 586.950 87.600 589.050 88.050 ;
        RECT 613.950 87.600 616.050 88.050 ;
        RECT 586.950 86.400 616.050 87.600 ;
        RECT 586.950 85.950 589.050 86.400 ;
        RECT 613.950 85.950 616.050 86.400 ;
        RECT 323.400 83.400 408.600 84.600 ;
        RECT 103.950 81.600 106.050 82.050 ;
        RECT 115.950 81.600 118.050 82.050 ;
        RECT 103.950 80.400 118.050 81.600 ;
        RECT 103.950 79.950 106.050 80.400 ;
        RECT 115.950 79.950 118.050 80.400 ;
        RECT 166.950 81.600 169.050 82.050 ;
        RECT 172.950 81.600 175.050 82.050 ;
        RECT 223.950 81.600 226.050 82.050 ;
        RECT 271.950 81.600 274.050 82.050 ;
        RECT 301.950 81.600 304.050 82.050 ;
        RECT 166.950 80.400 226.050 81.600 ;
        RECT 166.950 79.950 169.050 80.400 ;
        RECT 172.950 79.950 175.050 80.400 ;
        RECT 223.950 79.950 226.050 80.400 ;
        RECT 251.400 80.400 304.050 81.600 ;
        RECT 46.950 78.600 49.050 79.050 ;
        RECT 70.950 78.600 73.050 79.050 ;
        RECT 46.950 77.400 73.050 78.600 ;
        RECT 46.950 76.950 49.050 77.400 ;
        RECT 70.950 76.950 73.050 77.400 ;
        RECT 202.950 78.600 205.050 79.050 ;
        RECT 229.950 78.600 232.050 79.050 ;
        RECT 202.950 77.400 232.050 78.600 ;
        RECT 202.950 76.950 205.050 77.400 ;
        RECT 229.950 76.950 232.050 77.400 ;
        RECT 232.950 78.600 235.050 79.050 ;
        RECT 238.950 78.600 241.050 79.050 ;
        RECT 232.950 77.400 241.050 78.600 ;
        RECT 232.950 76.950 235.050 77.400 ;
        RECT 238.950 76.950 241.050 77.400 ;
        RECT 244.950 78.600 247.050 79.050 ;
        RECT 251.400 78.600 252.600 80.400 ;
        RECT 271.950 79.950 274.050 80.400 ;
        RECT 301.950 79.950 304.050 80.400 ;
        RECT 304.950 81.600 307.050 82.050 ;
        RECT 325.950 81.600 328.050 82.050 ;
        RECT 304.950 80.400 328.050 81.600 ;
        RECT 304.950 79.950 307.050 80.400 ;
        RECT 325.950 79.950 328.050 80.400 ;
        RECT 400.950 81.600 403.050 82.050 ;
        RECT 409.950 81.600 412.050 82.050 ;
        RECT 400.950 80.400 412.050 81.600 ;
        RECT 400.950 79.950 403.050 80.400 ;
        RECT 409.950 79.950 412.050 80.400 ;
        RECT 568.950 81.600 571.050 82.050 ;
        RECT 598.950 81.600 601.050 82.050 ;
        RECT 568.950 80.400 601.050 81.600 ;
        RECT 568.950 79.950 571.050 80.400 ;
        RECT 598.950 79.950 601.050 80.400 ;
        RECT 244.950 77.400 252.600 78.600 ;
        RECT 253.950 78.600 256.050 79.050 ;
        RECT 274.950 78.600 277.050 79.050 ;
        RECT 253.950 77.400 277.050 78.600 ;
        RECT 244.950 76.950 247.050 77.400 ;
        RECT 253.950 76.950 256.050 77.400 ;
        RECT 274.950 76.950 277.050 77.400 ;
        RECT 307.950 78.600 310.050 79.050 ;
        RECT 319.950 78.600 322.050 79.050 ;
        RECT 307.950 77.400 322.050 78.600 ;
        RECT 307.950 76.950 310.050 77.400 ;
        RECT 319.950 76.950 322.050 77.400 ;
        RECT 670.950 78.600 673.050 79.050 ;
        RECT 703.950 78.600 706.050 79.050 ;
        RECT 670.950 77.400 706.050 78.600 ;
        RECT 670.950 76.950 673.050 77.400 ;
        RECT 703.950 76.950 706.050 77.400 ;
        RECT 52.950 75.600 55.050 76.050 ;
        RECT 64.950 75.600 67.050 76.050 ;
        RECT 52.950 74.400 67.050 75.600 ;
        RECT 52.950 73.950 55.050 74.400 ;
        RECT 64.950 73.950 67.050 74.400 ;
        RECT 181.950 75.600 184.050 76.050 ;
        RECT 259.950 75.600 262.050 76.050 ;
        RECT 181.950 74.400 262.050 75.600 ;
        RECT 181.950 73.950 184.050 74.400 ;
        RECT 259.950 73.950 262.050 74.400 ;
        RECT 274.950 75.600 277.050 76.050 ;
        RECT 361.950 75.600 364.050 76.050 ;
        RECT 274.950 74.400 364.050 75.600 ;
        RECT 274.950 73.950 277.050 74.400 ;
        RECT 361.950 73.950 364.050 74.400 ;
        RECT 64.950 72.600 67.050 73.050 ;
        RECT 73.950 72.600 76.050 73.050 ;
        RECT 64.950 71.400 76.050 72.600 ;
        RECT 64.950 70.950 67.050 71.400 ;
        RECT 73.950 70.950 76.050 71.400 ;
        RECT 256.950 72.600 259.050 73.050 ;
        RECT 265.950 72.600 268.050 73.050 ;
        RECT 256.950 71.400 268.050 72.600 ;
        RECT 256.950 70.950 259.050 71.400 ;
        RECT 265.950 70.950 268.050 71.400 ;
        RECT 268.950 72.600 271.050 73.050 ;
        RECT 298.950 72.600 301.050 73.050 ;
        RECT 268.950 71.400 301.050 72.600 ;
        RECT 268.950 70.950 271.050 71.400 ;
        RECT 298.950 70.950 301.050 71.400 ;
        RECT 319.950 72.600 322.050 73.050 ;
        RECT 325.950 72.600 328.050 73.050 ;
        RECT 343.950 72.600 346.050 73.050 ;
        RECT 319.950 71.400 346.050 72.600 ;
        RECT 319.950 70.950 322.050 71.400 ;
        RECT 325.950 70.950 328.050 71.400 ;
        RECT 343.950 70.950 346.050 71.400 ;
        RECT 46.950 69.600 49.050 70.050 ;
        RECT 76.950 69.600 79.050 70.050 ;
        RECT 130.950 69.600 133.050 70.050 ;
        RECT 46.950 68.400 133.050 69.600 ;
        RECT 46.950 67.950 49.050 68.400 ;
        RECT 76.950 67.950 79.050 68.400 ;
        RECT 130.950 67.950 133.050 68.400 ;
        RECT 208.950 69.600 211.050 70.050 ;
        RECT 280.950 69.600 283.050 70.050 ;
        RECT 208.950 68.400 283.050 69.600 ;
        RECT 208.950 67.950 211.050 68.400 ;
        RECT 280.950 67.950 283.050 68.400 ;
        RECT 286.950 69.600 289.050 70.050 ;
        RECT 328.950 69.600 331.050 70.050 ;
        RECT 286.950 68.400 331.050 69.600 ;
        RECT 286.950 67.950 289.050 68.400 ;
        RECT 328.950 67.950 331.050 68.400 ;
        RECT 58.950 66.600 61.050 67.050 ;
        RECT 94.950 66.600 97.050 67.050 ;
        RECT 58.950 65.400 97.050 66.600 ;
        RECT 58.950 64.950 61.050 65.400 ;
        RECT 94.950 64.950 97.050 65.400 ;
        RECT 202.950 66.600 205.050 67.050 ;
        RECT 238.950 66.600 241.050 67.050 ;
        RECT 277.950 66.600 280.050 67.050 ;
        RECT 202.950 65.400 280.050 66.600 ;
        RECT 202.950 64.950 205.050 65.400 ;
        RECT 238.950 64.950 241.050 65.400 ;
        RECT 277.950 64.950 280.050 65.400 ;
        RECT 286.950 66.600 289.050 67.050 ;
        RECT 340.950 66.600 343.050 67.050 ;
        RECT 286.950 65.400 343.050 66.600 ;
        RECT 286.950 64.950 289.050 65.400 ;
        RECT 340.950 64.950 343.050 65.400 ;
        RECT 34.950 63.600 37.050 64.050 ;
        RECT 49.950 63.600 52.050 64.050 ;
        RECT 34.950 62.400 52.050 63.600 ;
        RECT 34.950 61.950 37.050 62.400 ;
        RECT 49.950 61.950 52.050 62.400 ;
        RECT 79.950 63.600 82.050 64.050 ;
        RECT 88.950 63.600 91.050 64.050 ;
        RECT 79.950 62.400 91.050 63.600 ;
        RECT 79.950 61.950 82.050 62.400 ;
        RECT 88.950 61.950 91.050 62.400 ;
        RECT 130.950 63.600 133.050 64.050 ;
        RECT 148.950 63.600 151.050 64.050 ;
        RECT 130.950 62.400 151.050 63.600 ;
        RECT 130.950 61.950 133.050 62.400 ;
        RECT 148.950 61.950 151.050 62.400 ;
        RECT 169.950 63.600 172.050 64.050 ;
        RECT 202.950 63.600 205.050 64.050 ;
        RECT 169.950 62.400 205.050 63.600 ;
        RECT 169.950 61.950 172.050 62.400 ;
        RECT 202.950 61.950 205.050 62.400 ;
        RECT 205.950 63.600 208.050 64.050 ;
        RECT 253.950 63.600 256.050 64.050 ;
        RECT 205.950 62.400 256.050 63.600 ;
        RECT 205.950 61.950 208.050 62.400 ;
        RECT 253.950 61.950 256.050 62.400 ;
        RECT 256.950 63.600 259.050 64.050 ;
        RECT 283.950 63.600 286.050 64.050 ;
        RECT 256.950 62.400 286.050 63.600 ;
        RECT 256.950 61.950 259.050 62.400 ;
        RECT 283.950 61.950 286.050 62.400 ;
        RECT 304.950 63.600 307.050 64.050 ;
        RECT 316.950 63.600 319.050 64.050 ;
        RECT 361.950 63.600 364.050 64.050 ;
        RECT 304.950 62.400 364.050 63.600 ;
        RECT 304.950 61.950 307.050 62.400 ;
        RECT 316.950 61.950 319.050 62.400 ;
        RECT 361.950 61.950 364.050 62.400 ;
        RECT 382.950 63.600 385.050 64.050 ;
        RECT 394.950 63.600 397.050 64.050 ;
        RECT 430.950 63.600 433.050 64.050 ;
        RECT 382.950 62.400 433.050 63.600 ;
        RECT 382.950 61.950 385.050 62.400 ;
        RECT 394.950 61.950 397.050 62.400 ;
        RECT 430.950 61.950 433.050 62.400 ;
        RECT 520.950 63.600 523.050 64.050 ;
        RECT 583.950 63.600 586.050 64.050 ;
        RECT 643.950 63.600 646.050 64.050 ;
        RECT 670.950 63.600 673.050 64.050 ;
        RECT 679.950 63.600 682.050 64.050 ;
        RECT 520.950 62.400 682.050 63.600 ;
        RECT 520.950 61.950 523.050 62.400 ;
        RECT 583.950 61.950 586.050 62.400 ;
        RECT 643.950 61.950 646.050 62.400 ;
        RECT 670.950 61.950 673.050 62.400 ;
        RECT 679.950 61.950 682.050 62.400 ;
        RECT 13.950 60.600 16.050 61.050 ;
        RECT 64.950 60.600 67.050 61.050 ;
        RECT 13.950 59.400 67.050 60.600 ;
        RECT 13.950 58.950 16.050 59.400 ;
        RECT 64.950 58.950 67.050 59.400 ;
        RECT 67.950 60.600 70.050 61.050 ;
        RECT 97.950 60.600 100.050 61.050 ;
        RECT 67.950 59.400 100.050 60.600 ;
        RECT 67.950 58.950 70.050 59.400 ;
        RECT 97.950 58.950 100.050 59.400 ;
        RECT 103.950 60.600 106.050 61.050 ;
        RECT 127.950 60.600 130.050 61.050 ;
        RECT 139.950 60.600 142.050 61.050 ;
        RECT 175.950 60.600 178.050 61.050 ;
        RECT 103.950 59.400 178.050 60.600 ;
        RECT 103.950 58.950 106.050 59.400 ;
        RECT 127.950 58.950 130.050 59.400 ;
        RECT 139.950 58.950 142.050 59.400 ;
        RECT 175.950 58.950 178.050 59.400 ;
        RECT 217.950 60.600 220.050 61.050 ;
        RECT 244.950 60.600 247.050 61.050 ;
        RECT 217.950 59.400 247.050 60.600 ;
        RECT 217.950 58.950 220.050 59.400 ;
        RECT 244.950 58.950 247.050 59.400 ;
        RECT 271.950 60.600 274.050 61.050 ;
        RECT 286.950 60.600 289.050 61.050 ;
        RECT 271.950 59.400 289.050 60.600 ;
        RECT 271.950 58.950 274.050 59.400 ;
        RECT 286.950 58.950 289.050 59.400 ;
        RECT 292.950 60.600 295.050 61.050 ;
        RECT 349.950 60.600 352.050 61.050 ;
        RECT 292.950 59.400 352.050 60.600 ;
        RECT 292.950 58.950 295.050 59.400 ;
        RECT 349.950 58.950 352.050 59.400 ;
        RECT 385.950 60.600 388.050 61.050 ;
        RECT 403.950 60.600 406.050 61.050 ;
        RECT 385.950 59.400 406.050 60.600 ;
        RECT 385.950 58.950 388.050 59.400 ;
        RECT 403.950 58.950 406.050 59.400 ;
        RECT 412.950 60.600 415.050 61.050 ;
        RECT 541.950 60.600 544.050 61.050 ;
        RECT 412.950 59.400 544.050 60.600 ;
        RECT 412.950 58.950 415.050 59.400 ;
        RECT 541.950 58.950 544.050 59.400 ;
        RECT 544.950 60.600 547.050 61.050 ;
        RECT 568.950 60.600 571.050 61.050 ;
        RECT 544.950 59.400 571.050 60.600 ;
        RECT 544.950 58.950 547.050 59.400 ;
        RECT 568.950 58.950 571.050 59.400 ;
        RECT 640.950 60.600 643.050 61.050 ;
        RECT 652.950 60.600 655.050 61.050 ;
        RECT 640.950 59.400 655.050 60.600 ;
        RECT 640.950 58.950 643.050 59.400 ;
        RECT 652.950 58.950 655.050 59.400 ;
        RECT 22.950 57.600 25.050 58.050 ;
        RECT 28.950 57.600 31.050 58.050 ;
        RECT 52.950 57.600 55.050 58.050 ;
        RECT 22.950 56.400 31.050 57.600 ;
        RECT 22.950 55.950 25.050 56.400 ;
        RECT 28.950 55.950 31.050 56.400 ;
        RECT 47.400 56.400 55.050 57.600 ;
        RECT 31.950 54.600 34.050 55.050 ;
        RECT 37.950 54.600 40.050 55.050 ;
        RECT 31.950 53.400 40.050 54.600 ;
        RECT 31.950 52.950 34.050 53.400 ;
        RECT 37.950 52.950 40.050 53.400 ;
        RECT 47.400 52.050 48.600 56.400 ;
        RECT 52.950 55.950 55.050 56.400 ;
        RECT 55.950 57.600 58.050 58.050 ;
        RECT 67.950 57.600 70.050 58.050 ;
        RECT 55.950 56.400 70.050 57.600 ;
        RECT 55.950 55.950 58.050 56.400 ;
        RECT 67.950 55.950 70.050 56.400 ;
        RECT 73.950 57.600 76.050 58.050 ;
        RECT 73.950 56.400 108.600 57.600 ;
        RECT 73.950 55.950 76.050 56.400 ;
        RECT 58.950 54.600 61.050 55.050 ;
        RECT 88.950 54.600 91.050 55.050 ;
        RECT 58.950 53.400 91.050 54.600 ;
        RECT 58.950 52.950 61.050 53.400 ;
        RECT 88.950 52.950 91.050 53.400 ;
        RECT 107.400 52.050 108.600 56.400 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 133.950 57.600 136.050 58.050 ;
        RECT 166.950 57.600 169.050 58.050 ;
        RECT 133.950 56.400 150.600 57.600 ;
        RECT 133.950 55.950 136.050 56.400 ;
        RECT 115.950 52.950 118.050 55.050 ;
        RECT 125.400 54.600 126.600 55.950 ;
        RECT 142.950 54.600 145.050 55.050 ;
        RECT 125.400 53.400 145.050 54.600 ;
        RECT 142.950 52.950 145.050 53.400 ;
        RECT 13.950 51.600 16.050 52.050 ;
        RECT 25.950 51.600 28.050 52.050 ;
        RECT 43.950 51.600 46.050 52.050 ;
        RECT 13.950 50.400 46.050 51.600 ;
        RECT 13.950 49.950 16.050 50.400 ;
        RECT 25.950 49.950 28.050 50.400 ;
        RECT 43.950 49.950 46.050 50.400 ;
        RECT 46.950 49.950 49.050 52.050 ;
        RECT 61.950 51.600 64.050 52.050 ;
        RECT 106.950 51.600 109.050 52.050 ;
        RECT 61.950 50.400 109.050 51.600 ;
        RECT 61.950 49.950 64.050 50.400 ;
        RECT 106.950 49.950 109.050 50.400 ;
        RECT 10.950 48.600 13.050 49.050 ;
        RECT 37.950 48.600 40.050 49.050 ;
        RECT 52.950 48.600 55.050 49.050 ;
        RECT 10.950 47.400 55.050 48.600 ;
        RECT 10.950 46.950 13.050 47.400 ;
        RECT 37.950 46.950 40.050 47.400 ;
        RECT 52.950 46.950 55.050 47.400 ;
        RECT 64.950 48.600 67.050 49.050 ;
        RECT 70.950 48.600 73.050 49.050 ;
        RECT 64.950 47.400 73.050 48.600 ;
        RECT 64.950 46.950 67.050 47.400 ;
        RECT 70.950 46.950 73.050 47.400 ;
        RECT 76.950 48.600 79.050 49.050 ;
        RECT 94.950 48.600 97.050 49.050 ;
        RECT 76.950 47.400 97.050 48.600 ;
        RECT 76.950 46.950 79.050 47.400 ;
        RECT 94.950 46.950 97.050 47.400 ;
        RECT 103.950 48.600 106.050 49.050 ;
        RECT 116.400 48.600 117.600 52.950 ;
        RECT 149.400 51.600 150.600 56.400 ;
        RECT 166.950 56.400 186.600 57.600 ;
        RECT 166.950 55.950 169.050 56.400 ;
        RECT 151.950 54.600 154.050 55.050 ;
        RECT 169.950 54.600 172.050 55.050 ;
        RECT 151.950 53.400 172.050 54.600 ;
        RECT 151.950 52.950 154.050 53.400 ;
        RECT 169.950 52.950 172.050 53.400 ;
        RECT 185.400 52.050 186.600 56.400 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 57.600 193.050 58.050 ;
        RECT 199.950 57.600 202.050 58.050 ;
        RECT 190.950 56.400 202.050 57.600 ;
        RECT 190.950 55.950 193.050 56.400 ;
        RECT 199.950 55.950 202.050 56.400 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 235.950 57.600 238.050 58.050 ;
        RECT 250.950 57.600 253.050 58.050 ;
        RECT 235.950 56.400 249.600 57.600 ;
        RECT 235.950 55.950 238.050 56.400 ;
        RECT 188.400 52.050 189.600 55.950 ;
        RECT 196.950 54.600 199.050 55.050 ;
        RECT 202.950 54.600 205.050 55.050 ;
        RECT 196.950 53.400 205.050 54.600 ;
        RECT 196.950 52.950 199.050 53.400 ;
        RECT 202.950 52.950 205.050 53.400 ;
        RECT 208.950 54.600 211.050 55.050 ;
        RECT 229.950 54.600 232.050 55.050 ;
        RECT 208.950 53.400 213.600 54.600 ;
        RECT 208.950 52.950 211.050 53.400 ;
        RECT 212.400 52.050 213.600 53.400 ;
        RECT 218.400 53.400 232.050 54.600 ;
        RECT 172.950 51.600 175.050 52.050 ;
        RECT 149.400 50.400 175.050 51.600 ;
        RECT 172.950 49.950 175.050 50.400 ;
        RECT 184.950 49.950 187.050 52.050 ;
        RECT 187.950 49.950 190.050 52.050 ;
        RECT 211.950 49.950 214.050 52.050 ;
        RECT 218.400 49.050 219.600 53.400 ;
        RECT 229.950 52.950 232.050 53.400 ;
        RECT 220.950 51.600 223.050 52.050 ;
        RECT 233.400 51.600 234.600 55.950 ;
        RECT 244.950 52.950 247.050 55.050 ;
        RECT 220.950 50.400 234.600 51.600 ;
        RECT 220.950 49.950 223.050 50.400 ;
        RECT 103.950 47.400 117.600 48.600 ;
        RECT 118.950 48.600 121.050 49.050 ;
        RECT 136.950 48.600 139.050 49.050 ;
        RECT 118.950 47.400 139.050 48.600 ;
        RECT 103.950 46.950 106.050 47.400 ;
        RECT 118.950 46.950 121.050 47.400 ;
        RECT 136.950 46.950 139.050 47.400 ;
        RECT 157.950 48.600 160.050 49.050 ;
        RECT 166.950 48.600 169.050 49.050 ;
        RECT 157.950 47.400 169.050 48.600 ;
        RECT 157.950 46.950 160.050 47.400 ;
        RECT 166.950 46.950 169.050 47.400 ;
        RECT 175.950 48.600 178.050 49.050 ;
        RECT 211.950 48.600 214.050 49.050 ;
        RECT 175.950 47.400 214.050 48.600 ;
        RECT 175.950 46.950 178.050 47.400 ;
        RECT 211.950 46.950 214.050 47.400 ;
        RECT 217.950 46.950 220.050 49.050 ;
        RECT 220.950 48.600 223.050 49.050 ;
        RECT 245.400 48.600 246.600 52.950 ;
        RECT 220.950 47.400 246.600 48.600 ;
        RECT 248.400 48.600 249.600 56.400 ;
        RECT 250.950 56.400 267.600 57.600 ;
        RECT 250.950 55.950 253.050 56.400 ;
        RECT 250.950 54.600 253.050 55.050 ;
        RECT 256.950 54.600 259.050 55.050 ;
        RECT 262.950 54.600 265.050 55.050 ;
        RECT 250.950 53.400 265.050 54.600 ;
        RECT 250.950 52.950 253.050 53.400 ;
        RECT 256.950 52.950 259.050 53.400 ;
        RECT 262.950 52.950 265.050 53.400 ;
        RECT 259.950 51.600 262.050 52.050 ;
        RECT 266.400 51.600 267.600 56.400 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 349.950 57.600 352.050 58.050 ;
        RECT 373.950 57.600 376.050 58.050 ;
        RECT 379.950 57.600 382.050 58.050 ;
        RECT 409.950 57.600 412.050 58.050 ;
        RECT 349.950 56.400 366.600 57.600 ;
        RECT 349.950 55.950 352.050 56.400 ;
        RECT 280.950 54.600 283.050 55.050 ;
        RECT 301.950 54.600 304.050 55.050 ;
        RECT 307.950 54.600 310.050 55.050 ;
        RECT 280.950 53.400 310.050 54.600 ;
        RECT 280.950 52.950 283.050 53.400 ;
        RECT 301.950 52.950 304.050 53.400 ;
        RECT 307.950 52.950 310.050 53.400 ;
        RECT 259.950 50.400 267.600 51.600 ;
        RECT 274.950 51.600 277.050 52.050 ;
        RECT 286.950 51.600 289.050 52.050 ;
        RECT 274.950 50.400 289.050 51.600 ;
        RECT 259.950 49.950 262.050 50.400 ;
        RECT 274.950 49.950 277.050 50.400 ;
        RECT 286.950 49.950 289.050 50.400 ;
        RECT 307.950 51.600 310.050 52.050 ;
        RECT 311.400 51.600 312.600 55.950 ;
        RECT 365.400 55.050 366.600 56.400 ;
        RECT 373.950 56.400 382.050 57.600 ;
        RECT 373.950 55.950 376.050 56.400 ;
        RECT 379.950 55.950 382.050 56.400 ;
        RECT 383.400 56.400 412.050 57.600 ;
        RECT 319.950 54.600 322.050 55.050 ;
        RECT 328.950 54.600 331.050 55.050 ;
        RECT 319.950 53.400 331.050 54.600 ;
        RECT 319.950 52.950 322.050 53.400 ;
        RECT 328.950 52.950 331.050 53.400 ;
        RECT 334.950 54.600 337.050 55.050 ;
        RECT 334.950 53.400 357.600 54.600 ;
        RECT 334.950 52.950 337.050 53.400 ;
        RECT 340.950 51.600 343.050 52.050 ;
        RECT 307.950 50.400 343.050 51.600 ;
        RECT 307.950 49.950 310.050 50.400 ;
        RECT 340.950 49.950 343.050 50.400 ;
        RECT 346.950 51.600 349.050 52.050 ;
        RECT 352.950 51.600 355.050 52.050 ;
        RECT 346.950 50.400 355.050 51.600 ;
        RECT 356.400 51.600 357.600 53.400 ;
        RECT 364.950 52.950 367.050 55.050 ;
        RECT 383.400 54.600 384.600 56.400 ;
        RECT 401.400 55.050 402.600 56.400 ;
        RECT 409.950 55.950 412.050 56.400 ;
        RECT 427.950 57.600 430.050 58.050 ;
        RECT 433.950 57.600 436.050 58.050 ;
        RECT 427.950 56.400 436.050 57.600 ;
        RECT 427.950 55.950 430.050 56.400 ;
        RECT 433.950 55.950 436.050 56.400 ;
        RECT 439.950 57.600 442.050 58.050 ;
        RECT 451.950 57.600 454.050 58.050 ;
        RECT 466.950 57.600 469.050 58.050 ;
        RECT 502.950 57.600 505.050 58.050 ;
        RECT 439.950 56.400 469.050 57.600 ;
        RECT 439.950 55.950 442.050 56.400 ;
        RECT 451.950 55.950 454.050 56.400 ;
        RECT 466.950 55.950 469.050 56.400 ;
        RECT 497.400 56.400 505.050 57.600 ;
        RECT 497.400 55.050 498.600 56.400 ;
        RECT 502.950 55.950 505.050 56.400 ;
        RECT 508.950 57.600 511.050 58.050 ;
        RECT 520.950 57.600 523.050 58.050 ;
        RECT 508.950 56.400 523.050 57.600 ;
        RECT 508.950 55.950 511.050 56.400 ;
        RECT 520.950 55.950 523.050 56.400 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 646.950 57.600 649.050 58.050 ;
        RECT 655.950 57.600 658.050 58.050 ;
        RECT 646.950 56.400 658.050 57.600 ;
        RECT 646.950 55.950 649.050 56.400 ;
        RECT 655.950 55.950 658.050 56.400 ;
        RECT 368.400 53.400 384.600 54.600 ;
        RECT 385.950 54.600 388.050 55.050 ;
        RECT 394.950 54.600 397.050 55.050 ;
        RECT 385.950 53.400 397.050 54.600 ;
        RECT 364.950 51.600 367.050 52.050 ;
        RECT 356.400 50.400 367.050 51.600 ;
        RECT 346.950 49.950 349.050 50.400 ;
        RECT 352.950 49.950 355.050 50.400 ;
        RECT 364.950 49.950 367.050 50.400 ;
        RECT 250.950 48.600 253.050 49.050 ;
        RECT 248.400 47.400 253.050 48.600 ;
        RECT 220.950 46.950 223.050 47.400 ;
        RECT 250.950 46.950 253.050 47.400 ;
        RECT 253.950 48.600 256.050 49.050 ;
        RECT 277.950 48.600 280.050 49.050 ;
        RECT 253.950 47.400 280.050 48.600 ;
        RECT 253.950 46.950 256.050 47.400 ;
        RECT 277.950 46.950 280.050 47.400 ;
        RECT 301.950 48.600 304.050 49.050 ;
        RECT 331.950 48.600 334.050 49.050 ;
        RECT 301.950 47.400 334.050 48.600 ;
        RECT 301.950 46.950 304.050 47.400 ;
        RECT 331.950 46.950 334.050 47.400 ;
        RECT 355.950 48.600 358.050 49.050 ;
        RECT 368.400 48.600 369.600 53.400 ;
        RECT 385.950 52.950 388.050 53.400 ;
        RECT 394.950 52.950 397.050 53.400 ;
        RECT 400.950 52.950 403.050 55.050 ;
        RECT 415.950 54.600 418.050 55.050 ;
        RECT 404.400 53.400 418.050 54.600 ;
        RECT 370.950 51.600 373.050 52.050 ;
        RECT 404.400 51.600 405.600 53.400 ;
        RECT 415.950 52.950 418.050 53.400 ;
        RECT 436.950 54.600 439.050 55.050 ;
        RECT 460.950 54.600 463.050 55.050 ;
        RECT 436.950 53.400 463.050 54.600 ;
        RECT 436.950 52.950 439.050 53.400 ;
        RECT 460.950 52.950 463.050 53.400 ;
        RECT 496.950 52.950 499.050 55.050 ;
        RECT 502.950 52.950 505.050 55.050 ;
        RECT 514.950 52.950 517.050 55.050 ;
        RECT 553.950 54.600 556.050 55.050 ;
        RECT 563.400 54.600 564.600 55.950 ;
        RECT 553.950 53.400 564.600 54.600 ;
        RECT 565.950 54.600 568.050 55.050 ;
        RECT 574.950 54.600 577.050 55.050 ;
        RECT 565.950 53.400 577.050 54.600 ;
        RECT 553.950 52.950 556.050 53.400 ;
        RECT 565.950 52.950 568.050 53.400 ;
        RECT 574.950 52.950 577.050 53.400 ;
        RECT 610.950 54.600 613.050 55.050 ;
        RECT 649.950 54.600 652.050 55.050 ;
        RECT 610.950 53.400 652.050 54.600 ;
        RECT 610.950 52.950 613.050 53.400 ;
        RECT 649.950 52.950 652.050 53.400 ;
        RECT 664.950 54.600 667.050 55.050 ;
        RECT 673.950 54.600 676.050 55.050 ;
        RECT 664.950 53.400 676.050 54.600 ;
        RECT 664.950 52.950 667.050 53.400 ;
        RECT 673.950 52.950 676.050 53.400 ;
        RECT 370.950 50.400 405.600 51.600 ;
        RECT 412.950 51.600 415.050 52.050 ;
        RECT 418.950 51.600 421.050 52.050 ;
        RECT 412.950 50.400 421.050 51.600 ;
        RECT 370.950 49.950 373.050 50.400 ;
        RECT 412.950 49.950 415.050 50.400 ;
        RECT 418.950 49.950 421.050 50.400 ;
        RECT 424.950 51.600 427.050 52.050 ;
        RECT 430.950 51.600 433.050 52.050 ;
        RECT 424.950 50.400 433.050 51.600 ;
        RECT 424.950 49.950 427.050 50.400 ;
        RECT 430.950 49.950 433.050 50.400 ;
        RECT 469.950 51.600 472.050 52.050 ;
        RECT 475.950 51.600 478.050 52.050 ;
        RECT 469.950 50.400 478.050 51.600 ;
        RECT 469.950 49.950 472.050 50.400 ;
        RECT 475.950 49.950 478.050 50.400 ;
        RECT 484.950 51.600 487.050 52.050 ;
        RECT 503.400 51.600 504.600 52.950 ;
        RECT 484.950 50.400 504.600 51.600 ;
        RECT 515.400 51.600 516.600 52.950 ;
        RECT 526.950 51.600 529.050 52.050 ;
        RECT 515.400 50.400 529.050 51.600 ;
        RECT 484.950 49.950 487.050 50.400 ;
        RECT 526.950 49.950 529.050 50.400 ;
        RECT 541.950 51.600 544.050 52.050 ;
        RECT 577.950 51.600 580.050 52.050 ;
        RECT 541.950 50.400 580.050 51.600 ;
        RECT 541.950 49.950 544.050 50.400 ;
        RECT 577.950 49.950 580.050 50.400 ;
        RECT 610.950 51.600 613.050 52.050 ;
        RECT 616.950 51.600 619.050 52.050 ;
        RECT 610.950 50.400 619.050 51.600 ;
        RECT 610.950 49.950 613.050 50.400 ;
        RECT 616.950 49.950 619.050 50.400 ;
        RECT 637.950 51.600 640.050 52.050 ;
        RECT 658.950 51.600 661.050 52.050 ;
        RECT 637.950 50.400 661.050 51.600 ;
        RECT 637.950 49.950 640.050 50.400 ;
        RECT 658.950 49.950 661.050 50.400 ;
        RECT 355.950 47.400 369.600 48.600 ;
        RECT 397.950 48.600 400.050 49.050 ;
        RECT 406.950 48.600 409.050 49.050 ;
        RECT 397.950 47.400 409.050 48.600 ;
        RECT 355.950 46.950 358.050 47.400 ;
        RECT 397.950 46.950 400.050 47.400 ;
        RECT 406.950 46.950 409.050 47.400 ;
        RECT 421.950 48.600 424.050 49.050 ;
        RECT 427.950 48.600 430.050 49.050 ;
        RECT 421.950 47.400 430.050 48.600 ;
        RECT 421.950 46.950 424.050 47.400 ;
        RECT 427.950 46.950 430.050 47.400 ;
        RECT 457.950 48.600 460.050 49.050 ;
        RECT 511.950 48.600 514.050 49.050 ;
        RECT 457.950 47.400 514.050 48.600 ;
        RECT 457.950 46.950 460.050 47.400 ;
        RECT 511.950 46.950 514.050 47.400 ;
        RECT 517.950 48.600 520.050 49.050 ;
        RECT 529.950 48.600 532.050 49.050 ;
        RECT 538.950 48.600 541.050 49.050 ;
        RECT 547.950 48.600 550.050 49.050 ;
        RECT 517.950 47.400 550.050 48.600 ;
        RECT 517.950 46.950 520.050 47.400 ;
        RECT 529.950 46.950 532.050 47.400 ;
        RECT 538.950 46.950 541.050 47.400 ;
        RECT 547.950 46.950 550.050 47.400 ;
        RECT 604.950 48.600 607.050 49.050 ;
        RECT 619.950 48.600 622.050 49.050 ;
        RECT 604.950 47.400 622.050 48.600 ;
        RECT 604.950 46.950 607.050 47.400 ;
        RECT 619.950 46.950 622.050 47.400 ;
        RECT 670.950 48.600 673.050 49.050 ;
        RECT 674.400 48.600 675.600 52.950 ;
        RECT 670.950 47.400 675.600 48.600 ;
        RECT 670.950 46.950 673.050 47.400 ;
        RECT 70.950 45.600 73.050 46.050 ;
        RECT 112.950 45.600 115.050 46.050 ;
        RECT 70.950 44.400 115.050 45.600 ;
        RECT 70.950 43.950 73.050 44.400 ;
        RECT 112.950 43.950 115.050 44.400 ;
        RECT 121.950 45.600 124.050 46.050 ;
        RECT 154.950 45.600 157.050 46.050 ;
        RECT 169.950 45.600 172.050 46.050 ;
        RECT 121.950 44.400 172.050 45.600 ;
        RECT 121.950 43.950 124.050 44.400 ;
        RECT 154.950 43.950 157.050 44.400 ;
        RECT 169.950 43.950 172.050 44.400 ;
        RECT 187.950 45.600 190.050 46.050 ;
        RECT 223.950 45.600 226.050 46.050 ;
        RECT 253.950 45.600 256.050 46.050 ;
        RECT 187.950 44.400 256.050 45.600 ;
        RECT 187.950 43.950 190.050 44.400 ;
        RECT 223.950 43.950 226.050 44.400 ;
        RECT 253.950 43.950 256.050 44.400 ;
        RECT 262.950 45.600 265.050 46.050 ;
        RECT 292.950 45.600 295.050 46.050 ;
        RECT 262.950 44.400 295.050 45.600 ;
        RECT 262.950 43.950 265.050 44.400 ;
        RECT 292.950 43.950 295.050 44.400 ;
        RECT 298.950 45.600 301.050 46.050 ;
        RECT 304.950 45.600 307.050 46.050 ;
        RECT 298.950 44.400 307.050 45.600 ;
        RECT 298.950 43.950 301.050 44.400 ;
        RECT 304.950 43.950 307.050 44.400 ;
        RECT 319.950 45.600 322.050 46.050 ;
        RECT 337.950 45.600 340.050 46.050 ;
        RECT 358.950 45.600 361.050 46.050 ;
        RECT 319.950 44.400 361.050 45.600 ;
        RECT 319.950 43.950 322.050 44.400 ;
        RECT 337.950 43.950 340.050 44.400 ;
        RECT 358.950 43.950 361.050 44.400 ;
        RECT 379.950 45.600 382.050 46.050 ;
        RECT 445.950 45.600 448.050 46.050 ;
        RECT 379.950 44.400 448.050 45.600 ;
        RECT 379.950 43.950 382.050 44.400 ;
        RECT 445.950 43.950 448.050 44.400 ;
        RECT 463.950 45.600 466.050 46.050 ;
        RECT 502.950 45.600 505.050 46.050 ;
        RECT 463.950 44.400 505.050 45.600 ;
        RECT 463.950 43.950 466.050 44.400 ;
        RECT 502.950 43.950 505.050 44.400 ;
        RECT 523.950 45.600 526.050 46.050 ;
        RECT 535.950 45.600 538.050 46.050 ;
        RECT 559.950 45.600 562.050 46.050 ;
        RECT 589.950 45.600 592.050 46.050 ;
        RECT 523.950 44.400 592.050 45.600 ;
        RECT 523.950 43.950 526.050 44.400 ;
        RECT 535.950 43.950 538.050 44.400 ;
        RECT 559.950 43.950 562.050 44.400 ;
        RECT 589.950 43.950 592.050 44.400 ;
        RECT 595.950 45.600 598.050 46.050 ;
        RECT 616.950 45.600 619.050 46.050 ;
        RECT 595.950 44.400 619.050 45.600 ;
        RECT 595.950 43.950 598.050 44.400 ;
        RECT 616.950 43.950 619.050 44.400 ;
        RECT 661.950 45.600 664.050 46.050 ;
        RECT 700.950 45.600 703.050 46.050 ;
        RECT 661.950 44.400 703.050 45.600 ;
        RECT 661.950 43.950 664.050 44.400 ;
        RECT 700.950 43.950 703.050 44.400 ;
        RECT 52.950 42.600 55.050 43.050 ;
        RECT 142.950 42.600 145.050 43.050 ;
        RECT 52.950 41.400 145.050 42.600 ;
        RECT 52.950 40.950 55.050 41.400 ;
        RECT 142.950 40.950 145.050 41.400 ;
        RECT 178.950 42.600 181.050 43.050 ;
        RECT 199.950 42.600 202.050 43.050 ;
        RECT 214.950 42.600 217.050 43.050 ;
        RECT 229.950 42.600 232.050 43.050 ;
        RECT 178.950 41.400 232.050 42.600 ;
        RECT 178.950 40.950 181.050 41.400 ;
        RECT 199.950 40.950 202.050 41.400 ;
        RECT 214.950 40.950 217.050 41.400 ;
        RECT 229.950 40.950 232.050 41.400 ;
        RECT 238.950 42.600 241.050 43.050 ;
        RECT 268.950 42.600 271.050 43.050 ;
        RECT 238.950 41.400 271.050 42.600 ;
        RECT 238.950 40.950 241.050 41.400 ;
        RECT 268.950 40.950 271.050 41.400 ;
        RECT 328.950 42.600 331.050 43.050 ;
        RECT 337.950 42.600 340.050 43.050 ;
        RECT 328.950 41.400 340.050 42.600 ;
        RECT 328.950 40.950 331.050 41.400 ;
        RECT 337.950 40.950 340.050 41.400 ;
        RECT 478.950 42.600 481.050 43.050 ;
        RECT 526.950 42.600 529.050 43.050 ;
        RECT 478.950 41.400 529.050 42.600 ;
        RECT 478.950 40.950 481.050 41.400 ;
        RECT 526.950 40.950 529.050 41.400 ;
        RECT 580.950 42.600 583.050 43.050 ;
        RECT 628.950 42.600 631.050 43.050 ;
        RECT 580.950 41.400 631.050 42.600 ;
        RECT 580.950 40.950 583.050 41.400 ;
        RECT 628.950 40.950 631.050 41.400 ;
        RECT 52.950 39.600 55.050 40.050 ;
        RECT 82.950 39.600 85.050 40.050 ;
        RECT 52.950 38.400 85.050 39.600 ;
        RECT 52.950 37.950 55.050 38.400 ;
        RECT 82.950 37.950 85.050 38.400 ;
        RECT 136.950 39.600 139.050 40.050 ;
        RECT 205.950 39.600 208.050 40.050 ;
        RECT 136.950 38.400 208.050 39.600 ;
        RECT 136.950 37.950 139.050 38.400 ;
        RECT 205.950 37.950 208.050 38.400 ;
        RECT 208.950 39.600 211.050 40.050 ;
        RECT 220.950 39.600 223.050 40.050 ;
        RECT 208.950 38.400 223.050 39.600 ;
        RECT 208.950 37.950 211.050 38.400 ;
        RECT 220.950 37.950 223.050 38.400 ;
        RECT 235.950 39.600 238.050 40.050 ;
        RECT 247.950 39.600 250.050 40.050 ;
        RECT 265.950 39.600 268.050 40.050 ;
        RECT 280.950 39.600 283.050 40.050 ;
        RECT 235.950 38.400 283.050 39.600 ;
        RECT 235.950 37.950 238.050 38.400 ;
        RECT 247.950 37.950 250.050 38.400 ;
        RECT 265.950 37.950 268.050 38.400 ;
        RECT 280.950 37.950 283.050 38.400 ;
        RECT 295.950 39.600 298.050 40.050 ;
        RECT 358.950 39.600 361.050 40.050 ;
        RECT 397.950 39.600 400.050 40.050 ;
        RECT 403.950 39.600 406.050 40.050 ;
        RECT 295.950 38.400 406.050 39.600 ;
        RECT 295.950 37.950 298.050 38.400 ;
        RECT 358.950 37.950 361.050 38.400 ;
        RECT 397.950 37.950 400.050 38.400 ;
        RECT 403.950 37.950 406.050 38.400 ;
        RECT 490.950 39.600 493.050 40.050 ;
        RECT 535.950 39.600 538.050 40.050 ;
        RECT 490.950 38.400 538.050 39.600 ;
        RECT 490.950 37.950 493.050 38.400 ;
        RECT 535.950 37.950 538.050 38.400 ;
        RECT 586.950 39.600 589.050 40.050 ;
        RECT 595.950 39.600 598.050 40.050 ;
        RECT 604.950 39.600 607.050 40.050 ;
        RECT 586.950 38.400 607.050 39.600 ;
        RECT 586.950 37.950 589.050 38.400 ;
        RECT 595.950 37.950 598.050 38.400 ;
        RECT 604.950 37.950 607.050 38.400 ;
        RECT 61.950 36.600 64.050 37.050 ;
        RECT 109.950 36.600 112.050 37.050 ;
        RECT 61.950 35.400 112.050 36.600 ;
        RECT 61.950 34.950 64.050 35.400 ;
        RECT 109.950 34.950 112.050 35.400 ;
        RECT 133.950 36.600 136.050 37.050 ;
        RECT 190.950 36.600 193.050 37.050 ;
        RECT 205.950 36.600 208.050 37.050 ;
        RECT 133.950 35.400 208.050 36.600 ;
        RECT 133.950 34.950 136.050 35.400 ;
        RECT 190.950 34.950 193.050 35.400 ;
        RECT 205.950 34.950 208.050 35.400 ;
        RECT 211.950 36.600 214.050 37.050 ;
        RECT 244.950 36.600 247.050 37.050 ;
        RECT 211.950 35.400 247.050 36.600 ;
        RECT 211.950 34.950 214.050 35.400 ;
        RECT 244.950 34.950 247.050 35.400 ;
        RECT 253.950 36.600 256.050 37.050 ;
        RECT 310.950 36.600 313.050 37.050 ;
        RECT 253.950 35.400 313.050 36.600 ;
        RECT 253.950 34.950 256.050 35.400 ;
        RECT 310.950 34.950 313.050 35.400 ;
        RECT 442.950 36.600 445.050 37.050 ;
        RECT 451.950 36.600 454.050 37.050 ;
        RECT 442.950 35.400 454.050 36.600 ;
        RECT 442.950 34.950 445.050 35.400 ;
        RECT 451.950 34.950 454.050 35.400 ;
        RECT 499.950 36.600 502.050 37.050 ;
        RECT 559.950 36.600 562.050 37.050 ;
        RECT 499.950 35.400 562.050 36.600 ;
        RECT 499.950 34.950 502.050 35.400 ;
        RECT 559.950 34.950 562.050 35.400 ;
        RECT 100.950 33.600 103.050 34.050 ;
        RECT 121.950 33.600 124.050 34.050 ;
        RECT 100.950 32.400 124.050 33.600 ;
        RECT 100.950 31.950 103.050 32.400 ;
        RECT 121.950 31.950 124.050 32.400 ;
        RECT 127.950 33.600 130.050 34.050 ;
        RECT 133.950 33.600 136.050 34.050 ;
        RECT 127.950 32.400 136.050 33.600 ;
        RECT 127.950 31.950 130.050 32.400 ;
        RECT 133.950 31.950 136.050 32.400 ;
        RECT 151.950 33.600 154.050 34.050 ;
        RECT 163.950 33.600 166.050 34.050 ;
        RECT 151.950 32.400 166.050 33.600 ;
        RECT 151.950 31.950 154.050 32.400 ;
        RECT 163.950 31.950 166.050 32.400 ;
        RECT 166.950 33.600 169.050 34.050 ;
        RECT 301.950 33.600 304.050 34.050 ;
        RECT 166.950 32.400 304.050 33.600 ;
        RECT 166.950 31.950 169.050 32.400 ;
        RECT 301.950 31.950 304.050 32.400 ;
        RECT 319.950 33.600 322.050 34.050 ;
        RECT 325.950 33.600 328.050 34.050 ;
        RECT 328.950 33.600 331.050 34.050 ;
        RECT 367.950 33.600 370.050 34.050 ;
        RECT 319.950 32.400 370.050 33.600 ;
        RECT 319.950 31.950 322.050 32.400 ;
        RECT 325.950 31.950 328.050 32.400 ;
        RECT 328.950 31.950 331.050 32.400 ;
        RECT 367.950 31.950 370.050 32.400 ;
        RECT 460.950 33.600 463.050 34.050 ;
        RECT 472.950 33.600 475.050 34.050 ;
        RECT 460.950 32.400 475.050 33.600 ;
        RECT 460.950 31.950 463.050 32.400 ;
        RECT 472.950 31.950 475.050 32.400 ;
        RECT 592.950 33.600 595.050 34.050 ;
        RECT 655.950 33.600 658.050 34.050 ;
        RECT 592.950 32.400 658.050 33.600 ;
        RECT 592.950 31.950 595.050 32.400 ;
        RECT 655.950 31.950 658.050 32.400 ;
        RECT 4.950 30.600 7.050 31.050 ;
        RECT 19.950 30.600 22.050 31.050 ;
        RECT 4.950 29.400 22.050 30.600 ;
        RECT 4.950 28.950 7.050 29.400 ;
        RECT 19.950 28.950 22.050 29.400 ;
        RECT 34.950 30.600 37.050 31.050 ;
        RECT 82.950 30.600 85.050 31.050 ;
        RECT 34.950 29.400 85.050 30.600 ;
        RECT 34.950 28.950 37.050 29.400 ;
        RECT 82.950 28.950 85.050 29.400 ;
        RECT 142.950 30.600 145.050 31.050 ;
        RECT 154.950 30.600 157.050 31.050 ;
        RECT 142.950 29.400 157.050 30.600 ;
        RECT 142.950 28.950 145.050 29.400 ;
        RECT 154.950 28.950 157.050 29.400 ;
        RECT 160.950 30.600 163.050 31.050 ;
        RECT 181.950 30.600 184.050 31.050 ;
        RECT 160.950 29.400 184.050 30.600 ;
        RECT 160.950 28.950 163.050 29.400 ;
        RECT 181.950 28.950 184.050 29.400 ;
        RECT 193.950 30.600 196.050 31.050 ;
        RECT 229.950 30.600 232.050 31.050 ;
        RECT 193.950 29.400 232.050 30.600 ;
        RECT 193.950 28.950 196.050 29.400 ;
        RECT 229.950 28.950 232.050 29.400 ;
        RECT 241.950 30.600 244.050 31.050 ;
        RECT 265.950 30.600 268.050 31.050 ;
        RECT 241.950 29.400 268.050 30.600 ;
        RECT 241.950 28.950 244.050 29.400 ;
        RECT 265.950 28.950 268.050 29.400 ;
        RECT 325.950 30.600 328.050 31.050 ;
        RECT 337.950 30.600 340.050 31.050 ;
        RECT 325.950 29.400 340.050 30.600 ;
        RECT 325.950 28.950 328.050 29.400 ;
        RECT 337.950 28.950 340.050 29.400 ;
        RECT 352.950 30.600 355.050 31.050 ;
        RECT 361.950 30.600 364.050 31.050 ;
        RECT 352.950 29.400 364.050 30.600 ;
        RECT 352.950 28.950 355.050 29.400 ;
        RECT 361.950 28.950 364.050 29.400 ;
        RECT 382.950 30.600 385.050 31.050 ;
        RECT 415.950 30.600 418.050 31.050 ;
        RECT 382.950 29.400 418.050 30.600 ;
        RECT 382.950 28.950 385.050 29.400 ;
        RECT 415.950 28.950 418.050 29.400 ;
        RECT 454.950 30.600 457.050 31.050 ;
        RECT 478.950 30.600 481.050 31.050 ;
        RECT 676.950 30.600 679.050 31.050 ;
        RECT 454.950 29.400 679.050 30.600 ;
        RECT 454.950 28.950 457.050 29.400 ;
        RECT 478.950 28.950 481.050 29.400 ;
        RECT 676.950 28.950 679.050 29.400 ;
        RECT 10.950 27.600 13.050 28.050 ;
        RECT 16.950 27.600 19.050 28.050 ;
        RECT 10.950 26.400 19.050 27.600 ;
        RECT 10.950 25.950 13.050 26.400 ;
        RECT 16.950 25.950 19.050 26.400 ;
        RECT 37.950 27.600 40.050 28.050 ;
        RECT 46.950 27.600 49.050 28.050 ;
        RECT 37.950 26.400 49.050 27.600 ;
        RECT 37.950 25.950 40.050 26.400 ;
        RECT 46.950 25.950 49.050 26.400 ;
        RECT 49.950 25.950 52.050 28.050 ;
        RECT 64.950 27.600 67.050 28.050 ;
        RECT 70.950 27.600 73.050 28.050 ;
        RECT 79.950 27.600 82.050 28.050 ;
        RECT 94.950 27.600 97.050 28.050 ;
        RECT 64.950 26.400 97.050 27.600 ;
        RECT 64.950 25.950 67.050 26.400 ;
        RECT 70.950 25.950 73.050 26.400 ;
        RECT 79.950 25.950 82.050 26.400 ;
        RECT 94.950 25.950 97.050 26.400 ;
        RECT 112.950 25.950 115.050 28.050 ;
        RECT 115.950 25.950 118.050 28.050 ;
        RECT 118.950 27.600 121.050 28.050 ;
        RECT 145.950 27.600 148.050 28.050 ;
        RECT 118.950 26.400 148.050 27.600 ;
        RECT 118.950 25.950 121.050 26.400 ;
        RECT 145.950 25.950 148.050 26.400 ;
        RECT 214.950 27.600 217.050 28.050 ;
        RECT 223.950 27.600 226.050 28.050 ;
        RECT 214.950 26.400 226.050 27.600 ;
        RECT 214.950 25.950 217.050 26.400 ;
        RECT 223.950 25.950 226.050 26.400 ;
        RECT 226.950 27.600 229.050 28.050 ;
        RECT 250.950 27.600 253.050 28.050 ;
        RECT 226.950 26.400 253.050 27.600 ;
        RECT 226.950 25.950 229.050 26.400 ;
        RECT 250.950 25.950 253.050 26.400 ;
        RECT 253.950 27.600 256.050 28.050 ;
        RECT 259.950 27.600 262.050 28.050 ;
        RECT 253.950 26.400 262.050 27.600 ;
        RECT 253.950 25.950 256.050 26.400 ;
        RECT 259.950 25.950 262.050 26.400 ;
        RECT 292.950 27.600 295.050 28.050 ;
        RECT 307.950 27.600 310.050 28.050 ;
        RECT 292.950 26.400 310.050 27.600 ;
        RECT 292.950 25.950 295.050 26.400 ;
        RECT 307.950 25.950 310.050 26.400 ;
        RECT 310.950 27.600 313.050 28.050 ;
        RECT 352.950 27.600 355.050 28.050 ;
        RECT 310.950 26.400 355.050 27.600 ;
        RECT 310.950 25.950 313.050 26.400 ;
        RECT 352.950 25.950 355.050 26.400 ;
        RECT 388.950 27.600 391.050 28.050 ;
        RECT 427.950 27.600 430.050 28.050 ;
        RECT 388.950 26.400 430.050 27.600 ;
        RECT 388.950 25.950 391.050 26.400 ;
        RECT 427.950 25.950 430.050 26.400 ;
        RECT 454.950 27.600 457.050 28.050 ;
        RECT 508.950 27.600 511.050 28.050 ;
        RECT 553.950 27.600 556.050 28.050 ;
        RECT 454.950 26.400 556.050 27.600 ;
        RECT 454.950 25.950 457.050 26.400 ;
        RECT 508.950 25.950 511.050 26.400 ;
        RECT 553.950 25.950 556.050 26.400 ;
        RECT 568.950 27.600 571.050 28.050 ;
        RECT 574.950 27.600 577.050 28.050 ;
        RECT 598.950 27.600 601.050 28.050 ;
        RECT 568.950 26.400 601.050 27.600 ;
        RECT 568.950 25.950 571.050 26.400 ;
        RECT 574.950 25.950 577.050 26.400 ;
        RECT 598.950 25.950 601.050 26.400 ;
        RECT 601.950 27.600 604.050 28.050 ;
        RECT 625.950 27.600 628.050 28.050 ;
        RECT 601.950 26.400 628.050 27.600 ;
        RECT 601.950 25.950 604.050 26.400 ;
        RECT 625.950 25.950 628.050 26.400 ;
        RECT 628.950 27.600 631.050 28.050 ;
        RECT 649.950 27.600 652.050 28.050 ;
        RECT 628.950 26.400 652.050 27.600 ;
        RECT 628.950 25.950 631.050 26.400 ;
        RECT 649.950 25.950 652.050 26.400 ;
        RECT 661.950 27.600 664.050 28.050 ;
        RECT 667.950 27.600 670.050 28.050 ;
        RECT 673.950 27.600 676.050 28.050 ;
        RECT 661.950 26.400 676.050 27.600 ;
        RECT 661.950 25.950 664.050 26.400 ;
        RECT 667.950 25.950 670.050 26.400 ;
        RECT 673.950 25.950 676.050 26.400 ;
        RECT 676.950 27.600 679.050 28.050 ;
        RECT 691.950 27.600 694.050 28.050 ;
        RECT 676.950 26.400 694.050 27.600 ;
        RECT 676.950 25.950 679.050 26.400 ;
        RECT 691.950 25.950 694.050 26.400 ;
        RECT 13.950 24.600 16.050 25.050 ;
        RECT 25.950 24.600 28.050 25.050 ;
        RECT 43.950 24.600 46.050 25.050 ;
        RECT 46.950 24.600 49.050 25.050 ;
        RECT 13.950 23.400 24.600 24.600 ;
        RECT 13.950 22.950 16.050 23.400 ;
        RECT 23.400 22.050 24.600 23.400 ;
        RECT 25.950 23.400 49.050 24.600 ;
        RECT 25.950 22.950 28.050 23.400 ;
        RECT 43.950 22.950 46.050 23.400 ;
        RECT 46.950 22.950 49.050 23.400 ;
        RECT 50.400 22.050 51.600 25.950 ;
        RECT 55.950 24.600 58.050 25.050 ;
        RECT 73.950 24.600 76.050 25.050 ;
        RECT 88.950 24.600 91.050 25.050 ;
        RECT 109.950 24.600 112.050 25.050 ;
        RECT 55.950 23.400 91.050 24.600 ;
        RECT 55.950 22.950 58.050 23.400 ;
        RECT 73.950 22.950 76.050 23.400 ;
        RECT 88.950 22.950 91.050 23.400 ;
        RECT 92.400 23.400 112.050 24.600 ;
        RECT 10.950 21.600 13.050 22.050 ;
        RECT 16.950 21.600 19.050 22.050 ;
        RECT 10.950 20.400 19.050 21.600 ;
        RECT 10.950 19.950 13.050 20.400 ;
        RECT 16.950 19.950 19.050 20.400 ;
        RECT 22.950 19.950 25.050 22.050 ;
        RECT 40.950 21.600 43.050 22.050 ;
        RECT 49.950 21.600 52.050 22.050 ;
        RECT 40.950 20.400 52.050 21.600 ;
        RECT 40.950 19.950 43.050 20.400 ;
        RECT 49.950 19.950 52.050 20.400 ;
        RECT 67.950 21.600 70.050 22.050 ;
        RECT 76.950 21.600 79.050 22.050 ;
        RECT 67.950 20.400 79.050 21.600 ;
        RECT 67.950 19.950 70.050 20.400 ;
        RECT 76.950 19.950 79.050 20.400 ;
        RECT 82.950 21.600 85.050 22.050 ;
        RECT 92.400 21.600 93.600 23.400 ;
        RECT 109.950 22.950 112.050 23.400 ;
        RECT 113.400 22.050 114.600 25.950 ;
        RECT 116.400 24.600 117.600 25.950 ;
        RECT 130.950 24.600 133.050 25.050 ;
        RECT 136.950 24.600 139.050 25.050 ;
        RECT 163.950 24.600 166.050 25.050 ;
        RECT 199.950 24.600 202.050 25.050 ;
        RECT 116.400 23.400 129.600 24.600 ;
        RECT 82.950 20.400 93.600 21.600 ;
        RECT 82.950 19.950 85.050 20.400 ;
        RECT 112.950 19.950 115.050 22.050 ;
        RECT 118.950 21.600 121.050 22.050 ;
        RECT 124.950 21.600 127.050 22.050 ;
        RECT 118.950 20.400 127.050 21.600 ;
        RECT 128.400 21.600 129.600 23.400 ;
        RECT 130.950 23.400 139.050 24.600 ;
        RECT 130.950 22.950 133.050 23.400 ;
        RECT 136.950 22.950 139.050 23.400 ;
        RECT 140.400 23.400 202.050 24.600 ;
        RECT 140.400 22.050 141.600 23.400 ;
        RECT 163.950 22.950 166.050 23.400 ;
        RECT 199.950 22.950 202.050 23.400 ;
        RECT 214.950 24.600 217.050 25.050 ;
        RECT 232.950 24.600 235.050 25.050 ;
        RECT 262.950 24.600 265.050 25.050 ;
        RECT 214.950 23.400 235.050 24.600 ;
        RECT 214.950 22.950 217.050 23.400 ;
        RECT 232.950 22.950 235.050 23.400 ;
        RECT 239.400 23.400 265.050 24.600 ;
        RECT 128.400 20.400 135.600 21.600 ;
        RECT 118.950 19.950 121.050 20.400 ;
        RECT 124.950 19.950 127.050 20.400 ;
        RECT 4.950 18.600 7.050 19.050 ;
        RECT 77.400 18.600 78.600 19.950 ;
        RECT 4.950 17.400 78.600 18.600 ;
        RECT 4.950 16.950 7.050 17.400 ;
        RECT 77.400 15.600 78.600 17.400 ;
        RECT 88.950 18.600 91.050 19.050 ;
        RECT 97.950 18.600 100.050 19.050 ;
        RECT 130.950 18.600 133.050 19.050 ;
        RECT 88.950 17.400 133.050 18.600 ;
        RECT 134.400 18.600 135.600 20.400 ;
        RECT 139.950 19.950 142.050 22.050 ;
        RECT 145.950 21.600 148.050 22.050 ;
        RECT 157.950 21.600 160.050 22.050 ;
        RECT 166.950 21.600 169.050 22.050 ;
        RECT 178.950 21.600 181.050 22.050 ;
        RECT 184.950 21.600 187.050 22.050 ;
        RECT 214.950 21.600 217.050 22.050 ;
        RECT 145.950 20.400 169.050 21.600 ;
        RECT 145.950 19.950 148.050 20.400 ;
        RECT 157.950 19.950 160.050 20.400 ;
        RECT 166.950 19.950 169.050 20.400 ;
        RECT 173.400 20.400 187.050 21.600 ;
        RECT 148.950 18.600 151.050 19.050 ;
        RECT 173.400 18.600 174.600 20.400 ;
        RECT 178.950 19.950 181.050 20.400 ;
        RECT 184.950 19.950 187.050 20.400 ;
        RECT 200.400 20.400 217.050 21.600 ;
        RECT 187.950 18.600 190.050 19.050 ;
        RECT 134.400 17.400 174.600 18.600 ;
        RECT 185.400 17.400 190.050 18.600 ;
        RECT 88.950 16.950 91.050 17.400 ;
        RECT 97.950 16.950 100.050 17.400 ;
        RECT 130.950 16.950 133.050 17.400 ;
        RECT 148.950 16.950 151.050 17.400 ;
        RECT 91.950 15.600 94.050 16.050 ;
        RECT 77.400 14.400 94.050 15.600 ;
        RECT 91.950 13.950 94.050 14.400 ;
        RECT 124.950 15.600 127.050 16.050 ;
        RECT 185.400 15.600 186.600 17.400 ;
        RECT 187.950 16.950 190.050 17.400 ;
        RECT 193.950 18.600 196.050 19.050 ;
        RECT 200.400 18.600 201.600 20.400 ;
        RECT 214.950 19.950 217.050 20.400 ;
        RECT 220.950 21.600 223.050 22.050 ;
        RECT 229.950 21.600 232.050 22.050 ;
        RECT 220.950 20.400 232.050 21.600 ;
        RECT 220.950 19.950 223.050 20.400 ;
        RECT 229.950 19.950 232.050 20.400 ;
        RECT 235.950 19.950 238.050 22.050 ;
        RECT 193.950 17.400 201.600 18.600 ;
        RECT 193.950 16.950 196.050 17.400 ;
        RECT 202.950 16.950 205.050 19.050 ;
        RECT 226.950 18.600 229.050 19.050 ;
        RECT 236.400 18.600 237.600 19.950 ;
        RECT 239.400 19.050 240.600 23.400 ;
        RECT 262.950 22.950 265.050 23.400 ;
        RECT 301.950 24.600 304.050 25.050 ;
        RECT 331.950 24.600 334.050 25.050 ;
        RECT 301.950 23.400 334.050 24.600 ;
        RECT 301.950 22.950 304.050 23.400 ;
        RECT 331.950 22.950 334.050 23.400 ;
        RECT 346.950 24.600 349.050 25.050 ;
        RECT 388.950 24.600 391.050 25.050 ;
        RECT 346.950 23.400 391.050 24.600 ;
        RECT 346.950 22.950 349.050 23.400 ;
        RECT 362.400 22.050 363.600 23.400 ;
        RECT 388.950 22.950 391.050 23.400 ;
        RECT 415.950 24.600 418.050 25.050 ;
        RECT 460.950 24.600 463.050 25.050 ;
        RECT 466.950 24.600 469.050 25.050 ;
        RECT 415.950 23.400 423.600 24.600 ;
        RECT 415.950 22.950 418.050 23.400 ;
        RECT 241.950 21.600 244.050 22.050 ;
        RECT 250.950 21.600 253.050 22.050 ;
        RECT 241.950 20.400 253.050 21.600 ;
        RECT 241.950 19.950 244.050 20.400 ;
        RECT 250.950 19.950 253.050 20.400 ;
        RECT 253.950 21.600 256.050 22.050 ;
        RECT 259.950 21.600 262.050 22.050 ;
        RECT 325.950 21.600 328.050 22.050 ;
        RECT 253.950 20.400 262.050 21.600 ;
        RECT 253.950 19.950 256.050 20.400 ;
        RECT 259.950 19.950 262.050 20.400 ;
        RECT 290.400 20.400 328.050 21.600 ;
        RECT 226.950 17.400 237.600 18.600 ;
        RECT 226.950 16.950 229.050 17.400 ;
        RECT 238.950 16.950 241.050 19.050 ;
        RECT 244.950 18.600 247.050 19.050 ;
        RECT 256.950 18.600 259.050 19.050 ;
        RECT 262.950 18.600 265.050 19.050 ;
        RECT 244.950 17.400 265.050 18.600 ;
        RECT 244.950 16.950 247.050 17.400 ;
        RECT 256.950 16.950 259.050 17.400 ;
        RECT 262.950 16.950 265.050 17.400 ;
        RECT 286.950 18.600 289.050 19.050 ;
        RECT 290.400 18.600 291.600 20.400 ;
        RECT 325.950 19.950 328.050 20.400 ;
        RECT 328.950 21.600 331.050 22.050 ;
        RECT 349.950 21.600 352.050 22.050 ;
        RECT 328.950 20.400 352.050 21.600 ;
        RECT 328.950 19.950 331.050 20.400 ;
        RECT 349.950 19.950 352.050 20.400 ;
        RECT 361.950 19.950 364.050 22.050 ;
        RECT 385.950 21.600 388.050 22.050 ;
        RECT 406.950 21.600 409.050 22.050 ;
        RECT 412.950 21.600 415.050 22.050 ;
        RECT 385.950 20.400 415.050 21.600 ;
        RECT 385.950 19.950 388.050 20.400 ;
        RECT 406.950 19.950 409.050 20.400 ;
        RECT 412.950 19.950 415.050 20.400 ;
        RECT 418.950 19.950 421.050 22.050 ;
        RECT 422.400 21.600 423.600 23.400 ;
        RECT 460.950 23.400 469.050 24.600 ;
        RECT 460.950 22.950 463.050 23.400 ;
        RECT 466.950 22.950 469.050 23.400 ;
        RECT 490.950 24.600 493.050 25.050 ;
        RECT 520.950 24.600 523.050 25.050 ;
        RECT 529.950 24.600 532.050 25.050 ;
        RECT 490.950 23.400 532.050 24.600 ;
        RECT 490.950 22.950 493.050 23.400 ;
        RECT 520.950 22.950 523.050 23.400 ;
        RECT 529.950 22.950 532.050 23.400 ;
        RECT 535.950 24.600 538.050 25.050 ;
        RECT 541.950 24.600 544.050 25.050 ;
        RECT 535.950 23.400 544.050 24.600 ;
        RECT 535.950 22.950 538.050 23.400 ;
        RECT 541.950 22.950 544.050 23.400 ;
        RECT 571.950 24.600 574.050 25.050 ;
        RECT 580.950 24.600 583.050 25.050 ;
        RECT 583.950 24.600 586.050 25.050 ;
        RECT 598.950 24.600 601.050 25.050 ;
        RECT 610.950 24.600 613.050 25.050 ;
        RECT 571.950 23.400 601.050 24.600 ;
        RECT 571.950 22.950 574.050 23.400 ;
        RECT 580.950 22.950 583.050 23.400 ;
        RECT 583.950 22.950 586.050 23.400 ;
        RECT 598.950 22.950 601.050 23.400 ;
        RECT 602.400 23.400 613.050 24.600 ;
        RECT 430.950 21.600 433.050 22.050 ;
        RECT 422.400 20.400 433.050 21.600 ;
        RECT 430.950 19.950 433.050 20.400 ;
        RECT 469.950 21.600 472.050 22.050 ;
        RECT 484.950 21.600 487.050 22.050 ;
        RECT 469.950 20.400 487.050 21.600 ;
        RECT 469.950 19.950 472.050 20.400 ;
        RECT 484.950 19.950 487.050 20.400 ;
        RECT 568.950 21.600 571.050 22.050 ;
        RECT 602.400 21.600 603.600 23.400 ;
        RECT 610.950 22.950 613.050 23.400 ;
        RECT 631.950 22.950 634.050 25.050 ;
        RECT 670.950 24.600 673.050 25.050 ;
        RECT 679.950 24.600 682.050 25.050 ;
        RECT 670.950 23.400 682.050 24.600 ;
        RECT 670.950 22.950 673.050 23.400 ;
        RECT 679.950 22.950 682.050 23.400 ;
        RECT 568.950 20.400 603.600 21.600 ;
        RECT 607.950 21.600 610.050 22.050 ;
        RECT 632.400 21.600 633.600 22.950 ;
        RECT 637.950 21.600 640.050 22.050 ;
        RECT 607.950 20.400 640.050 21.600 ;
        RECT 568.950 19.950 571.050 20.400 ;
        RECT 607.950 19.950 610.050 20.400 ;
        RECT 637.950 19.950 640.050 20.400 ;
        RECT 643.950 21.600 646.050 22.050 ;
        RECT 664.950 21.600 667.050 22.050 ;
        RECT 643.950 20.400 667.050 21.600 ;
        RECT 643.950 19.950 646.050 20.400 ;
        RECT 664.950 19.950 667.050 20.400 ;
        RECT 685.950 21.600 688.050 22.050 ;
        RECT 697.950 21.600 700.050 22.050 ;
        RECT 712.950 21.600 715.050 22.050 ;
        RECT 685.950 20.400 696.600 21.600 ;
        RECT 685.950 19.950 688.050 20.400 ;
        RECT 286.950 17.400 291.600 18.600 ;
        RECT 337.950 18.600 340.050 19.050 ;
        RECT 379.950 18.600 382.050 19.050 ;
        RECT 391.950 18.600 394.050 19.050 ;
        RECT 337.950 17.400 394.050 18.600 ;
        RECT 286.950 16.950 289.050 17.400 ;
        RECT 337.950 16.950 340.050 17.400 ;
        RECT 379.950 16.950 382.050 17.400 ;
        RECT 391.950 16.950 394.050 17.400 ;
        RECT 203.400 15.600 204.600 16.950 ;
        RECT 124.950 14.400 204.600 15.600 ;
        RECT 208.950 15.600 211.050 16.050 ;
        RECT 253.950 15.600 256.050 16.050 ;
        RECT 208.950 14.400 256.050 15.600 ;
        RECT 124.950 13.950 127.050 14.400 ;
        RECT 208.950 13.950 211.050 14.400 ;
        RECT 253.950 13.950 256.050 14.400 ;
        RECT 268.950 15.600 271.050 16.050 ;
        RECT 298.950 15.600 301.050 16.050 ;
        RECT 268.950 14.400 301.050 15.600 ;
        RECT 268.950 13.950 271.050 14.400 ;
        RECT 298.950 13.950 301.050 14.400 ;
        RECT 334.950 15.600 337.050 16.050 ;
        RECT 370.950 15.600 373.050 16.050 ;
        RECT 419.400 15.600 420.600 19.950 ;
        RECT 586.950 18.600 589.050 19.050 ;
        RECT 595.950 18.600 598.050 19.050 ;
        RECT 586.950 17.400 598.050 18.600 ;
        RECT 695.400 18.600 696.600 20.400 ;
        RECT 697.950 20.400 715.050 21.600 ;
        RECT 697.950 19.950 700.050 20.400 ;
        RECT 712.950 19.950 715.050 20.400 ;
        RECT 703.950 18.600 706.050 19.050 ;
        RECT 695.400 17.400 706.050 18.600 ;
        RECT 586.950 16.950 589.050 17.400 ;
        RECT 595.950 16.950 598.050 17.400 ;
        RECT 703.950 16.950 706.050 17.400 ;
        RECT 334.950 14.400 420.600 15.600 ;
        RECT 664.950 15.600 667.050 16.050 ;
        RECT 709.950 15.600 712.050 16.050 ;
        RECT 664.950 14.400 712.050 15.600 ;
        RECT 334.950 13.950 337.050 14.400 ;
        RECT 370.950 13.950 373.050 14.400 ;
        RECT 664.950 13.950 667.050 14.400 ;
        RECT 709.950 13.950 712.050 14.400 ;
        RECT 274.950 12.600 277.050 13.050 ;
        RECT 286.950 12.600 289.050 13.050 ;
        RECT 274.950 11.400 289.050 12.600 ;
        RECT 274.950 10.950 277.050 11.400 ;
        RECT 286.950 10.950 289.050 11.400 ;
        RECT 307.950 12.600 310.050 13.050 ;
        RECT 343.950 12.600 346.050 13.050 ;
        RECT 307.950 11.400 346.050 12.600 ;
        RECT 307.950 10.950 310.050 11.400 ;
        RECT 343.950 10.950 346.050 11.400 ;
        RECT 409.950 12.600 412.050 13.050 ;
        RECT 421.950 12.600 424.050 13.050 ;
        RECT 409.950 11.400 424.050 12.600 ;
        RECT 409.950 10.950 412.050 11.400 ;
        RECT 421.950 10.950 424.050 11.400 ;
        RECT 181.950 9.600 184.050 10.050 ;
        RECT 226.950 9.600 229.050 10.050 ;
        RECT 181.950 8.400 229.050 9.600 ;
        RECT 181.950 7.950 184.050 8.400 ;
        RECT 226.950 7.950 229.050 8.400 ;
  END
END fir_pe
END LIBRARY

