magic
tech scmos
magscale 1 2
timestamp 1727424219
<< nwell >>
rect -12 152 92 272
<< ntransistor >>
rect 20 14 24 34
rect 40 14 44 34
<< ptransistor >>
rect 20 166 24 246
rect 28 166 32 246
<< ndiffusion >>
rect 18 14 20 34
rect 24 14 26 34
rect 38 14 40 34
rect 44 14 46 34
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 28 246
rect 32 166 34 246
<< ndcontact >>
rect 6 14 18 34
rect 26 14 38 34
rect 46 14 58 34
<< pdcontact >>
rect 6 166 18 246
rect 34 166 46 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 20 246 24 250
rect 28 246 32 250
rect 20 149 24 166
rect 16 137 24 149
rect 20 34 24 137
rect 28 129 32 166
rect 28 117 44 129
rect 40 34 44 117
rect 20 10 24 14
rect 40 10 44 14
<< polycontact >>
rect 4 137 16 149
rect 44 117 56 129
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 6 246 18 252
rect 28 159 46 166
rect 3 123 17 137
rect 28 77 37 159
rect 43 103 57 117
rect 23 63 37 77
rect 26 34 34 63
rect 6 8 18 14
rect 46 8 58 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m1p >>
rect 3 123 17 137
rect 43 103 57 117
rect 23 63 37 77
<< labels >>
rlabel metal1 -6 252 86 268 0 vdd
port 3 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 3 123 17 137 0 A
port 0 nsew signal input
rlabel metal1 23 63 37 77 0 Y
port 2 nsew signal output
rlabel metal1 43 103 57 117 0 B
port 1 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
