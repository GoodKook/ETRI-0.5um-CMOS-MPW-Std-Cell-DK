magic
tech scmos
magscale 1 3
timestamp 1723012252
<< checkpaint >>
rect -56 -56 84 404
<< diffusion >>
rect 5 5 23 343
<< metal1 >>
rect 4 4 24 344
<< end >>
