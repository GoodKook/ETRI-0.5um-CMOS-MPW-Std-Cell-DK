magic
tech scmos
magscale 1 30
timestamp 1741148472
<< checkpaint >>
rect -1190 25645 3530 26220
rect -1190 -615 3786 25645
rect -1190 -1380 3530 -615
<< metal3 >>
rect 30 23400 1770 25060
rect 30 21100 1770 22760
rect 30 11290 1770 19100
rect 30 0 1770 7800
use IOFILLER10  IOFILLER10_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 400 0 1 0
box -35 0 1035 25060
<< end >>
