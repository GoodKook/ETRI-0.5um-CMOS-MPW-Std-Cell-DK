magic
tech scmos
magscale 1 2
timestamp 1701001990
<< checkpaint >>
rect -52 612 192 912
rect -53 312 275 612
rect 328 608 1232 912
rect 1368 608 1712 912
rect 328 552 1712 608
rect 1101 512 1397 552
rect -53 252 593 312
rect 1094 252 1393 348
rect 132 -48 593 252
<< error_s >>
rect 0 854 1592 866
rect 0 594 1600 606
rect 0 554 1246 566
rect 0 294 1246 306
rect 0 254 1344 266
rect 0 0 1344 6
rect 0 -6 784 0
rect 946 -6 1344 0
<< metal1 >>
rect -97 868 -37 953
rect -97 852 24 868
rect -97 568 -37 852
rect 1781 608 1841 943
rect 1466 592 1841 608
rect -97 552 21 568
rect 1141 552 1753 568
rect -97 268 -37 552
rect 1781 308 1841 592
rect 1134 292 1841 308
rect -97 252 28 268
rect -97 -47 -37 252
rect 1781 8 1841 292
rect 1292 -8 1841 8
rect 1781 -57 1841 -8
use AND2X1  AND2X1_0
timestamp 1700698000
transform 1 0 0 0 1 0
box -13 -8 94 272
use AND2X2  AND2X2_0
timestamp 1700698000
transform 1 0 92 0 1 0
box -12 -8 94 272
use AOI21X1  AOI21X1_0
timestamp 1700712373
transform 1 0 184 0 1 0
box -12 -8 92 272
use AOI22X1  AOI22X1_0
timestamp 1700712373
transform 1 0 276 0 1 0
box -14 -8 114 272
use BUFX2  BUFX2_0
timestamp 1700717866
transform 1 0 388 0 1 0
box -12 -8 72 272
use BUFX4  BUFX4_0
timestamp 1700717866
transform 1 0 460 0 1 0
box -13 -8 93 272
use CLKBUF1  CLKBUF1_0
timestamp 1700699651
transform 1 0 552 0 1 0
box -12 -8 192 272
use CLKBUF2  CLKBUF2_0
timestamp 1700698000
transform 1 0 738 0 1 0
box -12 -8 273 272
use CLKBUF3  CLKBUF3_0
timestamp 1700698000
transform 1 0 998 0 1 0
box -12 -8 353 272
use DFFNEGX1  DFFNEGX1_0
timestamp 1700717866
transform 1 0 0 0 1 300
box -13 -8 235 272
use DFFPOSX1  DFFPOSX1_0
timestamp 1700699651
transform 1 0 220 0 1 300
box -13 -8 253 272
use DFFSR  DFFSR_0
timestamp 1700698000
transform 1 0 460 0 1 300
box -12 -8 474 272
use FAX1  FAX1_0
timestamp 1700698000
transform 1 0 920 0 1 300
box -13 -8 313 272
use FILL  FILL_0
timestamp 1700315010
transform 1 0 1220 0 1 300
box -12 -8 32 272
use HAX1  HAX1_0
timestamp 1700698000
transform 1 0 1540 0 1 300
box -13 -8 213 272
use INVX1  INVX1_0
timestamp 1700712373
transform 1 0 0 0 1 600
box -12 -8 52 272
use INVX2  INVX2_0
timestamp 1700698000
transform 1 0 40 0 1 600
box -12 -8 52 272
use INVX4  INVX4_0
timestamp 1700715846
transform 1 0 80 0 1 600
box -12 -8 72 272
use INVX8  INVX8_0
timestamp 1700698000
transform 1 0 140 0 1 600
box -12 -8 114 272
use LATCH  LATCH_0
timestamp 1700698000
transform 1 0 240 0 1 600
box -12 -8 153 272
use MUX2X1  MUX2X1_0
timestamp 1700700889
transform 1 0 380 0 1 600
box -12 -8 114 272
use NAND2X1  NAND2X1_0
timestamp 1700712373
transform 1 0 480 0 1 600
box -12 -8 72 272
use NAND3X1  NAND3X1_0
timestamp 1700712373
transform 1 0 540 0 1 600
box -12 -8 92 272
use NOR2X1  NOR2X1_0
timestamp 1700712373
transform 1 0 620 0 1 600
box -12 -8 74 272
use NOR3X1  NOR3X1_0
timestamp 1700720714
transform 1 0 680 0 1 600
box -12 -8 172 272
use OAI21X1  OAI21X1_0
timestamp 1700726220
transform 1 0 840 0 1 600
box -12 -8 92 272
use OAI22X1  OAI22X1_0
timestamp 1700700889
transform 1 0 920 0 1 600
box -12 -8 112 272
use OR2X1  OR2X1_0
timestamp 1700717866
transform 1 0 1020 0 1 600
box -13 -8 93 272
use OR2X2  OR2X2_0
timestamp 1700708354
transform 1 0 1100 0 1 600
box -12 -8 92 272
use TBUFX1  TBUFX1_0
timestamp 1700498524
transform 1 0 1180 0 1 600
box -14 -8 113 272
use TBUFX2  TBUFX2_0
timestamp 1700347708
transform 1 0 1280 0 1 600
box -13 -8 153 272
use XNOR2X1  XNOR2X1_0
timestamp 1700717866
transform 1 0 1420 0 1 600
box -12 -8 132 272
use XOR2X1  XOR2X1_0
timestamp 1700717866
transform 1 0 1540 0 1 600
box -12 -8 132 272
<< labels >>
rlabel metal1 -73 921 -73 921 0 vdd
port 1 nsew power bidirectional abutment
rlabel metal1 1808 905 1808 905 0 gnd
port 2 nsew ground bidirectional abutment
<< end >>
