magic
tech scmos
magscale 1 3
timestamp 1555596690
<< checkpaint >>
rect -60 -60 330 330
<< nwell >>
rect 0 0 270 270
<< nsubstratendiff >>
rect 20 230 250 250
rect 20 40 40 230
rect 230 40 250 230
rect 20 20 250 40
<< metal1 >>
rect 20 230 250 250
rect 20 40 40 230
rect 230 40 250 230
rect 20 20 250 40
use ntap_CDNS_723012252911  ntap_CDNS_723012252911_0
timestamp 1555596690
transform 1 0 226 0 1 36
box 4 4 24 194
use ntap_CDNS_723012252911  ntap_CDNS_723012252911_1
timestamp 1555596690
transform 1 0 16 0 1 36
box 4 4 24 194
use ntap_CDNS_7230122529129  ntap_CDNS_7230122529129_0
timestamp 1555596690
transform 1 0 36 0 1 226
box 4 4 194 24
use ntap_CDNS_7230122529129  ntap_CDNS_7230122529129_1
timestamp 1555596690
transform 1 0 36 0 1 16
box 4 4 194 24
<< end >>
