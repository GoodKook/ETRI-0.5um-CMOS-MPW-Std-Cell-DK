magic
tech scmos
timestamp 1569139307
<< checkpaint >>
rect -21 -21 21 21
<< genericcontact >>
rect -1 -1 1 1
<< end >>
