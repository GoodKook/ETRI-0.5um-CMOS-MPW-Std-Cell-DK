magic
tech scmos
timestamp 1721969656
<< error_p >>
rect 33 126 33 132
<< nwell >>
rect -8 124 36 135
rect -8 96 36 124
<< ntransistor >>
rect 8 6 10 16
rect 18 6 20 16
<< ptransistor >>
rect 8 112 10 122
rect 18 112 20 122
<< ndiffusion >>
rect 7 6 8 16
rect 10 6 11 16
rect 17 6 18 16
rect 20 6 21 16
<< pdiffusion >>
rect 7 112 8 122
rect 10 112 11 122
rect 17 112 18 122
rect 20 112 21 122
<< ndcontact >>
rect 1 6 7 16
rect 11 6 17 16
rect 21 6 27 16
<< pdcontact >>
rect 1 112 7 122
rect 11 112 17 122
rect 21 112 27 122
<< psubstratepcontact >>
rect -5 -4 33 2
<< nsubstratencontact >>
rect -5 126 33 132
<< polysilicon >>
rect 8 122 10 124
rect 18 122 20 124
rect 8 39 10 112
rect 18 49 20 112
rect 8 37 20 39
rect 8 16 10 27
rect 18 16 20 37
rect 8 4 10 6
rect 18 4 20 6
<< polycontact >>
rect 14 43 20 49
rect 8 27 14 33
<< metal1 >>
rect -5 132 33 133
rect -5 125 33 126
rect 2 67 5 112
rect 13 60 16 112
rect 23 66 26 112
rect 13 43 14 49
rect 13 33 16 43
rect 14 27 16 33
rect -5 2 33 3
rect -5 -5 33 -4
<< m2contact >>
rect -2 60 5 67
rect 10 53 17 60
rect 23 59 30 66
rect 0 16 7 24
rect 10 16 17 24
rect 20 16 27 24
<< metal2 >>
rect 2 24 5 60
rect 13 24 16 53
rect 23 24 26 59
<< end >>
