magic
tech scmos
magscale 1 30
timestamp 1756369954
<< checkpaint >>
rect 9150 9150 180850 180850
<< metal1 >>
rect 144100 163300 148200 171100
rect 145550 147700 148200 163300
rect 143950 146000 169800 147700
rect 142700 145100 169800 146000
rect 140200 143600 169800 145100
rect 46700 141950 47900 142000
rect 46450 49950 47900 141950
rect 46450 46300 47940 49950
rect 166800 43900 169800 143600
rect 143300 42300 169800 43900
rect 146800 40100 169800 42300
rect 146800 26700 149700 40100
rect 143900 18900 149700 26700
<< m2contact >>
rect 142800 163300 144100 171100
rect 142700 146000 143950 147700
rect 130800 143600 140200 145100
rect 46450 45100 57900 46300
rect 142300 42300 143300 43900
rect 142700 18900 143900 26700
<< metal2 >>
rect 59800 145100 60200 145900
rect 48200 142230 48500 144800
rect 73300 144600 73700 145900
rect 44100 140600 45600 141000
rect 48210 140047 48315 142230
rect 50500 142200 50800 144300
rect 86800 144100 87200 145900
rect 52000 142200 52300 143800
rect 100300 143600 100700 145900
rect 53200 142230 53500 143300
rect 113800 143100 114200 145900
rect 54700 142250 55000 142800
rect 127300 142600 127700 145900
rect 130800 145100 140200 145800
rect 56010 142048 56115 142300
rect 44100 116300 46500 116700
rect 44100 102800 45700 103200
rect 45400 94600 45700 102800
rect 45400 89700 45700 92600
rect 44100 89300 45700 89700
rect 44100 75800 45900 76200
rect 44100 73100 46400 73500
rect 44100 59600 45800 60000
rect 45500 47300 45800 59600
rect 46100 47900 46400 73100
rect 101610 47900 101715 48057
rect 101500 47300 101800 47900
rect 102400 46700 102700 47900
rect 51200 44100 57900 45100
rect 62500 44100 62900 46400
rect 105400 46100 105700 47900
rect 76000 44100 76400 45800
rect 106600 45500 106900 47900
rect 89500 44100 89900 45200
rect 113800 44900 114100 47900
rect 117700 45700 118000 48000
rect 123200 46400 123500 47900
rect 123200 46100 130400 46400
rect 116500 45300 118000 45700
rect 103000 44100 103400 44600
rect 116500 44100 116900 45300
rect 130000 44100 130400 46100
<< m3contact >>
rect 141500 163300 142800 171100
rect 141450 146000 142700 147700
rect 48200 144800 48800 145100
rect 59600 144800 60200 145100
rect 50500 144300 51100 144600
rect 73100 144300 73700 144600
rect 45600 139500 45900 141000
rect 52000 143800 52600 144100
rect 86600 143800 87200 144100
rect 53200 143300 53800 143600
rect 100100 143300 100700 143600
rect 54700 142800 55300 143100
rect 113600 142800 114200 143100
rect 56000 142300 56600 142600
rect 127100 142300 127700 142600
rect 46500 116300 46800 117000
rect 45400 94000 45700 94600
rect 45400 92600 45700 93300
rect 45900 75800 46200 76500
rect 46100 47600 46700 47900
rect 99300 47600 100000 47900
rect 45500 47000 46100 47300
rect 101100 47000 101800 47300
rect 62500 46400 63200 46700
rect 102000 46400 102700 46700
rect 76000 45800 76700 46100
rect 105000 45800 105700 46100
rect 89500 45200 90200 45500
rect 106200 45200 106900 45500
rect 103000 44600 103700 44900
rect 113400 44600 114100 44900
rect 141500 42300 142300 43900
rect 141500 18900 142700 26700
<< metal3 >>
rect 48800 144800 59600 145100
rect 51100 144300 73100 144600
rect 52600 143800 86600 144100
rect 53800 143300 100100 143600
rect 55300 142800 113600 143100
rect 56600 142300 127100 142600
rect 45900 139500 47700 139800
rect 46500 129300 47800 129600
rect 46500 117000 46800 129300
rect 45700 94000 47800 94300
rect 45700 93000 47800 93300
rect 45900 85800 47800 86100
rect 45900 76500 46200 85800
rect 46700 47600 99300 47900
rect 46100 47000 101100 47300
rect 63200 46400 102000 46700
rect 76700 45800 105000 46100
rect 90200 45200 106200 45500
rect 103700 44600 113400 44900
use PIC  CLK ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1756352440
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use fir_hls_Core  fir_hls_Core_0
timestamp 1756369697
transform 1 0 47970 0 1 48170
box -930 -360 119730 94140
use PVSS  GND ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 129500 0 -1 171100
box 0 -9150 12000 25300
use IOFILLER18  IOFILLER18_6 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1741148472
transform 1 0 73845 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_7
timestamp 1741148472
transform 1 0 60345 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_8
timestamp 1741148472
transform 1 0 100845 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_9
timestamp 1741148472
transform 1 0 87345 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_10
timestamp 1741148472
transform 1 0 127845 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_11
timestamp 1741148472
transform 1 0 114345 0 1 18900
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_12
timestamp 1741148472
transform 0 1 18899 -1 0 75655
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_13
timestamp 1741148472
transform 0 1 18899 -1 0 62155
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_14
timestamp 1741148472
transform 0 1 18900 -1 0 102655
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_15
timestamp 1741148472
transform 0 1 18900 -1 0 89155
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_16
timestamp 1741148472
transform 1 0 73845 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_17
timestamp 1741148472
transform 0 1 18897 -1 0 116155
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_18
timestamp 1741148472
transform 0 1 18900 -1 0 129655
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_19
timestamp 1741148472
transform 1 0 60345 0 -1 171101
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_20
timestamp 1741148472
transform 1 0 100845 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_21
timestamp 1741148472
transform 1 0 87344 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_22
timestamp 1741148472
transform 1 0 127845 0 -1 171100
box 30 0 1770 25060
use IOFILLER18  IOFILLER18_23
timestamp 1741148472
transform 1 0 114345 0 -1 171100
box 30 0 1770 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use MY_LOGO  MY_LOGO_0
timestamp 1756367991
transform 1 0 -610 0 1 -230
box 152200 14900 178300 173120
use PAD_80__0  PAD_80_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1740657577
transform 0 -1 176000 1 0 135500
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_1
timestamp 1740657577
transform 0 -1 176000 1 0 122000
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_2
timestamp 1740657577
transform 0 -1 176000 1 0 108500
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_3
timestamp 1740657577
transform 0 -1 176000 1 0 95000
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_4
timestamp 1740657577
transform 0 -1 176000 1 0 81500
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_5
timestamp 1740657577
transform 0 -1 176000 1 0 68000
box -4250 -4250 4250 4900
use PAD_80__0  PAD_80_6
timestamp 1740657577
transform 0 -1 176000 1 0 54500
box -4250 -4250 4250 4900
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use POB8  READY ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PIC  RST
timestamp 1756352440
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PVDD  VDD ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 48500 0 1 18900
box 0 -9150 12000 25300
use PIC  X_0
timestamp 1756352440
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_1
timestamp 1756352440
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_2
timestamp 1756352440
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_3
timestamp 1756352440
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  X_4
timestamp 1756352440
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_5
timestamp 1756352440
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  X_6
timestamp 1756352440
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  X_7
timestamp 1756352440
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use POB8  Y_0
timestamp 1569139307
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_1
timestamp 1569139307
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use POB8  Y_2
timestamp 1569139307
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use POB8  Y_3
timestamp 1569139307
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_4
timestamp 1569139307
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_5
timestamp 1569139307
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_6
timestamp 1569139307
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use POB8  Y_7
timestamp 1569139307
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
<< end >>
