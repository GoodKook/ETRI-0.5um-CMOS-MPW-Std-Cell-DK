magic
tech scmos
magscale 1 2
timestamp 1702316108
<< nwell >>
rect -12 154 353 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
rect 78 14 82 54
rect 98 14 102 54
rect 118 14 122 54
rect 138 14 142 54
rect 158 14 162 54
rect 178 14 182 54
rect 198 14 202 54
rect 218 14 222 54
rect 238 14 242 54
rect 258 14 262 54
rect 278 14 282 54
rect 298 14 302 54
rect 318 14 322 54
<< ptransistor >>
rect 18 166 22 246
rect 38 166 42 246
rect 58 166 62 246
rect 78 166 82 246
rect 98 166 102 246
rect 118 166 122 246
rect 138 166 142 246
rect 158 166 162 246
rect 178 166 182 246
rect 198 166 202 246
rect 218 166 222 246
rect 238 166 242 246
rect 258 166 262 246
rect 278 166 282 246
rect 298 166 302 246
rect 318 166 322 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 14 24 54
rect 36 14 38 54
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
rect 76 14 78 54
rect 82 14 84 54
rect 96 14 98 54
rect 102 14 104 54
rect 116 14 118 54
rect 122 14 124 54
rect 136 14 138 54
rect 142 14 144 54
rect 156 14 158 54
rect 162 14 164 54
rect 176 14 178 54
rect 182 14 184 54
rect 196 14 198 54
rect 202 14 204 54
rect 216 14 218 54
rect 222 14 224 54
rect 236 14 238 54
rect 242 14 244 54
rect 256 14 258 54
rect 262 14 264 54
rect 276 14 278 54
rect 282 14 284 54
rect 296 14 298 54
rect 302 14 304 54
rect 316 14 318 54
rect 322 14 324 54
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 24 246
rect 36 166 38 246
rect 42 166 44 246
rect 56 166 58 246
rect 62 166 64 246
rect 76 166 78 246
rect 82 166 84 246
rect 96 166 98 246
rect 102 166 104 246
rect 116 166 118 246
rect 122 166 124 246
rect 136 166 138 246
rect 142 166 144 246
rect 156 166 158 246
rect 162 166 164 246
rect 176 166 178 246
rect 182 166 184 246
rect 196 166 198 246
rect 202 166 204 246
rect 216 166 218 246
rect 222 166 224 246
rect 236 166 238 246
rect 242 166 244 246
rect 256 166 258 246
rect 262 166 264 246
rect 276 166 278 246
rect 282 166 284 246
rect 296 166 298 246
rect 302 166 304 246
rect 316 166 318 246
rect 322 166 324 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 54
rect 44 14 56 54
rect 64 14 76 54
rect 84 14 96 54
rect 104 14 116 54
rect 124 14 136 54
rect 144 14 156 54
rect 164 14 176 54
rect 184 14 196 54
rect 204 14 216 54
rect 224 14 236 54
rect 244 14 256 54
rect 264 14 276 54
rect 284 14 296 54
rect 304 14 316 54
rect 324 14 336 54
<< pdcontact >>
rect 4 166 16 246
rect 24 166 36 246
rect 44 166 56 246
rect 64 166 76 246
rect 84 166 96 246
rect 104 166 116 246
rect 124 166 136 246
rect 144 166 156 246
rect 164 166 176 246
rect 184 166 196 246
rect 204 166 216 246
rect 224 166 236 246
rect 244 166 256 246
rect 264 166 276 246
rect 284 166 296 246
rect 304 166 316 246
rect 324 166 336 246
<< psubstratepcontact >>
rect -6 -6 346 6
<< nsubstratencontact >>
rect -6 254 346 266
<< polysilicon >>
rect 18 246 22 250
rect 38 246 42 250
rect 58 246 62 250
rect 78 246 82 250
rect 98 246 102 250
rect 118 246 122 250
rect 138 246 142 250
rect 158 246 162 250
rect 178 246 182 250
rect 198 246 202 250
rect 218 246 222 250
rect 238 246 242 250
rect 258 246 262 250
rect 278 246 282 250
rect 298 246 302 250
rect 318 246 322 250
rect 18 117 22 166
rect 38 117 42 166
rect 18 108 42 117
rect 18 54 22 108
rect 38 54 42 108
rect 58 120 62 166
rect 78 116 82 166
rect 70 108 82 116
rect 58 54 62 108
rect 78 54 82 108
rect 98 120 102 166
rect 118 116 122 166
rect 110 108 122 116
rect 98 54 102 108
rect 118 54 122 108
rect 138 120 142 166
rect 158 116 162 166
rect 150 108 162 116
rect 138 54 142 108
rect 158 54 162 108
rect 178 120 182 166
rect 198 116 202 166
rect 190 108 202 116
rect 178 54 182 108
rect 198 54 202 108
rect 218 120 222 166
rect 238 116 242 166
rect 230 108 242 116
rect 218 54 222 108
rect 238 54 242 108
rect 258 120 262 166
rect 278 116 282 166
rect 270 108 282 116
rect 258 54 262 108
rect 278 54 282 108
rect 298 107 302 166
rect 318 107 322 166
rect 310 99 322 107
rect 298 54 302 95
rect 318 54 322 99
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
rect 78 10 82 14
rect 98 10 102 14
rect 118 10 122 14
rect 138 10 142 14
rect 158 10 162 14
rect 178 10 182 14
rect 198 10 202 14
rect 218 10 222 14
rect 238 10 242 14
rect 258 10 262 14
rect 278 10 282 14
rect 298 10 302 14
rect 318 10 322 14
<< polycontact >>
rect 6 105 18 117
rect 58 108 70 120
rect 98 108 110 120
rect 138 108 150 120
rect 178 108 190 120
rect 218 108 230 120
rect 258 108 270 120
rect 298 95 310 107
<< metal1 >>
rect -6 266 346 268
rect -6 252 346 254
rect 4 246 16 252
rect 44 246 56 252
rect 84 246 96 252
rect 124 246 136 252
rect 164 246 176 252
rect 204 246 216 252
rect 244 246 256 252
rect 284 246 296 252
rect 324 246 336 252
rect 24 160 36 166
rect 64 160 76 166
rect 104 160 116 166
rect 144 160 156 166
rect 184 160 196 166
rect 224 160 236 166
rect 264 160 276 166
rect 24 152 47 160
rect 64 152 90 160
rect 104 152 130 160
rect 144 152 172 160
rect 184 152 206 160
rect 224 152 250 160
rect 264 152 290 160
rect 3 123 17 137
rect 6 117 17 123
rect 39 116 47 152
rect 39 108 58 116
rect 82 116 90 152
rect 82 108 98 116
rect 122 116 130 152
rect 122 108 138 116
rect 164 116 172 152
rect 164 108 178 116
rect 198 116 206 152
rect 198 108 218 116
rect 242 116 250 152
rect 242 108 258 116
rect 39 68 47 108
rect 82 68 90 108
rect 122 68 130 108
rect 164 68 172 108
rect 198 68 206 108
rect 242 68 250 108
rect 282 107 290 152
rect 306 137 316 166
rect 303 123 326 137
rect 282 99 298 107
rect 282 68 290 99
rect 319 68 326 123
rect 24 60 47 68
rect 64 60 90 68
rect 104 60 130 68
rect 144 60 172 68
rect 184 60 206 68
rect 224 60 250 68
rect 264 60 290 68
rect 304 60 326 68
rect 24 54 36 60
rect 64 54 76 60
rect 104 54 116 60
rect 144 54 156 60
rect 184 54 196 60
rect 224 54 236 60
rect 264 54 276 60
rect 304 54 316 60
rect 4 8 16 14
rect 44 8 56 14
rect 84 8 96 14
rect 124 8 136 14
rect 164 8 176 14
rect 204 8 216 14
rect 244 8 256 14
rect 284 8 296 14
rect 324 8 336 14
rect -6 6 346 8
rect -6 -8 346 -6
<< m1p >>
rect -6 252 346 268
rect 3 123 17 137
rect 303 123 317 137
rect -6 -8 346 8
<< labels >>
rlabel nsubstratencontact 170 260 170 260 0 vdd
port 3 nsew power bidirectional abutment
rlabel psubstratepcontact 170 0 170 0 0 gnd
port 4 nsew ground bidirectional abutment
rlabel metal1 10 131 10 131 0 A
port 1 nsew signal input
rlabel metal1 310 130 310 130 0 Y
port 2 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 340 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
