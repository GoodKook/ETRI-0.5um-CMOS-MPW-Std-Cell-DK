magic
tech scmos
magscale 1 2
timestamp 1702316108
<< nwell >>
rect -12 154 153 272
<< ntransistor >>
rect 22 14 26 54
rect 42 14 46 34
rect 54 14 58 34
rect 82 14 86 34
rect 92 14 96 34
rect 114 14 118 54
<< ptransistor >>
rect 22 166 26 246
rect 44 206 48 246
rect 54 206 58 246
rect 82 226 86 246
rect 92 226 96 246
rect 114 166 118 246
<< ndiffusion >>
rect 20 14 22 54
rect 26 14 28 54
rect 40 14 42 34
rect 46 14 54 34
rect 58 14 64 34
rect 76 14 82 34
rect 86 14 92 34
rect 96 14 100 34
rect 112 14 114 54
rect 118 14 120 54
<< pdiffusion >>
rect 20 166 22 246
rect 26 166 28 246
rect 40 206 44 246
rect 48 206 54 246
rect 58 206 62 246
rect 75 226 82 246
rect 86 226 92 246
rect 96 226 100 246
rect 112 166 114 246
rect 118 166 120 246
<< ndcontact >>
rect 8 14 20 54
rect 28 14 40 54
rect 64 14 76 34
rect 100 14 112 54
rect 120 14 132 54
<< pdcontact >>
rect 8 166 20 246
rect 28 166 40 246
rect 62 206 75 246
rect 100 166 112 246
rect 120 166 132 246
<< psubstratepcontact >>
rect -6 -6 146 6
<< nsubstratencontact >>
rect -6 254 146 266
<< polysilicon >>
rect 22 246 26 250
rect 44 246 48 250
rect 54 246 58 250
rect 82 246 86 250
rect 92 246 96 250
rect 114 246 118 250
rect 22 117 26 166
rect 44 161 48 206
rect 42 154 48 161
rect 22 54 26 105
rect 42 96 46 154
rect 54 148 58 206
rect 82 191 86 226
rect 74 187 86 191
rect 42 34 46 84
rect 60 78 64 136
rect 74 99 78 187
rect 92 99 96 226
rect 114 160 118 166
rect 116 148 118 160
rect 92 87 94 99
rect 60 74 86 78
rect 54 54 57 66
rect 54 34 58 54
rect 82 34 86 74
rect 92 34 96 87
rect 114 54 118 148
rect 22 10 26 14
rect 42 10 46 14
rect 54 10 58 14
rect 82 10 86 14
rect 92 10 96 14
rect 114 10 118 14
<< polycontact >>
rect 21 105 33 117
rect 54 136 66 148
rect 40 84 52 96
rect 104 148 116 160
rect 72 87 84 99
rect 94 87 106 99
rect 57 54 69 66
<< metal1 >>
rect -6 266 146 268
rect -6 252 146 254
rect 28 246 40 252
rect 100 246 112 252
rect 8 160 16 166
rect 8 154 58 160
rect 132 166 134 173
rect 78 154 104 160
rect 8 142 17 154
rect 50 148 58 154
rect 23 123 37 137
rect 50 136 54 148
rect 126 137 134 166
rect 83 127 97 137
rect 23 117 34 123
rect 33 105 34 117
rect 27 66 34 105
rect 45 121 97 127
rect 123 123 137 137
rect 45 96 52 121
rect 126 99 134 123
rect 106 87 134 99
rect 72 66 78 87
rect 27 60 57 66
rect 69 54 78 66
rect 126 54 134 87
rect 62 14 64 34
rect 132 45 134 54
rect 28 8 40 14
rect 100 8 112 14
rect -6 6 146 8
rect -6 -8 146 -6
<< m2contact >>
rect 64 192 78 206
rect 64 154 78 168
rect 3 128 17 142
rect 7 54 21 68
rect 64 34 78 48
<< metal2 >>
rect 64 168 72 192
rect 8 68 16 128
rect 64 48 72 154
<< m1p >>
rect -6 252 146 268
rect 23 123 37 137
rect 83 123 97 137
rect 123 123 137 137
rect -6 -8 146 8
<< labels >>
rlabel nsubstratencontact 70 260 70 260 0 vdd
port 4 nsew power bidirectional abutment
rlabel psubstratepcontact 70 0 70 0 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 30 131 30 131 0 CLK
port 2 nsew clock input
rlabel metal1 90 130 90 130 0 D
port 1 nsew signal input
rlabel metal1 130 133 130 133 0 Q
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 140 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
