magic
tech scmos
magscale 1 6
timestamp 1725338570
<< checkpaint >>
rect -82 334 190 386
rect -108 330 216 334
rect -108 -106 270 330
<< ntransistor >>
rect 49 14 59 214
<< ndiffusion >>
rect 46 14 49 214
rect 59 14 62 214
<< ndcontact >>
rect 12 14 46 214
rect 62 14 96 214
<< psubstratepcontact >>
rect 118 14 150 210
<< polysilicon >>
rect 49 214 59 234
rect 49 4 59 14
<< polycontact >>
rect 38 234 70 266
<< metal1 >>
rect 36 266 72 268
rect 36 234 38 266
rect 70 234 72 266
rect 36 232 72 234
rect 10 214 46 216
rect 10 14 12 214
rect 10 12 46 14
rect 62 214 98 216
rect 96 14 98 214
rect 62 12 98 14
rect 116 210 152 212
rect 116 14 118 210
rect 150 14 152 210
rect 116 12 152 14
<< end >>
