magic
tech scmos
magscale 1 30
timestamp 1709384323
<< nwell >>
rect 0 30150 12195 32010
rect 0 20350 12200 28350
rect 0 17350 12195 18550
<< ntransistor >>
rect 7965 33210 8015 33710
rect 8225 33210 8275 33710
rect 8485 33210 8535 33710
rect 8745 33210 8795 33710
rect 9305 33120 9355 33740
rect 10185 33120 10235 33740
rect 10775 33120 10825 33740
rect 11365 33120 11415 33740
rect 1190 10050 1260 16050
rect 2120 10050 2190 16050
rect 2450 10050 2520 16050
rect 3380 10050 3450 16050
rect 3710 10050 3780 16050
rect 4640 10050 4710 16050
rect 4970 10050 5040 16050
rect 5900 10050 5970 16050
rect 6230 10050 6300 16050
rect 7160 10050 7230 16050
rect 7490 10050 7560 16050
rect 8420 10050 8490 16050
rect 8750 10050 8820 16050
rect 9680 10050 9750 16050
rect 10010 10050 10080 16050
rect 10940 10050 11010 16050
<< ndiffusion >>
rect 7780 33610 7965 33710
rect 7780 33550 7830 33610
rect 7890 33550 7965 33610
rect 7780 33490 7965 33550
rect 7780 33430 7830 33490
rect 7890 33430 7965 33490
rect 7780 33370 7965 33430
rect 7780 33310 7830 33370
rect 7890 33310 7965 33370
rect 7780 33210 7965 33310
rect 8015 33610 8225 33710
rect 8015 33550 8090 33610
rect 8150 33550 8225 33610
rect 8015 33490 8225 33550
rect 8015 33430 8090 33490
rect 8150 33430 8225 33490
rect 8015 33370 8225 33430
rect 8015 33310 8090 33370
rect 8150 33310 8225 33370
rect 8015 33210 8225 33310
rect 8275 33610 8485 33710
rect 8275 33550 8350 33610
rect 8410 33550 8485 33610
rect 8275 33490 8485 33550
rect 8275 33430 8350 33490
rect 8410 33430 8485 33490
rect 8275 33370 8485 33430
rect 8275 33310 8350 33370
rect 8410 33310 8485 33370
rect 8275 33210 8485 33310
rect 8535 33610 8745 33710
rect 8535 33550 8610 33610
rect 8670 33550 8745 33610
rect 8535 33490 8745 33550
rect 8535 33430 8610 33490
rect 8670 33430 8745 33490
rect 8535 33370 8745 33430
rect 8535 33310 8610 33370
rect 8670 33310 8745 33370
rect 8535 33210 8745 33310
rect 8795 33610 8980 33710
rect 8795 33550 8870 33610
rect 8930 33550 8980 33610
rect 8795 33490 8980 33550
rect 8795 33430 8870 33490
rect 8930 33430 8980 33490
rect 8795 33370 8980 33430
rect 8795 33310 8870 33370
rect 8930 33310 8980 33370
rect 8795 33210 8980 33310
rect 9090 33530 9305 33740
rect 9090 33470 9150 33530
rect 9210 33470 9305 33530
rect 9090 33250 9305 33470
rect 9090 33190 9150 33250
rect 9210 33190 9305 33250
rect 9090 33120 9305 33190
rect 9355 33530 9570 33740
rect 9355 33470 9450 33530
rect 9510 33470 9570 33530
rect 9355 33250 9570 33470
rect 9355 33190 9450 33250
rect 9510 33190 9570 33250
rect 9355 33120 9570 33190
rect 9970 33530 10185 33740
rect 9970 33470 10030 33530
rect 10090 33470 10185 33530
rect 9970 33250 10185 33470
rect 9970 33190 10030 33250
rect 10090 33190 10185 33250
rect 9970 33120 10185 33190
rect 10235 33530 10450 33740
rect 10235 33470 10330 33530
rect 10390 33470 10450 33530
rect 10235 33250 10450 33470
rect 10235 33190 10330 33250
rect 10390 33190 10450 33250
rect 10235 33120 10450 33190
rect 10560 33530 10775 33740
rect 10560 33470 10620 33530
rect 10680 33470 10775 33530
rect 10560 33250 10775 33470
rect 10560 33190 10620 33250
rect 10680 33190 10775 33250
rect 10560 33120 10775 33190
rect 10825 33530 11040 33740
rect 10825 33470 10920 33530
rect 10980 33470 11040 33530
rect 10825 33250 11040 33470
rect 10825 33190 10920 33250
rect 10980 33190 11040 33250
rect 10825 33120 11040 33190
rect 11150 33530 11365 33740
rect 11150 33470 11210 33530
rect 11270 33470 11365 33530
rect 11150 33250 11365 33470
rect 11150 33190 11210 33250
rect 11270 33190 11365 33250
rect 11150 33120 11365 33190
rect 11415 33530 11630 33740
rect 11415 33470 11510 33530
rect 11570 33470 11630 33530
rect 11415 33250 11630 33470
rect 11415 33190 11510 33250
rect 11570 33190 11630 33250
rect 11415 33120 11630 33190
rect 930 10050 1190 16050
rect 1260 10050 2120 16050
rect 2190 10050 2450 16050
rect 2520 10050 3380 16050
rect 3450 10050 3710 16050
rect 3780 10050 4640 16050
rect 4710 10050 4970 16050
rect 5040 10050 5900 16050
rect 5970 10050 6230 16050
rect 6300 10050 7160 16050
rect 7230 10050 7490 16050
rect 7560 10050 8420 16050
rect 8490 10050 8750 16050
rect 8820 10050 9680 16050
rect 9750 10050 10010 16050
rect 10080 10050 10940 16050
rect 11010 10050 11270 16050
<< ndcontact >>
rect 7830 33550 7890 33610
rect 7830 33430 7890 33490
rect 7830 33310 7890 33370
rect 8090 33550 8150 33610
rect 8090 33430 8150 33490
rect 8090 33310 8150 33370
rect 8350 33550 8410 33610
rect 8350 33430 8410 33490
rect 8350 33310 8410 33370
rect 8610 33550 8670 33610
rect 8610 33430 8670 33490
rect 8610 33310 8670 33370
rect 8870 33550 8930 33610
rect 8870 33430 8930 33490
rect 8870 33310 8930 33370
rect 9150 33470 9210 33530
rect 9150 33190 9210 33250
rect 9450 33470 9510 33530
rect 9450 33190 9510 33250
rect 10030 33470 10090 33530
rect 10030 33190 10090 33250
rect 10330 33470 10390 33530
rect 10330 33190 10390 33250
rect 10620 33470 10680 33530
rect 10620 33190 10680 33250
rect 10920 33470 10980 33530
rect 10920 33190 10980 33250
rect 11210 33470 11270 33530
rect 11210 33190 11270 33250
rect 11510 33470 11570 33530
rect 11510 33190 11570 33250
<< psubstratepdiff >>
rect 100 34030 12100 34210
rect 100 32730 300 34030
rect 11900 32730 12100 34030
rect 100 32550 12100 32730
rect 8790 31270 9005 31340
rect 8790 31210 8850 31270
rect 8910 31210 9005 31270
rect 8790 30990 9005 31210
rect 8790 30930 8850 30990
rect 8910 30930 9005 30990
rect 8790 30720 9005 30930
rect 9055 31270 9305 31340
rect 9055 31210 9150 31270
rect 9210 31210 9305 31270
rect 9055 30990 9305 31210
rect 9055 30930 9150 30990
rect 9210 30930 9305 30990
rect 9055 30720 9305 30930
rect 9355 31270 9570 31340
rect 9355 31210 9450 31270
rect 9510 31210 9570 31270
rect 9355 30990 9570 31210
rect 9355 30930 9450 30990
rect 9510 30930 9570 30990
rect 9355 30720 9570 30930
rect 9670 31270 9885 31340
rect 9670 31210 9730 31270
rect 9790 31210 9885 31270
rect 9670 30990 9885 31210
rect 9670 30930 9730 30990
rect 9790 30930 9885 30990
rect 9670 30720 9885 30930
rect 9935 31270 10185 31340
rect 9935 31210 10030 31270
rect 10090 31210 10185 31270
rect 9935 30990 10185 31210
rect 9935 30930 10030 30990
rect 10090 30930 10185 30990
rect 9935 30720 10185 30930
rect 10235 31270 10485 31340
rect 10235 31210 10330 31270
rect 10390 31210 10485 31270
rect 10235 30990 10485 31210
rect 10235 30930 10330 30990
rect 10390 30930 10485 30990
rect 10235 30720 10485 30930
rect 10535 31270 10785 31340
rect 10535 31210 10630 31270
rect 10690 31210 10785 31270
rect 10535 30990 10785 31210
rect 10535 30930 10630 30990
rect 10690 30930 10785 30990
rect 10535 30720 10785 30930
rect 10835 31270 11085 31340
rect 10835 31210 10930 31270
rect 10990 31210 11085 31270
rect 10835 30990 11085 31210
rect 10835 30930 10930 30990
rect 10990 30930 11085 30990
rect 10835 30720 11085 30930
rect 11135 31270 11385 31340
rect 11135 31210 11230 31270
rect 11290 31210 11385 31270
rect 11135 30990 11385 31210
rect 11135 30930 11230 30990
rect 11290 30930 11385 30990
rect 11135 30720 11385 30930
rect 11435 31270 11650 31340
rect 11435 31210 11530 31270
rect 11590 31210 11650 31270
rect 11435 30990 11650 31210
rect 11435 30930 11530 30990
rect 11590 30930 11650 30990
rect 11435 30720 11650 30930
rect 100 28750 12100 29750
rect 930 21350 1190 27350
rect 1260 21350 2120 27350
rect 2190 21350 2450 27350
rect 2520 21350 3380 27350
rect 3450 21350 3710 27350
rect 3780 21350 4640 27350
rect 4710 21350 4970 27350
rect 5040 21350 5900 27350
rect 5970 21350 6230 27350
rect 6300 21350 7160 27350
rect 7230 21350 7490 27350
rect 7560 21350 8420 27350
rect 8490 21350 8750 27350
rect 8820 21350 9680 27350
rect 9750 21350 10010 27350
rect 10080 21350 10940 27350
rect 11010 21350 11270 27350
rect 100 18950 12100 19950
rect 100 16450 12100 16950
rect 100 9650 600 16450
rect 11600 9650 12100 16450
rect 100 9150 12100 9650
<< nsubstratendiff >>
rect 100 31730 12100 31910
rect 100 30430 300 31730
rect 11900 30430 12100 31730
rect 100 30250 12100 30430
rect 100 27750 12100 28250
rect 100 20950 600 27750
rect 11600 20950 12100 27750
rect 100 20450 12100 20950
rect 100 17450 12100 18450
<< psubstratepcontact >>
rect 8850 31210 8910 31270
rect 8850 30930 8910 30990
rect 9150 31210 9210 31270
rect 9150 30930 9210 30990
rect 9450 31210 9510 31270
rect 9450 30930 9510 30990
rect 9730 31210 9790 31270
rect 9730 30930 9790 30990
rect 10030 31210 10090 31270
rect 10030 30930 10090 30990
rect 10330 31210 10390 31270
rect 10330 30930 10390 30990
rect 10630 31210 10690 31270
rect 10630 30930 10690 30990
rect 10930 31210 10990 31270
rect 10930 30930 10990 30990
rect 11230 31210 11290 31270
rect 11230 30930 11290 30990
rect 11530 31210 11590 31270
rect 11530 30930 11590 30990
<< polysilicon >>
rect 7910 33920 8070 33970
rect 7910 33860 7960 33920
rect 8020 33860 8070 33920
rect 7910 33810 8070 33860
rect 8170 33920 8330 33970
rect 8170 33860 8220 33920
rect 8280 33860 8330 33920
rect 8170 33810 8330 33860
rect 8430 33920 8590 33970
rect 8430 33860 8480 33920
rect 8540 33860 8590 33920
rect 8430 33810 8590 33860
rect 8690 33920 8850 33970
rect 8690 33860 8740 33920
rect 8800 33860 8850 33920
rect 8690 33810 8850 33860
rect 7965 33710 8015 33810
rect 8225 33710 8275 33810
rect 8485 33710 8535 33810
rect 8745 33710 8795 33810
rect 9305 33740 9355 33790
rect 10185 33740 10235 33790
rect 10775 33740 10825 33790
rect 11365 33740 11415 33790
rect 7965 33160 8015 33210
rect 8225 33160 8275 33210
rect 8485 33160 8535 33210
rect 8745 33160 8795 33210
rect 9305 33000 9355 33120
rect 10185 33000 10235 33120
rect 10775 33000 10825 33120
rect 11365 33000 11415 33120
rect 9250 32950 9410 33000
rect 9250 32890 9300 32950
rect 9360 32890 9410 32950
rect 9250 32840 9410 32890
rect 10130 32950 10290 33000
rect 10130 32890 10180 32950
rect 10240 32890 10290 32950
rect 10130 32840 10290 32890
rect 10720 32950 10880 33000
rect 10720 32890 10770 32950
rect 10830 32890 10880 32950
rect 10720 32840 10880 32890
rect 11310 32950 11470 33000
rect 11310 32890 11360 32950
rect 11420 32890 11470 32950
rect 11310 32840 11470 32890
rect 8950 31570 9110 31620
rect 8950 31510 9000 31570
rect 9060 31510 9110 31570
rect 8950 31460 9110 31510
rect 9250 31570 9410 31620
rect 9250 31510 9300 31570
rect 9360 31510 9410 31570
rect 9250 31460 9410 31510
rect 9830 31570 9990 31620
rect 9830 31510 9880 31570
rect 9940 31510 9990 31570
rect 9830 31460 9990 31510
rect 10130 31570 10290 31620
rect 10130 31510 10180 31570
rect 10240 31510 10290 31570
rect 10130 31460 10290 31510
rect 10430 31570 10590 31620
rect 10430 31510 10480 31570
rect 10540 31510 10590 31570
rect 10430 31460 10590 31510
rect 10730 31570 10890 31620
rect 10730 31510 10780 31570
rect 10840 31510 10890 31570
rect 10730 31460 10890 31510
rect 11030 31570 11190 31620
rect 11030 31510 11080 31570
rect 11140 31510 11190 31570
rect 11030 31460 11190 31510
rect 11330 31570 11490 31620
rect 11330 31510 11380 31570
rect 11440 31510 11490 31570
rect 11330 31460 11490 31510
rect 9005 30670 9055 31460
rect 9305 30670 9355 31460
rect 9885 30670 9935 31460
rect 10185 30670 10235 31460
rect 10485 30670 10535 31460
rect 10785 30670 10835 31460
rect 11085 30670 11135 31460
rect 11385 30670 11435 31460
rect 1135 27450 1315 27630
rect 2065 27450 2245 27630
rect 2395 27450 2575 27630
rect 3325 27450 3505 27630
rect 3655 27450 3835 27630
rect 4585 27450 4765 27630
rect 4915 27450 5095 27630
rect 5845 27450 6025 27630
rect 6175 27450 6355 27630
rect 7105 27450 7285 27630
rect 7435 27450 7615 27630
rect 8365 27450 8545 27630
rect 8695 27450 8875 27630
rect 9625 27450 9805 27630
rect 9955 27450 10135 27630
rect 10885 27450 11065 27630
rect 1190 21250 1260 27450
rect 2120 21250 2190 27450
rect 2450 21250 2520 27450
rect 3380 21250 3450 27450
rect 3710 21250 3780 27450
rect 4640 21250 4710 27450
rect 4970 21250 5040 27450
rect 5900 21250 5970 27450
rect 6230 21250 6300 27450
rect 7160 21250 7230 27450
rect 7490 21250 7560 27450
rect 8420 21250 8490 27450
rect 8750 21250 8820 27450
rect 9680 21250 9750 27450
rect 10010 21250 10080 27450
rect 10940 21250 11010 27450
rect 1135 16150 1315 16330
rect 2065 16150 2245 16330
rect 2395 16150 2575 16330
rect 3325 16150 3505 16330
rect 3655 16150 3835 16330
rect 4585 16150 4765 16330
rect 4915 16150 5095 16330
rect 5845 16150 6025 16330
rect 6175 16150 6355 16330
rect 7105 16150 7285 16330
rect 7435 16150 7615 16330
rect 8365 16150 8545 16330
rect 8695 16150 8875 16330
rect 9625 16150 9805 16330
rect 9955 16150 10135 16330
rect 10885 16150 11065 16330
rect 1190 16050 1260 16150
rect 2120 16050 2190 16150
rect 2450 16050 2520 16150
rect 3380 16050 3450 16150
rect 3710 16050 3780 16150
rect 4640 16050 4710 16150
rect 4970 16050 5040 16150
rect 5900 16050 5970 16150
rect 6230 16050 6300 16150
rect 7160 16050 7230 16150
rect 7490 16050 7560 16150
rect 8420 16050 8490 16150
rect 8750 16050 8820 16150
rect 9680 16050 9750 16150
rect 10010 16050 10080 16150
rect 10940 16050 11010 16150
rect 1190 9950 1260 10050
rect 2120 9950 2190 10050
rect 2450 9950 2520 10050
rect 3380 9950 3450 10050
rect 3710 9950 3780 10050
rect 4640 9950 4710 10050
rect 4970 9950 5040 10050
rect 5900 9950 5970 10050
rect 6230 9950 6300 10050
rect 7160 9950 7230 10050
rect 7490 9950 7560 10050
rect 8420 9950 8490 10050
rect 8750 9950 8820 10050
rect 9680 9950 9750 10050
rect 10010 9950 10080 10050
rect 10940 9950 11010 10050
<< polycontact >>
rect 7960 33860 8020 33920
rect 8220 33860 8280 33920
rect 8480 33860 8540 33920
rect 8740 33860 8800 33920
rect 9300 32890 9360 32950
rect 10180 32890 10240 32950
rect 10770 32890 10830 32950
rect 11360 32890 11420 32950
rect 9000 31510 9060 31570
rect 9300 31510 9360 31570
rect 9880 31510 9940 31570
rect 10180 31510 10240 31570
rect 10480 31510 10540 31570
rect 10780 31510 10840 31570
rect 11080 31510 11140 31570
rect 11380 31510 11440 31570
<< genericcontact >>
rect 350 34090 410 34150
rect 470 34090 530 34150
rect 590 34090 650 34150
rect 710 34090 770 34150
rect 830 34090 890 34150
rect 950 34090 1010 34150
rect 1070 34090 1130 34150
rect 1190 34090 1250 34150
rect 1310 34090 1370 34150
rect 1430 34090 1490 34150
rect 1550 34090 1610 34150
rect 1670 34090 1730 34150
rect 1790 34090 1850 34150
rect 1910 34090 1970 34150
rect 2030 34090 2090 34150
rect 2150 34090 2210 34150
rect 2270 34090 2330 34150
rect 2390 34090 2450 34150
rect 2510 34090 2570 34150
rect 2630 34090 2690 34150
rect 2750 34090 2810 34150
rect 2870 34090 2930 34150
rect 2990 34090 3050 34150
rect 3110 34090 3170 34150
rect 3230 34090 3290 34150
rect 3350 34090 3410 34150
rect 3470 34090 3530 34150
rect 3590 34090 3650 34150
rect 3710 34090 3770 34150
rect 3830 34090 3890 34150
rect 3950 34090 4010 34150
rect 4070 34090 4130 34150
rect 4190 34090 4250 34150
rect 4310 34090 4370 34150
rect 4430 34090 4490 34150
rect 4550 34090 4610 34150
rect 4670 34090 4730 34150
rect 4790 34090 4850 34150
rect 4910 34090 4970 34150
rect 5030 34090 5090 34150
rect 5150 34090 5210 34150
rect 5270 34090 5330 34150
rect 5390 34090 5450 34150
rect 5510 34090 5570 34150
rect 5630 34090 5690 34150
rect 5750 34090 5810 34150
rect 5870 34090 5930 34150
rect 5990 34090 6050 34150
rect 6110 34090 6170 34150
rect 6230 34090 6290 34150
rect 6350 34090 6410 34150
rect 6470 34090 6530 34150
rect 6590 34090 6650 34150
rect 6710 34090 6770 34150
rect 6830 34090 6890 34150
rect 6950 34090 7010 34150
rect 7070 34090 7130 34150
rect 7190 34090 7250 34150
rect 7310 34090 7370 34150
rect 7430 34090 7490 34150
rect 7550 34090 7610 34150
rect 7670 34090 7730 34150
rect 7790 34090 7850 34150
rect 7910 34090 7970 34150
rect 8030 34090 8090 34150
rect 8150 34090 8210 34150
rect 8270 34090 8330 34150
rect 8390 34090 8450 34150
rect 8510 34090 8570 34150
rect 8630 34090 8690 34150
rect 8750 34090 8810 34150
rect 8870 34090 8930 34150
rect 8990 34090 9050 34150
rect 9110 34090 9170 34150
rect 9230 34090 9290 34150
rect 9350 34090 9410 34150
rect 9470 34090 9530 34150
rect 9590 34090 9650 34150
rect 9710 34090 9770 34150
rect 9830 34090 9890 34150
rect 9950 34090 10010 34150
rect 10070 34090 10130 34150
rect 10190 34090 10250 34150
rect 10310 34090 10370 34150
rect 10430 34090 10490 34150
rect 10550 34090 10610 34150
rect 10670 34090 10730 34150
rect 10790 34090 10850 34150
rect 10910 34090 10970 34150
rect 11030 34090 11090 34150
rect 11150 34090 11210 34150
rect 11270 34090 11330 34150
rect 11390 34090 11450 34150
rect 11510 34090 11570 34150
rect 11630 34090 11690 34150
rect 11750 34090 11810 34150
rect 170 33880 230 33940
rect 11970 33880 12030 33940
rect 170 33600 230 33660
rect 10330 33610 10390 33670
rect 10920 33610 10980 33670
rect 11970 33600 12030 33660
rect 170 33320 230 33380
rect 10330 33330 10390 33390
rect 10920 33330 10980 33390
rect 11970 33320 12030 33380
rect 170 33040 230 33100
rect 11970 33040 12030 33100
rect 170 32760 230 32820
rect 11970 32760 12030 32820
rect 350 32610 410 32670
rect 470 32610 530 32670
rect 590 32610 650 32670
rect 710 32610 770 32670
rect 830 32610 890 32670
rect 950 32610 1010 32670
rect 1070 32610 1130 32670
rect 1190 32610 1250 32670
rect 1310 32610 1370 32670
rect 1430 32610 1490 32670
rect 1550 32610 1610 32670
rect 1670 32610 1730 32670
rect 1790 32610 1850 32670
rect 1910 32610 1970 32670
rect 2030 32610 2090 32670
rect 2150 32610 2210 32670
rect 2270 32610 2330 32670
rect 2390 32610 2450 32670
rect 2510 32610 2570 32670
rect 2630 32610 2690 32670
rect 2750 32610 2810 32670
rect 2870 32610 2930 32670
rect 2990 32610 3050 32670
rect 3110 32610 3170 32670
rect 3230 32610 3290 32670
rect 3350 32610 3410 32670
rect 3470 32610 3530 32670
rect 3590 32610 3650 32670
rect 3710 32610 3770 32670
rect 3830 32610 3890 32670
rect 3950 32610 4010 32670
rect 4070 32610 4130 32670
rect 4190 32610 4250 32670
rect 4310 32610 4370 32670
rect 4430 32610 4490 32670
rect 4550 32610 4610 32670
rect 4670 32610 4730 32670
rect 4790 32610 4850 32670
rect 4910 32610 4970 32670
rect 5030 32610 5090 32670
rect 5150 32610 5210 32670
rect 5270 32610 5330 32670
rect 5390 32610 5450 32670
rect 5510 32610 5570 32670
rect 5630 32610 5690 32670
rect 5750 32610 5810 32670
rect 5870 32610 5930 32670
rect 5990 32610 6050 32670
rect 6110 32610 6170 32670
rect 6230 32610 6290 32670
rect 6350 32610 6410 32670
rect 6470 32610 6530 32670
rect 6590 32610 6650 32670
rect 6710 32610 6770 32670
rect 6830 32610 6890 32670
rect 6950 32610 7010 32670
rect 7070 32610 7130 32670
rect 7190 32610 7250 32670
rect 7310 32610 7370 32670
rect 7430 32610 7490 32670
rect 7550 32610 7610 32670
rect 7670 32610 7730 32670
rect 7790 32610 7850 32670
rect 7910 32610 7970 32670
rect 8030 32610 8090 32670
rect 8150 32610 8210 32670
rect 8270 32610 8330 32670
rect 8390 32610 8450 32670
rect 8510 32610 8570 32670
rect 8630 32610 8690 32670
rect 8750 32610 8810 32670
rect 8870 32610 8930 32670
rect 8990 32610 9050 32670
rect 9110 32610 9170 32670
rect 9230 32610 9290 32670
rect 9350 32610 9410 32670
rect 9470 32610 9530 32670
rect 9590 32610 9650 32670
rect 9710 32610 9770 32670
rect 9830 32610 9890 32670
rect 9950 32610 10010 32670
rect 10070 32610 10130 32670
rect 10190 32610 10250 32670
rect 10310 32610 10370 32670
rect 10430 32610 10490 32670
rect 10550 32610 10610 32670
rect 10670 32610 10730 32670
rect 10790 32610 10850 32670
rect 10910 32610 10970 32670
rect 11030 32610 11090 32670
rect 11150 32610 11210 32670
rect 11270 32610 11330 32670
rect 11390 32610 11450 32670
rect 11510 32610 11570 32670
rect 11630 32610 11690 32670
rect 11750 32610 11810 32670
rect 350 31790 410 31850
rect 470 31790 530 31850
rect 590 31790 650 31850
rect 710 31790 770 31850
rect 830 31790 890 31850
rect 950 31790 1010 31850
rect 1070 31790 1130 31850
rect 1190 31790 1250 31850
rect 1310 31790 1370 31850
rect 1430 31790 1490 31850
rect 1550 31790 1610 31850
rect 1670 31790 1730 31850
rect 1790 31790 1850 31850
rect 1910 31790 1970 31850
rect 2030 31790 2090 31850
rect 2150 31790 2210 31850
rect 2270 31790 2330 31850
rect 2390 31790 2450 31850
rect 2510 31790 2570 31850
rect 2630 31790 2690 31850
rect 2750 31790 2810 31850
rect 2870 31790 2930 31850
rect 2990 31790 3050 31850
rect 3110 31790 3170 31850
rect 3230 31790 3290 31850
rect 3350 31790 3410 31850
rect 3470 31790 3530 31850
rect 3590 31790 3650 31850
rect 3710 31790 3770 31850
rect 3830 31790 3890 31850
rect 3950 31790 4010 31850
rect 4070 31790 4130 31850
rect 4190 31790 4250 31850
rect 4310 31790 4370 31850
rect 4430 31790 4490 31850
rect 4550 31790 4610 31850
rect 4670 31790 4730 31850
rect 4790 31790 4850 31850
rect 4910 31790 4970 31850
rect 5030 31790 5090 31850
rect 5150 31790 5210 31850
rect 5270 31790 5330 31850
rect 5390 31790 5450 31850
rect 5510 31790 5570 31850
rect 5630 31790 5690 31850
rect 5750 31790 5810 31850
rect 5870 31790 5930 31850
rect 5990 31790 6050 31850
rect 6110 31790 6170 31850
rect 6230 31790 6290 31850
rect 6350 31790 6410 31850
rect 6470 31790 6530 31850
rect 6590 31790 6650 31850
rect 6710 31790 6770 31850
rect 6830 31790 6890 31850
rect 6950 31790 7010 31850
rect 7070 31790 7130 31850
rect 7190 31790 7250 31850
rect 7310 31790 7370 31850
rect 7430 31790 7490 31850
rect 7550 31790 7610 31850
rect 7670 31790 7730 31850
rect 7790 31790 7850 31850
rect 7910 31790 7970 31850
rect 8030 31790 8090 31850
rect 8150 31790 8210 31850
rect 8270 31790 8330 31850
rect 8390 31790 8450 31850
rect 8510 31790 8570 31850
rect 8630 31790 8690 31850
rect 8750 31790 8810 31850
rect 8870 31790 8930 31850
rect 8990 31790 9050 31850
rect 9110 31790 9170 31850
rect 9230 31790 9290 31850
rect 9350 31790 9410 31850
rect 9470 31790 9530 31850
rect 9590 31790 9650 31850
rect 9710 31790 9770 31850
rect 9830 31790 9890 31850
rect 9950 31790 10010 31850
rect 10070 31790 10130 31850
rect 10190 31790 10250 31850
rect 10310 31790 10370 31850
rect 10430 31790 10490 31850
rect 10550 31790 10610 31850
rect 10670 31790 10730 31850
rect 10790 31790 10850 31850
rect 10910 31790 10970 31850
rect 11030 31790 11090 31850
rect 11150 31790 11210 31850
rect 11270 31790 11330 31850
rect 11390 31790 11450 31850
rect 11510 31790 11570 31850
rect 11630 31790 11690 31850
rect 11750 31790 11810 31850
rect 170 31580 230 31640
rect 11970 31580 12030 31640
rect 170 31300 230 31360
rect 11970 31300 12030 31360
rect 5890 31085 5950 31145
rect 8350 31085 8410 31145
rect 170 31020 230 31080
rect 8850 31070 8910 31130
rect 9730 31070 9790 31130
rect 10330 31070 10390 31130
rect 10930 31070 10990 31130
rect 5890 30965 5950 31025
rect 8350 30965 8410 31025
rect 11970 31020 12030 31080
rect 170 30740 230 30800
rect 8850 30790 8910 30850
rect 9730 30790 9790 30850
rect 10330 30790 10390 30850
rect 10930 30790 10990 30850
rect 11970 30740 12030 30800
rect 170 30460 230 30520
rect 11970 30460 12030 30520
rect 350 30310 410 30370
rect 470 30310 530 30370
rect 590 30310 650 30370
rect 710 30310 770 30370
rect 830 30310 890 30370
rect 950 30310 1010 30370
rect 1070 30310 1130 30370
rect 1190 30310 1250 30370
rect 1310 30310 1370 30370
rect 1430 30310 1490 30370
rect 1550 30310 1610 30370
rect 1670 30310 1730 30370
rect 1790 30310 1850 30370
rect 1910 30310 1970 30370
rect 2030 30310 2090 30370
rect 2150 30310 2210 30370
rect 2270 30310 2330 30370
rect 2390 30310 2450 30370
rect 2510 30310 2570 30370
rect 2630 30310 2690 30370
rect 2750 30310 2810 30370
rect 2870 30310 2930 30370
rect 2990 30310 3050 30370
rect 3110 30310 3170 30370
rect 3230 30310 3290 30370
rect 3350 30310 3410 30370
rect 3470 30310 3530 30370
rect 3590 30310 3650 30370
rect 3710 30310 3770 30370
rect 3830 30310 3890 30370
rect 3950 30310 4010 30370
rect 4070 30310 4130 30370
rect 4190 30310 4250 30370
rect 4310 30310 4370 30370
rect 4430 30310 4490 30370
rect 4550 30310 4610 30370
rect 4670 30310 4730 30370
rect 4790 30310 4850 30370
rect 4910 30310 4970 30370
rect 5030 30310 5090 30370
rect 5150 30310 5210 30370
rect 5270 30310 5330 30370
rect 5390 30310 5450 30370
rect 5510 30310 5570 30370
rect 5630 30310 5690 30370
rect 5750 30310 5810 30370
rect 5870 30310 5930 30370
rect 5990 30310 6050 30370
rect 6110 30310 6170 30370
rect 6230 30310 6290 30370
rect 6350 30310 6410 30370
rect 6470 30310 6530 30370
rect 6590 30310 6650 30370
rect 6710 30310 6770 30370
rect 6830 30310 6890 30370
rect 6950 30310 7010 30370
rect 7070 30310 7130 30370
rect 7190 30310 7250 30370
rect 7310 30310 7370 30370
rect 7430 30310 7490 30370
rect 7550 30310 7610 30370
rect 7670 30310 7730 30370
rect 7790 30310 7850 30370
rect 7910 30310 7970 30370
rect 8030 30310 8090 30370
rect 8150 30310 8210 30370
rect 8270 30310 8330 30370
rect 8390 30310 8450 30370
rect 8510 30310 8570 30370
rect 8630 30310 8690 30370
rect 8750 30310 8810 30370
rect 8870 30310 8930 30370
rect 8990 30310 9050 30370
rect 9110 30310 9170 30370
rect 9230 30310 9290 30370
rect 9350 30310 9410 30370
rect 9470 30310 9530 30370
rect 9590 30310 9650 30370
rect 9710 30310 9770 30370
rect 9830 30310 9890 30370
rect 9950 30310 10010 30370
rect 10070 30310 10130 30370
rect 10190 30310 10250 30370
rect 10310 30310 10370 30370
rect 10430 30310 10490 30370
rect 10550 30310 10610 30370
rect 10670 30310 10730 30370
rect 10790 30310 10850 30370
rect 10910 30310 10970 30370
rect 11030 30310 11090 30370
rect 11150 30310 11210 30370
rect 11270 30310 11330 30370
rect 11390 30310 11450 30370
rect 11510 30310 11570 30370
rect 11630 30310 11690 30370
rect 11750 30310 11810 30370
rect 350 29575 410 29635
rect 530 29575 590 29635
rect 710 29575 770 29635
rect 890 29575 950 29635
rect 1070 29575 1130 29635
rect 1250 29575 1310 29635
rect 1430 29575 1490 29635
rect 1610 29575 1670 29635
rect 1790 29575 1850 29635
rect 1970 29575 2030 29635
rect 2150 29575 2210 29635
rect 2330 29575 2390 29635
rect 2510 29575 2570 29635
rect 2690 29575 2750 29635
rect 2870 29575 2930 29635
rect 3050 29575 3110 29635
rect 3230 29575 3290 29635
rect 3410 29575 3470 29635
rect 3590 29575 3650 29635
rect 3770 29575 3830 29635
rect 3950 29575 4010 29635
rect 4130 29575 4190 29635
rect 4310 29575 4370 29635
rect 4490 29575 4550 29635
rect 4670 29575 4730 29635
rect 5750 29575 5810 29635
rect 5930 29575 5990 29635
rect 6110 29575 6170 29635
rect 6290 29575 6350 29635
rect 6470 29575 6530 29635
rect 6650 29575 6710 29635
rect 6830 29575 6890 29635
rect 7010 29575 7070 29635
rect 7190 29575 7250 29635
rect 7370 29575 7430 29635
rect 7550 29575 7610 29635
rect 7730 29575 7790 29635
rect 8810 29575 8870 29635
rect 8990 29575 9050 29635
rect 9170 29575 9230 29635
rect 9350 29575 9410 29635
rect 9530 29575 9590 29635
rect 9710 29575 9770 29635
rect 9890 29575 9950 29635
rect 10070 29575 10130 29635
rect 10250 29575 10310 29635
rect 10430 29575 10490 29635
rect 10610 29575 10670 29635
rect 10790 29575 10850 29635
rect 10970 29575 11030 29635
rect 11150 29575 11210 29635
rect 11330 29575 11390 29635
rect 11510 29575 11570 29635
rect 11690 29575 11750 29635
rect 11870 29575 11930 29635
rect 350 29395 410 29455
rect 530 29395 590 29455
rect 710 29395 770 29455
rect 890 29395 950 29455
rect 1070 29395 1130 29455
rect 1250 29395 1310 29455
rect 1430 29395 1490 29455
rect 1610 29395 1670 29455
rect 1790 29395 1850 29455
rect 1970 29395 2030 29455
rect 2150 29395 2210 29455
rect 2330 29395 2390 29455
rect 2510 29395 2570 29455
rect 2690 29395 2750 29455
rect 2870 29395 2930 29455
rect 3050 29395 3110 29455
rect 3230 29395 3290 29455
rect 3410 29395 3470 29455
rect 3590 29395 3650 29455
rect 3770 29395 3830 29455
rect 3950 29395 4010 29455
rect 4130 29395 4190 29455
rect 4310 29395 4370 29455
rect 4490 29395 4550 29455
rect 4670 29395 4730 29455
rect 5750 29395 5810 29455
rect 5930 29395 5990 29455
rect 6110 29395 6170 29455
rect 6290 29395 6350 29455
rect 6470 29395 6530 29455
rect 6650 29395 6710 29455
rect 6830 29395 6890 29455
rect 7010 29395 7070 29455
rect 7190 29395 7250 29455
rect 7370 29395 7430 29455
rect 7550 29395 7610 29455
rect 7730 29395 7790 29455
rect 8810 29395 8870 29455
rect 8990 29395 9050 29455
rect 9170 29395 9230 29455
rect 9350 29395 9410 29455
rect 9530 29395 9590 29455
rect 9710 29395 9770 29455
rect 9890 29395 9950 29455
rect 10070 29395 10130 29455
rect 10250 29395 10310 29455
rect 10430 29395 10490 29455
rect 10610 29395 10670 29455
rect 10790 29395 10850 29455
rect 10970 29395 11030 29455
rect 11150 29395 11210 29455
rect 11330 29395 11390 29455
rect 11510 29395 11570 29455
rect 11690 29395 11750 29455
rect 11870 29395 11930 29455
rect 350 29215 410 29275
rect 530 29215 590 29275
rect 710 29215 770 29275
rect 890 29215 950 29275
rect 1070 29215 1130 29275
rect 1250 29215 1310 29275
rect 1430 29215 1490 29275
rect 1610 29215 1670 29275
rect 1790 29215 1850 29275
rect 1970 29215 2030 29275
rect 2150 29215 2210 29275
rect 2330 29215 2390 29275
rect 2510 29215 2570 29275
rect 2690 29215 2750 29275
rect 2870 29215 2930 29275
rect 3050 29215 3110 29275
rect 3230 29215 3290 29275
rect 3410 29215 3470 29275
rect 3590 29215 3650 29275
rect 3770 29215 3830 29275
rect 3950 29215 4010 29275
rect 4130 29215 4190 29275
rect 4310 29215 4370 29275
rect 4490 29215 4550 29275
rect 4670 29215 4730 29275
rect 5750 29215 5810 29275
rect 5930 29215 5990 29275
rect 6110 29215 6170 29275
rect 6290 29215 6350 29275
rect 6470 29215 6530 29275
rect 6650 29215 6710 29275
rect 6830 29215 6890 29275
rect 7010 29215 7070 29275
rect 7190 29215 7250 29275
rect 7370 29215 7430 29275
rect 7550 29215 7610 29275
rect 7730 29215 7790 29275
rect 8810 29215 8870 29275
rect 8990 29215 9050 29275
rect 9170 29215 9230 29275
rect 9350 29215 9410 29275
rect 9530 29215 9590 29275
rect 9710 29215 9770 29275
rect 9890 29215 9950 29275
rect 10070 29215 10130 29275
rect 10250 29215 10310 29275
rect 10430 29215 10490 29275
rect 10610 29215 10670 29275
rect 10790 29215 10850 29275
rect 10970 29215 11030 29275
rect 11150 29215 11210 29275
rect 11330 29215 11390 29275
rect 11510 29215 11570 29275
rect 11690 29215 11750 29275
rect 11870 29215 11930 29275
rect 350 29035 410 29095
rect 530 29035 590 29095
rect 710 29035 770 29095
rect 890 29035 950 29095
rect 1070 29035 1130 29095
rect 1250 29035 1310 29095
rect 1430 29035 1490 29095
rect 1610 29035 1670 29095
rect 1790 29035 1850 29095
rect 1970 29035 2030 29095
rect 2150 29035 2210 29095
rect 2330 29035 2390 29095
rect 2510 29035 2570 29095
rect 2690 29035 2750 29095
rect 2870 29035 2930 29095
rect 3050 29035 3110 29095
rect 3230 29035 3290 29095
rect 3410 29035 3470 29095
rect 3590 29035 3650 29095
rect 3770 29035 3830 29095
rect 3950 29035 4010 29095
rect 4130 29035 4190 29095
rect 4310 29035 4370 29095
rect 4490 29035 4550 29095
rect 4670 29035 4730 29095
rect 5750 29035 5810 29095
rect 5930 29035 5990 29095
rect 6110 29035 6170 29095
rect 6290 29035 6350 29095
rect 6470 29035 6530 29095
rect 6650 29035 6710 29095
rect 6830 29035 6890 29095
rect 7010 29035 7070 29095
rect 7190 29035 7250 29095
rect 7370 29035 7430 29095
rect 7550 29035 7610 29095
rect 7730 29035 7790 29095
rect 8810 29035 8870 29095
rect 8990 29035 9050 29095
rect 9170 29035 9230 29095
rect 9350 29035 9410 29095
rect 9530 29035 9590 29095
rect 9710 29035 9770 29095
rect 9890 29035 9950 29095
rect 10070 29035 10130 29095
rect 10250 29035 10310 29095
rect 10430 29035 10490 29095
rect 10610 29035 10670 29095
rect 10790 29035 10850 29095
rect 10970 29035 11030 29095
rect 11150 29035 11210 29095
rect 11330 29035 11390 29095
rect 11510 29035 11570 29095
rect 11690 29035 11750 29095
rect 11870 29035 11930 29095
rect 350 28855 410 28915
rect 530 28855 590 28915
rect 710 28855 770 28915
rect 890 28855 950 28915
rect 1070 28855 1130 28915
rect 1250 28855 1310 28915
rect 1430 28855 1490 28915
rect 1610 28855 1670 28915
rect 1790 28855 1850 28915
rect 1970 28855 2030 28915
rect 2150 28855 2210 28915
rect 2330 28855 2390 28915
rect 2510 28855 2570 28915
rect 2690 28855 2750 28915
rect 2870 28855 2930 28915
rect 3050 28855 3110 28915
rect 3230 28855 3290 28915
rect 3410 28855 3470 28915
rect 3590 28855 3650 28915
rect 3770 28855 3830 28915
rect 3950 28855 4010 28915
rect 4130 28855 4190 28915
rect 4310 28855 4370 28915
rect 4490 28855 4550 28915
rect 4670 28855 4730 28915
rect 5750 28855 5810 28915
rect 5930 28855 5990 28915
rect 6110 28855 6170 28915
rect 6290 28855 6350 28915
rect 6470 28855 6530 28915
rect 6650 28855 6710 28915
rect 6830 28855 6890 28915
rect 7010 28855 7070 28915
rect 7190 28855 7250 28915
rect 7370 28855 7430 28915
rect 7550 28855 7610 28915
rect 7730 28855 7790 28915
rect 8810 28855 8870 28915
rect 8990 28855 9050 28915
rect 9170 28855 9230 28915
rect 9350 28855 9410 28915
rect 9530 28855 9590 28915
rect 9710 28855 9770 28915
rect 9890 28855 9950 28915
rect 10070 28855 10130 28915
rect 10250 28855 10310 28915
rect 10430 28855 10490 28915
rect 10610 28855 10670 28915
rect 10790 28855 10850 28915
rect 10970 28855 11030 28915
rect 11150 28855 11210 28915
rect 11330 28855 11390 28915
rect 11510 28855 11570 28915
rect 11690 28855 11750 28915
rect 11870 28855 11930 28915
rect 320 28100 380 28160
rect 660 28090 720 28150
rect 780 28090 840 28150
rect 900 28090 960 28150
rect 1020 28090 1080 28150
rect 1140 28090 1200 28150
rect 1260 28090 1320 28150
rect 1380 28090 1440 28150
rect 1500 28090 1560 28150
rect 1620 28090 1680 28150
rect 1740 28090 1800 28150
rect 1860 28090 1920 28150
rect 1980 28090 2040 28150
rect 2100 28090 2160 28150
rect 2220 28090 2280 28150
rect 2340 28090 2400 28150
rect 2460 28090 2520 28150
rect 2580 28090 2640 28150
rect 2700 28090 2760 28150
rect 2820 28090 2880 28150
rect 2940 28090 3000 28150
rect 3060 28090 3120 28150
rect 3180 28090 3240 28150
rect 3300 28090 3360 28150
rect 3420 28090 3480 28150
rect 3540 28090 3600 28150
rect 3660 28090 3720 28150
rect 3780 28090 3840 28150
rect 3900 28090 3960 28150
rect 4020 28090 4080 28150
rect 4140 28090 4200 28150
rect 4260 28090 4320 28150
rect 4380 28090 4440 28150
rect 4500 28090 4560 28150
rect 4620 28090 4680 28150
rect 4740 28090 4800 28150
rect 4860 28090 4920 28150
rect 4980 28090 5040 28150
rect 5100 28090 5160 28150
rect 5220 28090 5280 28150
rect 5340 28090 5400 28150
rect 5460 28090 5520 28150
rect 5580 28090 5640 28150
rect 5700 28090 5760 28150
rect 5820 28090 5880 28150
rect 5940 28090 6000 28150
rect 6060 28090 6120 28150
rect 6180 28090 6240 28150
rect 6300 28090 6360 28150
rect 6420 28090 6480 28150
rect 6540 28090 6600 28150
rect 6660 28090 6720 28150
rect 6780 28090 6840 28150
rect 6900 28090 6960 28150
rect 7020 28090 7080 28150
rect 7140 28090 7200 28150
rect 7260 28090 7320 28150
rect 7380 28090 7440 28150
rect 7500 28090 7560 28150
rect 7620 28090 7680 28150
rect 7740 28090 7800 28150
rect 7860 28090 7920 28150
rect 7980 28090 8040 28150
rect 8100 28090 8160 28150
rect 8220 28090 8280 28150
rect 8340 28090 8400 28150
rect 8460 28090 8520 28150
rect 8580 28090 8640 28150
rect 8700 28090 8760 28150
rect 8820 28090 8880 28150
rect 8940 28090 9000 28150
rect 9060 28090 9120 28150
rect 9180 28090 9240 28150
rect 9300 28090 9360 28150
rect 9420 28090 9480 28150
rect 9540 28090 9600 28150
rect 9660 28090 9720 28150
rect 9780 28090 9840 28150
rect 9900 28090 9960 28150
rect 10020 28090 10080 28150
rect 10140 28090 10200 28150
rect 10260 28090 10320 28150
rect 10380 28090 10440 28150
rect 10500 28090 10560 28150
rect 10620 28090 10680 28150
rect 10740 28090 10800 28150
rect 10860 28090 10920 28150
rect 10980 28090 11040 28150
rect 11100 28090 11160 28150
rect 11220 28090 11280 28150
rect 11340 28090 11400 28150
rect 11460 28090 11520 28150
rect 11820 28100 11880 28160
rect 320 27920 380 27980
rect 660 27970 720 28030
rect 780 27970 840 28030
rect 900 27970 960 28030
rect 1020 27970 1080 28030
rect 1140 27970 1200 28030
rect 1260 27970 1320 28030
rect 1380 27970 1440 28030
rect 1500 27970 1560 28030
rect 1620 27970 1680 28030
rect 1740 27970 1800 28030
rect 1860 27970 1920 28030
rect 1980 27970 2040 28030
rect 2100 27970 2160 28030
rect 2220 27970 2280 28030
rect 2340 27970 2400 28030
rect 2460 27970 2520 28030
rect 2580 27970 2640 28030
rect 2700 27970 2760 28030
rect 2820 27970 2880 28030
rect 2940 27970 3000 28030
rect 3060 27970 3120 28030
rect 3180 27970 3240 28030
rect 3300 27970 3360 28030
rect 3420 27970 3480 28030
rect 3540 27970 3600 28030
rect 3660 27970 3720 28030
rect 3780 27970 3840 28030
rect 3900 27970 3960 28030
rect 4020 27970 4080 28030
rect 4140 27970 4200 28030
rect 4260 27970 4320 28030
rect 4380 27970 4440 28030
rect 4500 27970 4560 28030
rect 4620 27970 4680 28030
rect 4740 27970 4800 28030
rect 4860 27970 4920 28030
rect 4980 27970 5040 28030
rect 5100 27970 5160 28030
rect 5220 27970 5280 28030
rect 5340 27970 5400 28030
rect 5460 27970 5520 28030
rect 5580 27970 5640 28030
rect 5700 27970 5760 28030
rect 5820 27970 5880 28030
rect 5940 27970 6000 28030
rect 6060 27970 6120 28030
rect 6180 27970 6240 28030
rect 6300 27970 6360 28030
rect 6420 27970 6480 28030
rect 6540 27970 6600 28030
rect 6660 27970 6720 28030
rect 6780 27970 6840 28030
rect 6900 27970 6960 28030
rect 7020 27970 7080 28030
rect 7140 27970 7200 28030
rect 7260 27970 7320 28030
rect 7380 27970 7440 28030
rect 7500 27970 7560 28030
rect 7620 27970 7680 28030
rect 7740 27970 7800 28030
rect 7860 27970 7920 28030
rect 7980 27970 8040 28030
rect 8100 27970 8160 28030
rect 8220 27970 8280 28030
rect 8340 27970 8400 28030
rect 8460 27970 8520 28030
rect 8580 27970 8640 28030
rect 8700 27970 8760 28030
rect 8820 27970 8880 28030
rect 8940 27970 9000 28030
rect 9060 27970 9120 28030
rect 9180 27970 9240 28030
rect 9300 27970 9360 28030
rect 9420 27970 9480 28030
rect 9540 27970 9600 28030
rect 9660 27970 9720 28030
rect 9780 27970 9840 28030
rect 9900 27970 9960 28030
rect 10020 27970 10080 28030
rect 10140 27970 10200 28030
rect 10260 27970 10320 28030
rect 10380 27970 10440 28030
rect 10500 27970 10560 28030
rect 10620 27970 10680 28030
rect 10740 27970 10800 28030
rect 10860 27970 10920 28030
rect 10980 27970 11040 28030
rect 11100 27970 11160 28030
rect 11220 27970 11280 28030
rect 11340 27970 11400 28030
rect 11460 27970 11520 28030
rect 11820 27920 11880 27980
rect 660 27850 720 27910
rect 780 27850 840 27910
rect 900 27850 960 27910
rect 1020 27850 1080 27910
rect 1140 27850 1200 27910
rect 1260 27850 1320 27910
rect 1380 27850 1440 27910
rect 1500 27850 1560 27910
rect 1620 27850 1680 27910
rect 1740 27850 1800 27910
rect 1860 27850 1920 27910
rect 1980 27850 2040 27910
rect 2100 27850 2160 27910
rect 2220 27850 2280 27910
rect 2340 27850 2400 27910
rect 2460 27850 2520 27910
rect 2580 27850 2640 27910
rect 2700 27850 2760 27910
rect 2820 27850 2880 27910
rect 2940 27850 3000 27910
rect 3060 27850 3120 27910
rect 3180 27850 3240 27910
rect 3300 27850 3360 27910
rect 3420 27850 3480 27910
rect 3540 27850 3600 27910
rect 3660 27850 3720 27910
rect 3780 27850 3840 27910
rect 3900 27850 3960 27910
rect 4020 27850 4080 27910
rect 4140 27850 4200 27910
rect 4260 27850 4320 27910
rect 4380 27850 4440 27910
rect 4500 27850 4560 27910
rect 4620 27850 4680 27910
rect 4740 27850 4800 27910
rect 4860 27850 4920 27910
rect 4980 27850 5040 27910
rect 5100 27850 5160 27910
rect 5220 27850 5280 27910
rect 5340 27850 5400 27910
rect 5460 27850 5520 27910
rect 5580 27850 5640 27910
rect 5700 27850 5760 27910
rect 5820 27850 5880 27910
rect 5940 27850 6000 27910
rect 6060 27850 6120 27910
rect 6180 27850 6240 27910
rect 6300 27850 6360 27910
rect 6420 27850 6480 27910
rect 6540 27850 6600 27910
rect 6660 27850 6720 27910
rect 6780 27850 6840 27910
rect 6900 27850 6960 27910
rect 7020 27850 7080 27910
rect 7140 27850 7200 27910
rect 7260 27850 7320 27910
rect 7380 27850 7440 27910
rect 7500 27850 7560 27910
rect 7620 27850 7680 27910
rect 7740 27850 7800 27910
rect 7860 27850 7920 27910
rect 7980 27850 8040 27910
rect 8100 27850 8160 27910
rect 8220 27850 8280 27910
rect 8340 27850 8400 27910
rect 8460 27850 8520 27910
rect 8580 27850 8640 27910
rect 8700 27850 8760 27910
rect 8820 27850 8880 27910
rect 8940 27850 9000 27910
rect 9060 27850 9120 27910
rect 9180 27850 9240 27910
rect 9300 27850 9360 27910
rect 9420 27850 9480 27910
rect 9540 27850 9600 27910
rect 9660 27850 9720 27910
rect 9780 27850 9840 27910
rect 9900 27850 9960 27910
rect 10020 27850 10080 27910
rect 10140 27850 10200 27910
rect 10260 27850 10320 27910
rect 10380 27850 10440 27910
rect 10500 27850 10560 27910
rect 10620 27850 10680 27910
rect 10740 27850 10800 27910
rect 10860 27850 10920 27910
rect 10980 27850 11040 27910
rect 11100 27850 11160 27910
rect 11220 27850 11280 27910
rect 11340 27850 11400 27910
rect 11460 27850 11520 27910
rect 320 27740 380 27800
rect 11820 27740 11880 27800
rect 320 27560 380 27620
rect 1195 27510 1255 27570
rect 2125 27510 2185 27570
rect 2455 27510 2515 27570
rect 3385 27510 3445 27570
rect 3715 27510 3775 27570
rect 4645 27510 4705 27570
rect 4975 27510 5035 27570
rect 5905 27510 5965 27570
rect 6235 27510 6295 27570
rect 7165 27510 7225 27570
rect 7495 27510 7555 27570
rect 8425 27510 8485 27570
rect 8755 27510 8815 27570
rect 9685 27510 9745 27570
rect 10015 27510 10075 27570
rect 10945 27510 11005 27570
rect 11820 27560 11880 27620
rect 320 27380 380 27440
rect 11820 27380 11880 27440
rect 320 27200 380 27260
rect 11820 27200 11880 27260
rect 320 27020 380 27080
rect 11820 27020 11880 27080
rect 320 26840 380 26900
rect 1030 26840 1090 26900
rect 1660 26840 1720 26900
rect 2290 26840 2350 26900
rect 2920 26840 2980 26900
rect 3550 26840 3610 26900
rect 4180 26840 4240 26900
rect 4810 26840 4870 26900
rect 5440 26840 5500 26900
rect 6070 26840 6130 26900
rect 6700 26840 6760 26900
rect 7330 26840 7390 26900
rect 7960 26840 8020 26900
rect 8590 26840 8650 26900
rect 9220 26840 9280 26900
rect 9850 26840 9910 26900
rect 10480 26840 10540 26900
rect 11110 26840 11170 26900
rect 11820 26840 11880 26900
rect 320 26660 380 26720
rect 1030 26660 1090 26720
rect 1660 26660 1720 26720
rect 2290 26660 2350 26720
rect 2920 26660 2980 26720
rect 3550 26660 3610 26720
rect 4180 26660 4240 26720
rect 4810 26660 4870 26720
rect 5440 26660 5500 26720
rect 6070 26660 6130 26720
rect 6700 26660 6760 26720
rect 7330 26660 7390 26720
rect 7960 26660 8020 26720
rect 8590 26660 8650 26720
rect 9220 26660 9280 26720
rect 9850 26660 9910 26720
rect 10480 26660 10540 26720
rect 11110 26660 11170 26720
rect 11820 26660 11880 26720
rect 320 26480 380 26540
rect 1030 26480 1090 26540
rect 1660 26480 1720 26540
rect 2290 26480 2350 26540
rect 2920 26480 2980 26540
rect 3550 26480 3610 26540
rect 4180 26480 4240 26540
rect 4810 26480 4870 26540
rect 5440 26480 5500 26540
rect 6070 26480 6130 26540
rect 6700 26480 6760 26540
rect 7330 26480 7390 26540
rect 7960 26480 8020 26540
rect 8590 26480 8650 26540
rect 9220 26480 9280 26540
rect 9850 26480 9910 26540
rect 10480 26480 10540 26540
rect 11110 26480 11170 26540
rect 11820 26480 11880 26540
rect 320 26300 380 26360
rect 1030 26300 1090 26360
rect 1660 26300 1720 26360
rect 2290 26300 2350 26360
rect 2920 26300 2980 26360
rect 3550 26300 3610 26360
rect 4180 26300 4240 26360
rect 4810 26300 4870 26360
rect 5440 26300 5500 26360
rect 6070 26300 6130 26360
rect 6700 26300 6760 26360
rect 7330 26300 7390 26360
rect 7960 26300 8020 26360
rect 8590 26300 8650 26360
rect 9220 26300 9280 26360
rect 9850 26300 9910 26360
rect 10480 26300 10540 26360
rect 11110 26300 11170 26360
rect 11820 26300 11880 26360
rect 320 26120 380 26180
rect 1030 26120 1090 26180
rect 1660 26120 1720 26180
rect 2290 26120 2350 26180
rect 2920 26120 2980 26180
rect 3550 26120 3610 26180
rect 4180 26120 4240 26180
rect 4810 26120 4870 26180
rect 5440 26120 5500 26180
rect 6070 26120 6130 26180
rect 6700 26120 6760 26180
rect 7330 26120 7390 26180
rect 7960 26120 8020 26180
rect 8590 26120 8650 26180
rect 9220 26120 9280 26180
rect 9850 26120 9910 26180
rect 10480 26120 10540 26180
rect 11110 26120 11170 26180
rect 11820 26120 11880 26180
rect 320 25940 380 26000
rect 1030 25940 1090 26000
rect 1660 25940 1720 26000
rect 2290 25940 2350 26000
rect 2920 25940 2980 26000
rect 3550 25940 3610 26000
rect 4180 25940 4240 26000
rect 4810 25940 4870 26000
rect 5440 25940 5500 26000
rect 6070 25940 6130 26000
rect 6700 25940 6760 26000
rect 7330 25940 7390 26000
rect 7960 25940 8020 26000
rect 8590 25940 8650 26000
rect 9220 25940 9280 26000
rect 9850 25940 9910 26000
rect 10480 25940 10540 26000
rect 11110 25940 11170 26000
rect 11820 25940 11880 26000
rect 320 25760 380 25820
rect 1030 25760 1090 25820
rect 1660 25760 1720 25820
rect 2290 25760 2350 25820
rect 2920 25760 2980 25820
rect 3550 25760 3610 25820
rect 4180 25760 4240 25820
rect 4810 25760 4870 25820
rect 5440 25760 5500 25820
rect 6070 25760 6130 25820
rect 6700 25760 6760 25820
rect 7330 25760 7390 25820
rect 7960 25760 8020 25820
rect 8590 25760 8650 25820
rect 9220 25760 9280 25820
rect 9850 25760 9910 25820
rect 10480 25760 10540 25820
rect 11110 25760 11170 25820
rect 11820 25760 11880 25820
rect 320 25580 380 25640
rect 1030 25580 1090 25640
rect 1660 25580 1720 25640
rect 2290 25580 2350 25640
rect 2920 25580 2980 25640
rect 3550 25580 3610 25640
rect 4180 25580 4240 25640
rect 4810 25580 4870 25640
rect 5440 25580 5500 25640
rect 6070 25580 6130 25640
rect 6700 25580 6760 25640
rect 7330 25580 7390 25640
rect 7960 25580 8020 25640
rect 8590 25580 8650 25640
rect 9220 25580 9280 25640
rect 9850 25580 9910 25640
rect 10480 25580 10540 25640
rect 11110 25580 11170 25640
rect 11820 25580 11880 25640
rect 320 25400 380 25460
rect 1030 25400 1090 25460
rect 1660 25400 1720 25460
rect 2290 25400 2350 25460
rect 2920 25400 2980 25460
rect 3550 25400 3610 25460
rect 4180 25400 4240 25460
rect 4810 25400 4870 25460
rect 5440 25400 5500 25460
rect 6070 25400 6130 25460
rect 6700 25400 6760 25460
rect 7330 25400 7390 25460
rect 7960 25400 8020 25460
rect 8590 25400 8650 25460
rect 9220 25400 9280 25460
rect 9850 25400 9910 25460
rect 10480 25400 10540 25460
rect 11110 25400 11170 25460
rect 11820 25400 11880 25460
rect 320 25220 380 25280
rect 1030 25220 1090 25280
rect 1660 25220 1720 25280
rect 2290 25220 2350 25280
rect 2920 25220 2980 25280
rect 3550 25220 3610 25280
rect 4180 25220 4240 25280
rect 4810 25220 4870 25280
rect 5440 25220 5500 25280
rect 6070 25220 6130 25280
rect 6700 25220 6760 25280
rect 7330 25220 7390 25280
rect 7960 25220 8020 25280
rect 8590 25220 8650 25280
rect 9220 25220 9280 25280
rect 9850 25220 9910 25280
rect 10480 25220 10540 25280
rect 11110 25220 11170 25280
rect 11820 25220 11880 25280
rect 320 25040 380 25100
rect 1030 25040 1090 25100
rect 1660 25040 1720 25100
rect 2290 25040 2350 25100
rect 2920 25040 2980 25100
rect 3550 25040 3610 25100
rect 4180 25040 4240 25100
rect 4810 25040 4870 25100
rect 5440 25040 5500 25100
rect 6070 25040 6130 25100
rect 6700 25040 6760 25100
rect 7330 25040 7390 25100
rect 7960 25040 8020 25100
rect 8590 25040 8650 25100
rect 9220 25040 9280 25100
rect 9850 25040 9910 25100
rect 10480 25040 10540 25100
rect 11110 25040 11170 25100
rect 11820 25040 11880 25100
rect 320 24860 380 24920
rect 1030 24860 1090 24920
rect 1660 24860 1720 24920
rect 2290 24860 2350 24920
rect 2920 24860 2980 24920
rect 3550 24860 3610 24920
rect 4180 24860 4240 24920
rect 4810 24860 4870 24920
rect 5440 24860 5500 24920
rect 6070 24860 6130 24920
rect 6700 24860 6760 24920
rect 7330 24860 7390 24920
rect 7960 24860 8020 24920
rect 8590 24860 8650 24920
rect 9220 24860 9280 24920
rect 9850 24860 9910 24920
rect 10480 24860 10540 24920
rect 11110 24860 11170 24920
rect 11820 24860 11880 24920
rect 320 24680 380 24740
rect 1030 24680 1090 24740
rect 1660 24680 1720 24740
rect 2290 24680 2350 24740
rect 2920 24680 2980 24740
rect 3550 24680 3610 24740
rect 4180 24680 4240 24740
rect 4810 24680 4870 24740
rect 5440 24680 5500 24740
rect 6070 24680 6130 24740
rect 6700 24680 6760 24740
rect 7330 24680 7390 24740
rect 7960 24680 8020 24740
rect 8590 24680 8650 24740
rect 9220 24680 9280 24740
rect 9850 24680 9910 24740
rect 10480 24680 10540 24740
rect 11110 24680 11170 24740
rect 11820 24680 11880 24740
rect 320 24500 380 24560
rect 1030 24500 1090 24560
rect 1660 24500 1720 24560
rect 2290 24500 2350 24560
rect 2920 24500 2980 24560
rect 3550 24500 3610 24560
rect 4180 24500 4240 24560
rect 4810 24500 4870 24560
rect 5440 24500 5500 24560
rect 6070 24500 6130 24560
rect 6700 24500 6760 24560
rect 7330 24500 7390 24560
rect 7960 24500 8020 24560
rect 8590 24500 8650 24560
rect 9220 24500 9280 24560
rect 9850 24500 9910 24560
rect 10480 24500 10540 24560
rect 11110 24500 11170 24560
rect 11820 24500 11880 24560
rect 320 24320 380 24380
rect 1030 24320 1090 24380
rect 1660 24320 1720 24380
rect 2290 24320 2350 24380
rect 2920 24320 2980 24380
rect 3550 24320 3610 24380
rect 4180 24320 4240 24380
rect 4810 24320 4870 24380
rect 5440 24320 5500 24380
rect 6070 24320 6130 24380
rect 6700 24320 6760 24380
rect 7330 24320 7390 24380
rect 7960 24320 8020 24380
rect 8590 24320 8650 24380
rect 9220 24320 9280 24380
rect 9850 24320 9910 24380
rect 10480 24320 10540 24380
rect 11110 24320 11170 24380
rect 11820 24320 11880 24380
rect 320 24140 380 24200
rect 1030 24140 1090 24200
rect 1660 24140 1720 24200
rect 2290 24140 2350 24200
rect 2920 24140 2980 24200
rect 3550 24140 3610 24200
rect 4180 24140 4240 24200
rect 4810 24140 4870 24200
rect 5440 24140 5500 24200
rect 6070 24140 6130 24200
rect 6700 24140 6760 24200
rect 7330 24140 7390 24200
rect 7960 24140 8020 24200
rect 8590 24140 8650 24200
rect 9220 24140 9280 24200
rect 9850 24140 9910 24200
rect 10480 24140 10540 24200
rect 11110 24140 11170 24200
rect 11820 24140 11880 24200
rect 320 23960 380 24020
rect 1030 23960 1090 24020
rect 1660 23960 1720 24020
rect 2290 23960 2350 24020
rect 2920 23960 2980 24020
rect 3550 23960 3610 24020
rect 4180 23960 4240 24020
rect 4810 23960 4870 24020
rect 5440 23960 5500 24020
rect 6070 23960 6130 24020
rect 6700 23960 6760 24020
rect 7330 23960 7390 24020
rect 7960 23960 8020 24020
rect 8590 23960 8650 24020
rect 9220 23960 9280 24020
rect 9850 23960 9910 24020
rect 10480 23960 10540 24020
rect 11110 23960 11170 24020
rect 11820 23960 11880 24020
rect 320 23780 380 23840
rect 1030 23780 1090 23840
rect 1660 23780 1720 23840
rect 2290 23780 2350 23840
rect 2920 23780 2980 23840
rect 3550 23780 3610 23840
rect 4180 23780 4240 23840
rect 4810 23780 4870 23840
rect 5440 23780 5500 23840
rect 6070 23780 6130 23840
rect 6700 23780 6760 23840
rect 7330 23780 7390 23840
rect 7960 23780 8020 23840
rect 8590 23780 8650 23840
rect 9220 23780 9280 23840
rect 9850 23780 9910 23840
rect 10480 23780 10540 23840
rect 11110 23780 11170 23840
rect 11820 23780 11880 23840
rect 320 23600 380 23660
rect 1030 23600 1090 23660
rect 1660 23600 1720 23660
rect 2290 23600 2350 23660
rect 2920 23600 2980 23660
rect 3550 23600 3610 23660
rect 4180 23600 4240 23660
rect 4810 23600 4870 23660
rect 5440 23600 5500 23660
rect 6070 23600 6130 23660
rect 6700 23600 6760 23660
rect 7330 23600 7390 23660
rect 7960 23600 8020 23660
rect 8590 23600 8650 23660
rect 9220 23600 9280 23660
rect 9850 23600 9910 23660
rect 10480 23600 10540 23660
rect 11110 23600 11170 23660
rect 11820 23600 11880 23660
rect 320 23420 380 23480
rect 1030 23420 1090 23480
rect 1660 23420 1720 23480
rect 2290 23420 2350 23480
rect 2920 23420 2980 23480
rect 3550 23420 3610 23480
rect 4180 23420 4240 23480
rect 4810 23420 4870 23480
rect 5440 23420 5500 23480
rect 6070 23420 6130 23480
rect 6700 23420 6760 23480
rect 7330 23420 7390 23480
rect 7960 23420 8020 23480
rect 8590 23420 8650 23480
rect 9220 23420 9280 23480
rect 9850 23420 9910 23480
rect 10480 23420 10540 23480
rect 11110 23420 11170 23480
rect 11820 23420 11880 23480
rect 320 23240 380 23300
rect 1030 23240 1090 23300
rect 1660 23240 1720 23300
rect 2290 23240 2350 23300
rect 2920 23240 2980 23300
rect 3550 23240 3610 23300
rect 4180 23240 4240 23300
rect 4810 23240 4870 23300
rect 5440 23240 5500 23300
rect 6070 23240 6130 23300
rect 6700 23240 6760 23300
rect 7330 23240 7390 23300
rect 7960 23240 8020 23300
rect 8590 23240 8650 23300
rect 9220 23240 9280 23300
rect 9850 23240 9910 23300
rect 10480 23240 10540 23300
rect 11110 23240 11170 23300
rect 11820 23240 11880 23300
rect 320 23060 380 23120
rect 1030 23060 1090 23120
rect 1660 23060 1720 23120
rect 2290 23060 2350 23120
rect 2920 23060 2980 23120
rect 3550 23060 3610 23120
rect 4180 23060 4240 23120
rect 4810 23060 4870 23120
rect 5440 23060 5500 23120
rect 6070 23060 6130 23120
rect 6700 23060 6760 23120
rect 7330 23060 7390 23120
rect 7960 23060 8020 23120
rect 8590 23060 8650 23120
rect 9220 23060 9280 23120
rect 9850 23060 9910 23120
rect 10480 23060 10540 23120
rect 11110 23060 11170 23120
rect 11820 23060 11880 23120
rect 320 22880 380 22940
rect 1030 22880 1090 22940
rect 1660 22880 1720 22940
rect 2290 22880 2350 22940
rect 2920 22880 2980 22940
rect 3550 22880 3610 22940
rect 4180 22880 4240 22940
rect 4810 22880 4870 22940
rect 5440 22880 5500 22940
rect 6070 22880 6130 22940
rect 6700 22880 6760 22940
rect 7330 22880 7390 22940
rect 7960 22880 8020 22940
rect 8590 22880 8650 22940
rect 9220 22880 9280 22940
rect 9850 22880 9910 22940
rect 10480 22880 10540 22940
rect 11110 22880 11170 22940
rect 11820 22880 11880 22940
rect 320 22700 380 22760
rect 1030 22700 1090 22760
rect 1660 22700 1720 22760
rect 2290 22700 2350 22760
rect 2920 22700 2980 22760
rect 3550 22700 3610 22760
rect 4180 22700 4240 22760
rect 4810 22700 4870 22760
rect 5440 22700 5500 22760
rect 6070 22700 6130 22760
rect 6700 22700 6760 22760
rect 7330 22700 7390 22760
rect 7960 22700 8020 22760
rect 8590 22700 8650 22760
rect 9220 22700 9280 22760
rect 9850 22700 9910 22760
rect 10480 22700 10540 22760
rect 11110 22700 11170 22760
rect 11820 22700 11880 22760
rect 320 22520 380 22580
rect 1030 22520 1090 22580
rect 1660 22520 1720 22580
rect 2290 22520 2350 22580
rect 2920 22520 2980 22580
rect 3550 22520 3610 22580
rect 4180 22520 4240 22580
rect 4810 22520 4870 22580
rect 5440 22520 5500 22580
rect 6070 22520 6130 22580
rect 6700 22520 6760 22580
rect 7330 22520 7390 22580
rect 7960 22520 8020 22580
rect 8590 22520 8650 22580
rect 9220 22520 9280 22580
rect 9850 22520 9910 22580
rect 10480 22520 10540 22580
rect 11110 22520 11170 22580
rect 11820 22520 11880 22580
rect 320 22340 380 22400
rect 1030 22340 1090 22400
rect 1660 22340 1720 22400
rect 2290 22340 2350 22400
rect 2920 22340 2980 22400
rect 3550 22340 3610 22400
rect 4180 22340 4240 22400
rect 4810 22340 4870 22400
rect 5440 22340 5500 22400
rect 6070 22340 6130 22400
rect 6700 22340 6760 22400
rect 7330 22340 7390 22400
rect 7960 22340 8020 22400
rect 8590 22340 8650 22400
rect 9220 22340 9280 22400
rect 9850 22340 9910 22400
rect 10480 22340 10540 22400
rect 11110 22340 11170 22400
rect 11820 22340 11880 22400
rect 320 22160 380 22220
rect 1030 22160 1090 22220
rect 1660 22160 1720 22220
rect 2290 22160 2350 22220
rect 2920 22160 2980 22220
rect 3550 22160 3610 22220
rect 4180 22160 4240 22220
rect 4810 22160 4870 22220
rect 5440 22160 5500 22220
rect 6070 22160 6130 22220
rect 6700 22160 6760 22220
rect 7330 22160 7390 22220
rect 7960 22160 8020 22220
rect 8590 22160 8650 22220
rect 9220 22160 9280 22220
rect 9850 22160 9910 22220
rect 10480 22160 10540 22220
rect 11110 22160 11170 22220
rect 11820 22160 11880 22220
rect 320 21980 380 22040
rect 1030 21980 1090 22040
rect 1660 21980 1720 22040
rect 2290 21980 2350 22040
rect 2920 21980 2980 22040
rect 3550 21980 3610 22040
rect 4180 21980 4240 22040
rect 4810 21980 4870 22040
rect 5440 21980 5500 22040
rect 6070 21980 6130 22040
rect 6700 21980 6760 22040
rect 7330 21980 7390 22040
rect 7960 21980 8020 22040
rect 8590 21980 8650 22040
rect 9220 21980 9280 22040
rect 9850 21980 9910 22040
rect 10480 21980 10540 22040
rect 11110 21980 11170 22040
rect 11820 21980 11880 22040
rect 320 21800 380 21860
rect 1030 21800 1090 21860
rect 1660 21800 1720 21860
rect 2290 21800 2350 21860
rect 2920 21800 2980 21860
rect 3550 21800 3610 21860
rect 4180 21800 4240 21860
rect 4810 21800 4870 21860
rect 5440 21800 5500 21860
rect 6070 21800 6130 21860
rect 6700 21800 6760 21860
rect 7330 21800 7390 21860
rect 7960 21800 8020 21860
rect 8590 21800 8650 21860
rect 9220 21800 9280 21860
rect 9850 21800 9910 21860
rect 10480 21800 10540 21860
rect 11110 21800 11170 21860
rect 11820 21800 11880 21860
rect 320 21620 380 21680
rect 11820 21620 11880 21680
rect 320 21440 380 21500
rect 11820 21440 11880 21500
rect 320 21260 380 21320
rect 11820 21260 11880 21320
rect 320 21080 380 21140
rect 11820 21080 11880 21140
rect 320 20900 380 20960
rect 11820 20900 11880 20960
rect 660 20790 720 20850
rect 780 20790 840 20850
rect 900 20790 960 20850
rect 1020 20790 1080 20850
rect 1140 20790 1200 20850
rect 1260 20790 1320 20850
rect 1380 20790 1440 20850
rect 1500 20790 1560 20850
rect 1620 20790 1680 20850
rect 1740 20790 1800 20850
rect 1860 20790 1920 20850
rect 1980 20790 2040 20850
rect 2100 20790 2160 20850
rect 2220 20790 2280 20850
rect 2340 20790 2400 20850
rect 2460 20790 2520 20850
rect 2580 20790 2640 20850
rect 2700 20790 2760 20850
rect 2820 20790 2880 20850
rect 2940 20790 3000 20850
rect 3060 20790 3120 20850
rect 3180 20790 3240 20850
rect 3300 20790 3360 20850
rect 3420 20790 3480 20850
rect 3540 20790 3600 20850
rect 3660 20790 3720 20850
rect 3780 20790 3840 20850
rect 3900 20790 3960 20850
rect 4020 20790 4080 20850
rect 4140 20790 4200 20850
rect 4260 20790 4320 20850
rect 4380 20790 4440 20850
rect 4500 20790 4560 20850
rect 4620 20790 4680 20850
rect 4740 20790 4800 20850
rect 4860 20790 4920 20850
rect 4980 20790 5040 20850
rect 5100 20790 5160 20850
rect 5220 20790 5280 20850
rect 5340 20790 5400 20850
rect 5460 20790 5520 20850
rect 5580 20790 5640 20850
rect 5700 20790 5760 20850
rect 5820 20790 5880 20850
rect 5940 20790 6000 20850
rect 6060 20790 6120 20850
rect 6180 20790 6240 20850
rect 6300 20790 6360 20850
rect 6420 20790 6480 20850
rect 6540 20790 6600 20850
rect 6660 20790 6720 20850
rect 6780 20790 6840 20850
rect 6900 20790 6960 20850
rect 7020 20790 7080 20850
rect 7140 20790 7200 20850
rect 7260 20790 7320 20850
rect 7380 20790 7440 20850
rect 7500 20790 7560 20850
rect 7620 20790 7680 20850
rect 7740 20790 7800 20850
rect 7860 20790 7920 20850
rect 7980 20790 8040 20850
rect 8100 20790 8160 20850
rect 8220 20790 8280 20850
rect 8340 20790 8400 20850
rect 8460 20790 8520 20850
rect 8580 20790 8640 20850
rect 8700 20790 8760 20850
rect 8820 20790 8880 20850
rect 8940 20790 9000 20850
rect 9060 20790 9120 20850
rect 9180 20790 9240 20850
rect 9300 20790 9360 20850
rect 9420 20790 9480 20850
rect 9540 20790 9600 20850
rect 9660 20790 9720 20850
rect 9780 20790 9840 20850
rect 9900 20790 9960 20850
rect 10020 20790 10080 20850
rect 10140 20790 10200 20850
rect 10260 20790 10320 20850
rect 10380 20790 10440 20850
rect 10500 20790 10560 20850
rect 10620 20790 10680 20850
rect 10740 20790 10800 20850
rect 10860 20790 10920 20850
rect 10980 20790 11040 20850
rect 11100 20790 11160 20850
rect 11220 20790 11280 20850
rect 11340 20790 11400 20850
rect 11460 20790 11520 20850
rect 320 20720 380 20780
rect 660 20670 720 20730
rect 780 20670 840 20730
rect 900 20670 960 20730
rect 1020 20670 1080 20730
rect 1140 20670 1200 20730
rect 1260 20670 1320 20730
rect 1380 20670 1440 20730
rect 1500 20670 1560 20730
rect 1620 20670 1680 20730
rect 1740 20670 1800 20730
rect 1860 20670 1920 20730
rect 1980 20670 2040 20730
rect 2100 20670 2160 20730
rect 2220 20670 2280 20730
rect 2340 20670 2400 20730
rect 2460 20670 2520 20730
rect 2580 20670 2640 20730
rect 2700 20670 2760 20730
rect 2820 20670 2880 20730
rect 2940 20670 3000 20730
rect 3060 20670 3120 20730
rect 3180 20670 3240 20730
rect 3300 20670 3360 20730
rect 3420 20670 3480 20730
rect 3540 20670 3600 20730
rect 3660 20670 3720 20730
rect 3780 20670 3840 20730
rect 3900 20670 3960 20730
rect 4020 20670 4080 20730
rect 4140 20670 4200 20730
rect 4260 20670 4320 20730
rect 4380 20670 4440 20730
rect 4500 20670 4560 20730
rect 4620 20670 4680 20730
rect 4740 20670 4800 20730
rect 4860 20670 4920 20730
rect 4980 20670 5040 20730
rect 5100 20670 5160 20730
rect 5220 20670 5280 20730
rect 5340 20670 5400 20730
rect 5460 20670 5520 20730
rect 5580 20670 5640 20730
rect 5700 20670 5760 20730
rect 5820 20670 5880 20730
rect 5940 20670 6000 20730
rect 6060 20670 6120 20730
rect 6180 20670 6240 20730
rect 6300 20670 6360 20730
rect 6420 20670 6480 20730
rect 6540 20670 6600 20730
rect 6660 20670 6720 20730
rect 6780 20670 6840 20730
rect 6900 20670 6960 20730
rect 7020 20670 7080 20730
rect 7140 20670 7200 20730
rect 7260 20670 7320 20730
rect 7380 20670 7440 20730
rect 7500 20670 7560 20730
rect 7620 20670 7680 20730
rect 7740 20670 7800 20730
rect 7860 20670 7920 20730
rect 7980 20670 8040 20730
rect 8100 20670 8160 20730
rect 8220 20670 8280 20730
rect 8340 20670 8400 20730
rect 8460 20670 8520 20730
rect 8580 20670 8640 20730
rect 8700 20670 8760 20730
rect 8820 20670 8880 20730
rect 8940 20670 9000 20730
rect 9060 20670 9120 20730
rect 9180 20670 9240 20730
rect 9300 20670 9360 20730
rect 9420 20670 9480 20730
rect 9540 20670 9600 20730
rect 9660 20670 9720 20730
rect 9780 20670 9840 20730
rect 9900 20670 9960 20730
rect 10020 20670 10080 20730
rect 10140 20670 10200 20730
rect 10260 20670 10320 20730
rect 10380 20670 10440 20730
rect 10500 20670 10560 20730
rect 10620 20670 10680 20730
rect 10740 20670 10800 20730
rect 10860 20670 10920 20730
rect 10980 20670 11040 20730
rect 11100 20670 11160 20730
rect 11220 20670 11280 20730
rect 11340 20670 11400 20730
rect 11460 20670 11520 20730
rect 11820 20720 11880 20780
rect 320 20540 380 20600
rect 660 20550 720 20610
rect 780 20550 840 20610
rect 900 20550 960 20610
rect 1020 20550 1080 20610
rect 1140 20550 1200 20610
rect 1260 20550 1320 20610
rect 1380 20550 1440 20610
rect 1500 20550 1560 20610
rect 1620 20550 1680 20610
rect 1740 20550 1800 20610
rect 1860 20550 1920 20610
rect 1980 20550 2040 20610
rect 2100 20550 2160 20610
rect 2220 20550 2280 20610
rect 2340 20550 2400 20610
rect 2460 20550 2520 20610
rect 2580 20550 2640 20610
rect 2700 20550 2760 20610
rect 2820 20550 2880 20610
rect 2940 20550 3000 20610
rect 3060 20550 3120 20610
rect 3180 20550 3240 20610
rect 3300 20550 3360 20610
rect 3420 20550 3480 20610
rect 3540 20550 3600 20610
rect 3660 20550 3720 20610
rect 3780 20550 3840 20610
rect 3900 20550 3960 20610
rect 4020 20550 4080 20610
rect 4140 20550 4200 20610
rect 4260 20550 4320 20610
rect 4380 20550 4440 20610
rect 4500 20550 4560 20610
rect 4620 20550 4680 20610
rect 4740 20550 4800 20610
rect 4860 20550 4920 20610
rect 4980 20550 5040 20610
rect 5100 20550 5160 20610
rect 5220 20550 5280 20610
rect 5340 20550 5400 20610
rect 5460 20550 5520 20610
rect 5580 20550 5640 20610
rect 5700 20550 5760 20610
rect 5820 20550 5880 20610
rect 5940 20550 6000 20610
rect 6060 20550 6120 20610
rect 6180 20550 6240 20610
rect 6300 20550 6360 20610
rect 6420 20550 6480 20610
rect 6540 20550 6600 20610
rect 6660 20550 6720 20610
rect 6780 20550 6840 20610
rect 6900 20550 6960 20610
rect 7020 20550 7080 20610
rect 7140 20550 7200 20610
rect 7260 20550 7320 20610
rect 7380 20550 7440 20610
rect 7500 20550 7560 20610
rect 7620 20550 7680 20610
rect 7740 20550 7800 20610
rect 7860 20550 7920 20610
rect 7980 20550 8040 20610
rect 8100 20550 8160 20610
rect 8220 20550 8280 20610
rect 8340 20550 8400 20610
rect 8460 20550 8520 20610
rect 8580 20550 8640 20610
rect 8700 20550 8760 20610
rect 8820 20550 8880 20610
rect 8940 20550 9000 20610
rect 9060 20550 9120 20610
rect 9180 20550 9240 20610
rect 9300 20550 9360 20610
rect 9420 20550 9480 20610
rect 9540 20550 9600 20610
rect 9660 20550 9720 20610
rect 9780 20550 9840 20610
rect 9900 20550 9960 20610
rect 10020 20550 10080 20610
rect 10140 20550 10200 20610
rect 10260 20550 10320 20610
rect 10380 20550 10440 20610
rect 10500 20550 10560 20610
rect 10620 20550 10680 20610
rect 10740 20550 10800 20610
rect 10860 20550 10920 20610
rect 10980 20550 11040 20610
rect 11100 20550 11160 20610
rect 11220 20550 11280 20610
rect 11340 20550 11400 20610
rect 11460 20550 11520 20610
rect 11820 20540 11880 20600
rect 890 19765 950 19825
rect 1070 19765 1130 19825
rect 1250 19765 1310 19825
rect 1430 19765 1490 19825
rect 1610 19765 1670 19825
rect 1790 19765 1850 19825
rect 1970 19765 2030 19825
rect 2150 19765 2210 19825
rect 2330 19765 2390 19825
rect 2510 19765 2570 19825
rect 2690 19765 2750 19825
rect 2870 19765 2930 19825
rect 3050 19765 3110 19825
rect 3230 19765 3290 19825
rect 3410 19765 3470 19825
rect 3590 19765 3650 19825
rect 3770 19765 3830 19825
rect 3950 19765 4010 19825
rect 4130 19765 4190 19825
rect 4310 19765 4370 19825
rect 4490 19765 4550 19825
rect 4670 19765 4730 19825
rect 4850 19765 4910 19825
rect 5030 19765 5090 19825
rect 5210 19765 5270 19825
rect 5390 19765 5450 19825
rect 5570 19765 5630 19825
rect 5750 19765 5810 19825
rect 5930 19765 5990 19825
rect 6110 19765 6170 19825
rect 6290 19765 6350 19825
rect 6470 19765 6530 19825
rect 6650 19765 6710 19825
rect 6830 19765 6890 19825
rect 7010 19765 7070 19825
rect 7190 19765 7250 19825
rect 7370 19765 7430 19825
rect 7550 19765 7610 19825
rect 7730 19765 7790 19825
rect 7910 19765 7970 19825
rect 8090 19765 8150 19825
rect 8270 19765 8330 19825
rect 8450 19765 8510 19825
rect 8630 19765 8690 19825
rect 8810 19765 8870 19825
rect 8990 19765 9050 19825
rect 9170 19765 9230 19825
rect 9350 19765 9410 19825
rect 9530 19765 9590 19825
rect 9710 19765 9770 19825
rect 9890 19765 9950 19825
rect 10070 19765 10130 19825
rect 10250 19765 10310 19825
rect 10430 19765 10490 19825
rect 10610 19765 10670 19825
rect 10790 19765 10850 19825
rect 10970 19765 11030 19825
rect 11150 19765 11210 19825
rect 11330 19765 11390 19825
rect 11510 19765 11570 19825
rect 11690 19765 11750 19825
rect 11870 19765 11930 19825
rect 890 19585 950 19645
rect 1070 19585 1130 19645
rect 1250 19585 1310 19645
rect 1430 19585 1490 19645
rect 1610 19585 1670 19645
rect 1790 19585 1850 19645
rect 1970 19585 2030 19645
rect 2150 19585 2210 19645
rect 2330 19585 2390 19645
rect 2510 19585 2570 19645
rect 2690 19585 2750 19645
rect 2870 19585 2930 19645
rect 3050 19585 3110 19645
rect 3230 19585 3290 19645
rect 3410 19585 3470 19645
rect 3590 19585 3650 19645
rect 3770 19585 3830 19645
rect 3950 19585 4010 19645
rect 4130 19585 4190 19645
rect 4310 19585 4370 19645
rect 4490 19585 4550 19645
rect 4670 19585 4730 19645
rect 4850 19585 4910 19645
rect 5030 19585 5090 19645
rect 5210 19585 5270 19645
rect 5390 19585 5450 19645
rect 5570 19585 5630 19645
rect 5750 19585 5810 19645
rect 5930 19585 5990 19645
rect 6110 19585 6170 19645
rect 6290 19585 6350 19645
rect 6470 19585 6530 19645
rect 6650 19585 6710 19645
rect 6830 19585 6890 19645
rect 7010 19585 7070 19645
rect 7190 19585 7250 19645
rect 7370 19585 7430 19645
rect 7550 19585 7610 19645
rect 7730 19585 7790 19645
rect 7910 19585 7970 19645
rect 8090 19585 8150 19645
rect 8270 19585 8330 19645
rect 8450 19585 8510 19645
rect 8630 19585 8690 19645
rect 8810 19585 8870 19645
rect 8990 19585 9050 19645
rect 9170 19585 9230 19645
rect 9350 19585 9410 19645
rect 9530 19585 9590 19645
rect 9710 19585 9770 19645
rect 9890 19585 9950 19645
rect 10070 19585 10130 19645
rect 10250 19585 10310 19645
rect 10430 19585 10490 19645
rect 10610 19585 10670 19645
rect 10790 19585 10850 19645
rect 10970 19585 11030 19645
rect 11150 19585 11210 19645
rect 11330 19585 11390 19645
rect 11510 19585 11570 19645
rect 11690 19585 11750 19645
rect 11870 19585 11930 19645
rect 890 19405 950 19465
rect 1070 19405 1130 19465
rect 1250 19405 1310 19465
rect 1430 19405 1490 19465
rect 1610 19405 1670 19465
rect 1790 19405 1850 19465
rect 1970 19405 2030 19465
rect 2150 19405 2210 19465
rect 2330 19405 2390 19465
rect 2510 19405 2570 19465
rect 2690 19405 2750 19465
rect 2870 19405 2930 19465
rect 3050 19405 3110 19465
rect 3230 19405 3290 19465
rect 3410 19405 3470 19465
rect 3590 19405 3650 19465
rect 3770 19405 3830 19465
rect 3950 19405 4010 19465
rect 4130 19405 4190 19465
rect 4310 19405 4370 19465
rect 4490 19405 4550 19465
rect 4670 19405 4730 19465
rect 4850 19405 4910 19465
rect 5030 19405 5090 19465
rect 5210 19405 5270 19465
rect 5390 19405 5450 19465
rect 5570 19405 5630 19465
rect 5750 19405 5810 19465
rect 5930 19405 5990 19465
rect 6110 19405 6170 19465
rect 6290 19405 6350 19465
rect 6470 19405 6530 19465
rect 6650 19405 6710 19465
rect 6830 19405 6890 19465
rect 7010 19405 7070 19465
rect 7190 19405 7250 19465
rect 7370 19405 7430 19465
rect 7550 19405 7610 19465
rect 7730 19405 7790 19465
rect 7910 19405 7970 19465
rect 8090 19405 8150 19465
rect 8270 19405 8330 19465
rect 8450 19405 8510 19465
rect 8630 19405 8690 19465
rect 8810 19405 8870 19465
rect 8990 19405 9050 19465
rect 9170 19405 9230 19465
rect 9350 19405 9410 19465
rect 9530 19405 9590 19465
rect 9710 19405 9770 19465
rect 9890 19405 9950 19465
rect 10070 19405 10130 19465
rect 10250 19405 10310 19465
rect 10430 19405 10490 19465
rect 10610 19405 10670 19465
rect 10790 19405 10850 19465
rect 10970 19405 11030 19465
rect 11150 19405 11210 19465
rect 11330 19405 11390 19465
rect 11510 19405 11570 19465
rect 11690 19405 11750 19465
rect 11870 19405 11930 19465
rect 890 19225 950 19285
rect 1070 19225 1130 19285
rect 1250 19225 1310 19285
rect 1430 19225 1490 19285
rect 1610 19225 1670 19285
rect 1790 19225 1850 19285
rect 1970 19225 2030 19285
rect 2150 19225 2210 19285
rect 2330 19225 2390 19285
rect 2510 19225 2570 19285
rect 2690 19225 2750 19285
rect 2870 19225 2930 19285
rect 3050 19225 3110 19285
rect 3230 19225 3290 19285
rect 3410 19225 3470 19285
rect 3590 19225 3650 19285
rect 3770 19225 3830 19285
rect 3950 19225 4010 19285
rect 4130 19225 4190 19285
rect 4310 19225 4370 19285
rect 4490 19225 4550 19285
rect 4670 19225 4730 19285
rect 4850 19225 4910 19285
rect 5030 19225 5090 19285
rect 5210 19225 5270 19285
rect 5390 19225 5450 19285
rect 5570 19225 5630 19285
rect 5750 19225 5810 19285
rect 5930 19225 5990 19285
rect 6110 19225 6170 19285
rect 6290 19225 6350 19285
rect 6470 19225 6530 19285
rect 6650 19225 6710 19285
rect 6830 19225 6890 19285
rect 7010 19225 7070 19285
rect 7190 19225 7250 19285
rect 7370 19225 7430 19285
rect 7550 19225 7610 19285
rect 7730 19225 7790 19285
rect 7910 19225 7970 19285
rect 8090 19225 8150 19285
rect 8270 19225 8330 19285
rect 8450 19225 8510 19285
rect 8630 19225 8690 19285
rect 8810 19225 8870 19285
rect 8990 19225 9050 19285
rect 9170 19225 9230 19285
rect 9350 19225 9410 19285
rect 9530 19225 9590 19285
rect 9710 19225 9770 19285
rect 9890 19225 9950 19285
rect 10070 19225 10130 19285
rect 10250 19225 10310 19285
rect 10430 19225 10490 19285
rect 10610 19225 10670 19285
rect 10790 19225 10850 19285
rect 10970 19225 11030 19285
rect 11150 19225 11210 19285
rect 11330 19225 11390 19285
rect 11510 19225 11570 19285
rect 11690 19225 11750 19285
rect 11870 19225 11930 19285
rect 890 19045 950 19105
rect 1070 19045 1130 19105
rect 1250 19045 1310 19105
rect 1430 19045 1490 19105
rect 1610 19045 1670 19105
rect 1790 19045 1850 19105
rect 1970 19045 2030 19105
rect 2150 19045 2210 19105
rect 2330 19045 2390 19105
rect 2510 19045 2570 19105
rect 2690 19045 2750 19105
rect 2870 19045 2930 19105
rect 3050 19045 3110 19105
rect 3230 19045 3290 19105
rect 3410 19045 3470 19105
rect 3590 19045 3650 19105
rect 3770 19045 3830 19105
rect 3950 19045 4010 19105
rect 4130 19045 4190 19105
rect 4310 19045 4370 19105
rect 4490 19045 4550 19105
rect 4670 19045 4730 19105
rect 4850 19045 4910 19105
rect 5030 19045 5090 19105
rect 5210 19045 5270 19105
rect 5390 19045 5450 19105
rect 5570 19045 5630 19105
rect 5750 19045 5810 19105
rect 5930 19045 5990 19105
rect 6110 19045 6170 19105
rect 6290 19045 6350 19105
rect 6470 19045 6530 19105
rect 6650 19045 6710 19105
rect 6830 19045 6890 19105
rect 7010 19045 7070 19105
rect 7190 19045 7250 19105
rect 7370 19045 7430 19105
rect 7550 19045 7610 19105
rect 7730 19045 7790 19105
rect 7910 19045 7970 19105
rect 8090 19045 8150 19105
rect 8270 19045 8330 19105
rect 8450 19045 8510 19105
rect 8630 19045 8690 19105
rect 8810 19045 8870 19105
rect 8990 19045 9050 19105
rect 9170 19045 9230 19105
rect 9350 19045 9410 19105
rect 9530 19045 9590 19105
rect 9710 19045 9770 19105
rect 9890 19045 9950 19105
rect 10070 19045 10130 19105
rect 10250 19045 10310 19105
rect 10430 19045 10490 19105
rect 10610 19045 10670 19105
rect 10790 19045 10850 19105
rect 10970 19045 11030 19105
rect 11150 19045 11210 19105
rect 11330 19045 11390 19105
rect 11510 19045 11570 19105
rect 11690 19045 11750 19105
rect 11870 19045 11930 19105
rect 350 18295 410 18355
rect 530 18295 590 18355
rect 710 18295 770 18355
rect 890 18295 950 18355
rect 1070 18295 1130 18355
rect 1250 18295 1310 18355
rect 1430 18295 1490 18355
rect 1610 18295 1670 18355
rect 1790 18295 1850 18355
rect 1970 18295 2030 18355
rect 2150 18295 2210 18355
rect 2330 18295 2390 18355
rect 2510 18295 2570 18355
rect 2690 18295 2750 18355
rect 2870 18295 2930 18355
rect 3050 18295 3110 18355
rect 3230 18295 3290 18355
rect 3410 18295 3470 18355
rect 3590 18295 3650 18355
rect 3770 18295 3830 18355
rect 3950 18295 4010 18355
rect 4130 18295 4190 18355
rect 4310 18295 4370 18355
rect 4490 18295 4550 18355
rect 4670 18295 4730 18355
rect 4850 18295 4910 18355
rect 5030 18295 5090 18355
rect 5210 18295 5270 18355
rect 5390 18295 5450 18355
rect 5570 18295 5630 18355
rect 5750 18295 5810 18355
rect 5930 18295 5990 18355
rect 6110 18295 6170 18355
rect 6290 18295 6350 18355
rect 6470 18295 6530 18355
rect 6650 18295 6710 18355
rect 6830 18295 6890 18355
rect 7010 18295 7070 18355
rect 7190 18295 7250 18355
rect 7370 18295 7430 18355
rect 7550 18295 7610 18355
rect 7730 18295 7790 18355
rect 7910 18295 7970 18355
rect 8090 18295 8150 18355
rect 8270 18295 8330 18355
rect 8450 18295 8510 18355
rect 8630 18295 8690 18355
rect 8810 18295 8870 18355
rect 8990 18295 9050 18355
rect 9170 18295 9230 18355
rect 9350 18295 9410 18355
rect 9530 18295 9590 18355
rect 9710 18295 9770 18355
rect 9890 18295 9950 18355
rect 10070 18295 10130 18355
rect 10250 18295 10310 18355
rect 10430 18295 10490 18355
rect 10610 18295 10670 18355
rect 10790 18295 10850 18355
rect 10970 18295 11030 18355
rect 11150 18295 11210 18355
rect 11330 18295 11390 18355
rect 350 18115 410 18175
rect 530 18115 590 18175
rect 710 18115 770 18175
rect 890 18115 950 18175
rect 1070 18115 1130 18175
rect 1250 18115 1310 18175
rect 1430 18115 1490 18175
rect 1610 18115 1670 18175
rect 1790 18115 1850 18175
rect 1970 18115 2030 18175
rect 2150 18115 2210 18175
rect 2330 18115 2390 18175
rect 2510 18115 2570 18175
rect 2690 18115 2750 18175
rect 2870 18115 2930 18175
rect 3050 18115 3110 18175
rect 3230 18115 3290 18175
rect 3410 18115 3470 18175
rect 3590 18115 3650 18175
rect 3770 18115 3830 18175
rect 3950 18115 4010 18175
rect 4130 18115 4190 18175
rect 4310 18115 4370 18175
rect 4490 18115 4550 18175
rect 4670 18115 4730 18175
rect 4850 18115 4910 18175
rect 5030 18115 5090 18175
rect 5210 18115 5270 18175
rect 5390 18115 5450 18175
rect 5570 18115 5630 18175
rect 5750 18115 5810 18175
rect 5930 18115 5990 18175
rect 6110 18115 6170 18175
rect 6290 18115 6350 18175
rect 6470 18115 6530 18175
rect 6650 18115 6710 18175
rect 6830 18115 6890 18175
rect 7010 18115 7070 18175
rect 7190 18115 7250 18175
rect 7370 18115 7430 18175
rect 7550 18115 7610 18175
rect 7730 18115 7790 18175
rect 7910 18115 7970 18175
rect 8090 18115 8150 18175
rect 8270 18115 8330 18175
rect 8450 18115 8510 18175
rect 8630 18115 8690 18175
rect 8810 18115 8870 18175
rect 8990 18115 9050 18175
rect 9170 18115 9230 18175
rect 9350 18115 9410 18175
rect 9530 18115 9590 18175
rect 9710 18115 9770 18175
rect 9890 18115 9950 18175
rect 10070 18115 10130 18175
rect 10250 18115 10310 18175
rect 10430 18115 10490 18175
rect 10610 18115 10670 18175
rect 10790 18115 10850 18175
rect 10970 18115 11030 18175
rect 11150 18115 11210 18175
rect 11330 18115 11390 18175
rect 350 17935 410 17995
rect 530 17935 590 17995
rect 710 17935 770 17995
rect 890 17935 950 17995
rect 1070 17935 1130 17995
rect 1250 17935 1310 17995
rect 1430 17935 1490 17995
rect 1610 17935 1670 17995
rect 1790 17935 1850 17995
rect 1970 17935 2030 17995
rect 2150 17935 2210 17995
rect 2330 17935 2390 17995
rect 2510 17935 2570 17995
rect 2690 17935 2750 17995
rect 2870 17935 2930 17995
rect 3050 17935 3110 17995
rect 3230 17935 3290 17995
rect 3410 17935 3470 17995
rect 3590 17935 3650 17995
rect 3770 17935 3830 17995
rect 3950 17935 4010 17995
rect 4130 17935 4190 17995
rect 4310 17935 4370 17995
rect 4490 17935 4550 17995
rect 4670 17935 4730 17995
rect 4850 17935 4910 17995
rect 5030 17935 5090 17995
rect 5210 17935 5270 17995
rect 5390 17935 5450 17995
rect 5570 17935 5630 17995
rect 5750 17935 5810 17995
rect 5930 17935 5990 17995
rect 6110 17935 6170 17995
rect 6290 17935 6350 17995
rect 6470 17935 6530 17995
rect 6650 17935 6710 17995
rect 6830 17935 6890 17995
rect 7010 17935 7070 17995
rect 7190 17935 7250 17995
rect 7370 17935 7430 17995
rect 7550 17935 7610 17995
rect 7730 17935 7790 17995
rect 7910 17935 7970 17995
rect 8090 17935 8150 17995
rect 8270 17935 8330 17995
rect 8450 17935 8510 17995
rect 8630 17935 8690 17995
rect 8810 17935 8870 17995
rect 8990 17935 9050 17995
rect 9170 17935 9230 17995
rect 9350 17935 9410 17995
rect 9530 17935 9590 17995
rect 9710 17935 9770 17995
rect 9890 17935 9950 17995
rect 10070 17935 10130 17995
rect 10250 17935 10310 17995
rect 10430 17935 10490 17995
rect 10610 17935 10670 17995
rect 10790 17935 10850 17995
rect 10970 17935 11030 17995
rect 11150 17935 11210 17995
rect 11330 17935 11390 17995
rect 350 17755 410 17815
rect 530 17755 590 17815
rect 710 17755 770 17815
rect 890 17755 950 17815
rect 1070 17755 1130 17815
rect 1250 17755 1310 17815
rect 1430 17755 1490 17815
rect 1610 17755 1670 17815
rect 1790 17755 1850 17815
rect 1970 17755 2030 17815
rect 2150 17755 2210 17815
rect 2330 17755 2390 17815
rect 2510 17755 2570 17815
rect 2690 17755 2750 17815
rect 2870 17755 2930 17815
rect 3050 17755 3110 17815
rect 3230 17755 3290 17815
rect 3410 17755 3470 17815
rect 3590 17755 3650 17815
rect 3770 17755 3830 17815
rect 3950 17755 4010 17815
rect 4130 17755 4190 17815
rect 4310 17755 4370 17815
rect 4490 17755 4550 17815
rect 4670 17755 4730 17815
rect 4850 17755 4910 17815
rect 5030 17755 5090 17815
rect 5210 17755 5270 17815
rect 5390 17755 5450 17815
rect 5570 17755 5630 17815
rect 5750 17755 5810 17815
rect 5930 17755 5990 17815
rect 6110 17755 6170 17815
rect 6290 17755 6350 17815
rect 6470 17755 6530 17815
rect 6650 17755 6710 17815
rect 6830 17755 6890 17815
rect 7010 17755 7070 17815
rect 7190 17755 7250 17815
rect 7370 17755 7430 17815
rect 7550 17755 7610 17815
rect 7730 17755 7790 17815
rect 7910 17755 7970 17815
rect 8090 17755 8150 17815
rect 8270 17755 8330 17815
rect 8450 17755 8510 17815
rect 8630 17755 8690 17815
rect 8810 17755 8870 17815
rect 8990 17755 9050 17815
rect 9170 17755 9230 17815
rect 9350 17755 9410 17815
rect 9530 17755 9590 17815
rect 9710 17755 9770 17815
rect 9890 17755 9950 17815
rect 10070 17755 10130 17815
rect 10250 17755 10310 17815
rect 10430 17755 10490 17815
rect 10610 17755 10670 17815
rect 10790 17755 10850 17815
rect 10970 17755 11030 17815
rect 11150 17755 11210 17815
rect 11330 17755 11390 17815
rect 350 17575 410 17635
rect 530 17575 590 17635
rect 710 17575 770 17635
rect 890 17575 950 17635
rect 1070 17575 1130 17635
rect 1250 17575 1310 17635
rect 1430 17575 1490 17635
rect 1610 17575 1670 17635
rect 1790 17575 1850 17635
rect 1970 17575 2030 17635
rect 2150 17575 2210 17635
rect 2330 17575 2390 17635
rect 2510 17575 2570 17635
rect 2690 17575 2750 17635
rect 2870 17575 2930 17635
rect 3050 17575 3110 17635
rect 3230 17575 3290 17635
rect 3410 17575 3470 17635
rect 3590 17575 3650 17635
rect 3770 17575 3830 17635
rect 3950 17575 4010 17635
rect 4130 17575 4190 17635
rect 4310 17575 4370 17635
rect 4490 17575 4550 17635
rect 4670 17575 4730 17635
rect 4850 17575 4910 17635
rect 5030 17575 5090 17635
rect 5210 17575 5270 17635
rect 5390 17575 5450 17635
rect 5570 17575 5630 17635
rect 5750 17575 5810 17635
rect 5930 17575 5990 17635
rect 6110 17575 6170 17635
rect 6290 17575 6350 17635
rect 6470 17575 6530 17635
rect 6650 17575 6710 17635
rect 6830 17575 6890 17635
rect 7010 17575 7070 17635
rect 7190 17575 7250 17635
rect 7370 17575 7430 17635
rect 7550 17575 7610 17635
rect 7730 17575 7790 17635
rect 7910 17575 7970 17635
rect 8090 17575 8150 17635
rect 8270 17575 8330 17635
rect 8450 17575 8510 17635
rect 8630 17575 8690 17635
rect 8810 17575 8870 17635
rect 8990 17575 9050 17635
rect 9170 17575 9230 17635
rect 9350 17575 9410 17635
rect 9530 17575 9590 17635
rect 9710 17575 9770 17635
rect 9890 17575 9950 17635
rect 10070 17575 10130 17635
rect 10250 17575 10310 17635
rect 10430 17575 10490 17635
rect 10610 17575 10670 17635
rect 10790 17575 10850 17635
rect 10970 17575 11030 17635
rect 11150 17575 11210 17635
rect 11330 17575 11390 17635
rect 320 16800 380 16860
rect 660 16790 720 16850
rect 780 16790 840 16850
rect 900 16790 960 16850
rect 1020 16790 1080 16850
rect 1140 16790 1200 16850
rect 1260 16790 1320 16850
rect 1380 16790 1440 16850
rect 1500 16790 1560 16850
rect 1620 16790 1680 16850
rect 1740 16790 1800 16850
rect 1860 16790 1920 16850
rect 1980 16790 2040 16850
rect 2100 16790 2160 16850
rect 2220 16790 2280 16850
rect 2340 16790 2400 16850
rect 2460 16790 2520 16850
rect 2580 16790 2640 16850
rect 2700 16790 2760 16850
rect 2820 16790 2880 16850
rect 2940 16790 3000 16850
rect 3060 16790 3120 16850
rect 3180 16790 3240 16850
rect 3300 16790 3360 16850
rect 3420 16790 3480 16850
rect 3540 16790 3600 16850
rect 3660 16790 3720 16850
rect 3780 16790 3840 16850
rect 3900 16790 3960 16850
rect 4020 16790 4080 16850
rect 4140 16790 4200 16850
rect 4260 16790 4320 16850
rect 4380 16790 4440 16850
rect 4500 16790 4560 16850
rect 4620 16790 4680 16850
rect 4740 16790 4800 16850
rect 4860 16790 4920 16850
rect 4980 16790 5040 16850
rect 5100 16790 5160 16850
rect 5220 16790 5280 16850
rect 5340 16790 5400 16850
rect 5460 16790 5520 16850
rect 5580 16790 5640 16850
rect 5700 16790 5760 16850
rect 5820 16790 5880 16850
rect 5940 16790 6000 16850
rect 6060 16790 6120 16850
rect 6180 16790 6240 16850
rect 6300 16790 6360 16850
rect 6420 16790 6480 16850
rect 6540 16790 6600 16850
rect 6660 16790 6720 16850
rect 6780 16790 6840 16850
rect 6900 16790 6960 16850
rect 7020 16790 7080 16850
rect 7140 16790 7200 16850
rect 7260 16790 7320 16850
rect 7380 16790 7440 16850
rect 7500 16790 7560 16850
rect 7620 16790 7680 16850
rect 7740 16790 7800 16850
rect 7860 16790 7920 16850
rect 7980 16790 8040 16850
rect 8100 16790 8160 16850
rect 8220 16790 8280 16850
rect 8340 16790 8400 16850
rect 8460 16790 8520 16850
rect 8580 16790 8640 16850
rect 8700 16790 8760 16850
rect 8820 16790 8880 16850
rect 8940 16790 9000 16850
rect 9060 16790 9120 16850
rect 9180 16790 9240 16850
rect 9300 16790 9360 16850
rect 9420 16790 9480 16850
rect 9540 16790 9600 16850
rect 9660 16790 9720 16850
rect 9780 16790 9840 16850
rect 9900 16790 9960 16850
rect 10020 16790 10080 16850
rect 10140 16790 10200 16850
rect 10260 16790 10320 16850
rect 10380 16790 10440 16850
rect 10500 16790 10560 16850
rect 10620 16790 10680 16850
rect 10740 16790 10800 16850
rect 10860 16790 10920 16850
rect 10980 16790 11040 16850
rect 11100 16790 11160 16850
rect 11220 16790 11280 16850
rect 11340 16790 11400 16850
rect 11820 16800 11880 16860
rect 320 16620 380 16680
rect 660 16670 720 16730
rect 780 16670 840 16730
rect 900 16670 960 16730
rect 1020 16670 1080 16730
rect 1140 16670 1200 16730
rect 1260 16670 1320 16730
rect 1380 16670 1440 16730
rect 1500 16670 1560 16730
rect 1620 16670 1680 16730
rect 1740 16670 1800 16730
rect 1860 16670 1920 16730
rect 1980 16670 2040 16730
rect 2100 16670 2160 16730
rect 2220 16670 2280 16730
rect 2340 16670 2400 16730
rect 2460 16670 2520 16730
rect 2580 16670 2640 16730
rect 2700 16670 2760 16730
rect 2820 16670 2880 16730
rect 2940 16670 3000 16730
rect 3060 16670 3120 16730
rect 3180 16670 3240 16730
rect 3300 16670 3360 16730
rect 3420 16670 3480 16730
rect 3540 16670 3600 16730
rect 3660 16670 3720 16730
rect 3780 16670 3840 16730
rect 3900 16670 3960 16730
rect 4020 16670 4080 16730
rect 4140 16670 4200 16730
rect 4260 16670 4320 16730
rect 4380 16670 4440 16730
rect 4500 16670 4560 16730
rect 4620 16670 4680 16730
rect 4740 16670 4800 16730
rect 4860 16670 4920 16730
rect 4980 16670 5040 16730
rect 5100 16670 5160 16730
rect 5220 16670 5280 16730
rect 5340 16670 5400 16730
rect 5460 16670 5520 16730
rect 5580 16670 5640 16730
rect 5700 16670 5760 16730
rect 5820 16670 5880 16730
rect 5940 16670 6000 16730
rect 6060 16670 6120 16730
rect 6180 16670 6240 16730
rect 6300 16670 6360 16730
rect 6420 16670 6480 16730
rect 6540 16670 6600 16730
rect 6660 16670 6720 16730
rect 6780 16670 6840 16730
rect 6900 16670 6960 16730
rect 7020 16670 7080 16730
rect 7140 16670 7200 16730
rect 7260 16670 7320 16730
rect 7380 16670 7440 16730
rect 7500 16670 7560 16730
rect 7620 16670 7680 16730
rect 7740 16670 7800 16730
rect 7860 16670 7920 16730
rect 7980 16670 8040 16730
rect 8100 16670 8160 16730
rect 8220 16670 8280 16730
rect 8340 16670 8400 16730
rect 8460 16670 8520 16730
rect 8580 16670 8640 16730
rect 8700 16670 8760 16730
rect 8820 16670 8880 16730
rect 8940 16670 9000 16730
rect 9060 16670 9120 16730
rect 9180 16670 9240 16730
rect 9300 16670 9360 16730
rect 9420 16670 9480 16730
rect 9540 16670 9600 16730
rect 9660 16670 9720 16730
rect 9780 16670 9840 16730
rect 9900 16670 9960 16730
rect 10020 16670 10080 16730
rect 10140 16670 10200 16730
rect 10260 16670 10320 16730
rect 10380 16670 10440 16730
rect 10500 16670 10560 16730
rect 10620 16670 10680 16730
rect 10740 16670 10800 16730
rect 10860 16670 10920 16730
rect 10980 16670 11040 16730
rect 11100 16670 11160 16730
rect 11220 16670 11280 16730
rect 11340 16670 11400 16730
rect 11820 16620 11880 16680
rect 660 16550 720 16610
rect 780 16550 840 16610
rect 900 16550 960 16610
rect 1020 16550 1080 16610
rect 1140 16550 1200 16610
rect 1260 16550 1320 16610
rect 1380 16550 1440 16610
rect 1500 16550 1560 16610
rect 1620 16550 1680 16610
rect 1740 16550 1800 16610
rect 1860 16550 1920 16610
rect 1980 16550 2040 16610
rect 2100 16550 2160 16610
rect 2220 16550 2280 16610
rect 2340 16550 2400 16610
rect 2460 16550 2520 16610
rect 2580 16550 2640 16610
rect 2700 16550 2760 16610
rect 2820 16550 2880 16610
rect 2940 16550 3000 16610
rect 3060 16550 3120 16610
rect 3180 16550 3240 16610
rect 3300 16550 3360 16610
rect 3420 16550 3480 16610
rect 3540 16550 3600 16610
rect 3660 16550 3720 16610
rect 3780 16550 3840 16610
rect 3900 16550 3960 16610
rect 4020 16550 4080 16610
rect 4140 16550 4200 16610
rect 4260 16550 4320 16610
rect 4380 16550 4440 16610
rect 4500 16550 4560 16610
rect 4620 16550 4680 16610
rect 4740 16550 4800 16610
rect 4860 16550 4920 16610
rect 4980 16550 5040 16610
rect 5100 16550 5160 16610
rect 5220 16550 5280 16610
rect 5340 16550 5400 16610
rect 5460 16550 5520 16610
rect 5580 16550 5640 16610
rect 5700 16550 5760 16610
rect 5820 16550 5880 16610
rect 5940 16550 6000 16610
rect 6060 16550 6120 16610
rect 6180 16550 6240 16610
rect 6300 16550 6360 16610
rect 6420 16550 6480 16610
rect 6540 16550 6600 16610
rect 6660 16550 6720 16610
rect 6780 16550 6840 16610
rect 6900 16550 6960 16610
rect 7020 16550 7080 16610
rect 7140 16550 7200 16610
rect 7260 16550 7320 16610
rect 7380 16550 7440 16610
rect 7500 16550 7560 16610
rect 7620 16550 7680 16610
rect 7740 16550 7800 16610
rect 7860 16550 7920 16610
rect 7980 16550 8040 16610
rect 8100 16550 8160 16610
rect 8220 16550 8280 16610
rect 8340 16550 8400 16610
rect 8460 16550 8520 16610
rect 8580 16550 8640 16610
rect 8700 16550 8760 16610
rect 8820 16550 8880 16610
rect 8940 16550 9000 16610
rect 9060 16550 9120 16610
rect 9180 16550 9240 16610
rect 9300 16550 9360 16610
rect 9420 16550 9480 16610
rect 9540 16550 9600 16610
rect 9660 16550 9720 16610
rect 9780 16550 9840 16610
rect 9900 16550 9960 16610
rect 10020 16550 10080 16610
rect 10140 16550 10200 16610
rect 10260 16550 10320 16610
rect 10380 16550 10440 16610
rect 10500 16550 10560 16610
rect 10620 16550 10680 16610
rect 10740 16550 10800 16610
rect 10860 16550 10920 16610
rect 10980 16550 11040 16610
rect 11100 16550 11160 16610
rect 11220 16550 11280 16610
rect 11340 16550 11400 16610
rect 320 16440 380 16500
rect 11820 16440 11880 16500
rect 320 16260 380 16320
rect 1195 16210 1255 16270
rect 2125 16210 2185 16270
rect 2455 16210 2515 16270
rect 3385 16210 3445 16270
rect 3715 16210 3775 16270
rect 4645 16210 4705 16270
rect 4975 16210 5035 16270
rect 5905 16210 5965 16270
rect 6235 16210 6295 16270
rect 7165 16210 7225 16270
rect 7495 16210 7555 16270
rect 8425 16210 8485 16270
rect 8755 16210 8815 16270
rect 9685 16210 9745 16270
rect 10015 16210 10075 16270
rect 10945 16210 11005 16270
rect 11820 16260 11880 16320
rect 320 16080 380 16140
rect 11820 16080 11880 16140
rect 320 15900 380 15960
rect 11820 15900 11880 15960
rect 320 15720 380 15780
rect 11820 15720 11880 15780
rect 320 15540 380 15600
rect 1030 15540 1090 15600
rect 1660 15540 1720 15600
rect 2290 15540 2350 15600
rect 2920 15540 2980 15600
rect 3550 15540 3610 15600
rect 4180 15540 4240 15600
rect 4810 15540 4870 15600
rect 5440 15540 5500 15600
rect 6070 15540 6130 15600
rect 6700 15540 6760 15600
rect 7330 15540 7390 15600
rect 7960 15540 8020 15600
rect 8590 15540 8650 15600
rect 9220 15540 9280 15600
rect 9850 15540 9910 15600
rect 10480 15540 10540 15600
rect 11110 15540 11170 15600
rect 11820 15540 11880 15600
rect 320 15360 380 15420
rect 1030 15360 1090 15420
rect 1660 15360 1720 15420
rect 2290 15360 2350 15420
rect 2920 15360 2980 15420
rect 3550 15360 3610 15420
rect 4180 15360 4240 15420
rect 4810 15360 4870 15420
rect 5440 15360 5500 15420
rect 6070 15360 6130 15420
rect 6700 15360 6760 15420
rect 7330 15360 7390 15420
rect 7960 15360 8020 15420
rect 8590 15360 8650 15420
rect 9220 15360 9280 15420
rect 9850 15360 9910 15420
rect 10480 15360 10540 15420
rect 11110 15360 11170 15420
rect 11820 15360 11880 15420
rect 320 15180 380 15240
rect 1030 15180 1090 15240
rect 1660 15180 1720 15240
rect 2290 15180 2350 15240
rect 2920 15180 2980 15240
rect 3550 15180 3610 15240
rect 4180 15180 4240 15240
rect 4810 15180 4870 15240
rect 5440 15180 5500 15240
rect 6070 15180 6130 15240
rect 6700 15180 6760 15240
rect 7330 15180 7390 15240
rect 7960 15180 8020 15240
rect 8590 15180 8650 15240
rect 9220 15180 9280 15240
rect 9850 15180 9910 15240
rect 10480 15180 10540 15240
rect 11110 15180 11170 15240
rect 11820 15180 11880 15240
rect 320 15000 380 15060
rect 1030 15000 1090 15060
rect 1660 15000 1720 15060
rect 2290 15000 2350 15060
rect 2920 15000 2980 15060
rect 3550 15000 3610 15060
rect 4180 15000 4240 15060
rect 4810 15000 4870 15060
rect 5440 15000 5500 15060
rect 6070 15000 6130 15060
rect 6700 15000 6760 15060
rect 7330 15000 7390 15060
rect 7960 15000 8020 15060
rect 8590 15000 8650 15060
rect 9220 15000 9280 15060
rect 9850 15000 9910 15060
rect 10480 15000 10540 15060
rect 11110 15000 11170 15060
rect 11820 15000 11880 15060
rect 320 14820 380 14880
rect 1030 14820 1090 14880
rect 1660 14820 1720 14880
rect 2290 14820 2350 14880
rect 2920 14820 2980 14880
rect 3550 14820 3610 14880
rect 4180 14820 4240 14880
rect 4810 14820 4870 14880
rect 5440 14820 5500 14880
rect 6070 14820 6130 14880
rect 6700 14820 6760 14880
rect 7330 14820 7390 14880
rect 7960 14820 8020 14880
rect 8590 14820 8650 14880
rect 9220 14820 9280 14880
rect 9850 14820 9910 14880
rect 10480 14820 10540 14880
rect 11110 14820 11170 14880
rect 11820 14820 11880 14880
rect 320 14640 380 14700
rect 1030 14640 1090 14700
rect 1660 14640 1720 14700
rect 2290 14640 2350 14700
rect 2920 14640 2980 14700
rect 3550 14640 3610 14700
rect 4180 14640 4240 14700
rect 4810 14640 4870 14700
rect 5440 14640 5500 14700
rect 6070 14640 6130 14700
rect 6700 14640 6760 14700
rect 7330 14640 7390 14700
rect 7960 14640 8020 14700
rect 8590 14640 8650 14700
rect 9220 14640 9280 14700
rect 9850 14640 9910 14700
rect 10480 14640 10540 14700
rect 11110 14640 11170 14700
rect 11820 14640 11880 14700
rect 320 14460 380 14520
rect 1030 14460 1090 14520
rect 1660 14460 1720 14520
rect 2290 14460 2350 14520
rect 2920 14460 2980 14520
rect 3550 14460 3610 14520
rect 4180 14460 4240 14520
rect 4810 14460 4870 14520
rect 5440 14460 5500 14520
rect 6070 14460 6130 14520
rect 6700 14460 6760 14520
rect 7330 14460 7390 14520
rect 7960 14460 8020 14520
rect 8590 14460 8650 14520
rect 9220 14460 9280 14520
rect 9850 14460 9910 14520
rect 10480 14460 10540 14520
rect 11110 14460 11170 14520
rect 11820 14460 11880 14520
rect 320 14280 380 14340
rect 1030 14280 1090 14340
rect 1660 14280 1720 14340
rect 2290 14280 2350 14340
rect 2920 14280 2980 14340
rect 3550 14280 3610 14340
rect 4180 14280 4240 14340
rect 4810 14280 4870 14340
rect 5440 14280 5500 14340
rect 6070 14280 6130 14340
rect 6700 14280 6760 14340
rect 7330 14280 7390 14340
rect 7960 14280 8020 14340
rect 8590 14280 8650 14340
rect 9220 14280 9280 14340
rect 9850 14280 9910 14340
rect 10480 14280 10540 14340
rect 11110 14280 11170 14340
rect 11820 14280 11880 14340
rect 320 14100 380 14160
rect 1030 14100 1090 14160
rect 1660 14100 1720 14160
rect 2290 14100 2350 14160
rect 2920 14100 2980 14160
rect 3550 14100 3610 14160
rect 4180 14100 4240 14160
rect 4810 14100 4870 14160
rect 5440 14100 5500 14160
rect 6070 14100 6130 14160
rect 6700 14100 6760 14160
rect 7330 14100 7390 14160
rect 7960 14100 8020 14160
rect 8590 14100 8650 14160
rect 9220 14100 9280 14160
rect 9850 14100 9910 14160
rect 10480 14100 10540 14160
rect 11110 14100 11170 14160
rect 11820 14100 11880 14160
rect 320 13920 380 13980
rect 1030 13920 1090 13980
rect 1660 13920 1720 13980
rect 2290 13920 2350 13980
rect 2920 13920 2980 13980
rect 3550 13920 3610 13980
rect 4180 13920 4240 13980
rect 4810 13920 4870 13980
rect 5440 13920 5500 13980
rect 6070 13920 6130 13980
rect 6700 13920 6760 13980
rect 7330 13920 7390 13980
rect 7960 13920 8020 13980
rect 8590 13920 8650 13980
rect 9220 13920 9280 13980
rect 9850 13920 9910 13980
rect 10480 13920 10540 13980
rect 11110 13920 11170 13980
rect 11820 13920 11880 13980
rect 320 13740 380 13800
rect 1030 13740 1090 13800
rect 1660 13740 1720 13800
rect 2290 13740 2350 13800
rect 2920 13740 2980 13800
rect 3550 13740 3610 13800
rect 4180 13740 4240 13800
rect 4810 13740 4870 13800
rect 5440 13740 5500 13800
rect 6070 13740 6130 13800
rect 6700 13740 6760 13800
rect 7330 13740 7390 13800
rect 7960 13740 8020 13800
rect 8590 13740 8650 13800
rect 9220 13740 9280 13800
rect 9850 13740 9910 13800
rect 10480 13740 10540 13800
rect 11110 13740 11170 13800
rect 11820 13740 11880 13800
rect 320 13560 380 13620
rect 1030 13560 1090 13620
rect 1660 13560 1720 13620
rect 2290 13560 2350 13620
rect 2920 13560 2980 13620
rect 3550 13560 3610 13620
rect 4180 13560 4240 13620
rect 4810 13560 4870 13620
rect 5440 13560 5500 13620
rect 6070 13560 6130 13620
rect 6700 13560 6760 13620
rect 7330 13560 7390 13620
rect 7960 13560 8020 13620
rect 8590 13560 8650 13620
rect 9220 13560 9280 13620
rect 9850 13560 9910 13620
rect 10480 13560 10540 13620
rect 11110 13560 11170 13620
rect 11820 13560 11880 13620
rect 320 13380 380 13440
rect 1030 13380 1090 13440
rect 1660 13380 1720 13440
rect 2290 13380 2350 13440
rect 2920 13380 2980 13440
rect 3550 13380 3610 13440
rect 4180 13380 4240 13440
rect 4810 13380 4870 13440
rect 5440 13380 5500 13440
rect 6070 13380 6130 13440
rect 6700 13380 6760 13440
rect 7330 13380 7390 13440
rect 7960 13380 8020 13440
rect 8590 13380 8650 13440
rect 9220 13380 9280 13440
rect 9850 13380 9910 13440
rect 10480 13380 10540 13440
rect 11110 13380 11170 13440
rect 11820 13380 11880 13440
rect 320 13200 380 13260
rect 1030 13200 1090 13260
rect 1660 13200 1720 13260
rect 2290 13200 2350 13260
rect 2920 13200 2980 13260
rect 3550 13200 3610 13260
rect 4180 13200 4240 13260
rect 4810 13200 4870 13260
rect 5440 13200 5500 13260
rect 6070 13200 6130 13260
rect 6700 13200 6760 13260
rect 7330 13200 7390 13260
rect 7960 13200 8020 13260
rect 8590 13200 8650 13260
rect 9220 13200 9280 13260
rect 9850 13200 9910 13260
rect 10480 13200 10540 13260
rect 11110 13200 11170 13260
rect 11820 13200 11880 13260
rect 320 13020 380 13080
rect 1030 13020 1090 13080
rect 1660 13020 1720 13080
rect 2290 13020 2350 13080
rect 2920 13020 2980 13080
rect 3550 13020 3610 13080
rect 4180 13020 4240 13080
rect 4810 13020 4870 13080
rect 5440 13020 5500 13080
rect 6070 13020 6130 13080
rect 6700 13020 6760 13080
rect 7330 13020 7390 13080
rect 7960 13020 8020 13080
rect 8590 13020 8650 13080
rect 9220 13020 9280 13080
rect 9850 13020 9910 13080
rect 10480 13020 10540 13080
rect 11110 13020 11170 13080
rect 11820 13020 11880 13080
rect 320 12840 380 12900
rect 1030 12840 1090 12900
rect 1660 12840 1720 12900
rect 2290 12840 2350 12900
rect 2920 12840 2980 12900
rect 3550 12840 3610 12900
rect 4180 12840 4240 12900
rect 4810 12840 4870 12900
rect 5440 12840 5500 12900
rect 6070 12840 6130 12900
rect 6700 12840 6760 12900
rect 7330 12840 7390 12900
rect 7960 12840 8020 12900
rect 8590 12840 8650 12900
rect 9220 12840 9280 12900
rect 9850 12840 9910 12900
rect 10480 12840 10540 12900
rect 11110 12840 11170 12900
rect 11820 12840 11880 12900
rect 320 12660 380 12720
rect 1030 12660 1090 12720
rect 1660 12660 1720 12720
rect 2290 12660 2350 12720
rect 2920 12660 2980 12720
rect 3550 12660 3610 12720
rect 4180 12660 4240 12720
rect 4810 12660 4870 12720
rect 5440 12660 5500 12720
rect 6070 12660 6130 12720
rect 6700 12660 6760 12720
rect 7330 12660 7390 12720
rect 7960 12660 8020 12720
rect 8590 12660 8650 12720
rect 9220 12660 9280 12720
rect 9850 12660 9910 12720
rect 10480 12660 10540 12720
rect 11110 12660 11170 12720
rect 11820 12660 11880 12720
rect 320 12480 380 12540
rect 1030 12480 1090 12540
rect 1660 12480 1720 12540
rect 2290 12480 2350 12540
rect 2920 12480 2980 12540
rect 3550 12480 3610 12540
rect 4180 12480 4240 12540
rect 4810 12480 4870 12540
rect 5440 12480 5500 12540
rect 6070 12480 6130 12540
rect 6700 12480 6760 12540
rect 7330 12480 7390 12540
rect 7960 12480 8020 12540
rect 8590 12480 8650 12540
rect 9220 12480 9280 12540
rect 9850 12480 9910 12540
rect 10480 12480 10540 12540
rect 11110 12480 11170 12540
rect 11820 12480 11880 12540
rect 320 12300 380 12360
rect 1030 12300 1090 12360
rect 1660 12300 1720 12360
rect 2290 12300 2350 12360
rect 2920 12300 2980 12360
rect 3550 12300 3610 12360
rect 4180 12300 4240 12360
rect 4810 12300 4870 12360
rect 5440 12300 5500 12360
rect 6070 12300 6130 12360
rect 6700 12300 6760 12360
rect 7330 12300 7390 12360
rect 7960 12300 8020 12360
rect 8590 12300 8650 12360
rect 9220 12300 9280 12360
rect 9850 12300 9910 12360
rect 10480 12300 10540 12360
rect 11110 12300 11170 12360
rect 11820 12300 11880 12360
rect 320 12120 380 12180
rect 1030 12120 1090 12180
rect 1660 12120 1720 12180
rect 2290 12120 2350 12180
rect 2920 12120 2980 12180
rect 3550 12120 3610 12180
rect 4180 12120 4240 12180
rect 4810 12120 4870 12180
rect 5440 12120 5500 12180
rect 6070 12120 6130 12180
rect 6700 12120 6760 12180
rect 7330 12120 7390 12180
rect 7960 12120 8020 12180
rect 8590 12120 8650 12180
rect 9220 12120 9280 12180
rect 9850 12120 9910 12180
rect 10480 12120 10540 12180
rect 11110 12120 11170 12180
rect 11820 12120 11880 12180
rect 320 11940 380 12000
rect 1030 11940 1090 12000
rect 1660 11940 1720 12000
rect 2290 11940 2350 12000
rect 2920 11940 2980 12000
rect 3550 11940 3610 12000
rect 4180 11940 4240 12000
rect 4810 11940 4870 12000
rect 5440 11940 5500 12000
rect 6070 11940 6130 12000
rect 6700 11940 6760 12000
rect 7330 11940 7390 12000
rect 7960 11940 8020 12000
rect 8590 11940 8650 12000
rect 9220 11940 9280 12000
rect 9850 11940 9910 12000
rect 10480 11940 10540 12000
rect 11110 11940 11170 12000
rect 11820 11940 11880 12000
rect 320 11760 380 11820
rect 1030 11760 1090 11820
rect 1660 11760 1720 11820
rect 2290 11760 2350 11820
rect 2920 11760 2980 11820
rect 3550 11760 3610 11820
rect 4180 11760 4240 11820
rect 4810 11760 4870 11820
rect 5440 11760 5500 11820
rect 6070 11760 6130 11820
rect 6700 11760 6760 11820
rect 7330 11760 7390 11820
rect 7960 11760 8020 11820
rect 8590 11760 8650 11820
rect 9220 11760 9280 11820
rect 9850 11760 9910 11820
rect 10480 11760 10540 11820
rect 11110 11760 11170 11820
rect 11820 11760 11880 11820
rect 320 11580 380 11640
rect 1030 11580 1090 11640
rect 1660 11580 1720 11640
rect 2290 11580 2350 11640
rect 2920 11580 2980 11640
rect 3550 11580 3610 11640
rect 4180 11580 4240 11640
rect 4810 11580 4870 11640
rect 5440 11580 5500 11640
rect 6070 11580 6130 11640
rect 6700 11580 6760 11640
rect 7330 11580 7390 11640
rect 7960 11580 8020 11640
rect 8590 11580 8650 11640
rect 9220 11580 9280 11640
rect 9850 11580 9910 11640
rect 10480 11580 10540 11640
rect 11110 11580 11170 11640
rect 11820 11580 11880 11640
rect 320 11400 380 11460
rect 1030 11400 1090 11460
rect 1660 11400 1720 11460
rect 2290 11400 2350 11460
rect 2920 11400 2980 11460
rect 3550 11400 3610 11460
rect 4180 11400 4240 11460
rect 4810 11400 4870 11460
rect 5440 11400 5500 11460
rect 6070 11400 6130 11460
rect 6700 11400 6760 11460
rect 7330 11400 7390 11460
rect 7960 11400 8020 11460
rect 8590 11400 8650 11460
rect 9220 11400 9280 11460
rect 9850 11400 9910 11460
rect 10480 11400 10540 11460
rect 11110 11400 11170 11460
rect 11820 11400 11880 11460
rect 320 11220 380 11280
rect 1030 11220 1090 11280
rect 1660 11220 1720 11280
rect 2290 11220 2350 11280
rect 2920 11220 2980 11280
rect 3550 11220 3610 11280
rect 4180 11220 4240 11280
rect 4810 11220 4870 11280
rect 5440 11220 5500 11280
rect 6070 11220 6130 11280
rect 6700 11220 6760 11280
rect 7330 11220 7390 11280
rect 7960 11220 8020 11280
rect 8590 11220 8650 11280
rect 9220 11220 9280 11280
rect 9850 11220 9910 11280
rect 10480 11220 10540 11280
rect 11110 11220 11170 11280
rect 11820 11220 11880 11280
rect 320 11040 380 11100
rect 1030 11040 1090 11100
rect 1660 11040 1720 11100
rect 2290 11040 2350 11100
rect 2920 11040 2980 11100
rect 3550 11040 3610 11100
rect 4180 11040 4240 11100
rect 4810 11040 4870 11100
rect 5440 11040 5500 11100
rect 6070 11040 6130 11100
rect 6700 11040 6760 11100
rect 7330 11040 7390 11100
rect 7960 11040 8020 11100
rect 8590 11040 8650 11100
rect 9220 11040 9280 11100
rect 9850 11040 9910 11100
rect 10480 11040 10540 11100
rect 11110 11040 11170 11100
rect 11820 11040 11880 11100
rect 320 10860 380 10920
rect 1030 10860 1090 10920
rect 1660 10860 1720 10920
rect 2290 10860 2350 10920
rect 2920 10860 2980 10920
rect 3550 10860 3610 10920
rect 4180 10860 4240 10920
rect 4810 10860 4870 10920
rect 5440 10860 5500 10920
rect 6070 10860 6130 10920
rect 6700 10860 6760 10920
rect 7330 10860 7390 10920
rect 7960 10860 8020 10920
rect 8590 10860 8650 10920
rect 9220 10860 9280 10920
rect 9850 10860 9910 10920
rect 10480 10860 10540 10920
rect 11110 10860 11170 10920
rect 11820 10860 11880 10920
rect 320 10680 380 10740
rect 1030 10680 1090 10740
rect 1660 10680 1720 10740
rect 2290 10680 2350 10740
rect 2920 10680 2980 10740
rect 3550 10680 3610 10740
rect 4180 10680 4240 10740
rect 4810 10680 4870 10740
rect 5440 10680 5500 10740
rect 6070 10680 6130 10740
rect 6700 10680 6760 10740
rect 7330 10680 7390 10740
rect 7960 10680 8020 10740
rect 8590 10680 8650 10740
rect 9220 10680 9280 10740
rect 9850 10680 9910 10740
rect 10480 10680 10540 10740
rect 11110 10680 11170 10740
rect 11820 10680 11880 10740
rect 320 10500 380 10560
rect 1030 10500 1090 10560
rect 1660 10500 1720 10560
rect 2290 10500 2350 10560
rect 2920 10500 2980 10560
rect 3550 10500 3610 10560
rect 4180 10500 4240 10560
rect 4810 10500 4870 10560
rect 5440 10500 5500 10560
rect 6070 10500 6130 10560
rect 6700 10500 6760 10560
rect 7330 10500 7390 10560
rect 7960 10500 8020 10560
rect 8590 10500 8650 10560
rect 9220 10500 9280 10560
rect 9850 10500 9910 10560
rect 10480 10500 10540 10560
rect 11110 10500 11170 10560
rect 11820 10500 11880 10560
rect 320 10320 380 10380
rect 11820 10320 11880 10380
rect 320 10140 380 10200
rect 11820 10140 11880 10200
rect 320 9960 380 10020
rect 11820 9960 11880 10020
rect 320 9780 380 9840
rect 11820 9780 11880 9840
rect 320 9600 380 9660
rect 11820 9600 11880 9660
rect 660 9500 720 9560
rect 780 9500 840 9560
rect 900 9500 960 9560
rect 1020 9500 1080 9560
rect 1140 9500 1200 9560
rect 1260 9500 1320 9560
rect 1380 9500 1440 9560
rect 1500 9500 1560 9560
rect 1620 9500 1680 9560
rect 1740 9500 1800 9560
rect 1860 9500 1920 9560
rect 1980 9500 2040 9560
rect 2100 9500 2160 9560
rect 2220 9500 2280 9560
rect 2340 9500 2400 9560
rect 2460 9500 2520 9560
rect 2580 9500 2640 9560
rect 2700 9500 2760 9560
rect 2820 9500 2880 9560
rect 2940 9500 3000 9560
rect 3060 9500 3120 9560
rect 3180 9500 3240 9560
rect 3300 9500 3360 9560
rect 3420 9500 3480 9560
rect 3540 9500 3600 9560
rect 3660 9500 3720 9560
rect 3780 9500 3840 9560
rect 3900 9500 3960 9560
rect 4020 9500 4080 9560
rect 4140 9500 4200 9560
rect 4260 9500 4320 9560
rect 4380 9500 4440 9560
rect 4500 9500 4560 9560
rect 4620 9500 4680 9560
rect 4740 9500 4800 9560
rect 4860 9500 4920 9560
rect 4980 9500 5040 9560
rect 5100 9500 5160 9560
rect 5220 9500 5280 9560
rect 5340 9500 5400 9560
rect 5460 9500 5520 9560
rect 5580 9500 5640 9560
rect 5700 9500 5760 9560
rect 5820 9500 5880 9560
rect 5940 9500 6000 9560
rect 6060 9500 6120 9560
rect 6180 9500 6240 9560
rect 6300 9500 6360 9560
rect 6420 9500 6480 9560
rect 6540 9500 6600 9560
rect 6660 9500 6720 9560
rect 6780 9500 6840 9560
rect 6900 9500 6960 9560
rect 7020 9500 7080 9560
rect 7140 9500 7200 9560
rect 7260 9500 7320 9560
rect 7380 9500 7440 9560
rect 7500 9500 7560 9560
rect 7620 9500 7680 9560
rect 7740 9500 7800 9560
rect 7860 9500 7920 9560
rect 7980 9500 8040 9560
rect 8100 9500 8160 9560
rect 8220 9500 8280 9560
rect 8340 9500 8400 9560
rect 8460 9500 8520 9560
rect 8580 9500 8640 9560
rect 8700 9500 8760 9560
rect 8820 9500 8880 9560
rect 8940 9500 9000 9560
rect 9060 9500 9120 9560
rect 9180 9500 9240 9560
rect 9300 9500 9360 9560
rect 9420 9500 9480 9560
rect 9540 9500 9600 9560
rect 9660 9500 9720 9560
rect 9780 9500 9840 9560
rect 9900 9500 9960 9560
rect 10020 9500 10080 9560
rect 10140 9500 10200 9560
rect 10260 9500 10320 9560
rect 10380 9500 10440 9560
rect 10500 9500 10560 9560
rect 10620 9500 10680 9560
rect 10740 9500 10800 9560
rect 10860 9500 10920 9560
rect 10980 9500 11040 9560
rect 11100 9500 11160 9560
rect 11220 9500 11280 9560
rect 11340 9500 11400 9560
rect 320 9420 380 9480
rect 660 9380 720 9440
rect 780 9380 840 9440
rect 900 9380 960 9440
rect 1020 9380 1080 9440
rect 1140 9380 1200 9440
rect 1260 9380 1320 9440
rect 1380 9380 1440 9440
rect 1500 9380 1560 9440
rect 1620 9380 1680 9440
rect 1740 9380 1800 9440
rect 1860 9380 1920 9440
rect 1980 9380 2040 9440
rect 2100 9380 2160 9440
rect 2220 9380 2280 9440
rect 2340 9380 2400 9440
rect 2460 9380 2520 9440
rect 2580 9380 2640 9440
rect 2700 9380 2760 9440
rect 2820 9380 2880 9440
rect 2940 9380 3000 9440
rect 3060 9380 3120 9440
rect 3180 9380 3240 9440
rect 3300 9380 3360 9440
rect 3420 9380 3480 9440
rect 3540 9380 3600 9440
rect 3660 9380 3720 9440
rect 3780 9380 3840 9440
rect 3900 9380 3960 9440
rect 4020 9380 4080 9440
rect 4140 9380 4200 9440
rect 4260 9380 4320 9440
rect 4380 9380 4440 9440
rect 4500 9380 4560 9440
rect 4620 9380 4680 9440
rect 4740 9380 4800 9440
rect 4860 9380 4920 9440
rect 4980 9380 5040 9440
rect 5100 9380 5160 9440
rect 5220 9380 5280 9440
rect 5340 9380 5400 9440
rect 5460 9380 5520 9440
rect 5580 9380 5640 9440
rect 5700 9380 5760 9440
rect 5820 9380 5880 9440
rect 5940 9380 6000 9440
rect 6060 9380 6120 9440
rect 6180 9380 6240 9440
rect 6300 9380 6360 9440
rect 6420 9380 6480 9440
rect 6540 9380 6600 9440
rect 6660 9380 6720 9440
rect 6780 9380 6840 9440
rect 6900 9380 6960 9440
rect 7020 9380 7080 9440
rect 7140 9380 7200 9440
rect 7260 9380 7320 9440
rect 7380 9380 7440 9440
rect 7500 9380 7560 9440
rect 7620 9380 7680 9440
rect 7740 9380 7800 9440
rect 7860 9380 7920 9440
rect 7980 9380 8040 9440
rect 8100 9380 8160 9440
rect 8220 9380 8280 9440
rect 8340 9380 8400 9440
rect 8460 9380 8520 9440
rect 8580 9380 8640 9440
rect 8700 9380 8760 9440
rect 8820 9380 8880 9440
rect 8940 9380 9000 9440
rect 9060 9380 9120 9440
rect 9180 9380 9240 9440
rect 9300 9380 9360 9440
rect 9420 9380 9480 9440
rect 9540 9380 9600 9440
rect 9660 9380 9720 9440
rect 9780 9380 9840 9440
rect 9900 9380 9960 9440
rect 10020 9380 10080 9440
rect 10140 9380 10200 9440
rect 10260 9380 10320 9440
rect 10380 9380 10440 9440
rect 10500 9380 10560 9440
rect 10620 9380 10680 9440
rect 10740 9380 10800 9440
rect 10860 9380 10920 9440
rect 10980 9380 11040 9440
rect 11100 9380 11160 9440
rect 11220 9380 11280 9440
rect 11340 9380 11400 9440
rect 11820 9420 11880 9480
rect 320 9240 380 9300
rect 660 9260 720 9320
rect 780 9260 840 9320
rect 900 9260 960 9320
rect 1020 9260 1080 9320
rect 1140 9260 1200 9320
rect 1260 9260 1320 9320
rect 1380 9260 1440 9320
rect 1500 9260 1560 9320
rect 1620 9260 1680 9320
rect 1740 9260 1800 9320
rect 1860 9260 1920 9320
rect 1980 9260 2040 9320
rect 2100 9260 2160 9320
rect 2220 9260 2280 9320
rect 2340 9260 2400 9320
rect 2460 9260 2520 9320
rect 2580 9260 2640 9320
rect 2700 9260 2760 9320
rect 2820 9260 2880 9320
rect 2940 9260 3000 9320
rect 3060 9260 3120 9320
rect 3180 9260 3240 9320
rect 3300 9260 3360 9320
rect 3420 9260 3480 9320
rect 3540 9260 3600 9320
rect 3660 9260 3720 9320
rect 3780 9260 3840 9320
rect 3900 9260 3960 9320
rect 4020 9260 4080 9320
rect 4140 9260 4200 9320
rect 4260 9260 4320 9320
rect 4380 9260 4440 9320
rect 4500 9260 4560 9320
rect 4620 9260 4680 9320
rect 4740 9260 4800 9320
rect 4860 9260 4920 9320
rect 4980 9260 5040 9320
rect 5100 9260 5160 9320
rect 5220 9260 5280 9320
rect 5340 9260 5400 9320
rect 5460 9260 5520 9320
rect 5580 9260 5640 9320
rect 5700 9260 5760 9320
rect 5820 9260 5880 9320
rect 5940 9260 6000 9320
rect 6060 9260 6120 9320
rect 6180 9260 6240 9320
rect 6300 9260 6360 9320
rect 6420 9260 6480 9320
rect 6540 9260 6600 9320
rect 6660 9260 6720 9320
rect 6780 9260 6840 9320
rect 6900 9260 6960 9320
rect 7020 9260 7080 9320
rect 7140 9260 7200 9320
rect 7260 9260 7320 9320
rect 7380 9260 7440 9320
rect 7500 9260 7560 9320
rect 7620 9260 7680 9320
rect 7740 9260 7800 9320
rect 7860 9260 7920 9320
rect 7980 9260 8040 9320
rect 8100 9260 8160 9320
rect 8220 9260 8280 9320
rect 8340 9260 8400 9320
rect 8460 9260 8520 9320
rect 8580 9260 8640 9320
rect 8700 9260 8760 9320
rect 8820 9260 8880 9320
rect 8940 9260 9000 9320
rect 9060 9260 9120 9320
rect 9180 9260 9240 9320
rect 9300 9260 9360 9320
rect 9420 9260 9480 9320
rect 9540 9260 9600 9320
rect 9660 9260 9720 9320
rect 9780 9260 9840 9320
rect 9900 9260 9960 9320
rect 10020 9260 10080 9320
rect 10140 9260 10200 9320
rect 10260 9260 10320 9320
rect 10380 9260 10440 9320
rect 10500 9260 10560 9320
rect 10620 9260 10680 9320
rect 10740 9260 10800 9320
rect 10860 9260 10920 9320
rect 10980 9260 11040 9320
rect 11100 9260 11160 9320
rect 11220 9260 11280 9320
rect 11340 9260 11400 9320
rect 11820 9240 11880 9300
<< metal1 >>
rect 100 34030 12100 34210
rect 100 32730 300 34030
rect 7770 33920 8990 34030
rect 7770 33860 7960 33920
rect 8020 33860 8220 33920
rect 8280 33860 8480 33920
rect 8540 33860 8740 33920
rect 8800 33860 8990 33920
rect 7770 33800 8990 33860
rect 7770 33610 7950 33800
rect 7770 33550 7830 33610
rect 7890 33550 7950 33610
rect 7770 33490 7950 33550
rect 7770 33430 7830 33490
rect 7890 33430 7950 33490
rect 7770 33370 7950 33430
rect 7770 33310 7830 33370
rect 7890 33310 7950 33370
rect 7770 33200 7950 33310
rect 8030 33610 8210 33720
rect 8030 33550 8090 33610
rect 8150 33550 8210 33610
rect 8030 33490 8210 33550
rect 8030 33430 8090 33490
rect 8150 33430 8210 33490
rect 8030 33370 8210 33430
rect 8030 33310 8090 33370
rect 8150 33310 8210 33370
rect 8030 33105 8210 33310
rect 8290 33610 8470 33800
rect 8290 33550 8350 33610
rect 8410 33550 8470 33610
rect 8290 33490 8470 33550
rect 8290 33430 8350 33490
rect 8410 33430 8470 33490
rect 8290 33370 8470 33430
rect 8290 33310 8350 33370
rect 8410 33310 8470 33370
rect 8290 33200 8470 33310
rect 8550 33610 8730 33720
rect 8550 33550 8610 33610
rect 8670 33550 8730 33610
rect 8550 33490 8730 33550
rect 8550 33430 8610 33490
rect 8670 33430 8730 33490
rect 8550 33370 8730 33430
rect 8550 33310 8610 33370
rect 8670 33310 8730 33370
rect 8550 33105 8730 33310
rect 8810 33610 8990 33800
rect 10250 33830 11640 33950
rect 8810 33550 8870 33610
rect 8930 33550 8990 33610
rect 8810 33490 8990 33550
rect 8810 33430 8870 33490
rect 8930 33430 8990 33490
rect 8810 33370 8990 33430
rect 8810 33310 8870 33370
rect 8930 33310 8990 33370
rect 8810 33200 8990 33310
rect 9080 33530 9290 33750
rect 9080 33470 9150 33530
rect 9210 33470 9290 33530
rect 9080 33250 9290 33470
rect 9080 33190 9150 33250
rect 9210 33190 9290 33250
rect 9080 33110 9290 33190
rect 9370 33530 9580 33750
rect 9370 33470 9450 33530
rect 9510 33470 9580 33530
rect 9370 33250 9580 33470
rect 9370 33190 9450 33250
rect 9510 33190 9580 33250
rect 9370 33110 9580 33190
rect 9960 33530 10170 33750
rect 9960 33470 10030 33530
rect 10090 33470 10170 33530
rect 9960 33250 10170 33470
rect 9960 33190 10030 33250
rect 10090 33190 10170 33250
rect 9960 33110 10170 33190
rect 10250 33530 10460 33830
rect 10250 33470 10330 33530
rect 10390 33470 10460 33530
rect 10250 33250 10460 33470
rect 10250 33190 10330 33250
rect 10390 33190 10460 33250
rect 10250 33110 10460 33190
rect 10550 33530 10760 33750
rect 10550 33470 10620 33530
rect 10680 33470 10760 33530
rect 10550 33250 10760 33470
rect 10550 33190 10620 33250
rect 10680 33190 10760 33250
rect 10550 33110 10760 33190
rect 10840 33530 11050 33830
rect 10840 33470 10920 33530
rect 10980 33470 11050 33530
rect 10840 33250 11050 33470
rect 10840 33190 10920 33250
rect 10980 33190 11050 33250
rect 10840 33110 11050 33190
rect 11140 33530 11350 33750
rect 11140 33470 11210 33530
rect 11270 33470 11350 33530
rect 11140 33250 11350 33470
rect 11140 33190 11210 33250
rect 11270 33190 11350 33250
rect 11140 33110 11350 33190
rect 11430 33530 11640 33830
rect 11430 33470 11510 33530
rect 11570 33470 11640 33530
rect 11430 33250 11640 33470
rect 11430 33190 11510 33250
rect 11570 33190 11640 33250
rect 11430 33110 11640 33190
rect 8030 33042 8730 33105
rect 8030 32965 8170 33042
rect 8110 32962 8170 32965
rect 8250 32962 8370 33042
rect 8450 32962 8570 33042
rect 8650 32965 8730 33042
rect 8650 32962 8710 32965
rect 8110 32902 8710 32962
rect 8940 32950 9420 33030
rect 8940 32890 9300 32950
rect 9360 32890 9420 32950
rect 8940 32810 9420 32890
rect 10120 32950 11480 33030
rect 10120 32890 10180 32950
rect 10240 32890 10770 32950
rect 10830 32890 11360 32950
rect 11420 32890 11480 32950
rect 10120 32810 11480 32890
rect 11900 32730 12100 34030
rect 100 32550 12100 32730
rect 100 31730 12100 31910
rect 100 30430 300 31730
rect 8800 31570 9420 31650
rect 8800 31510 9000 31570
rect 9060 31510 9300 31570
rect 9360 31510 9420 31570
rect 8800 31450 9420 31510
rect 9820 31570 11500 31650
rect 9820 31510 9880 31570
rect 9940 31510 10180 31570
rect 10240 31510 10480 31570
rect 10540 31510 10780 31570
rect 10840 31510 11080 31570
rect 11140 31510 11380 31570
rect 11440 31510 11500 31570
rect 9820 31450 11500 31510
rect 8780 31270 8990 31350
rect 5830 31253 6010 31255
rect 8290 31253 8470 31255
rect 5830 30855 6998 31253
rect 5901 30853 6998 30855
rect 8111 30853 8631 31253
rect 8780 31210 8850 31270
rect 8910 31210 8990 31270
rect 8780 30990 8990 31210
rect 8780 30930 8850 30990
rect 8910 30930 8990 30990
rect 8780 30630 8990 30930
rect 9070 31270 9290 31350
rect 9070 31210 9150 31270
rect 9210 31210 9290 31270
rect 9070 30990 9290 31210
rect 9070 30930 9150 30990
rect 9210 30930 9290 30990
rect 9070 30710 9290 30930
rect 9370 31270 9580 31350
rect 9370 31210 9450 31270
rect 9510 31210 9580 31270
rect 9370 30990 9580 31210
rect 9370 30930 9450 30990
rect 9510 30930 9580 30990
rect 9370 30630 9580 30930
rect 8780 30510 9580 30630
rect 9660 31270 9870 31350
rect 9660 31210 9730 31270
rect 9790 31210 9870 31270
rect 9660 30990 9870 31210
rect 9660 30930 9730 30990
rect 9790 30930 9870 30990
rect 9660 30630 9870 30930
rect 9950 31270 10170 31350
rect 9950 31210 10030 31270
rect 10090 31210 10170 31270
rect 9950 30990 10170 31210
rect 9950 30930 10030 30990
rect 10090 30930 10170 30990
rect 9950 30710 10170 30930
rect 10250 31270 10460 31350
rect 10250 31210 10330 31270
rect 10390 31210 10460 31270
rect 10250 30990 10460 31210
rect 10250 30930 10330 30990
rect 10390 30930 10460 30990
rect 10250 30710 10460 30930
rect 10550 31270 10770 31350
rect 10550 31210 10630 31270
rect 10690 31210 10770 31270
rect 10550 30990 10770 31210
rect 10550 30930 10630 30990
rect 10690 30930 10770 30990
rect 10550 30710 10770 30930
rect 10850 31270 11060 31350
rect 10850 31210 10930 31270
rect 10990 31210 11060 31270
rect 10850 30990 11060 31210
rect 10850 30930 10930 30990
rect 10990 30930 11060 30990
rect 10850 30710 11060 30930
rect 11150 31270 11370 31350
rect 11150 31210 11230 31270
rect 11290 31210 11370 31270
rect 11150 30990 11370 31210
rect 11150 30930 11230 30990
rect 11290 30930 11370 30990
rect 11150 30710 11370 30930
rect 11450 31270 11660 31350
rect 11450 31210 11530 31270
rect 11590 31210 11660 31270
rect 11450 30990 11660 31210
rect 11450 30930 11530 30990
rect 11590 30930 11660 30990
rect 10250 30630 10470 30710
rect 10850 30630 11070 30710
rect 11450 30630 11660 30930
rect 9660 30510 11660 30630
rect 11900 30430 12100 31730
rect 100 30250 12100 30430
rect 100 28750 12100 29750
rect 100 27450 12100 28250
rect 100 20950 600 27450
rect 810 21350 1310 27350
rect 1390 21350 1990 27350
rect 2070 21350 2570 27350
rect 2650 21350 3250 27350
rect 3330 21350 3830 27350
rect 3910 21350 4510 27350
rect 4590 21350 5090 27350
rect 5170 21350 5770 27350
rect 5850 21350 6350 27350
rect 6430 21350 7030 27350
rect 7110 21350 7610 27350
rect 7690 21350 8290 27350
rect 8370 21350 8870 27350
rect 8950 21350 9550 27350
rect 9630 21350 10130 27350
rect 10210 21350 10810 27350
rect 10890 21350 11390 27350
rect 11600 20950 12100 27450
rect 100 20450 12100 20950
rect 100 18950 12100 19950
rect 100 17450 12100 18450
rect 100 16150 12100 16950
rect 100 9650 600 16150
rect 810 10050 1310 16050
rect 1390 10050 1990 16050
rect 2070 10050 2570 16050
rect 2650 10050 3250 16050
rect 3330 10050 3830 16050
rect 3910 10050 4510 16050
rect 4590 10050 5090 16050
rect 5170 10050 5770 16050
rect 5850 10050 6350 16050
rect 6430 10050 7030 16050
rect 7110 10050 7610 16050
rect 7690 10050 8290 16050
rect 8370 10050 8870 16050
rect 8950 10050 9550 16050
rect 9630 10050 10130 16050
rect 10210 10050 10810 16050
rect 10890 10050 11390 16050
rect 11600 9650 12100 16150
rect 100 9150 12100 9650
rect 1850 8250 10350 8500
rect 1850 250 2100 8250
rect 2200 8090 2400 8150
rect 2200 8010 2260 8090
rect 2340 8010 2400 8090
rect 2200 7950 2400 8010
rect 2600 8090 2800 8150
rect 2600 8010 2660 8090
rect 2740 8010 2800 8090
rect 2600 7950 2800 8010
rect 3000 8090 3200 8150
rect 3000 8010 3060 8090
rect 3140 8010 3200 8090
rect 3000 7950 3200 8010
rect 3400 8090 3600 8150
rect 3400 8010 3460 8090
rect 3540 8010 3600 8090
rect 3400 7950 3600 8010
rect 3800 8090 4000 8150
rect 3800 8010 3860 8090
rect 3940 8010 4000 8090
rect 3800 7950 4000 8010
rect 4200 8090 4400 8150
rect 4200 8010 4260 8090
rect 4340 8010 4400 8090
rect 4200 7950 4400 8010
rect 4600 8090 4800 8150
rect 4600 8010 4660 8090
rect 4740 8010 4800 8090
rect 4600 7950 4800 8010
rect 5000 8090 5200 8150
rect 5000 8010 5060 8090
rect 5140 8010 5200 8090
rect 5000 7950 5200 8010
rect 5400 8090 5600 8150
rect 5400 8010 5460 8090
rect 5540 8010 5600 8090
rect 5400 7950 5600 8010
rect 5800 8090 6000 8150
rect 5800 8010 5860 8090
rect 5940 8010 6000 8090
rect 5800 7950 6000 8010
rect 6200 8090 6400 8150
rect 6200 8010 6260 8090
rect 6340 8010 6400 8090
rect 6200 7950 6400 8010
rect 6600 8090 6800 8150
rect 6600 8010 6660 8090
rect 6740 8010 6800 8090
rect 6600 7950 6800 8010
rect 7000 8090 7200 8150
rect 7000 8010 7060 8090
rect 7140 8010 7200 8090
rect 7000 7950 7200 8010
rect 7400 8090 7600 8150
rect 7400 8010 7460 8090
rect 7540 8010 7600 8090
rect 7400 7950 7600 8010
rect 7800 8090 8000 8150
rect 7800 8010 7860 8090
rect 7940 8010 8000 8090
rect 7800 7950 8000 8010
rect 8200 8090 8400 8150
rect 8200 8010 8260 8090
rect 8340 8010 8400 8090
rect 8200 7950 8400 8010
rect 8600 8090 8800 8150
rect 8600 8010 8660 8090
rect 8740 8010 8800 8090
rect 8600 7950 8800 8010
rect 9000 8090 9200 8150
rect 9000 8010 9060 8090
rect 9140 8010 9200 8090
rect 9000 7950 9200 8010
rect 9400 8090 9600 8150
rect 9400 8010 9460 8090
rect 9540 8010 9600 8090
rect 9400 7950 9600 8010
rect 9800 8090 10000 8150
rect 9800 8010 9860 8090
rect 9940 8010 10000 8090
rect 9800 7950 10000 8010
rect 2200 7690 2400 7750
rect 2200 7610 2260 7690
rect 2340 7610 2400 7690
rect 2200 7550 2400 7610
rect 2600 7690 2800 7750
rect 2600 7610 2660 7690
rect 2740 7610 2800 7690
rect 2600 7550 2800 7610
rect 3000 7690 3200 7750
rect 3000 7610 3060 7690
rect 3140 7610 3200 7690
rect 3000 7550 3200 7610
rect 3400 7690 3600 7750
rect 3400 7610 3460 7690
rect 3540 7610 3600 7690
rect 3400 7550 3600 7610
rect 3800 7690 4000 7750
rect 3800 7610 3860 7690
rect 3940 7610 4000 7690
rect 3800 7550 4000 7610
rect 4200 7690 4400 7750
rect 4200 7610 4260 7690
rect 4340 7610 4400 7690
rect 4200 7550 4400 7610
rect 4600 7690 4800 7750
rect 4600 7610 4660 7690
rect 4740 7610 4800 7690
rect 4600 7550 4800 7610
rect 5000 7690 5200 7750
rect 5000 7610 5060 7690
rect 5140 7610 5200 7690
rect 5000 7550 5200 7610
rect 5400 7690 5600 7750
rect 5400 7610 5460 7690
rect 5540 7610 5600 7690
rect 5400 7550 5600 7610
rect 5800 7690 6000 7750
rect 5800 7610 5860 7690
rect 5940 7610 6000 7690
rect 5800 7550 6000 7610
rect 6200 7690 6400 7750
rect 6200 7610 6260 7690
rect 6340 7610 6400 7690
rect 6200 7550 6400 7610
rect 6600 7690 6800 7750
rect 6600 7610 6660 7690
rect 6740 7610 6800 7690
rect 6600 7550 6800 7610
rect 7000 7690 7200 7750
rect 7000 7610 7060 7690
rect 7140 7610 7200 7690
rect 7000 7550 7200 7610
rect 7400 7690 7600 7750
rect 7400 7610 7460 7690
rect 7540 7610 7600 7690
rect 7400 7550 7600 7610
rect 7800 7690 8000 7750
rect 7800 7610 7860 7690
rect 7940 7610 8000 7690
rect 7800 7550 8000 7610
rect 8200 7690 8400 7750
rect 8200 7610 8260 7690
rect 8340 7610 8400 7690
rect 8200 7550 8400 7610
rect 8600 7690 8800 7750
rect 8600 7610 8660 7690
rect 8740 7610 8800 7690
rect 8600 7550 8800 7610
rect 9000 7690 9200 7750
rect 9000 7610 9060 7690
rect 9140 7610 9200 7690
rect 9000 7550 9200 7610
rect 9400 7690 9600 7750
rect 9400 7610 9460 7690
rect 9540 7610 9600 7690
rect 9400 7550 9600 7610
rect 9800 7690 10000 7750
rect 9800 7610 9860 7690
rect 9940 7610 10000 7690
rect 9800 7550 10000 7610
rect 2200 7290 2400 7350
rect 2200 7210 2260 7290
rect 2340 7210 2400 7290
rect 2200 7150 2400 7210
rect 2600 7290 2800 7350
rect 2600 7210 2660 7290
rect 2740 7210 2800 7290
rect 2600 7150 2800 7210
rect 3000 7290 3200 7350
rect 3000 7210 3060 7290
rect 3140 7210 3200 7290
rect 3000 7150 3200 7210
rect 3400 7290 3600 7350
rect 3400 7210 3460 7290
rect 3540 7210 3600 7290
rect 3400 7150 3600 7210
rect 3800 7290 4000 7350
rect 3800 7210 3860 7290
rect 3940 7210 4000 7290
rect 3800 7150 4000 7210
rect 4200 7290 4400 7350
rect 4200 7210 4260 7290
rect 4340 7210 4400 7290
rect 4200 7150 4400 7210
rect 4600 7290 4800 7350
rect 4600 7210 4660 7290
rect 4740 7210 4800 7290
rect 4600 7150 4800 7210
rect 5000 7290 5200 7350
rect 5000 7210 5060 7290
rect 5140 7210 5200 7290
rect 5000 7150 5200 7210
rect 5400 7290 5600 7350
rect 5400 7210 5460 7290
rect 5540 7210 5600 7290
rect 5400 7150 5600 7210
rect 5800 7290 6000 7350
rect 5800 7210 5860 7290
rect 5940 7210 6000 7290
rect 5800 7150 6000 7210
rect 6200 7290 6400 7350
rect 6200 7210 6260 7290
rect 6340 7210 6400 7290
rect 6200 7150 6400 7210
rect 6600 7290 6800 7350
rect 6600 7210 6660 7290
rect 6740 7210 6800 7290
rect 6600 7150 6800 7210
rect 7000 7290 7200 7350
rect 7000 7210 7060 7290
rect 7140 7210 7200 7290
rect 7000 7150 7200 7210
rect 7400 7290 7600 7350
rect 7400 7210 7460 7290
rect 7540 7210 7600 7290
rect 7400 7150 7600 7210
rect 7800 7290 8000 7350
rect 7800 7210 7860 7290
rect 7940 7210 8000 7290
rect 7800 7150 8000 7210
rect 8200 7290 8400 7350
rect 8200 7210 8260 7290
rect 8340 7210 8400 7290
rect 8200 7150 8400 7210
rect 8600 7290 8800 7350
rect 8600 7210 8660 7290
rect 8740 7210 8800 7290
rect 8600 7150 8800 7210
rect 9000 7290 9200 7350
rect 9000 7210 9060 7290
rect 9140 7210 9200 7290
rect 9000 7150 9200 7210
rect 9400 7290 9600 7350
rect 9400 7210 9460 7290
rect 9540 7210 9600 7290
rect 9400 7150 9600 7210
rect 9800 7290 10000 7350
rect 9800 7210 9860 7290
rect 9940 7210 10000 7290
rect 9800 7150 10000 7210
rect 2200 6890 2400 6950
rect 2200 6810 2260 6890
rect 2340 6810 2400 6890
rect 2200 6750 2400 6810
rect 2600 6890 2800 6950
rect 2600 6810 2660 6890
rect 2740 6810 2800 6890
rect 2600 6750 2800 6810
rect 3000 6890 3200 6950
rect 3000 6810 3060 6890
rect 3140 6810 3200 6890
rect 3000 6750 3200 6810
rect 3400 6890 3600 6950
rect 3400 6810 3460 6890
rect 3540 6810 3600 6890
rect 3400 6750 3600 6810
rect 3800 6890 4000 6950
rect 3800 6810 3860 6890
rect 3940 6810 4000 6890
rect 3800 6750 4000 6810
rect 4200 6890 4400 6950
rect 4200 6810 4260 6890
rect 4340 6810 4400 6890
rect 4200 6750 4400 6810
rect 4600 6890 4800 6950
rect 4600 6810 4660 6890
rect 4740 6810 4800 6890
rect 4600 6750 4800 6810
rect 5000 6890 5200 6950
rect 5000 6810 5060 6890
rect 5140 6810 5200 6890
rect 5000 6750 5200 6810
rect 5400 6890 5600 6950
rect 5400 6810 5460 6890
rect 5540 6810 5600 6890
rect 5400 6750 5600 6810
rect 5800 6890 6000 6950
rect 5800 6810 5860 6890
rect 5940 6810 6000 6890
rect 5800 6750 6000 6810
rect 6200 6890 6400 6950
rect 6200 6810 6260 6890
rect 6340 6810 6400 6890
rect 6200 6750 6400 6810
rect 6600 6890 6800 6950
rect 6600 6810 6660 6890
rect 6740 6810 6800 6890
rect 6600 6750 6800 6810
rect 7000 6890 7200 6950
rect 7000 6810 7060 6890
rect 7140 6810 7200 6890
rect 7000 6750 7200 6810
rect 7400 6890 7600 6950
rect 7400 6810 7460 6890
rect 7540 6810 7600 6890
rect 7400 6750 7600 6810
rect 7800 6890 8000 6950
rect 7800 6810 7860 6890
rect 7940 6810 8000 6890
rect 7800 6750 8000 6810
rect 8200 6890 8400 6950
rect 8200 6810 8260 6890
rect 8340 6810 8400 6890
rect 8200 6750 8400 6810
rect 8600 6890 8800 6950
rect 8600 6810 8660 6890
rect 8740 6810 8800 6890
rect 8600 6750 8800 6810
rect 9000 6890 9200 6950
rect 9000 6810 9060 6890
rect 9140 6810 9200 6890
rect 9000 6750 9200 6810
rect 9400 6890 9600 6950
rect 9400 6810 9460 6890
rect 9540 6810 9600 6890
rect 9400 6750 9600 6810
rect 9800 6890 10000 6950
rect 9800 6810 9860 6890
rect 9940 6810 10000 6890
rect 9800 6750 10000 6810
rect 2200 6490 2400 6550
rect 2200 6410 2260 6490
rect 2340 6410 2400 6490
rect 2200 6350 2400 6410
rect 2600 6490 2800 6550
rect 2600 6410 2660 6490
rect 2740 6410 2800 6490
rect 2600 6350 2800 6410
rect 3000 6490 3200 6550
rect 3000 6410 3060 6490
rect 3140 6410 3200 6490
rect 3000 6350 3200 6410
rect 3400 6490 3600 6550
rect 3400 6410 3460 6490
rect 3540 6410 3600 6490
rect 3400 6350 3600 6410
rect 3800 6490 4000 6550
rect 3800 6410 3860 6490
rect 3940 6410 4000 6490
rect 3800 6350 4000 6410
rect 4200 6490 4400 6550
rect 4200 6410 4260 6490
rect 4340 6410 4400 6490
rect 4200 6350 4400 6410
rect 4600 6490 4800 6550
rect 4600 6410 4660 6490
rect 4740 6410 4800 6490
rect 4600 6350 4800 6410
rect 5000 6490 5200 6550
rect 5000 6410 5060 6490
rect 5140 6410 5200 6490
rect 5000 6350 5200 6410
rect 5400 6490 5600 6550
rect 5400 6410 5460 6490
rect 5540 6410 5600 6490
rect 5400 6350 5600 6410
rect 5800 6490 6000 6550
rect 5800 6410 5860 6490
rect 5940 6410 6000 6490
rect 5800 6350 6000 6410
rect 6200 6490 6400 6550
rect 6200 6410 6260 6490
rect 6340 6410 6400 6490
rect 6200 6350 6400 6410
rect 6600 6490 6800 6550
rect 6600 6410 6660 6490
rect 6740 6410 6800 6490
rect 6600 6350 6800 6410
rect 7000 6490 7200 6550
rect 7000 6410 7060 6490
rect 7140 6410 7200 6490
rect 7000 6350 7200 6410
rect 7400 6490 7600 6550
rect 7400 6410 7460 6490
rect 7540 6410 7600 6490
rect 7400 6350 7600 6410
rect 7800 6490 8000 6550
rect 7800 6410 7860 6490
rect 7940 6410 8000 6490
rect 7800 6350 8000 6410
rect 8200 6490 8400 6550
rect 8200 6410 8260 6490
rect 8340 6410 8400 6490
rect 8200 6350 8400 6410
rect 8600 6490 8800 6550
rect 8600 6410 8660 6490
rect 8740 6410 8800 6490
rect 8600 6350 8800 6410
rect 9000 6490 9200 6550
rect 9000 6410 9060 6490
rect 9140 6410 9200 6490
rect 9000 6350 9200 6410
rect 9400 6490 9600 6550
rect 9400 6410 9460 6490
rect 9540 6410 9600 6490
rect 9400 6350 9600 6410
rect 9800 6490 10000 6550
rect 9800 6410 9860 6490
rect 9940 6410 10000 6490
rect 9800 6350 10000 6410
rect 2200 6090 2400 6150
rect 2200 6010 2260 6090
rect 2340 6010 2400 6090
rect 2200 5950 2400 6010
rect 2600 6090 2800 6150
rect 2600 6010 2660 6090
rect 2740 6010 2800 6090
rect 2600 5950 2800 6010
rect 3000 6090 3200 6150
rect 3000 6010 3060 6090
rect 3140 6010 3200 6090
rect 3000 5950 3200 6010
rect 3400 6090 3600 6150
rect 3400 6010 3460 6090
rect 3540 6010 3600 6090
rect 3400 5950 3600 6010
rect 3800 6090 4000 6150
rect 3800 6010 3860 6090
rect 3940 6010 4000 6090
rect 3800 5950 4000 6010
rect 4200 6090 4400 6150
rect 4200 6010 4260 6090
rect 4340 6010 4400 6090
rect 4200 5950 4400 6010
rect 4600 6090 4800 6150
rect 4600 6010 4660 6090
rect 4740 6010 4800 6090
rect 4600 5950 4800 6010
rect 5000 6090 5200 6150
rect 5000 6010 5060 6090
rect 5140 6010 5200 6090
rect 5000 5950 5200 6010
rect 5400 6090 5600 6150
rect 5400 6010 5460 6090
rect 5540 6010 5600 6090
rect 5400 5950 5600 6010
rect 5800 6090 6000 6150
rect 5800 6010 5860 6090
rect 5940 6010 6000 6090
rect 5800 5950 6000 6010
rect 6200 6090 6400 6150
rect 6200 6010 6260 6090
rect 6340 6010 6400 6090
rect 6200 5950 6400 6010
rect 6600 6090 6800 6150
rect 6600 6010 6660 6090
rect 6740 6010 6800 6090
rect 6600 5950 6800 6010
rect 7000 6090 7200 6150
rect 7000 6010 7060 6090
rect 7140 6010 7200 6090
rect 7000 5950 7200 6010
rect 7400 6090 7600 6150
rect 7400 6010 7460 6090
rect 7540 6010 7600 6090
rect 7400 5950 7600 6010
rect 7800 6090 8000 6150
rect 7800 6010 7860 6090
rect 7940 6010 8000 6090
rect 7800 5950 8000 6010
rect 8200 6090 8400 6150
rect 8200 6010 8260 6090
rect 8340 6010 8400 6090
rect 8200 5950 8400 6010
rect 8600 6090 8800 6150
rect 8600 6010 8660 6090
rect 8740 6010 8800 6090
rect 8600 5950 8800 6010
rect 9000 6090 9200 6150
rect 9000 6010 9060 6090
rect 9140 6010 9200 6090
rect 9000 5950 9200 6010
rect 9400 6090 9600 6150
rect 9400 6010 9460 6090
rect 9540 6010 9600 6090
rect 9400 5950 9600 6010
rect 9800 6090 10000 6150
rect 9800 6010 9860 6090
rect 9940 6010 10000 6090
rect 9800 5950 10000 6010
rect 2200 5690 2400 5750
rect 2200 5610 2260 5690
rect 2340 5610 2400 5690
rect 2200 5550 2400 5610
rect 2600 5690 2800 5750
rect 2600 5610 2660 5690
rect 2740 5610 2800 5690
rect 2600 5550 2800 5610
rect 3000 5690 3200 5750
rect 3000 5610 3060 5690
rect 3140 5610 3200 5690
rect 3000 5550 3200 5610
rect 3400 5690 3600 5750
rect 3400 5610 3460 5690
rect 3540 5610 3600 5690
rect 3400 5550 3600 5610
rect 3800 5690 4000 5750
rect 3800 5610 3860 5690
rect 3940 5610 4000 5690
rect 3800 5550 4000 5610
rect 4200 5690 4400 5750
rect 4200 5610 4260 5690
rect 4340 5610 4400 5690
rect 4200 5550 4400 5610
rect 4600 5690 4800 5750
rect 4600 5610 4660 5690
rect 4740 5610 4800 5690
rect 4600 5550 4800 5610
rect 5000 5690 5200 5750
rect 5000 5610 5060 5690
rect 5140 5610 5200 5690
rect 5000 5550 5200 5610
rect 5400 5690 5600 5750
rect 5400 5610 5460 5690
rect 5540 5610 5600 5690
rect 5400 5550 5600 5610
rect 5800 5690 6000 5750
rect 5800 5610 5860 5690
rect 5940 5610 6000 5690
rect 5800 5550 6000 5610
rect 6200 5690 6400 5750
rect 6200 5610 6260 5690
rect 6340 5610 6400 5690
rect 6200 5550 6400 5610
rect 6600 5690 6800 5750
rect 6600 5610 6660 5690
rect 6740 5610 6800 5690
rect 6600 5550 6800 5610
rect 7000 5690 7200 5750
rect 7000 5610 7060 5690
rect 7140 5610 7200 5690
rect 7000 5550 7200 5610
rect 7400 5690 7600 5750
rect 7400 5610 7460 5690
rect 7540 5610 7600 5690
rect 7400 5550 7600 5610
rect 7800 5690 8000 5750
rect 7800 5610 7860 5690
rect 7940 5610 8000 5690
rect 7800 5550 8000 5610
rect 8200 5690 8400 5750
rect 8200 5610 8260 5690
rect 8340 5610 8400 5690
rect 8200 5550 8400 5610
rect 8600 5690 8800 5750
rect 8600 5610 8660 5690
rect 8740 5610 8800 5690
rect 8600 5550 8800 5610
rect 9000 5690 9200 5750
rect 9000 5610 9060 5690
rect 9140 5610 9200 5690
rect 9000 5550 9200 5610
rect 9400 5690 9600 5750
rect 9400 5610 9460 5690
rect 9540 5610 9600 5690
rect 9400 5550 9600 5610
rect 9800 5690 10000 5750
rect 9800 5610 9860 5690
rect 9940 5610 10000 5690
rect 9800 5550 10000 5610
rect 2200 5290 2400 5350
rect 2200 5210 2260 5290
rect 2340 5210 2400 5290
rect 2200 5150 2400 5210
rect 2600 5290 2800 5350
rect 2600 5210 2660 5290
rect 2740 5210 2800 5290
rect 2600 5150 2800 5210
rect 3000 5290 3200 5350
rect 3000 5210 3060 5290
rect 3140 5210 3200 5290
rect 3000 5150 3200 5210
rect 3400 5290 3600 5350
rect 3400 5210 3460 5290
rect 3540 5210 3600 5290
rect 3400 5150 3600 5210
rect 3800 5290 4000 5350
rect 3800 5210 3860 5290
rect 3940 5210 4000 5290
rect 3800 5150 4000 5210
rect 4200 5290 4400 5350
rect 4200 5210 4260 5290
rect 4340 5210 4400 5290
rect 4200 5150 4400 5210
rect 4600 5290 4800 5350
rect 4600 5210 4660 5290
rect 4740 5210 4800 5290
rect 4600 5150 4800 5210
rect 5000 5290 5200 5350
rect 5000 5210 5060 5290
rect 5140 5210 5200 5290
rect 5000 5150 5200 5210
rect 5400 5290 5600 5350
rect 5400 5210 5460 5290
rect 5540 5210 5600 5290
rect 5400 5150 5600 5210
rect 5800 5290 6000 5350
rect 5800 5210 5860 5290
rect 5940 5210 6000 5290
rect 5800 5150 6000 5210
rect 6200 5290 6400 5350
rect 6200 5210 6260 5290
rect 6340 5210 6400 5290
rect 6200 5150 6400 5210
rect 6600 5290 6800 5350
rect 6600 5210 6660 5290
rect 6740 5210 6800 5290
rect 6600 5150 6800 5210
rect 7000 5290 7200 5350
rect 7000 5210 7060 5290
rect 7140 5210 7200 5290
rect 7000 5150 7200 5210
rect 7400 5290 7600 5350
rect 7400 5210 7460 5290
rect 7540 5210 7600 5290
rect 7400 5150 7600 5210
rect 7800 5290 8000 5350
rect 7800 5210 7860 5290
rect 7940 5210 8000 5290
rect 7800 5150 8000 5210
rect 8200 5290 8400 5350
rect 8200 5210 8260 5290
rect 8340 5210 8400 5290
rect 8200 5150 8400 5210
rect 8600 5290 8800 5350
rect 8600 5210 8660 5290
rect 8740 5210 8800 5290
rect 8600 5150 8800 5210
rect 9000 5290 9200 5350
rect 9000 5210 9060 5290
rect 9140 5210 9200 5290
rect 9000 5150 9200 5210
rect 9400 5290 9600 5350
rect 9400 5210 9460 5290
rect 9540 5210 9600 5290
rect 9400 5150 9600 5210
rect 9800 5290 10000 5350
rect 9800 5210 9860 5290
rect 9940 5210 10000 5290
rect 9800 5150 10000 5210
rect 2200 4890 2400 4950
rect 2200 4810 2260 4890
rect 2340 4810 2400 4890
rect 2200 4750 2400 4810
rect 2600 4890 2800 4950
rect 2600 4810 2660 4890
rect 2740 4810 2800 4890
rect 2600 4750 2800 4810
rect 3000 4890 3200 4950
rect 3000 4810 3060 4890
rect 3140 4810 3200 4890
rect 3000 4750 3200 4810
rect 3400 4890 3600 4950
rect 3400 4810 3460 4890
rect 3540 4810 3600 4890
rect 3400 4750 3600 4810
rect 3800 4890 4000 4950
rect 3800 4810 3860 4890
rect 3940 4810 4000 4890
rect 3800 4750 4000 4810
rect 4200 4890 4400 4950
rect 4200 4810 4260 4890
rect 4340 4810 4400 4890
rect 4200 4750 4400 4810
rect 4600 4890 4800 4950
rect 4600 4810 4660 4890
rect 4740 4810 4800 4890
rect 4600 4750 4800 4810
rect 5000 4890 5200 4950
rect 5000 4810 5060 4890
rect 5140 4810 5200 4890
rect 5000 4750 5200 4810
rect 5400 4890 5600 4950
rect 5400 4810 5460 4890
rect 5540 4810 5600 4890
rect 5400 4750 5600 4810
rect 5800 4890 6000 4950
rect 5800 4810 5860 4890
rect 5940 4810 6000 4890
rect 5800 4750 6000 4810
rect 6200 4890 6400 4950
rect 6200 4810 6260 4890
rect 6340 4810 6400 4890
rect 6200 4750 6400 4810
rect 6600 4890 6800 4950
rect 6600 4810 6660 4890
rect 6740 4810 6800 4890
rect 6600 4750 6800 4810
rect 7000 4890 7200 4950
rect 7000 4810 7060 4890
rect 7140 4810 7200 4890
rect 7000 4750 7200 4810
rect 7400 4890 7600 4950
rect 7400 4810 7460 4890
rect 7540 4810 7600 4890
rect 7400 4750 7600 4810
rect 7800 4890 8000 4950
rect 7800 4810 7860 4890
rect 7940 4810 8000 4890
rect 7800 4750 8000 4810
rect 8200 4890 8400 4950
rect 8200 4810 8260 4890
rect 8340 4810 8400 4890
rect 8200 4750 8400 4810
rect 8600 4890 8800 4950
rect 8600 4810 8660 4890
rect 8740 4810 8800 4890
rect 8600 4750 8800 4810
rect 9000 4890 9200 4950
rect 9000 4810 9060 4890
rect 9140 4810 9200 4890
rect 9000 4750 9200 4810
rect 9400 4890 9600 4950
rect 9400 4810 9460 4890
rect 9540 4810 9600 4890
rect 9400 4750 9600 4810
rect 9800 4890 10000 4950
rect 9800 4810 9860 4890
rect 9940 4810 10000 4890
rect 9800 4750 10000 4810
rect 2200 4490 2400 4550
rect 2200 4410 2260 4490
rect 2340 4410 2400 4490
rect 2200 4350 2400 4410
rect 2600 4490 2800 4550
rect 2600 4410 2660 4490
rect 2740 4410 2800 4490
rect 2600 4350 2800 4410
rect 3000 4490 3200 4550
rect 3000 4410 3060 4490
rect 3140 4410 3200 4490
rect 3000 4350 3200 4410
rect 3400 4490 3600 4550
rect 3400 4410 3460 4490
rect 3540 4410 3600 4490
rect 3400 4350 3600 4410
rect 3800 4490 4000 4550
rect 3800 4410 3860 4490
rect 3940 4410 4000 4490
rect 3800 4350 4000 4410
rect 4200 4490 4400 4550
rect 4200 4410 4260 4490
rect 4340 4410 4400 4490
rect 4200 4350 4400 4410
rect 4600 4490 4800 4550
rect 4600 4410 4660 4490
rect 4740 4410 4800 4490
rect 4600 4350 4800 4410
rect 5000 4490 5200 4550
rect 5000 4410 5060 4490
rect 5140 4410 5200 4490
rect 5000 4350 5200 4410
rect 5400 4490 5600 4550
rect 5400 4410 5460 4490
rect 5540 4410 5600 4490
rect 5400 4350 5600 4410
rect 5800 4490 6000 4550
rect 5800 4410 5860 4490
rect 5940 4410 6000 4490
rect 5800 4350 6000 4410
rect 6200 4490 6400 4550
rect 6200 4410 6260 4490
rect 6340 4410 6400 4490
rect 6200 4350 6400 4410
rect 6600 4490 6800 4550
rect 6600 4410 6660 4490
rect 6740 4410 6800 4490
rect 6600 4350 6800 4410
rect 7000 4490 7200 4550
rect 7000 4410 7060 4490
rect 7140 4410 7200 4490
rect 7000 4350 7200 4410
rect 7400 4490 7600 4550
rect 7400 4410 7460 4490
rect 7540 4410 7600 4490
rect 7400 4350 7600 4410
rect 7800 4490 8000 4550
rect 7800 4410 7860 4490
rect 7940 4410 8000 4490
rect 7800 4350 8000 4410
rect 8200 4490 8400 4550
rect 8200 4410 8260 4490
rect 8340 4410 8400 4490
rect 8200 4350 8400 4410
rect 8600 4490 8800 4550
rect 8600 4410 8660 4490
rect 8740 4410 8800 4490
rect 8600 4350 8800 4410
rect 9000 4490 9200 4550
rect 9000 4410 9060 4490
rect 9140 4410 9200 4490
rect 9000 4350 9200 4410
rect 9400 4490 9600 4550
rect 9400 4410 9460 4490
rect 9540 4410 9600 4490
rect 9400 4350 9600 4410
rect 9800 4490 10000 4550
rect 9800 4410 9860 4490
rect 9940 4410 10000 4490
rect 9800 4350 10000 4410
rect 2200 4090 2400 4150
rect 2200 4010 2260 4090
rect 2340 4010 2400 4090
rect 2200 3950 2400 4010
rect 2600 4090 2800 4150
rect 2600 4010 2660 4090
rect 2740 4010 2800 4090
rect 2600 3950 2800 4010
rect 3000 4090 3200 4150
rect 3000 4010 3060 4090
rect 3140 4010 3200 4090
rect 3000 3950 3200 4010
rect 3400 4090 3600 4150
rect 3400 4010 3460 4090
rect 3540 4010 3600 4090
rect 3400 3950 3600 4010
rect 3800 4090 4000 4150
rect 3800 4010 3860 4090
rect 3940 4010 4000 4090
rect 3800 3950 4000 4010
rect 4200 4090 4400 4150
rect 4200 4010 4260 4090
rect 4340 4010 4400 4090
rect 4200 3950 4400 4010
rect 4600 4090 4800 4150
rect 4600 4010 4660 4090
rect 4740 4010 4800 4090
rect 4600 3950 4800 4010
rect 5000 4090 5200 4150
rect 5000 4010 5060 4090
rect 5140 4010 5200 4090
rect 5000 3950 5200 4010
rect 5400 4090 5600 4150
rect 5400 4010 5460 4090
rect 5540 4010 5600 4090
rect 5400 3950 5600 4010
rect 5800 4090 6000 4150
rect 5800 4010 5860 4090
rect 5940 4010 6000 4090
rect 5800 3950 6000 4010
rect 6200 4090 6400 4150
rect 6200 4010 6260 4090
rect 6340 4010 6400 4090
rect 6200 3950 6400 4010
rect 6600 4090 6800 4150
rect 6600 4010 6660 4090
rect 6740 4010 6800 4090
rect 6600 3950 6800 4010
rect 7000 4090 7200 4150
rect 7000 4010 7060 4090
rect 7140 4010 7200 4090
rect 7000 3950 7200 4010
rect 7400 4090 7600 4150
rect 7400 4010 7460 4090
rect 7540 4010 7600 4090
rect 7400 3950 7600 4010
rect 7800 4090 8000 4150
rect 7800 4010 7860 4090
rect 7940 4010 8000 4090
rect 7800 3950 8000 4010
rect 8200 4090 8400 4150
rect 8200 4010 8260 4090
rect 8340 4010 8400 4090
rect 8200 3950 8400 4010
rect 8600 4090 8800 4150
rect 8600 4010 8660 4090
rect 8740 4010 8800 4090
rect 8600 3950 8800 4010
rect 9000 4090 9200 4150
rect 9000 4010 9060 4090
rect 9140 4010 9200 4090
rect 9000 3950 9200 4010
rect 9400 4090 9600 4150
rect 9400 4010 9460 4090
rect 9540 4010 9600 4090
rect 9400 3950 9600 4010
rect 9800 4090 10000 4150
rect 9800 4010 9860 4090
rect 9940 4010 10000 4090
rect 9800 3950 10000 4010
rect 2200 3690 2400 3750
rect 2200 3610 2260 3690
rect 2340 3610 2400 3690
rect 2200 3550 2400 3610
rect 2600 3690 2800 3750
rect 2600 3610 2660 3690
rect 2740 3610 2800 3690
rect 2600 3550 2800 3610
rect 3000 3690 3200 3750
rect 3000 3610 3060 3690
rect 3140 3610 3200 3690
rect 3000 3550 3200 3610
rect 3400 3690 3600 3750
rect 3400 3610 3460 3690
rect 3540 3610 3600 3690
rect 3400 3550 3600 3610
rect 3800 3690 4000 3750
rect 3800 3610 3860 3690
rect 3940 3610 4000 3690
rect 3800 3550 4000 3610
rect 4200 3690 4400 3750
rect 4200 3610 4260 3690
rect 4340 3610 4400 3690
rect 4200 3550 4400 3610
rect 4600 3690 4800 3750
rect 4600 3610 4660 3690
rect 4740 3610 4800 3690
rect 4600 3550 4800 3610
rect 5000 3690 5200 3750
rect 5000 3610 5060 3690
rect 5140 3610 5200 3690
rect 5000 3550 5200 3610
rect 5400 3690 5600 3750
rect 5400 3610 5460 3690
rect 5540 3610 5600 3690
rect 5400 3550 5600 3610
rect 5800 3690 6000 3750
rect 5800 3610 5860 3690
rect 5940 3610 6000 3690
rect 5800 3550 6000 3610
rect 6200 3690 6400 3750
rect 6200 3610 6260 3690
rect 6340 3610 6400 3690
rect 6200 3550 6400 3610
rect 6600 3690 6800 3750
rect 6600 3610 6660 3690
rect 6740 3610 6800 3690
rect 6600 3550 6800 3610
rect 7000 3690 7200 3750
rect 7000 3610 7060 3690
rect 7140 3610 7200 3690
rect 7000 3550 7200 3610
rect 7400 3690 7600 3750
rect 7400 3610 7460 3690
rect 7540 3610 7600 3690
rect 7400 3550 7600 3610
rect 7800 3690 8000 3750
rect 7800 3610 7860 3690
rect 7940 3610 8000 3690
rect 7800 3550 8000 3610
rect 8200 3690 8400 3750
rect 8200 3610 8260 3690
rect 8340 3610 8400 3690
rect 8200 3550 8400 3610
rect 8600 3690 8800 3750
rect 8600 3610 8660 3690
rect 8740 3610 8800 3690
rect 8600 3550 8800 3610
rect 9000 3690 9200 3750
rect 9000 3610 9060 3690
rect 9140 3610 9200 3690
rect 9000 3550 9200 3610
rect 9400 3690 9600 3750
rect 9400 3610 9460 3690
rect 9540 3610 9600 3690
rect 9400 3550 9600 3610
rect 9800 3690 10000 3750
rect 9800 3610 9860 3690
rect 9940 3610 10000 3690
rect 9800 3550 10000 3610
rect 2200 3290 2400 3350
rect 2200 3210 2260 3290
rect 2340 3210 2400 3290
rect 2200 3150 2400 3210
rect 2600 3290 2800 3350
rect 2600 3210 2660 3290
rect 2740 3210 2800 3290
rect 2600 3150 2800 3210
rect 3000 3290 3200 3350
rect 3000 3210 3060 3290
rect 3140 3210 3200 3290
rect 3000 3150 3200 3210
rect 3400 3290 3600 3350
rect 3400 3210 3460 3290
rect 3540 3210 3600 3290
rect 3400 3150 3600 3210
rect 3800 3290 4000 3350
rect 3800 3210 3860 3290
rect 3940 3210 4000 3290
rect 3800 3150 4000 3210
rect 4200 3290 4400 3350
rect 4200 3210 4260 3290
rect 4340 3210 4400 3290
rect 4200 3150 4400 3210
rect 4600 3290 4800 3350
rect 4600 3210 4660 3290
rect 4740 3210 4800 3290
rect 4600 3150 4800 3210
rect 5000 3290 5200 3350
rect 5000 3210 5060 3290
rect 5140 3210 5200 3290
rect 5000 3150 5200 3210
rect 5400 3290 5600 3350
rect 5400 3210 5460 3290
rect 5540 3210 5600 3290
rect 5400 3150 5600 3210
rect 5800 3290 6000 3350
rect 5800 3210 5860 3290
rect 5940 3210 6000 3290
rect 5800 3150 6000 3210
rect 6200 3290 6400 3350
rect 6200 3210 6260 3290
rect 6340 3210 6400 3290
rect 6200 3150 6400 3210
rect 6600 3290 6800 3350
rect 6600 3210 6660 3290
rect 6740 3210 6800 3290
rect 6600 3150 6800 3210
rect 7000 3290 7200 3350
rect 7000 3210 7060 3290
rect 7140 3210 7200 3290
rect 7000 3150 7200 3210
rect 7400 3290 7600 3350
rect 7400 3210 7460 3290
rect 7540 3210 7600 3290
rect 7400 3150 7600 3210
rect 7800 3290 8000 3350
rect 7800 3210 7860 3290
rect 7940 3210 8000 3290
rect 7800 3150 8000 3210
rect 8200 3290 8400 3350
rect 8200 3210 8260 3290
rect 8340 3210 8400 3290
rect 8200 3150 8400 3210
rect 8600 3290 8800 3350
rect 8600 3210 8660 3290
rect 8740 3210 8800 3290
rect 8600 3150 8800 3210
rect 9000 3290 9200 3350
rect 9000 3210 9060 3290
rect 9140 3210 9200 3290
rect 9000 3150 9200 3210
rect 9400 3290 9600 3350
rect 9400 3210 9460 3290
rect 9540 3210 9600 3290
rect 9400 3150 9600 3210
rect 9800 3290 10000 3350
rect 9800 3210 9860 3290
rect 9940 3210 10000 3290
rect 9800 3150 10000 3210
rect 2200 2890 2400 2950
rect 2200 2810 2260 2890
rect 2340 2810 2400 2890
rect 2200 2750 2400 2810
rect 2600 2890 2800 2950
rect 2600 2810 2660 2890
rect 2740 2810 2800 2890
rect 2600 2750 2800 2810
rect 3000 2890 3200 2950
rect 3000 2810 3060 2890
rect 3140 2810 3200 2890
rect 3000 2750 3200 2810
rect 3400 2890 3600 2950
rect 3400 2810 3460 2890
rect 3540 2810 3600 2890
rect 3400 2750 3600 2810
rect 3800 2890 4000 2950
rect 3800 2810 3860 2890
rect 3940 2810 4000 2890
rect 3800 2750 4000 2810
rect 4200 2890 4400 2950
rect 4200 2810 4260 2890
rect 4340 2810 4400 2890
rect 4200 2750 4400 2810
rect 4600 2890 4800 2950
rect 4600 2810 4660 2890
rect 4740 2810 4800 2890
rect 4600 2750 4800 2810
rect 5000 2890 5200 2950
rect 5000 2810 5060 2890
rect 5140 2810 5200 2890
rect 5000 2750 5200 2810
rect 5400 2890 5600 2950
rect 5400 2810 5460 2890
rect 5540 2810 5600 2890
rect 5400 2750 5600 2810
rect 5800 2890 6000 2950
rect 5800 2810 5860 2890
rect 5940 2810 6000 2890
rect 5800 2750 6000 2810
rect 6200 2890 6400 2950
rect 6200 2810 6260 2890
rect 6340 2810 6400 2890
rect 6200 2750 6400 2810
rect 6600 2890 6800 2950
rect 6600 2810 6660 2890
rect 6740 2810 6800 2890
rect 6600 2750 6800 2810
rect 7000 2890 7200 2950
rect 7000 2810 7060 2890
rect 7140 2810 7200 2890
rect 7000 2750 7200 2810
rect 7400 2890 7600 2950
rect 7400 2810 7460 2890
rect 7540 2810 7600 2890
rect 7400 2750 7600 2810
rect 7800 2890 8000 2950
rect 7800 2810 7860 2890
rect 7940 2810 8000 2890
rect 7800 2750 8000 2810
rect 8200 2890 8400 2950
rect 8200 2810 8260 2890
rect 8340 2810 8400 2890
rect 8200 2750 8400 2810
rect 8600 2890 8800 2950
rect 8600 2810 8660 2890
rect 8740 2810 8800 2890
rect 8600 2750 8800 2810
rect 9000 2890 9200 2950
rect 9000 2810 9060 2890
rect 9140 2810 9200 2890
rect 9000 2750 9200 2810
rect 9400 2890 9600 2950
rect 9400 2810 9460 2890
rect 9540 2810 9600 2890
rect 9400 2750 9600 2810
rect 9800 2890 10000 2950
rect 9800 2810 9860 2890
rect 9940 2810 10000 2890
rect 9800 2750 10000 2810
rect 2200 2490 2400 2550
rect 2200 2410 2260 2490
rect 2340 2410 2400 2490
rect 2200 2350 2400 2410
rect 2600 2490 2800 2550
rect 2600 2410 2660 2490
rect 2740 2410 2800 2490
rect 2600 2350 2800 2410
rect 3000 2490 3200 2550
rect 3000 2410 3060 2490
rect 3140 2410 3200 2490
rect 3000 2350 3200 2410
rect 3400 2490 3600 2550
rect 3400 2410 3460 2490
rect 3540 2410 3600 2490
rect 3400 2350 3600 2410
rect 3800 2490 4000 2550
rect 3800 2410 3860 2490
rect 3940 2410 4000 2490
rect 3800 2350 4000 2410
rect 4200 2490 4400 2550
rect 4200 2410 4260 2490
rect 4340 2410 4400 2490
rect 4200 2350 4400 2410
rect 4600 2490 4800 2550
rect 4600 2410 4660 2490
rect 4740 2410 4800 2490
rect 4600 2350 4800 2410
rect 5000 2490 5200 2550
rect 5000 2410 5060 2490
rect 5140 2410 5200 2490
rect 5000 2350 5200 2410
rect 5400 2490 5600 2550
rect 5400 2410 5460 2490
rect 5540 2410 5600 2490
rect 5400 2350 5600 2410
rect 5800 2490 6000 2550
rect 5800 2410 5860 2490
rect 5940 2410 6000 2490
rect 5800 2350 6000 2410
rect 6200 2490 6400 2550
rect 6200 2410 6260 2490
rect 6340 2410 6400 2490
rect 6200 2350 6400 2410
rect 6600 2490 6800 2550
rect 6600 2410 6660 2490
rect 6740 2410 6800 2490
rect 6600 2350 6800 2410
rect 7000 2490 7200 2550
rect 7000 2410 7060 2490
rect 7140 2410 7200 2490
rect 7000 2350 7200 2410
rect 7400 2490 7600 2550
rect 7400 2410 7460 2490
rect 7540 2410 7600 2490
rect 7400 2350 7600 2410
rect 7800 2490 8000 2550
rect 7800 2410 7860 2490
rect 7940 2410 8000 2490
rect 7800 2350 8000 2410
rect 8200 2490 8400 2550
rect 8200 2410 8260 2490
rect 8340 2410 8400 2490
rect 8200 2350 8400 2410
rect 8600 2490 8800 2550
rect 8600 2410 8660 2490
rect 8740 2410 8800 2490
rect 8600 2350 8800 2410
rect 9000 2490 9200 2550
rect 9000 2410 9060 2490
rect 9140 2410 9200 2490
rect 9000 2350 9200 2410
rect 9400 2490 9600 2550
rect 9400 2410 9460 2490
rect 9540 2410 9600 2490
rect 9400 2350 9600 2410
rect 9800 2490 10000 2550
rect 9800 2410 9860 2490
rect 9940 2410 10000 2490
rect 9800 2350 10000 2410
rect 2200 2090 2400 2150
rect 2200 2010 2260 2090
rect 2340 2010 2400 2090
rect 2200 1950 2400 2010
rect 2600 2090 2800 2150
rect 2600 2010 2660 2090
rect 2740 2010 2800 2090
rect 2600 1950 2800 2010
rect 3000 2090 3200 2150
rect 3000 2010 3060 2090
rect 3140 2010 3200 2090
rect 3000 1950 3200 2010
rect 3400 2090 3600 2150
rect 3400 2010 3460 2090
rect 3540 2010 3600 2090
rect 3400 1950 3600 2010
rect 3800 2090 4000 2150
rect 3800 2010 3860 2090
rect 3940 2010 4000 2090
rect 3800 1950 4000 2010
rect 4200 2090 4400 2150
rect 4200 2010 4260 2090
rect 4340 2010 4400 2090
rect 4200 1950 4400 2010
rect 4600 2090 4800 2150
rect 4600 2010 4660 2090
rect 4740 2010 4800 2090
rect 4600 1950 4800 2010
rect 5000 2090 5200 2150
rect 5000 2010 5060 2090
rect 5140 2010 5200 2090
rect 5000 1950 5200 2010
rect 5400 2090 5600 2150
rect 5400 2010 5460 2090
rect 5540 2010 5600 2090
rect 5400 1950 5600 2010
rect 5800 2090 6000 2150
rect 5800 2010 5860 2090
rect 5940 2010 6000 2090
rect 5800 1950 6000 2010
rect 6200 2090 6400 2150
rect 6200 2010 6260 2090
rect 6340 2010 6400 2090
rect 6200 1950 6400 2010
rect 6600 2090 6800 2150
rect 6600 2010 6660 2090
rect 6740 2010 6800 2090
rect 6600 1950 6800 2010
rect 7000 2090 7200 2150
rect 7000 2010 7060 2090
rect 7140 2010 7200 2090
rect 7000 1950 7200 2010
rect 7400 2090 7600 2150
rect 7400 2010 7460 2090
rect 7540 2010 7600 2090
rect 7400 1950 7600 2010
rect 7800 2090 8000 2150
rect 7800 2010 7860 2090
rect 7940 2010 8000 2090
rect 7800 1950 8000 2010
rect 8200 2090 8400 2150
rect 8200 2010 8260 2090
rect 8340 2010 8400 2090
rect 8200 1950 8400 2010
rect 8600 2090 8800 2150
rect 8600 2010 8660 2090
rect 8740 2010 8800 2090
rect 8600 1950 8800 2010
rect 9000 2090 9200 2150
rect 9000 2010 9060 2090
rect 9140 2010 9200 2090
rect 9000 1950 9200 2010
rect 9400 2090 9600 2150
rect 9400 2010 9460 2090
rect 9540 2010 9600 2090
rect 9400 1950 9600 2010
rect 9800 2090 10000 2150
rect 9800 2010 9860 2090
rect 9940 2010 10000 2090
rect 9800 1950 10000 2010
rect 2200 1690 2400 1750
rect 2200 1610 2260 1690
rect 2340 1610 2400 1690
rect 2200 1550 2400 1610
rect 2600 1690 2800 1750
rect 2600 1610 2660 1690
rect 2740 1610 2800 1690
rect 2600 1550 2800 1610
rect 3000 1690 3200 1750
rect 3000 1610 3060 1690
rect 3140 1610 3200 1690
rect 3000 1550 3200 1610
rect 3400 1690 3600 1750
rect 3400 1610 3460 1690
rect 3540 1610 3600 1690
rect 3400 1550 3600 1610
rect 3800 1690 4000 1750
rect 3800 1610 3860 1690
rect 3940 1610 4000 1690
rect 3800 1550 4000 1610
rect 4200 1690 4400 1750
rect 4200 1610 4260 1690
rect 4340 1610 4400 1690
rect 4200 1550 4400 1610
rect 4600 1690 4800 1750
rect 4600 1610 4660 1690
rect 4740 1610 4800 1690
rect 4600 1550 4800 1610
rect 5000 1690 5200 1750
rect 5000 1610 5060 1690
rect 5140 1610 5200 1690
rect 5000 1550 5200 1610
rect 5400 1690 5600 1750
rect 5400 1610 5460 1690
rect 5540 1610 5600 1690
rect 5400 1550 5600 1610
rect 5800 1690 6000 1750
rect 5800 1610 5860 1690
rect 5940 1610 6000 1690
rect 5800 1550 6000 1610
rect 6200 1690 6400 1750
rect 6200 1610 6260 1690
rect 6340 1610 6400 1690
rect 6200 1550 6400 1610
rect 6600 1690 6800 1750
rect 6600 1610 6660 1690
rect 6740 1610 6800 1690
rect 6600 1550 6800 1610
rect 7000 1690 7200 1750
rect 7000 1610 7060 1690
rect 7140 1610 7200 1690
rect 7000 1550 7200 1610
rect 7400 1690 7600 1750
rect 7400 1610 7460 1690
rect 7540 1610 7600 1690
rect 7400 1550 7600 1610
rect 7800 1690 8000 1750
rect 7800 1610 7860 1690
rect 7940 1610 8000 1690
rect 7800 1550 8000 1610
rect 8200 1690 8400 1750
rect 8200 1610 8260 1690
rect 8340 1610 8400 1690
rect 8200 1550 8400 1610
rect 8600 1690 8800 1750
rect 8600 1610 8660 1690
rect 8740 1610 8800 1690
rect 8600 1550 8800 1610
rect 9000 1690 9200 1750
rect 9000 1610 9060 1690
rect 9140 1610 9200 1690
rect 9000 1550 9200 1610
rect 9400 1690 9600 1750
rect 9400 1610 9460 1690
rect 9540 1610 9600 1690
rect 9400 1550 9600 1610
rect 9800 1690 10000 1750
rect 9800 1610 9860 1690
rect 9940 1610 10000 1690
rect 9800 1550 10000 1610
rect 2200 1290 2400 1350
rect 2200 1210 2260 1290
rect 2340 1210 2400 1290
rect 2200 1150 2400 1210
rect 2600 1290 2800 1350
rect 2600 1210 2660 1290
rect 2740 1210 2800 1290
rect 2600 1150 2800 1210
rect 3000 1290 3200 1350
rect 3000 1210 3060 1290
rect 3140 1210 3200 1290
rect 3000 1150 3200 1210
rect 3400 1290 3600 1350
rect 3400 1210 3460 1290
rect 3540 1210 3600 1290
rect 3400 1150 3600 1210
rect 3800 1290 4000 1350
rect 3800 1210 3860 1290
rect 3940 1210 4000 1290
rect 3800 1150 4000 1210
rect 4200 1290 4400 1350
rect 4200 1210 4260 1290
rect 4340 1210 4400 1290
rect 4200 1150 4400 1210
rect 4600 1290 4800 1350
rect 4600 1210 4660 1290
rect 4740 1210 4800 1290
rect 4600 1150 4800 1210
rect 5000 1290 5200 1350
rect 5000 1210 5060 1290
rect 5140 1210 5200 1290
rect 5000 1150 5200 1210
rect 5400 1290 5600 1350
rect 5400 1210 5460 1290
rect 5540 1210 5600 1290
rect 5400 1150 5600 1210
rect 5800 1290 6000 1350
rect 5800 1210 5860 1290
rect 5940 1210 6000 1290
rect 5800 1150 6000 1210
rect 6200 1290 6400 1350
rect 6200 1210 6260 1290
rect 6340 1210 6400 1290
rect 6200 1150 6400 1210
rect 6600 1290 6800 1350
rect 6600 1210 6660 1290
rect 6740 1210 6800 1290
rect 6600 1150 6800 1210
rect 7000 1290 7200 1350
rect 7000 1210 7060 1290
rect 7140 1210 7200 1290
rect 7000 1150 7200 1210
rect 7400 1290 7600 1350
rect 7400 1210 7460 1290
rect 7540 1210 7600 1290
rect 7400 1150 7600 1210
rect 7800 1290 8000 1350
rect 7800 1210 7860 1290
rect 7940 1210 8000 1290
rect 7800 1150 8000 1210
rect 8200 1290 8400 1350
rect 8200 1210 8260 1290
rect 8340 1210 8400 1290
rect 8200 1150 8400 1210
rect 8600 1290 8800 1350
rect 8600 1210 8660 1290
rect 8740 1210 8800 1290
rect 8600 1150 8800 1210
rect 9000 1290 9200 1350
rect 9000 1210 9060 1290
rect 9140 1210 9200 1290
rect 9000 1150 9200 1210
rect 9400 1290 9600 1350
rect 9400 1210 9460 1290
rect 9540 1210 9600 1290
rect 9400 1150 9600 1210
rect 9800 1290 10000 1350
rect 9800 1210 9860 1290
rect 9940 1210 10000 1290
rect 9800 1150 10000 1210
rect 2200 890 2400 950
rect 2200 810 2260 890
rect 2340 810 2400 890
rect 2200 750 2400 810
rect 2600 890 2800 950
rect 2600 810 2660 890
rect 2740 810 2800 890
rect 2600 750 2800 810
rect 3000 890 3200 950
rect 3000 810 3060 890
rect 3140 810 3200 890
rect 3000 750 3200 810
rect 3400 890 3600 950
rect 3400 810 3460 890
rect 3540 810 3600 890
rect 3400 750 3600 810
rect 3800 890 4000 950
rect 3800 810 3860 890
rect 3940 810 4000 890
rect 3800 750 4000 810
rect 4200 890 4400 950
rect 4200 810 4260 890
rect 4340 810 4400 890
rect 4200 750 4400 810
rect 4600 890 4800 950
rect 4600 810 4660 890
rect 4740 810 4800 890
rect 4600 750 4800 810
rect 5000 890 5200 950
rect 5000 810 5060 890
rect 5140 810 5200 890
rect 5000 750 5200 810
rect 5400 890 5600 950
rect 5400 810 5460 890
rect 5540 810 5600 890
rect 5400 750 5600 810
rect 5800 890 6000 950
rect 5800 810 5860 890
rect 5940 810 6000 890
rect 5800 750 6000 810
rect 6200 890 6400 950
rect 6200 810 6260 890
rect 6340 810 6400 890
rect 6200 750 6400 810
rect 6600 890 6800 950
rect 6600 810 6660 890
rect 6740 810 6800 890
rect 6600 750 6800 810
rect 7000 890 7200 950
rect 7000 810 7060 890
rect 7140 810 7200 890
rect 7000 750 7200 810
rect 7400 890 7600 950
rect 7400 810 7460 890
rect 7540 810 7600 890
rect 7400 750 7600 810
rect 7800 890 8000 950
rect 7800 810 7860 890
rect 7940 810 8000 890
rect 7800 750 8000 810
rect 8200 890 8400 950
rect 8200 810 8260 890
rect 8340 810 8400 890
rect 8200 750 8400 810
rect 8600 890 8800 950
rect 8600 810 8660 890
rect 8740 810 8800 890
rect 8600 750 8800 810
rect 9000 890 9200 950
rect 9000 810 9060 890
rect 9140 810 9200 890
rect 9000 750 9200 810
rect 9400 890 9600 950
rect 9400 810 9460 890
rect 9540 810 9600 890
rect 9400 750 9600 810
rect 9800 890 10000 950
rect 9800 810 9860 890
rect 9940 810 10000 890
rect 9800 750 10000 810
rect 2200 490 2400 550
rect 2200 410 2260 490
rect 2340 410 2400 490
rect 2200 350 2400 410
rect 2600 490 2800 550
rect 2600 410 2660 490
rect 2740 410 2800 490
rect 2600 350 2800 410
rect 3000 490 3200 550
rect 3000 410 3060 490
rect 3140 410 3200 490
rect 3000 350 3200 410
rect 3400 490 3600 550
rect 3400 410 3460 490
rect 3540 410 3600 490
rect 3400 350 3600 410
rect 3800 490 4000 550
rect 3800 410 3860 490
rect 3940 410 4000 490
rect 3800 350 4000 410
rect 4200 490 4400 550
rect 4200 410 4260 490
rect 4340 410 4400 490
rect 4200 350 4400 410
rect 4600 490 4800 550
rect 4600 410 4660 490
rect 4740 410 4800 490
rect 4600 350 4800 410
rect 5000 490 5200 550
rect 5000 410 5060 490
rect 5140 410 5200 490
rect 5000 350 5200 410
rect 5400 490 5600 550
rect 5400 410 5460 490
rect 5540 410 5600 490
rect 5400 350 5600 410
rect 5800 490 6000 550
rect 5800 410 5860 490
rect 5940 410 6000 490
rect 5800 350 6000 410
rect 6200 490 6400 550
rect 6200 410 6260 490
rect 6340 410 6400 490
rect 6200 350 6400 410
rect 6600 490 6800 550
rect 6600 410 6660 490
rect 6740 410 6800 490
rect 6600 350 6800 410
rect 7000 490 7200 550
rect 7000 410 7060 490
rect 7140 410 7200 490
rect 7000 350 7200 410
rect 7400 490 7600 550
rect 7400 410 7460 490
rect 7540 410 7600 490
rect 7400 350 7600 410
rect 7800 490 8000 550
rect 7800 410 7860 490
rect 7940 410 8000 490
rect 7800 350 8000 410
rect 8200 490 8400 550
rect 8200 410 8260 490
rect 8340 410 8400 490
rect 8200 350 8400 410
rect 8600 490 8800 550
rect 8600 410 8660 490
rect 8740 410 8800 490
rect 8600 350 8800 410
rect 9000 490 9200 550
rect 9000 410 9060 490
rect 9140 410 9200 490
rect 9000 350 9200 410
rect 9400 490 9600 550
rect 9400 410 9460 490
rect 9540 410 9600 490
rect 9400 350 9600 410
rect 9800 490 10000 550
rect 9800 410 9860 490
rect 9940 410 10000 490
rect 9800 350 10000 410
rect 10100 250 10350 8250
rect 1850 0 10350 250
<< m2contact >>
rect 8170 32962 8250 33042
rect 8370 32962 8450 33042
rect 8570 32962 8650 33042
rect 2260 8010 2340 8090
rect 2660 8010 2740 8090
rect 3060 8010 3140 8090
rect 3460 8010 3540 8090
rect 3860 8010 3940 8090
rect 4260 8010 4340 8090
rect 4660 8010 4740 8090
rect 5060 8010 5140 8090
rect 5460 8010 5540 8090
rect 5860 8010 5940 8090
rect 6260 8010 6340 8090
rect 6660 8010 6740 8090
rect 7060 8010 7140 8090
rect 7460 8010 7540 8090
rect 7860 8010 7940 8090
rect 8260 8010 8340 8090
rect 8660 8010 8740 8090
rect 9060 8010 9140 8090
rect 9460 8010 9540 8090
rect 9860 8010 9940 8090
rect 2260 7610 2340 7690
rect 2660 7610 2740 7690
rect 3060 7610 3140 7690
rect 3460 7610 3540 7690
rect 3860 7610 3940 7690
rect 4260 7610 4340 7690
rect 4660 7610 4740 7690
rect 5060 7610 5140 7690
rect 5460 7610 5540 7690
rect 5860 7610 5940 7690
rect 6260 7610 6340 7690
rect 6660 7610 6740 7690
rect 7060 7610 7140 7690
rect 7460 7610 7540 7690
rect 7860 7610 7940 7690
rect 8260 7610 8340 7690
rect 8660 7610 8740 7690
rect 9060 7610 9140 7690
rect 9460 7610 9540 7690
rect 9860 7610 9940 7690
rect 2260 7210 2340 7290
rect 2660 7210 2740 7290
rect 3060 7210 3140 7290
rect 3460 7210 3540 7290
rect 3860 7210 3940 7290
rect 4260 7210 4340 7290
rect 4660 7210 4740 7290
rect 5060 7210 5140 7290
rect 5460 7210 5540 7290
rect 5860 7210 5940 7290
rect 6260 7210 6340 7290
rect 6660 7210 6740 7290
rect 7060 7210 7140 7290
rect 7460 7210 7540 7290
rect 7860 7210 7940 7290
rect 8260 7210 8340 7290
rect 8660 7210 8740 7290
rect 9060 7210 9140 7290
rect 9460 7210 9540 7290
rect 9860 7210 9940 7290
rect 2260 6810 2340 6890
rect 2660 6810 2740 6890
rect 3060 6810 3140 6890
rect 3460 6810 3540 6890
rect 3860 6810 3940 6890
rect 4260 6810 4340 6890
rect 4660 6810 4740 6890
rect 5060 6810 5140 6890
rect 5460 6810 5540 6890
rect 5860 6810 5940 6890
rect 6260 6810 6340 6890
rect 6660 6810 6740 6890
rect 7060 6810 7140 6890
rect 7460 6810 7540 6890
rect 7860 6810 7940 6890
rect 8260 6810 8340 6890
rect 8660 6810 8740 6890
rect 9060 6810 9140 6890
rect 9460 6810 9540 6890
rect 9860 6810 9940 6890
rect 2260 6410 2340 6490
rect 2660 6410 2740 6490
rect 3060 6410 3140 6490
rect 3460 6410 3540 6490
rect 3860 6410 3940 6490
rect 4260 6410 4340 6490
rect 4660 6410 4740 6490
rect 5060 6410 5140 6490
rect 5460 6410 5540 6490
rect 5860 6410 5940 6490
rect 6260 6410 6340 6490
rect 6660 6410 6740 6490
rect 7060 6410 7140 6490
rect 7460 6410 7540 6490
rect 7860 6410 7940 6490
rect 8260 6410 8340 6490
rect 8660 6410 8740 6490
rect 9060 6410 9140 6490
rect 9460 6410 9540 6490
rect 9860 6410 9940 6490
rect 2260 6010 2340 6090
rect 2660 6010 2740 6090
rect 3060 6010 3140 6090
rect 3460 6010 3540 6090
rect 3860 6010 3940 6090
rect 4260 6010 4340 6090
rect 4660 6010 4740 6090
rect 5060 6010 5140 6090
rect 5460 6010 5540 6090
rect 5860 6010 5940 6090
rect 6260 6010 6340 6090
rect 6660 6010 6740 6090
rect 7060 6010 7140 6090
rect 7460 6010 7540 6090
rect 7860 6010 7940 6090
rect 8260 6010 8340 6090
rect 8660 6010 8740 6090
rect 9060 6010 9140 6090
rect 9460 6010 9540 6090
rect 9860 6010 9940 6090
rect 2260 5610 2340 5690
rect 2660 5610 2740 5690
rect 3060 5610 3140 5690
rect 3460 5610 3540 5690
rect 3860 5610 3940 5690
rect 4260 5610 4340 5690
rect 4660 5610 4740 5690
rect 5060 5610 5140 5690
rect 5460 5610 5540 5690
rect 5860 5610 5940 5690
rect 6260 5610 6340 5690
rect 6660 5610 6740 5690
rect 7060 5610 7140 5690
rect 7460 5610 7540 5690
rect 7860 5610 7940 5690
rect 8260 5610 8340 5690
rect 8660 5610 8740 5690
rect 9060 5610 9140 5690
rect 9460 5610 9540 5690
rect 9860 5610 9940 5690
rect 2260 5210 2340 5290
rect 2660 5210 2740 5290
rect 3060 5210 3140 5290
rect 3460 5210 3540 5290
rect 3860 5210 3940 5290
rect 4260 5210 4340 5290
rect 4660 5210 4740 5290
rect 5060 5210 5140 5290
rect 5460 5210 5540 5290
rect 5860 5210 5940 5290
rect 6260 5210 6340 5290
rect 6660 5210 6740 5290
rect 7060 5210 7140 5290
rect 7460 5210 7540 5290
rect 7860 5210 7940 5290
rect 8260 5210 8340 5290
rect 8660 5210 8740 5290
rect 9060 5210 9140 5290
rect 9460 5210 9540 5290
rect 9860 5210 9940 5290
rect 2260 4810 2340 4890
rect 2660 4810 2740 4890
rect 3060 4810 3140 4890
rect 3460 4810 3540 4890
rect 3860 4810 3940 4890
rect 4260 4810 4340 4890
rect 4660 4810 4740 4890
rect 5060 4810 5140 4890
rect 5460 4810 5540 4890
rect 5860 4810 5940 4890
rect 6260 4810 6340 4890
rect 6660 4810 6740 4890
rect 7060 4810 7140 4890
rect 7460 4810 7540 4890
rect 7860 4810 7940 4890
rect 8260 4810 8340 4890
rect 8660 4810 8740 4890
rect 9060 4810 9140 4890
rect 9460 4810 9540 4890
rect 9860 4810 9940 4890
rect 2260 4410 2340 4490
rect 2660 4410 2740 4490
rect 3060 4410 3140 4490
rect 3460 4410 3540 4490
rect 3860 4410 3940 4490
rect 4260 4410 4340 4490
rect 4660 4410 4740 4490
rect 5060 4410 5140 4490
rect 5460 4410 5540 4490
rect 5860 4410 5940 4490
rect 6260 4410 6340 4490
rect 6660 4410 6740 4490
rect 7060 4410 7140 4490
rect 7460 4410 7540 4490
rect 7860 4410 7940 4490
rect 8260 4410 8340 4490
rect 8660 4410 8740 4490
rect 9060 4410 9140 4490
rect 9460 4410 9540 4490
rect 9860 4410 9940 4490
rect 2260 4010 2340 4090
rect 2660 4010 2740 4090
rect 3060 4010 3140 4090
rect 3460 4010 3540 4090
rect 3860 4010 3940 4090
rect 4260 4010 4340 4090
rect 4660 4010 4740 4090
rect 5060 4010 5140 4090
rect 5460 4010 5540 4090
rect 5860 4010 5940 4090
rect 6260 4010 6340 4090
rect 6660 4010 6740 4090
rect 7060 4010 7140 4090
rect 7460 4010 7540 4090
rect 7860 4010 7940 4090
rect 8260 4010 8340 4090
rect 8660 4010 8740 4090
rect 9060 4010 9140 4090
rect 9460 4010 9540 4090
rect 9860 4010 9940 4090
rect 2260 3610 2340 3690
rect 2660 3610 2740 3690
rect 3060 3610 3140 3690
rect 3460 3610 3540 3690
rect 3860 3610 3940 3690
rect 4260 3610 4340 3690
rect 4660 3610 4740 3690
rect 5060 3610 5140 3690
rect 5460 3610 5540 3690
rect 5860 3610 5940 3690
rect 6260 3610 6340 3690
rect 6660 3610 6740 3690
rect 7060 3610 7140 3690
rect 7460 3610 7540 3690
rect 7860 3610 7940 3690
rect 8260 3610 8340 3690
rect 8660 3610 8740 3690
rect 9060 3610 9140 3690
rect 9460 3610 9540 3690
rect 9860 3610 9940 3690
rect 2260 3210 2340 3290
rect 2660 3210 2740 3290
rect 3060 3210 3140 3290
rect 3460 3210 3540 3290
rect 3860 3210 3940 3290
rect 4260 3210 4340 3290
rect 4660 3210 4740 3290
rect 5060 3210 5140 3290
rect 5460 3210 5540 3290
rect 5860 3210 5940 3290
rect 6260 3210 6340 3290
rect 6660 3210 6740 3290
rect 7060 3210 7140 3290
rect 7460 3210 7540 3290
rect 7860 3210 7940 3290
rect 8260 3210 8340 3290
rect 8660 3210 8740 3290
rect 9060 3210 9140 3290
rect 9460 3210 9540 3290
rect 9860 3210 9940 3290
rect 2260 2810 2340 2890
rect 2660 2810 2740 2890
rect 3060 2810 3140 2890
rect 3460 2810 3540 2890
rect 3860 2810 3940 2890
rect 4260 2810 4340 2890
rect 4660 2810 4740 2890
rect 5060 2810 5140 2890
rect 5460 2810 5540 2890
rect 5860 2810 5940 2890
rect 6260 2810 6340 2890
rect 6660 2810 6740 2890
rect 7060 2810 7140 2890
rect 7460 2810 7540 2890
rect 7860 2810 7940 2890
rect 8260 2810 8340 2890
rect 8660 2810 8740 2890
rect 9060 2810 9140 2890
rect 9460 2810 9540 2890
rect 9860 2810 9940 2890
rect 2260 2410 2340 2490
rect 2660 2410 2740 2490
rect 3060 2410 3140 2490
rect 3460 2410 3540 2490
rect 3860 2410 3940 2490
rect 4260 2410 4340 2490
rect 4660 2410 4740 2490
rect 5060 2410 5140 2490
rect 5460 2410 5540 2490
rect 5860 2410 5940 2490
rect 6260 2410 6340 2490
rect 6660 2410 6740 2490
rect 7060 2410 7140 2490
rect 7460 2410 7540 2490
rect 7860 2410 7940 2490
rect 8260 2410 8340 2490
rect 8660 2410 8740 2490
rect 9060 2410 9140 2490
rect 9460 2410 9540 2490
rect 9860 2410 9940 2490
rect 2260 2010 2340 2090
rect 2660 2010 2740 2090
rect 3060 2010 3140 2090
rect 3460 2010 3540 2090
rect 3860 2010 3940 2090
rect 4260 2010 4340 2090
rect 4660 2010 4740 2090
rect 5060 2010 5140 2090
rect 5460 2010 5540 2090
rect 5860 2010 5940 2090
rect 6260 2010 6340 2090
rect 6660 2010 6740 2090
rect 7060 2010 7140 2090
rect 7460 2010 7540 2090
rect 7860 2010 7940 2090
rect 8260 2010 8340 2090
rect 8660 2010 8740 2090
rect 9060 2010 9140 2090
rect 9460 2010 9540 2090
rect 9860 2010 9940 2090
rect 2260 1610 2340 1690
rect 2660 1610 2740 1690
rect 3060 1610 3140 1690
rect 3460 1610 3540 1690
rect 3860 1610 3940 1690
rect 4260 1610 4340 1690
rect 4660 1610 4740 1690
rect 5060 1610 5140 1690
rect 5460 1610 5540 1690
rect 5860 1610 5940 1690
rect 6260 1610 6340 1690
rect 6660 1610 6740 1690
rect 7060 1610 7140 1690
rect 7460 1610 7540 1690
rect 7860 1610 7940 1690
rect 8260 1610 8340 1690
rect 8660 1610 8740 1690
rect 9060 1610 9140 1690
rect 9460 1610 9540 1690
rect 9860 1610 9940 1690
rect 2260 1210 2340 1290
rect 2660 1210 2740 1290
rect 3060 1210 3140 1290
rect 3460 1210 3540 1290
rect 3860 1210 3940 1290
rect 4260 1210 4340 1290
rect 4660 1210 4740 1290
rect 5060 1210 5140 1290
rect 5460 1210 5540 1290
rect 5860 1210 5940 1290
rect 6260 1210 6340 1290
rect 6660 1210 6740 1290
rect 7060 1210 7140 1290
rect 7460 1210 7540 1290
rect 7860 1210 7940 1290
rect 8260 1210 8340 1290
rect 8660 1210 8740 1290
rect 9060 1210 9140 1290
rect 9460 1210 9540 1290
rect 9860 1210 9940 1290
rect 2260 810 2340 890
rect 2660 810 2740 890
rect 3060 810 3140 890
rect 3460 810 3540 890
rect 3860 810 3940 890
rect 4260 810 4340 890
rect 4660 810 4740 890
rect 5060 810 5140 890
rect 5460 810 5540 890
rect 5860 810 5940 890
rect 6260 810 6340 890
rect 6660 810 6740 890
rect 7060 810 7140 890
rect 7460 810 7540 890
rect 7860 810 7940 890
rect 8260 810 8340 890
rect 8660 810 8740 890
rect 9060 810 9140 890
rect 9460 810 9540 890
rect 9860 810 9940 890
rect 2260 410 2340 490
rect 2660 410 2740 490
rect 3060 410 3140 490
rect 3460 410 3540 490
rect 3860 410 3940 490
rect 4260 410 4340 490
rect 4660 410 4740 490
rect 5060 410 5140 490
rect 5460 410 5540 490
rect 5860 410 5940 490
rect 6260 410 6340 490
rect 6660 410 6740 490
rect 7060 410 7140 490
rect 7460 410 7540 490
rect 7860 410 7940 490
rect 8260 410 8340 490
rect 8660 410 8740 490
rect 9060 410 9140 490
rect 9460 410 9540 490
rect 9860 410 9940 490
<< metal2 >>
rect 11400 34310 11720 34450
rect 100 32550 300 34210
rect 11470 33750 11650 34310
rect 9080 33110 9280 33750
rect 9380 33350 9580 33750
rect 9380 33110 9720 33350
rect 9960 33110 10160 33750
rect 10550 33110 10750 33750
rect 11140 33110 11340 33750
rect 11440 33110 11800 33750
rect 8110 33042 8710 33102
rect 100 30250 300 31910
rect 100 20450 500 28250
rect 800 21350 1320 27350
rect 160 16950 500 19950
rect 100 9150 500 16950
rect 810 10050 1310 16050
rect 1420 9850 1960 27350
rect 2060 21350 2580 27350
rect 2070 10050 2570 16050
rect 2680 9850 3220 27350
rect 3320 21350 3840 27350
rect 3330 10050 3830 16050
rect 3940 9850 4480 27350
rect 4580 21350 5100 27350
rect 4590 10050 5090 16050
rect 5200 9850 5740 27350
rect 5840 21350 6360 27350
rect 5850 10050 6350 16050
rect 6460 9850 7000 31253
rect 7560 29750 7925 33005
rect 8110 32962 8170 33042
rect 8250 32962 8370 33042
rect 8450 32962 8570 33042
rect 8650 32962 8710 33042
rect 8110 32235 8710 32962
rect 8940 32810 9420 33010
rect 9180 32235 9320 32810
rect 8110 32010 9320 32235
rect 8110 30853 8631 32010
rect 9180 31650 9320 32010
rect 9520 32230 9720 33110
rect 10120 32810 11480 33010
rect 10590 32230 10730 32810
rect 9520 32010 10730 32230
rect 8800 31450 9420 31650
rect 9520 31350 9720 32010
rect 10590 31650 10730 32010
rect 9820 31450 11500 31650
rect 11600 31350 11800 33110
rect 11900 32550 12100 34210
rect 9080 30710 9280 31350
rect 9380 31110 9720 31350
rect 9380 30710 9580 31110
rect 9960 30710 10160 31350
rect 10560 30710 10760 31350
rect 11160 30710 11360 31350
rect 11460 30710 11800 31350
rect 11900 30250 12100 31910
rect 7560 28730 8810 29750
rect 7100 21350 7620 27350
rect 7110 10050 7610 16050
rect 7720 9850 8260 27350
rect 8360 21350 8880 27350
rect 8370 10050 8870 16050
rect 8980 9850 9520 27350
rect 9620 21350 10140 27350
rect 9630 10050 10130 16050
rect 10240 9850 10780 27350
rect 10880 21350 11400 27350
rect 11600 20450 12100 28250
rect 11600 17450 12040 20450
rect 10890 10050 11390 16050
rect 1420 9150 10780 9850
rect 11600 9150 12100 16950
rect 1850 8250 10350 9150
rect 1850 250 2100 8250
rect 2200 8090 2400 8150
rect 2200 8010 2260 8090
rect 2340 8010 2400 8090
rect 2200 7950 2400 8010
rect 2600 8090 2800 8150
rect 2600 8010 2660 8090
rect 2740 8010 2800 8090
rect 2600 7950 2800 8010
rect 3000 8090 3200 8150
rect 3000 8010 3060 8090
rect 3140 8010 3200 8090
rect 3000 7950 3200 8010
rect 3400 8090 3600 8150
rect 3400 8010 3460 8090
rect 3540 8010 3600 8090
rect 3400 7950 3600 8010
rect 3800 8090 4000 8150
rect 3800 8010 3860 8090
rect 3940 8010 4000 8090
rect 3800 7950 4000 8010
rect 4200 8090 4400 8150
rect 4200 8010 4260 8090
rect 4340 8010 4400 8090
rect 4200 7950 4400 8010
rect 4600 8090 4800 8150
rect 4600 8010 4660 8090
rect 4740 8010 4800 8090
rect 4600 7950 4800 8010
rect 5000 8090 5200 8150
rect 5000 8010 5060 8090
rect 5140 8010 5200 8090
rect 5000 7950 5200 8010
rect 5400 8090 5600 8150
rect 5400 8010 5460 8090
rect 5540 8010 5600 8090
rect 5400 7950 5600 8010
rect 5800 8090 6000 8150
rect 5800 8010 5860 8090
rect 5940 8010 6000 8090
rect 5800 7950 6000 8010
rect 6200 8090 6400 8150
rect 6200 8010 6260 8090
rect 6340 8010 6400 8090
rect 6200 7950 6400 8010
rect 6600 8090 6800 8150
rect 6600 8010 6660 8090
rect 6740 8010 6800 8090
rect 6600 7950 6800 8010
rect 7000 8090 7200 8150
rect 7000 8010 7060 8090
rect 7140 8010 7200 8090
rect 7000 7950 7200 8010
rect 7400 8090 7600 8150
rect 7400 8010 7460 8090
rect 7540 8010 7600 8090
rect 7400 7950 7600 8010
rect 7800 8090 8000 8150
rect 7800 8010 7860 8090
rect 7940 8010 8000 8090
rect 7800 7950 8000 8010
rect 8200 8090 8400 8150
rect 8200 8010 8260 8090
rect 8340 8010 8400 8090
rect 8200 7950 8400 8010
rect 8600 8090 8800 8150
rect 8600 8010 8660 8090
rect 8740 8010 8800 8090
rect 8600 7950 8800 8010
rect 9000 8090 9200 8150
rect 9000 8010 9060 8090
rect 9140 8010 9200 8090
rect 9000 7950 9200 8010
rect 9400 8090 9600 8150
rect 9400 8010 9460 8090
rect 9540 8010 9600 8090
rect 9400 7950 9600 8010
rect 9800 8090 10000 8150
rect 9800 8010 9860 8090
rect 9940 8010 10000 8090
rect 9800 7950 10000 8010
rect 2400 7890 2600 7950
rect 2400 7810 2460 7890
rect 2540 7810 2600 7890
rect 2400 7750 2600 7810
rect 2800 7890 3000 7950
rect 2800 7810 2860 7890
rect 2940 7810 3000 7890
rect 2800 7750 3000 7810
rect 3200 7890 3400 7950
rect 3200 7810 3260 7890
rect 3340 7810 3400 7890
rect 3200 7750 3400 7810
rect 3600 7890 3800 7950
rect 3600 7810 3660 7890
rect 3740 7810 3800 7890
rect 3600 7750 3800 7810
rect 4000 7890 4200 7950
rect 4000 7810 4060 7890
rect 4140 7810 4200 7890
rect 4000 7750 4200 7810
rect 4400 7890 4600 7950
rect 4400 7810 4460 7890
rect 4540 7810 4600 7890
rect 4400 7750 4600 7810
rect 4800 7890 5000 7950
rect 4800 7810 4860 7890
rect 4940 7810 5000 7890
rect 4800 7750 5000 7810
rect 5200 7890 5400 7950
rect 5200 7810 5260 7890
rect 5340 7810 5400 7890
rect 5200 7750 5400 7810
rect 5600 7890 5800 7950
rect 5600 7810 5660 7890
rect 5740 7810 5800 7890
rect 5600 7750 5800 7810
rect 6000 7890 6200 7950
rect 6000 7810 6060 7890
rect 6140 7810 6200 7890
rect 6000 7750 6200 7810
rect 6400 7890 6600 7950
rect 6400 7810 6460 7890
rect 6540 7810 6600 7890
rect 6400 7750 6600 7810
rect 6800 7890 7000 7950
rect 6800 7810 6860 7890
rect 6940 7810 7000 7890
rect 6800 7750 7000 7810
rect 7200 7890 7400 7950
rect 7200 7810 7260 7890
rect 7340 7810 7400 7890
rect 7200 7750 7400 7810
rect 7600 7890 7800 7950
rect 7600 7810 7660 7890
rect 7740 7810 7800 7890
rect 7600 7750 7800 7810
rect 8000 7890 8200 7950
rect 8000 7810 8060 7890
rect 8140 7810 8200 7890
rect 8000 7750 8200 7810
rect 8400 7890 8600 7950
rect 8400 7810 8460 7890
rect 8540 7810 8600 7890
rect 8400 7750 8600 7810
rect 8800 7890 9000 7950
rect 8800 7810 8860 7890
rect 8940 7810 9000 7890
rect 8800 7750 9000 7810
rect 9200 7890 9400 7950
rect 9200 7810 9260 7890
rect 9340 7810 9400 7890
rect 9200 7750 9400 7810
rect 9600 7890 9800 7950
rect 9600 7810 9660 7890
rect 9740 7810 9800 7890
rect 9600 7750 9800 7810
rect 2200 7690 2400 7750
rect 2200 7610 2260 7690
rect 2340 7610 2400 7690
rect 2200 7550 2400 7610
rect 2600 7690 2800 7750
rect 2600 7610 2660 7690
rect 2740 7610 2800 7690
rect 2600 7550 2800 7610
rect 3000 7690 3200 7750
rect 3000 7610 3060 7690
rect 3140 7610 3200 7690
rect 3000 7550 3200 7610
rect 3400 7690 3600 7750
rect 3400 7610 3460 7690
rect 3540 7610 3600 7690
rect 3400 7550 3600 7610
rect 3800 7690 4000 7750
rect 3800 7610 3860 7690
rect 3940 7610 4000 7690
rect 3800 7550 4000 7610
rect 4200 7690 4400 7750
rect 4200 7610 4260 7690
rect 4340 7610 4400 7690
rect 4200 7550 4400 7610
rect 4600 7690 4800 7750
rect 4600 7610 4660 7690
rect 4740 7610 4800 7690
rect 4600 7550 4800 7610
rect 5000 7690 5200 7750
rect 5000 7610 5060 7690
rect 5140 7610 5200 7690
rect 5000 7550 5200 7610
rect 5400 7690 5600 7750
rect 5400 7610 5460 7690
rect 5540 7610 5600 7690
rect 5400 7550 5600 7610
rect 5800 7690 6000 7750
rect 5800 7610 5860 7690
rect 5940 7610 6000 7690
rect 5800 7550 6000 7610
rect 6200 7690 6400 7750
rect 6200 7610 6260 7690
rect 6340 7610 6400 7690
rect 6200 7550 6400 7610
rect 6600 7690 6800 7750
rect 6600 7610 6660 7690
rect 6740 7610 6800 7690
rect 6600 7550 6800 7610
rect 7000 7690 7200 7750
rect 7000 7610 7060 7690
rect 7140 7610 7200 7690
rect 7000 7550 7200 7610
rect 7400 7690 7600 7750
rect 7400 7610 7460 7690
rect 7540 7610 7600 7690
rect 7400 7550 7600 7610
rect 7800 7690 8000 7750
rect 7800 7610 7860 7690
rect 7940 7610 8000 7690
rect 7800 7550 8000 7610
rect 8200 7690 8400 7750
rect 8200 7610 8260 7690
rect 8340 7610 8400 7690
rect 8200 7550 8400 7610
rect 8600 7690 8800 7750
rect 8600 7610 8660 7690
rect 8740 7610 8800 7690
rect 8600 7550 8800 7610
rect 9000 7690 9200 7750
rect 9000 7610 9060 7690
rect 9140 7610 9200 7690
rect 9000 7550 9200 7610
rect 9400 7690 9600 7750
rect 9400 7610 9460 7690
rect 9540 7610 9600 7690
rect 9400 7550 9600 7610
rect 9800 7690 10000 7750
rect 9800 7610 9860 7690
rect 9940 7610 10000 7690
rect 9800 7550 10000 7610
rect 2400 7490 2600 7550
rect 2400 7410 2460 7490
rect 2540 7410 2600 7490
rect 2400 7350 2600 7410
rect 2800 7490 3000 7550
rect 2800 7410 2860 7490
rect 2940 7410 3000 7490
rect 2800 7350 3000 7410
rect 3200 7490 3400 7550
rect 3200 7410 3260 7490
rect 3340 7410 3400 7490
rect 3200 7350 3400 7410
rect 3600 7490 3800 7550
rect 3600 7410 3660 7490
rect 3740 7410 3800 7490
rect 3600 7350 3800 7410
rect 4000 7490 4200 7550
rect 4000 7410 4060 7490
rect 4140 7410 4200 7490
rect 4000 7350 4200 7410
rect 4400 7490 4600 7550
rect 4400 7410 4460 7490
rect 4540 7410 4600 7490
rect 4400 7350 4600 7410
rect 4800 7490 5000 7550
rect 4800 7410 4860 7490
rect 4940 7410 5000 7490
rect 4800 7350 5000 7410
rect 5200 7490 5400 7550
rect 5200 7410 5260 7490
rect 5340 7410 5400 7490
rect 5200 7350 5400 7410
rect 5600 7490 5800 7550
rect 5600 7410 5660 7490
rect 5740 7410 5800 7490
rect 5600 7350 5800 7410
rect 6000 7490 6200 7550
rect 6000 7410 6060 7490
rect 6140 7410 6200 7490
rect 6000 7350 6200 7410
rect 6400 7490 6600 7550
rect 6400 7410 6460 7490
rect 6540 7410 6600 7490
rect 6400 7350 6600 7410
rect 6800 7490 7000 7550
rect 6800 7410 6860 7490
rect 6940 7410 7000 7490
rect 6800 7350 7000 7410
rect 7200 7490 7400 7550
rect 7200 7410 7260 7490
rect 7340 7410 7400 7490
rect 7200 7350 7400 7410
rect 7600 7490 7800 7550
rect 7600 7410 7660 7490
rect 7740 7410 7800 7490
rect 7600 7350 7800 7410
rect 8000 7490 8200 7550
rect 8000 7410 8060 7490
rect 8140 7410 8200 7490
rect 8000 7350 8200 7410
rect 8400 7490 8600 7550
rect 8400 7410 8460 7490
rect 8540 7410 8600 7490
rect 8400 7350 8600 7410
rect 8800 7490 9000 7550
rect 8800 7410 8860 7490
rect 8940 7410 9000 7490
rect 8800 7350 9000 7410
rect 9200 7490 9400 7550
rect 9200 7410 9260 7490
rect 9340 7410 9400 7490
rect 9200 7350 9400 7410
rect 9600 7490 9800 7550
rect 9600 7410 9660 7490
rect 9740 7410 9800 7490
rect 9600 7350 9800 7410
rect 2200 7290 2400 7350
rect 2200 7210 2260 7290
rect 2340 7210 2400 7290
rect 2200 7150 2400 7210
rect 2600 7290 2800 7350
rect 2600 7210 2660 7290
rect 2740 7210 2800 7290
rect 2600 7150 2800 7210
rect 3000 7290 3200 7350
rect 3000 7210 3060 7290
rect 3140 7210 3200 7290
rect 3000 7150 3200 7210
rect 3400 7290 3600 7350
rect 3400 7210 3460 7290
rect 3540 7210 3600 7290
rect 3400 7150 3600 7210
rect 3800 7290 4000 7350
rect 3800 7210 3860 7290
rect 3940 7210 4000 7290
rect 3800 7150 4000 7210
rect 4200 7290 4400 7350
rect 4200 7210 4260 7290
rect 4340 7210 4400 7290
rect 4200 7150 4400 7210
rect 4600 7290 4800 7350
rect 4600 7210 4660 7290
rect 4740 7210 4800 7290
rect 4600 7150 4800 7210
rect 5000 7290 5200 7350
rect 5000 7210 5060 7290
rect 5140 7210 5200 7290
rect 5000 7150 5200 7210
rect 5400 7290 5600 7350
rect 5400 7210 5460 7290
rect 5540 7210 5600 7290
rect 5400 7150 5600 7210
rect 5800 7290 6000 7350
rect 5800 7210 5860 7290
rect 5940 7210 6000 7290
rect 5800 7150 6000 7210
rect 6200 7290 6400 7350
rect 6200 7210 6260 7290
rect 6340 7210 6400 7290
rect 6200 7150 6400 7210
rect 6600 7290 6800 7350
rect 6600 7210 6660 7290
rect 6740 7210 6800 7290
rect 6600 7150 6800 7210
rect 7000 7290 7200 7350
rect 7000 7210 7060 7290
rect 7140 7210 7200 7290
rect 7000 7150 7200 7210
rect 7400 7290 7600 7350
rect 7400 7210 7460 7290
rect 7540 7210 7600 7290
rect 7400 7150 7600 7210
rect 7800 7290 8000 7350
rect 7800 7210 7860 7290
rect 7940 7210 8000 7290
rect 7800 7150 8000 7210
rect 8200 7290 8400 7350
rect 8200 7210 8260 7290
rect 8340 7210 8400 7290
rect 8200 7150 8400 7210
rect 8600 7290 8800 7350
rect 8600 7210 8660 7290
rect 8740 7210 8800 7290
rect 8600 7150 8800 7210
rect 9000 7290 9200 7350
rect 9000 7210 9060 7290
rect 9140 7210 9200 7290
rect 9000 7150 9200 7210
rect 9400 7290 9600 7350
rect 9400 7210 9460 7290
rect 9540 7210 9600 7290
rect 9400 7150 9600 7210
rect 9800 7290 10000 7350
rect 9800 7210 9860 7290
rect 9940 7210 10000 7290
rect 9800 7150 10000 7210
rect 2400 7090 2600 7150
rect 2400 7010 2460 7090
rect 2540 7010 2600 7090
rect 2400 6950 2600 7010
rect 2800 7090 3000 7150
rect 2800 7010 2860 7090
rect 2940 7010 3000 7090
rect 2800 6950 3000 7010
rect 3200 7090 3400 7150
rect 3200 7010 3260 7090
rect 3340 7010 3400 7090
rect 3200 6950 3400 7010
rect 3600 7090 3800 7150
rect 3600 7010 3660 7090
rect 3740 7010 3800 7090
rect 3600 6950 3800 7010
rect 4000 7090 4200 7150
rect 4000 7010 4060 7090
rect 4140 7010 4200 7090
rect 4000 6950 4200 7010
rect 4400 7090 4600 7150
rect 4400 7010 4460 7090
rect 4540 7010 4600 7090
rect 4400 6950 4600 7010
rect 4800 7090 5000 7150
rect 4800 7010 4860 7090
rect 4940 7010 5000 7090
rect 4800 6950 5000 7010
rect 5200 7090 5400 7150
rect 5200 7010 5260 7090
rect 5340 7010 5400 7090
rect 5200 6950 5400 7010
rect 5600 7090 5800 7150
rect 5600 7010 5660 7090
rect 5740 7010 5800 7090
rect 5600 6950 5800 7010
rect 6000 7090 6200 7150
rect 6000 7010 6060 7090
rect 6140 7010 6200 7090
rect 6000 6950 6200 7010
rect 6400 7090 6600 7150
rect 6400 7010 6460 7090
rect 6540 7010 6600 7090
rect 6400 6950 6600 7010
rect 6800 7090 7000 7150
rect 6800 7010 6860 7090
rect 6940 7010 7000 7090
rect 6800 6950 7000 7010
rect 7200 7090 7400 7150
rect 7200 7010 7260 7090
rect 7340 7010 7400 7090
rect 7200 6950 7400 7010
rect 7600 7090 7800 7150
rect 7600 7010 7660 7090
rect 7740 7010 7800 7090
rect 7600 6950 7800 7010
rect 8000 7090 8200 7150
rect 8000 7010 8060 7090
rect 8140 7010 8200 7090
rect 8000 6950 8200 7010
rect 8400 7090 8600 7150
rect 8400 7010 8460 7090
rect 8540 7010 8600 7090
rect 8400 6950 8600 7010
rect 8800 7090 9000 7150
rect 8800 7010 8860 7090
rect 8940 7010 9000 7090
rect 8800 6950 9000 7010
rect 9200 7090 9400 7150
rect 9200 7010 9260 7090
rect 9340 7010 9400 7090
rect 9200 6950 9400 7010
rect 9600 7090 9800 7150
rect 9600 7010 9660 7090
rect 9740 7010 9800 7090
rect 9600 6950 9800 7010
rect 2200 6890 2400 6950
rect 2200 6810 2260 6890
rect 2340 6810 2400 6890
rect 2200 6750 2400 6810
rect 2600 6890 2800 6950
rect 2600 6810 2660 6890
rect 2740 6810 2800 6890
rect 2600 6750 2800 6810
rect 3000 6890 3200 6950
rect 3000 6810 3060 6890
rect 3140 6810 3200 6890
rect 3000 6750 3200 6810
rect 3400 6890 3600 6950
rect 3400 6810 3460 6890
rect 3540 6810 3600 6890
rect 3400 6750 3600 6810
rect 3800 6890 4000 6950
rect 3800 6810 3860 6890
rect 3940 6810 4000 6890
rect 3800 6750 4000 6810
rect 4200 6890 4400 6950
rect 4200 6810 4260 6890
rect 4340 6810 4400 6890
rect 4200 6750 4400 6810
rect 4600 6890 4800 6950
rect 4600 6810 4660 6890
rect 4740 6810 4800 6890
rect 4600 6750 4800 6810
rect 5000 6890 5200 6950
rect 5000 6810 5060 6890
rect 5140 6810 5200 6890
rect 5000 6750 5200 6810
rect 5400 6890 5600 6950
rect 5400 6810 5460 6890
rect 5540 6810 5600 6890
rect 5400 6750 5600 6810
rect 5800 6890 6000 6950
rect 5800 6810 5860 6890
rect 5940 6810 6000 6890
rect 5800 6750 6000 6810
rect 6200 6890 6400 6950
rect 6200 6810 6260 6890
rect 6340 6810 6400 6890
rect 6200 6750 6400 6810
rect 6600 6890 6800 6950
rect 6600 6810 6660 6890
rect 6740 6810 6800 6890
rect 6600 6750 6800 6810
rect 7000 6890 7200 6950
rect 7000 6810 7060 6890
rect 7140 6810 7200 6890
rect 7000 6750 7200 6810
rect 7400 6890 7600 6950
rect 7400 6810 7460 6890
rect 7540 6810 7600 6890
rect 7400 6750 7600 6810
rect 7800 6890 8000 6950
rect 7800 6810 7860 6890
rect 7940 6810 8000 6890
rect 7800 6750 8000 6810
rect 8200 6890 8400 6950
rect 8200 6810 8260 6890
rect 8340 6810 8400 6890
rect 8200 6750 8400 6810
rect 8600 6890 8800 6950
rect 8600 6810 8660 6890
rect 8740 6810 8800 6890
rect 8600 6750 8800 6810
rect 9000 6890 9200 6950
rect 9000 6810 9060 6890
rect 9140 6810 9200 6890
rect 9000 6750 9200 6810
rect 9400 6890 9600 6950
rect 9400 6810 9460 6890
rect 9540 6810 9600 6890
rect 9400 6750 9600 6810
rect 9800 6890 10000 6950
rect 9800 6810 9860 6890
rect 9940 6810 10000 6890
rect 9800 6750 10000 6810
rect 2400 6690 2600 6750
rect 2400 6610 2460 6690
rect 2540 6610 2600 6690
rect 2400 6550 2600 6610
rect 2800 6690 3000 6750
rect 2800 6610 2860 6690
rect 2940 6610 3000 6690
rect 2800 6550 3000 6610
rect 3200 6690 3400 6750
rect 3200 6610 3260 6690
rect 3340 6610 3400 6690
rect 3200 6550 3400 6610
rect 3600 6690 3800 6750
rect 3600 6610 3660 6690
rect 3740 6610 3800 6690
rect 3600 6550 3800 6610
rect 4000 6690 4200 6750
rect 4000 6610 4060 6690
rect 4140 6610 4200 6690
rect 4000 6550 4200 6610
rect 4400 6690 4600 6750
rect 4400 6610 4460 6690
rect 4540 6610 4600 6690
rect 4400 6550 4600 6610
rect 4800 6690 5000 6750
rect 4800 6610 4860 6690
rect 4940 6610 5000 6690
rect 4800 6550 5000 6610
rect 5200 6690 5400 6750
rect 5200 6610 5260 6690
rect 5340 6610 5400 6690
rect 5200 6550 5400 6610
rect 5600 6690 5800 6750
rect 5600 6610 5660 6690
rect 5740 6610 5800 6690
rect 5600 6550 5800 6610
rect 6000 6690 6200 6750
rect 6000 6610 6060 6690
rect 6140 6610 6200 6690
rect 6000 6550 6200 6610
rect 6400 6690 6600 6750
rect 6400 6610 6460 6690
rect 6540 6610 6600 6690
rect 6400 6550 6600 6610
rect 6800 6690 7000 6750
rect 6800 6610 6860 6690
rect 6940 6610 7000 6690
rect 6800 6550 7000 6610
rect 7200 6690 7400 6750
rect 7200 6610 7260 6690
rect 7340 6610 7400 6690
rect 7200 6550 7400 6610
rect 7600 6690 7800 6750
rect 7600 6610 7660 6690
rect 7740 6610 7800 6690
rect 7600 6550 7800 6610
rect 8000 6690 8200 6750
rect 8000 6610 8060 6690
rect 8140 6610 8200 6690
rect 8000 6550 8200 6610
rect 8400 6690 8600 6750
rect 8400 6610 8460 6690
rect 8540 6610 8600 6690
rect 8400 6550 8600 6610
rect 8800 6690 9000 6750
rect 8800 6610 8860 6690
rect 8940 6610 9000 6690
rect 8800 6550 9000 6610
rect 9200 6690 9400 6750
rect 9200 6610 9260 6690
rect 9340 6610 9400 6690
rect 9200 6550 9400 6610
rect 9600 6690 9800 6750
rect 9600 6610 9660 6690
rect 9740 6610 9800 6690
rect 9600 6550 9800 6610
rect 2200 6490 2400 6550
rect 2200 6410 2260 6490
rect 2340 6410 2400 6490
rect 2200 6350 2400 6410
rect 2600 6490 2800 6550
rect 2600 6410 2660 6490
rect 2740 6410 2800 6490
rect 2600 6350 2800 6410
rect 3000 6490 3200 6550
rect 3000 6410 3060 6490
rect 3140 6410 3200 6490
rect 3000 6350 3200 6410
rect 3400 6490 3600 6550
rect 3400 6410 3460 6490
rect 3540 6410 3600 6490
rect 3400 6350 3600 6410
rect 3800 6490 4000 6550
rect 3800 6410 3860 6490
rect 3940 6410 4000 6490
rect 3800 6350 4000 6410
rect 4200 6490 4400 6550
rect 4200 6410 4260 6490
rect 4340 6410 4400 6490
rect 4200 6350 4400 6410
rect 4600 6490 4800 6550
rect 4600 6410 4660 6490
rect 4740 6410 4800 6490
rect 4600 6350 4800 6410
rect 5000 6490 5200 6550
rect 5000 6410 5060 6490
rect 5140 6410 5200 6490
rect 5000 6350 5200 6410
rect 5400 6490 5600 6550
rect 5400 6410 5460 6490
rect 5540 6410 5600 6490
rect 5400 6350 5600 6410
rect 5800 6490 6000 6550
rect 5800 6410 5860 6490
rect 5940 6410 6000 6490
rect 5800 6350 6000 6410
rect 6200 6490 6400 6550
rect 6200 6410 6260 6490
rect 6340 6410 6400 6490
rect 6200 6350 6400 6410
rect 6600 6490 6800 6550
rect 6600 6410 6660 6490
rect 6740 6410 6800 6490
rect 6600 6350 6800 6410
rect 7000 6490 7200 6550
rect 7000 6410 7060 6490
rect 7140 6410 7200 6490
rect 7000 6350 7200 6410
rect 7400 6490 7600 6550
rect 7400 6410 7460 6490
rect 7540 6410 7600 6490
rect 7400 6350 7600 6410
rect 7800 6490 8000 6550
rect 7800 6410 7860 6490
rect 7940 6410 8000 6490
rect 7800 6350 8000 6410
rect 8200 6490 8400 6550
rect 8200 6410 8260 6490
rect 8340 6410 8400 6490
rect 8200 6350 8400 6410
rect 8600 6490 8800 6550
rect 8600 6410 8660 6490
rect 8740 6410 8800 6490
rect 8600 6350 8800 6410
rect 9000 6490 9200 6550
rect 9000 6410 9060 6490
rect 9140 6410 9200 6490
rect 9000 6350 9200 6410
rect 9400 6490 9600 6550
rect 9400 6410 9460 6490
rect 9540 6410 9600 6490
rect 9400 6350 9600 6410
rect 9800 6490 10000 6550
rect 9800 6410 9860 6490
rect 9940 6410 10000 6490
rect 9800 6350 10000 6410
rect 2400 6290 2600 6350
rect 2400 6210 2460 6290
rect 2540 6210 2600 6290
rect 2400 6150 2600 6210
rect 2800 6290 3000 6350
rect 2800 6210 2860 6290
rect 2940 6210 3000 6290
rect 2800 6150 3000 6210
rect 3200 6290 3400 6350
rect 3200 6210 3260 6290
rect 3340 6210 3400 6290
rect 3200 6150 3400 6210
rect 3600 6290 3800 6350
rect 3600 6210 3660 6290
rect 3740 6210 3800 6290
rect 3600 6150 3800 6210
rect 4000 6290 4200 6350
rect 4000 6210 4060 6290
rect 4140 6210 4200 6290
rect 4000 6150 4200 6210
rect 4400 6290 4600 6350
rect 4400 6210 4460 6290
rect 4540 6210 4600 6290
rect 4400 6150 4600 6210
rect 4800 6290 5000 6350
rect 4800 6210 4860 6290
rect 4940 6210 5000 6290
rect 4800 6150 5000 6210
rect 5200 6290 5400 6350
rect 5200 6210 5260 6290
rect 5340 6210 5400 6290
rect 5200 6150 5400 6210
rect 5600 6290 5800 6350
rect 5600 6210 5660 6290
rect 5740 6210 5800 6290
rect 5600 6150 5800 6210
rect 6000 6290 6200 6350
rect 6000 6210 6060 6290
rect 6140 6210 6200 6290
rect 6000 6150 6200 6210
rect 6400 6290 6600 6350
rect 6400 6210 6460 6290
rect 6540 6210 6600 6290
rect 6400 6150 6600 6210
rect 6800 6290 7000 6350
rect 6800 6210 6860 6290
rect 6940 6210 7000 6290
rect 6800 6150 7000 6210
rect 7200 6290 7400 6350
rect 7200 6210 7260 6290
rect 7340 6210 7400 6290
rect 7200 6150 7400 6210
rect 7600 6290 7800 6350
rect 7600 6210 7660 6290
rect 7740 6210 7800 6290
rect 7600 6150 7800 6210
rect 8000 6290 8200 6350
rect 8000 6210 8060 6290
rect 8140 6210 8200 6290
rect 8000 6150 8200 6210
rect 8400 6290 8600 6350
rect 8400 6210 8460 6290
rect 8540 6210 8600 6290
rect 8400 6150 8600 6210
rect 8800 6290 9000 6350
rect 8800 6210 8860 6290
rect 8940 6210 9000 6290
rect 8800 6150 9000 6210
rect 9200 6290 9400 6350
rect 9200 6210 9260 6290
rect 9340 6210 9400 6290
rect 9200 6150 9400 6210
rect 9600 6290 9800 6350
rect 9600 6210 9660 6290
rect 9740 6210 9800 6290
rect 9600 6150 9800 6210
rect 2200 6090 2400 6150
rect 2200 6010 2260 6090
rect 2340 6010 2400 6090
rect 2200 5950 2400 6010
rect 2600 6090 2800 6150
rect 2600 6010 2660 6090
rect 2740 6010 2800 6090
rect 2600 5950 2800 6010
rect 3000 6090 3200 6150
rect 3000 6010 3060 6090
rect 3140 6010 3200 6090
rect 3000 5950 3200 6010
rect 3400 6090 3600 6150
rect 3400 6010 3460 6090
rect 3540 6010 3600 6090
rect 3400 5950 3600 6010
rect 3800 6090 4000 6150
rect 3800 6010 3860 6090
rect 3940 6010 4000 6090
rect 3800 5950 4000 6010
rect 4200 6090 4400 6150
rect 4200 6010 4260 6090
rect 4340 6010 4400 6090
rect 4200 5950 4400 6010
rect 4600 6090 4800 6150
rect 4600 6010 4660 6090
rect 4740 6010 4800 6090
rect 4600 5950 4800 6010
rect 5000 6090 5200 6150
rect 5000 6010 5060 6090
rect 5140 6010 5200 6090
rect 5000 5950 5200 6010
rect 5400 6090 5600 6150
rect 5400 6010 5460 6090
rect 5540 6010 5600 6090
rect 5400 5950 5600 6010
rect 5800 6090 6000 6150
rect 5800 6010 5860 6090
rect 5940 6010 6000 6090
rect 5800 5950 6000 6010
rect 6200 6090 6400 6150
rect 6200 6010 6260 6090
rect 6340 6010 6400 6090
rect 6200 5950 6400 6010
rect 6600 6090 6800 6150
rect 6600 6010 6660 6090
rect 6740 6010 6800 6090
rect 6600 5950 6800 6010
rect 7000 6090 7200 6150
rect 7000 6010 7060 6090
rect 7140 6010 7200 6090
rect 7000 5950 7200 6010
rect 7400 6090 7600 6150
rect 7400 6010 7460 6090
rect 7540 6010 7600 6090
rect 7400 5950 7600 6010
rect 7800 6090 8000 6150
rect 7800 6010 7860 6090
rect 7940 6010 8000 6090
rect 7800 5950 8000 6010
rect 8200 6090 8400 6150
rect 8200 6010 8260 6090
rect 8340 6010 8400 6090
rect 8200 5950 8400 6010
rect 8600 6090 8800 6150
rect 8600 6010 8660 6090
rect 8740 6010 8800 6090
rect 8600 5950 8800 6010
rect 9000 6090 9200 6150
rect 9000 6010 9060 6090
rect 9140 6010 9200 6090
rect 9000 5950 9200 6010
rect 9400 6090 9600 6150
rect 9400 6010 9460 6090
rect 9540 6010 9600 6090
rect 9400 5950 9600 6010
rect 9800 6090 10000 6150
rect 9800 6010 9860 6090
rect 9940 6010 10000 6090
rect 9800 5950 10000 6010
rect 2400 5890 2600 5950
rect 2400 5810 2460 5890
rect 2540 5810 2600 5890
rect 2400 5750 2600 5810
rect 2800 5890 3000 5950
rect 2800 5810 2860 5890
rect 2940 5810 3000 5890
rect 2800 5750 3000 5810
rect 3200 5890 3400 5950
rect 3200 5810 3260 5890
rect 3340 5810 3400 5890
rect 3200 5750 3400 5810
rect 3600 5890 3800 5950
rect 3600 5810 3660 5890
rect 3740 5810 3800 5890
rect 3600 5750 3800 5810
rect 4000 5890 4200 5950
rect 4000 5810 4060 5890
rect 4140 5810 4200 5890
rect 4000 5750 4200 5810
rect 4400 5890 4600 5950
rect 4400 5810 4460 5890
rect 4540 5810 4600 5890
rect 4400 5750 4600 5810
rect 4800 5890 5000 5950
rect 4800 5810 4860 5890
rect 4940 5810 5000 5890
rect 4800 5750 5000 5810
rect 5200 5890 5400 5950
rect 5200 5810 5260 5890
rect 5340 5810 5400 5890
rect 5200 5750 5400 5810
rect 5600 5890 5800 5950
rect 5600 5810 5660 5890
rect 5740 5810 5800 5890
rect 5600 5750 5800 5810
rect 6000 5890 6200 5950
rect 6000 5810 6060 5890
rect 6140 5810 6200 5890
rect 6000 5750 6200 5810
rect 6400 5890 6600 5950
rect 6400 5810 6460 5890
rect 6540 5810 6600 5890
rect 6400 5750 6600 5810
rect 6800 5890 7000 5950
rect 6800 5810 6860 5890
rect 6940 5810 7000 5890
rect 6800 5750 7000 5810
rect 7200 5890 7400 5950
rect 7200 5810 7260 5890
rect 7340 5810 7400 5890
rect 7200 5750 7400 5810
rect 7600 5890 7800 5950
rect 7600 5810 7660 5890
rect 7740 5810 7800 5890
rect 7600 5750 7800 5810
rect 8000 5890 8200 5950
rect 8000 5810 8060 5890
rect 8140 5810 8200 5890
rect 8000 5750 8200 5810
rect 8400 5890 8600 5950
rect 8400 5810 8460 5890
rect 8540 5810 8600 5890
rect 8400 5750 8600 5810
rect 8800 5890 9000 5950
rect 8800 5810 8860 5890
rect 8940 5810 9000 5890
rect 8800 5750 9000 5810
rect 9200 5890 9400 5950
rect 9200 5810 9260 5890
rect 9340 5810 9400 5890
rect 9200 5750 9400 5810
rect 9600 5890 9800 5950
rect 9600 5810 9660 5890
rect 9740 5810 9800 5890
rect 9600 5750 9800 5810
rect 2200 5690 2400 5750
rect 2200 5610 2260 5690
rect 2340 5610 2400 5690
rect 2200 5550 2400 5610
rect 2600 5690 2800 5750
rect 2600 5610 2660 5690
rect 2740 5610 2800 5690
rect 2600 5550 2800 5610
rect 3000 5690 3200 5750
rect 3000 5610 3060 5690
rect 3140 5610 3200 5690
rect 3000 5550 3200 5610
rect 3400 5690 3600 5750
rect 3400 5610 3460 5690
rect 3540 5610 3600 5690
rect 3400 5550 3600 5610
rect 3800 5690 4000 5750
rect 3800 5610 3860 5690
rect 3940 5610 4000 5690
rect 3800 5550 4000 5610
rect 4200 5690 4400 5750
rect 4200 5610 4260 5690
rect 4340 5610 4400 5690
rect 4200 5550 4400 5610
rect 4600 5690 4800 5750
rect 4600 5610 4660 5690
rect 4740 5610 4800 5690
rect 4600 5550 4800 5610
rect 5000 5690 5200 5750
rect 5000 5610 5060 5690
rect 5140 5610 5200 5690
rect 5000 5550 5200 5610
rect 5400 5690 5600 5750
rect 5400 5610 5460 5690
rect 5540 5610 5600 5690
rect 5400 5550 5600 5610
rect 5800 5690 6000 5750
rect 5800 5610 5860 5690
rect 5940 5610 6000 5690
rect 5800 5550 6000 5610
rect 6200 5690 6400 5750
rect 6200 5610 6260 5690
rect 6340 5610 6400 5690
rect 6200 5550 6400 5610
rect 6600 5690 6800 5750
rect 6600 5610 6660 5690
rect 6740 5610 6800 5690
rect 6600 5550 6800 5610
rect 7000 5690 7200 5750
rect 7000 5610 7060 5690
rect 7140 5610 7200 5690
rect 7000 5550 7200 5610
rect 7400 5690 7600 5750
rect 7400 5610 7460 5690
rect 7540 5610 7600 5690
rect 7400 5550 7600 5610
rect 7800 5690 8000 5750
rect 7800 5610 7860 5690
rect 7940 5610 8000 5690
rect 7800 5550 8000 5610
rect 8200 5690 8400 5750
rect 8200 5610 8260 5690
rect 8340 5610 8400 5690
rect 8200 5550 8400 5610
rect 8600 5690 8800 5750
rect 8600 5610 8660 5690
rect 8740 5610 8800 5690
rect 8600 5550 8800 5610
rect 9000 5690 9200 5750
rect 9000 5610 9060 5690
rect 9140 5610 9200 5690
rect 9000 5550 9200 5610
rect 9400 5690 9600 5750
rect 9400 5610 9460 5690
rect 9540 5610 9600 5690
rect 9400 5550 9600 5610
rect 9800 5690 10000 5750
rect 9800 5610 9860 5690
rect 9940 5610 10000 5690
rect 9800 5550 10000 5610
rect 2400 5490 2600 5550
rect 2400 5410 2460 5490
rect 2540 5410 2600 5490
rect 2400 5350 2600 5410
rect 2800 5490 3000 5550
rect 2800 5410 2860 5490
rect 2940 5410 3000 5490
rect 2800 5350 3000 5410
rect 3200 5490 3400 5550
rect 3200 5410 3260 5490
rect 3340 5410 3400 5490
rect 3200 5350 3400 5410
rect 3600 5490 3800 5550
rect 3600 5410 3660 5490
rect 3740 5410 3800 5490
rect 3600 5350 3800 5410
rect 4000 5490 4200 5550
rect 4000 5410 4060 5490
rect 4140 5410 4200 5490
rect 4000 5350 4200 5410
rect 4400 5490 4600 5550
rect 4400 5410 4460 5490
rect 4540 5410 4600 5490
rect 4400 5350 4600 5410
rect 4800 5490 5000 5550
rect 4800 5410 4860 5490
rect 4940 5410 5000 5490
rect 4800 5350 5000 5410
rect 5200 5490 5400 5550
rect 5200 5410 5260 5490
rect 5340 5410 5400 5490
rect 5200 5350 5400 5410
rect 5600 5490 5800 5550
rect 5600 5410 5660 5490
rect 5740 5410 5800 5490
rect 5600 5350 5800 5410
rect 6000 5490 6200 5550
rect 6000 5410 6060 5490
rect 6140 5410 6200 5490
rect 6000 5350 6200 5410
rect 6400 5490 6600 5550
rect 6400 5410 6460 5490
rect 6540 5410 6600 5490
rect 6400 5350 6600 5410
rect 6800 5490 7000 5550
rect 6800 5410 6860 5490
rect 6940 5410 7000 5490
rect 6800 5350 7000 5410
rect 7200 5490 7400 5550
rect 7200 5410 7260 5490
rect 7340 5410 7400 5490
rect 7200 5350 7400 5410
rect 7600 5490 7800 5550
rect 7600 5410 7660 5490
rect 7740 5410 7800 5490
rect 7600 5350 7800 5410
rect 8000 5490 8200 5550
rect 8000 5410 8060 5490
rect 8140 5410 8200 5490
rect 8000 5350 8200 5410
rect 8400 5490 8600 5550
rect 8400 5410 8460 5490
rect 8540 5410 8600 5490
rect 8400 5350 8600 5410
rect 8800 5490 9000 5550
rect 8800 5410 8860 5490
rect 8940 5410 9000 5490
rect 8800 5350 9000 5410
rect 9200 5490 9400 5550
rect 9200 5410 9260 5490
rect 9340 5410 9400 5490
rect 9200 5350 9400 5410
rect 9600 5490 9800 5550
rect 9600 5410 9660 5490
rect 9740 5410 9800 5490
rect 9600 5350 9800 5410
rect 2200 5290 2400 5350
rect 2200 5210 2260 5290
rect 2340 5210 2400 5290
rect 2200 5150 2400 5210
rect 2600 5290 2800 5350
rect 2600 5210 2660 5290
rect 2740 5210 2800 5290
rect 2600 5150 2800 5210
rect 3000 5290 3200 5350
rect 3000 5210 3060 5290
rect 3140 5210 3200 5290
rect 3000 5150 3200 5210
rect 3400 5290 3600 5350
rect 3400 5210 3460 5290
rect 3540 5210 3600 5290
rect 3400 5150 3600 5210
rect 3800 5290 4000 5350
rect 3800 5210 3860 5290
rect 3940 5210 4000 5290
rect 3800 5150 4000 5210
rect 4200 5290 4400 5350
rect 4200 5210 4260 5290
rect 4340 5210 4400 5290
rect 4200 5150 4400 5210
rect 4600 5290 4800 5350
rect 4600 5210 4660 5290
rect 4740 5210 4800 5290
rect 4600 5150 4800 5210
rect 5000 5290 5200 5350
rect 5000 5210 5060 5290
rect 5140 5210 5200 5290
rect 5000 5150 5200 5210
rect 5400 5290 5600 5350
rect 5400 5210 5460 5290
rect 5540 5210 5600 5290
rect 5400 5150 5600 5210
rect 5800 5290 6000 5350
rect 5800 5210 5860 5290
rect 5940 5210 6000 5290
rect 5800 5150 6000 5210
rect 6200 5290 6400 5350
rect 6200 5210 6260 5290
rect 6340 5210 6400 5290
rect 6200 5150 6400 5210
rect 6600 5290 6800 5350
rect 6600 5210 6660 5290
rect 6740 5210 6800 5290
rect 6600 5150 6800 5210
rect 7000 5290 7200 5350
rect 7000 5210 7060 5290
rect 7140 5210 7200 5290
rect 7000 5150 7200 5210
rect 7400 5290 7600 5350
rect 7400 5210 7460 5290
rect 7540 5210 7600 5290
rect 7400 5150 7600 5210
rect 7800 5290 8000 5350
rect 7800 5210 7860 5290
rect 7940 5210 8000 5290
rect 7800 5150 8000 5210
rect 8200 5290 8400 5350
rect 8200 5210 8260 5290
rect 8340 5210 8400 5290
rect 8200 5150 8400 5210
rect 8600 5290 8800 5350
rect 8600 5210 8660 5290
rect 8740 5210 8800 5290
rect 8600 5150 8800 5210
rect 9000 5290 9200 5350
rect 9000 5210 9060 5290
rect 9140 5210 9200 5290
rect 9000 5150 9200 5210
rect 9400 5290 9600 5350
rect 9400 5210 9460 5290
rect 9540 5210 9600 5290
rect 9400 5150 9600 5210
rect 9800 5290 10000 5350
rect 9800 5210 9860 5290
rect 9940 5210 10000 5290
rect 9800 5150 10000 5210
rect 2400 5090 2600 5150
rect 2400 5010 2460 5090
rect 2540 5010 2600 5090
rect 2400 4950 2600 5010
rect 2800 5090 3000 5150
rect 2800 5010 2860 5090
rect 2940 5010 3000 5090
rect 2800 4950 3000 5010
rect 3200 5090 3400 5150
rect 3200 5010 3260 5090
rect 3340 5010 3400 5090
rect 3200 4950 3400 5010
rect 3600 5090 3800 5150
rect 3600 5010 3660 5090
rect 3740 5010 3800 5090
rect 3600 4950 3800 5010
rect 4000 5090 4200 5150
rect 4000 5010 4060 5090
rect 4140 5010 4200 5090
rect 4000 4950 4200 5010
rect 4400 5090 4600 5150
rect 4400 5010 4460 5090
rect 4540 5010 4600 5090
rect 4400 4950 4600 5010
rect 4800 5090 5000 5150
rect 4800 5010 4860 5090
rect 4940 5010 5000 5090
rect 4800 4950 5000 5010
rect 5200 5090 5400 5150
rect 5200 5010 5260 5090
rect 5340 5010 5400 5090
rect 5200 4950 5400 5010
rect 5600 5090 5800 5150
rect 5600 5010 5660 5090
rect 5740 5010 5800 5090
rect 5600 4950 5800 5010
rect 6000 5090 6200 5150
rect 6000 5010 6060 5090
rect 6140 5010 6200 5090
rect 6000 4950 6200 5010
rect 6400 5090 6600 5150
rect 6400 5010 6460 5090
rect 6540 5010 6600 5090
rect 6400 4950 6600 5010
rect 6800 5090 7000 5150
rect 6800 5010 6860 5090
rect 6940 5010 7000 5090
rect 6800 4950 7000 5010
rect 7200 5090 7400 5150
rect 7200 5010 7260 5090
rect 7340 5010 7400 5090
rect 7200 4950 7400 5010
rect 7600 5090 7800 5150
rect 7600 5010 7660 5090
rect 7740 5010 7800 5090
rect 7600 4950 7800 5010
rect 8000 5090 8200 5150
rect 8000 5010 8060 5090
rect 8140 5010 8200 5090
rect 8000 4950 8200 5010
rect 8400 5090 8600 5150
rect 8400 5010 8460 5090
rect 8540 5010 8600 5090
rect 8400 4950 8600 5010
rect 8800 5090 9000 5150
rect 8800 5010 8860 5090
rect 8940 5010 9000 5090
rect 8800 4950 9000 5010
rect 9200 5090 9400 5150
rect 9200 5010 9260 5090
rect 9340 5010 9400 5090
rect 9200 4950 9400 5010
rect 9600 5090 9800 5150
rect 9600 5010 9660 5090
rect 9740 5010 9800 5090
rect 9600 4950 9800 5010
rect 2200 4890 2400 4950
rect 2200 4810 2260 4890
rect 2340 4810 2400 4890
rect 2200 4750 2400 4810
rect 2600 4890 2800 4950
rect 2600 4810 2660 4890
rect 2740 4810 2800 4890
rect 2600 4750 2800 4810
rect 3000 4890 3200 4950
rect 3000 4810 3060 4890
rect 3140 4810 3200 4890
rect 3000 4750 3200 4810
rect 3400 4890 3600 4950
rect 3400 4810 3460 4890
rect 3540 4810 3600 4890
rect 3400 4750 3600 4810
rect 3800 4890 4000 4950
rect 3800 4810 3860 4890
rect 3940 4810 4000 4890
rect 3800 4750 4000 4810
rect 4200 4890 4400 4950
rect 4200 4810 4260 4890
rect 4340 4810 4400 4890
rect 4200 4750 4400 4810
rect 4600 4890 4800 4950
rect 4600 4810 4660 4890
rect 4740 4810 4800 4890
rect 4600 4750 4800 4810
rect 5000 4890 5200 4950
rect 5000 4810 5060 4890
rect 5140 4810 5200 4890
rect 5000 4750 5200 4810
rect 5400 4890 5600 4950
rect 5400 4810 5460 4890
rect 5540 4810 5600 4890
rect 5400 4750 5600 4810
rect 5800 4890 6000 4950
rect 5800 4810 5860 4890
rect 5940 4810 6000 4890
rect 5800 4750 6000 4810
rect 6200 4890 6400 4950
rect 6200 4810 6260 4890
rect 6340 4810 6400 4890
rect 6200 4750 6400 4810
rect 6600 4890 6800 4950
rect 6600 4810 6660 4890
rect 6740 4810 6800 4890
rect 6600 4750 6800 4810
rect 7000 4890 7200 4950
rect 7000 4810 7060 4890
rect 7140 4810 7200 4890
rect 7000 4750 7200 4810
rect 7400 4890 7600 4950
rect 7400 4810 7460 4890
rect 7540 4810 7600 4890
rect 7400 4750 7600 4810
rect 7800 4890 8000 4950
rect 7800 4810 7860 4890
rect 7940 4810 8000 4890
rect 7800 4750 8000 4810
rect 8200 4890 8400 4950
rect 8200 4810 8260 4890
rect 8340 4810 8400 4890
rect 8200 4750 8400 4810
rect 8600 4890 8800 4950
rect 8600 4810 8660 4890
rect 8740 4810 8800 4890
rect 8600 4750 8800 4810
rect 9000 4890 9200 4950
rect 9000 4810 9060 4890
rect 9140 4810 9200 4890
rect 9000 4750 9200 4810
rect 9400 4890 9600 4950
rect 9400 4810 9460 4890
rect 9540 4810 9600 4890
rect 9400 4750 9600 4810
rect 9800 4890 10000 4950
rect 9800 4810 9860 4890
rect 9940 4810 10000 4890
rect 9800 4750 10000 4810
rect 2400 4690 2600 4750
rect 2400 4610 2460 4690
rect 2540 4610 2600 4690
rect 2400 4550 2600 4610
rect 2800 4690 3000 4750
rect 2800 4610 2860 4690
rect 2940 4610 3000 4690
rect 2800 4550 3000 4610
rect 3200 4690 3400 4750
rect 3200 4610 3260 4690
rect 3340 4610 3400 4690
rect 3200 4550 3400 4610
rect 3600 4690 3800 4750
rect 3600 4610 3660 4690
rect 3740 4610 3800 4690
rect 3600 4550 3800 4610
rect 4000 4690 4200 4750
rect 4000 4610 4060 4690
rect 4140 4610 4200 4690
rect 4000 4550 4200 4610
rect 4400 4690 4600 4750
rect 4400 4610 4460 4690
rect 4540 4610 4600 4690
rect 4400 4550 4600 4610
rect 4800 4690 5000 4750
rect 4800 4610 4860 4690
rect 4940 4610 5000 4690
rect 4800 4550 5000 4610
rect 5200 4690 5400 4750
rect 5200 4610 5260 4690
rect 5340 4610 5400 4690
rect 5200 4550 5400 4610
rect 5600 4690 5800 4750
rect 5600 4610 5660 4690
rect 5740 4610 5800 4690
rect 5600 4550 5800 4610
rect 6000 4690 6200 4750
rect 6000 4610 6060 4690
rect 6140 4610 6200 4690
rect 6000 4550 6200 4610
rect 6400 4690 6600 4750
rect 6400 4610 6460 4690
rect 6540 4610 6600 4690
rect 6400 4550 6600 4610
rect 6800 4690 7000 4750
rect 6800 4610 6860 4690
rect 6940 4610 7000 4690
rect 6800 4550 7000 4610
rect 7200 4690 7400 4750
rect 7200 4610 7260 4690
rect 7340 4610 7400 4690
rect 7200 4550 7400 4610
rect 7600 4690 7800 4750
rect 7600 4610 7660 4690
rect 7740 4610 7800 4690
rect 7600 4550 7800 4610
rect 8000 4690 8200 4750
rect 8000 4610 8060 4690
rect 8140 4610 8200 4690
rect 8000 4550 8200 4610
rect 8400 4690 8600 4750
rect 8400 4610 8460 4690
rect 8540 4610 8600 4690
rect 8400 4550 8600 4610
rect 8800 4690 9000 4750
rect 8800 4610 8860 4690
rect 8940 4610 9000 4690
rect 8800 4550 9000 4610
rect 9200 4690 9400 4750
rect 9200 4610 9260 4690
rect 9340 4610 9400 4690
rect 9200 4550 9400 4610
rect 9600 4690 9800 4750
rect 9600 4610 9660 4690
rect 9740 4610 9800 4690
rect 9600 4550 9800 4610
rect 2200 4490 2400 4550
rect 2200 4410 2260 4490
rect 2340 4410 2400 4490
rect 2200 4350 2400 4410
rect 2600 4490 2800 4550
rect 2600 4410 2660 4490
rect 2740 4410 2800 4490
rect 2600 4350 2800 4410
rect 3000 4490 3200 4550
rect 3000 4410 3060 4490
rect 3140 4410 3200 4490
rect 3000 4350 3200 4410
rect 3400 4490 3600 4550
rect 3400 4410 3460 4490
rect 3540 4410 3600 4490
rect 3400 4350 3600 4410
rect 3800 4490 4000 4550
rect 3800 4410 3860 4490
rect 3940 4410 4000 4490
rect 3800 4350 4000 4410
rect 4200 4490 4400 4550
rect 4200 4410 4260 4490
rect 4340 4410 4400 4490
rect 4200 4350 4400 4410
rect 4600 4490 4800 4550
rect 4600 4410 4660 4490
rect 4740 4410 4800 4490
rect 4600 4350 4800 4410
rect 5000 4490 5200 4550
rect 5000 4410 5060 4490
rect 5140 4410 5200 4490
rect 5000 4350 5200 4410
rect 5400 4490 5600 4550
rect 5400 4410 5460 4490
rect 5540 4410 5600 4490
rect 5400 4350 5600 4410
rect 5800 4490 6000 4550
rect 5800 4410 5860 4490
rect 5940 4410 6000 4490
rect 5800 4350 6000 4410
rect 6200 4490 6400 4550
rect 6200 4410 6260 4490
rect 6340 4410 6400 4490
rect 6200 4350 6400 4410
rect 6600 4490 6800 4550
rect 6600 4410 6660 4490
rect 6740 4410 6800 4490
rect 6600 4350 6800 4410
rect 7000 4490 7200 4550
rect 7000 4410 7060 4490
rect 7140 4410 7200 4490
rect 7000 4350 7200 4410
rect 7400 4490 7600 4550
rect 7400 4410 7460 4490
rect 7540 4410 7600 4490
rect 7400 4350 7600 4410
rect 7800 4490 8000 4550
rect 7800 4410 7860 4490
rect 7940 4410 8000 4490
rect 7800 4350 8000 4410
rect 8200 4490 8400 4550
rect 8200 4410 8260 4490
rect 8340 4410 8400 4490
rect 8200 4350 8400 4410
rect 8600 4490 8800 4550
rect 8600 4410 8660 4490
rect 8740 4410 8800 4490
rect 8600 4350 8800 4410
rect 9000 4490 9200 4550
rect 9000 4410 9060 4490
rect 9140 4410 9200 4490
rect 9000 4350 9200 4410
rect 9400 4490 9600 4550
rect 9400 4410 9460 4490
rect 9540 4410 9600 4490
rect 9400 4350 9600 4410
rect 9800 4490 10000 4550
rect 9800 4410 9860 4490
rect 9940 4410 10000 4490
rect 9800 4350 10000 4410
rect 2400 4290 2600 4350
rect 2400 4210 2460 4290
rect 2540 4210 2600 4290
rect 2400 4150 2600 4210
rect 2800 4290 3000 4350
rect 2800 4210 2860 4290
rect 2940 4210 3000 4290
rect 2800 4150 3000 4210
rect 3200 4290 3400 4350
rect 3200 4210 3260 4290
rect 3340 4210 3400 4290
rect 3200 4150 3400 4210
rect 3600 4290 3800 4350
rect 3600 4210 3660 4290
rect 3740 4210 3800 4290
rect 3600 4150 3800 4210
rect 4000 4290 4200 4350
rect 4000 4210 4060 4290
rect 4140 4210 4200 4290
rect 4000 4150 4200 4210
rect 4400 4290 4600 4350
rect 4400 4210 4460 4290
rect 4540 4210 4600 4290
rect 4400 4150 4600 4210
rect 4800 4290 5000 4350
rect 4800 4210 4860 4290
rect 4940 4210 5000 4290
rect 4800 4150 5000 4210
rect 5200 4290 5400 4350
rect 5200 4210 5260 4290
rect 5340 4210 5400 4290
rect 5200 4150 5400 4210
rect 5600 4290 5800 4350
rect 5600 4210 5660 4290
rect 5740 4210 5800 4290
rect 5600 4150 5800 4210
rect 6000 4290 6200 4350
rect 6000 4210 6060 4290
rect 6140 4210 6200 4290
rect 6000 4150 6200 4210
rect 6400 4290 6600 4350
rect 6400 4210 6460 4290
rect 6540 4210 6600 4290
rect 6400 4150 6600 4210
rect 6800 4290 7000 4350
rect 6800 4210 6860 4290
rect 6940 4210 7000 4290
rect 6800 4150 7000 4210
rect 7200 4290 7400 4350
rect 7200 4210 7260 4290
rect 7340 4210 7400 4290
rect 7200 4150 7400 4210
rect 7600 4290 7800 4350
rect 7600 4210 7660 4290
rect 7740 4210 7800 4290
rect 7600 4150 7800 4210
rect 8000 4290 8200 4350
rect 8000 4210 8060 4290
rect 8140 4210 8200 4290
rect 8000 4150 8200 4210
rect 8400 4290 8600 4350
rect 8400 4210 8460 4290
rect 8540 4210 8600 4290
rect 8400 4150 8600 4210
rect 8800 4290 9000 4350
rect 8800 4210 8860 4290
rect 8940 4210 9000 4290
rect 8800 4150 9000 4210
rect 9200 4290 9400 4350
rect 9200 4210 9260 4290
rect 9340 4210 9400 4290
rect 9200 4150 9400 4210
rect 9600 4290 9800 4350
rect 9600 4210 9660 4290
rect 9740 4210 9800 4290
rect 9600 4150 9800 4210
rect 2200 4090 2400 4150
rect 2200 4010 2260 4090
rect 2340 4010 2400 4090
rect 2200 3950 2400 4010
rect 2600 4090 2800 4150
rect 2600 4010 2660 4090
rect 2740 4010 2800 4090
rect 2600 3950 2800 4010
rect 3000 4090 3200 4150
rect 3000 4010 3060 4090
rect 3140 4010 3200 4090
rect 3000 3950 3200 4010
rect 3400 4090 3600 4150
rect 3400 4010 3460 4090
rect 3540 4010 3600 4090
rect 3400 3950 3600 4010
rect 3800 4090 4000 4150
rect 3800 4010 3860 4090
rect 3940 4010 4000 4090
rect 3800 3950 4000 4010
rect 4200 4090 4400 4150
rect 4200 4010 4260 4090
rect 4340 4010 4400 4090
rect 4200 3950 4400 4010
rect 4600 4090 4800 4150
rect 4600 4010 4660 4090
rect 4740 4010 4800 4090
rect 4600 3950 4800 4010
rect 5000 4090 5200 4150
rect 5000 4010 5060 4090
rect 5140 4010 5200 4090
rect 5000 3950 5200 4010
rect 5400 4090 5600 4150
rect 5400 4010 5460 4090
rect 5540 4010 5600 4090
rect 5400 3950 5600 4010
rect 5800 4090 6000 4150
rect 5800 4010 5860 4090
rect 5940 4010 6000 4090
rect 5800 3950 6000 4010
rect 6200 4090 6400 4150
rect 6200 4010 6260 4090
rect 6340 4010 6400 4090
rect 6200 3950 6400 4010
rect 6600 4090 6800 4150
rect 6600 4010 6660 4090
rect 6740 4010 6800 4090
rect 6600 3950 6800 4010
rect 7000 4090 7200 4150
rect 7000 4010 7060 4090
rect 7140 4010 7200 4090
rect 7000 3950 7200 4010
rect 7400 4090 7600 4150
rect 7400 4010 7460 4090
rect 7540 4010 7600 4090
rect 7400 3950 7600 4010
rect 7800 4090 8000 4150
rect 7800 4010 7860 4090
rect 7940 4010 8000 4090
rect 7800 3950 8000 4010
rect 8200 4090 8400 4150
rect 8200 4010 8260 4090
rect 8340 4010 8400 4090
rect 8200 3950 8400 4010
rect 8600 4090 8800 4150
rect 8600 4010 8660 4090
rect 8740 4010 8800 4090
rect 8600 3950 8800 4010
rect 9000 4090 9200 4150
rect 9000 4010 9060 4090
rect 9140 4010 9200 4090
rect 9000 3950 9200 4010
rect 9400 4090 9600 4150
rect 9400 4010 9460 4090
rect 9540 4010 9600 4090
rect 9400 3950 9600 4010
rect 9800 4090 10000 4150
rect 9800 4010 9860 4090
rect 9940 4010 10000 4090
rect 9800 3950 10000 4010
rect 2400 3890 2600 3950
rect 2400 3810 2460 3890
rect 2540 3810 2600 3890
rect 2400 3750 2600 3810
rect 2800 3890 3000 3950
rect 2800 3810 2860 3890
rect 2940 3810 3000 3890
rect 2800 3750 3000 3810
rect 3200 3890 3400 3950
rect 3200 3810 3260 3890
rect 3340 3810 3400 3890
rect 3200 3750 3400 3810
rect 3600 3890 3800 3950
rect 3600 3810 3660 3890
rect 3740 3810 3800 3890
rect 3600 3750 3800 3810
rect 4000 3890 4200 3950
rect 4000 3810 4060 3890
rect 4140 3810 4200 3890
rect 4000 3750 4200 3810
rect 4400 3890 4600 3950
rect 4400 3810 4460 3890
rect 4540 3810 4600 3890
rect 4400 3750 4600 3810
rect 4800 3890 5000 3950
rect 4800 3810 4860 3890
rect 4940 3810 5000 3890
rect 4800 3750 5000 3810
rect 5200 3890 5400 3950
rect 5200 3810 5260 3890
rect 5340 3810 5400 3890
rect 5200 3750 5400 3810
rect 5600 3890 5800 3950
rect 5600 3810 5660 3890
rect 5740 3810 5800 3890
rect 5600 3750 5800 3810
rect 6000 3890 6200 3950
rect 6000 3810 6060 3890
rect 6140 3810 6200 3890
rect 6000 3750 6200 3810
rect 6400 3890 6600 3950
rect 6400 3810 6460 3890
rect 6540 3810 6600 3890
rect 6400 3750 6600 3810
rect 6800 3890 7000 3950
rect 6800 3810 6860 3890
rect 6940 3810 7000 3890
rect 6800 3750 7000 3810
rect 7200 3890 7400 3950
rect 7200 3810 7260 3890
rect 7340 3810 7400 3890
rect 7200 3750 7400 3810
rect 7600 3890 7800 3950
rect 7600 3810 7660 3890
rect 7740 3810 7800 3890
rect 7600 3750 7800 3810
rect 8000 3890 8200 3950
rect 8000 3810 8060 3890
rect 8140 3810 8200 3890
rect 8000 3750 8200 3810
rect 8400 3890 8600 3950
rect 8400 3810 8460 3890
rect 8540 3810 8600 3890
rect 8400 3750 8600 3810
rect 8800 3890 9000 3950
rect 8800 3810 8860 3890
rect 8940 3810 9000 3890
rect 8800 3750 9000 3810
rect 9200 3890 9400 3950
rect 9200 3810 9260 3890
rect 9340 3810 9400 3890
rect 9200 3750 9400 3810
rect 9600 3890 9800 3950
rect 9600 3810 9660 3890
rect 9740 3810 9800 3890
rect 9600 3750 9800 3810
rect 2200 3690 2400 3750
rect 2200 3610 2260 3690
rect 2340 3610 2400 3690
rect 2200 3550 2400 3610
rect 2600 3690 2800 3750
rect 2600 3610 2660 3690
rect 2740 3610 2800 3690
rect 2600 3550 2800 3610
rect 3000 3690 3200 3750
rect 3000 3610 3060 3690
rect 3140 3610 3200 3690
rect 3000 3550 3200 3610
rect 3400 3690 3600 3750
rect 3400 3610 3460 3690
rect 3540 3610 3600 3690
rect 3400 3550 3600 3610
rect 3800 3690 4000 3750
rect 3800 3610 3860 3690
rect 3940 3610 4000 3690
rect 3800 3550 4000 3610
rect 4200 3690 4400 3750
rect 4200 3610 4260 3690
rect 4340 3610 4400 3690
rect 4200 3550 4400 3610
rect 4600 3690 4800 3750
rect 4600 3610 4660 3690
rect 4740 3610 4800 3690
rect 4600 3550 4800 3610
rect 5000 3690 5200 3750
rect 5000 3610 5060 3690
rect 5140 3610 5200 3690
rect 5000 3550 5200 3610
rect 5400 3690 5600 3750
rect 5400 3610 5460 3690
rect 5540 3610 5600 3690
rect 5400 3550 5600 3610
rect 5800 3690 6000 3750
rect 5800 3610 5860 3690
rect 5940 3610 6000 3690
rect 5800 3550 6000 3610
rect 6200 3690 6400 3750
rect 6200 3610 6260 3690
rect 6340 3610 6400 3690
rect 6200 3550 6400 3610
rect 6600 3690 6800 3750
rect 6600 3610 6660 3690
rect 6740 3610 6800 3690
rect 6600 3550 6800 3610
rect 7000 3690 7200 3750
rect 7000 3610 7060 3690
rect 7140 3610 7200 3690
rect 7000 3550 7200 3610
rect 7400 3690 7600 3750
rect 7400 3610 7460 3690
rect 7540 3610 7600 3690
rect 7400 3550 7600 3610
rect 7800 3690 8000 3750
rect 7800 3610 7860 3690
rect 7940 3610 8000 3690
rect 7800 3550 8000 3610
rect 8200 3690 8400 3750
rect 8200 3610 8260 3690
rect 8340 3610 8400 3690
rect 8200 3550 8400 3610
rect 8600 3690 8800 3750
rect 8600 3610 8660 3690
rect 8740 3610 8800 3690
rect 8600 3550 8800 3610
rect 9000 3690 9200 3750
rect 9000 3610 9060 3690
rect 9140 3610 9200 3690
rect 9000 3550 9200 3610
rect 9400 3690 9600 3750
rect 9400 3610 9460 3690
rect 9540 3610 9600 3690
rect 9400 3550 9600 3610
rect 9800 3690 10000 3750
rect 9800 3610 9860 3690
rect 9940 3610 10000 3690
rect 9800 3550 10000 3610
rect 2400 3490 2600 3550
rect 2400 3410 2460 3490
rect 2540 3410 2600 3490
rect 2400 3350 2600 3410
rect 2800 3490 3000 3550
rect 2800 3410 2860 3490
rect 2940 3410 3000 3490
rect 2800 3350 3000 3410
rect 3200 3490 3400 3550
rect 3200 3410 3260 3490
rect 3340 3410 3400 3490
rect 3200 3350 3400 3410
rect 3600 3490 3800 3550
rect 3600 3410 3660 3490
rect 3740 3410 3800 3490
rect 3600 3350 3800 3410
rect 4000 3490 4200 3550
rect 4000 3410 4060 3490
rect 4140 3410 4200 3490
rect 4000 3350 4200 3410
rect 4400 3490 4600 3550
rect 4400 3410 4460 3490
rect 4540 3410 4600 3490
rect 4400 3350 4600 3410
rect 4800 3490 5000 3550
rect 4800 3410 4860 3490
rect 4940 3410 5000 3490
rect 4800 3350 5000 3410
rect 5200 3490 5400 3550
rect 5200 3410 5260 3490
rect 5340 3410 5400 3490
rect 5200 3350 5400 3410
rect 5600 3490 5800 3550
rect 5600 3410 5660 3490
rect 5740 3410 5800 3490
rect 5600 3350 5800 3410
rect 6000 3490 6200 3550
rect 6000 3410 6060 3490
rect 6140 3410 6200 3490
rect 6000 3350 6200 3410
rect 6400 3490 6600 3550
rect 6400 3410 6460 3490
rect 6540 3410 6600 3490
rect 6400 3350 6600 3410
rect 6800 3490 7000 3550
rect 6800 3410 6860 3490
rect 6940 3410 7000 3490
rect 6800 3350 7000 3410
rect 7200 3490 7400 3550
rect 7200 3410 7260 3490
rect 7340 3410 7400 3490
rect 7200 3350 7400 3410
rect 7600 3490 7800 3550
rect 7600 3410 7660 3490
rect 7740 3410 7800 3490
rect 7600 3350 7800 3410
rect 8000 3490 8200 3550
rect 8000 3410 8060 3490
rect 8140 3410 8200 3490
rect 8000 3350 8200 3410
rect 8400 3490 8600 3550
rect 8400 3410 8460 3490
rect 8540 3410 8600 3490
rect 8400 3350 8600 3410
rect 8800 3490 9000 3550
rect 8800 3410 8860 3490
rect 8940 3410 9000 3490
rect 8800 3350 9000 3410
rect 9200 3490 9400 3550
rect 9200 3410 9260 3490
rect 9340 3410 9400 3490
rect 9200 3350 9400 3410
rect 9600 3490 9800 3550
rect 9600 3410 9660 3490
rect 9740 3410 9800 3490
rect 9600 3350 9800 3410
rect 2200 3290 2400 3350
rect 2200 3210 2260 3290
rect 2340 3210 2400 3290
rect 2200 3150 2400 3210
rect 2600 3290 2800 3350
rect 2600 3210 2660 3290
rect 2740 3210 2800 3290
rect 2600 3150 2800 3210
rect 3000 3290 3200 3350
rect 3000 3210 3060 3290
rect 3140 3210 3200 3290
rect 3000 3150 3200 3210
rect 3400 3290 3600 3350
rect 3400 3210 3460 3290
rect 3540 3210 3600 3290
rect 3400 3150 3600 3210
rect 3800 3290 4000 3350
rect 3800 3210 3860 3290
rect 3940 3210 4000 3290
rect 3800 3150 4000 3210
rect 4200 3290 4400 3350
rect 4200 3210 4260 3290
rect 4340 3210 4400 3290
rect 4200 3150 4400 3210
rect 4600 3290 4800 3350
rect 4600 3210 4660 3290
rect 4740 3210 4800 3290
rect 4600 3150 4800 3210
rect 5000 3290 5200 3350
rect 5000 3210 5060 3290
rect 5140 3210 5200 3290
rect 5000 3150 5200 3210
rect 5400 3290 5600 3350
rect 5400 3210 5460 3290
rect 5540 3210 5600 3290
rect 5400 3150 5600 3210
rect 5800 3290 6000 3350
rect 5800 3210 5860 3290
rect 5940 3210 6000 3290
rect 5800 3150 6000 3210
rect 6200 3290 6400 3350
rect 6200 3210 6260 3290
rect 6340 3210 6400 3290
rect 6200 3150 6400 3210
rect 6600 3290 6800 3350
rect 6600 3210 6660 3290
rect 6740 3210 6800 3290
rect 6600 3150 6800 3210
rect 7000 3290 7200 3350
rect 7000 3210 7060 3290
rect 7140 3210 7200 3290
rect 7000 3150 7200 3210
rect 7400 3290 7600 3350
rect 7400 3210 7460 3290
rect 7540 3210 7600 3290
rect 7400 3150 7600 3210
rect 7800 3290 8000 3350
rect 7800 3210 7860 3290
rect 7940 3210 8000 3290
rect 7800 3150 8000 3210
rect 8200 3290 8400 3350
rect 8200 3210 8260 3290
rect 8340 3210 8400 3290
rect 8200 3150 8400 3210
rect 8600 3290 8800 3350
rect 8600 3210 8660 3290
rect 8740 3210 8800 3290
rect 8600 3150 8800 3210
rect 9000 3290 9200 3350
rect 9000 3210 9060 3290
rect 9140 3210 9200 3290
rect 9000 3150 9200 3210
rect 9400 3290 9600 3350
rect 9400 3210 9460 3290
rect 9540 3210 9600 3290
rect 9400 3150 9600 3210
rect 9800 3290 10000 3350
rect 9800 3210 9860 3290
rect 9940 3210 10000 3290
rect 9800 3150 10000 3210
rect 2400 3090 2600 3150
rect 2400 3010 2460 3090
rect 2540 3010 2600 3090
rect 2400 2950 2600 3010
rect 2800 3090 3000 3150
rect 2800 3010 2860 3090
rect 2940 3010 3000 3090
rect 2800 2950 3000 3010
rect 3200 3090 3400 3150
rect 3200 3010 3260 3090
rect 3340 3010 3400 3090
rect 3200 2950 3400 3010
rect 3600 3090 3800 3150
rect 3600 3010 3660 3090
rect 3740 3010 3800 3090
rect 3600 2950 3800 3010
rect 4000 3090 4200 3150
rect 4000 3010 4060 3090
rect 4140 3010 4200 3090
rect 4000 2950 4200 3010
rect 4400 3090 4600 3150
rect 4400 3010 4460 3090
rect 4540 3010 4600 3090
rect 4400 2950 4600 3010
rect 4800 3090 5000 3150
rect 4800 3010 4860 3090
rect 4940 3010 5000 3090
rect 4800 2950 5000 3010
rect 5200 3090 5400 3150
rect 5200 3010 5260 3090
rect 5340 3010 5400 3090
rect 5200 2950 5400 3010
rect 5600 3090 5800 3150
rect 5600 3010 5660 3090
rect 5740 3010 5800 3090
rect 5600 2950 5800 3010
rect 6000 3090 6200 3150
rect 6000 3010 6060 3090
rect 6140 3010 6200 3090
rect 6000 2950 6200 3010
rect 6400 3090 6600 3150
rect 6400 3010 6460 3090
rect 6540 3010 6600 3090
rect 6400 2950 6600 3010
rect 6800 3090 7000 3150
rect 6800 3010 6860 3090
rect 6940 3010 7000 3090
rect 6800 2950 7000 3010
rect 7200 3090 7400 3150
rect 7200 3010 7260 3090
rect 7340 3010 7400 3090
rect 7200 2950 7400 3010
rect 7600 3090 7800 3150
rect 7600 3010 7660 3090
rect 7740 3010 7800 3090
rect 7600 2950 7800 3010
rect 8000 3090 8200 3150
rect 8000 3010 8060 3090
rect 8140 3010 8200 3090
rect 8000 2950 8200 3010
rect 8400 3090 8600 3150
rect 8400 3010 8460 3090
rect 8540 3010 8600 3090
rect 8400 2950 8600 3010
rect 8800 3090 9000 3150
rect 8800 3010 8860 3090
rect 8940 3010 9000 3090
rect 8800 2950 9000 3010
rect 9200 3090 9400 3150
rect 9200 3010 9260 3090
rect 9340 3010 9400 3090
rect 9200 2950 9400 3010
rect 9600 3090 9800 3150
rect 9600 3010 9660 3090
rect 9740 3010 9800 3090
rect 9600 2950 9800 3010
rect 2200 2890 2400 2950
rect 2200 2810 2260 2890
rect 2340 2810 2400 2890
rect 2200 2750 2400 2810
rect 2600 2890 2800 2950
rect 2600 2810 2660 2890
rect 2740 2810 2800 2890
rect 2600 2750 2800 2810
rect 3000 2890 3200 2950
rect 3000 2810 3060 2890
rect 3140 2810 3200 2890
rect 3000 2750 3200 2810
rect 3400 2890 3600 2950
rect 3400 2810 3460 2890
rect 3540 2810 3600 2890
rect 3400 2750 3600 2810
rect 3800 2890 4000 2950
rect 3800 2810 3860 2890
rect 3940 2810 4000 2890
rect 3800 2750 4000 2810
rect 4200 2890 4400 2950
rect 4200 2810 4260 2890
rect 4340 2810 4400 2890
rect 4200 2750 4400 2810
rect 4600 2890 4800 2950
rect 4600 2810 4660 2890
rect 4740 2810 4800 2890
rect 4600 2750 4800 2810
rect 5000 2890 5200 2950
rect 5000 2810 5060 2890
rect 5140 2810 5200 2890
rect 5000 2750 5200 2810
rect 5400 2890 5600 2950
rect 5400 2810 5460 2890
rect 5540 2810 5600 2890
rect 5400 2750 5600 2810
rect 5800 2890 6000 2950
rect 5800 2810 5860 2890
rect 5940 2810 6000 2890
rect 5800 2750 6000 2810
rect 6200 2890 6400 2950
rect 6200 2810 6260 2890
rect 6340 2810 6400 2890
rect 6200 2750 6400 2810
rect 6600 2890 6800 2950
rect 6600 2810 6660 2890
rect 6740 2810 6800 2890
rect 6600 2750 6800 2810
rect 7000 2890 7200 2950
rect 7000 2810 7060 2890
rect 7140 2810 7200 2890
rect 7000 2750 7200 2810
rect 7400 2890 7600 2950
rect 7400 2810 7460 2890
rect 7540 2810 7600 2890
rect 7400 2750 7600 2810
rect 7800 2890 8000 2950
rect 7800 2810 7860 2890
rect 7940 2810 8000 2890
rect 7800 2750 8000 2810
rect 8200 2890 8400 2950
rect 8200 2810 8260 2890
rect 8340 2810 8400 2890
rect 8200 2750 8400 2810
rect 8600 2890 8800 2950
rect 8600 2810 8660 2890
rect 8740 2810 8800 2890
rect 8600 2750 8800 2810
rect 9000 2890 9200 2950
rect 9000 2810 9060 2890
rect 9140 2810 9200 2890
rect 9000 2750 9200 2810
rect 9400 2890 9600 2950
rect 9400 2810 9460 2890
rect 9540 2810 9600 2890
rect 9400 2750 9600 2810
rect 9800 2890 10000 2950
rect 9800 2810 9860 2890
rect 9940 2810 10000 2890
rect 9800 2750 10000 2810
rect 2400 2690 2600 2750
rect 2400 2610 2460 2690
rect 2540 2610 2600 2690
rect 2400 2550 2600 2610
rect 2800 2690 3000 2750
rect 2800 2610 2860 2690
rect 2940 2610 3000 2690
rect 2800 2550 3000 2610
rect 3200 2690 3400 2750
rect 3200 2610 3260 2690
rect 3340 2610 3400 2690
rect 3200 2550 3400 2610
rect 3600 2690 3800 2750
rect 3600 2610 3660 2690
rect 3740 2610 3800 2690
rect 3600 2550 3800 2610
rect 4000 2690 4200 2750
rect 4000 2610 4060 2690
rect 4140 2610 4200 2690
rect 4000 2550 4200 2610
rect 4400 2690 4600 2750
rect 4400 2610 4460 2690
rect 4540 2610 4600 2690
rect 4400 2550 4600 2610
rect 4800 2690 5000 2750
rect 4800 2610 4860 2690
rect 4940 2610 5000 2690
rect 4800 2550 5000 2610
rect 5200 2690 5400 2750
rect 5200 2610 5260 2690
rect 5340 2610 5400 2690
rect 5200 2550 5400 2610
rect 5600 2690 5800 2750
rect 5600 2610 5660 2690
rect 5740 2610 5800 2690
rect 5600 2550 5800 2610
rect 6000 2690 6200 2750
rect 6000 2610 6060 2690
rect 6140 2610 6200 2690
rect 6000 2550 6200 2610
rect 6400 2690 6600 2750
rect 6400 2610 6460 2690
rect 6540 2610 6600 2690
rect 6400 2550 6600 2610
rect 6800 2690 7000 2750
rect 6800 2610 6860 2690
rect 6940 2610 7000 2690
rect 6800 2550 7000 2610
rect 7200 2690 7400 2750
rect 7200 2610 7260 2690
rect 7340 2610 7400 2690
rect 7200 2550 7400 2610
rect 7600 2690 7800 2750
rect 7600 2610 7660 2690
rect 7740 2610 7800 2690
rect 7600 2550 7800 2610
rect 8000 2690 8200 2750
rect 8000 2610 8060 2690
rect 8140 2610 8200 2690
rect 8000 2550 8200 2610
rect 8400 2690 8600 2750
rect 8400 2610 8460 2690
rect 8540 2610 8600 2690
rect 8400 2550 8600 2610
rect 8800 2690 9000 2750
rect 8800 2610 8860 2690
rect 8940 2610 9000 2690
rect 8800 2550 9000 2610
rect 9200 2690 9400 2750
rect 9200 2610 9260 2690
rect 9340 2610 9400 2690
rect 9200 2550 9400 2610
rect 9600 2690 9800 2750
rect 9600 2610 9660 2690
rect 9740 2610 9800 2690
rect 9600 2550 9800 2610
rect 2200 2490 2400 2550
rect 2200 2410 2260 2490
rect 2340 2410 2400 2490
rect 2200 2350 2400 2410
rect 2600 2490 2800 2550
rect 2600 2410 2660 2490
rect 2740 2410 2800 2490
rect 2600 2350 2800 2410
rect 3000 2490 3200 2550
rect 3000 2410 3060 2490
rect 3140 2410 3200 2490
rect 3000 2350 3200 2410
rect 3400 2490 3600 2550
rect 3400 2410 3460 2490
rect 3540 2410 3600 2490
rect 3400 2350 3600 2410
rect 3800 2490 4000 2550
rect 3800 2410 3860 2490
rect 3940 2410 4000 2490
rect 3800 2350 4000 2410
rect 4200 2490 4400 2550
rect 4200 2410 4260 2490
rect 4340 2410 4400 2490
rect 4200 2350 4400 2410
rect 4600 2490 4800 2550
rect 4600 2410 4660 2490
rect 4740 2410 4800 2490
rect 4600 2350 4800 2410
rect 5000 2490 5200 2550
rect 5000 2410 5060 2490
rect 5140 2410 5200 2490
rect 5000 2350 5200 2410
rect 5400 2490 5600 2550
rect 5400 2410 5460 2490
rect 5540 2410 5600 2490
rect 5400 2350 5600 2410
rect 5800 2490 6000 2550
rect 5800 2410 5860 2490
rect 5940 2410 6000 2490
rect 5800 2350 6000 2410
rect 6200 2490 6400 2550
rect 6200 2410 6260 2490
rect 6340 2410 6400 2490
rect 6200 2350 6400 2410
rect 6600 2490 6800 2550
rect 6600 2410 6660 2490
rect 6740 2410 6800 2490
rect 6600 2350 6800 2410
rect 7000 2490 7200 2550
rect 7000 2410 7060 2490
rect 7140 2410 7200 2490
rect 7000 2350 7200 2410
rect 7400 2490 7600 2550
rect 7400 2410 7460 2490
rect 7540 2410 7600 2490
rect 7400 2350 7600 2410
rect 7800 2490 8000 2550
rect 7800 2410 7860 2490
rect 7940 2410 8000 2490
rect 7800 2350 8000 2410
rect 8200 2490 8400 2550
rect 8200 2410 8260 2490
rect 8340 2410 8400 2490
rect 8200 2350 8400 2410
rect 8600 2490 8800 2550
rect 8600 2410 8660 2490
rect 8740 2410 8800 2490
rect 8600 2350 8800 2410
rect 9000 2490 9200 2550
rect 9000 2410 9060 2490
rect 9140 2410 9200 2490
rect 9000 2350 9200 2410
rect 9400 2490 9600 2550
rect 9400 2410 9460 2490
rect 9540 2410 9600 2490
rect 9400 2350 9600 2410
rect 9800 2490 10000 2550
rect 9800 2410 9860 2490
rect 9940 2410 10000 2490
rect 9800 2350 10000 2410
rect 2400 2290 2600 2350
rect 2400 2210 2460 2290
rect 2540 2210 2600 2290
rect 2400 2150 2600 2210
rect 2800 2290 3000 2350
rect 2800 2210 2860 2290
rect 2940 2210 3000 2290
rect 2800 2150 3000 2210
rect 3200 2290 3400 2350
rect 3200 2210 3260 2290
rect 3340 2210 3400 2290
rect 3200 2150 3400 2210
rect 3600 2290 3800 2350
rect 3600 2210 3660 2290
rect 3740 2210 3800 2290
rect 3600 2150 3800 2210
rect 4000 2290 4200 2350
rect 4000 2210 4060 2290
rect 4140 2210 4200 2290
rect 4000 2150 4200 2210
rect 4400 2290 4600 2350
rect 4400 2210 4460 2290
rect 4540 2210 4600 2290
rect 4400 2150 4600 2210
rect 4800 2290 5000 2350
rect 4800 2210 4860 2290
rect 4940 2210 5000 2290
rect 4800 2150 5000 2210
rect 5200 2290 5400 2350
rect 5200 2210 5260 2290
rect 5340 2210 5400 2290
rect 5200 2150 5400 2210
rect 5600 2290 5800 2350
rect 5600 2210 5660 2290
rect 5740 2210 5800 2290
rect 5600 2150 5800 2210
rect 6000 2290 6200 2350
rect 6000 2210 6060 2290
rect 6140 2210 6200 2290
rect 6000 2150 6200 2210
rect 6400 2290 6600 2350
rect 6400 2210 6460 2290
rect 6540 2210 6600 2290
rect 6400 2150 6600 2210
rect 6800 2290 7000 2350
rect 6800 2210 6860 2290
rect 6940 2210 7000 2290
rect 6800 2150 7000 2210
rect 7200 2290 7400 2350
rect 7200 2210 7260 2290
rect 7340 2210 7400 2290
rect 7200 2150 7400 2210
rect 7600 2290 7800 2350
rect 7600 2210 7660 2290
rect 7740 2210 7800 2290
rect 7600 2150 7800 2210
rect 8000 2290 8200 2350
rect 8000 2210 8060 2290
rect 8140 2210 8200 2290
rect 8000 2150 8200 2210
rect 8400 2290 8600 2350
rect 8400 2210 8460 2290
rect 8540 2210 8600 2290
rect 8400 2150 8600 2210
rect 8800 2290 9000 2350
rect 8800 2210 8860 2290
rect 8940 2210 9000 2290
rect 8800 2150 9000 2210
rect 9200 2290 9400 2350
rect 9200 2210 9260 2290
rect 9340 2210 9400 2290
rect 9200 2150 9400 2210
rect 9600 2290 9800 2350
rect 9600 2210 9660 2290
rect 9740 2210 9800 2290
rect 9600 2150 9800 2210
rect 2200 2090 2400 2150
rect 2200 2010 2260 2090
rect 2340 2010 2400 2090
rect 2200 1950 2400 2010
rect 2600 2090 2800 2150
rect 2600 2010 2660 2090
rect 2740 2010 2800 2090
rect 2600 1950 2800 2010
rect 3000 2090 3200 2150
rect 3000 2010 3060 2090
rect 3140 2010 3200 2090
rect 3000 1950 3200 2010
rect 3400 2090 3600 2150
rect 3400 2010 3460 2090
rect 3540 2010 3600 2090
rect 3400 1950 3600 2010
rect 3800 2090 4000 2150
rect 3800 2010 3860 2090
rect 3940 2010 4000 2090
rect 3800 1950 4000 2010
rect 4200 2090 4400 2150
rect 4200 2010 4260 2090
rect 4340 2010 4400 2090
rect 4200 1950 4400 2010
rect 4600 2090 4800 2150
rect 4600 2010 4660 2090
rect 4740 2010 4800 2090
rect 4600 1950 4800 2010
rect 5000 2090 5200 2150
rect 5000 2010 5060 2090
rect 5140 2010 5200 2090
rect 5000 1950 5200 2010
rect 5400 2090 5600 2150
rect 5400 2010 5460 2090
rect 5540 2010 5600 2090
rect 5400 1950 5600 2010
rect 5800 2090 6000 2150
rect 5800 2010 5860 2090
rect 5940 2010 6000 2090
rect 5800 1950 6000 2010
rect 6200 2090 6400 2150
rect 6200 2010 6260 2090
rect 6340 2010 6400 2090
rect 6200 1950 6400 2010
rect 6600 2090 6800 2150
rect 6600 2010 6660 2090
rect 6740 2010 6800 2090
rect 6600 1950 6800 2010
rect 7000 2090 7200 2150
rect 7000 2010 7060 2090
rect 7140 2010 7200 2090
rect 7000 1950 7200 2010
rect 7400 2090 7600 2150
rect 7400 2010 7460 2090
rect 7540 2010 7600 2090
rect 7400 1950 7600 2010
rect 7800 2090 8000 2150
rect 7800 2010 7860 2090
rect 7940 2010 8000 2090
rect 7800 1950 8000 2010
rect 8200 2090 8400 2150
rect 8200 2010 8260 2090
rect 8340 2010 8400 2090
rect 8200 1950 8400 2010
rect 8600 2090 8800 2150
rect 8600 2010 8660 2090
rect 8740 2010 8800 2090
rect 8600 1950 8800 2010
rect 9000 2090 9200 2150
rect 9000 2010 9060 2090
rect 9140 2010 9200 2090
rect 9000 1950 9200 2010
rect 9400 2090 9600 2150
rect 9400 2010 9460 2090
rect 9540 2010 9600 2090
rect 9400 1950 9600 2010
rect 9800 2090 10000 2150
rect 9800 2010 9860 2090
rect 9940 2010 10000 2090
rect 9800 1950 10000 2010
rect 2400 1890 2600 1950
rect 2400 1810 2460 1890
rect 2540 1810 2600 1890
rect 2400 1750 2600 1810
rect 2800 1890 3000 1950
rect 2800 1810 2860 1890
rect 2940 1810 3000 1890
rect 2800 1750 3000 1810
rect 3200 1890 3400 1950
rect 3200 1810 3260 1890
rect 3340 1810 3400 1890
rect 3200 1750 3400 1810
rect 3600 1890 3800 1950
rect 3600 1810 3660 1890
rect 3740 1810 3800 1890
rect 3600 1750 3800 1810
rect 4000 1890 4200 1950
rect 4000 1810 4060 1890
rect 4140 1810 4200 1890
rect 4000 1750 4200 1810
rect 4400 1890 4600 1950
rect 4400 1810 4460 1890
rect 4540 1810 4600 1890
rect 4400 1750 4600 1810
rect 4800 1890 5000 1950
rect 4800 1810 4860 1890
rect 4940 1810 5000 1890
rect 4800 1750 5000 1810
rect 5200 1890 5400 1950
rect 5200 1810 5260 1890
rect 5340 1810 5400 1890
rect 5200 1750 5400 1810
rect 5600 1890 5800 1950
rect 5600 1810 5660 1890
rect 5740 1810 5800 1890
rect 5600 1750 5800 1810
rect 6000 1890 6200 1950
rect 6000 1810 6060 1890
rect 6140 1810 6200 1890
rect 6000 1750 6200 1810
rect 6400 1890 6600 1950
rect 6400 1810 6460 1890
rect 6540 1810 6600 1890
rect 6400 1750 6600 1810
rect 6800 1890 7000 1950
rect 6800 1810 6860 1890
rect 6940 1810 7000 1890
rect 6800 1750 7000 1810
rect 7200 1890 7400 1950
rect 7200 1810 7260 1890
rect 7340 1810 7400 1890
rect 7200 1750 7400 1810
rect 7600 1890 7800 1950
rect 7600 1810 7660 1890
rect 7740 1810 7800 1890
rect 7600 1750 7800 1810
rect 8000 1890 8200 1950
rect 8000 1810 8060 1890
rect 8140 1810 8200 1890
rect 8000 1750 8200 1810
rect 8400 1890 8600 1950
rect 8400 1810 8460 1890
rect 8540 1810 8600 1890
rect 8400 1750 8600 1810
rect 8800 1890 9000 1950
rect 8800 1810 8860 1890
rect 8940 1810 9000 1890
rect 8800 1750 9000 1810
rect 9200 1890 9400 1950
rect 9200 1810 9260 1890
rect 9340 1810 9400 1890
rect 9200 1750 9400 1810
rect 9600 1890 9800 1950
rect 9600 1810 9660 1890
rect 9740 1810 9800 1890
rect 9600 1750 9800 1810
rect 2200 1690 2400 1750
rect 2200 1610 2260 1690
rect 2340 1610 2400 1690
rect 2200 1550 2400 1610
rect 2600 1690 2800 1750
rect 2600 1610 2660 1690
rect 2740 1610 2800 1690
rect 2600 1550 2800 1610
rect 3000 1690 3200 1750
rect 3000 1610 3060 1690
rect 3140 1610 3200 1690
rect 3000 1550 3200 1610
rect 3400 1690 3600 1750
rect 3400 1610 3460 1690
rect 3540 1610 3600 1690
rect 3400 1550 3600 1610
rect 3800 1690 4000 1750
rect 3800 1610 3860 1690
rect 3940 1610 4000 1690
rect 3800 1550 4000 1610
rect 4200 1690 4400 1750
rect 4200 1610 4260 1690
rect 4340 1610 4400 1690
rect 4200 1550 4400 1610
rect 4600 1690 4800 1750
rect 4600 1610 4660 1690
rect 4740 1610 4800 1690
rect 4600 1550 4800 1610
rect 5000 1690 5200 1750
rect 5000 1610 5060 1690
rect 5140 1610 5200 1690
rect 5000 1550 5200 1610
rect 5400 1690 5600 1750
rect 5400 1610 5460 1690
rect 5540 1610 5600 1690
rect 5400 1550 5600 1610
rect 5800 1690 6000 1750
rect 5800 1610 5860 1690
rect 5940 1610 6000 1690
rect 5800 1550 6000 1610
rect 6200 1690 6400 1750
rect 6200 1610 6260 1690
rect 6340 1610 6400 1690
rect 6200 1550 6400 1610
rect 6600 1690 6800 1750
rect 6600 1610 6660 1690
rect 6740 1610 6800 1690
rect 6600 1550 6800 1610
rect 7000 1690 7200 1750
rect 7000 1610 7060 1690
rect 7140 1610 7200 1690
rect 7000 1550 7200 1610
rect 7400 1690 7600 1750
rect 7400 1610 7460 1690
rect 7540 1610 7600 1690
rect 7400 1550 7600 1610
rect 7800 1690 8000 1750
rect 7800 1610 7860 1690
rect 7940 1610 8000 1690
rect 7800 1550 8000 1610
rect 8200 1690 8400 1750
rect 8200 1610 8260 1690
rect 8340 1610 8400 1690
rect 8200 1550 8400 1610
rect 8600 1690 8800 1750
rect 8600 1610 8660 1690
rect 8740 1610 8800 1690
rect 8600 1550 8800 1610
rect 9000 1690 9200 1750
rect 9000 1610 9060 1690
rect 9140 1610 9200 1690
rect 9000 1550 9200 1610
rect 9400 1690 9600 1750
rect 9400 1610 9460 1690
rect 9540 1610 9600 1690
rect 9400 1550 9600 1610
rect 9800 1690 10000 1750
rect 9800 1610 9860 1690
rect 9940 1610 10000 1690
rect 9800 1550 10000 1610
rect 2400 1490 2600 1550
rect 2400 1410 2460 1490
rect 2540 1410 2600 1490
rect 2400 1350 2600 1410
rect 2800 1490 3000 1550
rect 2800 1410 2860 1490
rect 2940 1410 3000 1490
rect 2800 1350 3000 1410
rect 3200 1490 3400 1550
rect 3200 1410 3260 1490
rect 3340 1410 3400 1490
rect 3200 1350 3400 1410
rect 3600 1490 3800 1550
rect 3600 1410 3660 1490
rect 3740 1410 3800 1490
rect 3600 1350 3800 1410
rect 4000 1490 4200 1550
rect 4000 1410 4060 1490
rect 4140 1410 4200 1490
rect 4000 1350 4200 1410
rect 4400 1490 4600 1550
rect 4400 1410 4460 1490
rect 4540 1410 4600 1490
rect 4400 1350 4600 1410
rect 4800 1490 5000 1550
rect 4800 1410 4860 1490
rect 4940 1410 5000 1490
rect 4800 1350 5000 1410
rect 5200 1490 5400 1550
rect 5200 1410 5260 1490
rect 5340 1410 5400 1490
rect 5200 1350 5400 1410
rect 5600 1490 5800 1550
rect 5600 1410 5660 1490
rect 5740 1410 5800 1490
rect 5600 1350 5800 1410
rect 6000 1490 6200 1550
rect 6000 1410 6060 1490
rect 6140 1410 6200 1490
rect 6000 1350 6200 1410
rect 6400 1490 6600 1550
rect 6400 1410 6460 1490
rect 6540 1410 6600 1490
rect 6400 1350 6600 1410
rect 6800 1490 7000 1550
rect 6800 1410 6860 1490
rect 6940 1410 7000 1490
rect 6800 1350 7000 1410
rect 7200 1490 7400 1550
rect 7200 1410 7260 1490
rect 7340 1410 7400 1490
rect 7200 1350 7400 1410
rect 7600 1490 7800 1550
rect 7600 1410 7660 1490
rect 7740 1410 7800 1490
rect 7600 1350 7800 1410
rect 8000 1490 8200 1550
rect 8000 1410 8060 1490
rect 8140 1410 8200 1490
rect 8000 1350 8200 1410
rect 8400 1490 8600 1550
rect 8400 1410 8460 1490
rect 8540 1410 8600 1490
rect 8400 1350 8600 1410
rect 8800 1490 9000 1550
rect 8800 1410 8860 1490
rect 8940 1410 9000 1490
rect 8800 1350 9000 1410
rect 9200 1490 9400 1550
rect 9200 1410 9260 1490
rect 9340 1410 9400 1490
rect 9200 1350 9400 1410
rect 9600 1490 9800 1550
rect 9600 1410 9660 1490
rect 9740 1410 9800 1490
rect 9600 1350 9800 1410
rect 2200 1290 2400 1350
rect 2200 1210 2260 1290
rect 2340 1210 2400 1290
rect 2200 1150 2400 1210
rect 2600 1290 2800 1350
rect 2600 1210 2660 1290
rect 2740 1210 2800 1290
rect 2600 1150 2800 1210
rect 3000 1290 3200 1350
rect 3000 1210 3060 1290
rect 3140 1210 3200 1290
rect 3000 1150 3200 1210
rect 3400 1290 3600 1350
rect 3400 1210 3460 1290
rect 3540 1210 3600 1290
rect 3400 1150 3600 1210
rect 3800 1290 4000 1350
rect 3800 1210 3860 1290
rect 3940 1210 4000 1290
rect 3800 1150 4000 1210
rect 4200 1290 4400 1350
rect 4200 1210 4260 1290
rect 4340 1210 4400 1290
rect 4200 1150 4400 1210
rect 4600 1290 4800 1350
rect 4600 1210 4660 1290
rect 4740 1210 4800 1290
rect 4600 1150 4800 1210
rect 5000 1290 5200 1350
rect 5000 1210 5060 1290
rect 5140 1210 5200 1290
rect 5000 1150 5200 1210
rect 5400 1290 5600 1350
rect 5400 1210 5460 1290
rect 5540 1210 5600 1290
rect 5400 1150 5600 1210
rect 5800 1290 6000 1350
rect 5800 1210 5860 1290
rect 5940 1210 6000 1290
rect 5800 1150 6000 1210
rect 6200 1290 6400 1350
rect 6200 1210 6260 1290
rect 6340 1210 6400 1290
rect 6200 1150 6400 1210
rect 6600 1290 6800 1350
rect 6600 1210 6660 1290
rect 6740 1210 6800 1290
rect 6600 1150 6800 1210
rect 7000 1290 7200 1350
rect 7000 1210 7060 1290
rect 7140 1210 7200 1290
rect 7000 1150 7200 1210
rect 7400 1290 7600 1350
rect 7400 1210 7460 1290
rect 7540 1210 7600 1290
rect 7400 1150 7600 1210
rect 7800 1290 8000 1350
rect 7800 1210 7860 1290
rect 7940 1210 8000 1290
rect 7800 1150 8000 1210
rect 8200 1290 8400 1350
rect 8200 1210 8260 1290
rect 8340 1210 8400 1290
rect 8200 1150 8400 1210
rect 8600 1290 8800 1350
rect 8600 1210 8660 1290
rect 8740 1210 8800 1290
rect 8600 1150 8800 1210
rect 9000 1290 9200 1350
rect 9000 1210 9060 1290
rect 9140 1210 9200 1290
rect 9000 1150 9200 1210
rect 9400 1290 9600 1350
rect 9400 1210 9460 1290
rect 9540 1210 9600 1290
rect 9400 1150 9600 1210
rect 9800 1290 10000 1350
rect 9800 1210 9860 1290
rect 9940 1210 10000 1290
rect 9800 1150 10000 1210
rect 2400 1090 2600 1150
rect 2400 1010 2460 1090
rect 2540 1010 2600 1090
rect 2400 950 2600 1010
rect 2800 1090 3000 1150
rect 2800 1010 2860 1090
rect 2940 1010 3000 1090
rect 2800 950 3000 1010
rect 3200 1090 3400 1150
rect 3200 1010 3260 1090
rect 3340 1010 3400 1090
rect 3200 950 3400 1010
rect 3600 1090 3800 1150
rect 3600 1010 3660 1090
rect 3740 1010 3800 1090
rect 3600 950 3800 1010
rect 4000 1090 4200 1150
rect 4000 1010 4060 1090
rect 4140 1010 4200 1090
rect 4000 950 4200 1010
rect 4400 1090 4600 1150
rect 4400 1010 4460 1090
rect 4540 1010 4600 1090
rect 4400 950 4600 1010
rect 4800 1090 5000 1150
rect 4800 1010 4860 1090
rect 4940 1010 5000 1090
rect 4800 950 5000 1010
rect 5200 1090 5400 1150
rect 5200 1010 5260 1090
rect 5340 1010 5400 1090
rect 5200 950 5400 1010
rect 5600 1090 5800 1150
rect 5600 1010 5660 1090
rect 5740 1010 5800 1090
rect 5600 950 5800 1010
rect 6000 1090 6200 1150
rect 6000 1010 6060 1090
rect 6140 1010 6200 1090
rect 6000 950 6200 1010
rect 6400 1090 6600 1150
rect 6400 1010 6460 1090
rect 6540 1010 6600 1090
rect 6400 950 6600 1010
rect 6800 1090 7000 1150
rect 6800 1010 6860 1090
rect 6940 1010 7000 1090
rect 6800 950 7000 1010
rect 7200 1090 7400 1150
rect 7200 1010 7260 1090
rect 7340 1010 7400 1090
rect 7200 950 7400 1010
rect 7600 1090 7800 1150
rect 7600 1010 7660 1090
rect 7740 1010 7800 1090
rect 7600 950 7800 1010
rect 8000 1090 8200 1150
rect 8000 1010 8060 1090
rect 8140 1010 8200 1090
rect 8000 950 8200 1010
rect 8400 1090 8600 1150
rect 8400 1010 8460 1090
rect 8540 1010 8600 1090
rect 8400 950 8600 1010
rect 8800 1090 9000 1150
rect 8800 1010 8860 1090
rect 8940 1010 9000 1090
rect 8800 950 9000 1010
rect 9200 1090 9400 1150
rect 9200 1010 9260 1090
rect 9340 1010 9400 1090
rect 9200 950 9400 1010
rect 9600 1090 9800 1150
rect 9600 1010 9660 1090
rect 9740 1010 9800 1090
rect 9600 950 9800 1010
rect 2200 890 2400 950
rect 2200 810 2260 890
rect 2340 810 2400 890
rect 2200 750 2400 810
rect 2600 890 2800 950
rect 2600 810 2660 890
rect 2740 810 2800 890
rect 2600 750 2800 810
rect 3000 890 3200 950
rect 3000 810 3060 890
rect 3140 810 3200 890
rect 3000 750 3200 810
rect 3400 890 3600 950
rect 3400 810 3460 890
rect 3540 810 3600 890
rect 3400 750 3600 810
rect 3800 890 4000 950
rect 3800 810 3860 890
rect 3940 810 4000 890
rect 3800 750 4000 810
rect 4200 890 4400 950
rect 4200 810 4260 890
rect 4340 810 4400 890
rect 4200 750 4400 810
rect 4600 890 4800 950
rect 4600 810 4660 890
rect 4740 810 4800 890
rect 4600 750 4800 810
rect 5000 890 5200 950
rect 5000 810 5060 890
rect 5140 810 5200 890
rect 5000 750 5200 810
rect 5400 890 5600 950
rect 5400 810 5460 890
rect 5540 810 5600 890
rect 5400 750 5600 810
rect 5800 890 6000 950
rect 5800 810 5860 890
rect 5940 810 6000 890
rect 5800 750 6000 810
rect 6200 890 6400 950
rect 6200 810 6260 890
rect 6340 810 6400 890
rect 6200 750 6400 810
rect 6600 890 6800 950
rect 6600 810 6660 890
rect 6740 810 6800 890
rect 6600 750 6800 810
rect 7000 890 7200 950
rect 7000 810 7060 890
rect 7140 810 7200 890
rect 7000 750 7200 810
rect 7400 890 7600 950
rect 7400 810 7460 890
rect 7540 810 7600 890
rect 7400 750 7600 810
rect 7800 890 8000 950
rect 7800 810 7860 890
rect 7940 810 8000 890
rect 7800 750 8000 810
rect 8200 890 8400 950
rect 8200 810 8260 890
rect 8340 810 8400 890
rect 8200 750 8400 810
rect 8600 890 8800 950
rect 8600 810 8660 890
rect 8740 810 8800 890
rect 8600 750 8800 810
rect 9000 890 9200 950
rect 9000 810 9060 890
rect 9140 810 9200 890
rect 9000 750 9200 810
rect 9400 890 9600 950
rect 9400 810 9460 890
rect 9540 810 9600 890
rect 9400 750 9600 810
rect 9800 890 10000 950
rect 9800 810 9860 890
rect 9940 810 10000 890
rect 9800 750 10000 810
rect 2400 690 2600 750
rect 2400 610 2460 690
rect 2540 610 2600 690
rect 2400 550 2600 610
rect 2800 690 3000 750
rect 2800 610 2860 690
rect 2940 610 3000 690
rect 2800 550 3000 610
rect 3200 690 3400 750
rect 3200 610 3260 690
rect 3340 610 3400 690
rect 3200 550 3400 610
rect 3600 690 3800 750
rect 3600 610 3660 690
rect 3740 610 3800 690
rect 3600 550 3800 610
rect 4000 690 4200 750
rect 4000 610 4060 690
rect 4140 610 4200 690
rect 4000 550 4200 610
rect 4400 690 4600 750
rect 4400 610 4460 690
rect 4540 610 4600 690
rect 4400 550 4600 610
rect 4800 690 5000 750
rect 4800 610 4860 690
rect 4940 610 5000 690
rect 4800 550 5000 610
rect 5200 690 5400 750
rect 5200 610 5260 690
rect 5340 610 5400 690
rect 5200 550 5400 610
rect 5600 690 5800 750
rect 5600 610 5660 690
rect 5740 610 5800 690
rect 5600 550 5800 610
rect 6000 690 6200 750
rect 6000 610 6060 690
rect 6140 610 6200 690
rect 6000 550 6200 610
rect 6400 690 6600 750
rect 6400 610 6460 690
rect 6540 610 6600 690
rect 6400 550 6600 610
rect 6800 690 7000 750
rect 6800 610 6860 690
rect 6940 610 7000 690
rect 6800 550 7000 610
rect 7200 690 7400 750
rect 7200 610 7260 690
rect 7340 610 7400 690
rect 7200 550 7400 610
rect 7600 690 7800 750
rect 7600 610 7660 690
rect 7740 610 7800 690
rect 7600 550 7800 610
rect 8000 690 8200 750
rect 8000 610 8060 690
rect 8140 610 8200 690
rect 8000 550 8200 610
rect 8400 690 8600 750
rect 8400 610 8460 690
rect 8540 610 8600 690
rect 8400 550 8600 610
rect 8800 690 9000 750
rect 8800 610 8860 690
rect 8940 610 9000 690
rect 8800 550 9000 610
rect 9200 690 9400 750
rect 9200 610 9260 690
rect 9340 610 9400 690
rect 9200 550 9400 610
rect 9600 690 9800 750
rect 9600 610 9660 690
rect 9740 610 9800 690
rect 9600 550 9800 610
rect 2200 490 2400 550
rect 2200 410 2260 490
rect 2340 410 2400 490
rect 2200 350 2400 410
rect 2600 490 2800 550
rect 2600 410 2660 490
rect 2740 410 2800 490
rect 2600 350 2800 410
rect 3000 490 3200 550
rect 3000 410 3060 490
rect 3140 410 3200 490
rect 3000 350 3200 410
rect 3400 490 3600 550
rect 3400 410 3460 490
rect 3540 410 3600 490
rect 3400 350 3600 410
rect 3800 490 4000 550
rect 3800 410 3860 490
rect 3940 410 4000 490
rect 3800 350 4000 410
rect 4200 490 4400 550
rect 4200 410 4260 490
rect 4340 410 4400 490
rect 4200 350 4400 410
rect 4600 490 4800 550
rect 4600 410 4660 490
rect 4740 410 4800 490
rect 4600 350 4800 410
rect 5000 490 5200 550
rect 5000 410 5060 490
rect 5140 410 5200 490
rect 5000 350 5200 410
rect 5400 490 5600 550
rect 5400 410 5460 490
rect 5540 410 5600 490
rect 5400 350 5600 410
rect 5800 490 6000 550
rect 5800 410 5860 490
rect 5940 410 6000 490
rect 5800 350 6000 410
rect 6200 490 6400 550
rect 6200 410 6260 490
rect 6340 410 6400 490
rect 6200 350 6400 410
rect 6600 490 6800 550
rect 6600 410 6660 490
rect 6740 410 6800 490
rect 6600 350 6800 410
rect 7000 490 7200 550
rect 7000 410 7060 490
rect 7140 410 7200 490
rect 7000 350 7200 410
rect 7400 490 7600 550
rect 7400 410 7460 490
rect 7540 410 7600 490
rect 7400 350 7600 410
rect 7800 490 8000 550
rect 7800 410 7860 490
rect 7940 410 8000 490
rect 7800 350 8000 410
rect 8200 490 8400 550
rect 8200 410 8260 490
rect 8340 410 8400 490
rect 8200 350 8400 410
rect 8600 490 8800 550
rect 8600 410 8660 490
rect 8740 410 8800 490
rect 8600 350 8800 410
rect 9000 490 9200 550
rect 9000 410 9060 490
rect 9140 410 9200 490
rect 9000 350 9200 410
rect 9400 490 9600 550
rect 9400 410 9460 490
rect 9540 410 9600 490
rect 9400 350 9600 410
rect 9800 490 10000 550
rect 9800 410 9860 490
rect 9940 410 10000 490
rect 9800 350 10000 410
rect 10100 250 10350 8250
rect 1850 0 10350 250
<< gv1 >>
rect 160 33730 240 33810
rect 11960 33730 12040 33810
rect 9140 33600 9220 33680
rect 9440 33600 9520 33680
rect 10020 33600 10100 33680
rect 10610 33600 10690 33680
rect 11200 33600 11280 33680
rect 11500 33600 11580 33680
rect 160 33450 240 33530
rect 11960 33450 12040 33530
rect 9140 33320 9220 33400
rect 9440 33320 9520 33400
rect 10020 33320 10100 33400
rect 10610 33320 10690 33400
rect 11200 33320 11280 33400
rect 11500 33320 11580 33400
rect 160 33170 240 33250
rect 11960 33170 12040 33250
rect 160 32890 240 32970
rect 9000 32870 9080 32950
rect 9160 32870 9240 32950
rect 10360 32870 10440 32950
rect 10540 32870 10620 32950
rect 10960 32870 11040 32950
rect 11140 32870 11220 32950
rect 11960 32890 12040 32970
rect 160 32610 240 32690
rect 11960 32610 12040 32690
rect 8860 31510 8940 31590
rect 9140 31510 9220 31590
rect 10020 31510 10100 31590
rect 10320 31510 10400 31590
rect 10620 31510 10700 31590
rect 10920 31510 11000 31590
rect 11230 31510 11310 31590
rect 160 31430 240 31510
rect 11960 31430 12040 31510
rect 160 31150 240 31230
rect 6596 31088 6676 31168
rect 6756 31088 6836 31168
rect 8201 31088 8281 31168
rect 8471 31088 8551 31168
rect 11960 31150 12040 31230
rect 9140 31060 9220 31140
rect 9440 31060 9520 31140
rect 10020 31060 10100 31140
rect 10620 31060 10700 31140
rect 11220 31060 11300 31140
rect 11520 31060 11600 31140
rect 160 30870 240 30950
rect 6596 30928 6676 31008
rect 6756 30928 6836 31008
rect 8201 30928 8281 31008
rect 8471 30928 8551 31008
rect 11960 30870 12040 30950
rect 9140 30780 9220 30860
rect 9440 30780 9520 30860
rect 10020 30780 10100 30860
rect 10620 30780 10700 30860
rect 11220 30780 11300 30860
rect 11520 30780 11600 30860
rect 160 30590 240 30670
rect 11960 30590 12040 30670
rect 160 30310 240 30390
rect 11960 30310 12040 30390
rect 7885 29565 7965 29645
rect 8065 29565 8145 29645
rect 8245 29565 8325 29645
rect 8425 29565 8505 29645
rect 8605 29565 8685 29645
rect 7885 29385 7965 29465
rect 8065 29385 8145 29465
rect 8245 29385 8325 29465
rect 8425 29385 8505 29465
rect 8605 29385 8685 29465
rect 7885 29205 7965 29285
rect 8065 29205 8145 29285
rect 8245 29205 8325 29285
rect 8425 29205 8505 29285
rect 8605 29205 8685 29285
rect 7885 29025 7965 29105
rect 8065 29025 8145 29105
rect 8245 29025 8325 29105
rect 8425 29025 8505 29105
rect 8605 29025 8685 29105
rect 7885 28845 7965 28925
rect 8065 28845 8145 28925
rect 8245 28845 8325 28925
rect 8425 28845 8505 28925
rect 8605 28845 8685 28925
rect 160 28090 240 28170
rect 11660 28090 11740 28170
rect 11960 28090 12040 28170
rect 160 27910 240 27990
rect 11660 27910 11740 27990
rect 11960 27910 12040 27990
rect 160 27730 240 27810
rect 11660 27730 11740 27810
rect 11960 27730 12040 27810
rect 160 27550 240 27630
rect 11660 27550 11740 27630
rect 11960 27550 12040 27630
rect 160 27370 240 27450
rect 11660 27370 11740 27450
rect 11960 27370 12040 27450
rect 160 27190 240 27270
rect 870 27190 950 27270
rect 1170 27190 1250 27270
rect 1490 27190 1570 27270
rect 1810 27190 1890 27270
rect 2130 27190 2210 27270
rect 2430 27190 2510 27270
rect 2750 27190 2830 27270
rect 3070 27190 3150 27270
rect 3390 27190 3470 27270
rect 3690 27190 3770 27270
rect 4010 27190 4090 27270
rect 4330 27190 4410 27270
rect 4650 27190 4730 27270
rect 4950 27190 5030 27270
rect 5270 27190 5350 27270
rect 5590 27190 5670 27270
rect 5910 27190 5990 27270
rect 6210 27190 6290 27270
rect 6530 27190 6610 27270
rect 6850 27190 6930 27270
rect 7170 27190 7250 27270
rect 7470 27190 7550 27270
rect 7790 27190 7870 27270
rect 8110 27190 8190 27270
rect 8430 27190 8510 27270
rect 8730 27190 8810 27270
rect 9050 27190 9130 27270
rect 9370 27190 9450 27270
rect 9690 27190 9770 27270
rect 9990 27190 10070 27270
rect 10310 27190 10390 27270
rect 10630 27190 10710 27270
rect 10950 27190 11030 27270
rect 11250 27190 11330 27270
rect 11660 27190 11740 27270
rect 11960 27190 12040 27270
rect 160 27010 240 27090
rect 870 27010 950 27090
rect 1170 27010 1250 27090
rect 1490 27010 1570 27090
rect 1810 27010 1890 27090
rect 2130 27010 2210 27090
rect 2430 27010 2510 27090
rect 2750 27010 2830 27090
rect 3070 27010 3150 27090
rect 3390 27010 3470 27090
rect 3690 27010 3770 27090
rect 4010 27010 4090 27090
rect 4330 27010 4410 27090
rect 4650 27010 4730 27090
rect 4950 27010 5030 27090
rect 5270 27010 5350 27090
rect 5590 27010 5670 27090
rect 5910 27010 5990 27090
rect 6210 27010 6290 27090
rect 6530 27010 6610 27090
rect 6850 27010 6930 27090
rect 7170 27010 7250 27090
rect 7470 27010 7550 27090
rect 7790 27010 7870 27090
rect 8110 27010 8190 27090
rect 8430 27010 8510 27090
rect 8730 27010 8810 27090
rect 9050 27010 9130 27090
rect 9370 27010 9450 27090
rect 9690 27010 9770 27090
rect 9990 27010 10070 27090
rect 10310 27010 10390 27090
rect 10630 27010 10710 27090
rect 10950 27010 11030 27090
rect 11250 27010 11330 27090
rect 11660 27010 11740 27090
rect 11960 27010 12040 27090
rect 160 26830 240 26910
rect 870 26830 950 26910
rect 1170 26830 1250 26910
rect 1490 26830 1570 26910
rect 1810 26830 1890 26910
rect 2130 26830 2210 26910
rect 2430 26830 2510 26910
rect 2750 26830 2830 26910
rect 3070 26830 3150 26910
rect 3390 26830 3470 26910
rect 3690 26830 3770 26910
rect 4010 26830 4090 26910
rect 4330 26830 4410 26910
rect 4650 26830 4730 26910
rect 4950 26830 5030 26910
rect 5270 26830 5350 26910
rect 5590 26830 5670 26910
rect 5910 26830 5990 26910
rect 6210 26830 6290 26910
rect 6530 26830 6610 26910
rect 6850 26830 6930 26910
rect 7170 26830 7250 26910
rect 7470 26830 7550 26910
rect 7790 26830 7870 26910
rect 8110 26830 8190 26910
rect 8430 26830 8510 26910
rect 8730 26830 8810 26910
rect 9050 26830 9130 26910
rect 9370 26830 9450 26910
rect 9690 26830 9770 26910
rect 9990 26830 10070 26910
rect 10310 26830 10390 26910
rect 10630 26830 10710 26910
rect 10950 26830 11030 26910
rect 11250 26830 11330 26910
rect 11660 26830 11740 26910
rect 11960 26830 12040 26910
rect 160 26650 240 26730
rect 870 26650 950 26730
rect 1170 26650 1250 26730
rect 1490 26650 1570 26730
rect 1810 26650 1890 26730
rect 2130 26650 2210 26730
rect 2430 26650 2510 26730
rect 2750 26650 2830 26730
rect 3070 26650 3150 26730
rect 3390 26650 3470 26730
rect 3690 26650 3770 26730
rect 4010 26650 4090 26730
rect 4330 26650 4410 26730
rect 4650 26650 4730 26730
rect 4950 26650 5030 26730
rect 5270 26650 5350 26730
rect 5590 26650 5670 26730
rect 5910 26650 5990 26730
rect 6210 26650 6290 26730
rect 6530 26650 6610 26730
rect 6850 26650 6930 26730
rect 7170 26650 7250 26730
rect 7470 26650 7550 26730
rect 7790 26650 7870 26730
rect 8110 26650 8190 26730
rect 8430 26650 8510 26730
rect 8730 26650 8810 26730
rect 9050 26650 9130 26730
rect 9370 26650 9450 26730
rect 9690 26650 9770 26730
rect 9990 26650 10070 26730
rect 10310 26650 10390 26730
rect 10630 26650 10710 26730
rect 10950 26650 11030 26730
rect 11250 26650 11330 26730
rect 11660 26650 11740 26730
rect 11960 26650 12040 26730
rect 160 26470 240 26550
rect 870 26470 950 26550
rect 1170 26470 1250 26550
rect 1490 26470 1570 26550
rect 1810 26470 1890 26550
rect 2130 26470 2210 26550
rect 2430 26470 2510 26550
rect 2750 26470 2830 26550
rect 3070 26470 3150 26550
rect 3390 26470 3470 26550
rect 3690 26470 3770 26550
rect 4010 26470 4090 26550
rect 4330 26470 4410 26550
rect 4650 26470 4730 26550
rect 4950 26470 5030 26550
rect 5270 26470 5350 26550
rect 5590 26470 5670 26550
rect 5910 26470 5990 26550
rect 6210 26470 6290 26550
rect 6530 26470 6610 26550
rect 6850 26470 6930 26550
rect 7170 26470 7250 26550
rect 7470 26470 7550 26550
rect 7790 26470 7870 26550
rect 8110 26470 8190 26550
rect 8430 26470 8510 26550
rect 8730 26470 8810 26550
rect 9050 26470 9130 26550
rect 9370 26470 9450 26550
rect 9690 26470 9770 26550
rect 9990 26470 10070 26550
rect 10310 26470 10390 26550
rect 10630 26470 10710 26550
rect 10950 26470 11030 26550
rect 11250 26470 11330 26550
rect 11660 26470 11740 26550
rect 11960 26470 12040 26550
rect 160 26290 240 26370
rect 870 26290 950 26370
rect 1170 26290 1250 26370
rect 1490 26290 1570 26370
rect 1810 26290 1890 26370
rect 2130 26290 2210 26370
rect 2430 26290 2510 26370
rect 2750 26290 2830 26370
rect 3070 26290 3150 26370
rect 3390 26290 3470 26370
rect 3690 26290 3770 26370
rect 4010 26290 4090 26370
rect 4330 26290 4410 26370
rect 4650 26290 4730 26370
rect 4950 26290 5030 26370
rect 5270 26290 5350 26370
rect 5590 26290 5670 26370
rect 5910 26290 5990 26370
rect 6210 26290 6290 26370
rect 6530 26290 6610 26370
rect 6850 26290 6930 26370
rect 7170 26290 7250 26370
rect 7470 26290 7550 26370
rect 7790 26290 7870 26370
rect 8110 26290 8190 26370
rect 8430 26290 8510 26370
rect 8730 26290 8810 26370
rect 9050 26290 9130 26370
rect 9370 26290 9450 26370
rect 9690 26290 9770 26370
rect 9990 26290 10070 26370
rect 10310 26290 10390 26370
rect 10630 26290 10710 26370
rect 10950 26290 11030 26370
rect 11250 26290 11330 26370
rect 11660 26290 11740 26370
rect 11960 26290 12040 26370
rect 160 26110 240 26190
rect 870 26110 950 26190
rect 1170 26110 1250 26190
rect 1490 26110 1570 26190
rect 1810 26110 1890 26190
rect 2130 26110 2210 26190
rect 2430 26110 2510 26190
rect 2750 26110 2830 26190
rect 3070 26110 3150 26190
rect 3390 26110 3470 26190
rect 3690 26110 3770 26190
rect 4010 26110 4090 26190
rect 4330 26110 4410 26190
rect 4650 26110 4730 26190
rect 4950 26110 5030 26190
rect 5270 26110 5350 26190
rect 5590 26110 5670 26190
rect 5910 26110 5990 26190
rect 6210 26110 6290 26190
rect 6530 26110 6610 26190
rect 6850 26110 6930 26190
rect 7170 26110 7250 26190
rect 7470 26110 7550 26190
rect 7790 26110 7870 26190
rect 8110 26110 8190 26190
rect 8430 26110 8510 26190
rect 8730 26110 8810 26190
rect 9050 26110 9130 26190
rect 9370 26110 9450 26190
rect 9690 26110 9770 26190
rect 9990 26110 10070 26190
rect 10310 26110 10390 26190
rect 10630 26110 10710 26190
rect 10950 26110 11030 26190
rect 11250 26110 11330 26190
rect 11660 26110 11740 26190
rect 11960 26110 12040 26190
rect 160 25930 240 26010
rect 870 25930 950 26010
rect 1170 25930 1250 26010
rect 1490 25930 1570 26010
rect 1810 25930 1890 26010
rect 2130 25930 2210 26010
rect 2430 25930 2510 26010
rect 2750 25930 2830 26010
rect 3070 25930 3150 26010
rect 3390 25930 3470 26010
rect 3690 25930 3770 26010
rect 4010 25930 4090 26010
rect 4330 25930 4410 26010
rect 4650 25930 4730 26010
rect 4950 25930 5030 26010
rect 5270 25930 5350 26010
rect 5590 25930 5670 26010
rect 5910 25930 5990 26010
rect 6210 25930 6290 26010
rect 6530 25930 6610 26010
rect 6850 25930 6930 26010
rect 7170 25930 7250 26010
rect 7470 25930 7550 26010
rect 7790 25930 7870 26010
rect 8110 25930 8190 26010
rect 8430 25930 8510 26010
rect 8730 25930 8810 26010
rect 9050 25930 9130 26010
rect 9370 25930 9450 26010
rect 9690 25930 9770 26010
rect 9990 25930 10070 26010
rect 10310 25930 10390 26010
rect 10630 25930 10710 26010
rect 10950 25930 11030 26010
rect 11250 25930 11330 26010
rect 11660 25930 11740 26010
rect 11960 25930 12040 26010
rect 160 25750 240 25830
rect 870 25750 950 25830
rect 1170 25750 1250 25830
rect 1490 25750 1570 25830
rect 1810 25750 1890 25830
rect 2130 25750 2210 25830
rect 2430 25750 2510 25830
rect 2750 25750 2830 25830
rect 3070 25750 3150 25830
rect 3390 25750 3470 25830
rect 3690 25750 3770 25830
rect 4010 25750 4090 25830
rect 4330 25750 4410 25830
rect 4650 25750 4730 25830
rect 4950 25750 5030 25830
rect 5270 25750 5350 25830
rect 5590 25750 5670 25830
rect 5910 25750 5990 25830
rect 6210 25750 6290 25830
rect 6530 25750 6610 25830
rect 6850 25750 6930 25830
rect 7170 25750 7250 25830
rect 7470 25750 7550 25830
rect 7790 25750 7870 25830
rect 8110 25750 8190 25830
rect 8430 25750 8510 25830
rect 8730 25750 8810 25830
rect 9050 25750 9130 25830
rect 9370 25750 9450 25830
rect 9690 25750 9770 25830
rect 9990 25750 10070 25830
rect 10310 25750 10390 25830
rect 10630 25750 10710 25830
rect 10950 25750 11030 25830
rect 11250 25750 11330 25830
rect 11660 25750 11740 25830
rect 11960 25750 12040 25830
rect 160 25570 240 25650
rect 870 25570 950 25650
rect 1170 25570 1250 25650
rect 1490 25570 1570 25650
rect 1810 25570 1890 25650
rect 2130 25570 2210 25650
rect 2430 25570 2510 25650
rect 2750 25570 2830 25650
rect 3070 25570 3150 25650
rect 3390 25570 3470 25650
rect 3690 25570 3770 25650
rect 4010 25570 4090 25650
rect 4330 25570 4410 25650
rect 4650 25570 4730 25650
rect 4950 25570 5030 25650
rect 5270 25570 5350 25650
rect 5590 25570 5670 25650
rect 5910 25570 5990 25650
rect 6210 25570 6290 25650
rect 6530 25570 6610 25650
rect 6850 25570 6930 25650
rect 7170 25570 7250 25650
rect 7470 25570 7550 25650
rect 7790 25570 7870 25650
rect 8110 25570 8190 25650
rect 8430 25570 8510 25650
rect 8730 25570 8810 25650
rect 9050 25570 9130 25650
rect 9370 25570 9450 25650
rect 9690 25570 9770 25650
rect 9990 25570 10070 25650
rect 10310 25570 10390 25650
rect 10630 25570 10710 25650
rect 10950 25570 11030 25650
rect 11250 25570 11330 25650
rect 11660 25570 11740 25650
rect 11960 25570 12040 25650
rect 160 25390 240 25470
rect 870 25390 950 25470
rect 1170 25390 1250 25470
rect 1490 25390 1570 25470
rect 1810 25390 1890 25470
rect 2130 25390 2210 25470
rect 2430 25390 2510 25470
rect 2750 25390 2830 25470
rect 3070 25390 3150 25470
rect 3390 25390 3470 25470
rect 3690 25390 3770 25470
rect 4010 25390 4090 25470
rect 4330 25390 4410 25470
rect 4650 25390 4730 25470
rect 4950 25390 5030 25470
rect 5270 25390 5350 25470
rect 5590 25390 5670 25470
rect 5910 25390 5990 25470
rect 6210 25390 6290 25470
rect 6530 25390 6610 25470
rect 6850 25390 6930 25470
rect 7170 25390 7250 25470
rect 7470 25390 7550 25470
rect 7790 25390 7870 25470
rect 8110 25390 8190 25470
rect 8430 25390 8510 25470
rect 8730 25390 8810 25470
rect 9050 25390 9130 25470
rect 9370 25390 9450 25470
rect 9690 25390 9770 25470
rect 9990 25390 10070 25470
rect 10310 25390 10390 25470
rect 10630 25390 10710 25470
rect 10950 25390 11030 25470
rect 11250 25390 11330 25470
rect 11660 25390 11740 25470
rect 11960 25390 12040 25470
rect 160 25210 240 25290
rect 870 25210 950 25290
rect 1170 25210 1250 25290
rect 1490 25210 1570 25290
rect 1810 25210 1890 25290
rect 2130 25210 2210 25290
rect 2430 25210 2510 25290
rect 2750 25210 2830 25290
rect 3070 25210 3150 25290
rect 3390 25210 3470 25290
rect 3690 25210 3770 25290
rect 4010 25210 4090 25290
rect 4330 25210 4410 25290
rect 4650 25210 4730 25290
rect 4950 25210 5030 25290
rect 5270 25210 5350 25290
rect 5590 25210 5670 25290
rect 5910 25210 5990 25290
rect 6210 25210 6290 25290
rect 6530 25210 6610 25290
rect 6850 25210 6930 25290
rect 7170 25210 7250 25290
rect 7470 25210 7550 25290
rect 7790 25210 7870 25290
rect 8110 25210 8190 25290
rect 8430 25210 8510 25290
rect 8730 25210 8810 25290
rect 9050 25210 9130 25290
rect 9370 25210 9450 25290
rect 9690 25210 9770 25290
rect 9990 25210 10070 25290
rect 10310 25210 10390 25290
rect 10630 25210 10710 25290
rect 10950 25210 11030 25290
rect 11250 25210 11330 25290
rect 11660 25210 11740 25290
rect 11960 25210 12040 25290
rect 160 25030 240 25110
rect 870 25030 950 25110
rect 1170 25030 1250 25110
rect 1490 25030 1570 25110
rect 1810 25030 1890 25110
rect 2130 25030 2210 25110
rect 2430 25030 2510 25110
rect 2750 25030 2830 25110
rect 3070 25030 3150 25110
rect 3390 25030 3470 25110
rect 3690 25030 3770 25110
rect 4010 25030 4090 25110
rect 4330 25030 4410 25110
rect 4650 25030 4730 25110
rect 4950 25030 5030 25110
rect 5270 25030 5350 25110
rect 5590 25030 5670 25110
rect 5910 25030 5990 25110
rect 6210 25030 6290 25110
rect 6530 25030 6610 25110
rect 6850 25030 6930 25110
rect 7170 25030 7250 25110
rect 7470 25030 7550 25110
rect 7790 25030 7870 25110
rect 8110 25030 8190 25110
rect 8430 25030 8510 25110
rect 8730 25030 8810 25110
rect 9050 25030 9130 25110
rect 9370 25030 9450 25110
rect 9690 25030 9770 25110
rect 9990 25030 10070 25110
rect 10310 25030 10390 25110
rect 10630 25030 10710 25110
rect 10950 25030 11030 25110
rect 11250 25030 11330 25110
rect 11660 25030 11740 25110
rect 11960 25030 12040 25110
rect 160 24850 240 24930
rect 870 24850 950 24930
rect 1170 24850 1250 24930
rect 1490 24850 1570 24930
rect 1810 24850 1890 24930
rect 2130 24850 2210 24930
rect 2430 24850 2510 24930
rect 2750 24850 2830 24930
rect 3070 24850 3150 24930
rect 3390 24850 3470 24930
rect 3690 24850 3770 24930
rect 4010 24850 4090 24930
rect 4330 24850 4410 24930
rect 4650 24850 4730 24930
rect 4950 24850 5030 24930
rect 5270 24850 5350 24930
rect 5590 24850 5670 24930
rect 5910 24850 5990 24930
rect 6210 24850 6290 24930
rect 6530 24850 6610 24930
rect 6850 24850 6930 24930
rect 7170 24850 7250 24930
rect 7470 24850 7550 24930
rect 7790 24850 7870 24930
rect 8110 24850 8190 24930
rect 8430 24850 8510 24930
rect 8730 24850 8810 24930
rect 9050 24850 9130 24930
rect 9370 24850 9450 24930
rect 9690 24850 9770 24930
rect 9990 24850 10070 24930
rect 10310 24850 10390 24930
rect 10630 24850 10710 24930
rect 10950 24850 11030 24930
rect 11250 24850 11330 24930
rect 11660 24850 11740 24930
rect 11960 24850 12040 24930
rect 160 24670 240 24750
rect 870 24670 950 24750
rect 1170 24670 1250 24750
rect 1490 24670 1570 24750
rect 1810 24670 1890 24750
rect 2130 24670 2210 24750
rect 2430 24670 2510 24750
rect 2750 24670 2830 24750
rect 3070 24670 3150 24750
rect 3390 24670 3470 24750
rect 3690 24670 3770 24750
rect 4010 24670 4090 24750
rect 4330 24670 4410 24750
rect 4650 24670 4730 24750
rect 4950 24670 5030 24750
rect 5270 24670 5350 24750
rect 5590 24670 5670 24750
rect 5910 24670 5990 24750
rect 6210 24670 6290 24750
rect 6530 24670 6610 24750
rect 6850 24670 6930 24750
rect 7170 24670 7250 24750
rect 7470 24670 7550 24750
rect 7790 24670 7870 24750
rect 8110 24670 8190 24750
rect 8430 24670 8510 24750
rect 8730 24670 8810 24750
rect 9050 24670 9130 24750
rect 9370 24670 9450 24750
rect 9690 24670 9770 24750
rect 9990 24670 10070 24750
rect 10310 24670 10390 24750
rect 10630 24670 10710 24750
rect 10950 24670 11030 24750
rect 11250 24670 11330 24750
rect 11660 24670 11740 24750
rect 11960 24670 12040 24750
rect 160 24490 240 24570
rect 870 24490 950 24570
rect 1170 24490 1250 24570
rect 1490 24490 1570 24570
rect 1810 24490 1890 24570
rect 2130 24490 2210 24570
rect 2430 24490 2510 24570
rect 2750 24490 2830 24570
rect 3070 24490 3150 24570
rect 3390 24490 3470 24570
rect 3690 24490 3770 24570
rect 4010 24490 4090 24570
rect 4330 24490 4410 24570
rect 4650 24490 4730 24570
rect 4950 24490 5030 24570
rect 5270 24490 5350 24570
rect 5590 24490 5670 24570
rect 5910 24490 5990 24570
rect 6210 24490 6290 24570
rect 6530 24490 6610 24570
rect 6850 24490 6930 24570
rect 7170 24490 7250 24570
rect 7470 24490 7550 24570
rect 7790 24490 7870 24570
rect 8110 24490 8190 24570
rect 8430 24490 8510 24570
rect 8730 24490 8810 24570
rect 9050 24490 9130 24570
rect 9370 24490 9450 24570
rect 9690 24490 9770 24570
rect 9990 24490 10070 24570
rect 10310 24490 10390 24570
rect 10630 24490 10710 24570
rect 10950 24490 11030 24570
rect 11250 24490 11330 24570
rect 11660 24490 11740 24570
rect 11960 24490 12040 24570
rect 160 24310 240 24390
rect 870 24310 950 24390
rect 1170 24310 1250 24390
rect 1490 24310 1570 24390
rect 1810 24310 1890 24390
rect 2130 24310 2210 24390
rect 2430 24310 2510 24390
rect 2750 24310 2830 24390
rect 3070 24310 3150 24390
rect 3390 24310 3470 24390
rect 3690 24310 3770 24390
rect 4010 24310 4090 24390
rect 4330 24310 4410 24390
rect 4650 24310 4730 24390
rect 4950 24310 5030 24390
rect 5270 24310 5350 24390
rect 5590 24310 5670 24390
rect 5910 24310 5990 24390
rect 6210 24310 6290 24390
rect 6530 24310 6610 24390
rect 6850 24310 6930 24390
rect 7170 24310 7250 24390
rect 7470 24310 7550 24390
rect 7790 24310 7870 24390
rect 8110 24310 8190 24390
rect 8430 24310 8510 24390
rect 8730 24310 8810 24390
rect 9050 24310 9130 24390
rect 9370 24310 9450 24390
rect 9690 24310 9770 24390
rect 9990 24310 10070 24390
rect 10310 24310 10390 24390
rect 10630 24310 10710 24390
rect 10950 24310 11030 24390
rect 11250 24310 11330 24390
rect 11660 24310 11740 24390
rect 11960 24310 12040 24390
rect 160 24130 240 24210
rect 870 24130 950 24210
rect 1170 24130 1250 24210
rect 1490 24130 1570 24210
rect 1810 24130 1890 24210
rect 2130 24130 2210 24210
rect 2430 24130 2510 24210
rect 2750 24130 2830 24210
rect 3070 24130 3150 24210
rect 3390 24130 3470 24210
rect 3690 24130 3770 24210
rect 4010 24130 4090 24210
rect 4330 24130 4410 24210
rect 4650 24130 4730 24210
rect 4950 24130 5030 24210
rect 5270 24130 5350 24210
rect 5590 24130 5670 24210
rect 5910 24130 5990 24210
rect 6210 24130 6290 24210
rect 6530 24130 6610 24210
rect 6850 24130 6930 24210
rect 7170 24130 7250 24210
rect 7470 24130 7550 24210
rect 7790 24130 7870 24210
rect 8110 24130 8190 24210
rect 8430 24130 8510 24210
rect 8730 24130 8810 24210
rect 9050 24130 9130 24210
rect 9370 24130 9450 24210
rect 9690 24130 9770 24210
rect 9990 24130 10070 24210
rect 10310 24130 10390 24210
rect 10630 24130 10710 24210
rect 10950 24130 11030 24210
rect 11250 24130 11330 24210
rect 11660 24130 11740 24210
rect 11960 24130 12040 24210
rect 160 23950 240 24030
rect 870 23950 950 24030
rect 1170 23950 1250 24030
rect 1490 23950 1570 24030
rect 1810 23950 1890 24030
rect 2130 23950 2210 24030
rect 2430 23950 2510 24030
rect 2750 23950 2830 24030
rect 3070 23950 3150 24030
rect 3390 23950 3470 24030
rect 3690 23950 3770 24030
rect 4010 23950 4090 24030
rect 4330 23950 4410 24030
rect 4650 23950 4730 24030
rect 4950 23950 5030 24030
rect 5270 23950 5350 24030
rect 5590 23950 5670 24030
rect 5910 23950 5990 24030
rect 6210 23950 6290 24030
rect 6530 23950 6610 24030
rect 6850 23950 6930 24030
rect 7170 23950 7250 24030
rect 7470 23950 7550 24030
rect 7790 23950 7870 24030
rect 8110 23950 8190 24030
rect 8430 23950 8510 24030
rect 8730 23950 8810 24030
rect 9050 23950 9130 24030
rect 9370 23950 9450 24030
rect 9690 23950 9770 24030
rect 9990 23950 10070 24030
rect 10310 23950 10390 24030
rect 10630 23950 10710 24030
rect 10950 23950 11030 24030
rect 11250 23950 11330 24030
rect 11660 23950 11740 24030
rect 11960 23950 12040 24030
rect 160 23770 240 23850
rect 870 23770 950 23850
rect 1170 23770 1250 23850
rect 1490 23770 1570 23850
rect 1810 23770 1890 23850
rect 2130 23770 2210 23850
rect 2430 23770 2510 23850
rect 2750 23770 2830 23850
rect 3070 23770 3150 23850
rect 3390 23770 3470 23850
rect 3690 23770 3770 23850
rect 4010 23770 4090 23850
rect 4330 23770 4410 23850
rect 4650 23770 4730 23850
rect 4950 23770 5030 23850
rect 5270 23770 5350 23850
rect 5590 23770 5670 23850
rect 5910 23770 5990 23850
rect 6210 23770 6290 23850
rect 6530 23770 6610 23850
rect 6850 23770 6930 23850
rect 7170 23770 7250 23850
rect 7470 23770 7550 23850
rect 7790 23770 7870 23850
rect 8110 23770 8190 23850
rect 8430 23770 8510 23850
rect 8730 23770 8810 23850
rect 9050 23770 9130 23850
rect 9370 23770 9450 23850
rect 9690 23770 9770 23850
rect 9990 23770 10070 23850
rect 10310 23770 10390 23850
rect 10630 23770 10710 23850
rect 10950 23770 11030 23850
rect 11250 23770 11330 23850
rect 11660 23770 11740 23850
rect 11960 23770 12040 23850
rect 160 23590 240 23670
rect 870 23590 950 23670
rect 1170 23590 1250 23670
rect 1490 23590 1570 23670
rect 1810 23590 1890 23670
rect 2130 23590 2210 23670
rect 2430 23590 2510 23670
rect 2750 23590 2830 23670
rect 3070 23590 3150 23670
rect 3390 23590 3470 23670
rect 3690 23590 3770 23670
rect 4010 23590 4090 23670
rect 4330 23590 4410 23670
rect 4650 23590 4730 23670
rect 4950 23590 5030 23670
rect 5270 23590 5350 23670
rect 5590 23590 5670 23670
rect 5910 23590 5990 23670
rect 6210 23590 6290 23670
rect 6530 23590 6610 23670
rect 6850 23590 6930 23670
rect 7170 23590 7250 23670
rect 7470 23590 7550 23670
rect 7790 23590 7870 23670
rect 8110 23590 8190 23670
rect 8430 23590 8510 23670
rect 8730 23590 8810 23670
rect 9050 23590 9130 23670
rect 9370 23590 9450 23670
rect 9690 23590 9770 23670
rect 9990 23590 10070 23670
rect 10310 23590 10390 23670
rect 10630 23590 10710 23670
rect 10950 23590 11030 23670
rect 11250 23590 11330 23670
rect 11660 23590 11740 23670
rect 11960 23590 12040 23670
rect 160 23410 240 23490
rect 870 23410 950 23490
rect 1170 23410 1250 23490
rect 1490 23410 1570 23490
rect 1810 23410 1890 23490
rect 2130 23410 2210 23490
rect 2430 23410 2510 23490
rect 2750 23410 2830 23490
rect 3070 23410 3150 23490
rect 3390 23410 3470 23490
rect 3690 23410 3770 23490
rect 4010 23410 4090 23490
rect 4330 23410 4410 23490
rect 4650 23410 4730 23490
rect 4950 23410 5030 23490
rect 5270 23410 5350 23490
rect 5590 23410 5670 23490
rect 5910 23410 5990 23490
rect 6210 23410 6290 23490
rect 6530 23410 6610 23490
rect 6850 23410 6930 23490
rect 7170 23410 7250 23490
rect 7470 23410 7550 23490
rect 7790 23410 7870 23490
rect 8110 23410 8190 23490
rect 8430 23410 8510 23490
rect 8730 23410 8810 23490
rect 9050 23410 9130 23490
rect 9370 23410 9450 23490
rect 9690 23410 9770 23490
rect 9990 23410 10070 23490
rect 10310 23410 10390 23490
rect 10630 23410 10710 23490
rect 10950 23410 11030 23490
rect 11250 23410 11330 23490
rect 11660 23410 11740 23490
rect 11960 23410 12040 23490
rect 160 23230 240 23310
rect 870 23230 950 23310
rect 1170 23230 1250 23310
rect 1490 23230 1570 23310
rect 1810 23230 1890 23310
rect 2130 23230 2210 23310
rect 2430 23230 2510 23310
rect 2750 23230 2830 23310
rect 3070 23230 3150 23310
rect 3390 23230 3470 23310
rect 3690 23230 3770 23310
rect 4010 23230 4090 23310
rect 4330 23230 4410 23310
rect 4650 23230 4730 23310
rect 4950 23230 5030 23310
rect 5270 23230 5350 23310
rect 5590 23230 5670 23310
rect 5910 23230 5990 23310
rect 6210 23230 6290 23310
rect 6530 23230 6610 23310
rect 6850 23230 6930 23310
rect 7170 23230 7250 23310
rect 7470 23230 7550 23310
rect 7790 23230 7870 23310
rect 8110 23230 8190 23310
rect 8430 23230 8510 23310
rect 8730 23230 8810 23310
rect 9050 23230 9130 23310
rect 9370 23230 9450 23310
rect 9690 23230 9770 23310
rect 9990 23230 10070 23310
rect 10310 23230 10390 23310
rect 10630 23230 10710 23310
rect 10950 23230 11030 23310
rect 11250 23230 11330 23310
rect 11660 23230 11740 23310
rect 11960 23230 12040 23310
rect 160 23050 240 23130
rect 870 23050 950 23130
rect 1170 23050 1250 23130
rect 1490 23050 1570 23130
rect 1810 23050 1890 23130
rect 2130 23050 2210 23130
rect 2430 23050 2510 23130
rect 2750 23050 2830 23130
rect 3070 23050 3150 23130
rect 3390 23050 3470 23130
rect 3690 23050 3770 23130
rect 4010 23050 4090 23130
rect 4330 23050 4410 23130
rect 4650 23050 4730 23130
rect 4950 23050 5030 23130
rect 5270 23050 5350 23130
rect 5590 23050 5670 23130
rect 5910 23050 5990 23130
rect 6210 23050 6290 23130
rect 6530 23050 6610 23130
rect 6850 23050 6930 23130
rect 7170 23050 7250 23130
rect 7470 23050 7550 23130
rect 7790 23050 7870 23130
rect 8110 23050 8190 23130
rect 8430 23050 8510 23130
rect 8730 23050 8810 23130
rect 9050 23050 9130 23130
rect 9370 23050 9450 23130
rect 9690 23050 9770 23130
rect 9990 23050 10070 23130
rect 10310 23050 10390 23130
rect 10630 23050 10710 23130
rect 10950 23050 11030 23130
rect 11250 23050 11330 23130
rect 11660 23050 11740 23130
rect 11960 23050 12040 23130
rect 160 22870 240 22950
rect 870 22870 950 22950
rect 1170 22870 1250 22950
rect 1490 22870 1570 22950
rect 1810 22870 1890 22950
rect 2130 22870 2210 22950
rect 2430 22870 2510 22950
rect 2750 22870 2830 22950
rect 3070 22870 3150 22950
rect 3390 22870 3470 22950
rect 3690 22870 3770 22950
rect 4010 22870 4090 22950
rect 4330 22870 4410 22950
rect 4650 22870 4730 22950
rect 4950 22870 5030 22950
rect 5270 22870 5350 22950
rect 5590 22870 5670 22950
rect 5910 22870 5990 22950
rect 6210 22870 6290 22950
rect 6530 22870 6610 22950
rect 6850 22870 6930 22950
rect 7170 22870 7250 22950
rect 7470 22870 7550 22950
rect 7790 22870 7870 22950
rect 8110 22870 8190 22950
rect 8430 22870 8510 22950
rect 8730 22870 8810 22950
rect 9050 22870 9130 22950
rect 9370 22870 9450 22950
rect 9690 22870 9770 22950
rect 9990 22870 10070 22950
rect 10310 22870 10390 22950
rect 10630 22870 10710 22950
rect 10950 22870 11030 22950
rect 11250 22870 11330 22950
rect 11660 22870 11740 22950
rect 11960 22870 12040 22950
rect 160 22690 240 22770
rect 870 22690 950 22770
rect 1170 22690 1250 22770
rect 1490 22690 1570 22770
rect 1810 22690 1890 22770
rect 2130 22690 2210 22770
rect 2430 22690 2510 22770
rect 2750 22690 2830 22770
rect 3070 22690 3150 22770
rect 3390 22690 3470 22770
rect 3690 22690 3770 22770
rect 4010 22690 4090 22770
rect 4330 22690 4410 22770
rect 4650 22690 4730 22770
rect 4950 22690 5030 22770
rect 5270 22690 5350 22770
rect 5590 22690 5670 22770
rect 5910 22690 5990 22770
rect 6210 22690 6290 22770
rect 6530 22690 6610 22770
rect 6850 22690 6930 22770
rect 7170 22690 7250 22770
rect 7470 22690 7550 22770
rect 7790 22690 7870 22770
rect 8110 22690 8190 22770
rect 8430 22690 8510 22770
rect 8730 22690 8810 22770
rect 9050 22690 9130 22770
rect 9370 22690 9450 22770
rect 9690 22690 9770 22770
rect 9990 22690 10070 22770
rect 10310 22690 10390 22770
rect 10630 22690 10710 22770
rect 10950 22690 11030 22770
rect 11250 22690 11330 22770
rect 11660 22690 11740 22770
rect 11960 22690 12040 22770
rect 160 22510 240 22590
rect 870 22510 950 22590
rect 1170 22510 1250 22590
rect 1490 22510 1570 22590
rect 1810 22510 1890 22590
rect 2130 22510 2210 22590
rect 2430 22510 2510 22590
rect 2750 22510 2830 22590
rect 3070 22510 3150 22590
rect 3390 22510 3470 22590
rect 3690 22510 3770 22590
rect 4010 22510 4090 22590
rect 4330 22510 4410 22590
rect 4650 22510 4730 22590
rect 4950 22510 5030 22590
rect 5270 22510 5350 22590
rect 5590 22510 5670 22590
rect 5910 22510 5990 22590
rect 6210 22510 6290 22590
rect 6530 22510 6610 22590
rect 6850 22510 6930 22590
rect 7170 22510 7250 22590
rect 7470 22510 7550 22590
rect 7790 22510 7870 22590
rect 8110 22510 8190 22590
rect 8430 22510 8510 22590
rect 8730 22510 8810 22590
rect 9050 22510 9130 22590
rect 9370 22510 9450 22590
rect 9690 22510 9770 22590
rect 9990 22510 10070 22590
rect 10310 22510 10390 22590
rect 10630 22510 10710 22590
rect 10950 22510 11030 22590
rect 11250 22510 11330 22590
rect 11660 22510 11740 22590
rect 11960 22510 12040 22590
rect 160 22330 240 22410
rect 870 22330 950 22410
rect 1170 22330 1250 22410
rect 1490 22330 1570 22410
rect 1810 22330 1890 22410
rect 2130 22330 2210 22410
rect 2430 22330 2510 22410
rect 2750 22330 2830 22410
rect 3070 22330 3150 22410
rect 3390 22330 3470 22410
rect 3690 22330 3770 22410
rect 4010 22330 4090 22410
rect 4330 22330 4410 22410
rect 4650 22330 4730 22410
rect 4950 22330 5030 22410
rect 5270 22330 5350 22410
rect 5590 22330 5670 22410
rect 5910 22330 5990 22410
rect 6210 22330 6290 22410
rect 6530 22330 6610 22410
rect 6850 22330 6930 22410
rect 7170 22330 7250 22410
rect 7470 22330 7550 22410
rect 7790 22330 7870 22410
rect 8110 22330 8190 22410
rect 8430 22330 8510 22410
rect 8730 22330 8810 22410
rect 9050 22330 9130 22410
rect 9370 22330 9450 22410
rect 9690 22330 9770 22410
rect 9990 22330 10070 22410
rect 10310 22330 10390 22410
rect 10630 22330 10710 22410
rect 10950 22330 11030 22410
rect 11250 22330 11330 22410
rect 11660 22330 11740 22410
rect 11960 22330 12040 22410
rect 160 22150 240 22230
rect 870 22150 950 22230
rect 1170 22150 1250 22230
rect 1490 22150 1570 22230
rect 1810 22150 1890 22230
rect 2130 22150 2210 22230
rect 2430 22150 2510 22230
rect 2750 22150 2830 22230
rect 3070 22150 3150 22230
rect 3390 22150 3470 22230
rect 3690 22150 3770 22230
rect 4010 22150 4090 22230
rect 4330 22150 4410 22230
rect 4650 22150 4730 22230
rect 4950 22150 5030 22230
rect 5270 22150 5350 22230
rect 5590 22150 5670 22230
rect 5910 22150 5990 22230
rect 6210 22150 6290 22230
rect 6530 22150 6610 22230
rect 6850 22150 6930 22230
rect 7170 22150 7250 22230
rect 7470 22150 7550 22230
rect 7790 22150 7870 22230
rect 8110 22150 8190 22230
rect 8430 22150 8510 22230
rect 8730 22150 8810 22230
rect 9050 22150 9130 22230
rect 9370 22150 9450 22230
rect 9690 22150 9770 22230
rect 9990 22150 10070 22230
rect 10310 22150 10390 22230
rect 10630 22150 10710 22230
rect 10950 22150 11030 22230
rect 11250 22150 11330 22230
rect 11660 22150 11740 22230
rect 11960 22150 12040 22230
rect 160 21970 240 22050
rect 870 21970 950 22050
rect 1170 21970 1250 22050
rect 1490 21970 1570 22050
rect 1810 21970 1890 22050
rect 2130 21970 2210 22050
rect 2430 21970 2510 22050
rect 2750 21970 2830 22050
rect 3070 21970 3150 22050
rect 3390 21970 3470 22050
rect 3690 21970 3770 22050
rect 4010 21970 4090 22050
rect 4330 21970 4410 22050
rect 4650 21970 4730 22050
rect 4950 21970 5030 22050
rect 5270 21970 5350 22050
rect 5590 21970 5670 22050
rect 5910 21970 5990 22050
rect 6210 21970 6290 22050
rect 6530 21970 6610 22050
rect 6850 21970 6930 22050
rect 7170 21970 7250 22050
rect 7470 21970 7550 22050
rect 7790 21970 7870 22050
rect 8110 21970 8190 22050
rect 8430 21970 8510 22050
rect 8730 21970 8810 22050
rect 9050 21970 9130 22050
rect 9370 21970 9450 22050
rect 9690 21970 9770 22050
rect 9990 21970 10070 22050
rect 10310 21970 10390 22050
rect 10630 21970 10710 22050
rect 10950 21970 11030 22050
rect 11250 21970 11330 22050
rect 11660 21970 11740 22050
rect 11960 21970 12040 22050
rect 160 21790 240 21870
rect 870 21790 950 21870
rect 1170 21790 1250 21870
rect 1490 21790 1570 21870
rect 1810 21790 1890 21870
rect 2130 21790 2210 21870
rect 2430 21790 2510 21870
rect 2750 21790 2830 21870
rect 3070 21790 3150 21870
rect 3390 21790 3470 21870
rect 3690 21790 3770 21870
rect 4010 21790 4090 21870
rect 4330 21790 4410 21870
rect 4650 21790 4730 21870
rect 4950 21790 5030 21870
rect 5270 21790 5350 21870
rect 5590 21790 5670 21870
rect 5910 21790 5990 21870
rect 6210 21790 6290 21870
rect 6530 21790 6610 21870
rect 6850 21790 6930 21870
rect 7170 21790 7250 21870
rect 7470 21790 7550 21870
rect 7790 21790 7870 21870
rect 8110 21790 8190 21870
rect 8430 21790 8510 21870
rect 8730 21790 8810 21870
rect 9050 21790 9130 21870
rect 9370 21790 9450 21870
rect 9690 21790 9770 21870
rect 9990 21790 10070 21870
rect 10310 21790 10390 21870
rect 10630 21790 10710 21870
rect 10950 21790 11030 21870
rect 11250 21790 11330 21870
rect 11660 21790 11740 21870
rect 11960 21790 12040 21870
rect 160 21610 240 21690
rect 870 21610 950 21690
rect 1170 21610 1250 21690
rect 1490 21610 1570 21690
rect 1810 21610 1890 21690
rect 2130 21610 2210 21690
rect 2430 21610 2510 21690
rect 2750 21610 2830 21690
rect 3070 21610 3150 21690
rect 3390 21610 3470 21690
rect 3690 21610 3770 21690
rect 4010 21610 4090 21690
rect 4330 21610 4410 21690
rect 4650 21610 4730 21690
rect 4950 21610 5030 21690
rect 5270 21610 5350 21690
rect 5590 21610 5670 21690
rect 5910 21610 5990 21690
rect 6210 21610 6290 21690
rect 6530 21610 6610 21690
rect 6850 21610 6930 21690
rect 7170 21610 7250 21690
rect 7470 21610 7550 21690
rect 7790 21610 7870 21690
rect 8110 21610 8190 21690
rect 8430 21610 8510 21690
rect 8730 21610 8810 21690
rect 9050 21610 9130 21690
rect 9370 21610 9450 21690
rect 9690 21610 9770 21690
rect 9990 21610 10070 21690
rect 10310 21610 10390 21690
rect 10630 21610 10710 21690
rect 10950 21610 11030 21690
rect 11250 21610 11330 21690
rect 11660 21610 11740 21690
rect 11960 21610 12040 21690
rect 160 21430 240 21510
rect 870 21430 950 21510
rect 1170 21430 1250 21510
rect 1490 21430 1570 21510
rect 1810 21430 1890 21510
rect 2130 21430 2210 21510
rect 2430 21430 2510 21510
rect 2750 21430 2830 21510
rect 3070 21430 3150 21510
rect 3390 21430 3470 21510
rect 3690 21430 3770 21510
rect 4010 21430 4090 21510
rect 4330 21430 4410 21510
rect 4650 21430 4730 21510
rect 4950 21430 5030 21510
rect 5270 21430 5350 21510
rect 5590 21430 5670 21510
rect 5910 21430 5990 21510
rect 6210 21430 6290 21510
rect 6530 21430 6610 21510
rect 6850 21430 6930 21510
rect 7170 21430 7250 21510
rect 7470 21430 7550 21510
rect 7790 21430 7870 21510
rect 8110 21430 8190 21510
rect 8430 21430 8510 21510
rect 8730 21430 8810 21510
rect 9050 21430 9130 21510
rect 9370 21430 9450 21510
rect 9690 21430 9770 21510
rect 9990 21430 10070 21510
rect 10310 21430 10390 21510
rect 10630 21430 10710 21510
rect 10950 21430 11030 21510
rect 11250 21430 11330 21510
rect 11660 21430 11740 21510
rect 11960 21430 12040 21510
rect 160 21250 240 21330
rect 11660 21250 11740 21330
rect 11960 21250 12040 21330
rect 160 21070 240 21150
rect 11660 21070 11740 21150
rect 11960 21070 12040 21150
rect 160 20890 240 20970
rect 11660 20890 11740 20970
rect 11960 20890 12040 20970
rect 160 20710 240 20790
rect 11660 20710 11740 20790
rect 11960 20710 12040 20790
rect 160 20530 240 20610
rect 11660 20530 11740 20610
rect 11960 20530 12040 20610
rect 285 19740 365 19820
rect 285 19580 365 19660
rect 285 19420 365 19500
rect 285 19260 365 19340
rect 285 19100 365 19180
rect 11685 18285 11765 18365
rect 11865 18285 11945 18365
rect 11685 18105 11765 18185
rect 11865 18105 11945 18185
rect 11685 17925 11765 18005
rect 11865 17925 11945 18005
rect 11685 17745 11765 17825
rect 11865 17745 11945 17825
rect 11685 17565 11765 17645
rect 11865 17565 11945 17645
rect 160 16790 240 16870
rect 11660 16790 11740 16870
rect 11960 16790 12040 16870
rect 160 16610 240 16690
rect 11660 16610 11740 16690
rect 11960 16610 12040 16690
rect 160 16430 240 16510
rect 11660 16430 11740 16510
rect 11960 16430 12040 16510
rect 160 16250 240 16330
rect 11660 16250 11740 16330
rect 11960 16250 12040 16330
rect 160 16070 240 16150
rect 11660 16070 11740 16150
rect 11960 16070 12040 16150
rect 160 15890 240 15970
rect 870 15890 950 15970
rect 1170 15890 1250 15970
rect 1510 15890 1590 15970
rect 1810 15890 1890 15970
rect 2130 15890 2210 15970
rect 2430 15890 2510 15970
rect 2770 15890 2850 15970
rect 3070 15890 3150 15970
rect 3390 15890 3470 15970
rect 3690 15890 3770 15970
rect 4030 15890 4110 15970
rect 4330 15890 4410 15970
rect 4650 15890 4730 15970
rect 4950 15890 5030 15970
rect 5290 15890 5370 15970
rect 5590 15890 5670 15970
rect 5910 15890 5990 15970
rect 6210 15890 6290 15970
rect 6550 15890 6630 15970
rect 6850 15890 6930 15970
rect 7170 15890 7250 15970
rect 7470 15890 7550 15970
rect 7810 15890 7890 15970
rect 8110 15890 8190 15970
rect 8430 15890 8510 15970
rect 8730 15890 8810 15970
rect 9070 15890 9150 15970
rect 9370 15890 9450 15970
rect 9690 15890 9770 15970
rect 9990 15890 10070 15970
rect 10330 15890 10410 15970
rect 10630 15890 10710 15970
rect 10950 15890 11030 15970
rect 11250 15890 11330 15970
rect 11660 15890 11740 15970
rect 11960 15890 12040 15970
rect 160 15710 240 15790
rect 870 15710 950 15790
rect 1170 15710 1250 15790
rect 1510 15710 1590 15790
rect 1810 15710 1890 15790
rect 2130 15710 2210 15790
rect 2430 15710 2510 15790
rect 2770 15710 2850 15790
rect 3070 15710 3150 15790
rect 3390 15710 3470 15790
rect 3690 15710 3770 15790
rect 4030 15710 4110 15790
rect 4330 15710 4410 15790
rect 4650 15710 4730 15790
rect 4950 15710 5030 15790
rect 5290 15710 5370 15790
rect 5590 15710 5670 15790
rect 5910 15710 5990 15790
rect 6210 15710 6290 15790
rect 6550 15710 6630 15790
rect 6850 15710 6930 15790
rect 7170 15710 7250 15790
rect 7470 15710 7550 15790
rect 7810 15710 7890 15790
rect 8110 15710 8190 15790
rect 8430 15710 8510 15790
rect 8730 15710 8810 15790
rect 9070 15710 9150 15790
rect 9370 15710 9450 15790
rect 9690 15710 9770 15790
rect 9990 15710 10070 15790
rect 10330 15710 10410 15790
rect 10630 15710 10710 15790
rect 10950 15710 11030 15790
rect 11250 15710 11330 15790
rect 11660 15710 11740 15790
rect 11960 15710 12040 15790
rect 160 15530 240 15610
rect 870 15530 950 15610
rect 1170 15530 1250 15610
rect 1510 15530 1590 15610
rect 1810 15530 1890 15610
rect 2130 15530 2210 15610
rect 2430 15530 2510 15610
rect 2770 15530 2850 15610
rect 3070 15530 3150 15610
rect 3390 15530 3470 15610
rect 3690 15530 3770 15610
rect 4030 15530 4110 15610
rect 4330 15530 4410 15610
rect 4650 15530 4730 15610
rect 4950 15530 5030 15610
rect 5290 15530 5370 15610
rect 5590 15530 5670 15610
rect 5910 15530 5990 15610
rect 6210 15530 6290 15610
rect 6550 15530 6630 15610
rect 6850 15530 6930 15610
rect 7170 15530 7250 15610
rect 7470 15530 7550 15610
rect 7810 15530 7890 15610
rect 8110 15530 8190 15610
rect 8430 15530 8510 15610
rect 8730 15530 8810 15610
rect 9070 15530 9150 15610
rect 9370 15530 9450 15610
rect 9690 15530 9770 15610
rect 9990 15530 10070 15610
rect 10330 15530 10410 15610
rect 10630 15530 10710 15610
rect 10950 15530 11030 15610
rect 11250 15530 11330 15610
rect 11660 15530 11740 15610
rect 11960 15530 12040 15610
rect 160 15350 240 15430
rect 870 15350 950 15430
rect 1170 15350 1250 15430
rect 1510 15350 1590 15430
rect 1810 15350 1890 15430
rect 2130 15350 2210 15430
rect 2430 15350 2510 15430
rect 2770 15350 2850 15430
rect 3070 15350 3150 15430
rect 3390 15350 3470 15430
rect 3690 15350 3770 15430
rect 4030 15350 4110 15430
rect 4330 15350 4410 15430
rect 4650 15350 4730 15430
rect 4950 15350 5030 15430
rect 5290 15350 5370 15430
rect 5590 15350 5670 15430
rect 5910 15350 5990 15430
rect 6210 15350 6290 15430
rect 6550 15350 6630 15430
rect 6850 15350 6930 15430
rect 7170 15350 7250 15430
rect 7470 15350 7550 15430
rect 7810 15350 7890 15430
rect 8110 15350 8190 15430
rect 8430 15350 8510 15430
rect 8730 15350 8810 15430
rect 9070 15350 9150 15430
rect 9370 15350 9450 15430
rect 9690 15350 9770 15430
rect 9990 15350 10070 15430
rect 10330 15350 10410 15430
rect 10630 15350 10710 15430
rect 10950 15350 11030 15430
rect 11250 15350 11330 15430
rect 11660 15350 11740 15430
rect 11960 15350 12040 15430
rect 160 15170 240 15250
rect 870 15170 950 15250
rect 1170 15170 1250 15250
rect 1510 15170 1590 15250
rect 1810 15170 1890 15250
rect 2130 15170 2210 15250
rect 2430 15170 2510 15250
rect 2770 15170 2850 15250
rect 3070 15170 3150 15250
rect 3390 15170 3470 15250
rect 3690 15170 3770 15250
rect 4030 15170 4110 15250
rect 4330 15170 4410 15250
rect 4650 15170 4730 15250
rect 4950 15170 5030 15250
rect 5290 15170 5370 15250
rect 5590 15170 5670 15250
rect 5910 15170 5990 15250
rect 6210 15170 6290 15250
rect 6550 15170 6630 15250
rect 6850 15170 6930 15250
rect 7170 15170 7250 15250
rect 7470 15170 7550 15250
rect 7810 15170 7890 15250
rect 8110 15170 8190 15250
rect 8430 15170 8510 15250
rect 8730 15170 8810 15250
rect 9070 15170 9150 15250
rect 9370 15170 9450 15250
rect 9690 15170 9770 15250
rect 9990 15170 10070 15250
rect 10330 15170 10410 15250
rect 10630 15170 10710 15250
rect 10950 15170 11030 15250
rect 11250 15170 11330 15250
rect 11660 15170 11740 15250
rect 11960 15170 12040 15250
rect 160 14990 240 15070
rect 870 14990 950 15070
rect 1170 14990 1250 15070
rect 1510 14990 1590 15070
rect 1810 14990 1890 15070
rect 2130 14990 2210 15070
rect 2430 14990 2510 15070
rect 2770 14990 2850 15070
rect 3070 14990 3150 15070
rect 3390 14990 3470 15070
rect 3690 14990 3770 15070
rect 4030 14990 4110 15070
rect 4330 14990 4410 15070
rect 4650 14990 4730 15070
rect 4950 14990 5030 15070
rect 5290 14990 5370 15070
rect 5590 14990 5670 15070
rect 5910 14990 5990 15070
rect 6210 14990 6290 15070
rect 6550 14990 6630 15070
rect 6850 14990 6930 15070
rect 7170 14990 7250 15070
rect 7470 14990 7550 15070
rect 7810 14990 7890 15070
rect 8110 14990 8190 15070
rect 8430 14990 8510 15070
rect 8730 14990 8810 15070
rect 9070 14990 9150 15070
rect 9370 14990 9450 15070
rect 9690 14990 9770 15070
rect 9990 14990 10070 15070
rect 10330 14990 10410 15070
rect 10630 14990 10710 15070
rect 10950 14990 11030 15070
rect 11250 14990 11330 15070
rect 11660 14990 11740 15070
rect 11960 14990 12040 15070
rect 160 14810 240 14890
rect 870 14810 950 14890
rect 1170 14810 1250 14890
rect 1510 14810 1590 14890
rect 1810 14810 1890 14890
rect 2130 14810 2210 14890
rect 2430 14810 2510 14890
rect 2770 14810 2850 14890
rect 3070 14810 3150 14890
rect 3390 14810 3470 14890
rect 3690 14810 3770 14890
rect 4030 14810 4110 14890
rect 4330 14810 4410 14890
rect 4650 14810 4730 14890
rect 4950 14810 5030 14890
rect 5290 14810 5370 14890
rect 5590 14810 5670 14890
rect 5910 14810 5990 14890
rect 6210 14810 6290 14890
rect 6550 14810 6630 14890
rect 6850 14810 6930 14890
rect 7170 14810 7250 14890
rect 7470 14810 7550 14890
rect 7810 14810 7890 14890
rect 8110 14810 8190 14890
rect 8430 14810 8510 14890
rect 8730 14810 8810 14890
rect 9070 14810 9150 14890
rect 9370 14810 9450 14890
rect 9690 14810 9770 14890
rect 9990 14810 10070 14890
rect 10330 14810 10410 14890
rect 10630 14810 10710 14890
rect 10950 14810 11030 14890
rect 11250 14810 11330 14890
rect 11660 14810 11740 14890
rect 11960 14810 12040 14890
rect 160 14630 240 14710
rect 870 14630 950 14710
rect 1170 14630 1250 14710
rect 1510 14630 1590 14710
rect 1810 14630 1890 14710
rect 2130 14630 2210 14710
rect 2430 14630 2510 14710
rect 2770 14630 2850 14710
rect 3070 14630 3150 14710
rect 3390 14630 3470 14710
rect 3690 14630 3770 14710
rect 4030 14630 4110 14710
rect 4330 14630 4410 14710
rect 4650 14630 4730 14710
rect 4950 14630 5030 14710
rect 5290 14630 5370 14710
rect 5590 14630 5670 14710
rect 5910 14630 5990 14710
rect 6210 14630 6290 14710
rect 6550 14630 6630 14710
rect 6850 14630 6930 14710
rect 7170 14630 7250 14710
rect 7470 14630 7550 14710
rect 7810 14630 7890 14710
rect 8110 14630 8190 14710
rect 8430 14630 8510 14710
rect 8730 14630 8810 14710
rect 9070 14630 9150 14710
rect 9370 14630 9450 14710
rect 9690 14630 9770 14710
rect 9990 14630 10070 14710
rect 10330 14630 10410 14710
rect 10630 14630 10710 14710
rect 10950 14630 11030 14710
rect 11250 14630 11330 14710
rect 11660 14630 11740 14710
rect 11960 14630 12040 14710
rect 160 14450 240 14530
rect 870 14450 950 14530
rect 1170 14450 1250 14530
rect 1510 14450 1590 14530
rect 1810 14450 1890 14530
rect 2130 14450 2210 14530
rect 2430 14450 2510 14530
rect 2770 14450 2850 14530
rect 3070 14450 3150 14530
rect 3390 14450 3470 14530
rect 3690 14450 3770 14530
rect 4030 14450 4110 14530
rect 4330 14450 4410 14530
rect 4650 14450 4730 14530
rect 4950 14450 5030 14530
rect 5290 14450 5370 14530
rect 5590 14450 5670 14530
rect 5910 14450 5990 14530
rect 6210 14450 6290 14530
rect 6550 14450 6630 14530
rect 6850 14450 6930 14530
rect 7170 14450 7250 14530
rect 7470 14450 7550 14530
rect 7810 14450 7890 14530
rect 8110 14450 8190 14530
rect 8430 14450 8510 14530
rect 8730 14450 8810 14530
rect 9070 14450 9150 14530
rect 9370 14450 9450 14530
rect 9690 14450 9770 14530
rect 9990 14450 10070 14530
rect 10330 14450 10410 14530
rect 10630 14450 10710 14530
rect 10950 14450 11030 14530
rect 11250 14450 11330 14530
rect 11660 14450 11740 14530
rect 11960 14450 12040 14530
rect 160 14270 240 14350
rect 870 14270 950 14350
rect 1170 14270 1250 14350
rect 1510 14270 1590 14350
rect 1810 14270 1890 14350
rect 2130 14270 2210 14350
rect 2430 14270 2510 14350
rect 2770 14270 2850 14350
rect 3070 14270 3150 14350
rect 3390 14270 3470 14350
rect 3690 14270 3770 14350
rect 4030 14270 4110 14350
rect 4330 14270 4410 14350
rect 4650 14270 4730 14350
rect 4950 14270 5030 14350
rect 5290 14270 5370 14350
rect 5590 14270 5670 14350
rect 5910 14270 5990 14350
rect 6210 14270 6290 14350
rect 6550 14270 6630 14350
rect 6850 14270 6930 14350
rect 7170 14270 7250 14350
rect 7470 14270 7550 14350
rect 7810 14270 7890 14350
rect 8110 14270 8190 14350
rect 8430 14270 8510 14350
rect 8730 14270 8810 14350
rect 9070 14270 9150 14350
rect 9370 14270 9450 14350
rect 9690 14270 9770 14350
rect 9990 14270 10070 14350
rect 10330 14270 10410 14350
rect 10630 14270 10710 14350
rect 10950 14270 11030 14350
rect 11250 14270 11330 14350
rect 11660 14270 11740 14350
rect 11960 14270 12040 14350
rect 160 14090 240 14170
rect 870 14090 950 14170
rect 1170 14090 1250 14170
rect 1510 14090 1590 14170
rect 1810 14090 1890 14170
rect 2130 14090 2210 14170
rect 2430 14090 2510 14170
rect 2770 14090 2850 14170
rect 3070 14090 3150 14170
rect 3390 14090 3470 14170
rect 3690 14090 3770 14170
rect 4030 14090 4110 14170
rect 4330 14090 4410 14170
rect 4650 14090 4730 14170
rect 4950 14090 5030 14170
rect 5290 14090 5370 14170
rect 5590 14090 5670 14170
rect 5910 14090 5990 14170
rect 6210 14090 6290 14170
rect 6550 14090 6630 14170
rect 6850 14090 6930 14170
rect 7170 14090 7250 14170
rect 7470 14090 7550 14170
rect 7810 14090 7890 14170
rect 8110 14090 8190 14170
rect 8430 14090 8510 14170
rect 8730 14090 8810 14170
rect 9070 14090 9150 14170
rect 9370 14090 9450 14170
rect 9690 14090 9770 14170
rect 9990 14090 10070 14170
rect 10330 14090 10410 14170
rect 10630 14090 10710 14170
rect 10950 14090 11030 14170
rect 11250 14090 11330 14170
rect 11660 14090 11740 14170
rect 11960 14090 12040 14170
rect 160 13910 240 13990
rect 870 13910 950 13990
rect 1170 13910 1250 13990
rect 1510 13910 1590 13990
rect 1810 13910 1890 13990
rect 2130 13910 2210 13990
rect 2430 13910 2510 13990
rect 2770 13910 2850 13990
rect 3070 13910 3150 13990
rect 3390 13910 3470 13990
rect 3690 13910 3770 13990
rect 4030 13910 4110 13990
rect 4330 13910 4410 13990
rect 4650 13910 4730 13990
rect 4950 13910 5030 13990
rect 5290 13910 5370 13990
rect 5590 13910 5670 13990
rect 5910 13910 5990 13990
rect 6210 13910 6290 13990
rect 6550 13910 6630 13990
rect 6850 13910 6930 13990
rect 7170 13910 7250 13990
rect 7470 13910 7550 13990
rect 7810 13910 7890 13990
rect 8110 13910 8190 13990
rect 8430 13910 8510 13990
rect 8730 13910 8810 13990
rect 9070 13910 9150 13990
rect 9370 13910 9450 13990
rect 9690 13910 9770 13990
rect 9990 13910 10070 13990
rect 10330 13910 10410 13990
rect 10630 13910 10710 13990
rect 10950 13910 11030 13990
rect 11250 13910 11330 13990
rect 11660 13910 11740 13990
rect 11960 13910 12040 13990
rect 160 13730 240 13810
rect 870 13730 950 13810
rect 1170 13730 1250 13810
rect 1510 13730 1590 13810
rect 1810 13730 1890 13810
rect 2130 13730 2210 13810
rect 2430 13730 2510 13810
rect 2770 13730 2850 13810
rect 3070 13730 3150 13810
rect 3390 13730 3470 13810
rect 3690 13730 3770 13810
rect 4030 13730 4110 13810
rect 4330 13730 4410 13810
rect 4650 13730 4730 13810
rect 4950 13730 5030 13810
rect 5290 13730 5370 13810
rect 5590 13730 5670 13810
rect 5910 13730 5990 13810
rect 6210 13730 6290 13810
rect 6550 13730 6630 13810
rect 6850 13730 6930 13810
rect 7170 13730 7250 13810
rect 7470 13730 7550 13810
rect 7810 13730 7890 13810
rect 8110 13730 8190 13810
rect 8430 13730 8510 13810
rect 8730 13730 8810 13810
rect 9070 13730 9150 13810
rect 9370 13730 9450 13810
rect 9690 13730 9770 13810
rect 9990 13730 10070 13810
rect 10330 13730 10410 13810
rect 10630 13730 10710 13810
rect 10950 13730 11030 13810
rect 11250 13730 11330 13810
rect 11660 13730 11740 13810
rect 11960 13730 12040 13810
rect 160 13550 240 13630
rect 870 13550 950 13630
rect 1170 13550 1250 13630
rect 1510 13550 1590 13630
rect 1810 13550 1890 13630
rect 2130 13550 2210 13630
rect 2430 13550 2510 13630
rect 2770 13550 2850 13630
rect 3070 13550 3150 13630
rect 3390 13550 3470 13630
rect 3690 13550 3770 13630
rect 4030 13550 4110 13630
rect 4330 13550 4410 13630
rect 4650 13550 4730 13630
rect 4950 13550 5030 13630
rect 5290 13550 5370 13630
rect 5590 13550 5670 13630
rect 5910 13550 5990 13630
rect 6210 13550 6290 13630
rect 6550 13550 6630 13630
rect 6850 13550 6930 13630
rect 7170 13550 7250 13630
rect 7470 13550 7550 13630
rect 7810 13550 7890 13630
rect 8110 13550 8190 13630
rect 8430 13550 8510 13630
rect 8730 13550 8810 13630
rect 9070 13550 9150 13630
rect 9370 13550 9450 13630
rect 9690 13550 9770 13630
rect 9990 13550 10070 13630
rect 10330 13550 10410 13630
rect 10630 13550 10710 13630
rect 10950 13550 11030 13630
rect 11250 13550 11330 13630
rect 11660 13550 11740 13630
rect 11960 13550 12040 13630
rect 160 13370 240 13450
rect 870 13370 950 13450
rect 1170 13370 1250 13450
rect 1510 13370 1590 13450
rect 1810 13370 1890 13450
rect 2130 13370 2210 13450
rect 2430 13370 2510 13450
rect 2770 13370 2850 13450
rect 3070 13370 3150 13450
rect 3390 13370 3470 13450
rect 3690 13370 3770 13450
rect 4030 13370 4110 13450
rect 4330 13370 4410 13450
rect 4650 13370 4730 13450
rect 4950 13370 5030 13450
rect 5290 13370 5370 13450
rect 5590 13370 5670 13450
rect 5910 13370 5990 13450
rect 6210 13370 6290 13450
rect 6550 13370 6630 13450
rect 6850 13370 6930 13450
rect 7170 13370 7250 13450
rect 7470 13370 7550 13450
rect 7810 13370 7890 13450
rect 8110 13370 8190 13450
rect 8430 13370 8510 13450
rect 8730 13370 8810 13450
rect 9070 13370 9150 13450
rect 9370 13370 9450 13450
rect 9690 13370 9770 13450
rect 9990 13370 10070 13450
rect 10330 13370 10410 13450
rect 10630 13370 10710 13450
rect 10950 13370 11030 13450
rect 11250 13370 11330 13450
rect 11660 13370 11740 13450
rect 11960 13370 12040 13450
rect 160 13190 240 13270
rect 870 13190 950 13270
rect 1170 13190 1250 13270
rect 1510 13190 1590 13270
rect 1810 13190 1890 13270
rect 2130 13190 2210 13270
rect 2430 13190 2510 13270
rect 2770 13190 2850 13270
rect 3070 13190 3150 13270
rect 3390 13190 3470 13270
rect 3690 13190 3770 13270
rect 4030 13190 4110 13270
rect 4330 13190 4410 13270
rect 4650 13190 4730 13270
rect 4950 13190 5030 13270
rect 5290 13190 5370 13270
rect 5590 13190 5670 13270
rect 5910 13190 5990 13270
rect 6210 13190 6290 13270
rect 6550 13190 6630 13270
rect 6850 13190 6930 13270
rect 7170 13190 7250 13270
rect 7470 13190 7550 13270
rect 7810 13190 7890 13270
rect 8110 13190 8190 13270
rect 8430 13190 8510 13270
rect 8730 13190 8810 13270
rect 9070 13190 9150 13270
rect 9370 13190 9450 13270
rect 9690 13190 9770 13270
rect 9990 13190 10070 13270
rect 10330 13190 10410 13270
rect 10630 13190 10710 13270
rect 10950 13190 11030 13270
rect 11250 13190 11330 13270
rect 11660 13190 11740 13270
rect 11960 13190 12040 13270
rect 160 13010 240 13090
rect 870 13010 950 13090
rect 1170 13010 1250 13090
rect 1510 13010 1590 13090
rect 1810 13010 1890 13090
rect 2130 13010 2210 13090
rect 2430 13010 2510 13090
rect 2770 13010 2850 13090
rect 3070 13010 3150 13090
rect 3390 13010 3470 13090
rect 3690 13010 3770 13090
rect 4030 13010 4110 13090
rect 4330 13010 4410 13090
rect 4650 13010 4730 13090
rect 4950 13010 5030 13090
rect 5290 13010 5370 13090
rect 5590 13010 5670 13090
rect 5910 13010 5990 13090
rect 6210 13010 6290 13090
rect 6550 13010 6630 13090
rect 6850 13010 6930 13090
rect 7170 13010 7250 13090
rect 7470 13010 7550 13090
rect 7810 13010 7890 13090
rect 8110 13010 8190 13090
rect 8430 13010 8510 13090
rect 8730 13010 8810 13090
rect 9070 13010 9150 13090
rect 9370 13010 9450 13090
rect 9690 13010 9770 13090
rect 9990 13010 10070 13090
rect 10330 13010 10410 13090
rect 10630 13010 10710 13090
rect 10950 13010 11030 13090
rect 11250 13010 11330 13090
rect 11660 13010 11740 13090
rect 11960 13010 12040 13090
rect 160 12830 240 12910
rect 870 12830 950 12910
rect 1170 12830 1250 12910
rect 1510 12830 1590 12910
rect 1810 12830 1890 12910
rect 2130 12830 2210 12910
rect 2430 12830 2510 12910
rect 2770 12830 2850 12910
rect 3070 12830 3150 12910
rect 3390 12830 3470 12910
rect 3690 12830 3770 12910
rect 4030 12830 4110 12910
rect 4330 12830 4410 12910
rect 4650 12830 4730 12910
rect 4950 12830 5030 12910
rect 5290 12830 5370 12910
rect 5590 12830 5670 12910
rect 5910 12830 5990 12910
rect 6210 12830 6290 12910
rect 6550 12830 6630 12910
rect 6850 12830 6930 12910
rect 7170 12830 7250 12910
rect 7470 12830 7550 12910
rect 7810 12830 7890 12910
rect 8110 12830 8190 12910
rect 8430 12830 8510 12910
rect 8730 12830 8810 12910
rect 9070 12830 9150 12910
rect 9370 12830 9450 12910
rect 9690 12830 9770 12910
rect 9990 12830 10070 12910
rect 10330 12830 10410 12910
rect 10630 12830 10710 12910
rect 10950 12830 11030 12910
rect 11250 12830 11330 12910
rect 11660 12830 11740 12910
rect 11960 12830 12040 12910
rect 160 12650 240 12730
rect 870 12650 950 12730
rect 1170 12650 1250 12730
rect 1510 12650 1590 12730
rect 1810 12650 1890 12730
rect 2130 12650 2210 12730
rect 2430 12650 2510 12730
rect 2770 12650 2850 12730
rect 3070 12650 3150 12730
rect 3390 12650 3470 12730
rect 3690 12650 3770 12730
rect 4030 12650 4110 12730
rect 4330 12650 4410 12730
rect 4650 12650 4730 12730
rect 4950 12650 5030 12730
rect 5290 12650 5370 12730
rect 5590 12650 5670 12730
rect 5910 12650 5990 12730
rect 6210 12650 6290 12730
rect 6550 12650 6630 12730
rect 6850 12650 6930 12730
rect 7170 12650 7250 12730
rect 7470 12650 7550 12730
rect 7810 12650 7890 12730
rect 8110 12650 8190 12730
rect 8430 12650 8510 12730
rect 8730 12650 8810 12730
rect 9070 12650 9150 12730
rect 9370 12650 9450 12730
rect 9690 12650 9770 12730
rect 9990 12650 10070 12730
rect 10330 12650 10410 12730
rect 10630 12650 10710 12730
rect 10950 12650 11030 12730
rect 11250 12650 11330 12730
rect 11660 12650 11740 12730
rect 11960 12650 12040 12730
rect 160 12470 240 12550
rect 870 12470 950 12550
rect 1170 12470 1250 12550
rect 1510 12470 1590 12550
rect 1810 12470 1890 12550
rect 2130 12470 2210 12550
rect 2430 12470 2510 12550
rect 2770 12470 2850 12550
rect 3070 12470 3150 12550
rect 3390 12470 3470 12550
rect 3690 12470 3770 12550
rect 4030 12470 4110 12550
rect 4330 12470 4410 12550
rect 4650 12470 4730 12550
rect 4950 12470 5030 12550
rect 5290 12470 5370 12550
rect 5590 12470 5670 12550
rect 5910 12470 5990 12550
rect 6210 12470 6290 12550
rect 6550 12470 6630 12550
rect 6850 12470 6930 12550
rect 7170 12470 7250 12550
rect 7470 12470 7550 12550
rect 7810 12470 7890 12550
rect 8110 12470 8190 12550
rect 8430 12470 8510 12550
rect 8730 12470 8810 12550
rect 9070 12470 9150 12550
rect 9370 12470 9450 12550
rect 9690 12470 9770 12550
rect 9990 12470 10070 12550
rect 10330 12470 10410 12550
rect 10630 12470 10710 12550
rect 10950 12470 11030 12550
rect 11250 12470 11330 12550
rect 11660 12470 11740 12550
rect 11960 12470 12040 12550
rect 160 12290 240 12370
rect 870 12290 950 12370
rect 1170 12290 1250 12370
rect 1510 12290 1590 12370
rect 1810 12290 1890 12370
rect 2130 12290 2210 12370
rect 2430 12290 2510 12370
rect 2770 12290 2850 12370
rect 3070 12290 3150 12370
rect 3390 12290 3470 12370
rect 3690 12290 3770 12370
rect 4030 12290 4110 12370
rect 4330 12290 4410 12370
rect 4650 12290 4730 12370
rect 4950 12290 5030 12370
rect 5290 12290 5370 12370
rect 5590 12290 5670 12370
rect 5910 12290 5990 12370
rect 6210 12290 6290 12370
rect 6550 12290 6630 12370
rect 6850 12290 6930 12370
rect 7170 12290 7250 12370
rect 7470 12290 7550 12370
rect 7810 12290 7890 12370
rect 8110 12290 8190 12370
rect 8430 12290 8510 12370
rect 8730 12290 8810 12370
rect 9070 12290 9150 12370
rect 9370 12290 9450 12370
rect 9690 12290 9770 12370
rect 9990 12290 10070 12370
rect 10330 12290 10410 12370
rect 10630 12290 10710 12370
rect 10950 12290 11030 12370
rect 11250 12290 11330 12370
rect 11660 12290 11740 12370
rect 11960 12290 12040 12370
rect 160 12110 240 12190
rect 870 12110 950 12190
rect 1170 12110 1250 12190
rect 1510 12110 1590 12190
rect 1810 12110 1890 12190
rect 2130 12110 2210 12190
rect 2430 12110 2510 12190
rect 2770 12110 2850 12190
rect 3070 12110 3150 12190
rect 3390 12110 3470 12190
rect 3690 12110 3770 12190
rect 4030 12110 4110 12190
rect 4330 12110 4410 12190
rect 4650 12110 4730 12190
rect 4950 12110 5030 12190
rect 5290 12110 5370 12190
rect 5590 12110 5670 12190
rect 5910 12110 5990 12190
rect 6210 12110 6290 12190
rect 6550 12110 6630 12190
rect 6850 12110 6930 12190
rect 7170 12110 7250 12190
rect 7470 12110 7550 12190
rect 7810 12110 7890 12190
rect 8110 12110 8190 12190
rect 8430 12110 8510 12190
rect 8730 12110 8810 12190
rect 9070 12110 9150 12190
rect 9370 12110 9450 12190
rect 9690 12110 9770 12190
rect 9990 12110 10070 12190
rect 10330 12110 10410 12190
rect 10630 12110 10710 12190
rect 10950 12110 11030 12190
rect 11250 12110 11330 12190
rect 11660 12110 11740 12190
rect 11960 12110 12040 12190
rect 160 11930 240 12010
rect 870 11930 950 12010
rect 1170 11930 1250 12010
rect 1510 11930 1590 12010
rect 1810 11930 1890 12010
rect 2130 11930 2210 12010
rect 2430 11930 2510 12010
rect 2770 11930 2850 12010
rect 3070 11930 3150 12010
rect 3390 11930 3470 12010
rect 3690 11930 3770 12010
rect 4030 11930 4110 12010
rect 4330 11930 4410 12010
rect 4650 11930 4730 12010
rect 4950 11930 5030 12010
rect 5290 11930 5370 12010
rect 5590 11930 5670 12010
rect 5910 11930 5990 12010
rect 6210 11930 6290 12010
rect 6550 11930 6630 12010
rect 6850 11930 6930 12010
rect 7170 11930 7250 12010
rect 7470 11930 7550 12010
rect 7810 11930 7890 12010
rect 8110 11930 8190 12010
rect 8430 11930 8510 12010
rect 8730 11930 8810 12010
rect 9070 11930 9150 12010
rect 9370 11930 9450 12010
rect 9690 11930 9770 12010
rect 9990 11930 10070 12010
rect 10330 11930 10410 12010
rect 10630 11930 10710 12010
rect 10950 11930 11030 12010
rect 11250 11930 11330 12010
rect 11660 11930 11740 12010
rect 11960 11930 12040 12010
rect 160 11750 240 11830
rect 870 11750 950 11830
rect 1170 11750 1250 11830
rect 1510 11750 1590 11830
rect 1810 11750 1890 11830
rect 2130 11750 2210 11830
rect 2430 11750 2510 11830
rect 2770 11750 2850 11830
rect 3070 11750 3150 11830
rect 3390 11750 3470 11830
rect 3690 11750 3770 11830
rect 4030 11750 4110 11830
rect 4330 11750 4410 11830
rect 4650 11750 4730 11830
rect 4950 11750 5030 11830
rect 5290 11750 5370 11830
rect 5590 11750 5670 11830
rect 5910 11750 5990 11830
rect 6210 11750 6290 11830
rect 6550 11750 6630 11830
rect 6850 11750 6930 11830
rect 7170 11750 7250 11830
rect 7470 11750 7550 11830
rect 7810 11750 7890 11830
rect 8110 11750 8190 11830
rect 8430 11750 8510 11830
rect 8730 11750 8810 11830
rect 9070 11750 9150 11830
rect 9370 11750 9450 11830
rect 9690 11750 9770 11830
rect 9990 11750 10070 11830
rect 10330 11750 10410 11830
rect 10630 11750 10710 11830
rect 10950 11750 11030 11830
rect 11250 11750 11330 11830
rect 11660 11750 11740 11830
rect 11960 11750 12040 11830
rect 160 11570 240 11650
rect 870 11570 950 11650
rect 1170 11570 1250 11650
rect 1510 11570 1590 11650
rect 1810 11570 1890 11650
rect 2130 11570 2210 11650
rect 2430 11570 2510 11650
rect 2770 11570 2850 11650
rect 3070 11570 3150 11650
rect 3390 11570 3470 11650
rect 3690 11570 3770 11650
rect 4030 11570 4110 11650
rect 4330 11570 4410 11650
rect 4650 11570 4730 11650
rect 4950 11570 5030 11650
rect 5290 11570 5370 11650
rect 5590 11570 5670 11650
rect 5910 11570 5990 11650
rect 6210 11570 6290 11650
rect 6550 11570 6630 11650
rect 6850 11570 6930 11650
rect 7170 11570 7250 11650
rect 7470 11570 7550 11650
rect 7810 11570 7890 11650
rect 8110 11570 8190 11650
rect 8430 11570 8510 11650
rect 8730 11570 8810 11650
rect 9070 11570 9150 11650
rect 9370 11570 9450 11650
rect 9690 11570 9770 11650
rect 9990 11570 10070 11650
rect 10330 11570 10410 11650
rect 10630 11570 10710 11650
rect 10950 11570 11030 11650
rect 11250 11570 11330 11650
rect 11660 11570 11740 11650
rect 11960 11570 12040 11650
rect 160 11390 240 11470
rect 870 11390 950 11470
rect 1170 11390 1250 11470
rect 1510 11390 1590 11470
rect 1810 11390 1890 11470
rect 2130 11390 2210 11470
rect 2430 11390 2510 11470
rect 2770 11390 2850 11470
rect 3070 11390 3150 11470
rect 3390 11390 3470 11470
rect 3690 11390 3770 11470
rect 4030 11390 4110 11470
rect 4330 11390 4410 11470
rect 4650 11390 4730 11470
rect 4950 11390 5030 11470
rect 5290 11390 5370 11470
rect 5590 11390 5670 11470
rect 5910 11390 5990 11470
rect 6210 11390 6290 11470
rect 6550 11390 6630 11470
rect 6850 11390 6930 11470
rect 7170 11390 7250 11470
rect 7470 11390 7550 11470
rect 7810 11390 7890 11470
rect 8110 11390 8190 11470
rect 8430 11390 8510 11470
rect 8730 11390 8810 11470
rect 9070 11390 9150 11470
rect 9370 11390 9450 11470
rect 9690 11390 9770 11470
rect 9990 11390 10070 11470
rect 10330 11390 10410 11470
rect 10630 11390 10710 11470
rect 10950 11390 11030 11470
rect 11250 11390 11330 11470
rect 11660 11390 11740 11470
rect 11960 11390 12040 11470
rect 160 11210 240 11290
rect 870 11210 950 11290
rect 1170 11210 1250 11290
rect 1510 11210 1590 11290
rect 1810 11210 1890 11290
rect 2130 11210 2210 11290
rect 2430 11210 2510 11290
rect 2770 11210 2850 11290
rect 3070 11210 3150 11290
rect 3390 11210 3470 11290
rect 3690 11210 3770 11290
rect 4030 11210 4110 11290
rect 4330 11210 4410 11290
rect 4650 11210 4730 11290
rect 4950 11210 5030 11290
rect 5290 11210 5370 11290
rect 5590 11210 5670 11290
rect 5910 11210 5990 11290
rect 6210 11210 6290 11290
rect 6550 11210 6630 11290
rect 6850 11210 6930 11290
rect 7170 11210 7250 11290
rect 7470 11210 7550 11290
rect 7810 11210 7890 11290
rect 8110 11210 8190 11290
rect 8430 11210 8510 11290
rect 8730 11210 8810 11290
rect 9070 11210 9150 11290
rect 9370 11210 9450 11290
rect 9690 11210 9770 11290
rect 9990 11210 10070 11290
rect 10330 11210 10410 11290
rect 10630 11210 10710 11290
rect 10950 11210 11030 11290
rect 11250 11210 11330 11290
rect 11660 11210 11740 11290
rect 11960 11210 12040 11290
rect 160 11030 240 11110
rect 870 11030 950 11110
rect 1170 11030 1250 11110
rect 1510 11030 1590 11110
rect 1810 11030 1890 11110
rect 2130 11030 2210 11110
rect 2430 11030 2510 11110
rect 2770 11030 2850 11110
rect 3070 11030 3150 11110
rect 3390 11030 3470 11110
rect 3690 11030 3770 11110
rect 4030 11030 4110 11110
rect 4330 11030 4410 11110
rect 4650 11030 4730 11110
rect 4950 11030 5030 11110
rect 5290 11030 5370 11110
rect 5590 11030 5670 11110
rect 5910 11030 5990 11110
rect 6210 11030 6290 11110
rect 6550 11030 6630 11110
rect 6850 11030 6930 11110
rect 7170 11030 7250 11110
rect 7470 11030 7550 11110
rect 7810 11030 7890 11110
rect 8110 11030 8190 11110
rect 8430 11030 8510 11110
rect 8730 11030 8810 11110
rect 9070 11030 9150 11110
rect 9370 11030 9450 11110
rect 9690 11030 9770 11110
rect 9990 11030 10070 11110
rect 10330 11030 10410 11110
rect 10630 11030 10710 11110
rect 10950 11030 11030 11110
rect 11250 11030 11330 11110
rect 11660 11030 11740 11110
rect 11960 11030 12040 11110
rect 160 10850 240 10930
rect 870 10850 950 10930
rect 1170 10850 1250 10930
rect 1510 10850 1590 10930
rect 1810 10850 1890 10930
rect 2130 10850 2210 10930
rect 2430 10850 2510 10930
rect 2770 10850 2850 10930
rect 3070 10850 3150 10930
rect 3390 10850 3470 10930
rect 3690 10850 3770 10930
rect 4030 10850 4110 10930
rect 4330 10850 4410 10930
rect 4650 10850 4730 10930
rect 4950 10850 5030 10930
rect 5290 10850 5370 10930
rect 5590 10850 5670 10930
rect 5910 10850 5990 10930
rect 6210 10850 6290 10930
rect 6550 10850 6630 10930
rect 6850 10850 6930 10930
rect 7170 10850 7250 10930
rect 7470 10850 7550 10930
rect 7810 10850 7890 10930
rect 8110 10850 8190 10930
rect 8430 10850 8510 10930
rect 8730 10850 8810 10930
rect 9070 10850 9150 10930
rect 9370 10850 9450 10930
rect 9690 10850 9770 10930
rect 9990 10850 10070 10930
rect 10330 10850 10410 10930
rect 10630 10850 10710 10930
rect 10950 10850 11030 10930
rect 11250 10850 11330 10930
rect 11660 10850 11740 10930
rect 11960 10850 12040 10930
rect 160 10670 240 10750
rect 870 10670 950 10750
rect 1170 10670 1250 10750
rect 1510 10670 1590 10750
rect 1810 10670 1890 10750
rect 2130 10670 2210 10750
rect 2430 10670 2510 10750
rect 2770 10670 2850 10750
rect 3070 10670 3150 10750
rect 3390 10670 3470 10750
rect 3690 10670 3770 10750
rect 4030 10670 4110 10750
rect 4330 10670 4410 10750
rect 4650 10670 4730 10750
rect 4950 10670 5030 10750
rect 5290 10670 5370 10750
rect 5590 10670 5670 10750
rect 5910 10670 5990 10750
rect 6210 10670 6290 10750
rect 6550 10670 6630 10750
rect 6850 10670 6930 10750
rect 7170 10670 7250 10750
rect 7470 10670 7550 10750
rect 7810 10670 7890 10750
rect 8110 10670 8190 10750
rect 8430 10670 8510 10750
rect 8730 10670 8810 10750
rect 9070 10670 9150 10750
rect 9370 10670 9450 10750
rect 9690 10670 9770 10750
rect 9990 10670 10070 10750
rect 10330 10670 10410 10750
rect 10630 10670 10710 10750
rect 10950 10670 11030 10750
rect 11250 10670 11330 10750
rect 11660 10670 11740 10750
rect 11960 10670 12040 10750
rect 160 10490 240 10570
rect 870 10490 950 10570
rect 1170 10490 1250 10570
rect 1510 10490 1590 10570
rect 1810 10490 1890 10570
rect 2130 10490 2210 10570
rect 2430 10490 2510 10570
rect 2770 10490 2850 10570
rect 3070 10490 3150 10570
rect 3390 10490 3470 10570
rect 3690 10490 3770 10570
rect 4030 10490 4110 10570
rect 4330 10490 4410 10570
rect 4650 10490 4730 10570
rect 4950 10490 5030 10570
rect 5290 10490 5370 10570
rect 5590 10490 5670 10570
rect 5910 10490 5990 10570
rect 6210 10490 6290 10570
rect 6550 10490 6630 10570
rect 6850 10490 6930 10570
rect 7170 10490 7250 10570
rect 7470 10490 7550 10570
rect 7810 10490 7890 10570
rect 8110 10490 8190 10570
rect 8430 10490 8510 10570
rect 8730 10490 8810 10570
rect 9070 10490 9150 10570
rect 9370 10490 9450 10570
rect 9690 10490 9770 10570
rect 9990 10490 10070 10570
rect 10330 10490 10410 10570
rect 10630 10490 10710 10570
rect 10950 10490 11030 10570
rect 11250 10490 11330 10570
rect 11660 10490 11740 10570
rect 11960 10490 12040 10570
rect 160 10310 240 10390
rect 870 10310 950 10390
rect 1170 10310 1250 10390
rect 1510 10310 1590 10390
rect 1810 10310 1890 10390
rect 2130 10310 2210 10390
rect 2430 10310 2510 10390
rect 2770 10310 2850 10390
rect 3070 10310 3150 10390
rect 3390 10310 3470 10390
rect 3690 10310 3770 10390
rect 4030 10310 4110 10390
rect 4330 10310 4410 10390
rect 4650 10310 4730 10390
rect 4950 10310 5030 10390
rect 5290 10310 5370 10390
rect 5590 10310 5670 10390
rect 5910 10310 5990 10390
rect 6210 10310 6290 10390
rect 6550 10310 6630 10390
rect 6850 10310 6930 10390
rect 7170 10310 7250 10390
rect 7470 10310 7550 10390
rect 7810 10310 7890 10390
rect 8110 10310 8190 10390
rect 8430 10310 8510 10390
rect 8730 10310 8810 10390
rect 9070 10310 9150 10390
rect 9370 10310 9450 10390
rect 9690 10310 9770 10390
rect 9990 10310 10070 10390
rect 10330 10310 10410 10390
rect 10630 10310 10710 10390
rect 10950 10310 11030 10390
rect 11250 10310 11330 10390
rect 11660 10310 11740 10390
rect 11960 10310 12040 10390
rect 160 10130 240 10210
rect 870 10130 950 10210
rect 1170 10130 1250 10210
rect 1510 10130 1590 10210
rect 1810 10130 1890 10210
rect 2130 10130 2210 10210
rect 2430 10130 2510 10210
rect 2770 10130 2850 10210
rect 3070 10130 3150 10210
rect 3390 10130 3470 10210
rect 3690 10130 3770 10210
rect 4030 10130 4110 10210
rect 4330 10130 4410 10210
rect 4650 10130 4730 10210
rect 4950 10130 5030 10210
rect 5290 10130 5370 10210
rect 5590 10130 5670 10210
rect 5910 10130 5990 10210
rect 6210 10130 6290 10210
rect 6550 10130 6630 10210
rect 6850 10130 6930 10210
rect 7170 10130 7250 10210
rect 7470 10130 7550 10210
rect 7810 10130 7890 10210
rect 8110 10130 8190 10210
rect 8430 10130 8510 10210
rect 8730 10130 8810 10210
rect 9070 10130 9150 10210
rect 9370 10130 9450 10210
rect 9690 10130 9770 10210
rect 9990 10130 10070 10210
rect 10330 10130 10410 10210
rect 10630 10130 10710 10210
rect 10950 10130 11030 10210
rect 11250 10130 11330 10210
rect 11660 10130 11740 10210
rect 11960 10130 12040 10210
rect 160 9950 240 10030
rect 11660 9950 11740 10030
rect 11960 9950 12040 10030
rect 160 9770 240 9850
rect 11660 9770 11740 9850
rect 11960 9770 12040 9850
rect 160 9590 240 9670
rect 11660 9590 11740 9670
rect 11960 9590 12040 9670
rect 160 9410 240 9490
rect 11660 9410 11740 9490
rect 11960 9410 12040 9490
rect 160 9230 240 9310
rect 11660 9230 11740 9310
rect 11960 9230 12040 9310
<< m3contact >>
rect 2460 7810 2540 7890
rect 2860 7810 2940 7890
rect 3260 7810 3340 7890
rect 3660 7810 3740 7890
rect 4060 7810 4140 7890
rect 4460 7810 4540 7890
rect 4860 7810 4940 7890
rect 5260 7810 5340 7890
rect 5660 7810 5740 7890
rect 6060 7810 6140 7890
rect 6460 7810 6540 7890
rect 6860 7810 6940 7890
rect 7260 7810 7340 7890
rect 7660 7810 7740 7890
rect 8060 7810 8140 7890
rect 8460 7810 8540 7890
rect 8860 7810 8940 7890
rect 9260 7810 9340 7890
rect 9660 7810 9740 7890
rect 2460 7410 2540 7490
rect 2860 7410 2940 7490
rect 3260 7410 3340 7490
rect 3660 7410 3740 7490
rect 4060 7410 4140 7490
rect 4460 7410 4540 7490
rect 4860 7410 4940 7490
rect 5260 7410 5340 7490
rect 5660 7410 5740 7490
rect 6060 7410 6140 7490
rect 6460 7410 6540 7490
rect 6860 7410 6940 7490
rect 7260 7410 7340 7490
rect 7660 7410 7740 7490
rect 8060 7410 8140 7490
rect 8460 7410 8540 7490
rect 8860 7410 8940 7490
rect 9260 7410 9340 7490
rect 9660 7410 9740 7490
rect 2460 7010 2540 7090
rect 2860 7010 2940 7090
rect 3260 7010 3340 7090
rect 3660 7010 3740 7090
rect 4060 7010 4140 7090
rect 4460 7010 4540 7090
rect 4860 7010 4940 7090
rect 5260 7010 5340 7090
rect 5660 7010 5740 7090
rect 6060 7010 6140 7090
rect 6460 7010 6540 7090
rect 6860 7010 6940 7090
rect 7260 7010 7340 7090
rect 7660 7010 7740 7090
rect 8060 7010 8140 7090
rect 8460 7010 8540 7090
rect 8860 7010 8940 7090
rect 9260 7010 9340 7090
rect 9660 7010 9740 7090
rect 2460 6610 2540 6690
rect 2860 6610 2940 6690
rect 3260 6610 3340 6690
rect 3660 6610 3740 6690
rect 4060 6610 4140 6690
rect 4460 6610 4540 6690
rect 4860 6610 4940 6690
rect 5260 6610 5340 6690
rect 5660 6610 5740 6690
rect 6060 6610 6140 6690
rect 6460 6610 6540 6690
rect 6860 6610 6940 6690
rect 7260 6610 7340 6690
rect 7660 6610 7740 6690
rect 8060 6610 8140 6690
rect 8460 6610 8540 6690
rect 8860 6610 8940 6690
rect 9260 6610 9340 6690
rect 9660 6610 9740 6690
rect 2460 6210 2540 6290
rect 2860 6210 2940 6290
rect 3260 6210 3340 6290
rect 3660 6210 3740 6290
rect 4060 6210 4140 6290
rect 4460 6210 4540 6290
rect 4860 6210 4940 6290
rect 5260 6210 5340 6290
rect 5660 6210 5740 6290
rect 6060 6210 6140 6290
rect 6460 6210 6540 6290
rect 6860 6210 6940 6290
rect 7260 6210 7340 6290
rect 7660 6210 7740 6290
rect 8060 6210 8140 6290
rect 8460 6210 8540 6290
rect 8860 6210 8940 6290
rect 9260 6210 9340 6290
rect 9660 6210 9740 6290
rect 2460 5810 2540 5890
rect 2860 5810 2940 5890
rect 3260 5810 3340 5890
rect 3660 5810 3740 5890
rect 4060 5810 4140 5890
rect 4460 5810 4540 5890
rect 4860 5810 4940 5890
rect 5260 5810 5340 5890
rect 5660 5810 5740 5890
rect 6060 5810 6140 5890
rect 6460 5810 6540 5890
rect 6860 5810 6940 5890
rect 7260 5810 7340 5890
rect 7660 5810 7740 5890
rect 8060 5810 8140 5890
rect 8460 5810 8540 5890
rect 8860 5810 8940 5890
rect 9260 5810 9340 5890
rect 9660 5810 9740 5890
rect 2460 5410 2540 5490
rect 2860 5410 2940 5490
rect 3260 5410 3340 5490
rect 3660 5410 3740 5490
rect 4060 5410 4140 5490
rect 4460 5410 4540 5490
rect 4860 5410 4940 5490
rect 5260 5410 5340 5490
rect 5660 5410 5740 5490
rect 6060 5410 6140 5490
rect 6460 5410 6540 5490
rect 6860 5410 6940 5490
rect 7260 5410 7340 5490
rect 7660 5410 7740 5490
rect 8060 5410 8140 5490
rect 8460 5410 8540 5490
rect 8860 5410 8940 5490
rect 9260 5410 9340 5490
rect 9660 5410 9740 5490
rect 2460 5010 2540 5090
rect 2860 5010 2940 5090
rect 3260 5010 3340 5090
rect 3660 5010 3740 5090
rect 4060 5010 4140 5090
rect 4460 5010 4540 5090
rect 4860 5010 4940 5090
rect 5260 5010 5340 5090
rect 5660 5010 5740 5090
rect 6060 5010 6140 5090
rect 6460 5010 6540 5090
rect 6860 5010 6940 5090
rect 7260 5010 7340 5090
rect 7660 5010 7740 5090
rect 8060 5010 8140 5090
rect 8460 5010 8540 5090
rect 8860 5010 8940 5090
rect 9260 5010 9340 5090
rect 9660 5010 9740 5090
rect 2460 4610 2540 4690
rect 2860 4610 2940 4690
rect 3260 4610 3340 4690
rect 3660 4610 3740 4690
rect 4060 4610 4140 4690
rect 4460 4610 4540 4690
rect 4860 4610 4940 4690
rect 5260 4610 5340 4690
rect 5660 4610 5740 4690
rect 6060 4610 6140 4690
rect 6460 4610 6540 4690
rect 6860 4610 6940 4690
rect 7260 4610 7340 4690
rect 7660 4610 7740 4690
rect 8060 4610 8140 4690
rect 8460 4610 8540 4690
rect 8860 4610 8940 4690
rect 9260 4610 9340 4690
rect 9660 4610 9740 4690
rect 2460 4210 2540 4290
rect 2860 4210 2940 4290
rect 3260 4210 3340 4290
rect 3660 4210 3740 4290
rect 4060 4210 4140 4290
rect 4460 4210 4540 4290
rect 4860 4210 4940 4290
rect 5260 4210 5340 4290
rect 5660 4210 5740 4290
rect 6060 4210 6140 4290
rect 6460 4210 6540 4290
rect 6860 4210 6940 4290
rect 7260 4210 7340 4290
rect 7660 4210 7740 4290
rect 8060 4210 8140 4290
rect 8460 4210 8540 4290
rect 8860 4210 8940 4290
rect 9260 4210 9340 4290
rect 9660 4210 9740 4290
rect 2460 3810 2540 3890
rect 2860 3810 2940 3890
rect 3260 3810 3340 3890
rect 3660 3810 3740 3890
rect 4060 3810 4140 3890
rect 4460 3810 4540 3890
rect 4860 3810 4940 3890
rect 5260 3810 5340 3890
rect 5660 3810 5740 3890
rect 6060 3810 6140 3890
rect 6460 3810 6540 3890
rect 6860 3810 6940 3890
rect 7260 3810 7340 3890
rect 7660 3810 7740 3890
rect 8060 3810 8140 3890
rect 8460 3810 8540 3890
rect 8860 3810 8940 3890
rect 9260 3810 9340 3890
rect 9660 3810 9740 3890
rect 2460 3410 2540 3490
rect 2860 3410 2940 3490
rect 3260 3410 3340 3490
rect 3660 3410 3740 3490
rect 4060 3410 4140 3490
rect 4460 3410 4540 3490
rect 4860 3410 4940 3490
rect 5260 3410 5340 3490
rect 5660 3410 5740 3490
rect 6060 3410 6140 3490
rect 6460 3410 6540 3490
rect 6860 3410 6940 3490
rect 7260 3410 7340 3490
rect 7660 3410 7740 3490
rect 8060 3410 8140 3490
rect 8460 3410 8540 3490
rect 8860 3410 8940 3490
rect 9260 3410 9340 3490
rect 9660 3410 9740 3490
rect 2460 3010 2540 3090
rect 2860 3010 2940 3090
rect 3260 3010 3340 3090
rect 3660 3010 3740 3090
rect 4060 3010 4140 3090
rect 4460 3010 4540 3090
rect 4860 3010 4940 3090
rect 5260 3010 5340 3090
rect 5660 3010 5740 3090
rect 6060 3010 6140 3090
rect 6460 3010 6540 3090
rect 6860 3010 6940 3090
rect 7260 3010 7340 3090
rect 7660 3010 7740 3090
rect 8060 3010 8140 3090
rect 8460 3010 8540 3090
rect 8860 3010 8940 3090
rect 9260 3010 9340 3090
rect 9660 3010 9740 3090
rect 2460 2610 2540 2690
rect 2860 2610 2940 2690
rect 3260 2610 3340 2690
rect 3660 2610 3740 2690
rect 4060 2610 4140 2690
rect 4460 2610 4540 2690
rect 4860 2610 4940 2690
rect 5260 2610 5340 2690
rect 5660 2610 5740 2690
rect 6060 2610 6140 2690
rect 6460 2610 6540 2690
rect 6860 2610 6940 2690
rect 7260 2610 7340 2690
rect 7660 2610 7740 2690
rect 8060 2610 8140 2690
rect 8460 2610 8540 2690
rect 8860 2610 8940 2690
rect 9260 2610 9340 2690
rect 9660 2610 9740 2690
rect 2460 2210 2540 2290
rect 2860 2210 2940 2290
rect 3260 2210 3340 2290
rect 3660 2210 3740 2290
rect 4060 2210 4140 2290
rect 4460 2210 4540 2290
rect 4860 2210 4940 2290
rect 5260 2210 5340 2290
rect 5660 2210 5740 2290
rect 6060 2210 6140 2290
rect 6460 2210 6540 2290
rect 6860 2210 6940 2290
rect 7260 2210 7340 2290
rect 7660 2210 7740 2290
rect 8060 2210 8140 2290
rect 8460 2210 8540 2290
rect 8860 2210 8940 2290
rect 9260 2210 9340 2290
rect 9660 2210 9740 2290
rect 2460 1810 2540 1890
rect 2860 1810 2940 1890
rect 3260 1810 3340 1890
rect 3660 1810 3740 1890
rect 4060 1810 4140 1890
rect 4460 1810 4540 1890
rect 4860 1810 4940 1890
rect 5260 1810 5340 1890
rect 5660 1810 5740 1890
rect 6060 1810 6140 1890
rect 6460 1810 6540 1890
rect 6860 1810 6940 1890
rect 7260 1810 7340 1890
rect 7660 1810 7740 1890
rect 8060 1810 8140 1890
rect 8460 1810 8540 1890
rect 8860 1810 8940 1890
rect 9260 1810 9340 1890
rect 9660 1810 9740 1890
rect 2460 1410 2540 1490
rect 2860 1410 2940 1490
rect 3260 1410 3340 1490
rect 3660 1410 3740 1490
rect 4060 1410 4140 1490
rect 4460 1410 4540 1490
rect 4860 1410 4940 1490
rect 5260 1410 5340 1490
rect 5660 1410 5740 1490
rect 6060 1410 6140 1490
rect 6460 1410 6540 1490
rect 6860 1410 6940 1490
rect 7260 1410 7340 1490
rect 7660 1410 7740 1490
rect 8060 1410 8140 1490
rect 8460 1410 8540 1490
rect 8860 1410 8940 1490
rect 9260 1410 9340 1490
rect 9660 1410 9740 1490
rect 2460 1010 2540 1090
rect 2860 1010 2940 1090
rect 3260 1010 3340 1090
rect 3660 1010 3740 1090
rect 4060 1010 4140 1090
rect 4460 1010 4540 1090
rect 4860 1010 4940 1090
rect 5260 1010 5340 1090
rect 5660 1010 5740 1090
rect 6060 1010 6140 1090
rect 6460 1010 6540 1090
rect 6860 1010 6940 1090
rect 7260 1010 7340 1090
rect 7660 1010 7740 1090
rect 8060 1010 8140 1090
rect 8460 1010 8540 1090
rect 8860 1010 8940 1090
rect 9260 1010 9340 1090
rect 9660 1010 9740 1090
rect 2460 610 2540 690
rect 2860 610 2940 690
rect 3260 610 3340 690
rect 3660 610 3740 690
rect 4060 610 4140 690
rect 4460 610 4540 690
rect 4860 610 4940 690
rect 5260 610 5340 690
rect 5660 610 5740 690
rect 6060 610 6140 690
rect 6460 610 6540 690
rect 6860 610 6940 690
rect 7260 610 7340 690
rect 7660 610 7740 690
rect 8060 610 8140 690
rect 8460 610 8540 690
rect 8860 610 8940 690
rect 9260 610 9340 690
rect 9660 610 9740 690
<< metal3 >>
rect 100 32550 12100 34210
rect 100 30250 12100 31910
rect 100 20450 12100 28250
rect 100 9150 12100 16950
rect 1850 8250 10350 8500
rect 1850 250 2100 8250
rect 10100 250 10350 8250
rect 1850 0 10350 250
<< gv2 >>
rect 160 33870 240 33950
rect 11960 33870 12040 33950
rect 160 33590 240 33670
rect 11960 33590 12040 33670
rect 9140 33460 9220 33540
rect 10020 33460 10100 33540
rect 10610 33460 10690 33540
rect 11200 33460 11280 33540
rect 160 33310 240 33390
rect 11960 33310 12040 33390
rect 9140 33180 9220 33260
rect 10020 33180 10100 33260
rect 10610 33180 10690 33260
rect 11200 33180 11280 33260
rect 160 33030 240 33110
rect 11960 33030 12040 33110
rect 7625 32845 7705 32925
rect 7785 32845 7865 32925
rect 160 32750 240 32830
rect 11960 32750 12040 32830
rect 160 31570 240 31650
rect 11960 31570 12040 31650
rect 160 31290 240 31370
rect 11960 31290 12040 31370
rect 9140 31200 9220 31280
rect 10020 31200 10100 31280
rect 10620 31200 10700 31280
rect 11220 31200 11300 31280
rect 160 31010 240 31090
rect 11960 31010 12040 31090
rect 9140 30920 9220 31000
rect 10020 30920 10100 31000
rect 10620 30920 10700 31000
rect 11220 30920 11300 31000
rect 160 30730 240 30810
rect 11960 30730 12040 30810
rect 160 30450 240 30530
rect 11960 30450 12040 30530
rect 310 28090 390 28170
rect 11810 28090 11890 28170
rect 310 27910 390 27990
rect 11810 27910 11890 27990
rect 310 27730 390 27810
rect 11810 27730 11890 27810
rect 310 27550 390 27630
rect 11810 27550 11890 27630
rect 310 27370 390 27450
rect 11810 27370 11890 27450
rect 310 27190 390 27270
rect 1020 27190 1100 27270
rect 2280 27190 2360 27270
rect 3540 27190 3620 27270
rect 4800 27190 4880 27270
rect 6060 27190 6140 27270
rect 7320 27190 7400 27270
rect 8580 27190 8660 27270
rect 9840 27190 9920 27270
rect 11100 27190 11180 27270
rect 11810 27190 11890 27270
rect 310 27010 390 27090
rect 1020 27010 1100 27090
rect 2280 27010 2360 27090
rect 3540 27010 3620 27090
rect 4800 27010 4880 27090
rect 6060 27010 6140 27090
rect 7320 27010 7400 27090
rect 8580 27010 8660 27090
rect 9840 27010 9920 27090
rect 11100 27010 11180 27090
rect 11810 27010 11890 27090
rect 310 26830 390 26910
rect 1020 26830 1100 26910
rect 2280 26830 2360 26910
rect 3540 26830 3620 26910
rect 4800 26830 4880 26910
rect 6060 26830 6140 26910
rect 7320 26830 7400 26910
rect 8580 26830 8660 26910
rect 9840 26830 9920 26910
rect 11100 26830 11180 26910
rect 11810 26830 11890 26910
rect 310 26650 390 26730
rect 1020 26650 1100 26730
rect 2280 26650 2360 26730
rect 3540 26650 3620 26730
rect 4800 26650 4880 26730
rect 6060 26650 6140 26730
rect 7320 26650 7400 26730
rect 8580 26650 8660 26730
rect 9840 26650 9920 26730
rect 11100 26650 11180 26730
rect 11810 26650 11890 26730
rect 310 26470 390 26550
rect 1020 26470 1100 26550
rect 2280 26470 2360 26550
rect 3540 26470 3620 26550
rect 4800 26470 4880 26550
rect 6060 26470 6140 26550
rect 7320 26470 7400 26550
rect 8580 26470 8660 26550
rect 9840 26470 9920 26550
rect 11100 26470 11180 26550
rect 11810 26470 11890 26550
rect 310 26290 390 26370
rect 1020 26290 1100 26370
rect 2280 26290 2360 26370
rect 3540 26290 3620 26370
rect 4800 26290 4880 26370
rect 6060 26290 6140 26370
rect 7320 26290 7400 26370
rect 8580 26290 8660 26370
rect 9840 26290 9920 26370
rect 11100 26290 11180 26370
rect 11810 26290 11890 26370
rect 310 26110 390 26190
rect 1020 26110 1100 26190
rect 2280 26110 2360 26190
rect 3540 26110 3620 26190
rect 4800 26110 4880 26190
rect 6060 26110 6140 26190
rect 7320 26110 7400 26190
rect 8580 26110 8660 26190
rect 9840 26110 9920 26190
rect 11100 26110 11180 26190
rect 11810 26110 11890 26190
rect 310 25930 390 26010
rect 1020 25930 1100 26010
rect 2280 25930 2360 26010
rect 3540 25930 3620 26010
rect 4800 25930 4880 26010
rect 6060 25930 6140 26010
rect 7320 25930 7400 26010
rect 8580 25930 8660 26010
rect 9840 25930 9920 26010
rect 11100 25930 11180 26010
rect 11810 25930 11890 26010
rect 310 25750 390 25830
rect 1020 25750 1100 25830
rect 2280 25750 2360 25830
rect 3540 25750 3620 25830
rect 4800 25750 4880 25830
rect 6060 25750 6140 25830
rect 7320 25750 7400 25830
rect 8580 25750 8660 25830
rect 9840 25750 9920 25830
rect 11100 25750 11180 25830
rect 11810 25750 11890 25830
rect 310 25570 390 25650
rect 1020 25570 1100 25650
rect 2280 25570 2360 25650
rect 3540 25570 3620 25650
rect 4800 25570 4880 25650
rect 6060 25570 6140 25650
rect 7320 25570 7400 25650
rect 8580 25570 8660 25650
rect 9840 25570 9920 25650
rect 11100 25570 11180 25650
rect 11810 25570 11890 25650
rect 310 25390 390 25470
rect 1020 25390 1100 25470
rect 2280 25390 2360 25470
rect 3540 25390 3620 25470
rect 4800 25390 4880 25470
rect 6060 25390 6140 25470
rect 7320 25390 7400 25470
rect 8580 25390 8660 25470
rect 9840 25390 9920 25470
rect 11100 25390 11180 25470
rect 11810 25390 11890 25470
rect 310 25210 390 25290
rect 1020 25210 1100 25290
rect 2280 25210 2360 25290
rect 3540 25210 3620 25290
rect 4800 25210 4880 25290
rect 6060 25210 6140 25290
rect 7320 25210 7400 25290
rect 8580 25210 8660 25290
rect 9840 25210 9920 25290
rect 11100 25210 11180 25290
rect 11810 25210 11890 25290
rect 310 25030 390 25110
rect 1020 25030 1100 25110
rect 2280 25030 2360 25110
rect 3540 25030 3620 25110
rect 4800 25030 4880 25110
rect 6060 25030 6140 25110
rect 7320 25030 7400 25110
rect 8580 25030 8660 25110
rect 9840 25030 9920 25110
rect 11100 25030 11180 25110
rect 11810 25030 11890 25110
rect 310 24850 390 24930
rect 1020 24850 1100 24930
rect 2280 24850 2360 24930
rect 3540 24850 3620 24930
rect 4800 24850 4880 24930
rect 6060 24850 6140 24930
rect 7320 24850 7400 24930
rect 8580 24850 8660 24930
rect 9840 24850 9920 24930
rect 11100 24850 11180 24930
rect 11810 24850 11890 24930
rect 310 24670 390 24750
rect 1020 24670 1100 24750
rect 2280 24670 2360 24750
rect 3540 24670 3620 24750
rect 4800 24670 4880 24750
rect 6060 24670 6140 24750
rect 7320 24670 7400 24750
rect 8580 24670 8660 24750
rect 9840 24670 9920 24750
rect 11100 24670 11180 24750
rect 11810 24670 11890 24750
rect 310 24490 390 24570
rect 1020 24490 1100 24570
rect 2280 24490 2360 24570
rect 3540 24490 3620 24570
rect 4800 24490 4880 24570
rect 6060 24490 6140 24570
rect 7320 24490 7400 24570
rect 8580 24490 8660 24570
rect 9840 24490 9920 24570
rect 11100 24490 11180 24570
rect 11810 24490 11890 24570
rect 310 24310 390 24390
rect 1020 24310 1100 24390
rect 2280 24310 2360 24390
rect 3540 24310 3620 24390
rect 4800 24310 4880 24390
rect 6060 24310 6140 24390
rect 7320 24310 7400 24390
rect 8580 24310 8660 24390
rect 9840 24310 9920 24390
rect 11100 24310 11180 24390
rect 11810 24310 11890 24390
rect 310 24130 390 24210
rect 1020 24130 1100 24210
rect 2280 24130 2360 24210
rect 3540 24130 3620 24210
rect 4800 24130 4880 24210
rect 6060 24130 6140 24210
rect 7320 24130 7400 24210
rect 8580 24130 8660 24210
rect 9840 24130 9920 24210
rect 11100 24130 11180 24210
rect 11810 24130 11890 24210
rect 310 23950 390 24030
rect 1020 23950 1100 24030
rect 2280 23950 2360 24030
rect 3540 23950 3620 24030
rect 4800 23950 4880 24030
rect 6060 23950 6140 24030
rect 7320 23950 7400 24030
rect 8580 23950 8660 24030
rect 9840 23950 9920 24030
rect 11100 23950 11180 24030
rect 11810 23950 11890 24030
rect 310 23770 390 23850
rect 1020 23770 1100 23850
rect 2280 23770 2360 23850
rect 3540 23770 3620 23850
rect 4800 23770 4880 23850
rect 6060 23770 6140 23850
rect 7320 23770 7400 23850
rect 8580 23770 8660 23850
rect 9840 23770 9920 23850
rect 11100 23770 11180 23850
rect 11810 23770 11890 23850
rect 310 23590 390 23670
rect 1020 23590 1100 23670
rect 2280 23590 2360 23670
rect 3540 23590 3620 23670
rect 4800 23590 4880 23670
rect 6060 23590 6140 23670
rect 7320 23590 7400 23670
rect 8580 23590 8660 23670
rect 9840 23590 9920 23670
rect 11100 23590 11180 23670
rect 11810 23590 11890 23670
rect 310 23410 390 23490
rect 1020 23410 1100 23490
rect 2280 23410 2360 23490
rect 3540 23410 3620 23490
rect 4800 23410 4880 23490
rect 6060 23410 6140 23490
rect 7320 23410 7400 23490
rect 8580 23410 8660 23490
rect 9840 23410 9920 23490
rect 11100 23410 11180 23490
rect 11810 23410 11890 23490
rect 310 23230 390 23310
rect 1020 23230 1100 23310
rect 2280 23230 2360 23310
rect 3540 23230 3620 23310
rect 4800 23230 4880 23310
rect 6060 23230 6140 23310
rect 7320 23230 7400 23310
rect 8580 23230 8660 23310
rect 9840 23230 9920 23310
rect 11100 23230 11180 23310
rect 11810 23230 11890 23310
rect 310 23050 390 23130
rect 1020 23050 1100 23130
rect 2280 23050 2360 23130
rect 3540 23050 3620 23130
rect 4800 23050 4880 23130
rect 6060 23050 6140 23130
rect 7320 23050 7400 23130
rect 8580 23050 8660 23130
rect 9840 23050 9920 23130
rect 11100 23050 11180 23130
rect 11810 23050 11890 23130
rect 310 22870 390 22950
rect 1020 22870 1100 22950
rect 2280 22870 2360 22950
rect 3540 22870 3620 22950
rect 4800 22870 4880 22950
rect 6060 22870 6140 22950
rect 7320 22870 7400 22950
rect 8580 22870 8660 22950
rect 9840 22870 9920 22950
rect 11100 22870 11180 22950
rect 11810 22870 11890 22950
rect 310 22690 390 22770
rect 1020 22690 1100 22770
rect 2280 22690 2360 22770
rect 3540 22690 3620 22770
rect 4800 22690 4880 22770
rect 6060 22690 6140 22770
rect 7320 22690 7400 22770
rect 8580 22690 8660 22770
rect 9840 22690 9920 22770
rect 11100 22690 11180 22770
rect 11810 22690 11890 22770
rect 310 22510 390 22590
rect 1020 22510 1100 22590
rect 2280 22510 2360 22590
rect 3540 22510 3620 22590
rect 4800 22510 4880 22590
rect 6060 22510 6140 22590
rect 7320 22510 7400 22590
rect 8580 22510 8660 22590
rect 9840 22510 9920 22590
rect 11100 22510 11180 22590
rect 11810 22510 11890 22590
rect 310 22330 390 22410
rect 1020 22330 1100 22410
rect 2280 22330 2360 22410
rect 3540 22330 3620 22410
rect 4800 22330 4880 22410
rect 6060 22330 6140 22410
rect 7320 22330 7400 22410
rect 8580 22330 8660 22410
rect 9840 22330 9920 22410
rect 11100 22330 11180 22410
rect 11810 22330 11890 22410
rect 310 22150 390 22230
rect 1020 22150 1100 22230
rect 2280 22150 2360 22230
rect 3540 22150 3620 22230
rect 4800 22150 4880 22230
rect 6060 22150 6140 22230
rect 7320 22150 7400 22230
rect 8580 22150 8660 22230
rect 9840 22150 9920 22230
rect 11100 22150 11180 22230
rect 11810 22150 11890 22230
rect 310 21970 390 22050
rect 1020 21970 1100 22050
rect 2280 21970 2360 22050
rect 3540 21970 3620 22050
rect 4800 21970 4880 22050
rect 6060 21970 6140 22050
rect 7320 21970 7400 22050
rect 8580 21970 8660 22050
rect 9840 21970 9920 22050
rect 11100 21970 11180 22050
rect 11810 21970 11890 22050
rect 310 21790 390 21870
rect 1020 21790 1100 21870
rect 2280 21790 2360 21870
rect 3540 21790 3620 21870
rect 4800 21790 4880 21870
rect 6060 21790 6140 21870
rect 7320 21790 7400 21870
rect 8580 21790 8660 21870
rect 9840 21790 9920 21870
rect 11100 21790 11180 21870
rect 11810 21790 11890 21870
rect 310 21610 390 21690
rect 1020 21610 1100 21690
rect 2280 21610 2360 21690
rect 3540 21610 3620 21690
rect 4800 21610 4880 21690
rect 6060 21610 6140 21690
rect 7320 21610 7400 21690
rect 8580 21610 8660 21690
rect 9840 21610 9920 21690
rect 11100 21610 11180 21690
rect 11810 21610 11890 21690
rect 310 21430 390 21510
rect 1020 21430 1100 21510
rect 2280 21430 2360 21510
rect 3540 21430 3620 21510
rect 4800 21430 4880 21510
rect 6060 21430 6140 21510
rect 7320 21430 7400 21510
rect 8580 21430 8660 21510
rect 9840 21430 9920 21510
rect 11100 21430 11180 21510
rect 11810 21430 11890 21510
rect 310 21250 390 21330
rect 11810 21250 11890 21330
rect 310 21070 390 21150
rect 11810 21070 11890 21150
rect 310 20890 390 20970
rect 11810 20890 11890 20970
rect 310 20710 390 20790
rect 11810 20710 11890 20790
rect 310 20530 390 20610
rect 11810 20530 11890 20610
rect 310 16790 390 16870
rect 11810 16790 11890 16870
rect 310 16610 390 16690
rect 11810 16610 11890 16690
rect 310 16430 390 16510
rect 11810 16430 11890 16510
rect 310 16250 390 16330
rect 11810 16250 11890 16330
rect 310 16070 390 16150
rect 11810 16070 11890 16150
rect 310 15890 390 15970
rect 1020 15890 1100 15970
rect 2280 15890 2360 15970
rect 3540 15890 3620 15970
rect 4800 15890 4880 15970
rect 6060 15890 6140 15970
rect 7320 15890 7400 15970
rect 8580 15890 8660 15970
rect 9840 15890 9920 15970
rect 11100 15890 11180 15970
rect 11810 15890 11890 15970
rect 310 15710 390 15790
rect 1020 15710 1100 15790
rect 2280 15710 2360 15790
rect 3540 15710 3620 15790
rect 4800 15710 4880 15790
rect 6060 15710 6140 15790
rect 7320 15710 7400 15790
rect 8580 15710 8660 15790
rect 9840 15710 9920 15790
rect 11100 15710 11180 15790
rect 11810 15710 11890 15790
rect 310 15530 390 15610
rect 1020 15530 1100 15610
rect 2280 15530 2360 15610
rect 3540 15530 3620 15610
rect 4800 15530 4880 15610
rect 6060 15530 6140 15610
rect 7320 15530 7400 15610
rect 8580 15530 8660 15610
rect 9840 15530 9920 15610
rect 11100 15530 11180 15610
rect 11810 15530 11890 15610
rect 310 15350 390 15430
rect 1020 15350 1100 15430
rect 2280 15350 2360 15430
rect 3540 15350 3620 15430
rect 4800 15350 4880 15430
rect 6060 15350 6140 15430
rect 7320 15350 7400 15430
rect 8580 15350 8660 15430
rect 9840 15350 9920 15430
rect 11100 15350 11180 15430
rect 11810 15350 11890 15430
rect 310 15170 390 15250
rect 1020 15170 1100 15250
rect 2280 15170 2360 15250
rect 3540 15170 3620 15250
rect 4800 15170 4880 15250
rect 6060 15170 6140 15250
rect 7320 15170 7400 15250
rect 8580 15170 8660 15250
rect 9840 15170 9920 15250
rect 11100 15170 11180 15250
rect 11810 15170 11890 15250
rect 310 14990 390 15070
rect 1020 14990 1100 15070
rect 2280 14990 2360 15070
rect 3540 14990 3620 15070
rect 4800 14990 4880 15070
rect 6060 14990 6140 15070
rect 7320 14990 7400 15070
rect 8580 14990 8660 15070
rect 9840 14990 9920 15070
rect 11100 14990 11180 15070
rect 11810 14990 11890 15070
rect 310 14810 390 14890
rect 1020 14810 1100 14890
rect 2280 14810 2360 14890
rect 3540 14810 3620 14890
rect 4800 14810 4880 14890
rect 6060 14810 6140 14890
rect 7320 14810 7400 14890
rect 8580 14810 8660 14890
rect 9840 14810 9920 14890
rect 11100 14810 11180 14890
rect 11810 14810 11890 14890
rect 310 14630 390 14710
rect 1020 14630 1100 14710
rect 2280 14630 2360 14710
rect 3540 14630 3620 14710
rect 4800 14630 4880 14710
rect 6060 14630 6140 14710
rect 7320 14630 7400 14710
rect 8580 14630 8660 14710
rect 9840 14630 9920 14710
rect 11100 14630 11180 14710
rect 11810 14630 11890 14710
rect 310 14450 390 14530
rect 1020 14450 1100 14530
rect 2280 14450 2360 14530
rect 3540 14450 3620 14530
rect 4800 14450 4880 14530
rect 6060 14450 6140 14530
rect 7320 14450 7400 14530
rect 8580 14450 8660 14530
rect 9840 14450 9920 14530
rect 11100 14450 11180 14530
rect 11810 14450 11890 14530
rect 310 14270 390 14350
rect 1020 14270 1100 14350
rect 2280 14270 2360 14350
rect 3540 14270 3620 14350
rect 4800 14270 4880 14350
rect 6060 14270 6140 14350
rect 7320 14270 7400 14350
rect 8580 14270 8660 14350
rect 9840 14270 9920 14350
rect 11100 14270 11180 14350
rect 11810 14270 11890 14350
rect 310 14090 390 14170
rect 1020 14090 1100 14170
rect 2280 14090 2360 14170
rect 3540 14090 3620 14170
rect 4800 14090 4880 14170
rect 6060 14090 6140 14170
rect 7320 14090 7400 14170
rect 8580 14090 8660 14170
rect 9840 14090 9920 14170
rect 11100 14090 11180 14170
rect 11810 14090 11890 14170
rect 310 13910 390 13990
rect 1020 13910 1100 13990
rect 2280 13910 2360 13990
rect 3540 13910 3620 13990
rect 4800 13910 4880 13990
rect 6060 13910 6140 13990
rect 7320 13910 7400 13990
rect 8580 13910 8660 13990
rect 9840 13910 9920 13990
rect 11100 13910 11180 13990
rect 11810 13910 11890 13990
rect 310 13730 390 13810
rect 1020 13730 1100 13810
rect 2280 13730 2360 13810
rect 3540 13730 3620 13810
rect 4800 13730 4880 13810
rect 6060 13730 6140 13810
rect 7320 13730 7400 13810
rect 8580 13730 8660 13810
rect 9840 13730 9920 13810
rect 11100 13730 11180 13810
rect 11810 13730 11890 13810
rect 310 13550 390 13630
rect 1020 13550 1100 13630
rect 2280 13550 2360 13630
rect 3540 13550 3620 13630
rect 4800 13550 4880 13630
rect 6060 13550 6140 13630
rect 7320 13550 7400 13630
rect 8580 13550 8660 13630
rect 9840 13550 9920 13630
rect 11100 13550 11180 13630
rect 11810 13550 11890 13630
rect 310 13370 390 13450
rect 1020 13370 1100 13450
rect 2280 13370 2360 13450
rect 3540 13370 3620 13450
rect 4800 13370 4880 13450
rect 6060 13370 6140 13450
rect 7320 13370 7400 13450
rect 8580 13370 8660 13450
rect 9840 13370 9920 13450
rect 11100 13370 11180 13450
rect 11810 13370 11890 13450
rect 310 13190 390 13270
rect 1020 13190 1100 13270
rect 2280 13190 2360 13270
rect 3540 13190 3620 13270
rect 4800 13190 4880 13270
rect 6060 13190 6140 13270
rect 7320 13190 7400 13270
rect 8580 13190 8660 13270
rect 9840 13190 9920 13270
rect 11100 13190 11180 13270
rect 11810 13190 11890 13270
rect 310 13010 390 13090
rect 1020 13010 1100 13090
rect 2280 13010 2360 13090
rect 3540 13010 3620 13090
rect 4800 13010 4880 13090
rect 6060 13010 6140 13090
rect 7320 13010 7400 13090
rect 8580 13010 8660 13090
rect 9840 13010 9920 13090
rect 11100 13010 11180 13090
rect 11810 13010 11890 13090
rect 310 12830 390 12910
rect 1020 12830 1100 12910
rect 2280 12830 2360 12910
rect 3540 12830 3620 12910
rect 4800 12830 4880 12910
rect 6060 12830 6140 12910
rect 7320 12830 7400 12910
rect 8580 12830 8660 12910
rect 9840 12830 9920 12910
rect 11100 12830 11180 12910
rect 11810 12830 11890 12910
rect 310 12650 390 12730
rect 1020 12650 1100 12730
rect 2280 12650 2360 12730
rect 3540 12650 3620 12730
rect 4800 12650 4880 12730
rect 6060 12650 6140 12730
rect 7320 12650 7400 12730
rect 8580 12650 8660 12730
rect 9840 12650 9920 12730
rect 11100 12650 11180 12730
rect 11810 12650 11890 12730
rect 310 12470 390 12550
rect 1020 12470 1100 12550
rect 2280 12470 2360 12550
rect 3540 12470 3620 12550
rect 4800 12470 4880 12550
rect 6060 12470 6140 12550
rect 7320 12470 7400 12550
rect 8580 12470 8660 12550
rect 9840 12470 9920 12550
rect 11100 12470 11180 12550
rect 11810 12470 11890 12550
rect 310 12290 390 12370
rect 1020 12290 1100 12370
rect 2280 12290 2360 12370
rect 3540 12290 3620 12370
rect 4800 12290 4880 12370
rect 6060 12290 6140 12370
rect 7320 12290 7400 12370
rect 8580 12290 8660 12370
rect 9840 12290 9920 12370
rect 11100 12290 11180 12370
rect 11810 12290 11890 12370
rect 310 12110 390 12190
rect 1020 12110 1100 12190
rect 2280 12110 2360 12190
rect 3540 12110 3620 12190
rect 4800 12110 4880 12190
rect 6060 12110 6140 12190
rect 7320 12110 7400 12190
rect 8580 12110 8660 12190
rect 9840 12110 9920 12190
rect 11100 12110 11180 12190
rect 11810 12110 11890 12190
rect 310 11930 390 12010
rect 1020 11930 1100 12010
rect 2280 11930 2360 12010
rect 3540 11930 3620 12010
rect 4800 11930 4880 12010
rect 6060 11930 6140 12010
rect 7320 11930 7400 12010
rect 8580 11930 8660 12010
rect 9840 11930 9920 12010
rect 11100 11930 11180 12010
rect 11810 11930 11890 12010
rect 310 11750 390 11830
rect 1020 11750 1100 11830
rect 2280 11750 2360 11830
rect 3540 11750 3620 11830
rect 4800 11750 4880 11830
rect 6060 11750 6140 11830
rect 7320 11750 7400 11830
rect 8580 11750 8660 11830
rect 9840 11750 9920 11830
rect 11100 11750 11180 11830
rect 11810 11750 11890 11830
rect 310 11570 390 11650
rect 1020 11570 1100 11650
rect 2280 11570 2360 11650
rect 3540 11570 3620 11650
rect 4800 11570 4880 11650
rect 6060 11570 6140 11650
rect 7320 11570 7400 11650
rect 8580 11570 8660 11650
rect 9840 11570 9920 11650
rect 11100 11570 11180 11650
rect 11810 11570 11890 11650
rect 310 11390 390 11470
rect 1020 11390 1100 11470
rect 2280 11390 2360 11470
rect 3540 11390 3620 11470
rect 4800 11390 4880 11470
rect 6060 11390 6140 11470
rect 7320 11390 7400 11470
rect 8580 11390 8660 11470
rect 9840 11390 9920 11470
rect 11100 11390 11180 11470
rect 11810 11390 11890 11470
rect 310 11210 390 11290
rect 1020 11210 1100 11290
rect 2280 11210 2360 11290
rect 3540 11210 3620 11290
rect 4800 11210 4880 11290
rect 6060 11210 6140 11290
rect 7320 11210 7400 11290
rect 8580 11210 8660 11290
rect 9840 11210 9920 11290
rect 11100 11210 11180 11290
rect 11810 11210 11890 11290
rect 310 11030 390 11110
rect 1020 11030 1100 11110
rect 2280 11030 2360 11110
rect 3540 11030 3620 11110
rect 4800 11030 4880 11110
rect 6060 11030 6140 11110
rect 7320 11030 7400 11110
rect 8580 11030 8660 11110
rect 9840 11030 9920 11110
rect 11100 11030 11180 11110
rect 11810 11030 11890 11110
rect 310 10850 390 10930
rect 1020 10850 1100 10930
rect 2280 10850 2360 10930
rect 3540 10850 3620 10930
rect 4800 10850 4880 10930
rect 6060 10850 6140 10930
rect 7320 10850 7400 10930
rect 8580 10850 8660 10930
rect 9840 10850 9920 10930
rect 11100 10850 11180 10930
rect 11810 10850 11890 10930
rect 310 10670 390 10750
rect 1020 10670 1100 10750
rect 2280 10670 2360 10750
rect 3540 10670 3620 10750
rect 4800 10670 4880 10750
rect 6060 10670 6140 10750
rect 7320 10670 7400 10750
rect 8580 10670 8660 10750
rect 9840 10670 9920 10750
rect 11100 10670 11180 10750
rect 11810 10670 11890 10750
rect 310 10490 390 10570
rect 1020 10490 1100 10570
rect 2280 10490 2360 10570
rect 3540 10490 3620 10570
rect 4800 10490 4880 10570
rect 6060 10490 6140 10570
rect 7320 10490 7400 10570
rect 8580 10490 8660 10570
rect 9840 10490 9920 10570
rect 11100 10490 11180 10570
rect 11810 10490 11890 10570
rect 310 10310 390 10390
rect 1020 10310 1100 10390
rect 2280 10310 2360 10390
rect 3540 10310 3620 10390
rect 4800 10310 4880 10390
rect 6060 10310 6140 10390
rect 7320 10310 7400 10390
rect 8580 10310 8660 10390
rect 9840 10310 9920 10390
rect 11100 10310 11180 10390
rect 11810 10310 11890 10390
rect 310 10130 390 10210
rect 1020 10130 1100 10210
rect 2280 10130 2360 10210
rect 3540 10130 3620 10210
rect 4800 10130 4880 10210
rect 6060 10130 6140 10210
rect 7320 10130 7400 10210
rect 8580 10130 8660 10210
rect 9840 10130 9920 10210
rect 11100 10130 11180 10210
rect 11810 10130 11890 10210
rect 310 9950 390 10030
rect 11810 9950 11890 10030
rect 310 9770 390 9850
rect 11810 9770 11890 9850
rect 310 9590 390 9670
rect 11810 9590 11890 9670
rect 310 9410 390 9490
rect 11810 9410 11890 9490
rect 310 9230 390 9310
rect 11810 9230 11890 9310
<< pad >>
rect 2100 7890 10100 8250
rect 2100 7810 2460 7890
rect 2540 7810 2860 7890
rect 2940 7810 3260 7890
rect 3340 7810 3660 7890
rect 3740 7810 4060 7890
rect 4140 7810 4460 7890
rect 4540 7810 4860 7890
rect 4940 7810 5260 7890
rect 5340 7810 5660 7890
rect 5740 7810 6060 7890
rect 6140 7810 6460 7890
rect 6540 7810 6860 7890
rect 6940 7810 7260 7890
rect 7340 7810 7660 7890
rect 7740 7810 8060 7890
rect 8140 7810 8460 7890
rect 8540 7810 8860 7890
rect 8940 7810 9260 7890
rect 9340 7810 9660 7890
rect 9740 7810 10100 7890
rect 2100 7490 10100 7810
rect 2100 7410 2460 7490
rect 2540 7410 2860 7490
rect 2940 7410 3260 7490
rect 3340 7410 3660 7490
rect 3740 7410 4060 7490
rect 4140 7410 4460 7490
rect 4540 7410 4860 7490
rect 4940 7410 5260 7490
rect 5340 7410 5660 7490
rect 5740 7410 6060 7490
rect 6140 7410 6460 7490
rect 6540 7410 6860 7490
rect 6940 7410 7260 7490
rect 7340 7410 7660 7490
rect 7740 7410 8060 7490
rect 8140 7410 8460 7490
rect 8540 7410 8860 7490
rect 8940 7410 9260 7490
rect 9340 7410 9660 7490
rect 9740 7410 10100 7490
rect 2100 7090 10100 7410
rect 2100 7010 2460 7090
rect 2540 7010 2860 7090
rect 2940 7010 3260 7090
rect 3340 7010 3660 7090
rect 3740 7010 4060 7090
rect 4140 7010 4460 7090
rect 4540 7010 4860 7090
rect 4940 7010 5260 7090
rect 5340 7010 5660 7090
rect 5740 7010 6060 7090
rect 6140 7010 6460 7090
rect 6540 7010 6860 7090
rect 6940 7010 7260 7090
rect 7340 7010 7660 7090
rect 7740 7010 8060 7090
rect 8140 7010 8460 7090
rect 8540 7010 8860 7090
rect 8940 7010 9260 7090
rect 9340 7010 9660 7090
rect 9740 7010 10100 7090
rect 2100 6690 10100 7010
rect 2100 6610 2460 6690
rect 2540 6610 2860 6690
rect 2940 6610 3260 6690
rect 3340 6610 3660 6690
rect 3740 6610 4060 6690
rect 4140 6610 4460 6690
rect 4540 6610 4860 6690
rect 4940 6610 5260 6690
rect 5340 6610 5660 6690
rect 5740 6610 6060 6690
rect 6140 6610 6460 6690
rect 6540 6610 6860 6690
rect 6940 6610 7260 6690
rect 7340 6610 7660 6690
rect 7740 6610 8060 6690
rect 8140 6610 8460 6690
rect 8540 6610 8860 6690
rect 8940 6610 9260 6690
rect 9340 6610 9660 6690
rect 9740 6610 10100 6690
rect 2100 6290 10100 6610
rect 2100 6210 2460 6290
rect 2540 6210 2860 6290
rect 2940 6210 3260 6290
rect 3340 6210 3660 6290
rect 3740 6210 4060 6290
rect 4140 6210 4460 6290
rect 4540 6210 4860 6290
rect 4940 6210 5260 6290
rect 5340 6210 5660 6290
rect 5740 6210 6060 6290
rect 6140 6210 6460 6290
rect 6540 6210 6860 6290
rect 6940 6210 7260 6290
rect 7340 6210 7660 6290
rect 7740 6210 8060 6290
rect 8140 6210 8460 6290
rect 8540 6210 8860 6290
rect 8940 6210 9260 6290
rect 9340 6210 9660 6290
rect 9740 6210 10100 6290
rect 2100 5890 10100 6210
rect 2100 5810 2460 5890
rect 2540 5810 2860 5890
rect 2940 5810 3260 5890
rect 3340 5810 3660 5890
rect 3740 5810 4060 5890
rect 4140 5810 4460 5890
rect 4540 5810 4860 5890
rect 4940 5810 5260 5890
rect 5340 5810 5660 5890
rect 5740 5810 6060 5890
rect 6140 5810 6460 5890
rect 6540 5810 6860 5890
rect 6940 5810 7260 5890
rect 7340 5810 7660 5890
rect 7740 5810 8060 5890
rect 8140 5810 8460 5890
rect 8540 5810 8860 5890
rect 8940 5810 9260 5890
rect 9340 5810 9660 5890
rect 9740 5810 10100 5890
rect 2100 5490 10100 5810
rect 2100 5410 2460 5490
rect 2540 5410 2860 5490
rect 2940 5410 3260 5490
rect 3340 5410 3660 5490
rect 3740 5410 4060 5490
rect 4140 5410 4460 5490
rect 4540 5410 4860 5490
rect 4940 5410 5260 5490
rect 5340 5410 5660 5490
rect 5740 5410 6060 5490
rect 6140 5410 6460 5490
rect 6540 5410 6860 5490
rect 6940 5410 7260 5490
rect 7340 5410 7660 5490
rect 7740 5410 8060 5490
rect 8140 5410 8460 5490
rect 8540 5410 8860 5490
rect 8940 5410 9260 5490
rect 9340 5410 9660 5490
rect 9740 5410 10100 5490
rect 2100 5090 10100 5410
rect 2100 5010 2460 5090
rect 2540 5010 2860 5090
rect 2940 5010 3260 5090
rect 3340 5010 3660 5090
rect 3740 5010 4060 5090
rect 4140 5010 4460 5090
rect 4540 5010 4860 5090
rect 4940 5010 5260 5090
rect 5340 5010 5660 5090
rect 5740 5010 6060 5090
rect 6140 5010 6460 5090
rect 6540 5010 6860 5090
rect 6940 5010 7260 5090
rect 7340 5010 7660 5090
rect 7740 5010 8060 5090
rect 8140 5010 8460 5090
rect 8540 5010 8860 5090
rect 8940 5010 9260 5090
rect 9340 5010 9660 5090
rect 9740 5010 10100 5090
rect 2100 4690 10100 5010
rect 2100 4610 2460 4690
rect 2540 4610 2860 4690
rect 2940 4610 3260 4690
rect 3340 4610 3660 4690
rect 3740 4610 4060 4690
rect 4140 4610 4460 4690
rect 4540 4610 4860 4690
rect 4940 4610 5260 4690
rect 5340 4610 5660 4690
rect 5740 4610 6060 4690
rect 6140 4610 6460 4690
rect 6540 4610 6860 4690
rect 6940 4610 7260 4690
rect 7340 4610 7660 4690
rect 7740 4610 8060 4690
rect 8140 4610 8460 4690
rect 8540 4610 8860 4690
rect 8940 4610 9260 4690
rect 9340 4610 9660 4690
rect 9740 4610 10100 4690
rect 2100 4290 10100 4610
rect 2100 4210 2460 4290
rect 2540 4210 2860 4290
rect 2940 4210 3260 4290
rect 3340 4210 3660 4290
rect 3740 4210 4060 4290
rect 4140 4210 4460 4290
rect 4540 4210 4860 4290
rect 4940 4210 5260 4290
rect 5340 4210 5660 4290
rect 5740 4210 6060 4290
rect 6140 4210 6460 4290
rect 6540 4210 6860 4290
rect 6940 4210 7260 4290
rect 7340 4210 7660 4290
rect 7740 4210 8060 4290
rect 8140 4210 8460 4290
rect 8540 4210 8860 4290
rect 8940 4210 9260 4290
rect 9340 4210 9660 4290
rect 9740 4210 10100 4290
rect 2100 3890 10100 4210
rect 2100 3810 2460 3890
rect 2540 3810 2860 3890
rect 2940 3810 3260 3890
rect 3340 3810 3660 3890
rect 3740 3810 4060 3890
rect 4140 3810 4460 3890
rect 4540 3810 4860 3890
rect 4940 3810 5260 3890
rect 5340 3810 5660 3890
rect 5740 3810 6060 3890
rect 6140 3810 6460 3890
rect 6540 3810 6860 3890
rect 6940 3810 7260 3890
rect 7340 3810 7660 3890
rect 7740 3810 8060 3890
rect 8140 3810 8460 3890
rect 8540 3810 8860 3890
rect 8940 3810 9260 3890
rect 9340 3810 9660 3890
rect 9740 3810 10100 3890
rect 2100 3490 10100 3810
rect 2100 3410 2460 3490
rect 2540 3410 2860 3490
rect 2940 3410 3260 3490
rect 3340 3410 3660 3490
rect 3740 3410 4060 3490
rect 4140 3410 4460 3490
rect 4540 3410 4860 3490
rect 4940 3410 5260 3490
rect 5340 3410 5660 3490
rect 5740 3410 6060 3490
rect 6140 3410 6460 3490
rect 6540 3410 6860 3490
rect 6940 3410 7260 3490
rect 7340 3410 7660 3490
rect 7740 3410 8060 3490
rect 8140 3410 8460 3490
rect 8540 3410 8860 3490
rect 8940 3410 9260 3490
rect 9340 3410 9660 3490
rect 9740 3410 10100 3490
rect 2100 3090 10100 3410
rect 2100 3010 2460 3090
rect 2540 3010 2860 3090
rect 2940 3010 3260 3090
rect 3340 3010 3660 3090
rect 3740 3010 4060 3090
rect 4140 3010 4460 3090
rect 4540 3010 4860 3090
rect 4940 3010 5260 3090
rect 5340 3010 5660 3090
rect 5740 3010 6060 3090
rect 6140 3010 6460 3090
rect 6540 3010 6860 3090
rect 6940 3010 7260 3090
rect 7340 3010 7660 3090
rect 7740 3010 8060 3090
rect 8140 3010 8460 3090
rect 8540 3010 8860 3090
rect 8940 3010 9260 3090
rect 9340 3010 9660 3090
rect 9740 3010 10100 3090
rect 2100 2690 10100 3010
rect 2100 2610 2460 2690
rect 2540 2610 2860 2690
rect 2940 2610 3260 2690
rect 3340 2610 3660 2690
rect 3740 2610 4060 2690
rect 4140 2610 4460 2690
rect 4540 2610 4860 2690
rect 4940 2610 5260 2690
rect 5340 2610 5660 2690
rect 5740 2610 6060 2690
rect 6140 2610 6460 2690
rect 6540 2610 6860 2690
rect 6940 2610 7260 2690
rect 7340 2610 7660 2690
rect 7740 2610 8060 2690
rect 8140 2610 8460 2690
rect 8540 2610 8860 2690
rect 8940 2610 9260 2690
rect 9340 2610 9660 2690
rect 9740 2610 10100 2690
rect 2100 2290 10100 2610
rect 2100 2210 2460 2290
rect 2540 2210 2860 2290
rect 2940 2210 3260 2290
rect 3340 2210 3660 2290
rect 3740 2210 4060 2290
rect 4140 2210 4460 2290
rect 4540 2210 4860 2290
rect 4940 2210 5260 2290
rect 5340 2210 5660 2290
rect 5740 2210 6060 2290
rect 6140 2210 6460 2290
rect 6540 2210 6860 2290
rect 6940 2210 7260 2290
rect 7340 2210 7660 2290
rect 7740 2210 8060 2290
rect 8140 2210 8460 2290
rect 8540 2210 8860 2290
rect 8940 2210 9260 2290
rect 9340 2210 9660 2290
rect 9740 2210 10100 2290
rect 2100 1890 10100 2210
rect 2100 1810 2460 1890
rect 2540 1810 2860 1890
rect 2940 1810 3260 1890
rect 3340 1810 3660 1890
rect 3740 1810 4060 1890
rect 4140 1810 4460 1890
rect 4540 1810 4860 1890
rect 4940 1810 5260 1890
rect 5340 1810 5660 1890
rect 5740 1810 6060 1890
rect 6140 1810 6460 1890
rect 6540 1810 6860 1890
rect 6940 1810 7260 1890
rect 7340 1810 7660 1890
rect 7740 1810 8060 1890
rect 8140 1810 8460 1890
rect 8540 1810 8860 1890
rect 8940 1810 9260 1890
rect 9340 1810 9660 1890
rect 9740 1810 10100 1890
rect 2100 1490 10100 1810
rect 2100 1410 2460 1490
rect 2540 1410 2860 1490
rect 2940 1410 3260 1490
rect 3340 1410 3660 1490
rect 3740 1410 4060 1490
rect 4140 1410 4460 1490
rect 4540 1410 4860 1490
rect 4940 1410 5260 1490
rect 5340 1410 5660 1490
rect 5740 1410 6060 1490
rect 6140 1410 6460 1490
rect 6540 1410 6860 1490
rect 6940 1410 7260 1490
rect 7340 1410 7660 1490
rect 7740 1410 8060 1490
rect 8140 1410 8460 1490
rect 8540 1410 8860 1490
rect 8940 1410 9260 1490
rect 9340 1410 9660 1490
rect 9740 1410 10100 1490
rect 2100 1090 10100 1410
rect 2100 1010 2460 1090
rect 2540 1010 2860 1090
rect 2940 1010 3260 1090
rect 3340 1010 3660 1090
rect 3740 1010 4060 1090
rect 4140 1010 4460 1090
rect 4540 1010 4860 1090
rect 4940 1010 5260 1090
rect 5340 1010 5660 1090
rect 5740 1010 6060 1090
rect 6140 1010 6460 1090
rect 6540 1010 6860 1090
rect 6940 1010 7260 1090
rect 7340 1010 7660 1090
rect 7740 1010 8060 1090
rect 8140 1010 8460 1090
rect 8540 1010 8860 1090
rect 8940 1010 9260 1090
rect 9340 1010 9660 1090
rect 9740 1010 10100 1090
rect 2100 690 10100 1010
rect 2100 610 2460 690
rect 2540 610 2860 690
rect 2940 610 3260 690
rect 3340 610 3660 690
rect 3740 610 4060 690
rect 4140 610 4460 690
rect 4540 610 4860 690
rect 4940 610 5260 690
rect 5340 610 5660 690
rect 5740 610 6060 690
rect 6140 610 6460 690
rect 6540 610 6860 690
rect 6940 610 7260 690
rect 7340 610 7660 690
rect 7740 610 8060 690
rect 8140 610 8460 690
rect 8540 610 8860 690
rect 8940 610 9260 690
rect 9340 610 9660 690
rect 9740 610 10100 690
rect 2100 250 10100 610
<< labels >>
flabel space 6100 4250 6100 4250 0 FreeSans 5000 0 0 0 PIC_0.PAD
flabel m3p 100 24240 100 24240 0 FreeSans 5000 0 0 0 PIC_0.VDD
flabel m3p 100 30845 100 30845 0 FreeSans 5000 0 0 0 PIC_0.VDD
flabel m3p 100 33090 100 33090 0 FreeSans 5000 0 0 0 PIC_0.VSS
flabel m3p 100 12910 100 12910 0 FreeSans 5000 0 0 0 PIC_0.VSS
flabel m2p 11560 34450 11560 34450 0 FreeSans 2000 0 0 0 PIC_0.Y
<< end >>
