magic
tech scmos
magscale 1 2
timestamp 1702508443
<< nwell >>
rect -12 154 92 272
<< ntransistor >>
rect 18 14 22 54
rect 38 14 42 54
rect 58 14 62 54
<< ptransistor >>
rect 20 166 24 246
rect 34 166 38 246
rect 54 206 58 246
<< ndiffusion >>
rect 16 14 18 54
rect 22 42 38 54
rect 22 14 24 42
rect 36 14 38 42
rect 42 14 44 54
rect 56 14 58 54
rect 62 14 64 54
<< pdiffusion >>
rect 18 166 20 246
rect 24 166 34 246
rect 38 166 40 246
rect 52 206 54 246
rect 58 206 60 246
<< ndcontact >>
rect 4 14 16 54
rect 24 14 36 42
rect 44 14 56 54
rect 64 14 76 54
<< pdcontact >>
rect 6 166 18 246
rect 40 166 52 246
rect 60 206 72 246
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 254 86 266
<< polysilicon >>
rect 20 246 24 250
rect 34 246 38 250
rect 54 246 58 250
rect 54 184 58 206
rect 20 164 24 166
rect 12 160 24 164
rect 34 164 38 166
rect 34 160 42 164
rect 12 129 16 160
rect 12 66 16 117
rect 38 103 42 160
rect 36 91 42 103
rect 12 58 22 66
rect 18 54 22 58
rect 38 54 42 91
rect 60 74 64 184
rect 58 68 64 74
rect 58 54 62 68
rect 18 10 22 14
rect 38 10 42 14
rect 58 10 62 14
<< polycontact >>
rect 58 184 70 196
rect 4 117 16 129
rect 24 91 36 103
rect 64 91 76 103
<< metal1 >>
rect -6 266 86 268
rect -6 252 86 254
rect 6 246 18 252
rect 60 246 72 252
rect 52 166 56 176
rect 48 117 56 166
rect 48 74 56 103
rect 48 68 72 74
rect 4 54 56 57
rect 16 48 44 54
rect 64 54 72 68
rect 24 8 36 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
rect 43 103 57 117
rect 63 103 77 117
<< metal2 >>
rect 26 117 34 134
rect 66 117 74 134
rect 6 86 14 103
rect 46 86 54 103
<< m1p >>
rect -6 252 86 268
rect -6 -8 86 8
<< m2p >>
rect 26 119 34 134
rect 66 119 74 134
rect 6 86 14 101
rect 46 86 54 101
<< labels >>
rlabel metal2 10 90 10 90 5 A
port 1 n signal input
rlabel metal2 30 130 30 130 5 B
port 2 n signal input
rlabel metal2 70 132 70 132 1 C
port 3 n signal input
rlabel metal2 50 90 50 90 1 Y
port 4 n signal output
rlabel metal1 -6 252 86 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 86 8 0 gnd
port 6 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 80 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
