magic
tech scmos
magscale 1 3
timestamp 1725342160
<< diffusion >>
rect 31 221 219 239
rect 11 31 29 219
rect 77 77 173 173
rect 221 31 239 219
rect 31 11 219 29
<< ndiffusion >>
rect 75 173 175 175
rect 75 77 77 173
rect 173 77 175 173
rect 75 75 175 77
<< psubstratepdiff >>
rect 10 239 240 240
rect 10 221 31 239
rect 219 221 240 239
rect 10 220 240 221
rect 10 219 30 220
rect 10 31 11 219
rect 29 31 30 219
rect 220 219 240 220
rect 10 30 30 31
rect 220 31 221 219
rect 239 31 240 219
rect 220 30 240 31
rect 10 29 240 30
rect 10 11 31 29
rect 219 11 240 29
rect 10 10 240 11
<< metal1 >>
rect 10 220 240 240
rect 10 30 30 220
rect 75 75 175 175
rect 220 30 240 220
rect 10 10 240 30
<< end >>
