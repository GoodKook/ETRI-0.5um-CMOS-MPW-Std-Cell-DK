magic
tech scmos
timestamp 1727493435
<< nwell >>
rect -3 77 13 136
<< psubstratepcontact >>
rect 0 -3 10 3
<< nsubstratencontact >>
rect 0 127 10 133
<< metal1 >>
rect 0 133 10 134
rect 0 126 10 127
rect 0 3 10 4
rect 0 -4 10 -3
<< labels >>
rlabel metal1 0 133 10 134 0 vdd
port 0 nsew power bidirectional abutment
rlabel metal1 0 127 10 133 0 vdd
port 0 nsew power bidirectional abutment
rlabel metal1 0 126 10 127 0 vdd
port 0 nsew power bidirectional abutment
rlabel metal1 0 3 10 4 0 gnd
port 1 nsew ground bidirectional abutment
rlabel metal1 0 -3 10 3 0 gnd
port 1 nsew ground bidirectional abutment
rlabel metal1 0 -4 10 -3 0 gnd
port 1 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 10 130
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
