magic
tech scmos
magscale 1 3
timestamp 1725343477
<< checkpaint >>
rect -19 289 289 309
rect -39 285 309 289
rect -40 -15 310 285
rect -39 -19 309 -15
rect -19 -39 289 -19
<< nwell >>
rect 0 0 270 270
<< psubstratepdiff >>
rect 85 85 185 185
<< nsubstratendiff >>
rect 20 230 250 250
rect 20 40 40 230
rect 230 40 250 230
rect 20 20 250 40
<< genericcontact >>
rect 45 230 225 250
rect 20 45 40 225
rect 85 85 185 185
rect 230 45 250 225
rect 45 20 225 40
<< metal1 >>
rect 20 230 250 250
rect 20 40 40 230
rect 85 85 185 185
rect 230 40 250 230
rect 20 20 250 40
<< end >>
