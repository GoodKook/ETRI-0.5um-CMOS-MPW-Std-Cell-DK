magic
tech scmos
magscale 1 2
timestamp 1701862152
<< checkpaint >>
rect -14 142 74 159
rect -34 61 94 142
<< nwell >>
rect -12 152 74 272
<< ntransistor >>
rect 18 14 22 34
rect 38 14 42 34
<< ptransistor >>
rect 18 166 22 246
rect 32 166 36 246
<< ndiffusion >>
rect 16 14 18 34
rect 22 14 24 34
rect 36 14 38 34
rect 42 14 44 34
<< pdiffusion >>
rect 16 166 18 246
rect 22 166 32 246
rect 36 166 38 246
<< ndcontact >>
rect 4 14 16 34
rect 24 14 36 34
rect 44 14 56 34
<< pdcontact >>
rect 4 166 16 246
rect 38 166 50 246
<< psubstratepcontact >>
rect -6 -6 66 6
<< nsubstratencontact >>
rect -6 254 66 266
<< polysilicon >>
rect 18 246 22 250
rect 32 246 36 250
rect 18 129 22 166
rect 32 164 36 166
rect 32 160 42 164
rect 17 117 22 129
rect 18 34 22 117
rect 38 129 42 160
rect 38 117 44 129
rect 38 34 42 117
rect 18 10 22 14
rect 38 10 42 14
<< polycontact >>
rect 5 117 17 129
rect 44 117 56 129
<< metal1 >>
rect -6 266 66 268
rect -6 252 66 254
rect 4 246 16 252
rect 26 166 38 174
rect 26 117 32 166
rect 26 34 32 103
rect 4 8 16 14
rect 44 8 56 14
rect -6 6 66 8
rect -6 -8 66 -6
<< m2contact >>
rect 3 103 17 117
rect 23 103 37 117
rect 43 103 57 117
<< metal2 >>
rect 26 117 34 134
rect 6 86 14 103
rect 46 86 54 103
<< m1p >>
rect -6 252 66 268
rect -6 -8 66 8
<< m2p >>
rect 26 119 34 134
rect 6 86 14 101
rect 46 86 54 101
<< labels >>
rlabel metal2 10 90 10 90 1 A
port 1 n signal input
rlabel metal2 50 88 50 88 5 B
port 2 n signal input
rlabel metal2 30 130 30 130 1 Y
port 3 n signal output
rlabel metal1 -6 252 66 268 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal1 -6 -8 66 8 0 gnd
port 5 nsew ground bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 60 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
