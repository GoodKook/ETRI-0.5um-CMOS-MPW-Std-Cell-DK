* NGSPICE file created from DFFPOSX1.ext - technology: scmos

.subckt DFFPOSX1 D CLK Q vdd gnd
M1000 a_44_12# a_4_12# a_34_12# gnd nfet w=3u l=0.6u
+  ad=3.15p pd=5.1u as=1.35p ps=3.9u
M1001 vdd Q a_152_168# vdd pfet w=3u l=0.6u
+  ad=9.450001p pd=13.8u as=1.35p ps=3.9u
M1002 gnd a_68_8# a_62_12# gnd nfet w=3u l=0.6u
+  ad=3.15p pd=5.1u as=1.35p ps=3.9u
M1003 a_152_12# a_4_12# a_132_12# gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=3.6p ps=5.4u
M1004 a_68_8# a_44_12# vdd vdd pfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=5.4p ps=7.8u
M1005 a_152_168# CLK a_132_12# vdd pfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=6.750001p ps=8.400001u
M1006 gnd CLK a_4_12# gnd nfet w=6u l=0.6u
+  ad=4.95p pd=7.8u as=9p ps=15.000001u
M1007 a_62_148# a_4_12# a_44_12# vdd pfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=5.4p ps=7.8u
M1008 gnd Q a_152_12# gnd nfet w=3u l=0.6u
+  ad=4.95p pd=7.8u as=1.35p ps=3.9u
M1009 a_34_148# D vdd vdd pfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=9.900001p ps=13.8u
M1010 vdd a_68_8# a_62_148# vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=3.6p ps=7.2u
M1011 a_132_12# a_4_12# a_122_148# vdd pfet w=6u l=0.6u
+  ad=6.750001p pd=8.400001u as=2.7p ps=6.9u
M1012 a_68_8# a_44_12# gnd gnd nfet w=3u l=0.6u
+  ad=4.5p pd=9u as=3.15p ps=5.1u
M1013 a_44_12# CLK a_34_148# vdd pfet w=6u l=0.6u
+  ad=5.4p pd=7.8u as=3.6p ps=7.2u
M1014 a_122_12# a_68_8# gnd gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=4.5p ps=9u
M1015 a_122_148# a_68_8# vdd vdd pfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=9p ps=15.000001u
M1016 Q a_132_12# vdd vdd pfet w=12u l=0.6u
+  ad=18p pd=27.000002u as=9.450001p ps=13.8u
M1017 a_34_12# D gnd gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=4.95p ps=7.8u
M1018 a_132_12# CLK a_122_12# gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=1.35p ps=3.9u
M1019 Q a_132_12# gnd gnd nfet w=6u l=0.6u
+  ad=9p pd=15.000001u as=4.95p ps=7.8u
M1020 vdd CLK a_4_12# vdd pfet w=12u l=0.6u
+  ad=9.900001p pd=13.8u as=18p ps=27.000002u
M1021 a_62_12# CLK a_44_12# gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=3.15p ps=5.1u
.ends

