magic
tech scmos
magscale 1 2
timestamp 1728305047
<< nwell >>
rect -12 134 112 252
<< ntransistor >>
rect 22 14 26 74
rect 30 14 34 74
rect 38 14 42 74
<< ptransistor >>
rect 21 186 25 226
rect 41 186 45 226
rect 61 186 65 226
<< ndiffusion >>
rect 20 14 22 74
rect 26 14 30 74
rect 34 14 38 74
rect 42 72 56 74
rect 42 14 44 72
<< pdiffusion >>
rect 19 186 21 226
rect 25 186 27 226
rect 39 186 41 226
rect 45 190 47 226
rect 59 190 61 226
rect 45 186 61 190
rect 65 186 67 226
<< ndcontact >>
rect 8 14 20 74
rect 44 14 56 72
<< pdcontact >>
rect 7 186 19 226
rect 27 186 39 226
rect 47 190 59 226
rect 67 186 79 226
<< psubstratepcontact >>
rect -6 -6 106 6
<< nsubstratencontact >>
rect -6 234 106 246
<< polysilicon >>
rect 21 226 25 230
rect 41 226 45 230
rect 61 226 65 230
rect 21 178 25 186
rect 10 174 25 178
rect 41 174 45 186
rect 10 143 16 174
rect 30 170 45 174
rect 30 163 36 170
rect 16 131 26 143
rect 22 74 26 131
rect 30 74 34 151
rect 61 143 65 186
rect 38 131 45 143
rect 57 131 65 143
rect 38 74 42 131
rect 22 10 26 14
rect 30 10 34 14
rect 38 10 42 14
<< polycontact >>
rect 24 151 36 163
rect 4 131 16 143
rect 45 131 57 143
<< metal1 >>
rect -6 246 106 248
rect -6 232 106 234
rect 7 226 19 232
rect 47 226 59 232
rect 28 184 39 186
rect 67 184 75 186
rect 28 178 75 184
rect 68 123 75 178
rect 66 81 74 109
rect 44 72 74 81
rect 56 70 74 72
rect 8 8 20 14
rect -6 6 106 8
rect -6 -8 106 -6
<< m2contact >>
rect 23 137 37 151
rect 3 117 17 131
rect 43 117 57 131
rect 63 109 77 123
<< metal2 >>
rect 23 123 37 137
rect 3 103 17 117
rect 43 103 57 117
rect 63 123 77 137
<< m1p >>
rect -6 232 106 248
rect -6 -8 106 8
<< m2p >>
rect 23 123 37 137
rect 63 123 77 137
rect 3 103 17 117
rect 43 103 57 117
<< labels >>
rlabel metal1 -6 -8 106 8 0 gnd
port 5 nsew ground bidirectional abutment
rlabel metal1 -6 232 106 248 0 vdd
port 4 nsew power bidirectional abutment
rlabel metal2 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal2 23 123 37 137 0 B
port 1 nsew signal input
rlabel metal2 43 103 57 117 0 C
port 2 nsew signal input
rlabel metal2 63 123 77 137 0 Y
port 3 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 100 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
