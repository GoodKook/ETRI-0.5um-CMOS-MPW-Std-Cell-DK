VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO fir_pe
  CLASS BLOCK ;
  FOREIGN fir_pe ;
  ORIGIN 6.000 6.000 ;
  SIZE 888.000 BY 834.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 0.600 819.300 885.450 821.700 ;
        RECT 876.450 743.700 885.450 819.300 ;
        RECT 0.600 741.300 885.450 743.700 ;
        RECT 876.450 665.700 885.450 741.300 ;
        RECT 0.600 663.300 885.450 665.700 ;
        RECT 876.450 587.700 885.450 663.300 ;
        RECT 0.600 585.300 885.450 587.700 ;
        RECT 876.450 509.700 885.450 585.300 ;
        RECT 0.600 507.300 885.450 509.700 ;
        RECT 876.450 431.700 885.450 507.300 ;
        RECT 0.600 429.300 885.450 431.700 ;
        RECT 876.450 353.700 885.450 429.300 ;
        RECT 0.600 351.300 885.450 353.700 ;
        RECT 876.450 275.700 885.450 351.300 ;
        RECT 0.600 273.300 885.450 275.700 ;
        RECT 876.450 197.700 885.450 273.300 ;
        RECT 0.600 195.300 885.450 197.700 ;
        RECT 876.450 119.700 885.450 195.300 ;
        RECT 0.600 117.300 885.450 119.700 ;
        RECT 876.450 41.700 885.450 117.300 ;
        RECT 0.600 39.300 885.450 41.700 ;
        RECT 876.450 0.300 885.450 39.300 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.450 782.700 -0.450 821.700 ;
        RECT -9.450 780.300 875.400 782.700 ;
        RECT -9.450 704.700 -0.450 780.300 ;
        RECT -9.450 702.300 875.400 704.700 ;
        RECT -9.450 626.700 -0.450 702.300 ;
        RECT -9.450 624.300 875.400 626.700 ;
        RECT -9.450 548.700 -0.450 624.300 ;
        RECT -9.450 546.300 875.400 548.700 ;
        RECT -9.450 470.700 -0.450 546.300 ;
        RECT -9.450 468.300 875.400 470.700 ;
        RECT -9.450 392.700 -0.450 468.300 ;
        RECT -9.450 390.300 875.400 392.700 ;
        RECT -9.450 314.700 -0.450 390.300 ;
        RECT -9.450 312.300 875.400 314.700 ;
        RECT -9.450 236.700 -0.450 312.300 ;
        RECT -9.450 234.300 875.400 236.700 ;
        RECT -9.450 158.700 -0.450 234.300 ;
        RECT -9.450 156.300 875.400 158.700 ;
        RECT -9.450 80.700 -0.450 156.300 ;
        RECT -9.450 78.300 875.400 80.700 ;
        RECT -9.450 2.700 -0.450 78.300 ;
        RECT -9.450 0.300 875.400 2.700 ;
    END
  END vdd
  PIN Cin[5]
    PORT
      LAYER metal1 ;
        RECT 454.950 297.450 457.050 298.050 ;
        RECT 463.950 297.450 466.050 298.050 ;
        RECT 454.950 296.550 466.050 297.450 ;
        RECT 454.950 295.950 457.050 296.550 ;
        RECT 463.950 295.950 466.050 296.550 ;
        RECT 445.950 294.450 448.050 295.050 ;
        RECT 440.550 293.550 448.050 294.450 ;
        RECT 440.550 289.050 441.450 293.550 ;
        RECT 445.950 292.950 448.050 293.550 ;
        RECT 436.950 287.550 441.450 289.050 ;
        RECT 436.950 286.950 441.000 287.550 ;
        RECT 796.950 246.450 799.050 247.050 ;
        RECT 805.950 246.450 808.050 247.050 ;
        RECT 796.950 245.550 808.050 246.450 ;
        RECT 796.950 244.950 799.050 245.550 ;
        RECT 805.950 244.950 808.050 245.550 ;
      LAYER metal2 ;
        RECT 538.950 316.950 541.050 319.050 ;
        RECT 539.400 304.050 540.450 316.950 ;
        RECT 613.950 316.800 616.050 318.900 ;
        RECT 463.950 301.950 466.050 304.050 ;
        RECT 538.950 301.950 541.050 304.050 ;
        RECT 464.400 298.050 465.450 301.950 ;
        RECT 614.400 298.050 615.450 316.800 ;
        RECT 373.950 293.100 376.050 295.200 ;
        RECT 379.950 293.100 382.050 295.200 ;
        RECT 374.400 292.350 375.600 293.100 ;
        RECT 380.400 277.050 381.450 293.100 ;
        RECT 445.950 292.950 448.050 298.050 ;
        RECT 454.950 295.200 457.050 298.050 ;
        RECT 463.950 295.950 466.050 298.050 ;
        RECT 454.800 294.000 457.050 295.200 ;
        RECT 613.950 294.000 616.050 298.050 ;
        RECT 454.800 293.100 456.900 294.000 ;
        RECT 455.400 292.350 456.600 293.100 ;
        RECT 614.400 292.350 615.600 294.000 ;
        RECT 637.950 292.950 640.050 295.050 ;
        RECT 643.950 293.100 646.050 295.200 ;
        RECT 436.950 286.950 439.050 289.050 ;
        RECT 379.950 274.950 382.050 277.050 ;
        RECT 437.400 274.050 438.450 286.950 ;
        RECT 638.400 280.050 639.450 292.950 ;
        RECT 644.400 292.350 645.600 293.100 ;
        RECT 871.950 292.800 874.050 294.900 ;
        RECT 872.400 286.050 873.450 292.800 ;
        RECT 853.950 283.950 856.050 286.050 ;
        RECT 871.950 283.950 874.050 286.050 ;
        RECT 637.950 277.950 640.050 280.050 ;
        RECT 664.950 277.950 667.050 280.050 ;
        RECT 436.950 271.950 439.050 274.050 ;
        RECT 665.400 247.050 666.450 277.950 ;
        RECT 854.400 265.050 855.450 283.950 ;
        RECT 853.950 262.950 856.050 265.050 ;
        RECT 826.950 253.950 829.050 256.050 ;
        RECT 796.800 249.000 798.900 250.050 ;
        RECT 796.800 247.950 799.050 249.000 ;
        RECT 664.950 244.950 667.050 247.050 ;
        RECT 796.950 244.950 799.050 247.950 ;
        RECT 827.400 247.050 828.450 253.950 ;
        RECT 805.950 244.950 811.050 247.050 ;
        RECT 826.950 244.950 829.050 247.050 ;
      LAYER metal3 ;
        RECT 538.950 318.600 541.050 319.050 ;
        RECT 613.950 318.600 616.050 318.900 ;
        RECT 538.950 317.400 616.050 318.600 ;
        RECT 538.950 316.950 541.050 317.400 ;
        RECT 613.950 316.800 616.050 317.400 ;
        RECT 463.950 303.600 466.050 304.050 ;
        RECT 538.950 303.600 541.050 304.050 ;
        RECT 463.950 302.400 541.050 303.600 ;
        RECT 463.950 301.950 466.050 302.400 ;
        RECT 538.950 301.950 541.050 302.400 ;
        RECT 373.950 294.750 376.050 295.200 ;
        RECT 379.950 294.750 382.050 295.200 ;
        RECT 373.950 293.550 382.050 294.750 ;
        RECT 445.950 294.600 448.050 298.050 ;
        RECT 613.950 297.600 616.050 298.050 ;
        RECT 613.950 296.400 642.600 297.600 ;
        RECT 613.950 295.950 616.050 296.400 ;
        RECT 454.800 294.600 456.900 295.200 ;
        RECT 641.400 295.050 642.600 296.400 ;
        RECT 445.950 294.000 456.900 294.600 ;
        RECT 373.950 293.100 376.050 293.550 ;
        RECT 379.950 293.100 382.050 293.550 ;
        RECT 446.400 293.400 456.900 294.000 ;
        RECT 454.800 293.100 456.900 293.400 ;
        RECT 637.950 294.600 642.600 295.050 ;
        RECT 643.950 294.600 646.050 295.200 ;
        RECT 637.950 293.400 646.050 294.600 ;
        RECT 637.950 292.950 642.000 293.400 ;
        RECT 643.950 293.100 646.050 293.400 ;
        RECT 871.950 294.600 874.050 294.900 ;
        RECT 871.950 293.400 882.600 294.600 ;
        RECT 871.950 292.800 874.050 293.400 ;
        RECT 853.950 285.600 856.050 286.050 ;
        RECT 871.950 285.600 874.050 286.050 ;
        RECT 853.950 284.400 874.050 285.600 ;
        RECT 853.950 283.950 856.050 284.400 ;
        RECT 871.950 283.950 874.050 284.400 ;
        RECT 637.950 279.600 640.050 280.050 ;
        RECT 664.950 279.600 667.050 280.050 ;
        RECT 637.950 278.400 667.050 279.600 ;
        RECT 637.950 277.950 640.050 278.400 ;
        RECT 664.950 277.950 667.050 278.400 ;
        RECT 379.950 276.600 382.050 277.050 ;
        RECT 379.950 275.400 402.600 276.600 ;
        RECT 379.950 274.950 382.050 275.400 ;
        RECT 401.400 273.600 402.600 275.400 ;
        RECT 436.950 273.600 439.050 274.050 ;
        RECT 401.400 272.400 439.050 273.600 ;
        RECT 436.950 271.950 439.050 272.400 ;
        RECT 853.950 262.950 856.050 265.050 ;
        RECT 826.950 255.600 829.050 256.050 ;
        RECT 854.400 255.600 855.600 262.950 ;
        RECT 826.950 254.400 855.600 255.600 ;
        RECT 826.950 253.950 829.050 254.400 ;
        RECT 796.800 249.600 798.900 250.050 ;
        RECT 683.400 248.400 798.900 249.600 ;
        RECT 664.950 246.600 667.050 247.050 ;
        RECT 683.400 246.600 684.600 248.400 ;
        RECT 796.800 247.950 798.900 248.400 ;
        RECT 664.950 245.400 684.600 246.600 ;
        RECT 808.950 246.600 811.050 247.050 ;
        RECT 826.950 246.600 829.050 247.050 ;
        RECT 808.950 245.400 829.050 246.600 ;
        RECT 664.950 244.950 667.050 245.400 ;
        RECT 808.950 244.950 811.050 245.400 ;
        RECT 826.950 244.950 829.050 245.400 ;
    END
  END Cin[5]
  PIN Cin[4]
    PORT
      LAYER metal1 ;
        RECT 534.000 339.450 538.050 340.050 ;
        RECT 533.550 337.950 538.050 339.450 ;
        RECT 667.950 339.450 670.050 340.050 ;
        RECT 667.950 338.550 675.450 339.450 ;
        RECT 667.950 337.950 670.050 338.550 ;
        RECT 533.550 334.050 534.450 337.950 ;
        RECT 674.550 334.050 675.450 338.550 ;
        RECT 533.550 332.550 538.050 334.050 ;
        RECT 674.550 332.550 679.050 334.050 ;
        RECT 534.000 331.950 538.050 332.550 ;
        RECT 675.000 331.950 679.050 332.550 ;
        RECT 676.950 292.950 679.050 295.050 ;
        RECT 677.550 289.050 678.450 292.950 ;
        RECT 677.550 287.550 682.050 289.050 ;
        RECT 678.000 286.950 682.050 287.550 ;
      LAYER metal2 ;
        RECT 641.400 410.400 642.600 412.650 ;
        RECT 671.400 411.000 672.600 412.650 ;
        RECT 641.400 409.050 642.450 410.400 ;
        RECT 640.950 406.950 643.050 409.050 ;
        RECT 670.950 406.950 673.050 411.000 ;
        RECT 715.950 406.950 718.050 409.050 ;
        RECT 641.400 388.050 642.450 406.950 ;
        RECT 565.950 385.950 568.050 388.050 ;
        RECT 640.950 385.950 643.050 388.050 ;
        RECT 649.950 385.950 652.050 388.050 ;
        RECT 566.400 373.050 567.450 385.950 ;
        RECT 565.950 370.950 568.050 373.050 ;
        RECT 650.400 364.050 651.450 385.950 ;
        RECT 716.400 375.450 717.450 406.950 ;
        RECT 716.400 374.400 720.450 375.450 ;
        RECT 719.400 372.600 720.450 374.400 ;
        RECT 719.400 370.350 720.600 372.600 ;
        RECT 535.950 361.950 538.050 364.050 ;
        RECT 649.950 361.950 652.050 364.050 ;
        RECT 667.950 361.950 670.050 364.050 ;
        RECT 536.400 340.050 537.450 361.950 ;
        RECT 650.400 355.050 651.450 361.950 ;
        RECT 631.950 352.950 634.050 355.050 ;
        RECT 649.950 352.950 652.050 355.050 ;
        RECT 535.950 337.950 538.050 340.050 ;
        RECT 535.950 331.950 538.050 334.050 ;
        RECT 530.400 287.400 531.600 289.650 ;
        RECT 530.400 286.050 531.450 287.400 ;
        RECT 536.400 286.050 537.450 331.950 ;
        RECT 632.400 294.600 633.450 352.950 ;
        RECT 668.400 340.050 669.450 361.950 ;
        RECT 667.950 337.950 670.050 340.050 ;
        RECT 676.950 331.950 679.050 334.050 ;
        RECT 677.400 295.050 678.450 331.950 ;
        RECT 632.400 292.350 633.600 294.600 ;
        RECT 676.950 292.950 679.050 295.050 ;
        RECT 679.950 286.950 682.050 289.050 ;
        RECT 529.950 283.950 532.050 286.050 ;
        RECT 535.950 283.950 538.050 286.050 ;
        RECT 530.400 265.050 531.450 283.950 ;
        RECT 680.400 271.050 681.450 286.950 ;
        RECT 679.950 268.950 682.050 271.050 ;
        RECT 706.950 268.950 709.050 271.050 ;
        RECT 707.400 265.200 708.450 268.950 ;
        RECT 529.950 262.950 532.050 265.050 ;
        RECT 706.950 263.100 709.050 265.200 ;
        RECT 427.950 259.800 430.050 261.900 ;
        RECT 436.950 260.100 439.050 262.200 ;
        RECT 428.400 253.050 429.450 259.800 ;
        RECT 437.400 259.350 438.600 260.100 ;
        RECT 520.950 253.950 523.050 256.050 ;
        RECT 721.950 253.950 724.050 256.050 ;
        RECT 427.950 250.950 430.050 253.050 ;
        RECT 433.950 250.950 436.050 253.050 ;
        RECT 434.400 217.200 435.450 250.950 ;
        RECT 417.000 216.600 421.050 217.050 ;
        RECT 416.400 214.950 421.050 216.600 ;
        RECT 433.950 215.100 436.050 217.200 ;
        RECT 416.400 214.350 417.600 214.950 ;
        RECT 434.400 214.350 435.600 215.100 ;
        RECT 424.950 208.950 427.050 211.050 ;
        RECT 521.400 210.900 522.450 253.950 ;
        RECT 722.400 226.050 723.450 253.950 ;
        RECT 823.950 226.950 826.050 229.050 ;
        RECT 721.950 223.950 724.050 226.050 ;
        RECT 748.950 223.950 751.050 226.050 ;
        RECT 749.400 220.050 750.450 223.950 ;
        RECT 824.400 223.050 825.450 226.950 ;
        RECT 823.950 220.950 826.050 223.050 ;
        RECT 748.950 217.950 751.050 220.050 ;
        RECT 530.400 210.900 531.600 211.650 ;
        RECT 425.400 187.050 426.450 208.950 ;
        RECT 520.950 208.800 523.050 210.900 ;
        RECT 529.950 208.800 532.050 210.900 ;
        RECT 770.400 210.000 771.600 211.650 ;
        RECT 521.400 187.200 522.450 208.800 ;
        RECT 769.950 205.950 772.050 210.000 ;
        RECT 800.400 209.400 801.600 211.650 ;
        RECT 800.400 208.050 801.450 209.400 ;
        RECT 796.950 206.400 801.450 208.050 ;
        RECT 796.950 205.950 801.000 206.400 ;
        RECT 424.950 184.950 427.050 187.050 ;
        RECT 520.950 185.100 523.050 187.200 ;
      LAYER metal3 ;
        RECT 640.950 408.600 643.050 409.050 ;
        RECT 670.950 408.600 673.050 409.050 ;
        RECT 715.950 408.600 718.050 409.050 ;
        RECT 640.950 407.400 718.050 408.600 ;
        RECT 640.950 406.950 643.050 407.400 ;
        RECT 670.950 406.950 673.050 407.400 ;
        RECT 715.950 406.950 718.050 407.400 ;
        RECT 565.950 387.600 568.050 388.050 ;
        RECT 640.950 387.600 643.050 388.050 ;
        RECT 649.950 387.600 652.050 388.050 ;
        RECT 565.950 386.400 652.050 387.600 ;
        RECT 565.950 385.950 568.050 386.400 ;
        RECT 640.950 385.950 643.050 386.400 ;
        RECT 649.950 385.950 652.050 386.400 ;
        RECT 565.950 369.600 568.050 373.050 ;
        RECT 557.400 369.000 568.050 369.600 ;
        RECT 557.400 368.400 567.600 369.000 ;
        RECT 557.400 366.600 558.600 368.400 ;
        RECT 548.400 365.400 558.600 366.600 ;
        RECT 535.950 363.600 538.050 364.050 ;
        RECT 548.400 363.600 549.600 365.400 ;
        RECT 535.950 362.400 549.600 363.600 ;
        RECT 649.950 363.600 652.050 364.050 ;
        RECT 667.950 363.600 670.050 364.050 ;
        RECT 649.950 362.400 670.050 363.600 ;
        RECT 535.950 361.950 538.050 362.400 ;
        RECT 649.950 361.950 652.050 362.400 ;
        RECT 667.950 361.950 670.050 362.400 ;
        RECT 631.950 354.600 634.050 355.050 ;
        RECT 649.950 354.600 652.050 355.050 ;
        RECT 631.950 353.400 652.050 354.600 ;
        RECT 631.950 352.950 634.050 353.400 ;
        RECT 649.950 352.950 652.050 353.400 ;
        RECT 529.950 285.600 532.050 286.050 ;
        RECT 535.950 285.600 538.050 286.050 ;
        RECT 529.950 284.400 538.050 285.600 ;
        RECT 529.950 283.950 532.050 284.400 ;
        RECT 535.950 283.950 538.050 284.400 ;
        RECT 679.950 270.600 682.050 271.050 ;
        RECT 706.950 270.600 709.050 271.050 ;
        RECT 679.950 269.400 709.050 270.600 ;
        RECT 679.950 268.950 682.050 269.400 ;
        RECT 706.950 268.950 709.050 269.400 ;
        RECT 529.950 264.600 532.050 265.050 ;
        RECT 524.400 263.400 532.050 264.600 ;
        RECT 427.950 261.750 430.050 261.900 ;
        RECT 436.950 261.750 439.050 262.200 ;
        RECT 427.950 260.550 439.050 261.750 ;
        RECT 524.400 261.600 525.600 263.400 ;
        RECT 529.950 262.950 532.050 263.400 ;
        RECT 706.950 264.600 709.050 265.200 ;
        RECT 706.950 263.400 720.600 264.600 ;
        RECT 706.950 263.100 709.050 263.400 ;
        RECT 427.950 259.800 430.050 260.550 ;
        RECT 436.950 260.100 439.050 260.550 ;
        RECT 521.400 260.400 525.600 261.600 ;
        RECT 719.400 261.600 720.600 263.400 ;
        RECT 719.400 260.400 723.600 261.600 ;
        RECT 521.400 256.050 522.600 260.400 ;
        RECT 722.400 256.050 723.600 260.400 ;
        RECT 520.950 253.950 523.050 256.050 ;
        RECT 721.950 253.950 724.050 256.050 ;
        RECT 427.950 252.600 430.050 253.050 ;
        RECT 433.950 252.600 436.050 253.050 ;
        RECT 427.950 251.400 436.050 252.600 ;
        RECT 427.950 250.950 430.050 251.400 ;
        RECT 433.950 250.950 436.050 251.400 ;
        RECT 823.950 228.600 826.050 229.050 ;
        RECT 770.400 227.400 826.050 228.600 ;
        RECT 721.950 225.600 724.050 226.050 ;
        RECT 748.950 225.600 751.050 226.050 ;
        RECT 770.400 225.600 771.600 227.400 ;
        RECT 823.950 226.950 826.050 227.400 ;
        RECT 721.950 224.400 771.600 225.600 ;
        RECT 721.950 223.950 724.050 224.400 ;
        RECT 748.950 223.950 751.050 224.400 ;
        RECT 823.950 222.600 826.050 223.050 ;
        RECT 823.950 221.400 882.600 222.600 ;
        RECT 823.950 220.950 826.050 221.400 ;
        RECT 748.950 219.600 751.050 220.050 ;
        RECT 748.950 218.400 762.600 219.600 ;
        RECT 748.950 217.950 751.050 218.400 ;
        RECT 418.950 213.600 421.050 217.050 ;
        RECT 433.950 215.100 436.050 217.200 ;
        RECT 761.400 216.600 762.600 218.400 ;
        RECT 761.400 215.400 774.600 216.600 ;
        RECT 881.400 215.400 882.600 221.400 ;
        RECT 434.400 213.600 435.600 215.100 ;
        RECT 418.950 213.000 435.600 213.600 ;
        RECT 419.400 212.400 435.600 213.000 ;
        RECT 424.950 208.950 427.050 212.400 ;
        RECT 520.950 210.450 523.050 210.900 ;
        RECT 529.950 210.450 532.050 210.900 ;
        RECT 520.950 209.250 532.050 210.450 ;
        RECT 520.950 208.800 523.050 209.250 ;
        RECT 529.950 208.800 532.050 209.250 ;
        RECT 773.400 208.050 774.600 215.400 ;
        RECT 769.950 207.600 774.600 208.050 ;
        RECT 796.950 207.600 799.050 208.050 ;
        RECT 769.950 206.400 799.050 207.600 ;
        RECT 769.950 205.950 774.000 206.400 ;
        RECT 796.950 205.950 799.050 206.400 ;
        RECT 424.950 186.600 427.050 187.050 ;
        RECT 520.950 186.600 523.050 187.200 ;
        RECT 424.950 185.400 523.050 186.600 ;
        RECT 424.950 184.950 427.050 185.400 ;
        RECT 520.950 185.100 523.050 185.400 ;
    END
  END Cin[4]
  PIN Cin[3]
    PORT
      LAYER metal1 ;
        RECT 784.950 366.450 787.050 367.050 ;
        RECT 793.950 366.450 796.050 367.050 ;
        RECT 784.950 365.550 796.050 366.450 ;
        RECT 784.950 364.950 787.050 365.550 ;
        RECT 793.950 364.950 796.050 365.550 ;
        RECT 780.000 339.450 784.050 340.050 ;
        RECT 779.550 337.950 784.050 339.450 ;
        RECT 779.550 334.050 780.450 337.950 ;
        RECT 779.550 332.550 784.050 334.050 ;
        RECT 780.000 331.950 784.050 332.550 ;
        RECT 736.950 261.450 739.050 262.050 ;
        RECT 736.950 260.550 744.450 261.450 ;
        RECT 736.950 259.950 739.050 260.550 ;
        RECT 743.550 256.050 744.450 260.550 ;
        RECT 743.550 254.550 748.050 256.050 ;
        RECT 744.000 253.950 748.050 254.550 ;
        RECT 322.950 252.450 325.050 253.050 ;
        RECT 337.950 252.450 340.050 252.750 ;
        RECT 322.950 251.550 340.050 252.450 ;
        RECT 322.950 250.950 325.050 251.550 ;
        RECT 337.950 250.650 340.050 251.550 ;
        RECT 337.950 219.450 340.050 220.050 ;
        RECT 346.950 219.450 349.050 220.050 ;
        RECT 337.950 218.550 349.050 219.450 ;
        RECT 337.950 217.950 340.050 218.550 ;
        RECT 346.950 217.950 349.050 218.550 ;
      LAYER metal2 ;
        RECT 793.950 376.950 796.050 379.050 ;
        RECT 794.400 367.050 795.450 376.950 ;
        RECT 784.950 364.950 787.050 367.050 ;
        RECT 793.950 364.950 796.050 367.050 ;
        RECT 874.950 364.950 877.050 367.050 ;
        RECT 785.400 348.450 786.450 364.950 ;
        RECT 875.400 349.050 876.450 364.950 ;
        RECT 782.400 347.400 786.450 348.450 ;
        RECT 782.400 340.050 783.450 347.400 ;
        RECT 874.950 346.950 877.050 349.050 ;
        RECT 781.950 337.950 784.050 340.050 ;
        RECT 686.400 332.400 687.600 334.650 ;
        RECT 686.400 330.450 687.450 332.400 ;
        RECT 781.950 331.950 784.050 334.050 ;
        RECT 785.400 332.400 786.600 334.650 ;
        RECT 683.400 330.000 687.450 330.450 ;
        RECT 683.400 329.400 688.050 330.000 ;
        RECT 577.950 313.950 580.050 316.050 ;
        RECT 403.950 304.950 406.050 307.050 ;
        RECT 322.950 301.950 325.050 304.050 ;
        RECT 323.400 262.200 324.450 301.950 ;
        RECT 328.950 301.800 331.050 303.900 ;
        RECT 329.400 294.600 330.450 301.800 ;
        RECT 329.400 292.350 330.600 294.600 ;
        RECT 404.400 292.050 405.450 304.950 ;
        RECT 403.950 289.950 406.050 292.050 ;
        RECT 439.950 289.950 442.050 292.050 ;
        RECT 440.400 265.050 441.450 289.950 ;
        RECT 572.400 287.400 573.600 289.650 ;
        RECT 572.400 268.050 573.450 287.400 ;
        RECT 578.400 268.050 579.450 313.950 ;
        RECT 683.400 313.050 684.450 329.400 ;
        RECT 685.950 325.950 688.050 329.400 ;
        RECT 727.950 325.950 730.050 328.050 ;
        RECT 748.950 325.950 751.050 328.050 ;
        RECT 782.400 327.450 783.450 331.950 ;
        RECT 785.400 328.050 786.450 332.400 ;
        RECT 784.950 327.450 787.050 328.050 ;
        RECT 782.400 326.400 787.050 327.450 ;
        RECT 784.950 325.950 787.050 326.400 ;
        RECT 682.950 310.950 685.050 313.050 ;
        RECT 728.400 301.050 729.450 325.950 ;
        RECT 749.400 301.050 750.450 325.950 ;
        RECT 727.950 298.950 730.050 301.050 ;
        RECT 736.950 298.950 739.050 301.050 ;
        RECT 748.950 298.950 751.050 301.050 ;
        RECT 511.950 265.950 514.050 268.050 ;
        RECT 550.950 265.950 553.050 268.050 ;
        RECT 571.950 265.950 574.050 268.050 ;
        RECT 577.950 265.950 580.050 268.050 ;
        RECT 439.950 262.950 442.050 265.050 ;
        RECT 316.950 260.100 319.050 262.200 ;
        RECT 322.950 260.100 325.050 262.200 ;
        RECT 512.400 261.600 513.450 265.950 ;
        RECT 551.400 262.050 552.450 265.950 ;
        RECT 737.400 262.050 738.450 298.950 ;
        RECT 317.400 259.350 318.600 260.100 ;
        RECT 323.400 253.050 324.450 260.100 ;
        RECT 512.400 259.350 513.600 261.600 ;
        RECT 550.950 259.950 553.050 262.050 ;
        RECT 736.950 259.950 739.050 262.050 ;
        RECT 554.400 255.900 555.600 256.650 ;
        RECT 553.950 253.800 556.050 255.900 ;
        RECT 745.950 253.950 748.050 256.050 ;
        RECT 322.950 250.950 325.050 253.050 ;
        RECT 337.950 250.650 340.050 252.750 ;
        RECT 338.400 220.050 339.450 250.650 ;
        RECT 554.400 244.050 555.450 253.800 ;
        RECT 553.950 241.950 556.050 244.050 ;
        RECT 574.950 241.950 577.050 244.050 ;
        RECT 575.400 238.050 576.450 241.950 ;
        RECT 574.950 235.950 577.050 238.050 ;
        RECT 586.950 235.950 589.050 238.050 ;
        RECT 337.950 217.950 340.050 220.050 ;
        RECT 346.950 216.000 349.050 220.050 ;
        RECT 587.400 216.600 588.450 235.950 ;
        RECT 746.400 229.050 747.450 253.950 ;
        RECT 745.950 226.950 748.050 229.050 ;
        RECT 751.950 226.950 754.050 229.050 ;
        RECT 752.400 223.050 753.450 226.950 ;
        RECT 751.950 220.950 754.050 223.050 ;
        RECT 347.400 214.350 348.600 216.000 ;
        RECT 587.400 214.350 588.600 216.600 ;
        RECT 776.400 210.900 777.600 211.650 ;
        RECT 775.950 208.800 778.050 210.900 ;
      LAYER metal3 ;
        RECT 793.950 378.600 796.050 379.050 ;
        RECT 793.950 377.400 849.600 378.600 ;
        RECT 793.950 376.950 796.050 377.400 ;
        RECT 848.400 375.600 849.600 377.400 ;
        RECT 848.400 374.400 870.600 375.600 ;
        RECT 869.400 369.600 870.600 374.400 ;
        RECT 869.400 368.400 873.600 369.600 ;
        RECT 872.400 367.050 873.600 368.400 ;
        RECT 872.400 365.400 877.050 367.050 ;
        RECT 873.000 364.950 877.050 365.400 ;
        RECT 874.950 348.600 877.050 349.050 ;
        RECT 874.950 347.400 882.600 348.600 ;
        RECT 874.950 346.950 877.050 347.400 ;
        RECT 881.400 344.400 882.600 347.400 ;
        RECT 685.950 327.600 688.050 328.050 ;
        RECT 727.950 327.600 730.050 328.050 ;
        RECT 685.950 326.400 730.050 327.600 ;
        RECT 685.950 325.950 688.050 326.400 ;
        RECT 727.950 325.950 730.050 326.400 ;
        RECT 748.950 327.600 751.050 328.050 ;
        RECT 784.950 327.600 787.050 328.050 ;
        RECT 748.950 326.400 787.050 327.600 ;
        RECT 748.950 325.950 751.050 326.400 ;
        RECT 784.950 325.950 787.050 326.400 ;
        RECT 577.950 315.600 580.050 316.050 ;
        RECT 577.950 314.400 669.600 315.600 ;
        RECT 577.950 313.950 580.050 314.400 ;
        RECT 668.400 312.600 669.600 314.400 ;
        RECT 682.950 312.600 685.050 313.050 ;
        RECT 668.400 311.400 685.050 312.600 ;
        RECT 682.950 310.950 685.050 311.400 ;
        RECT 403.950 306.600 406.050 307.050 ;
        RECT 371.400 305.400 406.050 306.600 ;
        RECT 322.950 303.600 325.050 304.050 ;
        RECT 328.950 303.600 331.050 303.900 ;
        RECT 371.400 303.600 372.600 305.400 ;
        RECT 403.950 304.950 406.050 305.400 ;
        RECT 322.950 302.400 372.600 303.600 ;
        RECT 322.950 301.950 325.050 302.400 ;
        RECT 328.950 301.800 331.050 302.400 ;
        RECT 727.950 300.600 730.050 301.050 ;
        RECT 736.950 300.600 739.050 301.050 ;
        RECT 748.950 300.600 751.050 301.050 ;
        RECT 727.950 299.400 751.050 300.600 ;
        RECT 727.950 298.950 730.050 299.400 ;
        RECT 736.950 298.950 739.050 299.400 ;
        RECT 748.950 298.950 751.050 299.400 ;
        RECT 403.950 291.600 406.050 292.050 ;
        RECT 439.950 291.600 442.050 292.050 ;
        RECT 403.950 290.400 442.050 291.600 ;
        RECT 403.950 289.950 406.050 290.400 ;
        RECT 439.950 289.950 442.050 290.400 ;
        RECT 511.950 267.600 514.050 268.050 ;
        RECT 550.950 267.600 553.050 268.050 ;
        RECT 571.950 267.600 574.050 268.050 ;
        RECT 577.950 267.600 580.050 268.050 ;
        RECT 443.400 266.400 492.600 267.600 ;
        RECT 443.400 265.050 444.600 266.400 ;
        RECT 439.950 263.400 444.600 265.050 ;
        RECT 491.400 264.600 492.600 266.400 ;
        RECT 511.950 266.400 580.050 267.600 ;
        RECT 511.950 265.950 514.050 266.400 ;
        RECT 550.950 265.950 553.050 266.400 ;
        RECT 571.950 265.950 574.050 266.400 ;
        RECT 577.950 265.950 580.050 266.400 ;
        RECT 512.400 264.600 513.600 265.950 ;
        RECT 491.400 263.400 513.600 264.600 ;
        RECT 439.950 262.950 444.000 263.400 ;
        RECT 316.950 261.750 319.050 262.200 ;
        RECT 322.950 261.750 325.050 262.200 ;
        RECT 316.950 260.550 325.050 261.750 ;
        RECT 316.950 260.100 319.050 260.550 ;
        RECT 322.950 260.100 325.050 260.550 ;
        RECT 550.950 261.600 555.000 262.050 ;
        RECT 550.950 259.950 555.600 261.600 ;
        RECT 554.400 255.900 555.600 259.950 ;
        RECT 553.950 253.800 556.050 255.900 ;
        RECT 553.950 243.600 556.050 244.050 ;
        RECT 574.950 243.600 577.050 244.050 ;
        RECT 553.950 242.400 577.050 243.600 ;
        RECT 553.950 241.950 556.050 242.400 ;
        RECT 574.950 241.950 577.050 242.400 ;
        RECT 574.950 237.600 577.050 238.050 ;
        RECT 586.950 237.600 589.050 238.050 ;
        RECT 574.950 236.400 589.050 237.600 ;
        RECT 574.950 235.950 577.050 236.400 ;
        RECT 586.950 235.950 589.050 236.400 ;
        RECT 745.950 228.600 748.050 229.050 ;
        RECT 751.950 228.600 754.050 229.050 ;
        RECT 745.950 227.400 754.050 228.600 ;
        RECT 745.950 226.950 748.050 227.400 ;
        RECT 751.950 226.950 754.050 227.400 ;
        RECT 751.950 222.600 754.050 223.050 ;
        RECT 751.950 221.400 768.600 222.600 ;
        RECT 751.950 220.950 754.050 221.400 ;
        RECT 767.400 219.600 768.600 221.400 ;
        RECT 767.400 218.400 777.600 219.600 ;
        RECT 776.400 210.900 777.600 218.400 ;
        RECT 775.950 208.800 778.050 210.900 ;
    END
  END Cin[3]
  PIN Cin[2]
    PORT
      LAYER metal1 ;
        RECT 235.950 297.450 238.050 298.050 ;
        RECT 241.950 297.450 244.050 298.050 ;
        RECT 235.950 296.550 244.050 297.450 ;
        RECT 235.950 295.950 238.050 296.550 ;
        RECT 241.950 295.950 244.050 296.550 ;
        RECT 679.950 219.450 682.050 220.050 ;
        RECT 671.550 218.550 682.050 219.450 ;
        RECT 671.550 217.050 672.450 218.550 ;
        RECT 679.950 217.950 682.050 218.550 ;
        RECT 670.950 216.450 675.000 217.050 ;
        RECT 670.950 214.950 675.450 216.450 ;
        RECT 674.550 211.050 675.450 214.950 ;
        RECT 670.950 209.550 675.450 211.050 ;
        RECT 670.950 208.950 675.000 209.550 ;
        RECT 241.950 174.450 244.050 175.050 ;
        RECT 250.950 174.450 253.050 175.050 ;
        RECT 241.950 173.550 253.050 174.450 ;
        RECT 241.950 172.950 244.050 173.550 ;
        RECT 250.950 172.950 253.050 173.550 ;
        RECT 226.950 144.450 229.050 145.050 ;
        RECT 241.950 144.450 244.050 145.050 ;
        RECT 226.950 143.550 244.050 144.450 ;
        RECT 226.950 142.950 229.050 143.550 ;
        RECT 241.950 142.950 244.050 143.550 ;
        RECT 226.950 105.450 231.000 106.050 ;
        RECT 465.000 105.450 469.050 106.050 ;
        RECT 226.950 103.950 231.450 105.450 ;
        RECT 230.550 100.050 231.450 103.950 ;
        RECT 226.950 98.550 231.450 100.050 ;
        RECT 464.550 103.950 469.050 105.450 ;
        RECT 464.550 100.050 465.450 103.950 ;
        RECT 464.550 98.550 469.050 100.050 ;
        RECT 226.950 97.950 231.000 98.550 ;
        RECT 465.000 97.950 469.050 98.550 ;
      LAYER metal2 ;
        RECT 235.950 294.000 238.050 298.050 ;
        RECT 241.950 295.950 244.050 298.050 ;
        RECT 236.400 292.350 237.600 294.000 ;
        RECT 242.400 283.050 243.450 295.950 ;
        RECT 229.950 280.950 232.050 283.050 ;
        RECT 241.950 280.950 244.050 283.050 ;
        RECT 230.400 255.450 231.450 280.950 ;
        RECT 695.400 255.900 696.600 256.650 ;
        RECT 227.400 254.400 231.450 255.450 ;
        RECT 227.400 217.200 228.450 254.400 ;
        RECT 679.950 253.800 682.050 255.900 ;
        RECT 694.950 253.800 697.050 255.900 ;
        RECT 680.400 220.050 681.450 253.800 ;
        RECT 679.950 217.950 682.050 220.050 ;
        RECT 220.950 215.100 223.050 217.200 ;
        RECT 226.950 215.100 229.050 217.200 ;
        RECT 669.000 216.600 673.050 217.050 ;
        RECT 221.400 190.050 222.450 215.100 ;
        RECT 227.400 214.350 228.600 215.100 ;
        RECT 668.400 214.950 673.050 216.600 ;
        RECT 668.400 214.350 669.600 214.950 ;
        RECT 670.950 208.950 673.050 211.050 ;
        RECT 671.400 196.050 672.450 208.950 ;
        RECT 637.950 193.950 640.050 196.050 ;
        RECT 670.950 193.950 673.050 196.050 ;
        RECT 220.950 187.950 223.050 190.050 ;
        RECT 250.950 187.950 253.050 190.050 ;
        RECT 242.400 176.400 243.600 178.650 ;
        RECT 242.400 175.050 243.450 176.400 ;
        RECT 251.400 175.050 252.450 187.950 ;
        RECT 638.400 175.050 639.450 193.950 ;
        RECT 241.950 172.950 244.050 175.050 ;
        RECT 250.950 172.950 253.050 175.050 ;
        RECT 628.950 172.950 631.050 175.050 ;
        RECT 637.950 172.950 640.050 175.050 ;
        RECT 208.950 157.950 211.050 160.050 ;
        RECT 226.800 157.950 228.900 160.050 ;
        RECT 209.400 139.200 210.450 157.950 ;
        RECT 227.400 145.050 228.450 157.950 ;
        RECT 242.400 145.050 243.450 172.950 ;
        RECT 629.400 157.050 630.450 172.950 ;
        RECT 601.950 154.950 604.050 157.050 ;
        RECT 628.950 154.950 631.050 157.050 ;
        RECT 226.950 142.950 229.050 145.050 ;
        RECT 241.950 142.950 244.050 145.050 ;
        RECT 602.400 139.200 603.450 154.950 ;
        RECT 208.950 137.100 211.050 139.200 ;
        RECT 601.950 137.100 604.050 139.200 ;
        RECT 209.400 136.350 210.600 137.100 ;
        RECT 602.400 136.350 603.600 137.100 ;
        RECT 211.950 130.950 214.050 133.050 ;
        RECT 491.400 131.400 492.600 133.650 ;
        RECT 212.400 124.050 213.450 130.950 ;
        RECT 211.950 121.950 214.050 124.050 ;
        RECT 226.950 121.950 229.050 124.050 ;
        RECT 227.400 106.050 228.450 121.950 ;
        RECT 491.400 121.050 492.450 131.400 ;
        RECT 592.950 130.950 595.050 133.050 ;
        RECT 593.400 127.050 594.450 130.950 ;
        RECT 577.950 124.950 580.050 127.050 ;
        RECT 592.950 124.950 595.050 127.050 ;
        RECT 490.950 118.950 493.050 121.050 ;
        RECT 541.950 118.950 544.050 121.050 ;
        RECT 491.400 115.050 492.450 118.950 ;
        RECT 466.950 112.950 469.050 115.050 ;
        RECT 490.950 112.950 493.050 115.050 ;
        RECT 467.400 106.050 468.450 112.950 ;
        RECT 542.400 106.050 543.450 118.950 ;
        RECT 578.400 106.050 579.450 124.950 ;
        RECT 226.950 103.950 229.050 106.050 ;
        RECT 466.950 103.950 469.050 106.050 ;
        RECT 541.950 103.950 544.050 106.050 ;
        RECT 577.950 103.950 580.050 106.050 ;
        RECT 226.950 97.950 229.050 100.050 ;
        RECT 466.950 97.950 469.050 100.050 ;
        RECT 575.400 99.900 576.600 100.650 ;
        RECT 227.400 85.050 228.450 97.950 ;
        RECT 280.950 88.950 283.050 91.050 ;
        RECT 355.950 90.450 358.050 90.900 ;
        RECT 361.950 90.450 364.050 94.050 ;
        RECT 367.950 91.950 370.050 94.050 ;
        RECT 355.950 90.000 364.050 90.450 ;
        RECT 355.950 89.400 363.450 90.000 ;
        RECT 281.400 85.050 282.450 88.950 ;
        RECT 355.950 88.800 358.050 89.400 ;
        RECT 368.400 88.050 369.450 91.950 ;
        RECT 367.950 85.950 370.050 88.050 ;
        RECT 451.950 85.800 454.050 87.900 ;
        RECT 226.950 82.950 229.050 85.050 ;
        RECT 280.950 82.950 283.050 85.050 ;
        RECT 452.400 76.050 453.450 85.800 ;
        RECT 467.400 76.050 468.450 97.950 ;
        RECT 574.950 97.800 577.050 99.900 ;
        RECT 451.950 73.950 454.050 76.050 ;
        RECT 466.950 73.950 469.050 76.050 ;
        RECT 575.400 70.050 576.450 97.800 ;
        RECT 574.950 67.950 577.050 70.050 ;
        RECT 583.950 67.950 586.050 70.050 ;
        RECT 584.400 46.050 585.450 67.950 ;
        RECT 571.950 43.950 574.050 46.050 ;
        RECT 583.950 43.950 586.050 46.050 ;
        RECT 572.400 -2.550 573.450 43.950 ;
        RECT 572.400 -3.600 576.450 -2.550 ;
      LAYER metal3 ;
        RECT 229.950 282.600 232.050 283.050 ;
        RECT 241.950 282.600 244.050 283.050 ;
        RECT 229.950 281.400 244.050 282.600 ;
        RECT 229.950 280.950 232.050 281.400 ;
        RECT 241.950 280.950 244.050 281.400 ;
        RECT 679.950 255.450 682.050 255.900 ;
        RECT 694.950 255.450 697.050 255.900 ;
        RECT 679.950 254.250 697.050 255.450 ;
        RECT 679.950 253.800 682.050 254.250 ;
        RECT 694.950 253.800 697.050 254.250 ;
        RECT 220.950 216.750 223.050 217.200 ;
        RECT 226.950 216.750 229.050 217.200 ;
        RECT 220.950 215.550 229.050 216.750 ;
        RECT 220.950 215.100 223.050 215.550 ;
        RECT 226.950 215.100 229.050 215.550 ;
        RECT 637.950 195.600 640.050 196.050 ;
        RECT 670.950 195.600 673.050 196.050 ;
        RECT 637.950 194.400 673.050 195.600 ;
        RECT 637.950 193.950 640.050 194.400 ;
        RECT 670.950 193.950 673.050 194.400 ;
        RECT 220.950 189.600 223.050 190.050 ;
        RECT 250.950 189.600 253.050 190.050 ;
        RECT 220.950 188.400 253.050 189.600 ;
        RECT 220.950 187.950 223.050 188.400 ;
        RECT 250.950 187.950 253.050 188.400 ;
        RECT 628.950 174.600 631.050 175.050 ;
        RECT 637.950 174.600 640.050 175.050 ;
        RECT 628.950 173.400 640.050 174.600 ;
        RECT 628.950 172.950 631.050 173.400 ;
        RECT 637.950 172.950 640.050 173.400 ;
        RECT 208.950 159.600 211.050 160.050 ;
        RECT 226.800 159.600 228.900 160.050 ;
        RECT 208.950 158.400 228.900 159.600 ;
        RECT 208.950 157.950 211.050 158.400 ;
        RECT 226.800 157.950 228.900 158.400 ;
        RECT 601.950 156.600 604.050 157.050 ;
        RECT 628.950 156.600 631.050 157.050 ;
        RECT 601.950 155.400 631.050 156.600 ;
        RECT 601.950 154.950 604.050 155.400 ;
        RECT 628.950 154.950 631.050 155.400 ;
        RECT 208.950 137.100 211.050 139.200 ;
        RECT 601.950 137.100 604.050 139.200 ;
        RECT 209.400 133.050 210.600 137.100 ;
        RECT 602.400 135.600 603.600 137.100 ;
        RECT 596.400 134.400 603.600 135.600 ;
        RECT 596.400 133.050 597.600 134.400 ;
        RECT 209.400 131.400 214.050 133.050 ;
        RECT 210.000 130.950 214.050 131.400 ;
        RECT 592.950 131.400 597.600 133.050 ;
        RECT 592.950 130.950 597.000 131.400 ;
        RECT 577.950 126.600 580.050 127.050 ;
        RECT 592.950 126.600 595.050 127.050 ;
        RECT 577.950 125.400 595.050 126.600 ;
        RECT 577.950 124.950 580.050 125.400 ;
        RECT 592.950 124.950 595.050 125.400 ;
        RECT 211.950 123.600 214.050 124.050 ;
        RECT 226.950 123.600 229.050 124.050 ;
        RECT 211.950 122.400 229.050 123.600 ;
        RECT 211.950 121.950 214.050 122.400 ;
        RECT 226.950 121.950 229.050 122.400 ;
        RECT 490.950 120.600 493.050 121.050 ;
        RECT 541.950 120.600 544.050 121.050 ;
        RECT 490.950 119.400 544.050 120.600 ;
        RECT 490.950 118.950 493.050 119.400 ;
        RECT 541.950 118.950 544.050 119.400 ;
        RECT 466.950 114.600 469.050 115.050 ;
        RECT 490.950 114.600 493.050 115.050 ;
        RECT 466.950 113.400 493.050 114.600 ;
        RECT 466.950 112.950 469.050 113.400 ;
        RECT 490.950 112.950 493.050 113.400 ;
        RECT 541.950 105.600 544.050 106.050 ;
        RECT 576.000 105.600 580.050 106.050 ;
        RECT 541.950 104.400 580.050 105.600 ;
        RECT 541.950 103.950 544.050 104.400 ;
        RECT 575.400 103.950 580.050 104.400 ;
        RECT 575.400 99.900 576.600 103.950 ;
        RECT 574.950 97.800 577.050 99.900 ;
        RECT 361.950 93.600 364.050 94.050 ;
        RECT 367.950 93.600 370.050 94.050 ;
        RECT 361.950 92.400 370.050 93.600 ;
        RECT 361.950 91.950 364.050 92.400 ;
        RECT 367.950 91.950 370.050 92.400 ;
        RECT 280.950 90.600 283.050 91.050 ;
        RECT 355.950 90.600 358.050 90.900 ;
        RECT 280.950 89.400 358.050 90.600 ;
        RECT 280.950 88.950 283.050 89.400 ;
        RECT 355.950 88.800 358.050 89.400 ;
        RECT 367.950 87.600 370.050 88.050 ;
        RECT 451.950 87.600 454.050 87.900 ;
        RECT 367.950 86.400 454.050 87.600 ;
        RECT 367.950 85.950 370.050 86.400 ;
        RECT 451.950 85.800 454.050 86.400 ;
        RECT 226.950 84.600 229.050 85.050 ;
        RECT 280.950 84.600 283.050 85.050 ;
        RECT 226.950 83.400 283.050 84.600 ;
        RECT 226.950 82.950 229.050 83.400 ;
        RECT 280.950 82.950 283.050 83.400 ;
        RECT 451.950 75.600 454.050 76.050 ;
        RECT 466.950 75.600 469.050 76.050 ;
        RECT 451.950 74.400 469.050 75.600 ;
        RECT 451.950 73.950 454.050 74.400 ;
        RECT 466.950 73.950 469.050 74.400 ;
        RECT 574.950 69.600 577.050 70.050 ;
        RECT 583.950 69.600 586.050 70.050 ;
        RECT 574.950 68.400 586.050 69.600 ;
        RECT 574.950 67.950 577.050 68.400 ;
        RECT 583.950 67.950 586.050 68.400 ;
        RECT 571.950 45.600 574.050 46.050 ;
        RECT 583.950 45.600 586.050 46.050 ;
        RECT 571.950 44.400 586.050 45.600 ;
        RECT 571.950 43.950 574.050 44.400 ;
        RECT 583.950 43.950 586.050 44.400 ;
    END
  END Cin[2]
  PIN Cin[1]
    PORT
      LAYER metal1 ;
        RECT 415.950 105.450 420.000 106.050 ;
        RECT 415.950 103.950 420.450 105.450 ;
        RECT 419.550 100.050 420.450 103.950 ;
        RECT 419.550 98.550 424.050 100.050 ;
        RECT 420.000 97.950 424.050 98.550 ;
      LAYER metal2 ;
        RECT 439.950 244.800 442.050 246.900 ;
        RECT 466.950 244.950 469.050 247.050 ;
        RECT 403.950 238.950 406.050 241.050 ;
        RECT 293.400 209.400 294.600 211.650 ;
        RECT 404.400 210.450 405.450 238.950 ;
        RECT 440.400 238.050 441.450 244.800 ;
        RECT 467.400 238.050 468.450 244.950 ;
        RECT 439.950 235.950 442.050 238.050 ;
        RECT 466.950 235.950 469.050 238.050 ;
        RECT 538.950 235.950 541.050 238.050 ;
        RECT 539.400 210.900 540.450 235.950 ;
        RECT 548.400 210.900 549.600 211.650 ;
        RECT 401.400 209.400 405.450 210.450 ;
        RECT 293.400 205.050 294.450 209.400 ;
        RECT 292.950 202.950 295.050 205.050 ;
        RECT 370.950 202.950 373.050 205.050 ;
        RECT 293.400 196.050 294.450 202.950 ;
        RECT 262.950 193.950 265.050 196.050 ;
        RECT 292.950 193.950 295.050 196.050 ;
        RECT 263.400 183.600 264.450 193.950 ;
        RECT 371.400 190.050 372.450 202.950 ;
        RECT 401.400 193.050 402.450 209.400 ;
        RECT 538.950 208.800 541.050 210.900 ;
        RECT 547.950 208.800 550.050 210.900 ;
        RECT 400.800 190.950 402.900 193.050 ;
        RECT 370.950 187.950 373.050 190.050 ;
        RECT 401.400 183.600 402.450 190.950 ;
        RECT 263.400 181.350 264.600 183.600 ;
        RECT 401.400 183.450 402.600 183.600 ;
        RECT 398.400 182.400 402.600 183.450 ;
        RECT 398.400 141.450 399.450 182.400 ;
        RECT 401.400 181.350 402.600 182.400 ;
        RECT 398.400 140.400 402.450 141.450 ;
        RECT 401.400 133.050 402.450 140.400 ;
        RECT 400.950 130.950 403.050 133.050 ;
        RECT 415.950 130.950 418.050 133.050 ;
        RECT 416.400 106.050 417.450 130.950 ;
        RECT 415.950 103.950 418.050 106.050 ;
        RECT 421.950 97.950 424.050 100.050 ;
        RECT 422.400 73.050 423.450 97.950 ;
        RECT 421.950 70.950 424.050 73.050 ;
        RECT 448.950 70.950 451.050 73.050 ;
        RECT 449.400 4.050 450.450 70.950 ;
        RECT 403.950 1.950 406.050 4.050 ;
        RECT 448.950 1.950 451.050 4.050 ;
        RECT 404.400 -3.600 405.450 1.950 ;
      LAYER metal3 ;
        RECT 439.950 246.600 442.050 246.900 ;
        RECT 466.950 246.600 469.050 247.050 ;
        RECT 439.950 245.400 469.050 246.600 ;
        RECT 439.950 244.800 442.050 245.400 ;
        RECT 466.950 244.950 469.050 245.400 ;
        RECT 403.950 240.600 406.050 241.050 ;
        RECT 403.950 239.400 420.600 240.600 ;
        RECT 403.950 238.950 406.050 239.400 ;
        RECT 419.400 237.600 420.600 239.400 ;
        RECT 439.950 237.600 442.050 238.050 ;
        RECT 419.400 236.400 442.050 237.600 ;
        RECT 439.950 235.950 442.050 236.400 ;
        RECT 466.950 237.600 469.050 238.050 ;
        RECT 538.950 237.600 541.050 238.050 ;
        RECT 466.950 236.400 541.050 237.600 ;
        RECT 466.950 235.950 469.050 236.400 ;
        RECT 538.950 235.950 541.050 236.400 ;
        RECT 538.950 210.450 541.050 210.900 ;
        RECT 547.950 210.450 550.050 210.900 ;
        RECT 538.950 209.250 550.050 210.450 ;
        RECT 538.950 208.800 541.050 209.250 ;
        RECT 547.950 208.800 550.050 209.250 ;
        RECT 292.950 204.600 295.050 205.050 ;
        RECT 370.950 204.600 373.050 205.050 ;
        RECT 292.950 203.400 373.050 204.600 ;
        RECT 292.950 202.950 295.050 203.400 ;
        RECT 370.950 202.950 373.050 203.400 ;
        RECT 262.950 195.600 265.050 196.050 ;
        RECT 292.950 195.600 295.050 196.050 ;
        RECT 262.950 194.400 295.050 195.600 ;
        RECT 262.950 193.950 265.050 194.400 ;
        RECT 292.950 193.950 295.050 194.400 ;
        RECT 400.800 192.600 402.900 193.050 ;
        RECT 389.400 191.400 402.900 192.600 ;
        RECT 370.950 189.600 373.050 190.050 ;
        RECT 389.400 189.600 390.600 191.400 ;
        RECT 400.800 190.950 402.900 191.400 ;
        RECT 370.950 188.400 390.600 189.600 ;
        RECT 370.950 187.950 373.050 188.400 ;
        RECT 400.950 132.600 403.050 133.050 ;
        RECT 415.950 132.600 418.050 133.050 ;
        RECT 400.950 131.400 418.050 132.600 ;
        RECT 400.950 130.950 403.050 131.400 ;
        RECT 415.950 130.950 418.050 131.400 ;
        RECT 421.950 72.600 424.050 73.050 ;
        RECT 448.950 72.600 451.050 73.050 ;
        RECT 421.950 71.400 451.050 72.600 ;
        RECT 421.950 70.950 424.050 71.400 ;
        RECT 448.950 70.950 451.050 71.400 ;
        RECT 403.950 3.600 406.050 4.050 ;
        RECT 448.950 3.600 451.050 4.050 ;
        RECT 403.950 2.400 451.050 3.600 ;
        RECT 403.950 1.950 406.050 2.400 ;
        RECT 448.950 1.950 451.050 2.400 ;
    END
  END Cin[1]
  PIN Cin[0]
    PORT
      LAYER metal2 ;
        RECT 317.400 287.400 318.600 289.650 ;
        RECT 317.400 271.050 318.450 287.400 ;
        RECT 277.950 268.950 280.050 271.050 ;
        RECT 304.950 268.950 307.050 271.050 ;
        RECT 316.950 268.950 319.050 271.050 ;
        RECT 278.400 261.600 279.450 268.950 ;
        RECT 278.400 259.350 279.600 261.600 ;
        RECT 305.400 229.050 306.450 268.950 ;
        RECT 304.950 226.950 307.050 229.050 ;
        RECT 361.950 226.950 364.050 229.050 ;
        RECT 362.400 199.050 363.450 226.950 ;
        RECT 361.950 196.950 364.050 199.050 ;
        RECT 376.950 196.950 379.050 199.050 ;
        RECT 377.400 193.050 378.450 196.950 ;
        RECT 418.950 193.950 421.050 196.050 ;
        RECT 376.950 190.950 379.050 193.050 ;
        RECT 419.400 183.600 420.450 193.950 ;
        RECT 419.400 183.450 420.600 183.600 ;
        RECT 416.400 182.400 420.600 183.450 ;
        RECT 416.400 138.450 417.450 182.400 ;
        RECT 419.400 181.350 420.600 182.400 ;
        RECT 416.400 137.400 420.450 138.450 ;
        RECT 398.400 131.400 399.600 133.650 ;
        RECT 398.400 127.050 399.450 131.400 ;
        RECT 419.400 127.050 420.450 137.400 ;
        RECT 397.950 124.950 400.050 127.050 ;
        RECT 418.950 124.950 421.050 127.050 ;
        RECT 419.400 117.450 420.450 124.950 ;
        RECT 419.400 116.400 423.450 117.450 ;
        RECT 422.400 106.050 423.450 116.400 ;
        RECT 421.950 103.950 424.050 106.050 ;
        RECT 415.950 97.950 418.050 100.050 ;
        RECT 416.400 73.050 417.450 97.950 ;
        RECT 406.950 70.800 409.050 72.900 ;
        RECT 415.950 70.950 418.050 73.050 ;
        RECT 407.400 52.050 408.450 70.800 ;
        RECT 400.950 49.950 403.050 52.050 ;
        RECT 406.950 49.950 409.050 52.050 ;
        RECT 401.400 45.450 402.450 49.950 ;
        RECT 398.400 44.400 402.450 45.450 ;
        RECT 398.400 31.050 399.450 44.400 ;
        RECT 397.950 28.950 400.050 31.050 ;
        RECT 409.950 19.950 412.050 22.050 ;
        RECT 410.400 7.050 411.450 19.950 ;
        RECT 400.950 4.950 403.050 7.050 ;
        RECT 409.800 4.950 411.900 7.050 ;
        RECT 401.400 -2.550 402.450 4.950 ;
        RECT 398.400 -3.600 402.450 -2.550 ;
      LAYER metal3 ;
        RECT 277.950 270.600 280.050 271.050 ;
        RECT 304.950 270.600 307.050 271.050 ;
        RECT 316.950 270.600 319.050 271.050 ;
        RECT 277.950 269.400 319.050 270.600 ;
        RECT 277.950 268.950 280.050 269.400 ;
        RECT 304.950 268.950 307.050 269.400 ;
        RECT 316.950 268.950 319.050 269.400 ;
        RECT 304.950 228.600 307.050 229.050 ;
        RECT 361.950 228.600 364.050 229.050 ;
        RECT 304.950 227.400 364.050 228.600 ;
        RECT 304.950 226.950 307.050 227.400 ;
        RECT 361.950 226.950 364.050 227.400 ;
        RECT 361.950 198.600 364.050 199.050 ;
        RECT 376.950 198.600 379.050 199.050 ;
        RECT 361.950 197.400 379.050 198.600 ;
        RECT 361.950 196.950 364.050 197.400 ;
        RECT 376.950 196.950 379.050 197.400 ;
        RECT 418.950 195.600 421.050 196.050 ;
        RECT 386.400 194.400 421.050 195.600 ;
        RECT 376.950 192.600 379.050 193.050 ;
        RECT 386.400 192.600 387.600 194.400 ;
        RECT 418.950 193.950 421.050 194.400 ;
        RECT 376.950 191.400 387.600 192.600 ;
        RECT 376.950 190.950 379.050 191.400 ;
        RECT 397.950 126.600 400.050 127.050 ;
        RECT 418.950 126.600 421.050 127.050 ;
        RECT 397.950 125.400 421.050 126.600 ;
        RECT 397.950 124.950 400.050 125.400 ;
        RECT 418.950 124.950 421.050 125.400 ;
        RECT 421.950 105.600 424.050 106.050 ;
        RECT 416.400 104.400 424.050 105.600 ;
        RECT 416.400 100.050 417.600 104.400 ;
        RECT 421.950 103.950 424.050 104.400 ;
        RECT 415.950 97.950 418.050 100.050 ;
        RECT 406.950 72.600 409.050 72.900 ;
        RECT 415.950 72.600 418.050 73.050 ;
        RECT 406.950 71.400 418.050 72.600 ;
        RECT 406.950 70.800 409.050 71.400 ;
        RECT 415.950 70.950 418.050 71.400 ;
        RECT 400.950 51.600 403.050 52.050 ;
        RECT 406.950 51.600 409.050 52.050 ;
        RECT 400.950 50.400 409.050 51.600 ;
        RECT 400.950 49.950 403.050 50.400 ;
        RECT 406.950 49.950 409.050 50.400 ;
        RECT 397.950 30.600 402.000 31.050 ;
        RECT 397.950 28.950 402.600 30.600 ;
        RECT 401.400 27.600 402.600 28.950 ;
        RECT 401.400 26.400 411.600 27.600 ;
        RECT 410.400 22.050 411.600 26.400 ;
        RECT 409.950 19.950 412.050 22.050 ;
        RECT 400.950 6.600 403.050 7.050 ;
        RECT 409.800 6.600 411.900 7.050 ;
        RECT 400.950 5.400 411.900 6.600 ;
        RECT 400.950 4.950 403.050 5.400 ;
        RECT 409.800 4.950 411.900 5.400 ;
    END
  END Cin[0]
  PIN Rdy
    PORT
      LAYER metal2 ;
        RECT 14.400 411.000 15.600 412.650 ;
        RECT 13.950 406.950 16.050 411.000 ;
      LAYER metal3 ;
        RECT -3.600 408.600 -2.400 411.600 ;
        RECT 13.950 408.600 16.050 409.050 ;
        RECT -3.600 407.400 16.050 408.600 ;
        RECT 13.950 406.950 16.050 407.400 ;
    END
  END Rdy
  PIN Vld
    PORT
      LAYER metal2 ;
        RECT 10.950 449.100 13.050 451.200 ;
        RECT 11.400 448.350 12.600 449.100 ;
      LAYER metal3 ;
        RECT 10.950 450.600 13.050 451.200 ;
        RECT -3.600 449.400 13.050 450.600 ;
        RECT 10.950 449.100 13.050 449.400 ;
    END
  END Vld
  PIN Xin[3]
    PORT
      LAYER metal2 ;
        RECT 661.950 391.950 664.050 394.050 ;
        RECT 874.950 391.950 877.050 394.050 ;
        RECT 662.400 385.050 663.450 391.950 ;
        RECT 556.950 382.950 559.050 385.050 ;
        RECT 661.950 382.950 664.050 385.050 ;
        RECT 557.400 373.200 558.450 382.950 ;
        RECT 544.950 371.100 547.050 373.200 ;
        RECT 556.950 371.100 559.050 373.200 ;
        RECT 875.400 373.050 876.450 391.950 ;
        RECT 545.400 370.350 546.600 371.100 ;
        RECT 557.400 370.350 558.600 371.100 ;
        RECT 874.950 370.950 877.050 373.050 ;
      LAYER metal3 ;
        RECT 661.950 393.600 664.050 394.050 ;
        RECT 874.950 393.600 877.050 394.050 ;
        RECT 661.950 392.400 877.050 393.600 ;
        RECT 661.950 391.950 664.050 392.400 ;
        RECT 874.950 391.950 877.050 392.400 ;
        RECT 556.950 384.600 559.050 385.050 ;
        RECT 661.950 384.600 664.050 385.050 ;
        RECT 556.950 383.400 664.050 384.600 ;
        RECT 556.950 382.950 559.050 383.400 ;
        RECT 661.950 382.950 664.050 383.400 ;
        RECT 544.950 372.600 547.050 373.200 ;
        RECT 556.950 372.600 559.050 373.200 ;
        RECT 544.950 371.400 559.050 372.600 ;
        RECT 544.950 371.100 547.050 371.400 ;
        RECT 556.950 371.100 559.050 371.400 ;
        RECT 874.950 372.600 877.050 373.050 ;
        RECT 874.950 371.400 882.600 372.600 ;
        RECT 874.950 370.950 877.050 371.400 ;
    END
  END Xin[3]
  PIN Xin[2]
    PORT
      LAYER metal2 ;
        RECT 629.400 410.400 630.600 412.650 ;
        RECT 629.400 391.050 630.450 410.400 ;
        RECT 871.950 403.950 874.050 406.050 ;
        RECT 872.400 400.050 873.450 403.950 ;
        RECT 862.950 397.950 865.050 400.050 ;
        RECT 871.950 397.950 874.050 400.050 ;
        RECT 863.400 391.050 864.450 397.950 ;
        RECT 568.950 388.950 571.050 391.050 ;
        RECT 628.950 388.950 631.050 391.050 ;
        RECT 862.950 388.950 865.050 391.050 ;
        RECT 569.400 340.050 570.450 388.950 ;
        RECT 568.950 337.950 571.050 340.050 ;
        RECT 566.400 333.900 567.600 334.650 ;
        RECT 565.950 331.800 568.050 333.900 ;
      LAYER metal3 ;
        RECT 871.950 405.600 874.050 406.050 ;
        RECT 881.400 405.600 882.600 411.600 ;
        RECT 871.950 404.400 882.600 405.600 ;
        RECT 871.950 403.950 874.050 404.400 ;
        RECT 862.950 399.600 865.050 400.050 ;
        RECT 871.950 399.600 874.050 400.050 ;
        RECT 862.950 398.400 874.050 399.600 ;
        RECT 862.950 397.950 865.050 398.400 ;
        RECT 871.950 397.950 874.050 398.400 ;
        RECT 568.950 390.600 571.050 391.050 ;
        RECT 628.950 390.600 631.050 391.050 ;
        RECT 862.950 390.600 865.050 391.050 ;
        RECT 568.950 389.400 865.050 390.600 ;
        RECT 568.950 388.950 571.050 389.400 ;
        RECT 628.950 388.950 631.050 389.400 ;
        RECT 862.950 388.950 865.050 389.400 ;
        RECT 568.950 337.950 571.050 340.050 ;
        RECT 565.950 333.600 568.050 333.900 ;
        RECT 569.400 333.600 570.600 337.950 ;
        RECT 565.950 332.400 570.600 333.600 ;
        RECT 565.950 331.800 568.050 332.400 ;
    END
  END Xin[2]
  PIN Xin[1]
    PORT
      LAYER metal1 ;
        RECT 363.000 294.450 367.050 295.050 ;
        RECT 362.550 292.950 367.050 294.450 ;
        RECT 362.550 289.050 363.450 292.950 ;
        RECT 358.950 287.550 363.450 289.050 ;
        RECT 358.950 286.950 363.000 287.550 ;
      LAYER metal2 ;
        RECT 373.950 385.950 376.050 388.050 ;
        RECT 469.950 385.950 472.050 388.050 ;
        RECT 374.400 358.050 375.450 385.950 ;
        RECT 470.400 379.050 471.450 385.950 ;
        RECT 469.950 376.950 472.050 379.050 ;
        RECT 496.950 376.950 499.050 379.050 ;
        RECT 497.400 372.600 498.450 376.950 ;
        RECT 497.400 370.350 498.600 372.600 ;
        RECT 373.950 355.950 376.050 358.050 ;
        RECT 385.950 355.950 388.050 358.050 ;
        RECT 386.400 340.050 387.450 355.950 ;
        RECT 385.800 337.950 387.900 340.050 ;
        RECT 383.400 333.900 384.600 334.650 ;
        RECT 382.950 331.800 385.050 333.900 ;
        RECT 383.400 328.050 384.450 331.800 ;
        RECT 364.950 325.950 367.050 328.050 ;
        RECT 382.950 325.950 385.050 328.050 ;
        RECT 365.400 295.050 366.450 325.950 ;
        RECT 364.950 292.950 367.050 295.050 ;
        RECT 358.950 286.950 361.050 289.050 ;
        RECT 359.400 267.450 360.450 286.950 ;
        RECT 356.400 267.000 360.450 267.450 ;
        RECT 355.950 266.400 360.450 267.000 ;
        RECT 349.950 262.950 352.050 265.050 ;
        RECT 355.950 262.950 358.050 266.400 ;
        RECT 350.400 220.050 351.450 262.950 ;
        RECT 340.950 217.950 343.050 220.050 ;
        RECT 349.950 217.950 352.050 220.050 ;
        RECT 341.400 189.450 342.450 217.950 ;
        RECT 338.400 188.400 342.450 189.450 ;
        RECT 338.400 142.050 339.450 188.400 ;
        RECT 337.950 139.950 340.050 142.050 ;
        RECT 352.950 127.950 355.050 130.050 ;
        RECT 353.400 105.450 354.450 127.950 ;
        RECT 353.400 104.400 357.450 105.450 ;
        RECT 356.400 94.050 357.450 104.400 ;
        RECT 340.950 91.800 343.050 93.900 ;
        RECT 355.950 91.950 358.050 94.050 ;
        RECT 341.400 61.050 342.450 91.800 ;
        RECT 340.800 58.950 342.900 61.050 ;
        RECT 325.950 52.950 328.050 55.050 ;
        RECT 326.400 28.050 327.450 52.950 ;
        RECT 325.950 25.950 328.050 28.050 ;
        RECT 355.950 16.950 358.050 19.050 ;
        RECT 356.400 7.050 357.450 16.950 ;
        RECT 355.950 4.950 358.050 7.050 ;
        RECT 379.950 4.950 382.050 7.050 ;
        RECT 380.400 -3.600 381.450 4.950 ;
      LAYER metal3 ;
        RECT 373.950 387.600 376.050 388.050 ;
        RECT 469.950 387.600 472.050 388.050 ;
        RECT 373.950 386.400 472.050 387.600 ;
        RECT 373.950 385.950 376.050 386.400 ;
        RECT 469.950 385.950 472.050 386.400 ;
        RECT 469.950 378.600 472.050 379.050 ;
        RECT 496.950 378.600 499.050 379.050 ;
        RECT 469.950 377.400 499.050 378.600 ;
        RECT 469.950 376.950 472.050 377.400 ;
        RECT 496.950 376.950 499.050 377.400 ;
        RECT 373.950 357.600 376.050 358.050 ;
        RECT 385.950 357.600 388.050 358.050 ;
        RECT 373.950 356.400 388.050 357.600 ;
        RECT 373.950 355.950 376.050 356.400 ;
        RECT 385.950 355.950 388.050 356.400 ;
        RECT 384.000 339.600 387.900 340.050 ;
        RECT 383.400 337.950 387.900 339.600 ;
        RECT 383.400 333.900 384.600 337.950 ;
        RECT 382.950 331.800 385.050 333.900 ;
        RECT 364.950 327.600 367.050 328.050 ;
        RECT 382.950 327.600 385.050 328.050 ;
        RECT 364.950 326.400 385.050 327.600 ;
        RECT 364.950 325.950 367.050 326.400 ;
        RECT 382.950 325.950 385.050 326.400 ;
        RECT 349.950 264.600 352.050 265.050 ;
        RECT 355.950 264.600 358.050 265.050 ;
        RECT 349.950 263.400 358.050 264.600 ;
        RECT 349.950 262.950 352.050 263.400 ;
        RECT 355.950 262.950 358.050 263.400 ;
        RECT 340.950 219.600 343.050 220.050 ;
        RECT 349.950 219.600 352.050 220.050 ;
        RECT 340.950 218.400 352.050 219.600 ;
        RECT 340.950 217.950 343.050 218.400 ;
        RECT 349.950 217.950 352.050 218.400 ;
        RECT 337.950 138.600 340.050 142.050 ;
        RECT 337.950 138.000 348.600 138.600 ;
        RECT 338.400 137.400 348.600 138.000 ;
        RECT 347.400 129.600 348.600 137.400 ;
        RECT 352.950 129.600 355.050 130.050 ;
        RECT 347.400 128.400 355.050 129.600 ;
        RECT 352.950 127.950 355.050 128.400 ;
        RECT 340.950 93.600 343.050 93.900 ;
        RECT 355.950 93.600 358.050 94.050 ;
        RECT 340.950 92.400 358.050 93.600 ;
        RECT 340.950 91.800 343.050 92.400 ;
        RECT 355.950 91.950 358.050 92.400 ;
        RECT 340.800 60.600 342.900 61.050 ;
        RECT 332.400 59.400 342.900 60.600 ;
        RECT 332.400 57.600 333.600 59.400 ;
        RECT 340.800 58.950 342.900 59.400 ;
        RECT 326.400 57.000 333.600 57.600 ;
        RECT 325.950 56.400 333.600 57.000 ;
        RECT 325.950 52.950 328.050 56.400 ;
        RECT 325.950 27.600 328.050 28.050 ;
        RECT 325.950 26.400 336.600 27.600 ;
        RECT 325.950 25.950 328.050 26.400 ;
        RECT 335.400 18.600 336.600 26.400 ;
        RECT 355.950 18.600 358.050 19.050 ;
        RECT 335.400 17.400 358.050 18.600 ;
        RECT 355.950 16.950 358.050 17.400 ;
        RECT 355.950 6.600 358.050 7.050 ;
        RECT 379.950 6.600 382.050 7.050 ;
        RECT 355.950 5.400 382.050 6.600 ;
        RECT 355.950 4.950 358.050 5.400 ;
        RECT 379.950 4.950 382.050 5.400 ;
    END
  END Xin[1]
  PIN Xin[0]
    PORT
      LAYER metal1 ;
        RECT 423.000 216.450 427.050 217.050 ;
        RECT 422.550 214.950 427.050 216.450 ;
        RECT 422.550 211.050 423.450 214.950 ;
        RECT 418.950 209.550 423.450 211.050 ;
        RECT 418.950 208.950 423.000 209.550 ;
        RECT 406.950 138.450 409.050 139.050 ;
        RECT 401.550 137.550 409.050 138.450 ;
        RECT 401.550 129.900 402.450 137.550 ;
        RECT 406.950 136.950 409.050 137.550 ;
        RECT 400.950 127.800 403.050 129.900 ;
        RECT 418.950 63.450 421.050 64.050 ;
        RECT 418.950 62.550 429.450 63.450 ;
        RECT 418.950 61.950 421.050 62.550 ;
        RECT 428.550 55.050 429.450 62.550 ;
        RECT 424.950 53.550 429.450 55.050 ;
        RECT 424.950 52.950 429.000 53.550 ;
      LAYER metal2 ;
        RECT 409.950 371.100 412.050 373.200 ;
        RECT 410.400 370.350 411.600 371.100 ;
        RECT 415.950 370.950 418.050 373.050 ;
        RECT 421.950 371.100 424.050 373.200 ;
        RECT 416.400 346.050 417.450 370.950 ;
        RECT 422.400 370.350 423.600 371.100 ;
        RECT 415.950 343.950 418.050 346.050 ;
        RECT 424.950 343.950 427.050 346.050 ;
        RECT 425.400 217.050 426.450 343.950 ;
        RECT 424.950 214.950 427.050 217.050 ;
        RECT 418.950 208.950 421.050 211.050 ;
        RECT 419.400 202.050 420.450 208.950 ;
        RECT 412.950 199.800 415.050 201.900 ;
        RECT 418.950 199.950 421.050 202.050 ;
        RECT 413.400 142.050 414.450 199.800 ;
        RECT 406.950 136.950 409.050 142.050 ;
        RECT 412.950 139.950 415.050 142.050 ;
        RECT 400.950 127.800 403.050 129.900 ;
        RECT 401.400 106.050 402.450 127.800 ;
        RECT 400.950 103.950 403.050 106.050 ;
        RECT 400.950 97.950 403.050 100.050 ;
        RECT 401.400 67.050 402.450 97.950 ;
        RECT 400.950 64.950 403.050 67.050 ;
        RECT 418.950 61.950 421.050 67.050 ;
        RECT 424.950 52.950 427.050 55.050 ;
        RECT 425.400 27.450 426.450 52.950 ;
        RECT 425.400 26.400 429.450 27.450 ;
        RECT 428.400 -2.550 429.450 26.400 ;
        RECT 425.400 -3.600 429.450 -2.550 ;
      LAYER metal3 ;
        RECT 409.950 372.600 412.050 373.200 ;
        RECT 415.950 372.600 418.050 373.050 ;
        RECT 421.950 372.600 424.050 373.200 ;
        RECT 409.950 371.400 424.050 372.600 ;
        RECT 409.950 371.100 412.050 371.400 ;
        RECT 415.950 370.950 418.050 371.400 ;
        RECT 421.950 371.100 424.050 371.400 ;
        RECT 415.950 345.600 418.050 346.050 ;
        RECT 424.950 345.600 427.050 346.050 ;
        RECT 415.950 344.400 427.050 345.600 ;
        RECT 415.950 343.950 418.050 344.400 ;
        RECT 424.950 343.950 427.050 344.400 ;
        RECT 412.950 201.600 415.050 201.900 ;
        RECT 418.950 201.600 421.050 202.050 ;
        RECT 412.950 200.400 421.050 201.600 ;
        RECT 412.950 199.800 415.050 200.400 ;
        RECT 418.950 199.950 421.050 200.400 ;
        RECT 406.950 141.600 409.050 142.050 ;
        RECT 412.950 141.600 415.050 142.050 ;
        RECT 406.950 140.400 415.050 141.600 ;
        RECT 406.950 139.950 409.050 140.400 ;
        RECT 412.950 139.950 415.050 140.400 ;
        RECT 399.000 105.600 403.050 106.050 ;
        RECT 398.400 103.950 403.050 105.600 ;
        RECT 398.400 100.050 399.600 103.950 ;
        RECT 398.400 98.400 403.050 100.050 ;
        RECT 399.000 97.950 403.050 98.400 ;
        RECT 400.950 66.600 403.050 67.050 ;
        RECT 418.950 66.600 421.050 67.050 ;
        RECT 400.950 65.400 421.050 66.600 ;
        RECT 400.950 64.950 403.050 65.400 ;
        RECT 418.950 64.950 421.050 65.400 ;
    END
  END Xin[0]
  PIN Xout[3]
    PORT
      LAYER metal2 ;
        RECT 851.400 332.400 852.600 334.650 ;
        RECT 851.400 322.050 852.450 332.400 ;
        RECT 865.950 325.950 868.050 328.050 ;
        RECT 866.400 322.050 867.450 325.950 ;
        RECT 850.950 319.950 853.050 322.050 ;
        RECT 865.950 319.950 868.050 322.050 ;
      LAYER metal3 ;
        RECT 881.400 336.600 882.600 339.600 ;
        RECT 881.400 335.400 885.600 336.600 ;
        RECT 865.950 327.600 868.050 328.050 ;
        RECT 884.400 327.600 885.600 335.400 ;
        RECT 865.950 326.400 885.600 327.600 ;
        RECT 865.950 325.950 868.050 326.400 ;
        RECT 850.950 321.600 853.050 322.050 ;
        RECT 865.950 321.600 868.050 322.050 ;
        RECT 850.950 320.400 868.050 321.600 ;
        RECT 850.950 319.950 853.050 320.400 ;
        RECT 865.950 319.950 868.050 320.400 ;
    END
  END Xout[3]
  PIN Xout[2]
    PORT
      LAYER metal2 ;
        RECT 869.400 333.900 870.600 334.650 ;
        RECT 868.950 331.800 871.050 333.900 ;
      LAYER metal3 ;
        RECT 868.950 333.600 871.050 333.900 ;
        RECT 868.950 332.400 882.600 333.600 ;
        RECT 868.950 331.800 871.050 332.400 ;
    END
  END Xout[2]
  PIN Xout[1]
    PORT
      LAYER metal1 ;
        RECT 403.950 60.450 408.000 61.050 ;
        RECT 403.950 58.950 408.450 60.450 ;
        RECT 407.550 55.050 408.450 58.950 ;
        RECT 403.950 53.550 408.450 55.050 ;
        RECT 403.950 52.950 408.000 53.550 ;
        RECT 403.950 30.450 406.050 31.050 ;
        RECT 392.550 29.550 406.050 30.450 ;
        RECT 392.550 21.450 393.450 29.550 ;
        RECT 403.950 28.950 406.050 29.550 ;
        RECT 392.550 20.550 396.450 21.450 ;
        RECT 395.550 19.050 396.450 20.550 ;
        RECT 395.550 18.750 399.000 19.050 ;
        RECT 395.550 17.550 400.050 18.750 ;
        RECT 396.000 16.950 400.050 17.550 ;
        RECT 397.950 16.650 400.050 16.950 ;
      LAYER metal2 ;
        RECT 383.400 176.400 384.600 178.650 ;
        RECT 383.400 139.050 384.450 176.400 ;
        RECT 382.950 136.950 385.050 139.050 ;
        RECT 403.950 136.950 406.050 139.050 ;
        RECT 404.400 117.450 405.450 136.950 ;
        RECT 404.400 116.400 408.450 117.450 ;
        RECT 407.400 109.050 408.450 116.400 ;
        RECT 406.950 106.950 409.050 109.050 ;
        RECT 403.950 94.950 406.050 97.050 ;
        RECT 404.400 61.050 405.450 94.950 ;
        RECT 403.950 58.950 406.050 61.050 ;
        RECT 403.950 52.950 406.050 55.050 ;
        RECT 404.400 31.050 405.450 52.950 ;
        RECT 403.950 28.950 406.050 31.050 ;
        RECT 397.950 16.650 400.050 18.750 ;
        RECT 398.400 4.050 399.450 16.650 ;
        RECT 385.950 1.950 388.050 4.050 ;
        RECT 397.950 1.950 400.050 4.050 ;
        RECT 386.400 -3.600 387.450 1.950 ;
      LAYER metal3 ;
        RECT 382.950 138.600 385.050 139.050 ;
        RECT 403.950 138.600 406.050 139.050 ;
        RECT 382.950 137.400 406.050 138.600 ;
        RECT 382.950 136.950 385.050 137.400 ;
        RECT 403.950 136.950 406.050 137.400 ;
        RECT 406.950 106.950 409.050 109.050 ;
        RECT 407.400 97.050 408.600 106.950 ;
        RECT 403.950 95.400 408.600 97.050 ;
        RECT 403.950 94.950 408.000 95.400 ;
        RECT 385.950 3.600 388.050 4.050 ;
        RECT 397.950 3.600 400.050 4.050 ;
        RECT 385.950 2.400 400.050 3.600 ;
        RECT 385.950 1.950 388.050 2.400 ;
        RECT 397.950 1.950 400.050 2.400 ;
    END
  END Xout[1]
  PIN Xout[0]
    PORT
      LAYER metal1 ;
        RECT 346.950 108.450 349.050 109.200 ;
        RECT 341.550 107.550 349.050 108.450 ;
        RECT 341.550 100.050 342.450 107.550 ;
        RECT 346.950 107.100 349.050 107.550 ;
        RECT 341.550 98.550 346.050 100.050 ;
        RECT 342.000 97.950 346.050 98.550 ;
      LAYER metal2 ;
        RECT 371.400 176.400 372.600 178.650 ;
        RECT 371.400 160.050 372.450 176.400 ;
        RECT 346.950 157.950 349.050 160.050 ;
        RECT 370.950 157.950 373.050 160.050 ;
        RECT 347.400 109.200 348.450 157.950 ;
        RECT 346.950 107.100 349.050 109.200 ;
        RECT 343.950 97.950 346.050 100.050 ;
        RECT 344.400 82.050 345.450 97.950 ;
        RECT 343.950 79.950 346.050 82.050 ;
        RECT 361.950 79.950 364.050 82.050 ;
        RECT 362.400 61.050 363.450 79.950 ;
        RECT 361.950 58.950 364.050 61.050 ;
        RECT 361.950 52.950 364.050 55.050 ;
        RECT 362.400 43.050 363.450 52.950 ;
        RECT 349.950 40.950 352.050 43.050 ;
        RECT 361.950 40.950 364.050 43.050 ;
        RECT 350.400 4.050 351.450 40.950 ;
        RECT 349.950 1.950 352.050 4.050 ;
        RECT 367.950 1.950 370.050 4.050 ;
        RECT 368.400 -3.600 369.450 1.950 ;
      LAYER metal3 ;
        RECT 346.950 159.600 349.050 160.050 ;
        RECT 370.950 159.600 373.050 160.050 ;
        RECT 346.950 158.400 373.050 159.600 ;
        RECT 346.950 157.950 349.050 158.400 ;
        RECT 370.950 157.950 373.050 158.400 ;
        RECT 343.950 81.600 346.050 82.050 ;
        RECT 361.950 81.600 364.050 82.050 ;
        RECT 343.950 80.400 364.050 81.600 ;
        RECT 343.950 79.950 346.050 80.400 ;
        RECT 361.950 79.950 364.050 80.400 ;
        RECT 361.950 58.950 364.050 61.050 ;
        RECT 362.400 55.050 363.600 58.950 ;
        RECT 361.950 52.950 364.050 55.050 ;
        RECT 349.950 42.600 352.050 43.050 ;
        RECT 361.950 42.600 364.050 43.050 ;
        RECT 349.950 41.400 364.050 42.600 ;
        RECT 349.950 40.950 352.050 41.400 ;
        RECT 361.950 40.950 364.050 41.400 ;
        RECT 349.950 3.600 352.050 4.050 ;
        RECT 367.950 3.600 370.050 4.050 ;
        RECT 349.950 2.400 370.050 3.600 ;
        RECT 349.950 1.950 352.050 2.400 ;
        RECT 367.950 1.950 370.050 2.400 ;
    END
  END Xout[0]
  PIN Yin[3]
    PORT
      LAYER metal1 ;
        RECT 483.000 729.450 487.050 730.050 ;
        RECT 482.550 727.950 487.050 729.450 ;
        RECT 482.550 720.450 483.450 727.950 ;
        RECT 487.950 720.450 490.050 721.050 ;
        RECT 482.550 719.550 490.050 720.450 ;
        RECT 487.950 718.950 490.050 719.550 ;
      LAYER metal2 ;
        RECT 488.400 823.050 489.450 828.450 ;
        RECT 487.950 820.950 490.050 823.050 ;
        RECT 493.950 820.950 496.050 823.050 ;
        RECT 494.400 801.450 495.450 820.950 ;
        RECT 491.400 800.400 495.450 801.450 ;
        RECT 491.400 742.050 492.450 800.400 ;
        RECT 484.950 739.950 487.050 742.050 ;
        RECT 490.950 739.950 493.050 742.050 ;
        RECT 485.400 730.050 486.450 739.950 ;
        RECT 484.950 727.950 487.050 730.050 ;
        RECT 487.950 718.950 490.050 721.050 ;
        RECT 488.400 709.050 489.450 718.950 ;
        RECT 481.950 706.950 484.050 709.050 ;
        RECT 487.950 706.950 490.050 709.050 ;
        RECT 482.400 679.050 483.450 706.950 ;
        RECT 481.950 676.950 484.050 679.050 ;
        RECT 488.400 678.900 489.600 679.650 ;
        RECT 487.950 676.800 490.050 678.900 ;
      LAYER metal3 ;
        RECT 487.950 822.600 490.050 823.050 ;
        RECT 493.950 822.600 496.050 823.050 ;
        RECT 487.950 821.400 496.050 822.600 ;
        RECT 487.950 820.950 490.050 821.400 ;
        RECT 493.950 820.950 496.050 821.400 ;
        RECT 484.950 741.600 487.050 742.050 ;
        RECT 490.950 741.600 493.050 742.050 ;
        RECT 484.950 740.400 493.050 741.600 ;
        RECT 484.950 739.950 487.050 740.400 ;
        RECT 490.950 739.950 493.050 740.400 ;
        RECT 481.950 708.600 484.050 709.050 ;
        RECT 487.950 708.600 490.050 709.050 ;
        RECT 481.950 707.400 490.050 708.600 ;
        RECT 481.950 706.950 484.050 707.400 ;
        RECT 487.950 706.950 490.050 707.400 ;
        RECT 481.950 678.600 484.050 679.050 ;
        RECT 487.950 678.600 490.050 678.900 ;
        RECT 481.950 677.400 490.050 678.600 ;
        RECT 481.950 676.950 484.050 677.400 ;
        RECT 487.950 676.800 490.050 677.400 ;
    END
  END Yin[3]
  PIN Yin[2]
    PORT
      LAYER metal2 ;
        RECT 521.400 807.600 522.450 828.450 ;
        RECT 521.400 805.350 522.600 807.600 ;
    END
  END Yin[2]
  PIN Yin[1]
    PORT
      LAYER metal2 ;
        RECT 677.400 827.400 681.450 828.450 ;
        RECT 680.400 807.600 681.450 827.400 ;
        RECT 680.400 805.350 681.600 807.600 ;
    END
  END Yin[1]
  PIN Yin[0]
    PORT
      LAYER metal2 ;
        RECT 692.400 827.400 696.450 828.450 ;
        RECT 695.400 807.600 696.450 827.400 ;
        RECT 695.400 805.350 696.600 807.600 ;
    END
  END Yin[0]
  PIN Yout[3]
    PORT
      LAYER metal2 ;
        RECT 425.400 823.050 426.450 828.450 ;
        RECT 397.950 820.950 400.050 823.050 ;
        RECT 424.950 820.950 427.050 823.050 ;
        RECT 398.400 790.050 399.450 820.950 ;
        RECT 397.950 787.950 400.050 790.050 ;
        RECT 427.950 787.950 430.050 790.050 ;
        RECT 428.400 762.600 429.450 787.950 ;
        RECT 428.400 760.350 429.600 762.600 ;
      LAYER metal3 ;
        RECT 397.950 822.600 400.050 823.050 ;
        RECT 424.950 822.600 427.050 823.050 ;
        RECT 397.950 821.400 427.050 822.600 ;
        RECT 397.950 820.950 400.050 821.400 ;
        RECT 424.950 820.950 427.050 821.400 ;
        RECT 397.950 789.600 400.050 790.050 ;
        RECT 427.950 789.600 430.050 790.050 ;
        RECT 397.950 788.400 430.050 789.600 ;
        RECT 397.950 787.950 400.050 788.400 ;
        RECT 427.950 787.950 430.050 788.400 ;
    END
  END Yout[3]
  PIN Yout[2]
    PORT
      LAYER metal2 ;
        RECT 332.400 823.050 333.450 828.450 ;
        RECT 325.950 820.950 328.050 823.050 ;
        RECT 331.950 820.950 334.050 823.050 ;
        RECT 326.400 802.050 327.450 820.950 ;
        RECT 325.950 799.950 328.050 802.050 ;
        RECT 335.400 801.900 336.600 802.650 ;
        RECT 334.950 799.800 337.050 801.900 ;
      LAYER metal3 ;
        RECT 325.950 822.600 328.050 823.050 ;
        RECT 331.950 822.600 334.050 823.050 ;
        RECT 325.950 821.400 334.050 822.600 ;
        RECT 325.950 820.950 328.050 821.400 ;
        RECT 331.950 820.950 334.050 821.400 ;
        RECT 325.950 801.600 328.050 802.050 ;
        RECT 334.950 801.600 337.050 801.900 ;
        RECT 325.950 800.400 337.050 801.600 ;
        RECT 325.950 799.950 328.050 800.400 ;
        RECT 334.950 799.800 337.050 800.400 ;
    END
  END Yout[2]
  PIN Yout[1]
    PORT
      LAYER metal2 ;
        RECT 431.400 817.050 432.450 828.450 ;
        RECT 430.950 814.950 433.050 817.050 ;
        RECT 451.950 814.950 454.050 817.050 ;
        RECT 431.400 801.900 432.600 802.650 ;
        RECT 452.400 802.050 453.450 814.950 ;
        RECT 430.950 799.800 433.050 801.900 ;
        RECT 451.950 799.950 454.050 802.050 ;
      LAYER metal3 ;
        RECT 430.950 816.600 433.050 817.050 ;
        RECT 451.950 816.600 454.050 817.050 ;
        RECT 430.950 815.400 454.050 816.600 ;
        RECT 430.950 814.950 433.050 815.400 ;
        RECT 451.950 814.950 454.050 815.400 ;
        RECT 430.950 801.600 433.050 801.900 ;
        RECT 451.950 801.600 454.050 802.050 ;
        RECT 430.950 800.400 454.050 801.600 ;
        RECT 430.950 799.800 433.050 800.400 ;
        RECT 451.950 799.950 454.050 800.400 ;
    END
  END Yout[1]
  PIN Yout[0]
    PORT
      LAYER metal2 ;
        RECT 314.400 823.050 315.450 828.450 ;
        RECT 304.950 820.950 307.050 823.050 ;
        RECT 313.950 820.950 316.050 823.050 ;
        RECT 305.400 793.050 306.450 820.950 ;
        RECT 304.950 790.950 307.050 793.050 ;
        RECT 310.950 790.950 313.050 793.050 ;
        RECT 311.400 762.600 312.450 790.950 ;
        RECT 311.400 760.350 312.600 762.600 ;
      LAYER metal3 ;
        RECT 304.950 822.600 307.050 823.050 ;
        RECT 313.950 822.600 316.050 823.050 ;
        RECT 304.950 821.400 316.050 822.600 ;
        RECT 304.950 820.950 307.050 821.400 ;
        RECT 313.950 820.950 316.050 821.400 ;
        RECT 304.950 792.600 307.050 793.050 ;
        RECT 310.950 792.600 313.050 793.050 ;
        RECT 304.950 791.400 313.050 792.600 ;
        RECT 304.950 790.950 307.050 791.400 ;
        RECT 310.950 790.950 313.050 791.400 ;
    END
  END Yout[0]
  PIN clk
    PORT
      LAYER metal1 ;
        RECT 189.000 729.450 193.050 730.050 ;
        RECT 188.550 727.950 193.050 729.450 ;
        RECT 188.550 724.050 189.450 727.950 ;
        RECT 188.550 722.550 193.050 724.050 ;
        RECT 189.000 721.950 193.050 722.550 ;
      LAYER metal2 ;
        RECT 155.400 802.050 156.450 828.450 ;
        RECT 154.950 799.950 157.050 802.050 ;
        RECT 161.400 801.900 162.600 802.650 ;
        RECT 539.400 801.900 540.600 802.650 ;
        RECT 160.950 799.800 163.050 801.900 ;
        RECT 538.950 799.800 541.050 801.900 ;
        RECT 547.950 799.800 550.050 801.900 ;
        RECT 161.400 778.050 162.450 799.800 ;
        RECT 160.950 775.950 163.050 778.050 ;
        RECT 166.950 775.950 169.050 778.050 ;
        RECT 167.400 751.050 168.450 775.950 ;
        RECT 548.400 751.050 549.450 799.800 ;
        RECT 166.950 748.950 169.050 751.050 ;
        RECT 190.950 748.950 193.050 751.050 ;
        RECT 547.950 748.950 550.050 751.050 ;
        RECT 562.950 748.950 565.050 751.050 ;
        RECT 191.400 730.050 192.450 748.950 ;
        RECT 563.400 742.050 564.450 748.950 ;
        RECT 562.950 739.950 565.050 742.050 ;
        RECT 610.950 739.950 613.050 742.050 ;
        RECT 190.950 727.950 193.050 730.050 ;
        RECT 190.950 721.950 193.050 724.050 ;
        RECT 191.400 693.450 192.450 721.950 ;
        RECT 611.400 712.050 612.450 739.950 ;
        RECT 620.400 722.400 621.600 724.650 ;
        RECT 620.400 712.050 621.450 722.400 ;
        RECT 595.950 709.950 598.050 712.050 ;
        RECT 610.950 709.950 613.050 712.050 ;
        RECT 619.950 709.950 622.050 712.050 ;
        RECT 191.400 692.400 195.450 693.450 ;
        RECT 194.400 655.050 195.450 692.400 ;
        RECT 596.400 685.050 597.450 709.950 ;
        RECT 595.950 682.950 598.050 685.050 ;
        RECT 595.950 673.800 598.050 675.900 ;
        RECT 596.400 658.050 597.450 673.800 ;
        RECT 343.950 655.950 346.050 658.050 ;
        RECT 595.950 655.950 598.050 658.050 ;
        RECT 193.950 652.950 196.050 655.050 ;
        RECT 223.950 652.950 226.050 655.050 ;
        RECT 224.400 625.050 225.450 652.950 ;
        RECT 266.400 645.450 267.600 646.650 ;
        RECT 263.400 644.400 267.600 645.450 ;
        RECT 263.400 628.050 264.450 644.400 ;
        RECT 262.950 625.950 265.050 628.050 ;
        RECT 223.950 622.950 226.050 625.050 ;
        RECT 224.400 573.450 225.450 622.950 ;
        RECT 263.400 613.050 264.450 625.950 ;
        RECT 344.400 613.050 345.450 655.950 ;
        RECT 262.950 610.950 265.050 613.050 ;
        RECT 343.950 610.950 346.050 613.050 ;
        RECT 221.400 572.400 225.450 573.450 ;
        RECT 221.400 529.200 222.450 572.400 ;
        RECT 344.400 559.050 345.450 610.950 ;
        RECT 647.400 566.400 648.600 568.650 ;
        RECT 616.950 559.950 619.050 562.050 ;
        RECT 631.950 559.950 634.050 562.050 ;
        RECT 343.950 556.950 346.050 559.050 ;
        RECT 349.950 556.950 352.050 559.050 ;
        RECT 350.400 541.050 351.450 556.950 ;
        RECT 617.400 550.050 618.450 559.950 ;
        RECT 632.400 553.050 633.450 559.950 ;
        RECT 647.400 553.050 648.450 566.400 ;
        RECT 631.950 550.950 634.050 553.050 ;
        RECT 646.950 550.950 649.050 553.050 ;
        RECT 601.950 547.950 604.050 550.050 ;
        RECT 616.950 547.950 619.050 550.050 ;
        RECT 602.400 544.050 603.450 547.950 ;
        RECT 526.950 541.950 529.050 544.050 ;
        RECT 601.950 541.950 604.050 544.050 ;
        RECT 349.950 538.950 352.050 541.050 ;
        RECT 214.950 527.100 217.050 529.200 ;
        RECT 220.950 527.100 223.050 529.200 ;
        RECT 215.400 526.350 216.600 527.100 ;
        RECT 347.400 489.450 348.600 490.650 ;
        RECT 350.400 489.450 351.450 538.950 ;
        RECT 499.950 535.950 502.050 538.050 ;
        RECT 500.400 520.050 501.450 535.950 ;
        RECT 527.400 520.050 528.450 541.950 ;
        RECT 499.950 517.950 502.050 520.050 ;
        RECT 526.950 517.950 529.050 520.050 ;
        RECT 527.400 499.050 528.450 517.950 ;
        RECT 526.950 496.950 529.050 499.050 ;
        RECT 550.950 496.950 553.050 499.050 ;
        RECT 551.400 489.900 552.450 496.950 ;
        RECT 557.400 489.900 558.600 490.650 ;
        RECT 347.400 488.400 351.450 489.450 ;
        RECT 550.950 487.800 553.050 489.900 ;
        RECT 556.950 487.800 559.050 489.900 ;
      LAYER metal3 ;
        RECT 154.950 801.600 157.050 802.050 ;
        RECT 160.950 801.600 163.050 801.900 ;
        RECT 154.950 800.400 163.050 801.600 ;
        RECT 154.950 799.950 157.050 800.400 ;
        RECT 160.950 799.800 163.050 800.400 ;
        RECT 538.950 801.450 541.050 801.900 ;
        RECT 547.950 801.450 550.050 801.900 ;
        RECT 538.950 800.250 550.050 801.450 ;
        RECT 538.950 799.800 541.050 800.250 ;
        RECT 547.950 799.800 550.050 800.250 ;
        RECT 160.950 777.600 163.050 778.050 ;
        RECT 166.950 777.600 169.050 778.050 ;
        RECT 160.950 776.400 169.050 777.600 ;
        RECT 160.950 775.950 163.050 776.400 ;
        RECT 166.950 775.950 169.050 776.400 ;
        RECT 166.950 750.600 169.050 751.050 ;
        RECT 190.950 750.600 193.050 751.050 ;
        RECT 166.950 749.400 193.050 750.600 ;
        RECT 166.950 748.950 169.050 749.400 ;
        RECT 190.950 748.950 193.050 749.400 ;
        RECT 547.950 750.600 550.050 751.050 ;
        RECT 562.950 750.600 565.050 751.050 ;
        RECT 547.950 749.400 565.050 750.600 ;
        RECT 547.950 748.950 550.050 749.400 ;
        RECT 562.950 748.950 565.050 749.400 ;
        RECT 562.950 741.600 565.050 742.050 ;
        RECT 610.950 741.600 613.050 742.050 ;
        RECT 562.950 740.400 613.050 741.600 ;
        RECT 562.950 739.950 565.050 740.400 ;
        RECT 610.950 739.950 613.050 740.400 ;
        RECT 595.950 711.600 598.050 712.050 ;
        RECT 610.950 711.600 613.050 712.050 ;
        RECT 619.950 711.600 622.050 712.050 ;
        RECT 595.950 710.400 622.050 711.600 ;
        RECT 595.950 709.950 598.050 710.400 ;
        RECT 610.950 709.950 613.050 710.400 ;
        RECT 619.950 709.950 622.050 710.400 ;
        RECT 595.950 682.950 598.050 685.050 ;
        RECT 596.400 675.900 597.600 682.950 ;
        RECT 595.950 673.800 598.050 675.900 ;
        RECT 343.950 657.600 346.050 658.050 ;
        RECT 595.950 657.600 598.050 658.050 ;
        RECT 343.950 656.400 598.050 657.600 ;
        RECT 343.950 655.950 346.050 656.400 ;
        RECT 595.950 655.950 598.050 656.400 ;
        RECT 193.950 654.600 196.050 655.050 ;
        RECT 223.950 654.600 226.050 655.050 ;
        RECT 193.950 653.400 226.050 654.600 ;
        RECT 193.950 652.950 196.050 653.400 ;
        RECT 223.950 652.950 226.050 653.400 ;
        RECT 262.950 627.600 265.050 628.050 ;
        RECT 248.400 626.400 265.050 627.600 ;
        RECT 223.950 624.600 226.050 625.050 ;
        RECT 248.400 624.600 249.600 626.400 ;
        RECT 262.950 625.950 265.050 626.400 ;
        RECT 223.950 623.400 249.600 624.600 ;
        RECT 223.950 622.950 226.050 623.400 ;
        RECT 262.950 612.600 265.050 613.050 ;
        RECT 343.950 612.600 346.050 613.050 ;
        RECT 262.950 611.400 346.050 612.600 ;
        RECT 262.950 610.950 265.050 611.400 ;
        RECT 343.950 610.950 346.050 611.400 ;
        RECT 616.950 561.600 619.050 562.050 ;
        RECT 631.950 561.600 634.050 562.050 ;
        RECT 616.950 560.400 634.050 561.600 ;
        RECT 616.950 559.950 619.050 560.400 ;
        RECT 631.950 559.950 634.050 560.400 ;
        RECT 343.950 558.600 346.050 559.050 ;
        RECT 349.950 558.600 352.050 559.050 ;
        RECT 343.950 557.400 352.050 558.600 ;
        RECT 343.950 556.950 346.050 557.400 ;
        RECT 349.950 556.950 352.050 557.400 ;
        RECT 631.950 552.600 634.050 553.050 ;
        RECT 646.950 552.600 649.050 553.050 ;
        RECT 631.950 551.400 649.050 552.600 ;
        RECT 631.950 550.950 634.050 551.400 ;
        RECT 646.950 550.950 649.050 551.400 ;
        RECT 601.950 549.600 604.050 550.050 ;
        RECT 616.950 549.600 619.050 550.050 ;
        RECT 601.950 548.400 619.050 549.600 ;
        RECT 601.950 547.950 604.050 548.400 ;
        RECT 616.950 547.950 619.050 548.400 ;
        RECT 526.950 543.600 529.050 544.050 ;
        RECT 601.950 543.600 604.050 544.050 ;
        RECT 526.950 542.400 604.050 543.600 ;
        RECT 526.950 541.950 529.050 542.400 ;
        RECT 601.950 541.950 604.050 542.400 ;
        RECT 349.950 540.600 352.050 541.050 ;
        RECT 349.950 539.400 498.600 540.600 ;
        RECT 349.950 538.950 352.050 539.400 ;
        RECT 497.400 538.050 498.600 539.400 ;
        RECT 497.400 536.400 502.050 538.050 ;
        RECT 498.000 535.950 502.050 536.400 ;
        RECT 214.950 528.750 217.050 529.200 ;
        RECT 220.950 528.750 223.050 529.200 ;
        RECT 214.950 527.550 223.050 528.750 ;
        RECT 214.950 527.100 217.050 527.550 ;
        RECT 220.950 527.100 223.050 527.550 ;
        RECT 499.950 519.600 502.050 520.050 ;
        RECT 526.950 519.600 529.050 520.050 ;
        RECT 499.950 518.400 529.050 519.600 ;
        RECT 499.950 517.950 502.050 518.400 ;
        RECT 526.950 517.950 529.050 518.400 ;
        RECT 526.950 498.600 529.050 499.050 ;
        RECT 550.950 498.600 553.050 499.050 ;
        RECT 526.950 497.400 553.050 498.600 ;
        RECT 526.950 496.950 529.050 497.400 ;
        RECT 550.950 496.950 553.050 497.400 ;
        RECT 550.950 489.450 553.050 489.900 ;
        RECT 556.950 489.450 559.050 489.900 ;
        RECT 550.950 488.250 559.050 489.450 ;
        RECT 550.950 487.800 553.050 488.250 ;
        RECT 556.950 487.800 559.050 488.250 ;
    END
  END clk
  OBS
      LAYER metal1 ;
        RECT 3.150 814.200 4.950 818.400 ;
        RECT 2.550 812.400 4.950 814.200 ;
        RECT 6.150 812.400 7.950 819.000 ;
        RECT 10.950 816.300 12.750 818.400 ;
        RECT 9.150 815.400 12.750 816.300 ;
        RECT 15.450 815.400 17.250 819.000 ;
        RECT 18.750 815.400 20.550 818.400 ;
        RECT 21.750 815.400 23.550 819.000 ;
        RECT 26.250 815.400 28.050 818.400 ;
        RECT 8.850 814.800 12.750 815.400 ;
        RECT 8.850 813.300 10.950 814.800 ;
        RECT 18.750 814.500 19.800 815.400 ;
        RECT 2.550 797.700 3.450 812.400 ;
        RECT 11.850 811.800 13.650 813.600 ;
        RECT 14.850 813.450 19.800 814.500 ;
        RECT 14.850 812.700 16.650 813.450 ;
        RECT 26.250 813.300 28.650 815.400 ;
        RECT 31.350 812.400 33.150 819.000 ;
        RECT 34.650 812.400 36.450 818.400 ;
        RECT 47.100 815.400 48.900 818.400 ;
        RECT 50.100 815.400 51.900 819.000 ;
        RECT 11.850 810.000 12.900 811.800 ;
        RECT 22.050 810.000 23.850 810.600 ;
        RECT 11.850 808.800 23.850 810.000 ;
        RECT 4.950 807.600 12.900 808.800 ;
        RECT 4.950 805.050 6.750 807.600 ;
        RECT 11.100 807.000 12.900 807.600 ;
        RECT 8.100 805.800 9.900 806.400 ;
        RECT 4.950 802.950 7.050 805.050 ;
        RECT 8.100 804.600 16.200 805.800 ;
        RECT 14.100 802.950 16.200 804.600 ;
        RECT 12.450 797.700 14.250 798.000 ;
        RECT 2.550 797.100 14.250 797.700 ;
        RECT 2.550 796.500 20.850 797.100 ;
        RECT 2.550 795.600 3.450 796.500 ;
        RECT 12.450 796.200 20.850 796.500 ;
        RECT 2.550 793.800 4.950 795.600 ;
        RECT 3.150 783.600 4.950 793.800 ;
        RECT 6.150 783.000 7.950 795.600 ;
        RECT 17.250 794.700 19.050 795.300 ;
        RECT 11.250 793.500 19.050 794.700 ;
        RECT 19.950 794.100 20.850 796.200 ;
        RECT 22.950 796.200 23.850 808.800 ;
        RECT 35.250 805.050 36.450 812.400 ;
        RECT 47.700 805.050 48.900 815.400 ;
        RECT 53.550 812.400 55.350 818.400 ;
        RECT 56.850 812.400 58.650 819.000 ;
        RECT 61.950 815.400 63.750 818.400 ;
        RECT 66.450 815.400 68.250 819.000 ;
        RECT 69.450 815.400 71.250 818.400 ;
        RECT 72.750 815.400 74.550 819.000 ;
        RECT 77.250 816.300 79.050 818.400 ;
        RECT 77.250 815.400 80.850 816.300 ;
        RECT 61.350 813.300 63.750 815.400 ;
        RECT 70.200 814.500 71.250 815.400 ;
        RECT 77.250 814.800 81.150 815.400 ;
        RECT 70.200 813.450 75.150 814.500 ;
        RECT 73.350 812.700 75.150 813.450 ;
        RECT 53.550 805.050 54.750 812.400 ;
        RECT 76.350 811.800 78.150 813.600 ;
        RECT 79.050 813.300 81.150 814.800 ;
        RECT 82.050 812.400 83.850 819.000 ;
        RECT 85.050 814.200 86.850 818.400 ;
        RECT 85.050 812.400 87.450 814.200 ;
        RECT 66.150 810.000 67.950 810.600 ;
        RECT 77.100 810.000 78.150 811.800 ;
        RECT 66.150 808.800 78.150 810.000 ;
        RECT 30.150 803.250 36.450 805.050 ;
        RECT 31.950 802.950 36.450 803.250 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 49.950 802.950 52.050 805.050 ;
        RECT 53.550 803.250 59.850 805.050 ;
        RECT 53.550 802.950 58.050 803.250 ;
        RECT 26.550 800.100 28.650 800.400 ;
        RECT 32.550 800.100 34.350 800.250 ;
        RECT 26.550 798.900 34.350 800.100 ;
        RECT 26.550 798.300 28.650 798.900 ;
        RECT 32.550 798.450 34.350 798.900 ;
        RECT 22.950 795.300 27.750 796.200 ;
        RECT 35.250 795.600 36.450 802.950 ;
        RECT 26.550 794.400 27.750 795.300 ;
        RECT 23.850 794.100 25.650 794.400 ;
        RECT 11.250 792.600 13.350 793.500 ;
        RECT 19.950 793.200 25.650 794.100 ;
        RECT 23.850 792.600 25.650 793.200 ;
        RECT 26.550 792.600 29.550 794.400 ;
        RECT 11.550 783.600 13.350 792.600 ;
        RECT 15.450 791.550 17.250 792.300 ;
        RECT 20.250 791.550 22.050 792.300 ;
        RECT 15.450 790.500 22.050 791.550 ;
        RECT 16.350 783.000 18.150 789.600 ;
        RECT 19.350 783.600 21.150 790.500 ;
        RECT 26.550 789.600 28.650 791.700 ;
        RECT 22.350 783.000 24.150 789.600 ;
        RECT 26.850 783.600 28.650 789.600 ;
        RECT 31.650 783.000 33.450 795.600 ;
        RECT 34.650 783.600 36.450 795.600 ;
        RECT 47.700 789.600 48.900 802.950 ;
        RECT 50.100 801.150 51.900 802.950 ;
        RECT 53.550 795.600 54.750 802.950 ;
        RECT 55.650 800.100 57.450 800.250 ;
        RECT 61.350 800.100 63.450 800.400 ;
        RECT 55.650 798.900 63.450 800.100 ;
        RECT 55.650 798.450 57.450 798.900 ;
        RECT 61.350 798.300 63.450 798.900 ;
        RECT 66.150 796.200 67.050 808.800 ;
        RECT 77.100 807.600 85.050 808.800 ;
        RECT 77.100 807.000 78.900 807.600 ;
        RECT 80.100 805.800 81.900 806.400 ;
        RECT 73.800 804.600 81.900 805.800 ;
        RECT 83.250 805.050 85.050 807.600 ;
        RECT 73.800 802.950 75.900 804.600 ;
        RECT 82.950 802.950 85.050 805.050 ;
        RECT 75.750 797.700 77.550 798.000 ;
        RECT 86.550 797.700 87.450 812.400 ;
        RECT 98.100 813.300 99.900 818.400 ;
        RECT 101.100 814.200 102.900 819.000 ;
        RECT 104.100 813.300 105.900 818.400 ;
        RECT 98.100 811.950 105.900 813.300 ;
        RECT 107.100 812.400 108.900 818.400 ;
        RECT 119.400 812.400 121.200 819.000 ;
        RECT 107.100 810.300 108.300 812.400 ;
        RECT 124.500 811.200 126.300 818.400 ;
        RECT 140.100 812.400 141.900 819.000 ;
        RECT 143.100 811.500 144.900 818.400 ;
        RECT 146.100 812.400 147.900 819.000 ;
        RECT 149.100 811.500 150.900 818.400 ;
        RECT 152.100 812.400 153.900 819.000 ;
        RECT 155.100 811.500 156.900 818.400 ;
        RECT 158.100 812.400 159.900 819.000 ;
        RECT 161.100 811.500 162.900 818.400 ;
        RECT 164.100 812.400 165.900 819.000 ;
        RECT 168.150 814.200 169.950 818.400 ;
        RECT 167.550 812.400 169.950 814.200 ;
        RECT 171.150 812.400 172.950 819.000 ;
        RECT 175.950 816.300 177.750 818.400 ;
        RECT 174.150 815.400 177.750 816.300 ;
        RECT 180.450 815.400 182.250 819.000 ;
        RECT 183.750 815.400 185.550 818.400 ;
        RECT 186.750 815.400 188.550 819.000 ;
        RECT 191.250 815.400 193.050 818.400 ;
        RECT 173.850 814.800 177.750 815.400 ;
        RECT 173.850 813.300 175.950 814.800 ;
        RECT 183.750 814.500 184.800 815.400 ;
        RECT 104.700 809.400 108.300 810.300 ;
        RECT 122.100 810.300 126.300 811.200 ;
        RECT 142.050 810.300 144.900 811.500 ;
        RECT 147.000 810.300 150.900 811.500 ;
        RECT 153.000 810.300 156.900 811.500 ;
        RECT 159.000 810.300 162.900 811.500 ;
        RECT 101.100 805.050 102.900 806.850 ;
        RECT 104.700 805.050 105.900 809.400 ;
        RECT 107.100 805.050 108.900 806.850 ;
        RECT 119.250 805.050 121.050 806.850 ;
        RECT 122.100 805.050 123.300 810.300 ;
        RECT 125.100 805.050 126.900 806.850 ;
        RECT 142.050 805.050 143.100 810.300 ;
        RECT 147.000 809.400 148.200 810.300 ;
        RECT 153.000 809.400 154.200 810.300 ;
        RECT 159.000 809.400 160.200 810.300 ;
        RECT 144.000 808.200 148.200 809.400 ;
        RECT 144.000 807.600 145.800 808.200 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 100.950 802.950 103.050 805.050 ;
        RECT 103.950 802.950 106.050 805.050 ;
        RECT 106.950 802.950 109.050 805.050 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 142.050 802.950 145.200 805.050 ;
        RECT 98.100 801.150 99.900 802.950 ;
        RECT 75.750 797.100 87.450 797.700 ;
        RECT 47.100 783.600 48.900 789.600 ;
        RECT 50.100 783.000 51.900 789.600 ;
        RECT 53.550 783.600 55.350 795.600 ;
        RECT 56.550 783.000 58.350 795.600 ;
        RECT 62.250 795.300 67.050 796.200 ;
        RECT 69.150 796.500 87.450 797.100 ;
        RECT 69.150 796.200 77.550 796.500 ;
        RECT 62.250 794.400 63.450 795.300 ;
        RECT 60.450 792.600 63.450 794.400 ;
        RECT 64.350 794.100 66.150 794.400 ;
        RECT 69.150 794.100 70.050 796.200 ;
        RECT 86.550 795.600 87.450 796.500 ;
        RECT 104.700 795.600 105.900 802.950 ;
        RECT 64.350 793.200 70.050 794.100 ;
        RECT 70.950 794.700 72.750 795.300 ;
        RECT 70.950 793.500 78.750 794.700 ;
        RECT 64.350 792.600 66.150 793.200 ;
        RECT 76.650 792.600 78.750 793.500 ;
        RECT 61.350 789.600 63.450 791.700 ;
        RECT 67.950 791.550 69.750 792.300 ;
        RECT 72.750 791.550 74.550 792.300 ;
        RECT 67.950 790.500 74.550 791.550 ;
        RECT 61.350 783.600 63.150 789.600 ;
        RECT 65.850 783.000 67.650 789.600 ;
        RECT 68.850 783.600 70.650 790.500 ;
        RECT 71.850 783.000 73.650 789.600 ;
        RECT 76.650 783.600 78.450 792.600 ;
        RECT 82.050 783.000 83.850 795.600 ;
        RECT 85.050 793.800 87.450 795.600 ;
        RECT 85.050 783.600 86.850 793.800 ;
        RECT 98.400 783.000 100.200 795.600 ;
        RECT 103.500 794.100 105.900 795.600 ;
        RECT 103.500 783.600 105.300 794.100 ;
        RECT 106.200 791.100 108.000 792.900 ;
        RECT 122.100 789.600 123.300 802.950 ;
        RECT 142.050 797.700 143.100 802.950 ;
        RECT 147.000 797.700 148.200 808.200 ;
        RECT 150.000 808.200 154.200 809.400 ;
        RECT 150.000 807.600 151.800 808.200 ;
        RECT 153.000 797.700 154.200 808.200 ;
        RECT 156.000 808.200 160.200 809.400 ;
        RECT 156.000 807.600 157.800 808.200 ;
        RECT 159.000 797.700 160.200 808.200 ;
        RECT 161.400 805.050 163.200 806.850 ;
        RECT 161.100 802.950 163.200 805.050 ;
        RECT 167.550 797.700 168.450 812.400 ;
        RECT 176.850 811.800 178.650 813.600 ;
        RECT 179.850 813.450 184.800 814.500 ;
        RECT 179.850 812.700 181.650 813.450 ;
        RECT 191.250 813.300 193.650 815.400 ;
        RECT 196.350 812.400 198.150 819.000 ;
        RECT 199.650 812.400 201.450 818.400 ;
        RECT 212.100 815.400 213.900 819.000 ;
        RECT 215.100 815.400 216.900 818.400 ;
        RECT 176.850 810.000 177.900 811.800 ;
        RECT 187.050 810.000 188.850 810.600 ;
        RECT 176.850 808.800 188.850 810.000 ;
        RECT 169.950 807.600 177.900 808.800 ;
        RECT 169.950 805.050 171.750 807.600 ;
        RECT 176.100 807.000 177.900 807.600 ;
        RECT 173.100 805.800 174.900 806.400 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 173.100 804.600 181.200 805.800 ;
        RECT 179.100 802.950 181.200 804.600 ;
        RECT 177.450 797.700 179.250 798.000 ;
        RECT 142.050 796.500 144.900 797.700 ;
        RECT 147.000 796.500 150.900 797.700 ;
        RECT 153.000 796.500 156.900 797.700 ;
        RECT 159.000 796.500 162.900 797.700 ;
        RECT 106.500 783.000 108.300 789.600 ;
        RECT 119.100 783.000 120.900 789.600 ;
        RECT 122.100 783.600 123.900 789.600 ;
        RECT 125.100 783.000 126.900 789.600 ;
        RECT 140.100 783.000 141.900 795.600 ;
        RECT 143.100 783.600 144.900 796.500 ;
        RECT 146.100 783.000 147.900 795.600 ;
        RECT 149.100 783.600 150.900 796.500 ;
        RECT 152.100 783.000 153.900 795.600 ;
        RECT 155.100 783.600 156.900 796.500 ;
        RECT 158.100 783.000 159.900 795.600 ;
        RECT 161.100 783.600 162.900 796.500 ;
        RECT 167.550 797.100 179.250 797.700 ;
        RECT 167.550 796.500 185.850 797.100 ;
        RECT 167.550 795.600 168.450 796.500 ;
        RECT 177.450 796.200 185.850 796.500 ;
        RECT 164.100 783.000 165.900 795.600 ;
        RECT 167.550 793.800 169.950 795.600 ;
        RECT 168.150 783.600 169.950 793.800 ;
        RECT 171.150 783.000 172.950 795.600 ;
        RECT 182.250 794.700 184.050 795.300 ;
        RECT 176.250 793.500 184.050 794.700 ;
        RECT 184.950 794.100 185.850 796.200 ;
        RECT 187.950 796.200 188.850 808.800 ;
        RECT 200.250 805.050 201.450 812.400 ;
        RECT 215.100 805.050 216.300 815.400 ;
        RECT 227.100 813.300 228.900 818.400 ;
        RECT 230.100 814.200 231.900 819.000 ;
        RECT 233.100 813.300 234.900 818.400 ;
        RECT 227.100 811.950 234.900 813.300 ;
        RECT 236.100 812.400 237.900 818.400 ;
        RECT 248.400 812.400 250.200 819.000 ;
        RECT 217.950 810.450 220.050 811.050 ;
        RECT 223.950 810.450 226.050 811.050 ;
        RECT 217.950 809.550 226.050 810.450 ;
        RECT 236.100 810.300 237.300 812.400 ;
        RECT 253.500 811.200 255.300 818.400 ;
        RECT 266.400 812.400 268.200 819.000 ;
        RECT 271.500 811.200 273.300 818.400 ;
        RECT 288.600 814.200 290.400 818.400 ;
        RECT 217.950 808.950 220.050 809.550 ;
        RECT 223.950 808.950 226.050 809.550 ;
        RECT 233.700 809.400 237.300 810.300 ;
        RECT 251.100 810.300 255.300 811.200 ;
        RECT 269.100 810.300 273.300 811.200 ;
        RECT 287.700 812.400 290.400 814.200 ;
        RECT 291.600 812.400 293.400 819.000 ;
        RECT 230.100 805.050 231.900 806.850 ;
        RECT 233.700 805.050 234.900 809.400 ;
        RECT 236.100 805.050 237.900 806.850 ;
        RECT 248.250 805.050 250.050 806.850 ;
        RECT 251.100 805.050 252.300 810.300 ;
        RECT 254.100 805.050 255.900 806.850 ;
        RECT 266.250 805.050 268.050 806.850 ;
        RECT 269.100 805.050 270.300 810.300 ;
        RECT 272.100 805.050 273.900 806.850 ;
        RECT 287.700 805.050 288.600 812.400 ;
        RECT 289.500 810.600 291.300 811.500 ;
        RECT 296.100 810.600 297.900 818.400 ;
        RECT 289.500 809.700 297.900 810.600 ;
        RECT 308.100 812.400 309.900 818.400 ;
        RECT 311.100 813.000 312.900 819.000 ;
        RECT 317.700 818.400 318.900 819.000 ;
        RECT 314.100 815.400 315.900 818.400 ;
        RECT 317.100 815.400 318.900 818.400 ;
        RECT 329.100 815.400 330.900 818.400 ;
        RECT 195.150 803.250 201.450 805.050 ;
        RECT 196.950 802.950 201.450 803.250 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 226.950 802.950 229.050 805.050 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 287.100 802.950 289.200 805.050 ;
        RECT 290.400 802.950 292.500 805.050 ;
        RECT 191.550 800.100 193.650 800.400 ;
        RECT 197.550 800.100 199.350 800.250 ;
        RECT 191.550 798.900 199.350 800.100 ;
        RECT 191.550 798.300 193.650 798.900 ;
        RECT 197.550 798.450 199.350 798.900 ;
        RECT 187.950 795.300 192.750 796.200 ;
        RECT 200.250 795.600 201.450 802.950 ;
        RECT 212.100 801.150 213.900 802.950 ;
        RECT 191.550 794.400 192.750 795.300 ;
        RECT 188.850 794.100 190.650 794.400 ;
        RECT 176.250 792.600 178.350 793.500 ;
        RECT 184.950 793.200 190.650 794.100 ;
        RECT 188.850 792.600 190.650 793.200 ;
        RECT 191.550 792.600 194.550 794.400 ;
        RECT 176.550 783.600 178.350 792.600 ;
        RECT 180.450 791.550 182.250 792.300 ;
        RECT 185.250 791.550 187.050 792.300 ;
        RECT 180.450 790.500 187.050 791.550 ;
        RECT 181.350 783.000 183.150 789.600 ;
        RECT 184.350 783.600 186.150 790.500 ;
        RECT 191.550 789.600 193.650 791.700 ;
        RECT 187.350 783.000 189.150 789.600 ;
        RECT 191.850 783.600 193.650 789.600 ;
        RECT 196.650 783.000 198.450 795.600 ;
        RECT 199.650 783.600 201.450 795.600 ;
        RECT 215.100 789.600 216.300 802.950 ;
        RECT 227.100 801.150 228.900 802.950 ;
        RECT 233.700 795.600 234.900 802.950 ;
        RECT 212.100 783.000 213.900 789.600 ;
        RECT 215.100 783.600 216.900 789.600 ;
        RECT 227.400 783.000 229.200 795.600 ;
        RECT 232.500 794.100 234.900 795.600 ;
        RECT 232.500 783.600 234.300 794.100 ;
        RECT 235.200 791.100 237.000 792.900 ;
        RECT 251.100 789.600 252.300 802.950 ;
        RECT 253.950 792.450 256.050 793.050 ;
        RECT 265.950 792.450 268.050 792.900 ;
        RECT 253.950 791.550 268.050 792.450 ;
        RECT 253.950 790.950 256.050 791.550 ;
        RECT 265.950 790.800 268.050 791.550 ;
        RECT 269.100 789.600 270.300 802.950 ;
        RECT 287.700 795.600 288.600 802.950 ;
        RECT 291.000 801.150 292.800 802.950 ;
        RECT 235.500 783.000 237.300 789.600 ;
        RECT 248.100 783.000 249.900 789.600 ;
        RECT 251.100 783.600 252.900 789.600 ;
        RECT 254.100 783.000 255.900 789.600 ;
        RECT 266.100 783.000 267.900 789.600 ;
        RECT 269.100 783.600 270.900 789.600 ;
        RECT 272.100 783.000 273.900 789.600 ;
        RECT 287.100 783.600 288.900 795.600 ;
        RECT 290.100 783.000 291.900 795.000 ;
        RECT 294.000 789.600 294.900 809.700 ;
        RECT 295.950 805.050 297.750 806.850 ;
        RECT 308.100 805.050 309.000 812.400 ;
        RECT 314.700 811.200 315.600 815.400 ;
        RECT 310.200 810.300 315.600 811.200 ;
        RECT 329.100 811.500 330.300 815.400 ;
        RECT 332.100 812.400 333.900 819.000 ;
        RECT 335.100 812.400 336.900 818.400 ;
        RECT 339.150 814.200 340.950 818.400 ;
        RECT 329.100 810.600 334.800 811.500 ;
        RECT 310.200 809.400 312.300 810.300 ;
        RECT 295.800 802.950 297.900 805.050 ;
        RECT 308.100 802.950 310.200 805.050 ;
        RECT 309.000 795.600 310.200 802.950 ;
        RECT 311.400 798.900 312.300 809.400 ;
        RECT 333.000 809.700 334.800 810.600 ;
        RECT 316.800 805.050 318.600 806.850 ;
        RECT 313.500 802.950 315.600 805.050 ;
        RECT 316.800 802.950 318.900 805.050 ;
        RECT 329.400 802.950 331.500 805.050 ;
        RECT 313.200 801.150 315.000 802.950 ;
        RECT 329.400 801.150 331.200 802.950 ;
        RECT 311.100 798.300 312.900 798.900 ;
        RECT 333.000 798.300 333.900 809.700 ;
        RECT 335.700 805.050 336.900 812.400 ;
        RECT 334.800 802.950 336.900 805.050 ;
        RECT 311.100 797.100 318.900 798.300 ;
        RECT 333.000 797.400 334.800 798.300 ;
        RECT 317.700 795.600 318.900 797.100 ;
        RECT 309.000 794.100 311.400 795.600 ;
        RECT 293.100 783.600 294.900 789.600 ;
        RECT 296.100 783.000 297.900 789.600 ;
        RECT 309.600 783.600 311.400 794.100 ;
        RECT 312.600 783.000 314.400 795.600 ;
        RECT 317.100 783.600 318.900 795.600 ;
        RECT 329.100 796.500 334.800 797.400 ;
        RECT 329.100 789.600 330.300 796.500 ;
        RECT 335.700 795.600 336.900 802.950 ;
        RECT 329.100 783.600 330.900 789.600 ;
        RECT 332.100 783.000 333.900 793.800 ;
        RECT 335.100 783.600 336.900 795.600 ;
        RECT 338.550 812.400 340.950 814.200 ;
        RECT 342.150 812.400 343.950 819.000 ;
        RECT 346.950 816.300 348.750 818.400 ;
        RECT 345.150 815.400 348.750 816.300 ;
        RECT 351.450 815.400 353.250 819.000 ;
        RECT 354.750 815.400 356.550 818.400 ;
        RECT 357.750 815.400 359.550 819.000 ;
        RECT 362.250 815.400 364.050 818.400 ;
        RECT 344.850 814.800 348.750 815.400 ;
        RECT 344.850 813.300 346.950 814.800 ;
        RECT 354.750 814.500 355.800 815.400 ;
        RECT 338.550 797.700 339.450 812.400 ;
        RECT 347.850 811.800 349.650 813.600 ;
        RECT 350.850 813.450 355.800 814.500 ;
        RECT 350.850 812.700 352.650 813.450 ;
        RECT 362.250 813.300 364.650 815.400 ;
        RECT 367.350 812.400 369.150 819.000 ;
        RECT 370.650 812.400 372.450 818.400 ;
        RECT 383.100 815.400 384.900 819.000 ;
        RECT 386.100 815.400 387.900 818.400 ;
        RECT 389.100 815.400 390.900 819.000 ;
        RECT 404.700 815.400 406.500 819.000 ;
        RECT 347.850 810.000 348.900 811.800 ;
        RECT 358.050 810.000 359.850 810.600 ;
        RECT 347.850 808.800 359.850 810.000 ;
        RECT 340.950 807.600 348.900 808.800 ;
        RECT 340.950 805.050 342.750 807.600 ;
        RECT 347.100 807.000 348.900 807.600 ;
        RECT 344.100 805.800 345.900 806.400 ;
        RECT 340.950 802.950 343.050 805.050 ;
        RECT 344.100 804.600 352.200 805.800 ;
        RECT 350.100 802.950 352.200 804.600 ;
        RECT 348.450 797.700 350.250 798.000 ;
        RECT 338.550 797.100 350.250 797.700 ;
        RECT 338.550 796.500 356.850 797.100 ;
        RECT 338.550 795.600 339.450 796.500 ;
        RECT 348.450 796.200 356.850 796.500 ;
        RECT 338.550 793.800 340.950 795.600 ;
        RECT 339.150 783.600 340.950 793.800 ;
        RECT 342.150 783.000 343.950 795.600 ;
        RECT 353.250 794.700 355.050 795.300 ;
        RECT 347.250 793.500 355.050 794.700 ;
        RECT 355.950 794.100 356.850 796.200 ;
        RECT 358.950 796.200 359.850 808.800 ;
        RECT 371.250 805.050 372.450 812.400 ;
        RECT 386.400 805.050 387.300 815.400 ;
        RECT 407.700 813.600 409.500 818.400 ;
        RECT 404.400 812.400 409.500 813.600 ;
        RECT 412.200 812.400 414.000 819.000 ;
        RECT 425.100 815.400 426.900 818.400 ;
        RECT 404.400 805.050 405.300 812.400 ;
        RECT 425.100 811.500 426.300 815.400 ;
        RECT 428.100 812.400 429.900 819.000 ;
        RECT 431.100 812.400 432.900 818.400 ;
        RECT 435.150 814.200 436.950 818.400 ;
        RECT 406.950 810.450 409.050 811.050 ;
        RECT 421.950 810.450 424.050 811.050 ;
        RECT 425.100 810.600 430.800 811.500 ;
        RECT 406.950 809.550 424.050 810.450 ;
        RECT 406.950 808.950 409.050 809.550 ;
        RECT 421.950 808.950 424.050 809.550 ;
        RECT 429.000 809.700 430.800 810.600 ;
        RECT 406.950 805.050 408.750 806.850 ;
        RECT 413.100 805.050 414.900 806.850 ;
        RECT 366.150 803.250 372.450 805.050 ;
        RECT 367.950 802.950 372.450 803.250 ;
        RECT 382.950 802.950 385.050 805.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 403.950 802.950 406.050 805.050 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 425.400 802.950 427.500 805.050 ;
        RECT 362.550 800.100 364.650 800.400 ;
        RECT 368.550 800.100 370.350 800.250 ;
        RECT 362.550 798.900 370.350 800.100 ;
        RECT 362.550 798.300 364.650 798.900 ;
        RECT 368.550 798.450 370.350 798.900 ;
        RECT 358.950 795.300 363.750 796.200 ;
        RECT 371.250 795.600 372.450 802.950 ;
        RECT 383.250 801.150 385.050 802.950 ;
        RECT 386.400 795.600 387.300 802.950 ;
        RECT 389.100 801.150 390.900 802.950 ;
        RECT 404.400 795.600 405.300 802.950 ;
        RECT 409.950 801.150 411.750 802.950 ;
        RECT 425.400 801.150 427.200 802.950 ;
        RECT 429.000 798.300 429.900 809.700 ;
        RECT 431.700 805.050 432.900 812.400 ;
        RECT 430.800 802.950 432.900 805.050 ;
        RECT 429.000 797.400 430.800 798.300 ;
        RECT 425.100 796.500 430.800 797.400 ;
        RECT 362.550 794.400 363.750 795.300 ;
        RECT 359.850 794.100 361.650 794.400 ;
        RECT 347.250 792.600 349.350 793.500 ;
        RECT 355.950 793.200 361.650 794.100 ;
        RECT 359.850 792.600 361.650 793.200 ;
        RECT 362.550 792.600 365.550 794.400 ;
        RECT 347.550 783.600 349.350 792.600 ;
        RECT 351.450 791.550 353.250 792.300 ;
        RECT 356.250 791.550 358.050 792.300 ;
        RECT 351.450 790.500 358.050 791.550 ;
        RECT 352.350 783.000 354.150 789.600 ;
        RECT 355.350 783.600 357.150 790.500 ;
        RECT 362.550 789.600 364.650 791.700 ;
        RECT 358.350 783.000 360.150 789.600 ;
        RECT 362.850 783.600 364.650 789.600 ;
        RECT 367.650 783.000 369.450 795.600 ;
        RECT 370.650 783.600 372.450 795.600 ;
        RECT 383.100 783.000 384.900 795.600 ;
        RECT 386.400 794.400 390.000 795.600 ;
        RECT 388.200 783.600 390.000 794.400 ;
        RECT 404.100 783.600 405.900 795.600 ;
        RECT 407.100 794.700 414.900 795.600 ;
        RECT 407.100 783.600 408.900 794.700 ;
        RECT 410.100 783.000 411.900 793.800 ;
        RECT 413.100 783.600 414.900 794.700 ;
        RECT 425.100 789.600 426.300 796.500 ;
        RECT 431.700 795.600 432.900 802.950 ;
        RECT 425.100 783.600 426.900 789.600 ;
        RECT 428.100 783.000 429.900 793.800 ;
        RECT 431.100 783.600 432.900 795.600 ;
        RECT 434.550 812.400 436.950 814.200 ;
        RECT 438.150 812.400 439.950 819.000 ;
        RECT 442.950 816.300 444.750 818.400 ;
        RECT 441.150 815.400 444.750 816.300 ;
        RECT 447.450 815.400 449.250 819.000 ;
        RECT 450.750 815.400 452.550 818.400 ;
        RECT 453.750 815.400 455.550 819.000 ;
        RECT 458.250 815.400 460.050 818.400 ;
        RECT 440.850 814.800 444.750 815.400 ;
        RECT 440.850 813.300 442.950 814.800 ;
        RECT 450.750 814.500 451.800 815.400 ;
        RECT 434.550 797.700 435.450 812.400 ;
        RECT 443.850 811.800 445.650 813.600 ;
        RECT 446.850 813.450 451.800 814.500 ;
        RECT 446.850 812.700 448.650 813.450 ;
        RECT 458.250 813.300 460.650 815.400 ;
        RECT 463.350 812.400 465.150 819.000 ;
        RECT 466.650 812.400 468.450 818.400 ;
        RECT 443.850 810.000 444.900 811.800 ;
        RECT 454.050 810.000 455.850 810.600 ;
        RECT 443.850 808.800 455.850 810.000 ;
        RECT 436.950 807.600 444.900 808.800 ;
        RECT 436.950 805.050 438.750 807.600 ;
        RECT 443.100 807.000 444.900 807.600 ;
        RECT 440.100 805.800 441.900 806.400 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 440.100 804.600 448.200 805.800 ;
        RECT 446.100 802.950 448.200 804.600 ;
        RECT 444.450 797.700 446.250 798.000 ;
        RECT 434.550 797.100 446.250 797.700 ;
        RECT 434.550 796.500 452.850 797.100 ;
        RECT 434.550 795.600 435.450 796.500 ;
        RECT 444.450 796.200 452.850 796.500 ;
        RECT 434.550 793.800 436.950 795.600 ;
        RECT 435.150 783.600 436.950 793.800 ;
        RECT 438.150 783.000 439.950 795.600 ;
        RECT 449.250 794.700 451.050 795.300 ;
        RECT 443.250 793.500 451.050 794.700 ;
        RECT 451.950 794.100 452.850 796.200 ;
        RECT 454.950 796.200 455.850 808.800 ;
        RECT 467.250 805.050 468.450 812.400 ;
        RECT 472.950 811.950 478.050 814.050 ;
        RECT 479.100 813.300 480.900 818.400 ;
        RECT 482.100 814.200 483.900 819.000 ;
        RECT 485.100 813.300 486.900 818.400 ;
        RECT 479.100 811.950 486.900 813.300 ;
        RECT 488.100 812.400 489.900 818.400 ;
        RECT 500.400 812.400 502.200 819.000 ;
        RECT 488.100 810.300 489.300 812.400 ;
        RECT 505.500 811.200 507.300 818.400 ;
        RECT 521.100 815.400 522.900 819.000 ;
        RECT 524.100 815.400 525.900 818.400 ;
        RECT 485.700 809.400 489.300 810.300 ;
        RECT 503.100 810.300 507.300 811.200 ;
        RECT 482.100 805.050 483.900 806.850 ;
        RECT 485.700 805.050 486.900 809.400 ;
        RECT 495.000 807.450 499.050 808.050 ;
        RECT 488.100 805.050 489.900 806.850 ;
        RECT 494.550 805.950 499.050 807.450 ;
        RECT 462.150 803.250 468.450 805.050 ;
        RECT 463.950 802.950 468.450 803.250 ;
        RECT 478.950 802.950 481.050 805.050 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 458.550 800.100 460.650 800.400 ;
        RECT 464.550 800.100 466.350 800.250 ;
        RECT 458.550 798.900 466.350 800.100 ;
        RECT 458.550 798.300 460.650 798.900 ;
        RECT 464.550 798.450 466.350 798.900 ;
        RECT 454.950 795.300 459.750 796.200 ;
        RECT 467.250 795.600 468.450 802.950 ;
        RECT 479.100 801.150 480.900 802.950 ;
        RECT 485.700 795.600 486.900 802.950 ;
        RECT 494.550 801.450 495.450 805.950 ;
        RECT 500.250 805.050 502.050 806.850 ;
        RECT 503.100 805.050 504.300 810.300 ;
        RECT 506.100 805.050 507.900 806.850 ;
        RECT 524.100 805.050 525.300 815.400 ;
        RECT 536.100 812.400 537.900 819.000 ;
        RECT 539.100 811.500 540.900 818.400 ;
        RECT 542.100 812.400 543.900 819.000 ;
        RECT 545.100 811.500 546.900 818.400 ;
        RECT 548.100 812.400 549.900 819.000 ;
        RECT 551.100 811.500 552.900 818.400 ;
        RECT 554.100 812.400 555.900 819.000 ;
        RECT 557.100 811.500 558.900 818.400 ;
        RECT 560.100 812.400 561.900 819.000 ;
        RECT 572.400 812.400 574.200 819.000 ;
        RECT 539.100 810.300 543.000 811.500 ;
        RECT 545.100 810.300 549.000 811.500 ;
        RECT 551.100 810.300 555.000 811.500 ;
        RECT 557.100 810.300 559.950 811.500 ;
        RECT 577.500 811.200 579.300 818.400 ;
        RECT 541.800 809.400 543.000 810.300 ;
        RECT 547.800 809.400 549.000 810.300 ;
        RECT 553.800 809.400 555.000 810.300 ;
        RECT 541.800 808.200 546.000 809.400 ;
        RECT 538.800 805.050 540.600 806.850 ;
        RECT 499.950 802.950 502.050 805.050 ;
        RECT 502.950 802.950 505.050 805.050 ;
        RECT 505.950 802.950 508.050 805.050 ;
        RECT 520.950 802.950 523.050 805.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 538.800 802.950 540.900 805.050 ;
        RECT 491.550 800.550 495.450 801.450 ;
        RECT 491.550 799.050 492.450 800.550 ;
        RECT 487.950 797.550 492.450 799.050 ;
        RECT 487.950 796.950 492.000 797.550 ;
        RECT 458.550 794.400 459.750 795.300 ;
        RECT 455.850 794.100 457.650 794.400 ;
        RECT 443.250 792.600 445.350 793.500 ;
        RECT 451.950 793.200 457.650 794.100 ;
        RECT 455.850 792.600 457.650 793.200 ;
        RECT 458.550 792.600 461.550 794.400 ;
        RECT 443.550 783.600 445.350 792.600 ;
        RECT 447.450 791.550 449.250 792.300 ;
        RECT 452.250 791.550 454.050 792.300 ;
        RECT 447.450 790.500 454.050 791.550 ;
        RECT 448.350 783.000 450.150 789.600 ;
        RECT 451.350 783.600 453.150 790.500 ;
        RECT 458.550 789.600 460.650 791.700 ;
        RECT 454.350 783.000 456.150 789.600 ;
        RECT 458.850 783.600 460.650 789.600 ;
        RECT 463.650 783.000 465.450 795.600 ;
        RECT 466.650 783.600 468.450 795.600 ;
        RECT 479.400 783.000 481.200 795.600 ;
        RECT 484.500 794.100 486.900 795.600 ;
        RECT 484.500 783.600 486.300 794.100 ;
        RECT 487.200 791.100 489.000 792.900 ;
        RECT 503.100 789.600 504.300 802.950 ;
        RECT 521.100 801.150 522.900 802.950 ;
        RECT 524.100 789.600 525.300 802.950 ;
        RECT 541.800 797.700 543.000 808.200 ;
        RECT 544.200 807.600 546.000 808.200 ;
        RECT 547.800 808.200 552.000 809.400 ;
        RECT 547.800 797.700 549.000 808.200 ;
        RECT 550.200 807.600 552.000 808.200 ;
        RECT 553.800 808.200 558.000 809.400 ;
        RECT 553.800 797.700 555.000 808.200 ;
        RECT 556.200 807.600 558.000 808.200 ;
        RECT 558.900 805.050 559.950 810.300 ;
        RECT 575.100 810.300 579.300 811.200 ;
        RECT 581.550 812.400 583.350 818.400 ;
        RECT 584.850 812.400 586.650 819.000 ;
        RECT 589.950 815.400 591.750 818.400 ;
        RECT 594.450 815.400 596.250 819.000 ;
        RECT 597.450 815.400 599.250 818.400 ;
        RECT 600.750 815.400 602.550 819.000 ;
        RECT 605.250 816.300 607.050 818.400 ;
        RECT 605.250 815.400 608.850 816.300 ;
        RECT 589.350 813.300 591.750 815.400 ;
        RECT 598.200 814.500 599.250 815.400 ;
        RECT 605.250 814.800 609.150 815.400 ;
        RECT 598.200 813.450 603.150 814.500 ;
        RECT 601.350 812.700 603.150 813.450 ;
        RECT 572.250 805.050 574.050 806.850 ;
        RECT 575.100 805.050 576.300 810.300 ;
        RECT 578.100 805.050 579.900 806.850 ;
        RECT 581.550 805.050 582.750 812.400 ;
        RECT 604.350 811.800 606.150 813.600 ;
        RECT 607.050 813.300 609.150 814.800 ;
        RECT 610.050 812.400 611.850 819.000 ;
        RECT 613.050 814.200 614.850 818.400 ;
        RECT 626.100 815.400 627.900 818.400 ;
        RECT 629.100 815.400 630.900 819.000 ;
        RECT 613.050 812.400 615.450 814.200 ;
        RECT 594.150 810.000 595.950 810.600 ;
        RECT 605.100 810.000 606.150 811.800 ;
        RECT 594.150 808.800 606.150 810.000 ;
        RECT 556.800 802.950 559.950 805.050 ;
        RECT 571.950 802.950 574.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 581.550 803.250 587.850 805.050 ;
        RECT 581.550 802.950 586.050 803.250 ;
        RECT 558.900 797.700 559.950 802.950 ;
        RECT 539.100 796.500 543.000 797.700 ;
        RECT 545.100 796.500 549.000 797.700 ;
        RECT 551.100 796.500 555.000 797.700 ;
        RECT 557.100 796.500 559.950 797.700 ;
        RECT 487.500 783.000 489.300 789.600 ;
        RECT 500.100 783.000 501.900 789.600 ;
        RECT 503.100 783.600 504.900 789.600 ;
        RECT 506.100 783.000 507.900 789.600 ;
        RECT 521.100 783.000 522.900 789.600 ;
        RECT 524.100 783.600 525.900 789.600 ;
        RECT 536.100 783.000 537.900 795.600 ;
        RECT 539.100 783.600 540.900 796.500 ;
        RECT 542.100 783.000 543.900 795.600 ;
        RECT 545.100 783.600 546.900 796.500 ;
        RECT 548.100 783.000 549.900 795.600 ;
        RECT 551.100 783.600 552.900 796.500 ;
        RECT 554.100 783.000 555.900 795.600 ;
        RECT 557.100 783.600 558.900 796.500 ;
        RECT 560.100 783.000 561.900 795.600 ;
        RECT 575.100 789.600 576.300 802.950 ;
        RECT 581.550 795.600 582.750 802.950 ;
        RECT 583.650 800.100 585.450 800.250 ;
        RECT 589.350 800.100 591.450 800.400 ;
        RECT 583.650 798.900 591.450 800.100 ;
        RECT 583.650 798.450 585.450 798.900 ;
        RECT 589.350 798.300 591.450 798.900 ;
        RECT 594.150 796.200 595.050 808.800 ;
        RECT 605.100 807.600 613.050 808.800 ;
        RECT 605.100 807.000 606.900 807.600 ;
        RECT 608.100 805.800 609.900 806.400 ;
        RECT 601.800 804.600 609.900 805.800 ;
        RECT 611.250 805.050 613.050 807.600 ;
        RECT 601.800 802.950 603.900 804.600 ;
        RECT 610.950 802.950 613.050 805.050 ;
        RECT 603.750 797.700 605.550 798.000 ;
        RECT 614.550 797.700 615.450 812.400 ;
        RECT 626.700 805.050 627.900 815.400 ;
        RECT 632.550 812.400 634.350 818.400 ;
        RECT 635.850 812.400 637.650 819.000 ;
        RECT 640.950 815.400 642.750 818.400 ;
        RECT 645.450 815.400 647.250 819.000 ;
        RECT 648.450 815.400 650.250 818.400 ;
        RECT 651.750 815.400 653.550 819.000 ;
        RECT 656.250 816.300 658.050 818.400 ;
        RECT 656.250 815.400 659.850 816.300 ;
        RECT 640.350 813.300 642.750 815.400 ;
        RECT 649.200 814.500 650.250 815.400 ;
        RECT 656.250 814.800 660.150 815.400 ;
        RECT 649.200 813.450 654.150 814.500 ;
        RECT 652.350 812.700 654.150 813.450 ;
        RECT 632.550 805.050 633.750 812.400 ;
        RECT 655.350 811.800 657.150 813.600 ;
        RECT 658.050 813.300 660.150 814.800 ;
        RECT 661.050 812.400 662.850 819.000 ;
        RECT 664.050 814.200 665.850 818.400 ;
        RECT 677.100 815.400 678.900 818.400 ;
        RECT 680.100 815.400 681.900 819.000 ;
        RECT 692.100 815.400 693.900 818.400 ;
        RECT 695.100 815.400 696.900 819.000 ;
        RECT 664.050 812.400 666.450 814.200 ;
        RECT 645.150 810.000 646.950 810.600 ;
        RECT 656.100 810.000 657.150 811.800 ;
        RECT 645.150 808.800 657.150 810.000 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 632.550 803.250 638.850 805.050 ;
        RECT 632.550 802.950 637.050 803.250 ;
        RECT 603.750 797.100 615.450 797.700 ;
        RECT 572.100 783.000 573.900 789.600 ;
        RECT 575.100 783.600 576.900 789.600 ;
        RECT 578.100 783.000 579.900 789.600 ;
        RECT 581.550 783.600 583.350 795.600 ;
        RECT 584.550 783.000 586.350 795.600 ;
        RECT 590.250 795.300 595.050 796.200 ;
        RECT 597.150 796.500 615.450 797.100 ;
        RECT 597.150 796.200 605.550 796.500 ;
        RECT 590.250 794.400 591.450 795.300 ;
        RECT 588.450 792.600 591.450 794.400 ;
        RECT 592.350 794.100 594.150 794.400 ;
        RECT 597.150 794.100 598.050 796.200 ;
        RECT 614.550 795.600 615.450 796.500 ;
        RECT 592.350 793.200 598.050 794.100 ;
        RECT 598.950 794.700 600.750 795.300 ;
        RECT 598.950 793.500 606.750 794.700 ;
        RECT 592.350 792.600 594.150 793.200 ;
        RECT 604.650 792.600 606.750 793.500 ;
        RECT 589.350 789.600 591.450 791.700 ;
        RECT 595.950 791.550 597.750 792.300 ;
        RECT 600.750 791.550 602.550 792.300 ;
        RECT 595.950 790.500 602.550 791.550 ;
        RECT 589.350 783.600 591.150 789.600 ;
        RECT 593.850 783.000 595.650 789.600 ;
        RECT 596.850 783.600 598.650 790.500 ;
        RECT 599.850 783.000 601.650 789.600 ;
        RECT 604.650 783.600 606.450 792.600 ;
        RECT 610.050 783.000 611.850 795.600 ;
        RECT 613.050 793.800 615.450 795.600 ;
        RECT 613.050 783.600 614.850 793.800 ;
        RECT 626.700 789.600 627.900 802.950 ;
        RECT 629.100 801.150 630.900 802.950 ;
        RECT 632.550 795.600 633.750 802.950 ;
        RECT 634.650 800.100 636.450 800.250 ;
        RECT 640.350 800.100 642.450 800.400 ;
        RECT 634.650 798.900 642.450 800.100 ;
        RECT 634.650 798.450 636.450 798.900 ;
        RECT 640.350 798.300 642.450 798.900 ;
        RECT 645.150 796.200 646.050 808.800 ;
        RECT 656.100 807.600 664.050 808.800 ;
        RECT 656.100 807.000 657.900 807.600 ;
        RECT 659.100 805.800 660.900 806.400 ;
        RECT 652.800 804.600 660.900 805.800 ;
        RECT 662.250 805.050 664.050 807.600 ;
        RECT 652.800 802.950 654.900 804.600 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 654.750 797.700 656.550 798.000 ;
        RECT 665.550 797.700 666.450 812.400 ;
        RECT 677.700 805.050 678.900 815.400 ;
        RECT 692.700 805.050 693.900 815.400 ;
        RECT 707.700 812.400 709.500 819.000 ;
        RECT 712.200 812.400 714.000 818.400 ;
        RECT 716.700 812.400 718.500 819.000 ;
        RECT 731.700 815.400 733.500 819.000 ;
        RECT 734.700 813.600 736.500 818.400 ;
        RECT 731.400 812.400 736.500 813.600 ;
        RECT 739.200 812.400 741.000 819.000 ;
        RECT 755.100 818.400 756.300 819.000 ;
        RECT 755.100 815.400 756.900 818.400 ;
        RECT 758.100 815.400 759.900 818.400 ;
        RECT 707.250 805.050 709.050 806.850 ;
        RECT 713.100 805.050 714.300 812.400 ;
        RECT 719.100 805.050 720.900 806.850 ;
        RECT 731.400 805.050 732.300 812.400 ;
        RECT 758.400 811.200 759.300 815.400 ;
        RECT 761.100 813.000 762.900 819.000 ;
        RECT 764.100 812.400 765.900 818.400 ;
        RECT 758.400 810.300 763.800 811.200 ;
        RECT 761.700 809.400 763.800 810.300 ;
        RECT 733.950 805.050 735.750 806.850 ;
        RECT 740.100 805.050 741.900 806.850 ;
        RECT 755.400 805.050 757.200 806.850 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 694.950 802.950 697.050 805.050 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 736.950 802.950 739.050 805.050 ;
        RECT 739.950 802.950 742.050 805.050 ;
        RECT 755.100 802.950 757.200 805.050 ;
        RECT 758.400 802.950 760.500 805.050 ;
        RECT 654.750 797.100 666.450 797.700 ;
        RECT 626.100 783.600 627.900 789.600 ;
        RECT 629.100 783.000 630.900 789.600 ;
        RECT 632.550 783.600 634.350 795.600 ;
        RECT 635.550 783.000 637.350 795.600 ;
        RECT 641.250 795.300 646.050 796.200 ;
        RECT 648.150 796.500 666.450 797.100 ;
        RECT 648.150 796.200 656.550 796.500 ;
        RECT 641.250 794.400 642.450 795.300 ;
        RECT 639.450 792.600 642.450 794.400 ;
        RECT 643.350 794.100 645.150 794.400 ;
        RECT 648.150 794.100 649.050 796.200 ;
        RECT 665.550 795.600 666.450 796.500 ;
        RECT 643.350 793.200 649.050 794.100 ;
        RECT 649.950 794.700 651.750 795.300 ;
        RECT 649.950 793.500 657.750 794.700 ;
        RECT 643.350 792.600 645.150 793.200 ;
        RECT 655.650 792.600 657.750 793.500 ;
        RECT 640.350 789.600 642.450 791.700 ;
        RECT 646.950 791.550 648.750 792.300 ;
        RECT 651.750 791.550 653.550 792.300 ;
        RECT 646.950 790.500 653.550 791.550 ;
        RECT 640.350 783.600 642.150 789.600 ;
        RECT 644.850 783.000 646.650 789.600 ;
        RECT 647.850 783.600 649.650 790.500 ;
        RECT 650.850 783.000 652.650 789.600 ;
        RECT 655.650 783.600 657.450 792.600 ;
        RECT 661.050 783.000 662.850 795.600 ;
        RECT 664.050 793.800 666.450 795.600 ;
        RECT 664.050 783.600 665.850 793.800 ;
        RECT 677.700 789.600 678.900 802.950 ;
        RECT 680.100 801.150 681.900 802.950 ;
        RECT 692.700 789.600 693.900 802.950 ;
        RECT 695.100 801.150 696.900 802.950 ;
        RECT 710.250 801.150 712.050 802.950 ;
        RECT 713.100 797.400 714.000 802.950 ;
        RECT 716.100 801.150 717.900 802.950 ;
        RECT 713.100 796.500 717.900 797.400 ;
        RECT 707.100 794.400 714.900 795.300 ;
        RECT 677.100 783.600 678.900 789.600 ;
        RECT 680.100 783.000 681.900 789.600 ;
        RECT 692.100 783.600 693.900 789.600 ;
        RECT 695.100 783.000 696.900 789.600 ;
        RECT 707.100 783.600 708.900 794.400 ;
        RECT 710.100 783.000 711.900 793.500 ;
        RECT 713.100 784.500 714.900 794.400 ;
        RECT 716.100 785.400 717.900 796.500 ;
        RECT 731.400 795.600 732.300 802.950 ;
        RECT 736.950 801.150 738.750 802.950 ;
        RECT 759.000 801.150 760.800 802.950 ;
        RECT 761.700 798.900 762.600 809.400 ;
        RECT 765.000 805.050 765.900 812.400 ;
        RECT 776.100 813.300 777.900 818.400 ;
        RECT 779.100 814.200 780.900 819.000 ;
        RECT 782.100 813.300 783.900 818.400 ;
        RECT 776.100 811.950 783.900 813.300 ;
        RECT 785.100 812.400 786.900 818.400 ;
        RECT 797.100 815.400 798.900 818.400 ;
        RECT 800.100 815.400 801.900 819.000 ;
        RECT 785.100 810.300 786.300 812.400 ;
        RECT 782.700 809.400 786.300 810.300 ;
        RECT 779.100 805.050 780.900 806.850 ;
        RECT 782.700 805.050 783.900 809.400 ;
        RECT 785.100 805.050 786.900 806.850 ;
        RECT 797.700 805.050 798.900 815.400 ;
        RECT 812.100 810.600 813.900 818.400 ;
        RECT 816.600 812.400 818.400 819.000 ;
        RECT 819.600 814.200 821.400 818.400 ;
        RECT 833.100 815.400 834.900 819.000 ;
        RECT 836.100 815.400 837.900 818.400 ;
        RECT 839.100 815.400 840.900 819.000 ;
        RECT 819.600 812.400 822.300 814.200 ;
        RECT 818.700 810.600 820.500 811.500 ;
        RECT 812.100 809.700 820.500 810.600 ;
        RECT 812.250 805.050 814.050 806.850 ;
        RECT 763.800 802.950 765.900 805.050 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 796.950 802.950 799.050 805.050 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 812.100 802.950 814.200 805.050 ;
        RECT 761.100 798.300 762.900 798.900 ;
        RECT 755.100 797.100 762.900 798.300 ;
        RECT 755.100 795.600 756.300 797.100 ;
        RECT 763.800 795.600 765.000 802.950 ;
        RECT 776.100 801.150 777.900 802.950 ;
        RECT 782.700 795.600 783.900 802.950 ;
        RECT 719.100 784.500 720.900 795.600 ;
        RECT 713.100 783.600 720.900 784.500 ;
        RECT 731.100 783.600 732.900 795.600 ;
        RECT 734.100 794.700 741.900 795.600 ;
        RECT 734.100 783.600 735.900 794.700 ;
        RECT 737.100 783.000 738.900 793.800 ;
        RECT 740.100 783.600 741.900 794.700 ;
        RECT 755.100 783.600 756.900 795.600 ;
        RECT 759.600 783.000 761.400 795.600 ;
        RECT 762.600 794.100 765.000 795.600 ;
        RECT 762.600 783.600 764.400 794.100 ;
        RECT 776.400 783.000 778.200 795.600 ;
        RECT 781.500 794.100 783.900 795.600 ;
        RECT 781.500 783.600 783.300 794.100 ;
        RECT 784.200 791.100 786.000 792.900 ;
        RECT 797.700 789.600 798.900 802.950 ;
        RECT 800.100 801.150 801.900 802.950 ;
        RECT 799.950 798.450 802.050 799.050 ;
        RECT 811.950 798.450 814.050 799.050 ;
        RECT 799.950 797.550 814.050 798.450 ;
        RECT 799.950 796.950 802.050 797.550 ;
        RECT 811.950 796.950 814.050 797.550 ;
        RECT 815.100 789.600 816.000 809.700 ;
        RECT 821.400 805.050 822.300 812.400 ;
        RECT 836.400 805.050 837.300 815.400 ;
        RECT 851.700 811.200 853.500 818.400 ;
        RECT 856.800 812.400 858.600 819.000 ;
        RECT 851.700 810.300 855.900 811.200 ;
        RECT 851.100 805.050 852.900 806.850 ;
        RECT 854.700 805.050 855.900 810.300 ;
        RECT 856.950 805.050 858.750 806.850 ;
        RECT 817.500 802.950 819.600 805.050 ;
        RECT 820.800 802.950 822.900 805.050 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 856.950 802.950 859.050 805.050 ;
        RECT 817.200 801.150 819.000 802.950 ;
        RECT 821.400 795.600 822.300 802.950 ;
        RECT 833.250 801.150 835.050 802.950 ;
        RECT 836.400 795.600 837.300 802.950 ;
        RECT 839.100 801.150 840.900 802.950 ;
        RECT 784.500 783.000 786.300 789.600 ;
        RECT 797.100 783.600 798.900 789.600 ;
        RECT 800.100 783.000 801.900 789.600 ;
        RECT 812.100 783.000 813.900 789.600 ;
        RECT 815.100 783.600 816.900 789.600 ;
        RECT 818.100 783.000 819.900 795.000 ;
        RECT 821.100 783.600 822.900 795.600 ;
        RECT 833.100 783.000 834.900 795.600 ;
        RECT 836.400 794.400 840.000 795.600 ;
        RECT 838.200 783.600 840.000 794.400 ;
        RECT 854.700 789.600 855.900 802.950 ;
        RECT 851.100 783.000 852.900 789.600 ;
        RECT 854.100 783.600 855.900 789.600 ;
        RECT 857.100 783.000 858.900 789.600 ;
        RECT 14.400 767.400 16.200 780.000 ;
        RECT 19.500 768.900 21.300 779.400 ;
        RECT 22.500 773.400 24.300 780.000 ;
        RECT 35.100 773.400 36.900 780.000 ;
        RECT 38.100 773.400 39.900 779.400 ;
        RECT 41.100 773.400 42.900 780.000 ;
        RECT 22.200 770.100 24.000 771.900 ;
        RECT 19.500 767.400 21.900 768.900 ;
        RECT 9.000 762.450 13.050 763.050 ;
        RECT 8.550 760.950 13.050 762.450 ;
        RECT 8.550 757.050 9.450 760.950 ;
        RECT 14.100 760.050 15.900 761.850 ;
        RECT 20.700 760.050 21.900 767.400 ;
        RECT 38.700 760.050 39.900 773.400 ;
        RECT 56.100 767.400 57.900 780.000 ;
        RECT 61.200 768.600 63.000 779.400 ;
        RECT 59.400 767.400 63.000 768.600 ;
        RECT 74.400 767.400 76.200 780.000 ;
        RECT 79.500 768.900 81.300 779.400 ;
        RECT 82.500 773.400 84.300 780.000 ;
        RECT 82.200 770.100 84.000 771.900 ;
        RECT 87.150 769.200 88.950 779.400 ;
        RECT 79.500 767.400 81.900 768.900 ;
        RECT 56.250 760.050 58.050 761.850 ;
        RECT 59.400 760.050 60.300 767.400 ;
        RECT 62.100 760.050 63.900 761.850 ;
        RECT 74.100 760.050 75.900 761.850 ;
        RECT 80.700 760.050 81.900 767.400 ;
        RECT 86.550 767.400 88.950 769.200 ;
        RECT 90.150 767.400 91.950 780.000 ;
        RECT 95.550 770.400 97.350 779.400 ;
        RECT 100.350 773.400 102.150 780.000 ;
        RECT 103.350 772.500 105.150 779.400 ;
        RECT 106.350 773.400 108.150 780.000 ;
        RECT 110.850 773.400 112.650 779.400 ;
        RECT 99.450 771.450 106.050 772.500 ;
        RECT 99.450 770.700 101.250 771.450 ;
        RECT 104.250 770.700 106.050 771.450 ;
        RECT 110.550 771.300 112.650 773.400 ;
        RECT 95.250 769.500 97.350 770.400 ;
        RECT 107.850 769.800 109.650 770.400 ;
        RECT 95.250 768.300 103.050 769.500 ;
        RECT 101.250 767.700 103.050 768.300 ;
        RECT 103.950 768.900 109.650 769.800 ;
        RECT 86.550 766.500 87.450 767.400 ;
        RECT 103.950 766.800 104.850 768.900 ;
        RECT 107.850 768.600 109.650 768.900 ;
        RECT 110.550 768.600 113.550 770.400 ;
        RECT 110.550 767.700 111.750 768.600 ;
        RECT 96.450 766.500 104.850 766.800 ;
        RECT 86.550 765.900 104.850 766.500 ;
        RECT 106.950 766.800 111.750 767.700 ;
        RECT 115.650 767.400 117.450 780.000 ;
        RECT 118.650 767.400 120.450 779.400 ;
        RECT 131.100 773.400 132.900 780.000 ;
        RECT 134.100 773.400 135.900 779.400 ;
        RECT 137.100 773.400 138.900 780.000 ;
        RECT 149.100 778.500 156.900 779.400 ;
        RECT 86.550 765.300 98.250 765.900 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 22.950 757.950 25.050 760.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 73.950 757.950 76.050 760.050 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 8.550 755.550 13.050 757.050 ;
        RECT 17.100 756.150 18.900 757.950 ;
        RECT 9.000 754.950 13.050 755.550 ;
        RECT 20.700 753.600 21.900 757.950 ;
        RECT 23.100 756.150 24.900 757.950 ;
        RECT 35.100 756.150 36.900 757.950 ;
        RECT 20.700 752.700 24.300 753.600 ;
        RECT 38.700 752.700 39.900 757.950 ;
        RECT 40.950 756.150 42.750 757.950 ;
        RECT 14.100 749.700 21.900 751.050 ;
        RECT 14.100 744.600 15.900 749.700 ;
        RECT 17.100 744.000 18.900 748.800 ;
        RECT 20.100 744.600 21.900 749.700 ;
        RECT 23.100 750.600 24.300 752.700 ;
        RECT 35.700 751.800 39.900 752.700 ;
        RECT 23.100 744.600 24.900 750.600 ;
        RECT 35.700 744.600 37.500 751.800 ;
        RECT 40.800 744.000 42.600 750.600 ;
        RECT 59.400 747.600 60.300 757.950 ;
        RECT 77.100 756.150 78.900 757.950 ;
        RECT 80.700 753.600 81.900 757.950 ;
        RECT 83.100 756.150 84.900 757.950 ;
        RECT 80.700 752.700 84.300 753.600 ;
        RECT 74.100 749.700 81.900 751.050 ;
        RECT 56.100 744.000 57.900 747.600 ;
        RECT 59.100 744.600 60.900 747.600 ;
        RECT 62.100 744.000 63.900 747.600 ;
        RECT 74.100 744.600 75.900 749.700 ;
        RECT 77.100 744.000 78.900 748.800 ;
        RECT 80.100 744.600 81.900 749.700 ;
        RECT 83.100 750.600 84.300 752.700 ;
        RECT 86.550 750.600 87.450 765.300 ;
        RECT 96.450 765.000 98.250 765.300 ;
        RECT 88.950 757.950 91.050 760.050 ;
        RECT 98.100 758.400 100.200 760.050 ;
        RECT 88.950 755.400 90.750 757.950 ;
        RECT 92.100 757.200 100.200 758.400 ;
        RECT 92.100 756.600 93.900 757.200 ;
        RECT 95.100 755.400 96.900 756.000 ;
        RECT 88.950 754.200 96.900 755.400 ;
        RECT 106.950 754.200 107.850 766.800 ;
        RECT 110.550 764.100 112.650 764.700 ;
        RECT 116.550 764.100 118.350 764.550 ;
        RECT 110.550 762.900 118.350 764.100 ;
        RECT 110.550 762.600 112.650 762.900 ;
        RECT 116.550 762.750 118.350 762.900 ;
        RECT 119.250 760.050 120.450 767.400 ;
        RECT 134.100 760.050 135.300 773.400 ;
        RECT 149.100 767.400 150.900 778.500 ;
        RECT 152.100 766.500 153.900 777.600 ;
        RECT 155.100 768.600 156.900 778.500 ;
        RECT 158.100 769.500 159.900 780.000 ;
        RECT 161.100 768.600 162.900 779.400 ;
        RECT 155.100 767.700 162.900 768.600 ;
        RECT 176.100 778.500 183.900 779.400 ;
        RECT 176.100 767.400 177.900 778.500 ;
        RECT 179.100 766.500 180.900 777.600 ;
        RECT 182.100 768.600 183.900 778.500 ;
        RECT 185.100 769.500 186.900 780.000 ;
        RECT 188.100 768.600 189.900 779.400 ;
        RECT 192.150 769.200 193.950 779.400 ;
        RECT 182.100 767.700 189.900 768.600 ;
        RECT 191.550 767.400 193.950 769.200 ;
        RECT 195.150 767.400 196.950 780.000 ;
        RECT 200.550 770.400 202.350 779.400 ;
        RECT 205.350 773.400 207.150 780.000 ;
        RECT 208.350 772.500 210.150 779.400 ;
        RECT 211.350 773.400 213.150 780.000 ;
        RECT 215.850 773.400 217.650 779.400 ;
        RECT 204.450 771.450 211.050 772.500 ;
        RECT 204.450 770.700 206.250 771.450 ;
        RECT 209.250 770.700 211.050 771.450 ;
        RECT 215.550 771.300 217.650 773.400 ;
        RECT 200.250 769.500 202.350 770.400 ;
        RECT 212.850 769.800 214.650 770.400 ;
        RECT 200.250 768.300 208.050 769.500 ;
        RECT 206.250 767.700 208.050 768.300 ;
        RECT 208.950 768.900 214.650 769.800 ;
        RECT 191.550 766.500 192.450 767.400 ;
        RECT 208.950 766.800 209.850 768.900 ;
        RECT 212.850 768.600 214.650 768.900 ;
        RECT 215.550 768.600 218.550 770.400 ;
        RECT 215.550 767.700 216.750 768.600 ;
        RECT 201.450 766.500 209.850 766.800 ;
        RECT 152.100 765.600 156.900 766.500 ;
        RECT 179.100 765.600 183.900 766.500 ;
        RECT 152.100 760.050 153.900 761.850 ;
        RECT 156.000 760.050 156.900 765.600 ;
        RECT 157.950 760.050 159.750 761.850 ;
        RECT 179.100 760.050 180.900 761.850 ;
        RECT 183.000 760.050 183.900 765.600 ;
        RECT 191.550 765.900 209.850 766.500 ;
        RECT 211.950 766.800 216.750 767.700 ;
        RECT 220.650 767.400 222.450 780.000 ;
        RECT 223.650 767.400 225.450 779.400 ;
        RECT 236.700 773.400 238.500 780.000 ;
        RECT 237.000 770.100 238.800 771.900 ;
        RECT 239.700 768.900 241.500 779.400 ;
        RECT 191.550 765.300 203.250 765.900 ;
        RECT 184.950 760.050 186.750 761.850 ;
        RECT 115.950 759.750 120.450 760.050 ;
        RECT 114.150 757.950 120.450 759.750 ;
        RECT 130.950 757.950 133.050 760.050 ;
        RECT 133.950 757.950 136.050 760.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 154.950 757.950 157.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 178.950 757.950 181.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 95.850 753.000 107.850 754.200 ;
        RECT 95.850 751.200 96.900 753.000 ;
        RECT 106.050 752.400 107.850 753.000 ;
        RECT 83.100 744.600 84.900 750.600 ;
        RECT 86.550 748.800 88.950 750.600 ;
        RECT 87.150 744.600 88.950 748.800 ;
        RECT 90.150 744.000 91.950 750.600 ;
        RECT 92.850 748.200 94.950 749.700 ;
        RECT 95.850 749.400 97.650 751.200 ;
        RECT 119.250 750.600 120.450 757.950 ;
        RECT 131.250 756.150 133.050 757.950 ;
        RECT 134.100 752.700 135.300 757.950 ;
        RECT 137.100 756.150 138.900 757.950 ;
        RECT 149.100 756.150 150.900 757.950 ;
        RECT 134.100 751.800 138.300 752.700 ;
        RECT 98.850 749.550 100.650 750.300 ;
        RECT 98.850 748.500 103.800 749.550 ;
        RECT 92.850 747.600 96.750 748.200 ;
        RECT 102.750 747.600 103.800 748.500 ;
        RECT 110.250 747.600 112.650 749.700 ;
        RECT 93.150 746.700 96.750 747.600 ;
        RECT 94.950 744.600 96.750 746.700 ;
        RECT 99.450 744.000 101.250 747.600 ;
        RECT 102.750 744.600 104.550 747.600 ;
        RECT 105.750 744.000 107.550 747.600 ;
        RECT 110.250 744.600 112.050 747.600 ;
        RECT 115.350 744.000 117.150 750.600 ;
        RECT 118.650 744.600 120.450 750.600 ;
        RECT 131.400 744.000 133.200 750.600 ;
        RECT 136.500 744.600 138.300 751.800 ;
        RECT 155.700 750.600 156.900 757.950 ;
        RECT 160.950 756.150 162.750 757.950 ;
        RECT 176.100 756.150 177.900 757.950 ;
        RECT 182.700 750.600 183.900 757.950 ;
        RECT 187.950 756.150 189.750 757.950 ;
        RECT 191.550 750.600 192.450 765.300 ;
        RECT 201.450 765.000 203.250 765.300 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 203.100 758.400 205.200 760.050 ;
        RECT 193.950 755.400 195.750 757.950 ;
        RECT 197.100 757.200 205.200 758.400 ;
        RECT 197.100 756.600 198.900 757.200 ;
        RECT 200.100 755.400 201.900 756.000 ;
        RECT 193.950 754.200 201.900 755.400 ;
        RECT 211.950 754.200 212.850 766.800 ;
        RECT 215.550 764.100 217.650 764.700 ;
        RECT 221.550 764.100 223.350 764.550 ;
        RECT 215.550 762.900 223.350 764.100 ;
        RECT 215.550 762.600 217.650 762.900 ;
        RECT 221.550 762.750 223.350 762.900 ;
        RECT 224.250 760.050 225.450 767.400 ;
        RECT 239.100 767.400 241.500 768.900 ;
        RECT 244.800 767.400 246.600 780.000 ;
        RECT 257.100 773.400 258.900 780.000 ;
        RECT 260.100 773.400 261.900 779.400 ;
        RECT 263.100 773.400 264.900 780.000 ;
        RECT 239.100 760.050 240.300 767.400 ;
        RECT 247.950 762.450 250.050 766.050 ;
        RECT 247.950 762.000 252.450 762.450 ;
        RECT 245.100 760.050 246.900 761.850 ;
        RECT 248.550 761.550 252.450 762.000 ;
        RECT 220.950 759.750 225.450 760.050 ;
        RECT 219.150 757.950 225.450 759.750 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 200.850 753.000 212.850 754.200 ;
        RECT 200.850 751.200 201.900 753.000 ;
        RECT 211.050 752.400 212.850 753.000 ;
        RECT 151.500 744.000 153.300 750.600 ;
        RECT 156.000 744.600 157.800 750.600 ;
        RECT 160.500 744.000 162.300 750.600 ;
        RECT 178.500 744.000 180.300 750.600 ;
        RECT 183.000 744.600 184.800 750.600 ;
        RECT 187.500 744.000 189.300 750.600 ;
        RECT 191.550 748.800 193.950 750.600 ;
        RECT 192.150 744.600 193.950 748.800 ;
        RECT 195.150 744.000 196.950 750.600 ;
        RECT 197.850 748.200 199.950 749.700 ;
        RECT 200.850 749.400 202.650 751.200 ;
        RECT 224.250 750.600 225.450 757.950 ;
        RECT 236.100 756.150 237.900 757.950 ;
        RECT 239.100 753.600 240.300 757.950 ;
        RECT 242.100 756.150 243.900 757.950 ;
        RECT 251.550 756.450 252.450 761.550 ;
        RECT 260.700 760.050 261.900 773.400 ;
        RECT 276.000 768.600 277.800 779.400 ;
        RECT 276.000 767.400 279.600 768.600 ;
        RECT 281.100 767.400 282.900 780.000 ;
        RECT 293.100 773.400 294.900 780.000 ;
        RECT 296.100 773.400 297.900 779.400 ;
        RECT 275.100 760.050 276.900 761.850 ;
        RECT 278.700 760.050 279.600 767.400 ;
        RECT 280.950 760.050 282.750 761.850 ;
        RECT 286.950 760.950 289.050 763.050 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 251.550 756.000 255.450 756.450 ;
        RECT 257.100 756.150 258.900 757.950 ;
        RECT 251.550 755.550 256.050 756.000 ;
        RECT 236.700 752.700 240.300 753.600 ;
        RECT 236.700 750.600 237.900 752.700 ;
        RECT 253.950 751.950 256.050 755.550 ;
        RECT 260.700 752.700 261.900 757.950 ;
        RECT 262.950 756.150 264.750 757.950 ;
        RECT 257.700 751.800 261.900 752.700 ;
        RECT 203.850 749.550 205.650 750.300 ;
        RECT 203.850 748.500 208.800 749.550 ;
        RECT 197.850 747.600 201.750 748.200 ;
        RECT 207.750 747.600 208.800 748.500 ;
        RECT 215.250 747.600 217.650 749.700 ;
        RECT 198.150 746.700 201.750 747.600 ;
        RECT 199.950 744.600 201.750 746.700 ;
        RECT 204.450 744.000 206.250 747.600 ;
        RECT 207.750 744.600 209.550 747.600 ;
        RECT 210.750 744.000 212.550 747.600 ;
        RECT 215.250 744.600 217.050 747.600 ;
        RECT 220.350 744.000 222.150 750.600 ;
        RECT 223.650 744.600 225.450 750.600 ;
        RECT 236.100 744.600 237.900 750.600 ;
        RECT 239.100 749.700 246.900 751.050 ;
        RECT 239.100 744.600 240.900 749.700 ;
        RECT 242.100 744.000 243.900 748.800 ;
        RECT 245.100 744.600 246.900 749.700 ;
        RECT 257.700 744.600 259.500 751.800 ;
        RECT 262.800 744.000 264.600 750.600 ;
        RECT 278.700 747.600 279.600 757.950 ;
        RECT 287.550 757.050 288.450 760.950 ;
        RECT 293.100 760.050 294.900 761.850 ;
        RECT 296.100 760.050 297.300 773.400 ;
        RECT 311.100 767.400 312.900 779.400 ;
        RECT 314.100 769.200 315.900 780.000 ;
        RECT 317.100 773.400 318.900 779.400 ;
        RECT 329.700 773.400 331.500 780.000 ;
        RECT 311.100 760.050 312.300 767.400 ;
        RECT 317.700 766.500 318.900 773.400 ;
        RECT 330.000 770.100 331.800 771.900 ;
        RECT 332.700 768.900 334.500 779.400 ;
        RECT 313.200 765.600 318.900 766.500 ;
        RECT 332.100 767.400 334.500 768.900 ;
        RECT 337.800 767.400 339.600 780.000 ;
        RECT 350.700 773.400 352.500 780.000 ;
        RECT 351.000 770.100 352.800 771.900 ;
        RECT 353.700 768.900 355.500 779.400 ;
        RECT 353.100 767.400 355.500 768.900 ;
        RECT 358.800 767.400 360.600 780.000 ;
        RECT 372.000 768.600 373.800 779.400 ;
        RECT 372.000 767.400 375.600 768.600 ;
        RECT 377.100 767.400 378.900 780.000 ;
        RECT 389.700 773.400 391.500 780.000 ;
        RECT 390.000 770.100 391.800 771.900 ;
        RECT 392.700 768.900 394.500 779.400 ;
        RECT 392.100 767.400 394.500 768.900 ;
        RECT 397.800 767.400 399.600 780.000 ;
        RECT 410.100 767.400 411.900 780.000 ;
        RECT 415.200 768.600 417.000 779.400 ;
        RECT 413.400 767.400 417.000 768.600 ;
        RECT 428.100 767.400 429.900 779.400 ;
        RECT 431.100 769.200 432.900 780.000 ;
        RECT 434.100 773.400 435.900 779.400 ;
        RECT 313.200 764.700 315.000 765.600 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 311.100 757.950 313.200 760.050 ;
        RECT 283.950 754.950 292.050 757.050 ;
        RECT 296.100 747.600 297.300 757.950 ;
        RECT 311.100 750.600 312.300 757.950 ;
        RECT 314.100 753.300 315.000 764.700 ;
        RECT 316.800 760.050 318.600 761.850 ;
        RECT 332.100 760.050 333.300 767.400 ;
        RECT 338.100 760.050 339.900 761.850 ;
        RECT 353.100 760.050 354.300 767.400 ;
        RECT 359.100 760.050 360.900 761.850 ;
        RECT 371.100 760.050 372.900 761.850 ;
        RECT 374.700 760.050 375.600 767.400 ;
        RECT 376.950 760.050 378.750 761.850 ;
        RECT 392.100 760.050 393.300 767.400 ;
        RECT 398.100 760.050 399.900 761.850 ;
        RECT 410.250 760.050 412.050 761.850 ;
        RECT 413.400 760.050 414.300 767.400 ;
        RECT 416.100 760.050 417.900 761.850 ;
        RECT 428.100 760.050 429.300 767.400 ;
        RECT 434.700 766.500 435.900 773.400 ;
        RECT 446.400 767.400 448.200 780.000 ;
        RECT 451.500 768.900 453.300 779.400 ;
        RECT 454.500 773.400 456.300 780.000 ;
        RECT 467.100 773.400 468.900 780.000 ;
        RECT 470.100 773.400 471.900 779.400 ;
        RECT 473.100 773.400 474.900 780.000 ;
        RECT 454.200 770.100 456.000 771.900 ;
        RECT 451.500 767.400 453.900 768.900 ;
        RECT 430.200 765.600 435.900 766.500 ;
        RECT 430.200 764.700 432.000 765.600 ;
        RECT 316.500 757.950 318.600 760.050 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 355.950 757.950 358.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 391.950 757.950 394.050 760.050 ;
        RECT 394.950 757.950 397.050 760.050 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 412.950 757.950 415.050 760.050 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 428.100 757.950 430.200 760.050 ;
        RECT 329.100 756.150 330.900 757.950 ;
        RECT 332.100 753.600 333.300 757.950 ;
        RECT 335.100 756.150 336.900 757.950 ;
        RECT 350.100 756.150 351.900 757.950 ;
        RECT 353.100 753.600 354.300 757.950 ;
        RECT 356.100 756.150 357.900 757.950 ;
        RECT 313.200 752.400 315.000 753.300 ;
        RECT 329.700 752.700 333.300 753.600 ;
        RECT 350.700 752.700 354.300 753.600 ;
        RECT 313.200 751.500 318.900 752.400 ;
        RECT 275.100 744.000 276.900 747.600 ;
        RECT 278.100 744.600 279.900 747.600 ;
        RECT 281.100 744.000 282.900 747.600 ;
        RECT 293.100 744.000 294.900 747.600 ;
        RECT 296.100 744.600 297.900 747.600 ;
        RECT 311.100 744.600 312.900 750.600 ;
        RECT 314.100 744.000 315.900 750.600 ;
        RECT 317.700 747.600 318.900 751.500 ;
        RECT 329.700 750.600 330.900 752.700 ;
        RECT 317.100 744.600 318.900 747.600 ;
        RECT 329.100 744.600 330.900 750.600 ;
        RECT 332.100 749.700 339.900 751.050 ;
        RECT 350.700 750.600 351.900 752.700 ;
        RECT 332.100 744.600 333.900 749.700 ;
        RECT 335.100 744.000 336.900 748.800 ;
        RECT 338.100 744.600 339.900 749.700 ;
        RECT 350.100 744.600 351.900 750.600 ;
        RECT 353.100 749.700 360.900 751.050 ;
        RECT 353.100 744.600 354.900 749.700 ;
        RECT 356.100 744.000 357.900 748.800 ;
        RECT 359.100 744.600 360.900 749.700 ;
        RECT 374.700 747.600 375.600 757.950 ;
        RECT 389.100 756.150 390.900 757.950 ;
        RECT 392.100 753.600 393.300 757.950 ;
        RECT 395.100 756.150 396.900 757.950 ;
        RECT 389.700 752.700 393.300 753.600 ;
        RECT 389.700 750.600 390.900 752.700 ;
        RECT 371.100 744.000 372.900 747.600 ;
        RECT 374.100 744.600 375.900 747.600 ;
        RECT 377.100 744.000 378.900 747.600 ;
        RECT 389.100 744.600 390.900 750.600 ;
        RECT 392.100 749.700 399.900 751.050 ;
        RECT 392.100 744.600 393.900 749.700 ;
        RECT 395.100 744.000 396.900 748.800 ;
        RECT 398.100 744.600 399.900 749.700 ;
        RECT 413.400 747.600 414.300 757.950 ;
        RECT 428.100 750.600 429.300 757.950 ;
        RECT 431.100 753.300 432.000 764.700 ;
        RECT 433.800 760.050 435.600 761.850 ;
        RECT 446.100 760.050 447.900 761.850 ;
        RECT 452.700 760.050 453.900 767.400 ;
        RECT 470.100 760.050 471.300 773.400 ;
        RECT 476.550 767.400 478.350 779.400 ;
        RECT 479.550 767.400 481.350 780.000 ;
        RECT 484.350 773.400 486.150 779.400 ;
        RECT 488.850 773.400 490.650 780.000 ;
        RECT 484.350 771.300 486.450 773.400 ;
        RECT 491.850 772.500 493.650 779.400 ;
        RECT 494.850 773.400 496.650 780.000 ;
        RECT 490.950 771.450 497.550 772.500 ;
        RECT 490.950 770.700 492.750 771.450 ;
        RECT 495.750 770.700 497.550 771.450 ;
        RECT 499.650 770.400 501.450 779.400 ;
        RECT 483.450 768.600 486.450 770.400 ;
        RECT 487.350 769.800 489.150 770.400 ;
        RECT 487.350 768.900 493.050 769.800 ;
        RECT 499.650 769.500 501.750 770.400 ;
        RECT 487.350 768.600 489.150 768.900 ;
        RECT 485.250 767.700 486.450 768.600 ;
        RECT 476.550 760.050 477.750 767.400 ;
        RECT 485.250 766.800 490.050 767.700 ;
        RECT 478.650 764.100 480.450 764.550 ;
        RECT 484.350 764.100 486.450 764.700 ;
        RECT 478.650 762.900 486.450 764.100 ;
        RECT 478.650 762.750 480.450 762.900 ;
        RECT 484.350 762.600 486.450 762.900 ;
        RECT 433.500 757.950 435.600 760.050 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 454.950 757.950 457.050 760.050 ;
        RECT 466.950 757.950 469.050 760.050 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 476.550 759.750 481.050 760.050 ;
        RECT 476.550 757.950 482.850 759.750 ;
        RECT 449.100 756.150 450.900 757.950 ;
        RECT 430.200 752.400 432.000 753.300 ;
        RECT 452.700 753.600 453.900 757.950 ;
        RECT 455.100 756.150 456.900 757.950 ;
        RECT 467.250 756.150 469.050 757.950 ;
        RECT 452.700 752.700 456.300 753.600 ;
        RECT 430.200 751.500 435.900 752.400 ;
        RECT 410.100 744.000 411.900 747.600 ;
        RECT 413.100 744.600 414.900 747.600 ;
        RECT 416.100 744.000 417.900 747.600 ;
        RECT 428.100 744.600 429.900 750.600 ;
        RECT 431.100 744.000 432.900 750.600 ;
        RECT 434.700 747.600 435.900 751.500 ;
        RECT 434.100 744.600 435.900 747.600 ;
        RECT 446.100 749.700 453.900 751.050 ;
        RECT 446.100 744.600 447.900 749.700 ;
        RECT 449.100 744.000 450.900 748.800 ;
        RECT 452.100 744.600 453.900 749.700 ;
        RECT 455.100 750.600 456.300 752.700 ;
        RECT 470.100 752.700 471.300 757.950 ;
        RECT 473.100 756.150 474.900 757.950 ;
        RECT 470.100 751.800 474.300 752.700 ;
        RECT 455.100 744.600 456.900 750.600 ;
        RECT 467.400 744.000 469.200 750.600 ;
        RECT 472.500 744.600 474.300 751.800 ;
        RECT 476.550 750.600 477.750 757.950 ;
        RECT 489.150 754.200 490.050 766.800 ;
        RECT 492.150 766.800 493.050 768.900 ;
        RECT 493.950 768.300 501.750 769.500 ;
        RECT 493.950 767.700 495.750 768.300 ;
        RECT 505.050 767.400 506.850 780.000 ;
        RECT 508.050 769.200 509.850 779.400 ;
        RECT 513.150 769.200 514.950 779.400 ;
        RECT 508.050 767.400 510.450 769.200 ;
        RECT 492.150 766.500 500.550 766.800 ;
        RECT 509.550 766.500 510.450 767.400 ;
        RECT 492.150 765.900 510.450 766.500 ;
        RECT 498.750 765.300 510.450 765.900 ;
        RECT 498.750 765.000 500.550 765.300 ;
        RECT 496.800 758.400 498.900 760.050 ;
        RECT 496.800 757.200 504.900 758.400 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 503.100 756.600 504.900 757.200 ;
        RECT 500.100 755.400 501.900 756.000 ;
        RECT 506.250 755.400 508.050 757.950 ;
        RECT 500.100 754.200 508.050 755.400 ;
        RECT 489.150 753.000 501.150 754.200 ;
        RECT 489.150 752.400 490.950 753.000 ;
        RECT 500.100 751.200 501.150 753.000 ;
        RECT 476.550 744.600 478.350 750.600 ;
        RECT 479.850 744.000 481.650 750.600 ;
        RECT 484.350 747.600 486.750 749.700 ;
        RECT 496.350 749.550 498.150 750.300 ;
        RECT 493.200 748.500 498.150 749.550 ;
        RECT 499.350 749.400 501.150 751.200 ;
        RECT 509.550 750.600 510.450 765.300 ;
        RECT 493.200 747.600 494.250 748.500 ;
        RECT 502.050 748.200 504.150 749.700 ;
        RECT 500.250 747.600 504.150 748.200 ;
        RECT 484.950 744.600 486.750 747.600 ;
        RECT 489.450 744.000 491.250 747.600 ;
        RECT 492.450 744.600 494.250 747.600 ;
        RECT 495.750 744.000 497.550 747.600 ;
        RECT 500.250 746.700 503.850 747.600 ;
        RECT 500.250 744.600 502.050 746.700 ;
        RECT 505.050 744.000 506.850 750.600 ;
        RECT 508.050 748.800 510.450 750.600 ;
        RECT 512.550 767.400 514.950 769.200 ;
        RECT 516.150 767.400 517.950 780.000 ;
        RECT 521.550 770.400 523.350 779.400 ;
        RECT 526.350 773.400 528.150 780.000 ;
        RECT 529.350 772.500 531.150 779.400 ;
        RECT 532.350 773.400 534.150 780.000 ;
        RECT 536.850 773.400 538.650 779.400 ;
        RECT 525.450 771.450 532.050 772.500 ;
        RECT 525.450 770.700 527.250 771.450 ;
        RECT 530.250 770.700 532.050 771.450 ;
        RECT 536.550 771.300 538.650 773.400 ;
        RECT 521.250 769.500 523.350 770.400 ;
        RECT 533.850 769.800 535.650 770.400 ;
        RECT 521.250 768.300 529.050 769.500 ;
        RECT 527.250 767.700 529.050 768.300 ;
        RECT 529.950 768.900 535.650 769.800 ;
        RECT 512.550 766.500 513.450 767.400 ;
        RECT 529.950 766.800 530.850 768.900 ;
        RECT 533.850 768.600 535.650 768.900 ;
        RECT 536.550 768.600 539.550 770.400 ;
        RECT 536.550 767.700 537.750 768.600 ;
        RECT 522.450 766.500 530.850 766.800 ;
        RECT 512.550 765.900 530.850 766.500 ;
        RECT 532.950 766.800 537.750 767.700 ;
        RECT 541.650 767.400 543.450 780.000 ;
        RECT 544.650 767.400 546.450 779.400 ;
        RECT 557.100 773.400 558.900 779.400 ;
        RECT 560.100 773.400 561.900 780.000 ;
        RECT 575.700 773.400 577.500 780.000 ;
        RECT 512.550 765.300 524.250 765.900 ;
        RECT 512.550 750.600 513.450 765.300 ;
        RECT 522.450 765.000 524.250 765.300 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 524.100 758.400 526.200 760.050 ;
        RECT 514.950 755.400 516.750 757.950 ;
        RECT 518.100 757.200 526.200 758.400 ;
        RECT 518.100 756.600 519.900 757.200 ;
        RECT 521.100 755.400 522.900 756.000 ;
        RECT 514.950 754.200 522.900 755.400 ;
        RECT 532.950 754.200 533.850 766.800 ;
        RECT 536.550 764.100 538.650 764.700 ;
        RECT 542.550 764.100 544.350 764.550 ;
        RECT 536.550 762.900 544.350 764.100 ;
        RECT 536.550 762.600 538.650 762.900 ;
        RECT 542.550 762.750 544.350 762.900 ;
        RECT 545.250 760.050 546.450 767.400 ;
        RECT 557.700 760.050 558.900 773.400 ;
        RECT 576.000 770.100 577.800 771.900 ;
        RECT 578.700 768.900 580.500 779.400 ;
        RECT 578.100 767.400 580.500 768.900 ;
        RECT 583.800 767.400 585.600 780.000 ;
        RECT 596.100 773.400 597.900 780.000 ;
        RECT 599.100 773.400 600.900 779.400 ;
        RECT 602.100 773.400 603.900 780.000 ;
        RECT 560.100 760.050 561.900 761.850 ;
        RECT 578.100 760.050 579.300 767.400 ;
        RECT 584.100 760.050 585.900 761.850 ;
        RECT 599.700 760.050 600.900 773.400 ;
        RECT 605.550 767.400 607.350 779.400 ;
        RECT 608.550 767.400 610.350 780.000 ;
        RECT 613.350 773.400 615.150 779.400 ;
        RECT 617.850 773.400 619.650 780.000 ;
        RECT 613.350 771.300 615.450 773.400 ;
        RECT 620.850 772.500 622.650 779.400 ;
        RECT 623.850 773.400 625.650 780.000 ;
        RECT 619.950 771.450 626.550 772.500 ;
        RECT 619.950 770.700 621.750 771.450 ;
        RECT 624.750 770.700 626.550 771.450 ;
        RECT 628.650 770.400 630.450 779.400 ;
        RECT 612.450 768.600 615.450 770.400 ;
        RECT 616.350 769.800 618.150 770.400 ;
        RECT 616.350 768.900 622.050 769.800 ;
        RECT 628.650 769.500 630.750 770.400 ;
        RECT 616.350 768.600 618.150 768.900 ;
        RECT 614.250 767.700 615.450 768.600 ;
        RECT 605.550 760.050 606.750 767.400 ;
        RECT 614.250 766.800 619.050 767.700 ;
        RECT 607.650 764.100 609.450 764.550 ;
        RECT 613.350 764.100 615.450 764.700 ;
        RECT 607.650 762.900 615.450 764.100 ;
        RECT 607.650 762.750 609.450 762.900 ;
        RECT 613.350 762.600 615.450 762.900 ;
        RECT 541.950 759.750 546.450 760.050 ;
        RECT 540.150 757.950 546.450 759.750 ;
        RECT 556.950 757.950 559.050 760.050 ;
        RECT 559.950 757.950 562.050 760.050 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 577.950 757.950 580.050 760.050 ;
        RECT 580.950 757.950 583.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 605.550 759.750 610.050 760.050 ;
        RECT 605.550 757.950 611.850 759.750 ;
        RECT 521.850 753.000 533.850 754.200 ;
        RECT 521.850 751.200 522.900 753.000 ;
        RECT 532.050 752.400 533.850 753.000 ;
        RECT 512.550 748.800 514.950 750.600 ;
        RECT 508.050 744.600 509.850 748.800 ;
        RECT 513.150 744.600 514.950 748.800 ;
        RECT 516.150 744.000 517.950 750.600 ;
        RECT 518.850 748.200 520.950 749.700 ;
        RECT 521.850 749.400 523.650 751.200 ;
        RECT 545.250 750.600 546.450 757.950 ;
        RECT 524.850 749.550 526.650 750.300 ;
        RECT 524.850 748.500 529.800 749.550 ;
        RECT 518.850 747.600 522.750 748.200 ;
        RECT 528.750 747.600 529.800 748.500 ;
        RECT 536.250 747.600 538.650 749.700 ;
        RECT 519.150 746.700 522.750 747.600 ;
        RECT 520.950 744.600 522.750 746.700 ;
        RECT 525.450 744.000 527.250 747.600 ;
        RECT 528.750 744.600 530.550 747.600 ;
        RECT 531.750 744.000 533.550 747.600 ;
        RECT 536.250 744.600 538.050 747.600 ;
        RECT 541.350 744.000 543.150 750.600 ;
        RECT 544.650 744.600 546.450 750.600 ;
        RECT 557.700 747.600 558.900 757.950 ;
        RECT 575.100 756.150 576.900 757.950 ;
        RECT 578.100 753.600 579.300 757.950 ;
        RECT 581.100 756.150 582.900 757.950 ;
        RECT 596.100 756.150 597.900 757.950 ;
        RECT 575.700 752.700 579.300 753.600 ;
        RECT 599.700 752.700 600.900 757.950 ;
        RECT 601.950 756.150 603.750 757.950 ;
        RECT 575.700 750.600 576.900 752.700 ;
        RECT 596.700 751.800 600.900 752.700 ;
        RECT 557.100 744.600 558.900 747.600 ;
        RECT 560.100 744.000 561.900 747.600 ;
        RECT 575.100 744.600 576.900 750.600 ;
        RECT 578.100 749.700 585.900 751.050 ;
        RECT 578.100 744.600 579.900 749.700 ;
        RECT 581.100 744.000 582.900 748.800 ;
        RECT 584.100 744.600 585.900 749.700 ;
        RECT 596.700 744.600 598.500 751.800 ;
        RECT 605.550 750.600 606.750 757.950 ;
        RECT 618.150 754.200 619.050 766.800 ;
        RECT 621.150 766.800 622.050 768.900 ;
        RECT 622.950 768.300 630.750 769.500 ;
        RECT 622.950 767.700 624.750 768.300 ;
        RECT 634.050 767.400 635.850 780.000 ;
        RECT 637.050 769.200 638.850 779.400 ;
        RECT 650.700 773.400 652.500 780.000 ;
        RECT 651.000 770.100 652.800 771.900 ;
        RECT 637.050 767.400 639.450 769.200 ;
        RECT 653.700 768.900 655.500 779.400 ;
        RECT 621.150 766.500 629.550 766.800 ;
        RECT 638.550 766.500 639.450 767.400 ;
        RECT 621.150 765.900 639.450 766.500 ;
        RECT 627.750 765.300 639.450 765.900 ;
        RECT 627.750 765.000 629.550 765.300 ;
        RECT 625.800 758.400 627.900 760.050 ;
        RECT 625.800 757.200 633.900 758.400 ;
        RECT 634.950 757.950 637.050 760.050 ;
        RECT 632.100 756.600 633.900 757.200 ;
        RECT 629.100 755.400 630.900 756.000 ;
        RECT 635.250 755.400 637.050 757.950 ;
        RECT 629.100 754.200 637.050 755.400 ;
        RECT 618.150 753.000 630.150 754.200 ;
        RECT 618.150 752.400 619.950 753.000 ;
        RECT 629.100 751.200 630.150 753.000 ;
        RECT 601.800 744.000 603.600 750.600 ;
        RECT 605.550 744.600 607.350 750.600 ;
        RECT 608.850 744.000 610.650 750.600 ;
        RECT 613.350 747.600 615.750 749.700 ;
        RECT 625.350 749.550 627.150 750.300 ;
        RECT 622.200 748.500 627.150 749.550 ;
        RECT 628.350 749.400 630.150 751.200 ;
        RECT 638.550 750.600 639.450 765.300 ;
        RECT 653.100 767.400 655.500 768.900 ;
        RECT 658.800 767.400 660.600 780.000 ;
        RECT 672.000 768.600 673.800 779.400 ;
        RECT 672.000 767.400 675.600 768.600 ;
        RECT 677.100 767.400 678.900 780.000 ;
        RECT 689.100 773.400 690.900 780.000 ;
        RECT 692.100 773.400 693.900 779.400 ;
        RECT 707.700 773.400 709.500 780.000 ;
        RECT 653.100 760.050 654.300 767.400 ;
        RECT 659.100 760.050 660.900 761.850 ;
        RECT 671.100 760.050 672.900 761.850 ;
        RECT 674.700 760.050 675.600 767.400 ;
        RECT 676.950 760.050 678.750 761.850 ;
        RECT 689.100 760.050 690.900 761.850 ;
        RECT 692.100 760.050 693.300 773.400 ;
        RECT 708.000 770.100 709.800 771.900 ;
        RECT 710.700 768.900 712.500 779.400 ;
        RECT 710.100 767.400 712.500 768.900 ;
        RECT 715.800 767.400 717.600 780.000 ;
        RECT 728.100 773.400 729.900 779.400 ;
        RECT 731.100 773.400 732.900 780.000 ;
        RECT 743.100 773.400 744.900 779.400 ;
        RECT 746.100 773.400 747.900 780.000 ;
        RECT 710.100 760.050 711.300 767.400 ;
        RECT 712.950 765.450 715.050 766.050 ;
        RECT 724.950 765.450 727.050 766.050 ;
        RECT 712.950 764.550 727.050 765.450 ;
        RECT 712.950 763.950 715.050 764.550 ;
        RECT 724.950 763.950 727.050 764.550 ;
        RECT 716.100 760.050 717.900 761.850 ;
        RECT 728.700 760.050 729.900 773.400 ;
        RECT 731.100 760.050 732.900 761.850 ;
        RECT 743.700 760.050 744.900 773.400 ;
        RECT 758.100 767.400 759.900 779.400 ;
        RECT 761.100 768.300 762.900 779.400 ;
        RECT 764.100 769.200 765.900 780.000 ;
        RECT 767.100 768.300 768.900 779.400 ;
        RECT 761.100 767.400 768.900 768.300 ;
        RECT 780.000 768.600 781.800 779.400 ;
        RECT 780.000 767.400 783.600 768.600 ;
        RECT 785.100 767.400 786.900 780.000 ;
        RECT 797.100 767.400 798.900 780.000 ;
        RECT 802.200 768.600 804.000 779.400 ;
        RECT 800.400 767.400 804.000 768.600 ;
        RECT 815.400 767.400 817.200 780.000 ;
        RECT 820.500 768.900 822.300 779.400 ;
        RECT 823.500 773.400 825.300 780.000 ;
        RECT 823.200 770.100 825.000 771.900 ;
        RECT 828.150 769.200 829.950 779.400 ;
        RECT 820.500 767.400 822.900 768.900 ;
        RECT 746.100 760.050 747.900 761.850 ;
        RECT 758.400 760.050 759.300 767.400 ;
        RECT 763.950 760.050 765.750 761.850 ;
        RECT 779.100 760.050 780.900 761.850 ;
        RECT 782.700 760.050 783.600 767.400 ;
        RECT 784.950 760.050 786.750 761.850 ;
        RECT 797.250 760.050 799.050 761.850 ;
        RECT 800.400 760.050 801.300 767.400 ;
        RECT 803.100 760.050 804.900 761.850 ;
        RECT 815.100 760.050 816.900 761.850 ;
        RECT 821.700 760.050 822.900 767.400 ;
        RECT 827.550 767.400 829.950 769.200 ;
        RECT 831.150 767.400 832.950 780.000 ;
        RECT 836.550 770.400 838.350 779.400 ;
        RECT 841.350 773.400 843.150 780.000 ;
        RECT 844.350 772.500 846.150 779.400 ;
        RECT 847.350 773.400 849.150 780.000 ;
        RECT 851.850 773.400 853.650 779.400 ;
        RECT 840.450 771.450 847.050 772.500 ;
        RECT 840.450 770.700 842.250 771.450 ;
        RECT 845.250 770.700 847.050 771.450 ;
        RECT 851.550 771.300 853.650 773.400 ;
        RECT 836.250 769.500 838.350 770.400 ;
        RECT 848.850 769.800 850.650 770.400 ;
        RECT 836.250 768.300 844.050 769.500 ;
        RECT 842.250 767.700 844.050 768.300 ;
        RECT 844.950 768.900 850.650 769.800 ;
        RECT 827.550 766.500 828.450 767.400 ;
        RECT 844.950 766.800 845.850 768.900 ;
        RECT 848.850 768.600 850.650 768.900 ;
        RECT 851.550 768.600 854.550 770.400 ;
        RECT 851.550 767.700 852.750 768.600 ;
        RECT 837.450 766.500 845.850 766.800 ;
        RECT 827.550 765.900 845.850 766.500 ;
        RECT 847.950 766.800 852.750 767.700 ;
        RECT 856.650 767.400 858.450 780.000 ;
        RECT 859.650 767.400 861.450 779.400 ;
        RECT 827.550 765.300 839.250 765.900 ;
        RECT 649.950 757.950 652.050 760.050 ;
        RECT 652.950 757.950 655.050 760.050 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 688.950 757.950 691.050 760.050 ;
        RECT 691.950 757.950 694.050 760.050 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 715.950 757.950 718.050 760.050 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 742.950 757.950 745.050 760.050 ;
        RECT 745.950 757.950 748.050 760.050 ;
        RECT 757.950 757.950 760.050 760.050 ;
        RECT 760.950 757.950 763.050 760.050 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 784.950 757.950 787.050 760.050 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 650.100 756.150 651.900 757.950 ;
        RECT 653.100 753.600 654.300 757.950 ;
        RECT 656.100 756.150 657.900 757.950 ;
        RECT 650.700 752.700 654.300 753.600 ;
        RECT 650.700 750.600 651.900 752.700 ;
        RECT 622.200 747.600 623.250 748.500 ;
        RECT 631.050 748.200 633.150 749.700 ;
        RECT 629.250 747.600 633.150 748.200 ;
        RECT 613.950 744.600 615.750 747.600 ;
        RECT 618.450 744.000 620.250 747.600 ;
        RECT 621.450 744.600 623.250 747.600 ;
        RECT 624.750 744.000 626.550 747.600 ;
        RECT 629.250 746.700 632.850 747.600 ;
        RECT 629.250 744.600 631.050 746.700 ;
        RECT 634.050 744.000 635.850 750.600 ;
        RECT 637.050 748.800 639.450 750.600 ;
        RECT 637.050 744.600 638.850 748.800 ;
        RECT 650.100 744.600 651.900 750.600 ;
        RECT 653.100 749.700 660.900 751.050 ;
        RECT 653.100 744.600 654.900 749.700 ;
        RECT 656.100 744.000 657.900 748.800 ;
        RECT 659.100 744.600 660.900 749.700 ;
        RECT 674.700 747.600 675.600 757.950 ;
        RECT 692.100 747.600 693.300 757.950 ;
        RECT 707.100 756.150 708.900 757.950 ;
        RECT 710.100 753.600 711.300 757.950 ;
        RECT 713.100 756.150 714.900 757.950 ;
        RECT 707.700 752.700 711.300 753.600 ;
        RECT 707.700 750.600 708.900 752.700 ;
        RECT 671.100 744.000 672.900 747.600 ;
        RECT 674.100 744.600 675.900 747.600 ;
        RECT 677.100 744.000 678.900 747.600 ;
        RECT 689.100 744.000 690.900 747.600 ;
        RECT 692.100 744.600 693.900 747.600 ;
        RECT 707.100 744.600 708.900 750.600 ;
        RECT 710.100 749.700 717.900 751.050 ;
        RECT 710.100 744.600 711.900 749.700 ;
        RECT 713.100 744.000 714.900 748.800 ;
        RECT 716.100 744.600 717.900 749.700 ;
        RECT 728.700 747.600 729.900 757.950 ;
        RECT 743.700 747.600 744.900 757.950 ;
        RECT 758.400 750.600 759.300 757.950 ;
        RECT 760.950 756.150 762.750 757.950 ;
        RECT 767.100 756.150 768.900 757.950 ;
        RECT 758.400 749.400 763.500 750.600 ;
        RECT 728.100 744.600 729.900 747.600 ;
        RECT 731.100 744.000 732.900 747.600 ;
        RECT 743.100 744.600 744.900 747.600 ;
        RECT 746.100 744.000 747.900 747.600 ;
        RECT 758.700 744.000 760.500 747.600 ;
        RECT 761.700 744.600 763.500 749.400 ;
        RECT 766.200 744.000 768.000 750.600 ;
        RECT 782.700 747.600 783.600 757.950 ;
        RECT 800.400 747.600 801.300 757.950 ;
        RECT 818.100 756.150 819.900 757.950 ;
        RECT 821.700 753.600 822.900 757.950 ;
        RECT 824.100 756.150 825.900 757.950 ;
        RECT 821.700 752.700 825.300 753.600 ;
        RECT 815.100 749.700 822.900 751.050 ;
        RECT 779.100 744.000 780.900 747.600 ;
        RECT 782.100 744.600 783.900 747.600 ;
        RECT 785.100 744.000 786.900 747.600 ;
        RECT 797.100 744.000 798.900 747.600 ;
        RECT 800.100 744.600 801.900 747.600 ;
        RECT 803.100 744.000 804.900 747.600 ;
        RECT 815.100 744.600 816.900 749.700 ;
        RECT 818.100 744.000 819.900 748.800 ;
        RECT 821.100 744.600 822.900 749.700 ;
        RECT 824.100 750.600 825.300 752.700 ;
        RECT 827.550 750.600 828.450 765.300 ;
        RECT 837.450 765.000 839.250 765.300 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 839.100 758.400 841.200 760.050 ;
        RECT 829.950 755.400 831.750 757.950 ;
        RECT 833.100 757.200 841.200 758.400 ;
        RECT 833.100 756.600 834.900 757.200 ;
        RECT 836.100 755.400 837.900 756.000 ;
        RECT 829.950 754.200 837.900 755.400 ;
        RECT 847.950 754.200 848.850 766.800 ;
        RECT 851.550 764.100 853.650 764.700 ;
        RECT 857.550 764.100 859.350 764.550 ;
        RECT 851.550 762.900 859.350 764.100 ;
        RECT 851.550 762.600 853.650 762.900 ;
        RECT 857.550 762.750 859.350 762.900 ;
        RECT 860.250 760.050 861.450 767.400 ;
        RECT 856.950 759.750 861.450 760.050 ;
        RECT 855.150 757.950 861.450 759.750 ;
        RECT 836.850 753.000 848.850 754.200 ;
        RECT 836.850 751.200 837.900 753.000 ;
        RECT 847.050 752.400 848.850 753.000 ;
        RECT 824.100 744.600 825.900 750.600 ;
        RECT 827.550 748.800 829.950 750.600 ;
        RECT 828.150 744.600 829.950 748.800 ;
        RECT 831.150 744.000 832.950 750.600 ;
        RECT 833.850 748.200 835.950 749.700 ;
        RECT 836.850 749.400 838.650 751.200 ;
        RECT 860.250 750.600 861.450 757.950 ;
        RECT 839.850 749.550 841.650 750.300 ;
        RECT 839.850 748.500 844.800 749.550 ;
        RECT 833.850 747.600 837.750 748.200 ;
        RECT 843.750 747.600 844.800 748.500 ;
        RECT 851.250 747.600 853.650 749.700 ;
        RECT 834.150 746.700 837.750 747.600 ;
        RECT 835.950 744.600 837.750 746.700 ;
        RECT 840.450 744.000 842.250 747.600 ;
        RECT 843.750 744.600 845.550 747.600 ;
        RECT 846.750 744.000 848.550 747.600 ;
        RECT 851.250 744.600 853.050 747.600 ;
        RECT 856.350 744.000 858.150 750.600 ;
        RECT 859.650 744.600 861.450 750.600 ;
        RECT 11.400 734.400 13.200 741.000 ;
        RECT 16.500 733.200 18.300 740.400 ;
        RECT 29.100 737.400 30.900 741.000 ;
        RECT 32.100 737.400 33.900 740.400 ;
        RECT 35.100 737.400 36.900 741.000 ;
        RECT 14.100 732.300 18.300 733.200 ;
        RECT 11.250 727.050 13.050 728.850 ;
        RECT 14.100 727.050 15.300 732.300 ;
        RECT 17.100 727.050 18.900 728.850 ;
        RECT 32.700 727.050 33.600 737.400 ;
        RECT 47.100 735.300 48.900 740.400 ;
        RECT 50.100 736.200 51.900 741.000 ;
        RECT 53.100 735.300 54.900 740.400 ;
        RECT 47.100 733.950 54.900 735.300 ;
        RECT 56.100 734.400 57.900 740.400 ;
        RECT 68.400 734.400 70.200 741.000 ;
        RECT 56.100 732.300 57.300 734.400 ;
        RECT 73.500 733.200 75.300 740.400 ;
        RECT 86.100 737.400 87.900 741.000 ;
        RECT 89.100 737.400 90.900 740.400 ;
        RECT 92.100 737.400 93.900 741.000 ;
        RECT 53.700 731.400 57.300 732.300 ;
        RECT 71.100 732.300 75.300 733.200 ;
        RECT 50.100 727.050 51.900 728.850 ;
        RECT 53.700 727.050 54.900 731.400 ;
        RECT 56.100 727.050 57.900 728.850 ;
        RECT 68.250 727.050 70.050 728.850 ;
        RECT 71.100 727.050 72.300 732.300 ;
        RECT 74.100 727.050 75.900 728.850 ;
        RECT 89.400 727.050 90.300 737.400 ;
        RECT 104.100 734.400 105.900 740.400 ;
        RECT 104.700 732.300 105.900 734.400 ;
        RECT 107.100 735.300 108.900 740.400 ;
        RECT 110.100 736.200 111.900 741.000 ;
        RECT 113.100 735.300 114.900 740.400 ;
        RECT 125.100 737.400 126.900 740.400 ;
        RECT 128.100 737.400 129.900 741.000 ;
        RECT 107.100 733.950 114.900 735.300 ;
        RECT 104.700 731.400 108.300 732.300 ;
        RECT 104.100 727.050 105.900 728.850 ;
        RECT 107.100 727.050 108.300 731.400 ;
        RECT 110.100 727.050 111.900 728.850 ;
        RECT 125.700 727.050 126.900 737.400 ;
        RECT 131.550 734.400 133.350 740.400 ;
        RECT 134.850 734.400 136.650 741.000 ;
        RECT 139.950 737.400 141.750 740.400 ;
        RECT 144.450 737.400 146.250 741.000 ;
        RECT 147.450 737.400 149.250 740.400 ;
        RECT 150.750 737.400 152.550 741.000 ;
        RECT 155.250 738.300 157.050 740.400 ;
        RECT 155.250 737.400 158.850 738.300 ;
        RECT 139.350 735.300 141.750 737.400 ;
        RECT 148.200 736.500 149.250 737.400 ;
        RECT 155.250 736.800 159.150 737.400 ;
        RECT 148.200 735.450 153.150 736.500 ;
        RECT 151.350 734.700 153.150 735.450 ;
        RECT 131.550 727.050 132.750 734.400 ;
        RECT 154.350 733.800 156.150 735.600 ;
        RECT 157.050 735.300 159.150 736.800 ;
        RECT 160.050 734.400 161.850 741.000 ;
        RECT 163.050 736.200 164.850 740.400 ;
        RECT 176.100 737.400 177.900 741.000 ;
        RECT 179.100 737.400 180.900 740.400 ;
        RECT 182.100 737.400 183.900 741.000 ;
        RECT 194.700 737.400 196.500 741.000 ;
        RECT 163.050 734.400 165.450 736.200 ;
        RECT 144.150 732.000 145.950 732.600 ;
        RECT 155.100 732.000 156.150 733.800 ;
        RECT 144.150 730.800 156.150 732.000 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 28.950 724.950 31.050 727.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 46.950 724.950 49.050 727.050 ;
        RECT 49.950 724.950 52.050 727.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 67.950 724.950 70.050 727.050 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 91.950 724.950 94.050 727.050 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 131.550 725.250 137.850 727.050 ;
        RECT 131.550 724.950 136.050 725.250 ;
        RECT 14.100 711.600 15.300 724.950 ;
        RECT 29.100 723.150 30.900 724.950 ;
        RECT 16.950 720.450 19.050 721.050 ;
        RECT 28.950 720.450 31.050 721.050 ;
        RECT 16.950 719.550 31.050 720.450 ;
        RECT 16.950 718.950 19.050 719.550 ;
        RECT 28.950 718.950 31.050 719.550 ;
        RECT 32.700 717.600 33.600 724.950 ;
        RECT 34.950 723.150 36.750 724.950 ;
        RECT 47.100 723.150 48.900 724.950 ;
        RECT 53.700 717.600 54.900 724.950 ;
        RECT 30.000 716.400 33.600 717.600 ;
        RECT 11.100 705.000 12.900 711.600 ;
        RECT 14.100 705.600 15.900 711.600 ;
        RECT 17.100 705.000 18.900 711.600 ;
        RECT 30.000 705.600 31.800 716.400 ;
        RECT 35.100 705.000 36.900 717.600 ;
        RECT 47.400 705.000 49.200 717.600 ;
        RECT 52.500 716.100 54.900 717.600 ;
        RECT 52.500 705.600 54.300 716.100 ;
        RECT 55.200 713.100 57.000 714.900 ;
        RECT 71.100 711.600 72.300 724.950 ;
        RECT 86.250 723.150 88.050 724.950 ;
        RECT 89.400 717.600 90.300 724.950 ;
        RECT 92.100 723.150 93.900 724.950 ;
        RECT 107.100 717.600 108.300 724.950 ;
        RECT 113.100 723.150 114.900 724.950 ;
        RECT 55.500 705.000 57.300 711.600 ;
        RECT 68.100 705.000 69.900 711.600 ;
        RECT 71.100 705.600 72.900 711.600 ;
        RECT 74.100 705.000 75.900 711.600 ;
        RECT 86.100 705.000 87.900 717.600 ;
        RECT 89.400 716.400 93.000 717.600 ;
        RECT 91.200 705.600 93.000 716.400 ;
        RECT 107.100 716.100 109.500 717.600 ;
        RECT 105.000 713.100 106.800 714.900 ;
        RECT 104.700 705.000 106.500 711.600 ;
        RECT 107.700 705.600 109.500 716.100 ;
        RECT 112.800 705.000 114.600 717.600 ;
        RECT 125.700 711.600 126.900 724.950 ;
        RECT 128.100 723.150 129.900 724.950 ;
        RECT 131.550 717.600 132.750 724.950 ;
        RECT 133.650 722.100 135.450 722.250 ;
        RECT 139.350 722.100 141.450 722.400 ;
        RECT 133.650 720.900 141.450 722.100 ;
        RECT 133.650 720.450 135.450 720.900 ;
        RECT 139.350 720.300 141.450 720.900 ;
        RECT 144.150 718.200 145.050 730.800 ;
        RECT 155.100 729.600 163.050 730.800 ;
        RECT 155.100 729.000 156.900 729.600 ;
        RECT 158.100 727.800 159.900 728.400 ;
        RECT 151.800 726.600 159.900 727.800 ;
        RECT 161.250 727.050 163.050 729.600 ;
        RECT 151.800 724.950 153.900 726.600 ;
        RECT 160.950 724.950 163.050 727.050 ;
        RECT 153.750 719.700 155.550 720.000 ;
        RECT 164.550 719.700 165.450 734.400 ;
        RECT 166.950 732.450 169.050 736.050 ;
        RECT 175.950 732.450 178.050 733.050 ;
        RECT 166.950 732.000 178.050 732.450 ;
        RECT 167.550 731.550 178.050 732.000 ;
        RECT 175.950 730.950 178.050 731.550 ;
        RECT 166.950 729.450 169.050 729.900 ;
        RECT 172.950 729.450 175.050 730.050 ;
        RECT 166.950 728.550 175.050 729.450 ;
        RECT 166.950 727.800 169.050 728.550 ;
        RECT 172.950 727.950 175.050 728.550 ;
        RECT 179.700 727.050 180.600 737.400 ;
        RECT 197.700 735.600 199.500 740.400 ;
        RECT 194.400 734.400 199.500 735.600 ;
        RECT 202.200 734.400 204.000 741.000 ;
        RECT 215.100 737.400 216.900 741.000 ;
        RECT 218.100 737.400 219.900 740.400 ;
        RECT 194.400 727.050 195.300 734.400 ;
        RECT 210.000 729.450 214.050 730.050 ;
        RECT 196.950 727.050 198.750 728.850 ;
        RECT 203.100 727.050 204.900 728.850 ;
        RECT 209.550 727.950 214.050 729.450 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 181.950 724.950 184.050 727.050 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 202.950 724.950 205.050 727.050 ;
        RECT 176.100 723.150 177.900 724.950 ;
        RECT 153.750 719.100 165.450 719.700 ;
        RECT 125.100 705.600 126.900 711.600 ;
        RECT 128.100 705.000 129.900 711.600 ;
        RECT 131.550 705.600 133.350 717.600 ;
        RECT 134.550 705.000 136.350 717.600 ;
        RECT 140.250 717.300 145.050 718.200 ;
        RECT 147.150 718.500 165.450 719.100 ;
        RECT 147.150 718.200 155.550 718.500 ;
        RECT 140.250 716.400 141.450 717.300 ;
        RECT 138.450 714.600 141.450 716.400 ;
        RECT 142.350 716.100 144.150 716.400 ;
        RECT 147.150 716.100 148.050 718.200 ;
        RECT 164.550 717.600 165.450 718.500 ;
        RECT 179.700 717.600 180.600 724.950 ;
        RECT 181.950 723.150 183.750 724.950 ;
        RECT 194.400 717.600 195.300 724.950 ;
        RECT 199.950 723.150 201.750 724.950 ;
        RECT 199.950 720.450 202.050 721.050 ;
        RECT 209.550 720.450 210.450 727.950 ;
        RECT 218.100 727.050 219.300 737.400 ;
        RECT 230.100 734.400 231.900 740.400 ;
        RECT 230.700 732.300 231.900 734.400 ;
        RECT 233.100 735.300 234.900 740.400 ;
        RECT 236.100 736.200 237.900 741.000 ;
        RECT 239.100 735.300 240.900 740.400 ;
        RECT 233.100 733.950 240.900 735.300 ;
        RECT 251.100 735.300 252.900 740.400 ;
        RECT 254.100 736.200 255.900 741.000 ;
        RECT 257.100 735.300 258.900 740.400 ;
        RECT 251.100 733.950 258.900 735.300 ;
        RECT 260.100 734.400 261.900 740.400 ;
        RECT 275.100 737.400 276.900 741.000 ;
        RECT 278.100 737.400 279.900 740.400 ;
        RECT 281.100 737.400 282.900 741.000 ;
        RECT 260.100 732.300 261.300 734.400 ;
        RECT 230.700 731.400 234.300 732.300 ;
        RECT 230.100 727.050 231.900 728.850 ;
        RECT 233.100 727.050 234.300 731.400 ;
        RECT 257.700 731.400 261.300 732.300 ;
        RECT 236.100 727.050 237.900 728.850 ;
        RECT 254.100 727.050 255.900 728.850 ;
        RECT 257.700 727.050 258.900 731.400 ;
        RECT 260.100 727.050 261.900 728.850 ;
        RECT 278.700 727.050 279.600 737.400 ;
        RECT 293.100 734.400 294.900 740.400 ;
        RECT 296.100 735.300 297.900 741.000 ;
        RECT 300.600 734.400 302.400 740.400 ;
        RECT 305.100 735.300 306.900 741.000 ;
        RECT 308.100 734.400 309.900 740.400 ;
        RECT 320.100 734.400 321.900 740.400 ;
        RECT 293.700 732.600 294.900 734.400 ;
        RECT 300.900 732.900 302.100 734.400 ;
        RECT 305.100 733.500 309.900 734.400 ;
        RECT 293.700 731.700 300.000 732.600 ;
        RECT 297.900 729.600 300.000 731.700 ;
        RECT 293.400 727.050 295.200 728.850 ;
        RECT 298.200 727.800 300.000 729.600 ;
        RECT 300.900 730.800 303.900 732.900 ;
        RECT 305.100 732.300 307.200 733.500 ;
        RECT 320.700 732.300 321.900 734.400 ;
        RECT 323.100 735.300 324.900 740.400 ;
        RECT 326.100 736.200 327.900 741.000 ;
        RECT 329.100 735.300 330.900 740.400 ;
        RECT 341.100 737.400 342.900 740.400 ;
        RECT 344.100 737.400 345.900 741.000 ;
        RECT 323.100 733.950 330.900 735.300 ;
        RECT 320.700 731.400 324.300 732.300 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 229.950 724.950 232.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 280.950 724.950 283.050 727.050 ;
        RECT 293.100 726.300 295.200 727.050 ;
        RECT 293.100 724.950 300.000 726.300 ;
        RECT 215.100 723.150 216.900 724.950 ;
        RECT 199.950 719.550 210.450 720.450 ;
        RECT 199.950 718.950 202.050 719.550 ;
        RECT 142.350 715.200 148.050 716.100 ;
        RECT 148.950 716.700 150.750 717.300 ;
        RECT 148.950 715.500 156.750 716.700 ;
        RECT 142.350 714.600 144.150 715.200 ;
        RECT 154.650 714.600 156.750 715.500 ;
        RECT 139.350 711.600 141.450 713.700 ;
        RECT 145.950 713.550 147.750 714.300 ;
        RECT 150.750 713.550 152.550 714.300 ;
        RECT 145.950 712.500 152.550 713.550 ;
        RECT 139.350 705.600 141.150 711.600 ;
        RECT 143.850 705.000 145.650 711.600 ;
        RECT 146.850 705.600 148.650 712.500 ;
        RECT 149.850 705.000 151.650 711.600 ;
        RECT 154.650 705.600 156.450 714.600 ;
        RECT 160.050 705.000 161.850 717.600 ;
        RECT 163.050 715.800 165.450 717.600 ;
        RECT 177.000 716.400 180.600 717.600 ;
        RECT 163.050 705.600 164.850 715.800 ;
        RECT 177.000 705.600 178.800 716.400 ;
        RECT 182.100 705.000 183.900 717.600 ;
        RECT 194.100 705.600 195.900 717.600 ;
        RECT 197.100 716.700 204.900 717.600 ;
        RECT 197.100 705.600 198.900 716.700 ;
        RECT 200.100 705.000 201.900 715.800 ;
        RECT 203.100 705.600 204.900 716.700 ;
        RECT 218.100 711.600 219.300 724.950 ;
        RECT 233.100 717.600 234.300 724.950 ;
        RECT 239.100 723.150 240.900 724.950 ;
        RECT 251.100 723.150 252.900 724.950 ;
        RECT 257.700 717.600 258.900 724.950 ;
        RECT 275.100 723.150 276.900 724.950 ;
        RECT 278.700 717.600 279.600 724.950 ;
        RECT 280.950 723.150 282.750 724.950 ;
        RECT 298.200 724.500 300.000 724.950 ;
        RECT 300.900 725.100 302.100 730.800 ;
        RECT 303.000 727.800 305.100 729.900 ;
        RECT 303.300 726.000 305.100 727.800 ;
        RECT 320.100 727.050 321.900 728.850 ;
        RECT 323.100 727.050 324.300 731.400 ;
        RECT 326.100 727.050 327.900 728.850 ;
        RECT 341.700 727.050 342.900 737.400 ;
        RECT 356.100 735.300 357.900 740.400 ;
        RECT 359.100 736.200 360.900 741.000 ;
        RECT 362.100 735.300 363.900 740.400 ;
        RECT 356.100 733.950 363.900 735.300 ;
        RECT 365.100 734.400 366.900 740.400 ;
        RECT 377.400 734.400 379.200 741.000 ;
        RECT 365.100 732.300 366.300 734.400 ;
        RECT 382.500 733.200 384.300 740.400 ;
        RECT 395.100 734.400 396.900 740.400 ;
        RECT 398.100 734.400 399.900 741.000 ;
        RECT 410.100 737.400 411.900 740.400 ;
        RECT 413.100 737.400 414.900 741.000 ;
        RECT 362.700 731.400 366.300 732.300 ;
        RECT 380.100 732.300 384.300 733.200 ;
        RECT 359.100 727.050 360.900 728.850 ;
        RECT 362.700 727.050 363.900 731.400 ;
        RECT 365.100 727.050 366.900 728.850 ;
        RECT 377.250 727.050 379.050 728.850 ;
        RECT 380.100 727.050 381.300 732.300 ;
        RECT 383.100 727.050 384.900 728.850 ;
        RECT 395.700 727.050 396.900 734.400 ;
        RECT 398.100 727.050 399.900 728.850 ;
        RECT 410.700 727.050 411.900 737.400 ;
        RECT 425.100 735.000 426.900 740.400 ;
        RECT 428.100 735.900 429.900 741.000 ;
        RECT 431.100 739.500 438.900 740.400 ;
        RECT 431.100 735.000 432.900 739.500 ;
        RECT 425.100 734.100 432.900 735.000 ;
        RECT 434.100 734.400 435.900 738.600 ;
        RECT 437.100 734.400 438.900 739.500 ;
        RECT 449.100 734.400 450.900 740.400 ;
        RECT 434.400 732.900 435.300 734.400 ;
        RECT 430.950 731.700 435.300 732.900 ;
        RECT 436.950 732.450 439.050 733.200 ;
        RECT 428.250 727.050 430.050 728.850 ;
        RECT 300.900 724.200 303.300 725.100 ;
        RECT 301.800 724.050 303.300 724.200 ;
        RECT 307.800 724.950 309.900 727.050 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 382.950 724.950 385.050 727.050 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 409.950 724.950 412.050 727.050 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 427.950 724.950 430.050 727.050 ;
        RECT 430.950 727.050 432.000 731.700 ;
        RECT 436.950 731.550 444.450 732.450 ;
        RECT 436.950 731.100 439.050 731.550 ;
        RECT 433.950 727.050 435.750 728.850 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 436.950 724.950 439.050 727.050 ;
        RECT 297.000 721.500 300.900 723.300 ;
        RECT 298.800 721.200 300.900 721.500 ;
        RECT 301.800 721.950 303.900 724.050 ;
        RECT 307.800 723.150 309.600 724.950 ;
        RECT 301.800 720.000 302.700 721.950 ;
        RECT 295.500 717.600 297.600 719.700 ;
        RECT 301.200 718.950 302.700 720.000 ;
        RECT 301.200 717.600 302.400 718.950 ;
        RECT 233.100 716.100 235.500 717.600 ;
        RECT 231.000 713.100 232.800 714.900 ;
        RECT 215.100 705.000 216.900 711.600 ;
        RECT 218.100 705.600 219.900 711.600 ;
        RECT 230.700 705.000 232.500 711.600 ;
        RECT 233.700 705.600 235.500 716.100 ;
        RECT 238.800 705.000 240.600 717.600 ;
        RECT 251.400 705.000 253.200 717.600 ;
        RECT 256.500 716.100 258.900 717.600 ;
        RECT 276.000 716.400 279.600 717.600 ;
        RECT 256.500 705.600 258.300 716.100 ;
        RECT 259.200 713.100 261.000 714.900 ;
        RECT 259.500 705.000 261.300 711.600 ;
        RECT 276.000 705.600 277.800 716.400 ;
        RECT 281.100 705.000 282.900 717.600 ;
        RECT 293.100 716.700 297.600 717.600 ;
        RECT 293.100 705.600 294.900 716.700 ;
        RECT 296.100 705.000 297.900 715.500 ;
        RECT 300.600 705.600 302.400 717.600 ;
        RECT 305.100 717.600 307.200 718.500 ;
        RECT 323.100 717.600 324.300 724.950 ;
        RECT 329.100 723.150 330.900 724.950 ;
        RECT 305.100 716.400 309.900 717.600 ;
        RECT 305.100 705.000 306.900 715.500 ;
        RECT 308.100 705.600 309.900 716.400 ;
        RECT 323.100 716.100 325.500 717.600 ;
        RECT 321.000 713.100 322.800 714.900 ;
        RECT 320.700 705.000 322.500 711.600 ;
        RECT 323.700 705.600 325.500 716.100 ;
        RECT 328.800 705.000 330.600 717.600 ;
        RECT 341.700 711.600 342.900 724.950 ;
        RECT 344.100 723.150 345.900 724.950 ;
        RECT 356.100 723.150 357.900 724.950 ;
        RECT 362.700 717.600 363.900 724.950 ;
        RECT 341.100 705.600 342.900 711.600 ;
        RECT 344.100 705.000 345.900 711.600 ;
        RECT 356.400 705.000 358.200 717.600 ;
        RECT 361.500 716.100 363.900 717.600 ;
        RECT 361.500 705.600 363.300 716.100 ;
        RECT 364.200 713.100 366.000 714.900 ;
        RECT 380.100 711.600 381.300 724.950 ;
        RECT 395.700 717.600 396.900 724.950 ;
        RECT 364.500 705.000 366.300 711.600 ;
        RECT 377.100 705.000 378.900 711.600 ;
        RECT 380.100 705.600 381.900 711.600 ;
        RECT 383.100 705.000 384.900 711.600 ;
        RECT 395.100 705.600 396.900 717.600 ;
        RECT 398.100 705.000 399.900 717.600 ;
        RECT 410.700 711.600 411.900 724.950 ;
        RECT 413.100 723.150 414.900 724.950 ;
        RECT 425.100 723.150 426.900 724.950 ;
        RECT 430.950 717.600 432.000 724.950 ;
        RECT 436.950 723.150 438.750 724.950 ;
        RECT 443.550 724.050 444.450 731.550 ;
        RECT 449.700 732.300 450.900 734.400 ;
        RECT 452.100 735.300 453.900 740.400 ;
        RECT 455.100 736.200 456.900 741.000 ;
        RECT 458.100 735.300 459.900 740.400 ;
        RECT 470.100 737.400 471.900 741.000 ;
        RECT 473.100 737.400 474.900 740.400 ;
        RECT 488.100 737.400 489.900 741.000 ;
        RECT 491.100 737.400 492.900 740.400 ;
        RECT 494.100 737.400 495.900 741.000 ;
        RECT 452.100 733.950 459.900 735.300 ;
        RECT 463.950 735.450 466.050 736.050 ;
        RECT 469.950 735.450 472.050 736.050 ;
        RECT 463.950 734.550 472.050 735.450 ;
        RECT 463.950 733.950 466.050 734.550 ;
        RECT 469.950 733.950 472.050 734.550 ;
        RECT 449.700 731.400 453.300 732.300 ;
        RECT 449.100 727.050 450.900 728.850 ;
        RECT 452.100 727.050 453.300 731.400 ;
        RECT 465.000 729.450 469.050 730.050 ;
        RECT 455.100 727.050 456.900 728.850 ;
        RECT 464.550 727.950 469.050 729.450 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 451.950 724.950 454.050 727.050 ;
        RECT 454.950 724.950 457.050 727.050 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 439.950 722.550 444.450 724.050 ;
        RECT 439.950 721.950 444.000 722.550 ;
        RECT 452.100 717.600 453.300 724.950 ;
        RECT 458.100 723.150 459.900 724.950 ;
        RECT 464.550 724.050 465.450 727.950 ;
        RECT 473.100 727.050 474.300 737.400 ;
        RECT 491.700 727.050 492.600 737.400 ;
        RECT 506.100 731.400 507.900 741.000 ;
        RECT 512.700 732.000 514.500 740.400 ;
        RECT 527.700 733.200 529.500 740.400 ;
        RECT 532.800 734.400 534.600 741.000 ;
        RECT 545.100 734.400 546.900 740.400 ;
        RECT 527.700 732.300 531.900 733.200 ;
        RECT 512.700 730.800 516.000 732.000 ;
        RECT 506.100 727.050 507.900 728.850 ;
        RECT 512.100 727.050 513.900 728.850 ;
        RECT 515.100 727.050 516.000 730.800 ;
        RECT 527.100 727.050 528.900 728.850 ;
        RECT 530.700 727.050 531.900 732.300 ;
        RECT 545.700 732.300 546.900 734.400 ;
        RECT 548.100 735.300 549.900 740.400 ;
        RECT 551.100 736.200 552.900 741.000 ;
        RECT 554.100 735.300 555.900 740.400 ;
        RECT 566.100 737.400 567.900 740.400 ;
        RECT 569.100 737.400 570.900 741.000 ;
        RECT 548.100 733.950 555.900 735.300 ;
        RECT 545.700 731.400 549.300 732.300 ;
        RECT 540.000 729.450 544.050 730.050 ;
        RECT 532.950 727.050 534.750 728.850 ;
        RECT 539.550 727.950 544.050 729.450 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 487.950 724.950 490.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 464.550 722.550 469.050 724.050 ;
        RECT 470.100 723.150 471.900 724.950 ;
        RECT 465.000 721.950 469.050 722.550 ;
        RECT 410.100 705.600 411.900 711.600 ;
        RECT 413.100 705.000 414.900 711.600 ;
        RECT 425.100 705.000 426.900 717.600 ;
        RECT 429.600 705.600 432.900 717.600 ;
        RECT 435.600 705.000 437.400 717.600 ;
        RECT 452.100 716.100 454.500 717.600 ;
        RECT 450.000 713.100 451.800 714.900 ;
        RECT 449.700 705.000 451.500 711.600 ;
        RECT 452.700 705.600 454.500 716.100 ;
        RECT 457.800 705.000 459.600 717.600 ;
        RECT 473.100 711.600 474.300 724.950 ;
        RECT 488.100 723.150 489.900 724.950 ;
        RECT 491.700 717.600 492.600 724.950 ;
        RECT 493.950 723.150 495.750 724.950 ;
        RECT 509.100 723.150 510.900 724.950 ;
        RECT 489.000 716.400 492.600 717.600 ;
        RECT 470.100 705.000 471.900 711.600 ;
        RECT 473.100 705.600 474.900 711.600 ;
        RECT 489.000 705.600 490.800 716.400 ;
        RECT 494.100 705.000 495.900 717.600 ;
        RECT 515.100 712.800 516.000 724.950 ;
        RECT 509.400 711.900 516.000 712.800 ;
        RECT 509.400 711.600 510.900 711.900 ;
        RECT 506.100 705.000 507.900 711.600 ;
        RECT 509.100 705.600 510.900 711.600 ;
        RECT 515.100 711.600 516.000 711.900 ;
        RECT 530.700 711.600 531.900 724.950 ;
        RECT 539.550 724.050 540.450 727.950 ;
        RECT 545.100 727.050 546.900 728.850 ;
        RECT 548.100 727.050 549.300 731.400 ;
        RECT 551.100 727.050 552.900 728.850 ;
        RECT 566.700 727.050 567.900 737.400 ;
        RECT 572.550 734.400 574.350 740.400 ;
        RECT 575.850 734.400 577.650 741.000 ;
        RECT 580.950 737.400 582.750 740.400 ;
        RECT 585.450 737.400 587.250 741.000 ;
        RECT 588.450 737.400 590.250 740.400 ;
        RECT 591.750 737.400 593.550 741.000 ;
        RECT 596.250 738.300 598.050 740.400 ;
        RECT 596.250 737.400 599.850 738.300 ;
        RECT 580.350 735.300 582.750 737.400 ;
        RECT 589.200 736.500 590.250 737.400 ;
        RECT 596.250 736.800 600.150 737.400 ;
        RECT 589.200 735.450 594.150 736.500 ;
        RECT 592.350 734.700 594.150 735.450 ;
        RECT 572.550 727.050 573.750 734.400 ;
        RECT 595.350 733.800 597.150 735.600 ;
        RECT 598.050 735.300 600.150 736.800 ;
        RECT 601.050 734.400 602.850 741.000 ;
        RECT 604.050 736.200 605.850 740.400 ;
        RECT 604.050 734.400 606.450 736.200 ;
        RECT 617.100 734.400 618.900 741.000 ;
        RECT 585.150 732.000 586.950 732.600 ;
        RECT 596.100 732.000 597.150 733.800 ;
        RECT 585.150 730.800 597.150 732.000 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 572.550 725.250 578.850 727.050 ;
        RECT 572.550 724.950 577.050 725.250 ;
        RECT 535.950 722.550 540.450 724.050 ;
        RECT 535.950 721.950 540.000 722.550 ;
        RECT 548.100 717.600 549.300 724.950 ;
        RECT 554.100 723.150 555.900 724.950 ;
        RECT 548.100 716.100 550.500 717.600 ;
        RECT 546.000 713.100 547.800 714.900 ;
        RECT 512.100 705.000 513.900 711.000 ;
        RECT 515.100 705.600 516.900 711.600 ;
        RECT 527.100 705.000 528.900 711.600 ;
        RECT 530.100 705.600 531.900 711.600 ;
        RECT 533.100 705.000 534.900 711.600 ;
        RECT 545.700 705.000 547.500 711.600 ;
        RECT 548.700 705.600 550.500 716.100 ;
        RECT 553.800 705.000 555.600 717.600 ;
        RECT 566.700 711.600 567.900 724.950 ;
        RECT 569.100 723.150 570.900 724.950 ;
        RECT 572.550 717.600 573.750 724.950 ;
        RECT 574.650 722.100 576.450 722.250 ;
        RECT 580.350 722.100 582.450 722.400 ;
        RECT 574.650 720.900 582.450 722.100 ;
        RECT 574.650 720.450 576.450 720.900 ;
        RECT 580.350 720.300 582.450 720.900 ;
        RECT 585.150 718.200 586.050 730.800 ;
        RECT 596.100 729.600 604.050 730.800 ;
        RECT 596.100 729.000 597.900 729.600 ;
        RECT 599.100 727.800 600.900 728.400 ;
        RECT 592.800 726.600 600.900 727.800 ;
        RECT 602.250 727.050 604.050 729.600 ;
        RECT 592.800 724.950 594.900 726.600 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 594.750 719.700 596.550 720.000 ;
        RECT 605.550 719.700 606.450 734.400 ;
        RECT 620.100 733.500 621.900 740.400 ;
        RECT 623.100 734.400 624.900 741.000 ;
        RECT 626.100 733.500 627.900 740.400 ;
        RECT 629.100 734.400 630.900 741.000 ;
        RECT 632.100 733.500 633.900 740.400 ;
        RECT 635.100 734.400 636.900 741.000 ;
        RECT 638.100 733.500 639.900 740.400 ;
        RECT 641.100 734.400 642.900 741.000 ;
        RECT 653.700 737.400 655.500 741.000 ;
        RECT 656.700 735.600 658.500 740.400 ;
        RECT 653.400 734.400 658.500 735.600 ;
        RECT 661.200 734.400 663.000 741.000 ;
        RECT 674.100 737.400 675.900 740.400 ;
        RECT 677.100 737.400 678.900 741.000 ;
        RECT 620.100 732.300 624.000 733.500 ;
        RECT 626.100 732.300 630.000 733.500 ;
        RECT 632.100 732.300 636.000 733.500 ;
        RECT 638.100 732.300 640.950 733.500 ;
        RECT 622.800 731.400 624.000 732.300 ;
        RECT 628.800 731.400 630.000 732.300 ;
        RECT 634.800 731.400 636.000 732.300 ;
        RECT 622.800 730.200 627.000 731.400 ;
        RECT 619.800 727.050 621.600 728.850 ;
        RECT 619.800 724.950 621.900 727.050 ;
        RECT 622.800 719.700 624.000 730.200 ;
        RECT 625.200 729.600 627.000 730.200 ;
        RECT 628.800 730.200 633.000 731.400 ;
        RECT 628.800 719.700 630.000 730.200 ;
        RECT 631.200 729.600 633.000 730.200 ;
        RECT 634.800 730.200 639.000 731.400 ;
        RECT 634.800 719.700 636.000 730.200 ;
        RECT 637.200 729.600 639.000 730.200 ;
        RECT 639.900 727.050 640.950 732.300 ;
        RECT 653.400 727.050 654.300 734.400 ;
        RECT 655.950 727.050 657.750 728.850 ;
        RECT 662.100 727.050 663.900 728.850 ;
        RECT 674.700 727.050 675.900 737.400 ;
        RECT 689.100 734.400 690.900 740.400 ;
        RECT 689.700 732.300 690.900 734.400 ;
        RECT 692.100 735.300 693.900 740.400 ;
        RECT 695.100 736.200 696.900 741.000 ;
        RECT 698.100 735.300 699.900 740.400 ;
        RECT 710.100 737.400 711.900 741.000 ;
        RECT 713.100 737.400 714.900 740.400 ;
        RECT 716.100 737.400 717.900 741.000 ;
        RECT 692.100 733.950 699.900 735.300 ;
        RECT 689.700 731.400 693.300 732.300 ;
        RECT 689.100 727.050 690.900 728.850 ;
        RECT 692.100 727.050 693.300 731.400 ;
        RECT 695.100 727.050 696.900 728.850 ;
        RECT 713.700 727.050 714.600 737.400 ;
        RECT 720.150 736.200 721.950 740.400 ;
        RECT 719.550 734.400 721.950 736.200 ;
        RECT 723.150 734.400 724.950 741.000 ;
        RECT 727.950 738.300 729.750 740.400 ;
        RECT 726.150 737.400 729.750 738.300 ;
        RECT 732.450 737.400 734.250 741.000 ;
        RECT 735.750 737.400 737.550 740.400 ;
        RECT 738.750 737.400 740.550 741.000 ;
        RECT 743.250 737.400 745.050 740.400 ;
        RECT 725.850 736.800 729.750 737.400 ;
        RECT 725.850 735.300 727.950 736.800 ;
        RECT 735.750 736.500 736.800 737.400 ;
        RECT 637.800 724.950 640.950 727.050 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 688.950 724.950 691.050 727.050 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 712.950 724.950 715.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 639.900 719.700 640.950 724.950 ;
        RECT 594.750 719.100 606.450 719.700 ;
        RECT 566.100 705.600 567.900 711.600 ;
        RECT 569.100 705.000 570.900 711.600 ;
        RECT 572.550 705.600 574.350 717.600 ;
        RECT 575.550 705.000 577.350 717.600 ;
        RECT 581.250 717.300 586.050 718.200 ;
        RECT 588.150 718.500 606.450 719.100 ;
        RECT 588.150 718.200 596.550 718.500 ;
        RECT 581.250 716.400 582.450 717.300 ;
        RECT 579.450 714.600 582.450 716.400 ;
        RECT 583.350 716.100 585.150 716.400 ;
        RECT 588.150 716.100 589.050 718.200 ;
        RECT 605.550 717.600 606.450 718.500 ;
        RECT 620.100 718.500 624.000 719.700 ;
        RECT 626.100 718.500 630.000 719.700 ;
        RECT 632.100 718.500 636.000 719.700 ;
        RECT 638.100 718.500 640.950 719.700 ;
        RECT 583.350 715.200 589.050 716.100 ;
        RECT 589.950 716.700 591.750 717.300 ;
        RECT 589.950 715.500 597.750 716.700 ;
        RECT 583.350 714.600 585.150 715.200 ;
        RECT 595.650 714.600 597.750 715.500 ;
        RECT 580.350 711.600 582.450 713.700 ;
        RECT 586.950 713.550 588.750 714.300 ;
        RECT 591.750 713.550 593.550 714.300 ;
        RECT 586.950 712.500 593.550 713.550 ;
        RECT 580.350 705.600 582.150 711.600 ;
        RECT 584.850 705.000 586.650 711.600 ;
        RECT 587.850 705.600 589.650 712.500 ;
        RECT 590.850 705.000 592.650 711.600 ;
        RECT 595.650 705.600 597.450 714.600 ;
        RECT 601.050 705.000 602.850 717.600 ;
        RECT 604.050 715.800 606.450 717.600 ;
        RECT 604.050 705.600 605.850 715.800 ;
        RECT 617.100 705.000 618.900 717.600 ;
        RECT 620.100 705.600 621.900 718.500 ;
        RECT 623.100 705.000 624.900 717.600 ;
        RECT 626.100 705.600 627.900 718.500 ;
        RECT 629.100 705.000 630.900 717.600 ;
        RECT 632.100 705.600 633.900 718.500 ;
        RECT 635.100 705.000 636.900 717.600 ;
        RECT 638.100 705.600 639.900 718.500 ;
        RECT 653.400 717.600 654.300 724.950 ;
        RECT 658.950 723.150 660.750 724.950 ;
        RECT 641.100 705.000 642.900 717.600 ;
        RECT 653.100 705.600 654.900 717.600 ;
        RECT 656.100 716.700 663.900 717.600 ;
        RECT 656.100 705.600 657.900 716.700 ;
        RECT 659.100 705.000 660.900 715.800 ;
        RECT 662.100 705.600 663.900 716.700 ;
        RECT 674.700 711.600 675.900 724.950 ;
        RECT 677.100 723.150 678.900 724.950 ;
        RECT 692.100 717.600 693.300 724.950 ;
        RECT 698.100 723.150 699.900 724.950 ;
        RECT 710.100 723.150 711.900 724.950 ;
        RECT 713.700 717.600 714.600 724.950 ;
        RECT 715.950 723.150 717.750 724.950 ;
        RECT 719.550 719.700 720.450 734.400 ;
        RECT 728.850 733.800 730.650 735.600 ;
        RECT 731.850 735.450 736.800 736.500 ;
        RECT 731.850 734.700 733.650 735.450 ;
        RECT 743.250 735.300 745.650 737.400 ;
        RECT 748.350 734.400 750.150 741.000 ;
        RECT 751.650 734.400 753.450 740.400 ;
        RECT 764.100 737.400 765.900 741.000 ;
        RECT 767.100 737.400 768.900 740.400 ;
        RECT 770.100 737.400 771.900 741.000 ;
        RECT 782.100 737.400 783.900 740.400 ;
        RECT 785.100 737.400 786.900 741.000 ;
        RECT 797.100 737.400 798.900 741.000 ;
        RECT 800.100 737.400 801.900 740.400 ;
        RECT 728.850 732.000 729.900 733.800 ;
        RECT 739.050 732.000 740.850 732.600 ;
        RECT 728.850 730.800 740.850 732.000 ;
        RECT 721.950 729.600 729.900 730.800 ;
        RECT 721.950 727.050 723.750 729.600 ;
        RECT 728.100 729.000 729.900 729.600 ;
        RECT 725.100 727.800 726.900 728.400 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 725.100 726.600 733.200 727.800 ;
        RECT 731.100 724.950 733.200 726.600 ;
        RECT 729.450 719.700 731.250 720.000 ;
        RECT 719.550 719.100 731.250 719.700 ;
        RECT 719.550 718.500 737.850 719.100 ;
        RECT 719.550 717.600 720.450 718.500 ;
        RECT 729.450 718.200 737.850 718.500 ;
        RECT 692.100 716.100 694.500 717.600 ;
        RECT 690.000 713.100 691.800 714.900 ;
        RECT 674.100 705.600 675.900 711.600 ;
        RECT 677.100 705.000 678.900 711.600 ;
        RECT 689.700 705.000 691.500 711.600 ;
        RECT 692.700 705.600 694.500 716.100 ;
        RECT 697.800 705.000 699.600 717.600 ;
        RECT 711.000 716.400 714.600 717.600 ;
        RECT 711.000 705.600 712.800 716.400 ;
        RECT 716.100 705.000 717.900 717.600 ;
        RECT 719.550 715.800 721.950 717.600 ;
        RECT 720.150 705.600 721.950 715.800 ;
        RECT 723.150 705.000 724.950 717.600 ;
        RECT 734.250 716.700 736.050 717.300 ;
        RECT 728.250 715.500 736.050 716.700 ;
        RECT 736.950 716.100 737.850 718.200 ;
        RECT 739.950 718.200 740.850 730.800 ;
        RECT 752.250 727.050 753.450 734.400 ;
        RECT 767.400 727.050 768.300 737.400 ;
        RECT 782.700 727.050 783.900 737.400 ;
        RECT 800.100 727.050 801.300 737.400 ;
        RECT 804.150 736.200 805.950 740.400 ;
        RECT 803.550 734.400 805.950 736.200 ;
        RECT 807.150 734.400 808.950 741.000 ;
        RECT 811.950 738.300 813.750 740.400 ;
        RECT 810.150 737.400 813.750 738.300 ;
        RECT 816.450 737.400 818.250 741.000 ;
        RECT 819.750 737.400 821.550 740.400 ;
        RECT 822.750 737.400 824.550 741.000 ;
        RECT 827.250 737.400 829.050 740.400 ;
        RECT 809.850 736.800 813.750 737.400 ;
        RECT 809.850 735.300 811.950 736.800 ;
        RECT 819.750 736.500 820.800 737.400 ;
        RECT 747.150 725.250 753.450 727.050 ;
        RECT 748.950 724.950 753.450 725.250 ;
        RECT 763.950 724.950 766.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 781.950 724.950 784.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 743.550 722.100 745.650 722.400 ;
        RECT 749.550 722.100 751.350 722.250 ;
        RECT 743.550 720.900 751.350 722.100 ;
        RECT 743.550 720.300 745.650 720.900 ;
        RECT 749.550 720.450 751.350 720.900 ;
        RECT 739.950 717.300 744.750 718.200 ;
        RECT 752.250 717.600 753.450 724.950 ;
        RECT 764.250 723.150 766.050 724.950 ;
        RECT 767.400 717.600 768.300 724.950 ;
        RECT 770.100 723.150 771.900 724.950 ;
        RECT 743.550 716.400 744.750 717.300 ;
        RECT 740.850 716.100 742.650 716.400 ;
        RECT 728.250 714.600 730.350 715.500 ;
        RECT 736.950 715.200 742.650 716.100 ;
        RECT 740.850 714.600 742.650 715.200 ;
        RECT 743.550 714.600 746.550 716.400 ;
        RECT 728.550 705.600 730.350 714.600 ;
        RECT 732.450 713.550 734.250 714.300 ;
        RECT 737.250 713.550 739.050 714.300 ;
        RECT 732.450 712.500 739.050 713.550 ;
        RECT 733.350 705.000 735.150 711.600 ;
        RECT 736.350 705.600 738.150 712.500 ;
        RECT 743.550 711.600 745.650 713.700 ;
        RECT 739.350 705.000 741.150 711.600 ;
        RECT 743.850 705.600 745.650 711.600 ;
        RECT 748.650 705.000 750.450 717.600 ;
        RECT 751.650 705.600 753.450 717.600 ;
        RECT 764.100 705.000 765.900 717.600 ;
        RECT 767.400 716.400 771.000 717.600 ;
        RECT 769.200 705.600 771.000 716.400 ;
        RECT 782.700 711.600 783.900 724.950 ;
        RECT 785.100 723.150 786.900 724.950 ;
        RECT 797.100 723.150 798.900 724.950 ;
        RECT 800.100 711.600 801.300 724.950 ;
        RECT 803.550 719.700 804.450 734.400 ;
        RECT 812.850 733.800 814.650 735.600 ;
        RECT 815.850 735.450 820.800 736.500 ;
        RECT 815.850 734.700 817.650 735.450 ;
        RECT 827.250 735.300 829.650 737.400 ;
        RECT 832.350 734.400 834.150 741.000 ;
        RECT 835.650 734.400 837.450 740.400 ;
        RECT 848.400 734.400 850.200 741.000 ;
        RECT 812.850 732.000 813.900 733.800 ;
        RECT 823.050 732.000 824.850 732.600 ;
        RECT 812.850 730.800 824.850 732.000 ;
        RECT 805.950 729.600 813.900 730.800 ;
        RECT 805.950 727.050 807.750 729.600 ;
        RECT 812.100 729.000 813.900 729.600 ;
        RECT 809.100 727.800 810.900 728.400 ;
        RECT 805.950 724.950 808.050 727.050 ;
        RECT 809.100 726.600 817.200 727.800 ;
        RECT 815.100 724.950 817.200 726.600 ;
        RECT 813.450 719.700 815.250 720.000 ;
        RECT 803.550 719.100 815.250 719.700 ;
        RECT 803.550 718.500 821.850 719.100 ;
        RECT 803.550 717.600 804.450 718.500 ;
        RECT 813.450 718.200 821.850 718.500 ;
        RECT 803.550 715.800 805.950 717.600 ;
        RECT 782.100 705.600 783.900 711.600 ;
        RECT 785.100 705.000 786.900 711.600 ;
        RECT 797.100 705.000 798.900 711.600 ;
        RECT 800.100 705.600 801.900 711.600 ;
        RECT 804.150 705.600 805.950 715.800 ;
        RECT 807.150 705.000 808.950 717.600 ;
        RECT 818.250 716.700 820.050 717.300 ;
        RECT 812.250 715.500 820.050 716.700 ;
        RECT 820.950 716.100 821.850 718.200 ;
        RECT 823.950 718.200 824.850 730.800 ;
        RECT 836.250 727.050 837.450 734.400 ;
        RECT 853.500 733.200 855.300 740.400 ;
        RECT 866.100 737.400 867.900 741.000 ;
        RECT 869.100 737.400 870.900 740.400 ;
        RECT 856.950 735.450 859.050 735.900 ;
        RECT 865.950 735.450 868.050 736.050 ;
        RECT 856.950 734.550 868.050 735.450 ;
        RECT 856.950 733.800 859.050 734.550 ;
        RECT 865.950 733.950 868.050 734.550 ;
        RECT 851.100 732.300 855.300 733.200 ;
        RECT 848.250 727.050 850.050 728.850 ;
        RECT 851.100 727.050 852.300 732.300 ;
        RECT 856.950 729.450 861.000 730.050 ;
        RECT 854.100 727.050 855.900 728.850 ;
        RECT 856.950 727.950 861.450 729.450 ;
        RECT 831.150 725.250 837.450 727.050 ;
        RECT 832.950 724.950 837.450 725.250 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 827.550 722.100 829.650 722.400 ;
        RECT 833.550 722.100 835.350 722.250 ;
        RECT 827.550 720.900 835.350 722.100 ;
        RECT 827.550 720.300 829.650 720.900 ;
        RECT 833.550 720.450 835.350 720.900 ;
        RECT 823.950 717.300 828.750 718.200 ;
        RECT 836.250 717.600 837.450 724.950 ;
        RECT 827.550 716.400 828.750 717.300 ;
        RECT 824.850 716.100 826.650 716.400 ;
        RECT 812.250 714.600 814.350 715.500 ;
        RECT 820.950 715.200 826.650 716.100 ;
        RECT 824.850 714.600 826.650 715.200 ;
        RECT 827.550 714.600 830.550 716.400 ;
        RECT 812.550 705.600 814.350 714.600 ;
        RECT 816.450 713.550 818.250 714.300 ;
        RECT 821.250 713.550 823.050 714.300 ;
        RECT 816.450 712.500 823.050 713.550 ;
        RECT 817.350 705.000 819.150 711.600 ;
        RECT 820.350 705.600 822.150 712.500 ;
        RECT 827.550 711.600 829.650 713.700 ;
        RECT 823.350 705.000 825.150 711.600 ;
        RECT 827.850 705.600 829.650 711.600 ;
        RECT 832.650 705.000 834.450 717.600 ;
        RECT 835.650 705.600 837.450 717.600 ;
        RECT 851.100 711.600 852.300 724.950 ;
        RECT 860.550 724.050 861.450 727.950 ;
        RECT 869.100 727.050 870.300 737.400 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 856.950 722.550 861.450 724.050 ;
        RECT 866.100 723.150 867.900 724.950 ;
        RECT 856.950 721.950 861.000 722.550 ;
        RECT 869.100 711.600 870.300 724.950 ;
        RECT 848.100 705.000 849.900 711.600 ;
        RECT 851.100 705.600 852.900 711.600 ;
        RECT 854.100 705.000 855.900 711.600 ;
        RECT 866.100 705.000 867.900 711.600 ;
        RECT 869.100 705.600 870.900 711.600 ;
        RECT 14.100 695.400 15.900 702.000 ;
        RECT 17.100 695.400 18.900 701.400 ;
        RECT 14.100 682.050 15.900 683.850 ;
        RECT 17.100 682.050 18.300 695.400 ;
        RECT 30.000 690.600 31.800 701.400 ;
        RECT 30.000 689.400 33.600 690.600 ;
        RECT 35.100 689.400 36.900 702.000 ;
        RECT 47.100 695.400 48.900 702.000 ;
        RECT 50.100 695.400 51.900 701.400 ;
        RECT 53.100 695.400 54.900 702.000 ;
        RECT 65.100 695.400 66.900 702.000 ;
        RECT 68.100 695.400 69.900 701.400 ;
        RECT 71.100 695.400 72.900 702.000 ;
        RECT 29.100 682.050 30.900 683.850 ;
        RECT 32.700 682.050 33.600 689.400 ;
        RECT 34.950 682.050 36.750 683.850 ;
        RECT 50.100 682.050 51.300 695.400 ;
        RECT 68.700 682.050 69.900 695.400 ;
        RECT 83.400 689.400 85.200 702.000 ;
        RECT 88.500 690.900 90.300 701.400 ;
        RECT 91.500 695.400 93.300 702.000 ;
        RECT 104.100 695.400 105.900 702.000 ;
        RECT 107.100 695.400 108.900 701.400 ;
        RECT 110.100 695.400 111.900 702.000 ;
        RECT 91.200 692.100 93.000 693.900 ;
        RECT 88.500 689.400 90.900 690.900 ;
        RECT 83.100 682.050 84.900 683.850 ;
        RECT 89.700 682.050 90.900 689.400 ;
        RECT 107.700 682.050 108.900 695.400 ;
        RECT 114.150 691.200 115.950 701.400 ;
        RECT 113.550 689.400 115.950 691.200 ;
        RECT 117.150 689.400 118.950 702.000 ;
        RECT 122.550 692.400 124.350 701.400 ;
        RECT 127.350 695.400 129.150 702.000 ;
        RECT 130.350 694.500 132.150 701.400 ;
        RECT 133.350 695.400 135.150 702.000 ;
        RECT 137.850 695.400 139.650 701.400 ;
        RECT 126.450 693.450 133.050 694.500 ;
        RECT 126.450 692.700 128.250 693.450 ;
        RECT 131.250 692.700 133.050 693.450 ;
        RECT 137.550 693.300 139.650 695.400 ;
        RECT 122.250 691.500 124.350 692.400 ;
        RECT 134.850 691.800 136.650 692.400 ;
        RECT 122.250 690.300 130.050 691.500 ;
        RECT 128.250 689.700 130.050 690.300 ;
        RECT 130.950 690.900 136.650 691.800 ;
        RECT 113.550 688.500 114.450 689.400 ;
        RECT 130.950 688.800 131.850 690.900 ;
        RECT 134.850 690.600 136.650 690.900 ;
        RECT 137.550 690.600 140.550 692.400 ;
        RECT 137.550 689.700 138.750 690.600 ;
        RECT 123.450 688.500 131.850 688.800 ;
        RECT 113.550 687.900 131.850 688.500 ;
        RECT 133.950 688.800 138.750 689.700 ;
        RECT 142.650 689.400 144.450 702.000 ;
        RECT 145.650 689.400 147.450 701.400 ;
        RECT 158.100 695.400 159.900 702.000 ;
        RECT 161.100 695.400 162.900 701.400 ;
        RECT 164.100 695.400 165.900 702.000 ;
        RECT 113.550 687.300 125.250 687.900 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 28.950 679.950 31.050 682.050 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 67.950 679.950 70.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 91.950 679.950 94.050 682.050 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 17.100 669.600 18.300 679.950 ;
        RECT 32.700 669.600 33.600 679.950 ;
        RECT 47.250 678.150 49.050 679.950 ;
        RECT 50.100 674.700 51.300 679.950 ;
        RECT 53.100 678.150 54.900 679.950 ;
        RECT 65.100 678.150 66.900 679.950 ;
        RECT 68.700 674.700 69.900 679.950 ;
        RECT 70.950 678.150 72.750 679.950 ;
        RECT 86.100 678.150 87.900 679.950 ;
        RECT 89.700 675.600 90.900 679.950 ;
        RECT 92.100 678.150 93.900 679.950 ;
        RECT 104.100 678.150 105.900 679.950 ;
        RECT 89.700 674.700 93.300 675.600 ;
        RECT 107.700 674.700 108.900 679.950 ;
        RECT 109.950 678.150 111.750 679.950 ;
        RECT 50.100 673.800 54.300 674.700 ;
        RECT 14.100 666.000 15.900 669.600 ;
        RECT 17.100 666.600 18.900 669.600 ;
        RECT 29.100 666.000 30.900 669.600 ;
        RECT 32.100 666.600 33.900 669.600 ;
        RECT 35.100 666.000 36.900 669.600 ;
        RECT 47.400 666.000 49.200 672.600 ;
        RECT 52.500 666.600 54.300 673.800 ;
        RECT 65.700 673.800 69.900 674.700 ;
        RECT 65.700 666.600 67.500 673.800 ;
        RECT 70.800 666.000 72.600 672.600 ;
        RECT 83.100 671.700 90.900 673.050 ;
        RECT 83.100 666.600 84.900 671.700 ;
        RECT 86.100 666.000 87.900 670.800 ;
        RECT 89.100 666.600 90.900 671.700 ;
        RECT 92.100 672.600 93.300 674.700 ;
        RECT 104.700 673.800 108.900 674.700 ;
        RECT 92.100 666.600 93.900 672.600 ;
        RECT 104.700 666.600 106.500 673.800 ;
        RECT 113.550 672.600 114.450 687.300 ;
        RECT 123.450 687.000 125.250 687.300 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 125.100 680.400 127.200 682.050 ;
        RECT 115.950 677.400 117.750 679.950 ;
        RECT 119.100 679.200 127.200 680.400 ;
        RECT 119.100 678.600 120.900 679.200 ;
        RECT 122.100 677.400 123.900 678.000 ;
        RECT 115.950 676.200 123.900 677.400 ;
        RECT 133.950 676.200 134.850 688.800 ;
        RECT 137.550 686.100 139.650 686.700 ;
        RECT 143.550 686.100 145.350 686.550 ;
        RECT 137.550 684.900 145.350 686.100 ;
        RECT 137.550 684.600 139.650 684.900 ;
        RECT 143.550 684.750 145.350 684.900 ;
        RECT 146.250 682.050 147.450 689.400 ;
        RECT 161.700 682.050 162.900 695.400 ;
        RECT 176.100 689.400 177.900 702.000 ;
        RECT 179.100 688.500 180.900 701.400 ;
        RECT 182.100 689.400 183.900 702.000 ;
        RECT 185.100 689.400 186.900 701.400 ;
        RECT 188.100 689.400 189.900 702.000 ;
        RECT 200.100 689.400 201.900 701.400 ;
        RECT 203.100 691.200 204.900 702.000 ;
        RECT 206.100 695.400 207.900 701.400 ;
        RECT 218.100 695.400 219.900 701.400 ;
        RECT 221.100 695.400 222.900 702.000 ;
        RECT 185.100 688.500 186.300 689.400 ;
        RECT 179.100 687.600 186.300 688.500 ;
        RECT 179.100 682.050 180.900 683.850 ;
        RECT 185.100 682.050 186.300 687.600 ;
        RECT 200.100 682.050 201.300 689.400 ;
        RECT 206.700 688.500 207.900 695.400 ;
        RECT 202.200 687.600 207.900 688.500 ;
        RECT 202.200 686.700 204.000 687.600 ;
        RECT 142.950 681.750 147.450 682.050 ;
        RECT 141.150 679.950 147.450 681.750 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 179.100 679.950 181.200 682.050 ;
        RECT 185.100 679.950 187.200 682.050 ;
        RECT 200.100 679.950 202.200 682.050 ;
        RECT 122.850 675.000 134.850 676.200 ;
        RECT 122.850 673.200 123.900 675.000 ;
        RECT 133.050 674.400 134.850 675.000 ;
        RECT 109.800 666.000 111.600 672.600 ;
        RECT 113.550 670.800 115.950 672.600 ;
        RECT 114.150 666.600 115.950 670.800 ;
        RECT 117.150 666.000 118.950 672.600 ;
        RECT 119.850 670.200 121.950 671.700 ;
        RECT 122.850 671.400 124.650 673.200 ;
        RECT 146.250 672.600 147.450 679.950 ;
        RECT 158.100 678.150 159.900 679.950 ;
        RECT 161.700 674.700 162.900 679.950 ;
        RECT 163.950 678.150 165.750 679.950 ;
        RECT 185.100 674.700 186.300 679.950 ;
        RECT 125.850 671.550 127.650 672.300 ;
        RECT 125.850 670.500 130.800 671.550 ;
        RECT 119.850 669.600 123.750 670.200 ;
        RECT 129.750 669.600 130.800 670.500 ;
        RECT 137.250 669.600 139.650 671.700 ;
        RECT 120.150 668.700 123.750 669.600 ;
        RECT 121.950 666.600 123.750 668.700 ;
        RECT 126.450 666.000 128.250 669.600 ;
        RECT 129.750 666.600 131.550 669.600 ;
        RECT 132.750 666.000 134.550 669.600 ;
        RECT 137.250 666.600 139.050 669.600 ;
        RECT 142.350 666.000 144.150 672.600 ;
        RECT 145.650 666.600 147.450 672.600 ;
        RECT 158.700 673.800 162.900 674.700 ;
        RECT 158.700 666.600 160.500 673.800 ;
        RECT 179.100 673.500 186.300 674.700 ;
        RECT 179.100 672.600 180.300 673.500 ;
        RECT 185.100 672.600 186.300 673.500 ;
        RECT 200.100 672.600 201.300 679.950 ;
        RECT 203.100 675.300 204.000 686.700 ;
        RECT 205.800 682.050 207.600 683.850 ;
        RECT 218.700 682.050 219.900 695.400 ;
        RECT 234.000 690.600 235.800 701.400 ;
        RECT 234.000 689.400 237.600 690.600 ;
        RECT 239.100 689.400 240.900 702.000 ;
        RECT 251.100 695.400 252.900 702.000 ;
        RECT 254.100 695.400 255.900 701.400 ;
        RECT 223.950 684.450 228.000 685.050 ;
        RECT 221.100 682.050 222.900 683.850 ;
        RECT 223.950 682.950 228.450 684.450 ;
        RECT 205.500 679.950 207.600 682.050 ;
        RECT 217.950 679.950 220.050 682.050 ;
        RECT 220.950 679.950 223.050 682.050 ;
        RECT 202.200 674.400 204.000 675.300 ;
        RECT 202.200 673.500 207.900 674.400 ;
        RECT 163.800 666.000 165.600 672.600 ;
        RECT 176.100 666.000 177.900 672.600 ;
        RECT 179.100 666.600 180.900 672.600 ;
        RECT 182.100 666.000 183.900 672.600 ;
        RECT 185.100 666.600 186.900 672.600 ;
        RECT 188.100 666.000 189.900 672.600 ;
        RECT 200.100 666.600 201.900 672.600 ;
        RECT 203.100 666.000 204.900 672.600 ;
        RECT 206.700 669.600 207.900 673.500 ;
        RECT 218.700 669.600 219.900 679.950 ;
        RECT 227.550 679.050 228.450 682.950 ;
        RECT 233.100 682.050 234.900 683.850 ;
        RECT 236.700 682.050 237.600 689.400 ;
        RECT 241.950 684.450 244.050 688.050 ;
        RECT 241.950 684.000 246.450 684.450 ;
        RECT 238.950 682.050 240.750 683.850 ;
        RECT 242.550 683.550 246.450 684.000 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 238.950 679.950 241.050 682.050 ;
        RECT 227.550 677.550 232.050 679.050 ;
        RECT 228.000 676.950 232.050 677.550 ;
        RECT 236.700 669.600 237.600 679.950 ;
        RECT 245.550 679.050 246.450 683.550 ;
        RECT 251.100 682.050 252.900 683.850 ;
        RECT 254.100 682.050 255.300 695.400 ;
        RECT 266.400 689.400 268.200 702.000 ;
        RECT 271.500 690.900 273.300 701.400 ;
        RECT 274.500 695.400 276.300 702.000 ;
        RECT 274.200 692.100 276.000 693.900 ;
        RECT 271.500 689.400 273.900 690.900 ;
        RECT 287.100 689.400 288.900 702.000 ;
        RECT 292.200 690.600 294.000 701.400 ;
        RECT 308.100 695.400 309.900 702.000 ;
        RECT 311.100 695.400 312.900 701.400 ;
        RECT 314.100 695.400 315.900 702.000 ;
        RECT 290.400 689.400 294.000 690.600 ;
        RECT 259.950 687.450 262.050 688.050 ;
        RECT 268.950 687.450 271.050 688.050 ;
        RECT 259.950 686.550 271.050 687.450 ;
        RECT 259.950 685.950 262.050 686.550 ;
        RECT 268.950 685.950 271.050 686.550 ;
        RECT 256.950 684.450 261.000 685.050 ;
        RECT 256.950 682.950 261.450 684.450 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 245.550 677.550 250.050 679.050 ;
        RECT 246.000 676.950 250.050 677.550 ;
        RECT 254.100 669.600 255.300 679.950 ;
        RECT 260.550 678.900 261.450 682.950 ;
        RECT 266.100 682.050 267.900 683.850 ;
        RECT 272.700 682.050 273.900 689.400 ;
        RECT 287.250 682.050 289.050 683.850 ;
        RECT 290.400 682.050 291.300 689.400 ;
        RECT 293.100 682.050 294.900 683.850 ;
        RECT 311.700 682.050 312.900 695.400 ;
        RECT 318.150 691.200 319.950 701.400 ;
        RECT 317.550 689.400 319.950 691.200 ;
        RECT 321.150 689.400 322.950 702.000 ;
        RECT 326.550 692.400 328.350 701.400 ;
        RECT 331.350 695.400 333.150 702.000 ;
        RECT 334.350 694.500 336.150 701.400 ;
        RECT 337.350 695.400 339.150 702.000 ;
        RECT 341.850 695.400 343.650 701.400 ;
        RECT 330.450 693.450 337.050 694.500 ;
        RECT 330.450 692.700 332.250 693.450 ;
        RECT 335.250 692.700 337.050 693.450 ;
        RECT 341.550 693.300 343.650 695.400 ;
        RECT 326.250 691.500 328.350 692.400 ;
        RECT 338.850 691.800 340.650 692.400 ;
        RECT 326.250 690.300 334.050 691.500 ;
        RECT 332.250 689.700 334.050 690.300 ;
        RECT 334.950 690.900 340.650 691.800 ;
        RECT 317.550 688.500 318.450 689.400 ;
        RECT 334.950 688.800 335.850 690.900 ;
        RECT 338.850 690.600 340.650 690.900 ;
        RECT 341.550 690.600 344.550 692.400 ;
        RECT 341.550 689.700 342.750 690.600 ;
        RECT 327.450 688.500 335.850 688.800 ;
        RECT 317.550 687.900 335.850 688.500 ;
        RECT 337.950 688.800 342.750 689.700 ;
        RECT 346.650 689.400 348.450 702.000 ;
        RECT 349.650 689.400 351.450 701.400 ;
        RECT 362.100 695.400 363.900 702.000 ;
        RECT 365.100 695.400 366.900 701.400 ;
        RECT 368.100 695.400 369.900 702.000 ;
        RECT 380.700 695.400 382.500 702.000 ;
        RECT 317.550 687.300 329.250 687.900 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 268.950 679.950 271.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 274.950 679.950 277.050 682.050 ;
        RECT 286.950 679.950 289.050 682.050 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 259.950 676.800 262.050 678.900 ;
        RECT 269.100 678.150 270.900 679.950 ;
        RECT 272.700 675.600 273.900 679.950 ;
        RECT 275.100 678.150 276.900 679.950 ;
        RECT 272.700 674.700 276.300 675.600 ;
        RECT 266.100 671.700 273.900 673.050 ;
        RECT 206.100 666.600 207.900 669.600 ;
        RECT 218.100 666.600 219.900 669.600 ;
        RECT 221.100 666.000 222.900 669.600 ;
        RECT 233.100 666.000 234.900 669.600 ;
        RECT 236.100 666.600 237.900 669.600 ;
        RECT 239.100 666.000 240.900 669.600 ;
        RECT 251.100 666.000 252.900 669.600 ;
        RECT 254.100 666.600 255.900 669.600 ;
        RECT 266.100 666.600 267.900 671.700 ;
        RECT 269.100 666.000 270.900 670.800 ;
        RECT 272.100 666.600 273.900 671.700 ;
        RECT 275.100 672.600 276.300 674.700 ;
        RECT 275.100 666.600 276.900 672.600 ;
        RECT 290.400 669.600 291.300 679.950 ;
        RECT 308.100 678.150 309.900 679.950 ;
        RECT 311.700 674.700 312.900 679.950 ;
        RECT 313.950 678.150 315.750 679.950 ;
        RECT 308.700 673.800 312.900 674.700 ;
        RECT 287.100 666.000 288.900 669.600 ;
        RECT 290.100 666.600 291.900 669.600 ;
        RECT 293.100 666.000 294.900 669.600 ;
        RECT 308.700 666.600 310.500 673.800 ;
        RECT 317.550 672.600 318.450 687.300 ;
        RECT 327.450 687.000 329.250 687.300 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 329.100 680.400 331.200 682.050 ;
        RECT 319.950 677.400 321.750 679.950 ;
        RECT 323.100 679.200 331.200 680.400 ;
        RECT 323.100 678.600 324.900 679.200 ;
        RECT 326.100 677.400 327.900 678.000 ;
        RECT 319.950 676.200 327.900 677.400 ;
        RECT 337.950 676.200 338.850 688.800 ;
        RECT 341.550 686.100 343.650 686.700 ;
        RECT 347.550 686.100 349.350 686.550 ;
        RECT 341.550 684.900 349.350 686.100 ;
        RECT 341.550 684.600 343.650 684.900 ;
        RECT 347.550 684.750 349.350 684.900 ;
        RECT 350.250 682.050 351.450 689.400 ;
        RECT 352.950 687.450 355.050 688.050 ;
        RECT 361.950 687.450 364.050 688.050 ;
        RECT 352.950 686.550 364.050 687.450 ;
        RECT 352.950 685.950 355.050 686.550 ;
        RECT 361.950 685.950 364.050 686.550 ;
        RECT 365.100 682.050 366.300 695.400 ;
        RECT 381.000 692.100 382.800 693.900 ;
        RECT 383.700 690.900 385.500 701.400 ;
        RECT 383.100 689.400 385.500 690.900 ;
        RECT 388.800 689.400 390.600 702.000 ;
        RECT 401.700 695.400 403.500 702.000 ;
        RECT 402.000 692.100 403.800 693.900 ;
        RECT 404.700 690.900 406.500 701.400 ;
        RECT 404.100 689.400 406.500 690.900 ;
        RECT 409.800 689.400 411.600 702.000 ;
        RECT 425.100 689.400 426.900 701.400 ;
        RECT 428.100 690.000 429.900 702.000 ;
        RECT 431.100 695.400 432.900 701.400 ;
        RECT 434.100 695.400 435.900 702.000 ;
        RECT 383.100 682.050 384.300 689.400 ;
        RECT 385.950 687.450 388.050 688.050 ;
        RECT 400.950 687.450 403.050 688.200 ;
        RECT 385.950 686.550 403.050 687.450 ;
        RECT 385.950 685.950 388.050 686.550 ;
        RECT 400.950 686.100 403.050 686.550 ;
        RECT 389.100 682.050 390.900 683.850 ;
        RECT 404.100 682.050 405.300 689.400 ;
        RECT 410.100 682.050 411.900 683.850 ;
        RECT 425.700 682.050 426.600 689.400 ;
        RECT 429.000 682.050 430.800 683.850 ;
        RECT 346.950 681.750 351.450 682.050 ;
        RECT 345.150 679.950 351.450 681.750 ;
        RECT 361.950 679.950 364.050 682.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 379.950 679.950 382.050 682.050 ;
        RECT 382.950 679.950 385.050 682.050 ;
        RECT 385.950 679.950 388.050 682.050 ;
        RECT 388.950 679.950 391.050 682.050 ;
        RECT 400.950 679.950 403.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 406.950 679.950 409.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 425.100 679.950 427.200 682.050 ;
        RECT 428.400 679.950 430.500 682.050 ;
        RECT 326.850 675.000 338.850 676.200 ;
        RECT 326.850 673.200 327.900 675.000 ;
        RECT 337.050 674.400 338.850 675.000 ;
        RECT 313.800 666.000 315.600 672.600 ;
        RECT 317.550 670.800 319.950 672.600 ;
        RECT 318.150 666.600 319.950 670.800 ;
        RECT 321.150 666.000 322.950 672.600 ;
        RECT 323.850 670.200 325.950 671.700 ;
        RECT 326.850 671.400 328.650 673.200 ;
        RECT 350.250 672.600 351.450 679.950 ;
        RECT 362.250 678.150 364.050 679.950 ;
        RECT 365.100 674.700 366.300 679.950 ;
        RECT 368.100 678.150 369.900 679.950 ;
        RECT 380.100 678.150 381.900 679.950 ;
        RECT 383.100 675.600 384.300 679.950 ;
        RECT 386.100 678.150 387.900 679.950 ;
        RECT 401.100 678.150 402.900 679.950 ;
        RECT 404.100 675.600 405.300 679.950 ;
        RECT 407.100 678.150 408.900 679.950 ;
        RECT 380.700 674.700 384.300 675.600 ;
        RECT 401.700 674.700 405.300 675.600 ;
        RECT 365.100 673.800 369.300 674.700 ;
        RECT 357.000 672.900 361.050 673.050 ;
        RECT 329.850 671.550 331.650 672.300 ;
        RECT 329.850 670.500 334.800 671.550 ;
        RECT 323.850 669.600 327.750 670.200 ;
        RECT 333.750 669.600 334.800 670.500 ;
        RECT 341.250 669.600 343.650 671.700 ;
        RECT 324.150 668.700 327.750 669.600 ;
        RECT 325.950 666.600 327.750 668.700 ;
        RECT 330.450 666.000 332.250 669.600 ;
        RECT 333.750 666.600 335.550 669.600 ;
        RECT 336.750 666.000 338.550 669.600 ;
        RECT 341.250 666.600 343.050 669.600 ;
        RECT 346.350 666.000 348.150 672.600 ;
        RECT 349.650 666.600 351.450 672.600 ;
        RECT 355.950 670.950 361.050 672.900 ;
        RECT 355.950 670.800 358.050 670.950 ;
        RECT 362.400 666.000 364.200 672.600 ;
        RECT 367.500 666.600 369.300 673.800 ;
        RECT 380.700 672.600 381.900 674.700 ;
        RECT 380.100 666.600 381.900 672.600 ;
        RECT 383.100 671.700 390.900 673.050 ;
        RECT 401.700 672.600 402.900 674.700 ;
        RECT 383.100 666.600 384.900 671.700 ;
        RECT 386.100 666.000 387.900 670.800 ;
        RECT 389.100 666.600 390.900 671.700 ;
        RECT 401.100 666.600 402.900 672.600 ;
        RECT 404.100 671.700 411.900 673.050 ;
        RECT 404.100 666.600 405.900 671.700 ;
        RECT 407.100 666.000 408.900 670.800 ;
        RECT 410.100 666.600 411.900 671.700 ;
        RECT 425.700 672.600 426.600 679.950 ;
        RECT 432.000 675.300 432.900 695.400 ;
        RECT 446.100 689.400 447.900 701.400 ;
        RECT 449.100 691.200 450.900 702.000 ;
        RECT 452.100 695.400 453.900 701.400 ;
        RECT 446.100 682.050 447.300 689.400 ;
        RECT 452.700 688.500 453.900 695.400 ;
        RECT 467.400 689.400 469.200 702.000 ;
        RECT 472.500 690.900 474.300 701.400 ;
        RECT 475.500 695.400 477.300 702.000 ;
        RECT 488.100 695.400 489.900 702.000 ;
        RECT 491.100 695.400 492.900 701.400 ;
        RECT 503.100 695.400 504.900 702.000 ;
        RECT 506.100 695.400 507.900 701.400 ;
        RECT 509.100 695.400 510.900 702.000 ;
        RECT 524.700 695.400 526.500 702.000 ;
        RECT 475.200 692.100 477.000 693.900 ;
        RECT 472.500 689.400 474.900 690.900 ;
        RECT 448.200 687.600 453.900 688.500 ;
        RECT 448.200 686.700 450.000 687.600 ;
        RECT 433.800 679.950 435.900 682.050 ;
        RECT 446.100 679.950 448.200 682.050 ;
        RECT 433.950 678.150 435.750 679.950 ;
        RECT 427.500 674.400 435.900 675.300 ;
        RECT 427.500 673.500 429.300 674.400 ;
        RECT 425.700 670.800 428.400 672.600 ;
        RECT 426.600 666.600 428.400 670.800 ;
        RECT 429.600 666.000 431.400 672.600 ;
        RECT 434.100 666.600 435.900 674.400 ;
        RECT 446.100 672.600 447.300 679.950 ;
        RECT 449.100 675.300 450.000 686.700 ;
        RECT 451.800 682.050 453.600 683.850 ;
        RECT 467.100 682.050 468.900 683.850 ;
        RECT 473.700 682.050 474.900 689.400 ;
        RECT 480.000 684.900 483.000 685.050 ;
        RECT 478.950 684.450 483.000 684.900 ;
        RECT 478.950 682.950 483.450 684.450 ;
        RECT 478.950 682.800 481.050 682.950 ;
        RECT 451.500 679.950 453.600 682.050 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 472.950 679.950 475.050 682.050 ;
        RECT 475.950 679.950 478.050 682.050 ;
        RECT 470.100 678.150 471.900 679.950 ;
        RECT 448.200 674.400 450.000 675.300 ;
        RECT 473.700 675.600 474.900 679.950 ;
        RECT 476.100 678.150 477.900 679.950 ;
        RECT 482.550 679.050 483.450 682.950 ;
        RECT 488.100 682.050 489.900 683.850 ;
        RECT 491.100 682.050 492.300 695.400 ;
        RECT 506.100 682.050 507.300 695.400 ;
        RECT 525.000 692.100 526.800 693.900 ;
        RECT 527.700 690.900 529.500 701.400 ;
        RECT 527.100 689.400 529.500 690.900 ;
        RECT 532.800 689.400 534.600 702.000 ;
        RECT 536.550 689.400 538.350 701.400 ;
        RECT 539.550 689.400 541.350 702.000 ;
        RECT 544.350 695.400 546.150 701.400 ;
        RECT 548.850 695.400 550.650 702.000 ;
        RECT 544.350 693.300 546.450 695.400 ;
        RECT 551.850 694.500 553.650 701.400 ;
        RECT 554.850 695.400 556.650 702.000 ;
        RECT 550.950 693.450 557.550 694.500 ;
        RECT 550.950 692.700 552.750 693.450 ;
        RECT 555.750 692.700 557.550 693.450 ;
        RECT 559.650 692.400 561.450 701.400 ;
        RECT 543.450 690.600 546.450 692.400 ;
        RECT 547.350 691.800 549.150 692.400 ;
        RECT 547.350 690.900 553.050 691.800 ;
        RECT 559.650 691.500 561.750 692.400 ;
        RECT 547.350 690.600 549.150 690.900 ;
        RECT 545.250 689.700 546.450 690.600 ;
        RECT 519.000 684.450 523.050 685.050 ;
        RECT 518.550 682.950 523.050 684.450 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 490.950 679.950 493.050 682.050 ;
        RECT 502.950 679.950 505.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 508.950 679.950 511.050 682.050 ;
        RECT 478.950 677.550 483.450 679.050 ;
        RECT 478.950 676.950 483.000 677.550 ;
        RECT 473.700 674.700 477.300 675.600 ;
        RECT 448.200 673.500 453.900 674.400 ;
        RECT 446.100 666.600 447.900 672.600 ;
        RECT 449.100 666.000 450.900 672.600 ;
        RECT 452.700 669.600 453.900 673.500 ;
        RECT 452.100 666.600 453.900 669.600 ;
        RECT 467.100 671.700 474.900 673.050 ;
        RECT 467.100 666.600 468.900 671.700 ;
        RECT 470.100 666.000 471.900 670.800 ;
        RECT 473.100 666.600 474.900 671.700 ;
        RECT 476.100 672.600 477.300 674.700 ;
        RECT 476.100 666.600 477.900 672.600 ;
        RECT 491.100 669.600 492.300 679.950 ;
        RECT 503.250 678.150 505.050 679.950 ;
        RECT 506.100 674.700 507.300 679.950 ;
        RECT 509.100 678.150 510.900 679.950 ;
        RECT 511.950 678.450 514.050 679.050 ;
        RECT 518.550 678.450 519.450 682.950 ;
        RECT 527.100 682.050 528.300 689.400 ;
        RECT 533.100 682.050 534.900 683.850 ;
        RECT 536.550 682.050 537.750 689.400 ;
        RECT 545.250 688.800 550.050 689.700 ;
        RECT 538.650 686.100 540.450 686.550 ;
        RECT 544.350 686.100 546.450 686.700 ;
        RECT 538.650 684.900 546.450 686.100 ;
        RECT 538.650 684.750 540.450 684.900 ;
        RECT 544.350 684.600 546.450 684.900 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 526.950 679.950 529.050 682.050 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 536.550 681.750 541.050 682.050 ;
        RECT 536.550 679.950 542.850 681.750 ;
        RECT 511.950 677.550 519.450 678.450 ;
        RECT 524.100 678.150 525.900 679.950 ;
        RECT 511.950 676.950 514.050 677.550 ;
        RECT 527.100 675.600 528.300 679.950 ;
        RECT 530.100 678.150 531.900 679.950 ;
        RECT 524.700 674.700 528.300 675.600 ;
        RECT 506.100 673.800 510.300 674.700 ;
        RECT 488.100 666.000 489.900 669.600 ;
        RECT 491.100 666.600 492.900 669.600 ;
        RECT 503.400 666.000 505.200 672.600 ;
        RECT 508.500 666.600 510.300 673.800 ;
        RECT 524.700 672.600 525.900 674.700 ;
        RECT 524.100 666.600 525.900 672.600 ;
        RECT 527.100 671.700 534.900 673.050 ;
        RECT 527.100 666.600 528.900 671.700 ;
        RECT 530.100 666.000 531.900 670.800 ;
        RECT 533.100 666.600 534.900 671.700 ;
        RECT 536.550 672.600 537.750 679.950 ;
        RECT 549.150 676.200 550.050 688.800 ;
        RECT 552.150 688.800 553.050 690.900 ;
        RECT 553.950 690.300 561.750 691.500 ;
        RECT 553.950 689.700 555.750 690.300 ;
        RECT 565.050 689.400 566.850 702.000 ;
        RECT 568.050 691.200 569.850 701.400 ;
        RECT 568.050 689.400 570.450 691.200 ;
        RECT 582.000 690.600 583.800 701.400 ;
        RECT 582.000 689.400 585.600 690.600 ;
        RECT 587.100 689.400 588.900 702.000 ;
        RECT 600.000 690.600 601.800 701.400 ;
        RECT 600.000 689.400 603.600 690.600 ;
        RECT 605.100 689.400 606.900 702.000 ;
        RECT 617.100 690.300 618.900 701.400 ;
        RECT 620.100 691.500 621.900 702.000 ;
        RECT 617.100 689.400 621.600 690.300 ;
        RECT 624.600 689.400 626.400 701.400 ;
        RECT 629.100 691.500 630.900 702.000 ;
        RECT 632.100 690.600 633.900 701.400 ;
        RECT 644.100 695.400 645.900 701.400 ;
        RECT 647.100 695.400 648.900 702.000 ;
        RECT 659.100 695.400 660.900 702.000 ;
        RECT 662.100 695.400 663.900 701.400 ;
        RECT 665.100 695.400 666.900 702.000 ;
        RECT 552.150 688.500 560.550 688.800 ;
        RECT 569.550 688.500 570.450 689.400 ;
        RECT 552.150 687.900 570.450 688.500 ;
        RECT 558.750 687.300 570.450 687.900 ;
        RECT 558.750 687.000 560.550 687.300 ;
        RECT 556.800 680.400 558.900 682.050 ;
        RECT 556.800 679.200 564.900 680.400 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 563.100 678.600 564.900 679.200 ;
        RECT 560.100 677.400 561.900 678.000 ;
        RECT 566.250 677.400 568.050 679.950 ;
        RECT 560.100 676.200 568.050 677.400 ;
        RECT 549.150 675.000 561.150 676.200 ;
        RECT 549.150 674.400 550.950 675.000 ;
        RECT 560.100 673.200 561.150 675.000 ;
        RECT 536.550 666.600 538.350 672.600 ;
        RECT 539.850 666.000 541.650 672.600 ;
        RECT 544.350 669.600 546.750 671.700 ;
        RECT 556.350 671.550 558.150 672.300 ;
        RECT 553.200 670.500 558.150 671.550 ;
        RECT 559.350 671.400 561.150 673.200 ;
        RECT 569.550 672.600 570.450 687.300 ;
        RECT 581.100 682.050 582.900 683.850 ;
        RECT 584.700 682.050 585.600 689.400 ;
        RECT 589.950 684.450 594.000 685.050 ;
        RECT 586.950 682.050 588.750 683.850 ;
        RECT 589.950 682.950 594.450 684.450 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 553.200 669.600 554.250 670.500 ;
        RECT 562.050 670.200 564.150 671.700 ;
        RECT 560.250 669.600 564.150 670.200 ;
        RECT 544.950 666.600 546.750 669.600 ;
        RECT 549.450 666.000 551.250 669.600 ;
        RECT 552.450 666.600 554.250 669.600 ;
        RECT 555.750 666.000 557.550 669.600 ;
        RECT 560.250 668.700 563.850 669.600 ;
        RECT 560.250 666.600 562.050 668.700 ;
        RECT 565.050 666.000 566.850 672.600 ;
        RECT 568.050 670.800 570.450 672.600 ;
        RECT 568.050 666.600 569.850 670.800 ;
        RECT 584.700 669.600 585.600 679.950 ;
        RECT 593.550 679.050 594.450 682.950 ;
        RECT 599.100 682.050 600.900 683.850 ;
        RECT 602.700 682.050 603.600 689.400 ;
        RECT 619.500 687.300 621.600 689.400 ;
        RECT 625.200 688.050 626.400 689.400 ;
        RECT 629.100 689.400 633.900 690.600 ;
        RECT 629.100 688.500 631.200 689.400 ;
        RECT 625.200 687.000 626.700 688.050 ;
        RECT 622.800 685.500 624.900 685.800 ;
        RECT 604.950 682.050 606.750 683.850 ;
        RECT 621.000 683.700 624.900 685.500 ;
        RECT 625.800 685.050 626.700 687.000 ;
        RECT 625.800 682.950 627.900 685.050 ;
        RECT 634.950 684.450 637.050 685.050 ;
        RECT 640.950 684.450 643.050 685.050 ;
        RECT 625.800 682.800 627.300 682.950 ;
        RECT 622.200 682.050 624.000 682.500 ;
        RECT 598.950 679.950 601.050 682.050 ;
        RECT 601.950 679.950 604.050 682.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 617.100 680.700 624.000 682.050 ;
        RECT 624.900 681.900 627.300 682.800 ;
        RECT 631.800 682.050 633.600 683.850 ;
        RECT 634.950 683.550 643.050 684.450 ;
        RECT 634.950 682.950 637.050 683.550 ;
        RECT 640.950 682.950 643.050 683.550 ;
        RECT 644.700 682.050 645.900 695.400 ;
        RECT 647.100 682.050 648.900 683.850 ;
        RECT 662.700 682.050 663.900 695.400 ;
        RECT 664.950 690.450 667.050 691.050 ;
        RECT 676.950 690.450 679.050 691.050 ;
        RECT 664.950 689.550 679.050 690.450 ;
        RECT 664.950 688.950 667.050 689.550 ;
        RECT 676.950 688.950 679.050 689.550 ;
        RECT 680.400 689.400 682.200 702.000 ;
        RECT 685.500 690.900 687.300 701.400 ;
        RECT 688.500 695.400 690.300 702.000 ;
        RECT 688.200 692.100 690.000 693.900 ;
        RECT 685.500 689.400 687.900 690.900 ;
        RECT 702.000 690.600 703.800 701.400 ;
        RECT 702.000 689.400 705.600 690.600 ;
        RECT 707.100 689.400 708.900 702.000 ;
        RECT 719.100 689.400 720.900 702.000 ;
        RECT 724.200 690.600 726.000 701.400 ;
        RECT 722.400 689.400 726.000 690.600 ;
        RECT 737.100 689.400 738.900 701.400 ;
        RECT 740.100 690.300 741.900 701.400 ;
        RECT 743.100 691.200 744.900 702.000 ;
        RECT 746.100 690.300 747.900 701.400 ;
        RECT 740.100 689.400 747.900 690.300 ;
        RECT 761.100 689.400 762.900 702.000 ;
        RECT 766.200 690.600 768.000 701.400 ;
        RECT 771.150 691.200 772.950 701.400 ;
        RECT 764.400 689.400 768.000 690.600 ;
        RECT 770.550 689.400 772.950 691.200 ;
        RECT 774.150 689.400 775.950 702.000 ;
        RECT 779.550 692.400 781.350 701.400 ;
        RECT 784.350 695.400 786.150 702.000 ;
        RECT 787.350 694.500 789.150 701.400 ;
        RECT 790.350 695.400 792.150 702.000 ;
        RECT 794.850 695.400 796.650 701.400 ;
        RECT 783.450 693.450 790.050 694.500 ;
        RECT 783.450 692.700 785.250 693.450 ;
        RECT 788.250 692.700 790.050 693.450 ;
        RECT 794.550 693.300 796.650 695.400 ;
        RECT 779.250 691.500 781.350 692.400 ;
        RECT 791.850 691.800 793.650 692.400 ;
        RECT 779.250 690.300 787.050 691.500 ;
        RECT 785.250 689.700 787.050 690.300 ;
        RECT 787.950 690.900 793.650 691.800 ;
        RECT 682.950 687.450 685.050 688.050 ;
        RECT 677.550 686.550 685.050 687.450 ;
        RECT 667.950 684.450 672.000 685.050 ;
        RECT 677.550 684.450 678.450 686.550 ;
        RECT 682.950 685.950 685.050 686.550 ;
        RECT 667.950 682.950 672.450 684.450 ;
        RECT 617.100 679.950 619.200 680.700 ;
        RECT 593.550 677.550 598.050 679.050 ;
        RECT 594.000 676.950 598.050 677.550 ;
        RECT 586.950 672.450 589.050 673.050 ;
        RECT 598.950 672.450 601.050 673.050 ;
        RECT 586.950 671.550 601.050 672.450 ;
        RECT 586.950 670.950 589.050 671.550 ;
        RECT 598.950 670.950 601.050 671.550 ;
        RECT 602.700 669.600 603.600 679.950 ;
        RECT 617.400 678.150 619.200 679.950 ;
        RECT 622.200 677.400 624.000 679.200 ;
        RECT 621.900 675.300 624.000 677.400 ;
        RECT 617.700 674.400 624.000 675.300 ;
        RECT 624.900 676.200 626.100 681.900 ;
        RECT 627.300 679.200 629.100 681.000 ;
        RECT 631.800 679.950 633.900 682.050 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 661.950 679.950 664.050 682.050 ;
        RECT 664.950 679.950 667.050 682.050 ;
        RECT 627.000 677.100 629.100 679.200 ;
        RECT 617.700 672.600 618.900 674.400 ;
        RECT 624.900 674.100 627.900 676.200 ;
        RECT 624.900 672.600 626.100 674.100 ;
        RECT 629.100 673.500 631.200 674.700 ;
        RECT 629.100 672.600 633.900 673.500 ;
        RECT 581.100 666.000 582.900 669.600 ;
        RECT 584.100 666.600 585.900 669.600 ;
        RECT 587.100 666.000 588.900 669.600 ;
        RECT 599.100 666.000 600.900 669.600 ;
        RECT 602.100 666.600 603.900 669.600 ;
        RECT 605.100 666.000 606.900 669.600 ;
        RECT 617.100 666.600 618.900 672.600 ;
        RECT 620.100 666.000 621.900 671.700 ;
        RECT 624.600 666.600 626.400 672.600 ;
        RECT 629.100 666.000 630.900 671.700 ;
        RECT 632.100 666.600 633.900 672.600 ;
        RECT 644.700 669.600 645.900 679.950 ;
        RECT 659.100 678.150 660.900 679.950 ;
        RECT 662.700 674.700 663.900 679.950 ;
        RECT 664.950 678.150 666.750 679.950 ;
        RECT 659.700 673.800 663.900 674.700 ;
        RECT 664.950 675.450 667.050 676.050 ;
        RECT 671.550 675.450 672.450 682.950 ;
        RECT 674.550 683.550 678.450 684.450 ;
        RECT 674.550 679.050 675.450 683.550 ;
        RECT 680.100 682.050 681.900 683.850 ;
        RECT 686.700 682.050 687.900 689.400 ;
        RECT 701.100 682.050 702.900 683.850 ;
        RECT 704.700 682.050 705.600 689.400 ;
        RECT 706.950 682.050 708.750 683.850 ;
        RECT 719.250 682.050 721.050 683.850 ;
        RECT 722.400 682.050 723.300 689.400 ;
        RECT 732.000 684.450 736.050 685.050 ;
        RECT 725.100 682.050 726.900 683.850 ;
        RECT 731.550 682.950 736.050 684.450 ;
        RECT 679.950 679.950 682.050 682.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 688.950 679.950 691.050 682.050 ;
        RECT 700.950 679.950 703.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 718.950 679.950 721.050 682.050 ;
        RECT 721.950 679.950 724.050 682.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 674.550 677.550 679.050 679.050 ;
        RECT 683.100 678.150 684.900 679.950 ;
        RECT 675.000 676.950 679.050 677.550 ;
        RECT 664.950 674.550 672.450 675.450 ;
        RECT 686.700 675.600 687.900 679.950 ;
        RECT 689.100 678.150 690.900 679.950 ;
        RECT 686.700 674.700 690.300 675.600 ;
        RECT 664.950 673.950 667.050 674.550 ;
        RECT 644.100 666.600 645.900 669.600 ;
        RECT 647.100 666.000 648.900 669.600 ;
        RECT 659.700 666.600 661.500 673.800 ;
        RECT 664.800 666.000 666.600 672.600 ;
        RECT 680.100 671.700 687.900 673.050 ;
        RECT 680.100 666.600 681.900 671.700 ;
        RECT 683.100 666.000 684.900 670.800 ;
        RECT 686.100 666.600 687.900 671.700 ;
        RECT 689.100 672.600 690.300 674.700 ;
        RECT 689.100 666.600 690.900 672.600 ;
        RECT 704.700 669.600 705.600 679.950 ;
        RECT 722.400 669.600 723.300 679.950 ;
        RECT 731.550 679.050 732.450 682.950 ;
        RECT 737.400 682.050 738.300 689.400 ;
        RECT 742.950 682.050 744.750 683.850 ;
        RECT 761.250 682.050 763.050 683.850 ;
        RECT 764.400 682.050 765.300 689.400 ;
        RECT 770.550 688.500 771.450 689.400 ;
        RECT 787.950 688.800 788.850 690.900 ;
        RECT 791.850 690.600 793.650 690.900 ;
        RECT 794.550 690.600 797.550 692.400 ;
        RECT 794.550 689.700 795.750 690.600 ;
        RECT 780.450 688.500 788.850 688.800 ;
        RECT 770.550 687.900 788.850 688.500 ;
        RECT 790.950 688.800 795.750 689.700 ;
        RECT 799.650 689.400 801.450 702.000 ;
        RECT 802.650 689.400 804.450 701.400 ;
        RECT 816.000 690.600 817.800 701.400 ;
        RECT 816.000 689.400 819.600 690.600 ;
        RECT 821.100 689.400 822.900 702.000 ;
        RECT 833.100 695.400 834.900 702.000 ;
        RECT 836.100 695.400 837.900 701.400 ;
        RECT 848.100 695.400 849.900 702.000 ;
        RECT 851.100 695.400 852.900 701.400 ;
        RECT 854.100 695.400 855.900 702.000 ;
        RECT 770.550 687.300 782.250 687.900 ;
        RECT 767.100 682.050 768.900 683.850 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 731.550 677.550 736.050 679.050 ;
        RECT 732.000 676.950 736.050 677.550 ;
        RECT 737.400 672.600 738.300 679.950 ;
        RECT 739.950 678.150 741.750 679.950 ;
        RECT 746.100 678.150 747.900 679.950 ;
        RECT 737.400 671.400 742.500 672.600 ;
        RECT 701.100 666.000 702.900 669.600 ;
        RECT 704.100 666.600 705.900 669.600 ;
        RECT 707.100 666.000 708.900 669.600 ;
        RECT 719.100 666.000 720.900 669.600 ;
        RECT 722.100 666.600 723.900 669.600 ;
        RECT 725.100 666.000 726.900 669.600 ;
        RECT 737.700 666.000 739.500 669.600 ;
        RECT 740.700 666.600 742.500 671.400 ;
        RECT 745.200 666.000 747.000 672.600 ;
        RECT 751.950 672.450 754.050 673.050 ;
        RECT 760.950 672.450 763.050 673.050 ;
        RECT 751.950 671.550 763.050 672.450 ;
        RECT 751.950 670.950 754.050 671.550 ;
        RECT 760.950 670.950 763.050 671.550 ;
        RECT 764.400 669.600 765.300 679.950 ;
        RECT 770.550 672.600 771.450 687.300 ;
        RECT 780.450 687.000 782.250 687.300 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 782.100 680.400 784.200 682.050 ;
        RECT 772.950 677.400 774.750 679.950 ;
        RECT 776.100 679.200 784.200 680.400 ;
        RECT 776.100 678.600 777.900 679.200 ;
        RECT 779.100 677.400 780.900 678.000 ;
        RECT 772.950 676.200 780.900 677.400 ;
        RECT 790.950 676.200 791.850 688.800 ;
        RECT 794.550 686.100 796.650 686.700 ;
        RECT 800.550 686.100 802.350 686.550 ;
        RECT 794.550 684.900 802.350 686.100 ;
        RECT 794.550 684.600 796.650 684.900 ;
        RECT 800.550 684.750 802.350 684.900 ;
        RECT 803.250 682.050 804.450 689.400 ;
        RECT 815.100 682.050 816.900 683.850 ;
        RECT 818.700 682.050 819.600 689.400 ;
        RECT 820.950 682.050 822.750 683.850 ;
        RECT 833.100 682.050 834.900 683.850 ;
        RECT 836.100 682.050 837.300 695.400 ;
        RECT 843.000 684.450 847.050 685.050 ;
        RECT 842.550 682.950 847.050 684.450 ;
        RECT 799.950 681.750 804.450 682.050 ;
        RECT 798.150 679.950 804.450 681.750 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 820.950 679.950 823.050 682.050 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 779.850 675.000 791.850 676.200 ;
        RECT 779.850 673.200 780.900 675.000 ;
        RECT 790.050 674.400 791.850 675.000 ;
        RECT 770.550 670.800 772.950 672.600 ;
        RECT 761.100 666.000 762.900 669.600 ;
        RECT 764.100 666.600 765.900 669.600 ;
        RECT 767.100 666.000 768.900 669.600 ;
        RECT 771.150 666.600 772.950 670.800 ;
        RECT 774.150 666.000 775.950 672.600 ;
        RECT 776.850 670.200 778.950 671.700 ;
        RECT 779.850 671.400 781.650 673.200 ;
        RECT 803.250 672.600 804.450 679.950 ;
        RECT 782.850 671.550 784.650 672.300 ;
        RECT 782.850 670.500 787.800 671.550 ;
        RECT 776.850 669.600 780.750 670.200 ;
        RECT 786.750 669.600 787.800 670.500 ;
        RECT 794.250 669.600 796.650 671.700 ;
        RECT 777.150 668.700 780.750 669.600 ;
        RECT 778.950 666.600 780.750 668.700 ;
        RECT 783.450 666.000 785.250 669.600 ;
        RECT 786.750 666.600 788.550 669.600 ;
        RECT 789.750 666.000 791.550 669.600 ;
        RECT 794.250 666.600 796.050 669.600 ;
        RECT 799.350 666.000 801.150 672.600 ;
        RECT 802.650 666.600 804.450 672.600 ;
        RECT 818.700 669.600 819.600 679.950 ;
        RECT 836.100 669.600 837.300 679.950 ;
        RECT 842.550 679.050 843.450 682.950 ;
        RECT 851.700 682.050 852.900 695.400 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 850.950 679.950 853.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 838.950 677.550 843.450 679.050 ;
        RECT 848.100 678.150 849.900 679.950 ;
        RECT 838.950 676.950 843.000 677.550 ;
        RECT 851.700 674.700 852.900 679.950 ;
        RECT 853.950 678.150 855.750 679.950 ;
        RECT 848.700 673.800 852.900 674.700 ;
        RECT 815.100 666.000 816.900 669.600 ;
        RECT 818.100 666.600 819.900 669.600 ;
        RECT 821.100 666.000 822.900 669.600 ;
        RECT 833.100 666.000 834.900 669.600 ;
        RECT 836.100 666.600 837.900 669.600 ;
        RECT 848.700 666.600 850.500 673.800 ;
        RECT 853.800 666.000 855.600 672.600 ;
        RECT 11.700 655.200 13.500 662.400 ;
        RECT 16.800 656.400 18.600 663.000 ;
        RECT 29.100 659.400 30.900 662.400 ;
        RECT 32.100 659.400 33.900 663.000 ;
        RECT 11.700 654.300 15.900 655.200 ;
        RECT 11.100 649.050 12.900 650.850 ;
        RECT 14.700 649.050 15.900 654.300 ;
        RECT 16.950 649.050 18.750 650.850 ;
        RECT 29.700 649.050 30.900 659.400 ;
        RECT 44.700 655.200 46.500 662.400 ;
        RECT 49.800 656.400 51.600 663.000 ;
        RECT 62.100 659.400 63.900 663.000 ;
        RECT 65.100 659.400 66.900 662.400 ;
        RECT 68.100 659.400 69.900 663.000 ;
        RECT 44.700 654.300 48.900 655.200 ;
        RECT 34.950 651.450 39.000 652.050 ;
        RECT 34.950 649.950 39.450 651.450 ;
        RECT 10.950 646.950 13.050 649.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 28.950 646.950 31.050 649.050 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 14.700 633.600 15.900 646.950 ;
        RECT 29.700 633.600 30.900 646.950 ;
        RECT 32.100 645.150 33.900 646.950 ;
        RECT 38.550 646.050 39.450 649.950 ;
        RECT 44.100 649.050 45.900 650.850 ;
        RECT 47.700 649.050 48.900 654.300 ;
        RECT 49.950 649.050 51.750 650.850 ;
        RECT 65.700 649.050 66.600 659.400 ;
        RECT 80.100 656.400 81.900 662.400 ;
        RECT 80.700 654.300 81.900 656.400 ;
        RECT 83.100 657.300 84.900 662.400 ;
        RECT 86.100 658.200 87.900 663.000 ;
        RECT 89.100 657.300 90.900 662.400 ;
        RECT 101.100 659.400 102.900 662.400 ;
        RECT 104.100 659.400 105.900 663.000 ;
        RECT 83.100 655.950 90.900 657.300 ;
        RECT 80.700 653.400 84.300 654.300 ;
        RECT 80.100 649.050 81.900 650.850 ;
        RECT 83.100 649.050 84.300 653.400 ;
        RECT 91.950 651.450 96.000 652.050 ;
        RECT 86.100 649.050 87.900 650.850 ;
        RECT 91.950 649.950 96.450 651.450 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 46.950 646.950 49.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 67.950 646.950 70.050 649.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 88.950 646.950 91.050 649.050 ;
        RECT 38.550 644.550 43.050 646.050 ;
        RECT 39.000 643.950 43.050 644.550 ;
        RECT 47.700 633.600 48.900 646.950 ;
        RECT 62.100 645.150 63.900 646.950 ;
        RECT 65.700 639.600 66.600 646.950 ;
        RECT 67.950 645.150 69.750 646.950 ;
        RECT 83.100 639.600 84.300 646.950 ;
        RECT 89.100 645.150 90.900 646.950 ;
        RECT 95.550 646.050 96.450 649.950 ;
        RECT 101.700 649.050 102.900 659.400 ;
        RECT 107.550 656.400 109.350 662.400 ;
        RECT 110.850 656.400 112.650 663.000 ;
        RECT 115.950 659.400 117.750 662.400 ;
        RECT 120.450 659.400 122.250 663.000 ;
        RECT 123.450 659.400 125.250 662.400 ;
        RECT 126.750 659.400 128.550 663.000 ;
        RECT 131.250 660.300 133.050 662.400 ;
        RECT 131.250 659.400 134.850 660.300 ;
        RECT 115.350 657.300 117.750 659.400 ;
        RECT 124.200 658.500 125.250 659.400 ;
        RECT 131.250 658.800 135.150 659.400 ;
        RECT 124.200 657.450 129.150 658.500 ;
        RECT 127.350 656.700 129.150 657.450 ;
        RECT 107.550 649.050 108.750 656.400 ;
        RECT 130.350 655.800 132.150 657.600 ;
        RECT 133.050 657.300 135.150 658.800 ;
        RECT 136.050 656.400 137.850 663.000 ;
        RECT 139.050 658.200 140.850 662.400 ;
        RECT 139.050 656.400 141.450 658.200 ;
        RECT 152.400 656.400 154.200 663.000 ;
        RECT 120.150 654.000 121.950 654.600 ;
        RECT 131.100 654.000 132.150 655.800 ;
        RECT 120.150 652.800 132.150 654.000 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 107.550 647.250 113.850 649.050 ;
        RECT 107.550 646.950 112.050 647.250 ;
        RECT 95.550 644.550 100.050 646.050 ;
        RECT 96.000 643.950 100.050 644.550 ;
        RECT 63.000 638.400 66.600 639.600 ;
        RECT 11.100 627.000 12.900 633.600 ;
        RECT 14.100 627.600 15.900 633.600 ;
        RECT 17.100 627.000 18.900 633.600 ;
        RECT 29.100 627.600 30.900 633.600 ;
        RECT 32.100 627.000 33.900 633.600 ;
        RECT 44.100 627.000 45.900 633.600 ;
        RECT 47.100 627.600 48.900 633.600 ;
        RECT 50.100 627.000 51.900 633.600 ;
        RECT 63.000 627.600 64.800 638.400 ;
        RECT 68.100 627.000 69.900 639.600 ;
        RECT 83.100 638.100 85.500 639.600 ;
        RECT 81.000 635.100 82.800 636.900 ;
        RECT 80.700 627.000 82.500 633.600 ;
        RECT 83.700 627.600 85.500 638.100 ;
        RECT 88.800 627.000 90.600 639.600 ;
        RECT 101.700 633.600 102.900 646.950 ;
        RECT 104.100 645.150 105.900 646.950 ;
        RECT 107.550 639.600 108.750 646.950 ;
        RECT 109.650 644.100 111.450 644.250 ;
        RECT 115.350 644.100 117.450 644.400 ;
        RECT 109.650 642.900 117.450 644.100 ;
        RECT 109.650 642.450 111.450 642.900 ;
        RECT 115.350 642.300 117.450 642.900 ;
        RECT 120.150 640.200 121.050 652.800 ;
        RECT 131.100 651.600 139.050 652.800 ;
        RECT 131.100 651.000 132.900 651.600 ;
        RECT 134.100 649.800 135.900 650.400 ;
        RECT 127.800 648.600 135.900 649.800 ;
        RECT 137.250 649.050 139.050 651.600 ;
        RECT 127.800 646.950 129.900 648.600 ;
        RECT 136.950 646.950 139.050 649.050 ;
        RECT 129.750 641.700 131.550 642.000 ;
        RECT 140.550 641.700 141.450 656.400 ;
        RECT 157.500 655.200 159.300 662.400 ;
        RECT 142.950 654.450 145.050 655.050 ;
        RECT 151.950 654.450 154.050 655.050 ;
        RECT 142.950 653.550 154.050 654.450 ;
        RECT 142.950 652.950 145.050 653.550 ;
        RECT 151.950 652.950 154.050 653.550 ;
        RECT 155.100 654.300 159.300 655.200 ;
        RECT 161.550 656.400 163.350 662.400 ;
        RECT 164.850 656.400 166.650 663.000 ;
        RECT 169.950 659.400 171.750 662.400 ;
        RECT 174.450 659.400 176.250 663.000 ;
        RECT 177.450 659.400 179.250 662.400 ;
        RECT 180.750 659.400 182.550 663.000 ;
        RECT 185.250 660.300 187.050 662.400 ;
        RECT 185.250 659.400 188.850 660.300 ;
        RECT 169.350 657.300 171.750 659.400 ;
        RECT 178.200 658.500 179.250 659.400 ;
        RECT 185.250 658.800 189.150 659.400 ;
        RECT 178.200 657.450 183.150 658.500 ;
        RECT 181.350 656.700 183.150 657.450 ;
        RECT 152.250 649.050 154.050 650.850 ;
        RECT 155.100 649.050 156.300 654.300 ;
        RECT 158.100 649.050 159.900 650.850 ;
        RECT 161.550 649.050 162.750 656.400 ;
        RECT 184.350 655.800 186.150 657.600 ;
        RECT 187.050 657.300 189.150 658.800 ;
        RECT 190.050 656.400 191.850 663.000 ;
        RECT 193.050 658.200 194.850 662.400 ;
        RECT 193.050 656.400 195.450 658.200 ;
        RECT 206.100 656.400 207.900 662.400 ;
        RECT 174.150 654.000 175.950 654.600 ;
        RECT 185.100 654.000 186.150 655.800 ;
        RECT 174.150 652.800 186.150 654.000 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 154.950 646.950 157.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 161.550 647.250 167.850 649.050 ;
        RECT 161.550 646.950 166.050 647.250 ;
        RECT 129.750 641.100 141.450 641.700 ;
        RECT 101.100 627.600 102.900 633.600 ;
        RECT 104.100 627.000 105.900 633.600 ;
        RECT 107.550 627.600 109.350 639.600 ;
        RECT 110.550 627.000 112.350 639.600 ;
        RECT 116.250 639.300 121.050 640.200 ;
        RECT 123.150 640.500 141.450 641.100 ;
        RECT 123.150 640.200 131.550 640.500 ;
        RECT 116.250 638.400 117.450 639.300 ;
        RECT 114.450 636.600 117.450 638.400 ;
        RECT 118.350 638.100 120.150 638.400 ;
        RECT 123.150 638.100 124.050 640.200 ;
        RECT 140.550 639.600 141.450 640.500 ;
        RECT 118.350 637.200 124.050 638.100 ;
        RECT 124.950 638.700 126.750 639.300 ;
        RECT 124.950 637.500 132.750 638.700 ;
        RECT 118.350 636.600 120.150 637.200 ;
        RECT 130.650 636.600 132.750 637.500 ;
        RECT 115.350 633.600 117.450 635.700 ;
        RECT 121.950 635.550 123.750 636.300 ;
        RECT 126.750 635.550 128.550 636.300 ;
        RECT 121.950 634.500 128.550 635.550 ;
        RECT 115.350 627.600 117.150 633.600 ;
        RECT 119.850 627.000 121.650 633.600 ;
        RECT 122.850 627.600 124.650 634.500 ;
        RECT 125.850 627.000 127.650 633.600 ;
        RECT 130.650 627.600 132.450 636.600 ;
        RECT 136.050 627.000 137.850 639.600 ;
        RECT 139.050 637.800 141.450 639.600 ;
        RECT 139.050 627.600 140.850 637.800 ;
        RECT 155.100 633.600 156.300 646.950 ;
        RECT 161.550 639.600 162.750 646.950 ;
        RECT 163.650 644.100 165.450 644.250 ;
        RECT 169.350 644.100 171.450 644.400 ;
        RECT 163.650 642.900 171.450 644.100 ;
        RECT 163.650 642.450 165.450 642.900 ;
        RECT 169.350 642.300 171.450 642.900 ;
        RECT 174.150 640.200 175.050 652.800 ;
        RECT 185.100 651.600 193.050 652.800 ;
        RECT 185.100 651.000 186.900 651.600 ;
        RECT 188.100 649.800 189.900 650.400 ;
        RECT 181.800 648.600 189.900 649.800 ;
        RECT 191.250 649.050 193.050 651.600 ;
        RECT 181.800 646.950 183.900 648.600 ;
        RECT 190.950 646.950 193.050 649.050 ;
        RECT 183.750 641.700 185.550 642.000 ;
        RECT 194.550 641.700 195.450 656.400 ;
        RECT 206.700 654.300 207.900 656.400 ;
        RECT 209.100 657.300 210.900 662.400 ;
        RECT 212.100 658.200 213.900 663.000 ;
        RECT 215.100 657.300 216.900 662.400 ;
        RECT 209.100 655.950 216.900 657.300 ;
        RECT 227.100 656.400 228.900 662.400 ;
        RECT 230.100 656.400 231.900 663.000 ;
        RECT 233.100 659.400 234.900 662.400 ;
        RECT 206.700 653.400 210.300 654.300 ;
        RECT 206.100 649.050 207.900 650.850 ;
        RECT 209.100 649.050 210.300 653.400 ;
        RECT 212.100 649.050 213.900 650.850 ;
        RECT 227.100 649.050 228.300 656.400 ;
        RECT 233.700 655.500 234.900 659.400 ;
        RECT 245.100 656.400 246.900 663.000 ;
        RECT 248.100 655.500 249.900 662.400 ;
        RECT 251.100 656.400 252.900 663.000 ;
        RECT 254.100 655.500 255.900 662.400 ;
        RECT 257.100 656.400 258.900 663.000 ;
        RECT 260.100 655.500 261.900 662.400 ;
        RECT 263.100 656.400 264.900 663.000 ;
        RECT 266.100 655.500 267.900 662.400 ;
        RECT 269.100 656.400 270.900 663.000 ;
        RECT 282.000 656.400 283.800 663.000 ;
        RECT 286.500 657.600 288.300 662.400 ;
        RECT 289.500 659.400 291.300 663.000 ;
        RECT 302.100 659.400 303.900 663.000 ;
        RECT 305.100 659.400 306.900 662.400 ;
        RECT 286.500 656.400 291.600 657.600 ;
        RECT 229.200 654.600 234.900 655.500 ;
        RECT 229.200 653.700 231.000 654.600 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 208.950 646.950 211.050 649.050 ;
        RECT 211.950 646.950 214.050 649.050 ;
        RECT 214.950 646.950 217.050 649.050 ;
        RECT 227.100 646.950 229.200 649.050 ;
        RECT 183.750 641.100 195.450 641.700 ;
        RECT 152.100 627.000 153.900 633.600 ;
        RECT 155.100 627.600 156.900 633.600 ;
        RECT 158.100 627.000 159.900 633.600 ;
        RECT 161.550 627.600 163.350 639.600 ;
        RECT 164.550 627.000 166.350 639.600 ;
        RECT 170.250 639.300 175.050 640.200 ;
        RECT 177.150 640.500 195.450 641.100 ;
        RECT 196.950 642.450 199.050 643.050 ;
        RECT 205.950 642.450 208.050 643.050 ;
        RECT 196.950 641.550 208.050 642.450 ;
        RECT 196.950 640.950 199.050 641.550 ;
        RECT 205.950 640.950 208.050 641.550 ;
        RECT 177.150 640.200 185.550 640.500 ;
        RECT 170.250 638.400 171.450 639.300 ;
        RECT 168.450 636.600 171.450 638.400 ;
        RECT 172.350 638.100 174.150 638.400 ;
        RECT 177.150 638.100 178.050 640.200 ;
        RECT 194.550 639.600 195.450 640.500 ;
        RECT 172.350 637.200 178.050 638.100 ;
        RECT 178.950 638.700 180.750 639.300 ;
        RECT 178.950 637.500 186.750 638.700 ;
        RECT 172.350 636.600 174.150 637.200 ;
        RECT 184.650 636.600 186.750 637.500 ;
        RECT 169.350 633.600 171.450 635.700 ;
        RECT 175.950 635.550 177.750 636.300 ;
        RECT 180.750 635.550 182.550 636.300 ;
        RECT 175.950 634.500 182.550 635.550 ;
        RECT 169.350 627.600 171.150 633.600 ;
        RECT 173.850 627.000 175.650 633.600 ;
        RECT 176.850 627.600 178.650 634.500 ;
        RECT 179.850 627.000 181.650 633.600 ;
        RECT 184.650 627.600 186.450 636.600 ;
        RECT 190.050 627.000 191.850 639.600 ;
        RECT 193.050 637.800 195.450 639.600 ;
        RECT 209.100 639.600 210.300 646.950 ;
        RECT 215.100 645.150 216.900 646.950 ;
        RECT 227.100 639.600 228.300 646.950 ;
        RECT 230.100 642.300 231.000 653.700 ;
        RECT 247.050 654.300 249.900 655.500 ;
        RECT 252.000 654.300 255.900 655.500 ;
        RECT 258.000 654.300 261.900 655.500 ;
        RECT 264.000 654.300 267.900 655.500 ;
        RECT 247.050 649.050 248.100 654.300 ;
        RECT 252.000 653.400 253.200 654.300 ;
        RECT 258.000 653.400 259.200 654.300 ;
        RECT 264.000 653.400 265.200 654.300 ;
        RECT 249.000 652.200 253.200 653.400 ;
        RECT 249.000 651.600 250.800 652.200 ;
        RECT 232.500 646.950 234.600 649.050 ;
        RECT 232.800 645.150 234.600 646.950 ;
        RECT 247.050 646.950 250.200 649.050 ;
        RECT 229.200 641.400 231.000 642.300 ;
        RECT 247.050 641.700 248.100 646.950 ;
        RECT 252.000 641.700 253.200 652.200 ;
        RECT 255.000 652.200 259.200 653.400 ;
        RECT 255.000 651.600 256.800 652.200 ;
        RECT 258.000 641.700 259.200 652.200 ;
        RECT 261.000 652.200 265.200 653.400 ;
        RECT 261.000 651.600 262.800 652.200 ;
        RECT 264.000 641.700 265.200 652.200 ;
        RECT 266.400 649.050 268.200 650.850 ;
        RECT 281.100 649.050 282.900 650.850 ;
        RECT 287.250 649.050 289.050 650.850 ;
        RECT 290.700 649.050 291.600 656.400 ;
        RECT 305.100 649.050 306.300 659.400 ;
        RECT 308.550 656.400 310.350 662.400 ;
        RECT 311.850 656.400 313.650 663.000 ;
        RECT 316.950 659.400 318.750 662.400 ;
        RECT 321.450 659.400 323.250 663.000 ;
        RECT 324.450 659.400 326.250 662.400 ;
        RECT 327.750 659.400 329.550 663.000 ;
        RECT 332.250 660.300 334.050 662.400 ;
        RECT 332.250 659.400 335.850 660.300 ;
        RECT 316.350 657.300 318.750 659.400 ;
        RECT 325.200 658.500 326.250 659.400 ;
        RECT 332.250 658.800 336.150 659.400 ;
        RECT 325.200 657.450 330.150 658.500 ;
        RECT 328.350 656.700 330.150 657.450 ;
        RECT 308.550 649.050 309.750 656.400 ;
        RECT 331.350 655.800 333.150 657.600 ;
        RECT 334.050 657.300 336.150 658.800 ;
        RECT 337.050 656.400 338.850 663.000 ;
        RECT 340.050 658.200 341.850 662.400 ;
        RECT 340.050 656.400 342.450 658.200 ;
        RECT 356.100 656.400 357.900 662.400 ;
        RECT 321.150 654.000 322.950 654.600 ;
        RECT 332.100 654.000 333.150 655.800 ;
        RECT 321.150 652.800 333.150 654.000 ;
        RECT 266.100 646.950 268.200 649.050 ;
        RECT 280.950 646.950 283.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 301.950 646.950 304.050 649.050 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 308.550 647.250 314.850 649.050 ;
        RECT 308.550 646.950 313.050 647.250 ;
        RECT 284.250 645.150 286.050 646.950 ;
        RECT 271.950 642.450 274.050 643.050 ;
        RECT 286.950 642.450 289.050 643.050 ;
        RECT 229.200 640.500 234.900 641.400 ;
        RECT 247.050 640.500 249.900 641.700 ;
        RECT 252.000 640.500 255.900 641.700 ;
        RECT 258.000 640.500 261.900 641.700 ;
        RECT 264.000 640.500 267.900 641.700 ;
        RECT 271.950 641.550 289.050 642.450 ;
        RECT 271.950 640.950 274.050 641.550 ;
        RECT 286.950 640.950 289.050 641.550 ;
        RECT 209.100 638.100 211.500 639.600 ;
        RECT 193.050 627.600 194.850 637.800 ;
        RECT 207.000 635.100 208.800 636.900 ;
        RECT 206.700 627.000 208.500 633.600 ;
        RECT 209.700 627.600 211.500 638.100 ;
        RECT 214.800 627.000 216.600 639.600 ;
        RECT 227.100 627.600 228.900 639.600 ;
        RECT 230.100 627.000 231.900 637.800 ;
        RECT 233.700 633.600 234.900 640.500 ;
        RECT 233.100 627.600 234.900 633.600 ;
        RECT 245.100 627.000 246.900 639.600 ;
        RECT 248.100 627.600 249.900 640.500 ;
        RECT 251.100 627.000 252.900 639.600 ;
        RECT 254.100 627.600 255.900 640.500 ;
        RECT 257.100 627.000 258.900 639.600 ;
        RECT 260.100 627.600 261.900 640.500 ;
        RECT 263.100 627.000 264.900 639.600 ;
        RECT 266.100 627.600 267.900 640.500 ;
        RECT 290.700 639.600 291.600 646.950 ;
        RECT 302.100 645.150 303.900 646.950 ;
        RECT 269.100 627.000 270.900 639.600 ;
        RECT 281.100 638.700 288.900 639.600 ;
        RECT 281.100 627.600 282.900 638.700 ;
        RECT 284.100 627.000 285.900 637.800 ;
        RECT 287.100 627.600 288.900 638.700 ;
        RECT 290.100 627.600 291.900 639.600 ;
        RECT 305.100 633.600 306.300 646.950 ;
        RECT 308.550 639.600 309.750 646.950 ;
        RECT 310.650 644.100 312.450 644.250 ;
        RECT 316.350 644.100 318.450 644.400 ;
        RECT 310.650 642.900 318.450 644.100 ;
        RECT 310.650 642.450 312.450 642.900 ;
        RECT 316.350 642.300 318.450 642.900 ;
        RECT 321.150 640.200 322.050 652.800 ;
        RECT 332.100 651.600 340.050 652.800 ;
        RECT 332.100 651.000 333.900 651.600 ;
        RECT 335.100 649.800 336.900 650.400 ;
        RECT 328.800 648.600 336.900 649.800 ;
        RECT 338.250 649.050 340.050 651.600 ;
        RECT 328.800 646.950 330.900 648.600 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 330.750 641.700 332.550 642.000 ;
        RECT 341.550 641.700 342.450 656.400 ;
        RECT 356.700 654.300 357.900 656.400 ;
        RECT 359.100 657.300 360.900 662.400 ;
        RECT 362.100 658.200 363.900 663.000 ;
        RECT 365.100 657.300 366.900 662.400 ;
        RECT 359.100 655.950 366.900 657.300 ;
        RECT 377.400 656.400 379.200 663.000 ;
        RECT 382.500 655.200 384.300 662.400 ;
        RECT 395.100 656.400 396.900 662.400 ;
        RECT 380.100 654.300 384.300 655.200 ;
        RECT 395.700 654.300 396.900 656.400 ;
        RECT 398.100 657.300 399.900 662.400 ;
        RECT 401.100 658.200 402.900 663.000 ;
        RECT 404.100 657.300 405.900 662.400 ;
        RECT 419.100 659.400 420.900 663.000 ;
        RECT 422.100 659.400 423.900 662.400 ;
        RECT 425.100 659.400 426.900 663.000 ;
        RECT 398.100 655.950 405.900 657.300 ;
        RECT 356.700 653.400 360.300 654.300 ;
        RECT 356.100 649.050 357.900 650.850 ;
        RECT 359.100 649.050 360.300 653.400 ;
        RECT 362.100 649.050 363.900 650.850 ;
        RECT 377.250 649.050 379.050 650.850 ;
        RECT 380.100 649.050 381.300 654.300 ;
        RECT 395.700 653.400 399.300 654.300 ;
        RECT 383.100 649.050 384.900 650.850 ;
        RECT 395.100 649.050 396.900 650.850 ;
        RECT 398.100 649.050 399.300 653.400 ;
        RECT 401.100 649.050 402.900 650.850 ;
        RECT 422.400 649.050 423.300 659.400 ;
        RECT 429.150 658.200 430.950 662.400 ;
        RECT 428.550 656.400 430.950 658.200 ;
        RECT 432.150 656.400 433.950 663.000 ;
        RECT 436.950 660.300 438.750 662.400 ;
        RECT 435.150 659.400 438.750 660.300 ;
        RECT 441.450 659.400 443.250 663.000 ;
        RECT 444.750 659.400 446.550 662.400 ;
        RECT 447.750 659.400 449.550 663.000 ;
        RECT 452.250 659.400 454.050 662.400 ;
        RECT 434.850 658.800 438.750 659.400 ;
        RECT 434.850 657.300 436.950 658.800 ;
        RECT 444.750 658.500 445.800 659.400 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 376.950 646.950 379.050 649.050 ;
        RECT 379.950 646.950 382.050 649.050 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 394.950 646.950 397.050 649.050 ;
        RECT 397.950 646.950 400.050 649.050 ;
        RECT 400.950 646.950 403.050 649.050 ;
        RECT 403.950 646.950 406.050 649.050 ;
        RECT 418.950 646.950 421.050 649.050 ;
        RECT 421.950 646.950 424.050 649.050 ;
        RECT 424.950 646.950 427.050 649.050 ;
        RECT 330.750 641.100 342.450 641.700 ;
        RECT 302.100 627.000 303.900 633.600 ;
        RECT 305.100 627.600 306.900 633.600 ;
        RECT 308.550 627.600 310.350 639.600 ;
        RECT 311.550 627.000 313.350 639.600 ;
        RECT 317.250 639.300 322.050 640.200 ;
        RECT 324.150 640.500 342.450 641.100 ;
        RECT 324.150 640.200 332.550 640.500 ;
        RECT 317.250 638.400 318.450 639.300 ;
        RECT 315.450 636.600 318.450 638.400 ;
        RECT 319.350 638.100 321.150 638.400 ;
        RECT 324.150 638.100 325.050 640.200 ;
        RECT 341.550 639.600 342.450 640.500 ;
        RECT 319.350 637.200 325.050 638.100 ;
        RECT 325.950 638.700 327.750 639.300 ;
        RECT 325.950 637.500 333.750 638.700 ;
        RECT 319.350 636.600 321.150 637.200 ;
        RECT 331.650 636.600 333.750 637.500 ;
        RECT 316.350 633.600 318.450 635.700 ;
        RECT 322.950 635.550 324.750 636.300 ;
        RECT 327.750 635.550 329.550 636.300 ;
        RECT 322.950 634.500 329.550 635.550 ;
        RECT 316.350 627.600 318.150 633.600 ;
        RECT 320.850 627.000 322.650 633.600 ;
        RECT 323.850 627.600 325.650 634.500 ;
        RECT 326.850 627.000 328.650 633.600 ;
        RECT 331.650 627.600 333.450 636.600 ;
        RECT 337.050 627.000 338.850 639.600 ;
        RECT 340.050 637.800 342.450 639.600 ;
        RECT 359.100 639.600 360.300 646.950 ;
        RECT 365.100 645.150 366.900 646.950 ;
        RECT 359.100 638.100 361.500 639.600 ;
        RECT 340.050 627.600 341.850 637.800 ;
        RECT 357.000 635.100 358.800 636.900 ;
        RECT 356.700 627.000 358.500 633.600 ;
        RECT 359.700 627.600 361.500 638.100 ;
        RECT 364.800 627.000 366.600 639.600 ;
        RECT 380.100 633.600 381.300 646.950 ;
        RECT 398.100 639.600 399.300 646.950 ;
        RECT 404.100 645.150 405.900 646.950 ;
        RECT 419.250 645.150 421.050 646.950 ;
        RECT 422.400 639.600 423.300 646.950 ;
        RECT 425.100 645.150 426.900 646.950 ;
        RECT 428.550 641.700 429.450 656.400 ;
        RECT 437.850 655.800 439.650 657.600 ;
        RECT 440.850 657.450 445.800 658.500 ;
        RECT 440.850 656.700 442.650 657.450 ;
        RECT 452.250 657.300 454.650 659.400 ;
        RECT 457.350 656.400 459.150 663.000 ;
        RECT 460.650 656.400 462.450 662.400 ;
        RECT 473.400 656.400 475.200 663.000 ;
        RECT 437.850 654.000 438.900 655.800 ;
        RECT 448.050 654.000 449.850 654.600 ;
        RECT 437.850 652.800 449.850 654.000 ;
        RECT 430.950 651.600 438.900 652.800 ;
        RECT 430.950 649.050 432.750 651.600 ;
        RECT 437.100 651.000 438.900 651.600 ;
        RECT 434.100 649.800 435.900 650.400 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 434.100 648.600 442.200 649.800 ;
        RECT 440.100 646.950 442.200 648.600 ;
        RECT 438.450 641.700 440.250 642.000 ;
        RECT 428.550 641.100 440.250 641.700 ;
        RECT 428.550 640.500 446.850 641.100 ;
        RECT 428.550 639.600 429.450 640.500 ;
        RECT 438.450 640.200 446.850 640.500 ;
        RECT 398.100 638.100 400.500 639.600 ;
        RECT 396.000 635.100 397.800 636.900 ;
        RECT 377.100 627.000 378.900 633.600 ;
        RECT 380.100 627.600 381.900 633.600 ;
        RECT 383.100 627.000 384.900 633.600 ;
        RECT 395.700 627.000 397.500 633.600 ;
        RECT 398.700 627.600 400.500 638.100 ;
        RECT 403.800 627.000 405.600 639.600 ;
        RECT 419.100 627.000 420.900 639.600 ;
        RECT 422.400 638.400 426.000 639.600 ;
        RECT 424.200 627.600 426.000 638.400 ;
        RECT 428.550 637.800 430.950 639.600 ;
        RECT 429.150 627.600 430.950 637.800 ;
        RECT 432.150 627.000 433.950 639.600 ;
        RECT 443.250 638.700 445.050 639.300 ;
        RECT 437.250 637.500 445.050 638.700 ;
        RECT 445.950 638.100 446.850 640.200 ;
        RECT 448.950 640.200 449.850 652.800 ;
        RECT 461.250 649.050 462.450 656.400 ;
        RECT 478.500 655.200 480.300 662.400 ;
        RECT 492.000 656.400 493.800 663.000 ;
        RECT 496.500 657.600 498.300 662.400 ;
        RECT 499.500 659.400 501.300 663.000 ;
        RECT 504.150 658.200 505.950 662.400 ;
        RECT 496.500 656.400 501.600 657.600 ;
        RECT 476.100 654.300 480.300 655.200 ;
        RECT 473.250 649.050 475.050 650.850 ;
        RECT 476.100 649.050 477.300 654.300 ;
        RECT 479.100 649.050 480.900 650.850 ;
        RECT 491.100 649.050 492.900 650.850 ;
        RECT 497.250 649.050 499.050 650.850 ;
        RECT 500.700 649.050 501.600 656.400 ;
        RECT 503.550 656.400 505.950 658.200 ;
        RECT 507.150 656.400 508.950 663.000 ;
        RECT 511.950 660.300 513.750 662.400 ;
        RECT 510.150 659.400 513.750 660.300 ;
        RECT 516.450 659.400 518.250 663.000 ;
        RECT 519.750 659.400 521.550 662.400 ;
        RECT 522.750 659.400 524.550 663.000 ;
        RECT 527.250 659.400 529.050 662.400 ;
        RECT 509.850 658.800 513.750 659.400 ;
        RECT 509.850 657.300 511.950 658.800 ;
        RECT 519.750 658.500 520.800 659.400 ;
        RECT 456.150 647.250 462.450 649.050 ;
        RECT 457.950 646.950 462.450 647.250 ;
        RECT 472.950 646.950 475.050 649.050 ;
        RECT 475.950 646.950 478.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 490.950 646.950 493.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 496.950 646.950 499.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 452.550 644.100 454.650 644.400 ;
        RECT 458.550 644.100 460.350 644.250 ;
        RECT 452.550 642.900 460.350 644.100 ;
        RECT 452.550 642.300 454.650 642.900 ;
        RECT 458.550 642.450 460.350 642.900 ;
        RECT 448.950 639.300 453.750 640.200 ;
        RECT 461.250 639.600 462.450 646.950 ;
        RECT 466.950 642.450 469.050 643.050 ;
        RECT 472.950 642.450 475.050 643.050 ;
        RECT 466.950 641.550 475.050 642.450 ;
        RECT 466.950 640.950 469.050 641.550 ;
        RECT 472.950 640.950 475.050 641.550 ;
        RECT 452.550 638.400 453.750 639.300 ;
        RECT 449.850 638.100 451.650 638.400 ;
        RECT 437.250 636.600 439.350 637.500 ;
        RECT 445.950 637.200 451.650 638.100 ;
        RECT 449.850 636.600 451.650 637.200 ;
        RECT 452.550 636.600 455.550 638.400 ;
        RECT 437.550 627.600 439.350 636.600 ;
        RECT 441.450 635.550 443.250 636.300 ;
        RECT 446.250 635.550 448.050 636.300 ;
        RECT 441.450 634.500 448.050 635.550 ;
        RECT 442.350 627.000 444.150 633.600 ;
        RECT 445.350 627.600 447.150 634.500 ;
        RECT 452.550 633.600 454.650 635.700 ;
        RECT 448.350 627.000 450.150 633.600 ;
        RECT 452.850 627.600 454.650 633.600 ;
        RECT 457.650 627.000 459.450 639.600 ;
        RECT 460.650 627.600 462.450 639.600 ;
        RECT 476.100 633.600 477.300 646.950 ;
        RECT 494.250 645.150 496.050 646.950 ;
        RECT 500.700 639.600 501.600 646.950 ;
        RECT 503.550 641.700 504.450 656.400 ;
        RECT 512.850 655.800 514.650 657.600 ;
        RECT 515.850 657.450 520.800 658.500 ;
        RECT 515.850 656.700 517.650 657.450 ;
        RECT 527.250 657.300 529.650 659.400 ;
        RECT 532.350 656.400 534.150 663.000 ;
        RECT 535.650 656.400 537.450 662.400 ;
        RECT 548.100 659.400 549.900 663.000 ;
        RECT 551.100 659.400 552.900 662.400 ;
        RECT 554.100 659.400 555.900 663.000 ;
        RECT 512.850 654.000 513.900 655.800 ;
        RECT 523.050 654.000 524.850 654.600 ;
        RECT 512.850 652.800 524.850 654.000 ;
        RECT 505.950 651.600 513.900 652.800 ;
        RECT 505.950 649.050 507.750 651.600 ;
        RECT 512.100 651.000 513.900 651.600 ;
        RECT 509.100 649.800 510.900 650.400 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 509.100 648.600 517.200 649.800 ;
        RECT 515.100 646.950 517.200 648.600 ;
        RECT 513.450 641.700 515.250 642.000 ;
        RECT 503.550 641.100 515.250 641.700 ;
        RECT 503.550 640.500 521.850 641.100 ;
        RECT 503.550 639.600 504.450 640.500 ;
        RECT 513.450 640.200 521.850 640.500 ;
        RECT 491.100 638.700 498.900 639.600 ;
        RECT 473.100 627.000 474.900 633.600 ;
        RECT 476.100 627.600 477.900 633.600 ;
        RECT 479.100 627.000 480.900 633.600 ;
        RECT 491.100 627.600 492.900 638.700 ;
        RECT 494.100 627.000 495.900 637.800 ;
        RECT 497.100 627.600 498.900 638.700 ;
        RECT 500.100 627.600 501.900 639.600 ;
        RECT 503.550 637.800 505.950 639.600 ;
        RECT 504.150 627.600 505.950 637.800 ;
        RECT 507.150 627.000 508.950 639.600 ;
        RECT 518.250 638.700 520.050 639.300 ;
        RECT 512.250 637.500 520.050 638.700 ;
        RECT 520.950 638.100 521.850 640.200 ;
        RECT 523.950 640.200 524.850 652.800 ;
        RECT 536.250 649.050 537.450 656.400 ;
        RECT 551.700 649.050 552.600 659.400 ;
        RECT 566.100 657.300 567.900 662.400 ;
        RECT 569.100 658.200 570.900 663.000 ;
        RECT 572.100 657.300 573.900 662.400 ;
        RECT 566.100 655.950 573.900 657.300 ;
        RECT 575.100 656.400 576.900 662.400 ;
        RECT 587.100 657.300 588.900 662.400 ;
        RECT 590.100 658.200 591.900 663.000 ;
        RECT 593.100 657.300 594.900 662.400 ;
        RECT 575.100 654.300 576.300 656.400 ;
        RECT 587.100 655.950 594.900 657.300 ;
        RECT 596.100 656.400 597.900 662.400 ;
        RECT 596.100 654.300 597.300 656.400 ;
        RECT 608.700 655.200 610.500 662.400 ;
        RECT 613.800 656.400 615.600 663.000 ;
        RECT 617.550 656.400 619.350 662.400 ;
        RECT 620.850 656.400 622.650 663.000 ;
        RECT 625.950 659.400 627.750 662.400 ;
        RECT 630.450 659.400 632.250 663.000 ;
        RECT 633.450 659.400 635.250 662.400 ;
        RECT 636.750 659.400 638.550 663.000 ;
        RECT 641.250 660.300 643.050 662.400 ;
        RECT 641.250 659.400 644.850 660.300 ;
        RECT 625.350 657.300 627.750 659.400 ;
        RECT 634.200 658.500 635.250 659.400 ;
        RECT 641.250 658.800 645.150 659.400 ;
        RECT 634.200 657.450 639.150 658.500 ;
        RECT 637.350 656.700 639.150 657.450 ;
        RECT 608.700 654.300 612.900 655.200 ;
        RECT 572.700 653.400 576.300 654.300 ;
        RECT 593.700 653.400 597.300 654.300 ;
        RECT 569.100 649.050 570.900 650.850 ;
        RECT 572.700 649.050 573.900 653.400 ;
        RECT 575.100 649.050 576.900 650.850 ;
        RECT 590.100 649.050 591.900 650.850 ;
        RECT 593.700 649.050 594.900 653.400 ;
        RECT 603.000 651.450 607.050 652.050 ;
        RECT 596.100 649.050 597.900 650.850 ;
        RECT 602.550 649.950 607.050 651.450 ;
        RECT 531.150 647.250 537.450 649.050 ;
        RECT 532.950 646.950 537.450 647.250 ;
        RECT 547.950 646.950 550.050 649.050 ;
        RECT 550.950 646.950 553.050 649.050 ;
        RECT 553.950 646.950 556.050 649.050 ;
        RECT 565.950 646.950 568.050 649.050 ;
        RECT 568.950 646.950 571.050 649.050 ;
        RECT 571.950 646.950 574.050 649.050 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 589.950 646.950 592.050 649.050 ;
        RECT 592.950 646.950 595.050 649.050 ;
        RECT 595.950 646.950 598.050 649.050 ;
        RECT 527.550 644.100 529.650 644.400 ;
        RECT 533.550 644.100 535.350 644.250 ;
        RECT 527.550 642.900 535.350 644.100 ;
        RECT 527.550 642.300 529.650 642.900 ;
        RECT 533.550 642.450 535.350 642.900 ;
        RECT 523.950 639.300 528.750 640.200 ;
        RECT 536.250 639.600 537.450 646.950 ;
        RECT 548.100 645.150 549.900 646.950 ;
        RECT 551.700 639.600 552.600 646.950 ;
        RECT 553.950 645.150 555.750 646.950 ;
        RECT 566.100 645.150 567.900 646.950 ;
        RECT 572.700 639.600 573.900 646.950 ;
        RECT 587.100 645.150 588.900 646.950 ;
        RECT 593.700 639.600 594.900 646.950 ;
        RECT 602.550 646.050 603.450 649.950 ;
        RECT 608.100 649.050 609.900 650.850 ;
        RECT 611.700 649.050 612.900 654.300 ;
        RECT 613.950 649.050 615.750 650.850 ;
        RECT 617.550 649.050 618.750 656.400 ;
        RECT 640.350 655.800 642.150 657.600 ;
        RECT 643.050 657.300 645.150 658.800 ;
        RECT 646.050 656.400 647.850 663.000 ;
        RECT 649.050 658.200 650.850 662.400 ;
        RECT 649.050 656.400 651.450 658.200 ;
        RECT 630.150 654.000 631.950 654.600 ;
        RECT 641.100 654.000 642.150 655.800 ;
        RECT 630.150 652.800 642.150 654.000 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 610.950 646.950 613.050 649.050 ;
        RECT 613.950 646.950 616.050 649.050 ;
        RECT 617.550 647.250 623.850 649.050 ;
        RECT 617.550 646.950 622.050 647.250 ;
        RECT 598.950 644.550 603.450 646.050 ;
        RECT 598.950 643.950 603.000 644.550 ;
        RECT 527.550 638.400 528.750 639.300 ;
        RECT 524.850 638.100 526.650 638.400 ;
        RECT 512.250 636.600 514.350 637.500 ;
        RECT 520.950 637.200 526.650 638.100 ;
        RECT 524.850 636.600 526.650 637.200 ;
        RECT 527.550 636.600 530.550 638.400 ;
        RECT 512.550 627.600 514.350 636.600 ;
        RECT 516.450 635.550 518.250 636.300 ;
        RECT 521.250 635.550 523.050 636.300 ;
        RECT 516.450 634.500 523.050 635.550 ;
        RECT 517.350 627.000 519.150 633.600 ;
        RECT 520.350 627.600 522.150 634.500 ;
        RECT 527.550 633.600 529.650 635.700 ;
        RECT 523.350 627.000 525.150 633.600 ;
        RECT 527.850 627.600 529.650 633.600 ;
        RECT 532.650 627.000 534.450 639.600 ;
        RECT 535.650 627.600 537.450 639.600 ;
        RECT 549.000 638.400 552.600 639.600 ;
        RECT 549.000 627.600 550.800 638.400 ;
        RECT 554.100 627.000 555.900 639.600 ;
        RECT 566.400 627.000 568.200 639.600 ;
        RECT 571.500 638.100 573.900 639.600 ;
        RECT 571.500 627.600 573.300 638.100 ;
        RECT 574.200 635.100 576.000 636.900 ;
        RECT 574.500 627.000 576.300 633.600 ;
        RECT 587.400 627.000 589.200 639.600 ;
        RECT 592.500 638.100 594.900 639.600 ;
        RECT 595.950 639.450 598.050 640.050 ;
        RECT 607.950 639.450 610.050 639.900 ;
        RECT 595.950 638.550 610.050 639.450 ;
        RECT 592.500 627.600 594.300 638.100 ;
        RECT 595.950 637.950 598.050 638.550 ;
        RECT 607.950 637.800 610.050 638.550 ;
        RECT 595.200 635.100 597.000 636.900 ;
        RECT 611.700 633.600 612.900 646.950 ;
        RECT 617.550 639.600 618.750 646.950 ;
        RECT 619.650 644.100 621.450 644.250 ;
        RECT 625.350 644.100 627.450 644.400 ;
        RECT 619.650 642.900 627.450 644.100 ;
        RECT 619.650 642.450 621.450 642.900 ;
        RECT 625.350 642.300 627.450 642.900 ;
        RECT 630.150 640.200 631.050 652.800 ;
        RECT 641.100 651.600 649.050 652.800 ;
        RECT 641.100 651.000 642.900 651.600 ;
        RECT 644.100 649.800 645.900 650.400 ;
        RECT 637.800 648.600 645.900 649.800 ;
        RECT 647.250 649.050 649.050 651.600 ;
        RECT 637.800 646.950 639.900 648.600 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 639.750 641.700 641.550 642.000 ;
        RECT 650.550 641.700 651.450 656.400 ;
        RECT 662.700 655.200 664.500 662.400 ;
        RECT 667.800 656.400 669.600 663.000 ;
        RECT 672.150 658.200 673.950 662.400 ;
        RECT 671.550 656.400 673.950 658.200 ;
        RECT 675.150 656.400 676.950 663.000 ;
        RECT 679.950 660.300 681.750 662.400 ;
        RECT 678.150 659.400 681.750 660.300 ;
        RECT 684.450 659.400 686.250 663.000 ;
        RECT 687.750 659.400 689.550 662.400 ;
        RECT 690.750 659.400 692.550 663.000 ;
        RECT 695.250 659.400 697.050 662.400 ;
        RECT 677.850 658.800 681.750 659.400 ;
        RECT 677.850 657.300 679.950 658.800 ;
        RECT 687.750 658.500 688.800 659.400 ;
        RECT 662.700 654.300 666.900 655.200 ;
        RECT 662.100 649.050 663.900 650.850 ;
        RECT 665.700 649.050 666.900 654.300 ;
        RECT 667.950 649.050 669.750 650.850 ;
        RECT 661.950 646.950 664.050 649.050 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 639.750 641.100 651.450 641.700 ;
        RECT 595.500 627.000 597.300 633.600 ;
        RECT 608.100 627.000 609.900 633.600 ;
        RECT 611.100 627.600 612.900 633.600 ;
        RECT 614.100 627.000 615.900 633.600 ;
        RECT 617.550 627.600 619.350 639.600 ;
        RECT 620.550 627.000 622.350 639.600 ;
        RECT 626.250 639.300 631.050 640.200 ;
        RECT 633.150 640.500 651.450 641.100 ;
        RECT 633.150 640.200 641.550 640.500 ;
        RECT 626.250 638.400 627.450 639.300 ;
        RECT 624.450 636.600 627.450 638.400 ;
        RECT 628.350 638.100 630.150 638.400 ;
        RECT 633.150 638.100 634.050 640.200 ;
        RECT 650.550 639.600 651.450 640.500 ;
        RECT 628.350 637.200 634.050 638.100 ;
        RECT 634.950 638.700 636.750 639.300 ;
        RECT 634.950 637.500 642.750 638.700 ;
        RECT 628.350 636.600 630.150 637.200 ;
        RECT 640.650 636.600 642.750 637.500 ;
        RECT 625.350 633.600 627.450 635.700 ;
        RECT 631.950 635.550 633.750 636.300 ;
        RECT 636.750 635.550 638.550 636.300 ;
        RECT 631.950 634.500 638.550 635.550 ;
        RECT 625.350 627.600 627.150 633.600 ;
        RECT 629.850 627.000 631.650 633.600 ;
        RECT 632.850 627.600 634.650 634.500 ;
        RECT 635.850 627.000 637.650 633.600 ;
        RECT 640.650 627.600 642.450 636.600 ;
        RECT 646.050 627.000 647.850 639.600 ;
        RECT 649.050 637.800 651.450 639.600 ;
        RECT 649.050 627.600 650.850 637.800 ;
        RECT 665.700 633.600 666.900 646.950 ;
        RECT 671.550 641.700 672.450 656.400 ;
        RECT 680.850 655.800 682.650 657.600 ;
        RECT 683.850 657.450 688.800 658.500 ;
        RECT 683.850 656.700 685.650 657.450 ;
        RECT 695.250 657.300 697.650 659.400 ;
        RECT 700.350 656.400 702.150 663.000 ;
        RECT 703.650 656.400 705.450 662.400 ;
        RECT 716.100 659.400 717.900 662.400 ;
        RECT 719.100 659.400 720.900 663.000 ;
        RECT 731.100 659.400 732.900 663.000 ;
        RECT 734.100 659.400 735.900 662.400 ;
        RECT 737.100 659.400 738.900 663.000 ;
        RECT 752.100 659.400 753.900 662.400 ;
        RECT 755.100 659.400 756.900 663.000 ;
        RECT 680.850 654.000 681.900 655.800 ;
        RECT 691.050 654.000 692.850 654.600 ;
        RECT 680.850 652.800 692.850 654.000 ;
        RECT 673.950 651.600 681.900 652.800 ;
        RECT 673.950 649.050 675.750 651.600 ;
        RECT 680.100 651.000 681.900 651.600 ;
        RECT 677.100 649.800 678.900 650.400 ;
        RECT 673.950 646.950 676.050 649.050 ;
        RECT 677.100 648.600 685.200 649.800 ;
        RECT 683.100 646.950 685.200 648.600 ;
        RECT 681.450 641.700 683.250 642.000 ;
        RECT 671.550 641.100 683.250 641.700 ;
        RECT 671.550 640.500 689.850 641.100 ;
        RECT 671.550 639.600 672.450 640.500 ;
        RECT 681.450 640.200 689.850 640.500 ;
        RECT 671.550 637.800 673.950 639.600 ;
        RECT 662.100 627.000 663.900 633.600 ;
        RECT 665.100 627.600 666.900 633.600 ;
        RECT 668.100 627.000 669.900 633.600 ;
        RECT 672.150 627.600 673.950 637.800 ;
        RECT 675.150 627.000 676.950 639.600 ;
        RECT 686.250 638.700 688.050 639.300 ;
        RECT 680.250 637.500 688.050 638.700 ;
        RECT 688.950 638.100 689.850 640.200 ;
        RECT 691.950 640.200 692.850 652.800 ;
        RECT 704.250 649.050 705.450 656.400 ;
        RECT 716.700 649.050 717.900 659.400 ;
        RECT 734.400 649.050 735.300 659.400 ;
        RECT 747.000 651.450 751.050 652.050 ;
        RECT 746.550 649.950 751.050 651.450 ;
        RECT 699.150 647.250 705.450 649.050 ;
        RECT 700.950 646.950 705.450 647.250 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 695.550 644.100 697.650 644.400 ;
        RECT 701.550 644.100 703.350 644.250 ;
        RECT 695.550 642.900 703.350 644.100 ;
        RECT 695.550 642.300 697.650 642.900 ;
        RECT 701.550 642.450 703.350 642.900 ;
        RECT 691.950 639.300 696.750 640.200 ;
        RECT 704.250 639.600 705.450 646.950 ;
        RECT 695.550 638.400 696.750 639.300 ;
        RECT 692.850 638.100 694.650 638.400 ;
        RECT 680.250 636.600 682.350 637.500 ;
        RECT 688.950 637.200 694.650 638.100 ;
        RECT 692.850 636.600 694.650 637.200 ;
        RECT 695.550 636.600 698.550 638.400 ;
        RECT 680.550 627.600 682.350 636.600 ;
        RECT 684.450 635.550 686.250 636.300 ;
        RECT 689.250 635.550 691.050 636.300 ;
        RECT 684.450 634.500 691.050 635.550 ;
        RECT 685.350 627.000 687.150 633.600 ;
        RECT 688.350 627.600 690.150 634.500 ;
        RECT 695.550 633.600 697.650 635.700 ;
        RECT 691.350 627.000 693.150 633.600 ;
        RECT 695.850 627.600 697.650 633.600 ;
        RECT 700.650 627.000 702.450 639.600 ;
        RECT 703.650 627.600 705.450 639.600 ;
        RECT 716.700 633.600 717.900 646.950 ;
        RECT 719.100 645.150 720.900 646.950 ;
        RECT 731.250 645.150 733.050 646.950 ;
        RECT 734.400 639.600 735.300 646.950 ;
        RECT 737.100 645.150 738.900 646.950 ;
        RECT 736.950 642.450 739.050 643.050 ;
        RECT 746.550 642.450 747.450 649.950 ;
        RECT 752.700 649.050 753.900 659.400 ;
        RECT 767.700 655.200 769.500 662.400 ;
        RECT 772.800 656.400 774.600 663.000 ;
        RECT 785.400 656.400 787.200 663.000 ;
        RECT 790.500 655.200 792.300 662.400 ;
        RECT 803.100 661.500 810.900 662.400 ;
        RECT 803.100 656.400 804.900 661.500 ;
        RECT 806.100 656.400 807.900 660.600 ;
        RECT 809.100 657.000 810.900 661.500 ;
        RECT 812.100 657.900 813.900 663.000 ;
        RECT 815.100 657.000 816.900 662.400 ;
        RECT 819.150 658.200 820.950 662.400 ;
        RECT 767.700 654.300 771.900 655.200 ;
        RECT 767.100 649.050 768.900 650.850 ;
        RECT 770.700 649.050 771.900 654.300 ;
        RECT 788.100 654.300 792.300 655.200 ;
        RECT 806.700 654.900 807.600 656.400 ;
        RECT 809.100 656.100 816.900 657.000 ;
        RECT 818.550 656.400 820.950 658.200 ;
        RECT 822.150 656.400 823.950 663.000 ;
        RECT 826.950 660.300 828.750 662.400 ;
        RECT 825.150 659.400 828.750 660.300 ;
        RECT 831.450 659.400 833.250 663.000 ;
        RECT 834.750 659.400 836.550 662.400 ;
        RECT 837.750 659.400 839.550 663.000 ;
        RECT 842.250 659.400 844.050 662.400 ;
        RECT 824.850 658.800 828.750 659.400 ;
        RECT 824.850 657.300 826.950 658.800 ;
        RECT 834.750 658.500 835.800 659.400 ;
        RECT 775.950 651.450 780.000 652.050 ;
        RECT 772.950 649.050 774.750 650.850 ;
        RECT 775.950 649.950 780.450 651.450 ;
        RECT 751.950 646.950 754.050 649.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 766.950 646.950 769.050 649.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 736.950 641.550 747.450 642.450 ;
        RECT 736.950 640.950 739.050 641.550 ;
        RECT 716.100 627.600 717.900 633.600 ;
        RECT 719.100 627.000 720.900 633.600 ;
        RECT 731.100 627.000 732.900 639.600 ;
        RECT 734.400 638.400 738.000 639.600 ;
        RECT 736.200 627.600 738.000 638.400 ;
        RECT 752.700 633.600 753.900 646.950 ;
        RECT 755.100 645.150 756.900 646.950 ;
        RECT 770.700 633.600 771.900 646.950 ;
        RECT 779.550 646.050 780.450 649.950 ;
        RECT 785.250 649.050 787.050 650.850 ;
        RECT 788.100 649.050 789.300 654.300 ;
        RECT 806.700 653.700 811.050 654.900 ;
        RECT 791.100 649.050 792.900 650.850 ;
        RECT 806.250 649.050 808.050 650.850 ;
        RECT 810.000 649.050 811.050 653.700 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 802.950 646.950 805.050 649.050 ;
        RECT 805.950 646.950 808.050 649.050 ;
        RECT 808.950 646.950 811.050 649.050 ;
        RECT 811.950 649.050 813.750 650.850 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 779.550 644.550 784.050 646.050 ;
        RECT 780.000 643.950 784.050 644.550 ;
        RECT 772.950 642.450 775.050 642.750 ;
        RECT 778.950 642.450 781.050 643.050 ;
        RECT 772.950 641.550 781.050 642.450 ;
        RECT 772.950 640.650 775.050 641.550 ;
        RECT 778.950 640.950 781.050 641.550 ;
        RECT 788.100 633.600 789.300 646.950 ;
        RECT 803.250 645.150 805.050 646.950 ;
        RECT 810.000 639.600 811.050 646.950 ;
        RECT 815.100 645.150 816.900 646.950 ;
        RECT 818.550 641.700 819.450 656.400 ;
        RECT 827.850 655.800 829.650 657.600 ;
        RECT 830.850 657.450 835.800 658.500 ;
        RECT 830.850 656.700 832.650 657.450 ;
        RECT 842.250 657.300 844.650 659.400 ;
        RECT 847.350 656.400 849.150 663.000 ;
        RECT 850.650 656.400 852.450 662.400 ;
        RECT 827.850 654.000 828.900 655.800 ;
        RECT 838.050 654.000 839.850 654.600 ;
        RECT 827.850 652.800 839.850 654.000 ;
        RECT 820.950 651.600 828.900 652.800 ;
        RECT 820.950 649.050 822.750 651.600 ;
        RECT 827.100 651.000 828.900 651.600 ;
        RECT 824.100 649.800 825.900 650.400 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 824.100 648.600 832.200 649.800 ;
        RECT 830.100 646.950 832.200 648.600 ;
        RECT 828.450 641.700 830.250 642.000 ;
        RECT 818.550 641.100 830.250 641.700 ;
        RECT 818.550 640.500 836.850 641.100 ;
        RECT 818.550 639.600 819.450 640.500 ;
        RECT 828.450 640.200 836.850 640.500 ;
        RECT 752.100 627.600 753.900 633.600 ;
        RECT 755.100 627.000 756.900 633.600 ;
        RECT 767.100 627.000 768.900 633.600 ;
        RECT 770.100 627.600 771.900 633.600 ;
        RECT 773.100 627.000 774.900 633.600 ;
        RECT 785.100 627.000 786.900 633.600 ;
        RECT 788.100 627.600 789.900 633.600 ;
        RECT 791.100 627.000 792.900 633.600 ;
        RECT 804.600 627.000 806.400 639.600 ;
        RECT 809.100 627.600 812.400 639.600 ;
        RECT 815.100 627.000 816.900 639.600 ;
        RECT 818.550 637.800 820.950 639.600 ;
        RECT 819.150 627.600 820.950 637.800 ;
        RECT 822.150 627.000 823.950 639.600 ;
        RECT 833.250 638.700 835.050 639.300 ;
        RECT 827.250 637.500 835.050 638.700 ;
        RECT 835.950 638.100 836.850 640.200 ;
        RECT 838.950 640.200 839.850 652.800 ;
        RECT 851.250 649.050 852.450 656.400 ;
        RECT 853.950 657.450 858.000 658.050 ;
        RECT 853.950 655.950 858.450 657.450 ;
        RECT 846.150 647.250 852.450 649.050 ;
        RECT 847.950 646.950 852.450 647.250 ;
        RECT 842.550 644.100 844.650 644.400 ;
        RECT 848.550 644.100 850.350 644.250 ;
        RECT 842.550 642.900 850.350 644.100 ;
        RECT 842.550 642.300 844.650 642.900 ;
        RECT 848.550 642.450 850.350 642.900 ;
        RECT 838.950 639.300 843.750 640.200 ;
        RECT 851.250 639.600 852.450 646.950 ;
        RECT 857.550 645.450 858.450 655.950 ;
        RECT 865.500 654.000 867.300 662.400 ;
        RECT 864.000 652.800 867.300 654.000 ;
        RECT 872.100 653.400 873.900 663.000 ;
        RECT 864.000 649.050 864.900 652.800 ;
        RECT 866.100 649.050 867.900 650.850 ;
        RECT 872.100 649.050 873.900 650.850 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 857.550 644.550 861.450 645.450 ;
        RECT 842.550 638.400 843.750 639.300 ;
        RECT 839.850 638.100 841.650 638.400 ;
        RECT 827.250 636.600 829.350 637.500 ;
        RECT 835.950 637.200 841.650 638.100 ;
        RECT 839.850 636.600 841.650 637.200 ;
        RECT 842.550 636.600 845.550 638.400 ;
        RECT 827.550 627.600 829.350 636.600 ;
        RECT 831.450 635.550 833.250 636.300 ;
        RECT 836.250 635.550 838.050 636.300 ;
        RECT 831.450 634.500 838.050 635.550 ;
        RECT 832.350 627.000 834.150 633.600 ;
        RECT 835.350 627.600 837.150 634.500 ;
        RECT 842.550 633.600 844.650 635.700 ;
        RECT 838.350 627.000 840.150 633.600 ;
        RECT 842.850 627.600 844.650 633.600 ;
        RECT 847.650 627.000 849.450 639.600 ;
        RECT 850.650 627.600 852.450 639.600 ;
        RECT 860.550 636.900 861.450 644.550 ;
        RECT 859.950 634.800 862.050 636.900 ;
        RECT 864.000 634.800 864.900 646.950 ;
        RECT 869.100 645.150 870.900 646.950 ;
        RECT 864.000 633.900 870.600 634.800 ;
        RECT 864.000 633.600 864.900 633.900 ;
        RECT 863.100 627.600 864.900 633.600 ;
        RECT 869.100 633.600 870.600 633.900 ;
        RECT 866.100 627.000 867.900 633.000 ;
        RECT 869.100 627.600 870.900 633.600 ;
        RECT 872.100 627.000 873.900 633.600 ;
        RECT 14.100 617.400 15.900 624.000 ;
        RECT 17.100 617.400 18.900 623.400 ;
        RECT 14.100 601.950 16.200 604.050 ;
        RECT 14.250 600.150 16.050 601.950 ;
        RECT 17.100 597.300 18.000 617.400 ;
        RECT 20.100 612.000 21.900 624.000 ;
        RECT 23.100 611.400 24.900 623.400 ;
        RECT 35.100 617.400 36.900 624.000 ;
        RECT 38.100 617.400 39.900 623.400 ;
        RECT 41.100 617.400 42.900 624.000 ;
        RECT 53.100 617.400 54.900 624.000 ;
        RECT 56.100 617.400 57.900 623.400 ;
        RECT 19.200 604.050 21.000 605.850 ;
        RECT 23.400 604.050 24.300 611.400 ;
        RECT 38.100 604.050 39.300 617.400 ;
        RECT 48.000 606.450 52.050 607.050 ;
        RECT 47.550 604.950 52.050 606.450 ;
        RECT 19.500 601.950 21.600 604.050 ;
        RECT 22.800 601.950 24.900 604.050 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 14.100 596.400 22.500 597.300 ;
        RECT 14.100 588.600 15.900 596.400 ;
        RECT 20.700 595.500 22.500 596.400 ;
        RECT 23.400 594.600 24.300 601.950 ;
        RECT 35.250 600.150 37.050 601.950 ;
        RECT 38.100 596.700 39.300 601.950 ;
        RECT 41.100 600.150 42.900 601.950 ;
        RECT 47.550 601.050 48.450 604.950 ;
        RECT 53.100 604.050 54.900 605.850 ;
        RECT 56.100 604.050 57.300 617.400 ;
        RECT 69.000 612.600 70.800 623.400 ;
        RECT 69.000 611.400 72.600 612.600 ;
        RECT 74.100 611.400 75.900 624.000 ;
        RECT 86.100 617.400 87.900 624.000 ;
        RECT 89.100 617.400 90.900 623.400 ;
        RECT 58.950 606.450 63.000 607.050 ;
        RECT 58.950 604.950 63.450 606.450 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 43.950 599.550 48.450 601.050 ;
        RECT 43.950 598.950 48.000 599.550 ;
        RECT 38.100 595.800 42.300 596.700 ;
        RECT 18.600 588.000 20.400 594.600 ;
        RECT 21.600 592.800 24.300 594.600 ;
        RECT 21.600 588.600 23.400 592.800 ;
        RECT 35.400 588.000 37.200 594.600 ;
        RECT 40.500 588.600 42.300 595.800 ;
        RECT 56.100 591.600 57.300 601.950 ;
        RECT 62.550 600.450 63.450 604.950 ;
        RECT 68.100 604.050 69.900 605.850 ;
        RECT 71.700 604.050 72.600 611.400 ;
        RECT 73.950 609.450 76.050 610.050 ;
        RECT 82.950 609.450 85.050 610.050 ;
        RECT 73.950 608.550 85.050 609.450 ;
        RECT 73.950 607.950 76.050 608.550 ;
        RECT 82.950 607.950 85.050 608.550 ;
        RECT 73.950 604.050 75.750 605.850 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 70.950 601.950 73.050 604.050 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 86.100 601.950 88.200 604.050 ;
        RECT 62.550 599.550 66.450 600.450 ;
        RECT 65.550 598.050 66.450 599.550 ;
        RECT 65.550 596.550 70.050 598.050 ;
        RECT 66.000 595.950 70.050 596.550 ;
        RECT 71.700 591.600 72.600 601.950 ;
        RECT 86.250 600.150 88.050 601.950 ;
        RECT 89.100 597.300 90.000 617.400 ;
        RECT 92.100 612.000 93.900 624.000 ;
        RECT 95.100 611.400 96.900 623.400 ;
        RECT 108.600 612.900 110.400 623.400 ;
        RECT 108.000 611.400 110.400 612.900 ;
        RECT 111.600 611.400 113.400 624.000 ;
        RECT 116.100 611.400 117.900 623.400 ;
        RECT 128.100 617.400 129.900 624.000 ;
        RECT 131.100 617.400 132.900 623.400 ;
        RECT 134.100 617.400 135.900 624.000 ;
        RECT 91.200 604.050 93.000 605.850 ;
        RECT 95.400 604.050 96.300 611.400 ;
        RECT 108.000 604.050 109.200 611.400 ;
        RECT 116.700 609.900 117.900 611.400 ;
        RECT 110.100 608.700 117.900 609.900 ;
        RECT 110.100 608.100 111.900 608.700 ;
        RECT 91.500 601.950 93.600 604.050 ;
        RECT 94.800 601.950 96.900 604.050 ;
        RECT 107.100 601.950 109.200 604.050 ;
        RECT 86.100 596.400 94.500 597.300 ;
        RECT 53.100 588.000 54.900 591.600 ;
        RECT 56.100 588.600 57.900 591.600 ;
        RECT 68.100 588.000 69.900 591.600 ;
        RECT 71.100 588.600 72.900 591.600 ;
        RECT 74.100 588.000 75.900 591.600 ;
        RECT 86.100 588.600 87.900 596.400 ;
        RECT 92.700 595.500 94.500 596.400 ;
        RECT 95.400 594.600 96.300 601.950 ;
        RECT 90.600 588.000 92.400 594.600 ;
        RECT 93.600 592.800 96.300 594.600 ;
        RECT 107.100 594.600 108.000 601.950 ;
        RECT 110.400 597.600 111.300 608.100 ;
        RECT 112.200 604.050 114.000 605.850 ;
        RECT 131.700 604.050 132.900 617.400 ;
        RECT 137.550 611.400 139.350 623.400 ;
        RECT 140.550 611.400 142.350 624.000 ;
        RECT 145.350 617.400 147.150 623.400 ;
        RECT 149.850 617.400 151.650 624.000 ;
        RECT 145.350 615.300 147.450 617.400 ;
        RECT 152.850 616.500 154.650 623.400 ;
        RECT 155.850 617.400 157.650 624.000 ;
        RECT 151.950 615.450 158.550 616.500 ;
        RECT 151.950 614.700 153.750 615.450 ;
        RECT 156.750 614.700 158.550 615.450 ;
        RECT 160.650 614.400 162.450 623.400 ;
        RECT 144.450 612.600 147.450 614.400 ;
        RECT 148.350 613.800 150.150 614.400 ;
        RECT 148.350 612.900 154.050 613.800 ;
        RECT 160.650 613.500 162.750 614.400 ;
        RECT 148.350 612.600 150.150 612.900 ;
        RECT 146.250 611.700 147.450 612.600 ;
        RECT 137.550 604.050 138.750 611.400 ;
        RECT 146.250 610.800 151.050 611.700 ;
        RECT 139.650 608.100 141.450 608.550 ;
        RECT 145.350 608.100 147.450 608.700 ;
        RECT 139.650 606.900 147.450 608.100 ;
        RECT 139.650 606.750 141.450 606.900 ;
        RECT 145.350 606.600 147.450 606.900 ;
        RECT 112.500 601.950 114.600 604.050 ;
        RECT 115.800 601.950 117.900 604.050 ;
        RECT 127.950 601.950 130.050 604.050 ;
        RECT 130.950 601.950 133.050 604.050 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 137.550 603.750 142.050 604.050 ;
        RECT 137.550 601.950 143.850 603.750 ;
        RECT 115.800 600.150 117.600 601.950 ;
        RECT 128.100 600.150 129.900 601.950 ;
        RECT 109.200 596.700 111.300 597.600 ;
        RECT 131.700 596.700 132.900 601.950 ;
        RECT 133.950 600.150 135.750 601.950 ;
        RECT 109.200 595.800 114.600 596.700 ;
        RECT 93.600 588.600 95.400 592.800 ;
        RECT 107.100 588.600 108.900 594.600 ;
        RECT 110.100 588.000 111.900 594.000 ;
        RECT 113.700 591.600 114.600 595.800 ;
        RECT 128.700 595.800 132.900 596.700 ;
        RECT 113.100 588.600 114.900 591.600 ;
        RECT 116.100 588.600 117.900 591.600 ;
        RECT 128.700 588.600 130.500 595.800 ;
        RECT 137.550 594.600 138.750 601.950 ;
        RECT 150.150 598.200 151.050 610.800 ;
        RECT 153.150 610.800 154.050 612.900 ;
        RECT 154.950 612.300 162.750 613.500 ;
        RECT 154.950 611.700 156.750 612.300 ;
        RECT 166.050 611.400 167.850 624.000 ;
        RECT 169.050 613.200 170.850 623.400 ;
        RECT 182.100 617.400 183.900 624.000 ;
        RECT 185.100 617.400 186.900 623.400 ;
        RECT 169.050 611.400 171.450 613.200 ;
        RECT 153.150 610.500 161.550 610.800 ;
        RECT 170.550 610.500 171.450 611.400 ;
        RECT 153.150 609.900 171.450 610.500 ;
        RECT 159.750 609.300 171.450 609.900 ;
        RECT 159.750 609.000 161.550 609.300 ;
        RECT 157.800 602.400 159.900 604.050 ;
        RECT 157.800 601.200 165.900 602.400 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 164.100 600.600 165.900 601.200 ;
        RECT 161.100 599.400 162.900 600.000 ;
        RECT 167.250 599.400 169.050 601.950 ;
        RECT 161.100 598.200 169.050 599.400 ;
        RECT 150.150 597.000 162.150 598.200 ;
        RECT 150.150 596.400 151.950 597.000 ;
        RECT 161.100 595.200 162.150 597.000 ;
        RECT 116.700 588.000 117.900 588.600 ;
        RECT 133.800 588.000 135.600 594.600 ;
        RECT 137.550 588.600 139.350 594.600 ;
        RECT 140.850 588.000 142.650 594.600 ;
        RECT 145.350 591.600 147.750 593.700 ;
        RECT 157.350 593.550 159.150 594.300 ;
        RECT 154.200 592.500 159.150 593.550 ;
        RECT 160.350 593.400 162.150 595.200 ;
        RECT 170.550 594.600 171.450 609.300 ;
        RECT 182.100 604.050 183.900 605.850 ;
        RECT 185.100 604.050 186.300 617.400 ;
        RECT 188.550 611.400 190.350 623.400 ;
        RECT 191.550 611.400 193.350 624.000 ;
        RECT 196.350 617.400 198.150 623.400 ;
        RECT 200.850 617.400 202.650 624.000 ;
        RECT 196.350 615.300 198.450 617.400 ;
        RECT 203.850 616.500 205.650 623.400 ;
        RECT 206.850 617.400 208.650 624.000 ;
        RECT 202.950 615.450 209.550 616.500 ;
        RECT 202.950 614.700 204.750 615.450 ;
        RECT 207.750 614.700 209.550 615.450 ;
        RECT 211.650 614.400 213.450 623.400 ;
        RECT 195.450 612.600 198.450 614.400 ;
        RECT 199.350 613.800 201.150 614.400 ;
        RECT 199.350 612.900 205.050 613.800 ;
        RECT 211.650 613.500 213.750 614.400 ;
        RECT 199.350 612.600 201.150 612.900 ;
        RECT 197.250 611.700 198.450 612.600 ;
        RECT 188.550 604.050 189.750 611.400 ;
        RECT 197.250 610.800 202.050 611.700 ;
        RECT 190.650 608.100 192.450 608.550 ;
        RECT 196.350 608.100 198.450 608.700 ;
        RECT 190.650 606.900 198.450 608.100 ;
        RECT 190.650 606.750 192.450 606.900 ;
        RECT 196.350 606.600 198.450 606.900 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 188.550 603.750 193.050 604.050 ;
        RECT 188.550 601.950 194.850 603.750 ;
        RECT 154.200 591.600 155.250 592.500 ;
        RECT 163.050 592.200 165.150 593.700 ;
        RECT 161.250 591.600 165.150 592.200 ;
        RECT 145.950 588.600 147.750 591.600 ;
        RECT 150.450 588.000 152.250 591.600 ;
        RECT 153.450 588.600 155.250 591.600 ;
        RECT 156.750 588.000 158.550 591.600 ;
        RECT 161.250 590.700 164.850 591.600 ;
        RECT 161.250 588.600 163.050 590.700 ;
        RECT 166.050 588.000 167.850 594.600 ;
        RECT 169.050 592.800 171.450 594.600 ;
        RECT 169.050 588.600 170.850 592.800 ;
        RECT 185.100 591.600 186.300 601.950 ;
        RECT 188.550 594.600 189.750 601.950 ;
        RECT 201.150 598.200 202.050 610.800 ;
        RECT 204.150 610.800 205.050 612.900 ;
        RECT 205.950 612.300 213.750 613.500 ;
        RECT 205.950 611.700 207.750 612.300 ;
        RECT 217.050 611.400 218.850 624.000 ;
        RECT 220.050 613.200 221.850 623.400 ;
        RECT 220.050 611.400 222.450 613.200 ;
        RECT 233.400 611.400 235.200 624.000 ;
        RECT 238.500 612.900 240.300 623.400 ;
        RECT 241.500 617.400 243.300 624.000 ;
        RECT 241.200 614.100 243.000 615.900 ;
        RECT 246.150 613.200 247.950 623.400 ;
        RECT 238.500 611.400 240.900 612.900 ;
        RECT 204.150 610.500 212.550 610.800 ;
        RECT 221.550 610.500 222.450 611.400 ;
        RECT 204.150 609.900 222.450 610.500 ;
        RECT 210.750 609.300 222.450 609.900 ;
        RECT 210.750 609.000 212.550 609.300 ;
        RECT 208.800 602.400 210.900 604.050 ;
        RECT 208.800 601.200 216.900 602.400 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 215.100 600.600 216.900 601.200 ;
        RECT 212.100 599.400 213.900 600.000 ;
        RECT 218.250 599.400 220.050 601.950 ;
        RECT 212.100 598.200 220.050 599.400 ;
        RECT 201.150 597.000 213.150 598.200 ;
        RECT 201.150 596.400 202.950 597.000 ;
        RECT 212.100 595.200 213.150 597.000 ;
        RECT 182.100 588.000 183.900 591.600 ;
        RECT 185.100 588.600 186.900 591.600 ;
        RECT 188.550 588.600 190.350 594.600 ;
        RECT 191.850 588.000 193.650 594.600 ;
        RECT 196.350 591.600 198.750 593.700 ;
        RECT 208.350 593.550 210.150 594.300 ;
        RECT 205.200 592.500 210.150 593.550 ;
        RECT 211.350 593.400 213.150 595.200 ;
        RECT 221.550 594.600 222.450 609.300 ;
        RECT 233.100 604.050 234.900 605.850 ;
        RECT 239.700 604.050 240.900 611.400 ;
        RECT 245.550 611.400 247.950 613.200 ;
        RECT 249.150 611.400 250.950 624.000 ;
        RECT 254.550 614.400 256.350 623.400 ;
        RECT 259.350 617.400 261.150 624.000 ;
        RECT 262.350 616.500 264.150 623.400 ;
        RECT 265.350 617.400 267.150 624.000 ;
        RECT 269.850 617.400 271.650 623.400 ;
        RECT 258.450 615.450 265.050 616.500 ;
        RECT 258.450 614.700 260.250 615.450 ;
        RECT 263.250 614.700 265.050 615.450 ;
        RECT 269.550 615.300 271.650 617.400 ;
        RECT 254.250 613.500 256.350 614.400 ;
        RECT 266.850 613.800 268.650 614.400 ;
        RECT 254.250 612.300 262.050 613.500 ;
        RECT 260.250 611.700 262.050 612.300 ;
        RECT 262.950 612.900 268.650 613.800 ;
        RECT 245.550 610.500 246.450 611.400 ;
        RECT 262.950 610.800 263.850 612.900 ;
        RECT 266.850 612.600 268.650 612.900 ;
        RECT 269.550 612.600 272.550 614.400 ;
        RECT 269.550 611.700 270.750 612.600 ;
        RECT 255.450 610.500 263.850 610.800 ;
        RECT 245.550 609.900 263.850 610.500 ;
        RECT 265.950 610.800 270.750 611.700 ;
        RECT 274.650 611.400 276.450 624.000 ;
        RECT 277.650 611.400 279.450 623.400 ;
        RECT 290.100 612.600 291.900 623.400 ;
        RECT 293.100 613.500 294.900 624.000 ;
        RECT 296.100 622.500 303.900 623.400 ;
        RECT 296.100 612.600 297.900 622.500 ;
        RECT 290.100 611.700 297.900 612.600 ;
        RECT 245.550 609.300 257.250 609.900 ;
        RECT 232.950 601.950 235.050 604.050 ;
        RECT 235.950 601.950 238.050 604.050 ;
        RECT 238.950 601.950 241.050 604.050 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 236.100 600.150 237.900 601.950 ;
        RECT 239.700 597.600 240.900 601.950 ;
        RECT 242.100 600.150 243.900 601.950 ;
        RECT 239.700 596.700 243.300 597.600 ;
        RECT 205.200 591.600 206.250 592.500 ;
        RECT 214.050 592.200 216.150 593.700 ;
        RECT 212.250 591.600 216.150 592.200 ;
        RECT 196.950 588.600 198.750 591.600 ;
        RECT 201.450 588.000 203.250 591.600 ;
        RECT 204.450 588.600 206.250 591.600 ;
        RECT 207.750 588.000 209.550 591.600 ;
        RECT 212.250 590.700 215.850 591.600 ;
        RECT 212.250 588.600 214.050 590.700 ;
        RECT 217.050 588.000 218.850 594.600 ;
        RECT 220.050 592.800 222.450 594.600 ;
        RECT 233.100 593.700 240.900 595.050 ;
        RECT 220.050 588.600 221.850 592.800 ;
        RECT 233.100 588.600 234.900 593.700 ;
        RECT 236.100 588.000 237.900 592.800 ;
        RECT 239.100 588.600 240.900 593.700 ;
        RECT 242.100 594.600 243.300 596.700 ;
        RECT 245.550 594.600 246.450 609.300 ;
        RECT 255.450 609.000 257.250 609.300 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 257.100 602.400 259.200 604.050 ;
        RECT 247.950 599.400 249.750 601.950 ;
        RECT 251.100 601.200 259.200 602.400 ;
        RECT 251.100 600.600 252.900 601.200 ;
        RECT 254.100 599.400 255.900 600.000 ;
        RECT 247.950 598.200 255.900 599.400 ;
        RECT 265.950 598.200 266.850 610.800 ;
        RECT 269.550 608.100 271.650 608.700 ;
        RECT 275.550 608.100 277.350 608.550 ;
        RECT 269.550 606.900 277.350 608.100 ;
        RECT 269.550 606.600 271.650 606.900 ;
        RECT 275.550 606.750 277.350 606.900 ;
        RECT 278.250 604.050 279.450 611.400 ;
        RECT 299.100 610.500 300.900 621.600 ;
        RECT 302.100 611.400 303.900 622.500 ;
        RECT 305.550 611.400 307.350 623.400 ;
        RECT 308.550 611.400 310.350 624.000 ;
        RECT 313.350 617.400 315.150 623.400 ;
        RECT 317.850 617.400 319.650 624.000 ;
        RECT 313.350 615.300 315.450 617.400 ;
        RECT 320.850 616.500 322.650 623.400 ;
        RECT 323.850 617.400 325.650 624.000 ;
        RECT 319.950 615.450 326.550 616.500 ;
        RECT 319.950 614.700 321.750 615.450 ;
        RECT 324.750 614.700 326.550 615.450 ;
        RECT 328.650 614.400 330.450 623.400 ;
        RECT 312.450 612.600 315.450 614.400 ;
        RECT 316.350 613.800 318.150 614.400 ;
        RECT 316.350 612.900 322.050 613.800 ;
        RECT 328.650 613.500 330.750 614.400 ;
        RECT 316.350 612.600 318.150 612.900 ;
        RECT 314.250 611.700 315.450 612.600 ;
        RECT 296.100 609.600 300.900 610.500 ;
        RECT 293.250 604.050 295.050 605.850 ;
        RECT 296.100 604.050 297.000 609.600 ;
        RECT 299.100 604.050 300.900 605.850 ;
        RECT 305.550 604.050 306.750 611.400 ;
        RECT 314.250 610.800 319.050 611.700 ;
        RECT 307.650 608.100 309.450 608.550 ;
        RECT 313.350 608.100 315.450 608.700 ;
        RECT 307.650 606.900 315.450 608.100 ;
        RECT 307.650 606.750 309.450 606.900 ;
        RECT 313.350 606.600 315.450 606.900 ;
        RECT 274.950 603.750 279.450 604.050 ;
        RECT 273.150 601.950 279.450 603.750 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 305.550 603.750 310.050 604.050 ;
        RECT 305.550 601.950 311.850 603.750 ;
        RECT 254.850 597.000 266.850 598.200 ;
        RECT 254.850 595.200 255.900 597.000 ;
        RECT 265.050 596.400 266.850 597.000 ;
        RECT 242.100 588.600 243.900 594.600 ;
        RECT 245.550 592.800 247.950 594.600 ;
        RECT 246.150 588.600 247.950 592.800 ;
        RECT 249.150 588.000 250.950 594.600 ;
        RECT 251.850 592.200 253.950 593.700 ;
        RECT 254.850 593.400 256.650 595.200 ;
        RECT 278.250 594.600 279.450 601.950 ;
        RECT 290.250 600.150 292.050 601.950 ;
        RECT 296.100 594.600 297.300 601.950 ;
        RECT 302.100 600.150 303.900 601.950 ;
        RECT 305.550 594.600 306.750 601.950 ;
        RECT 318.150 598.200 319.050 610.800 ;
        RECT 321.150 610.800 322.050 612.900 ;
        RECT 322.950 612.300 330.750 613.500 ;
        RECT 322.950 611.700 324.750 612.300 ;
        RECT 334.050 611.400 335.850 624.000 ;
        RECT 337.050 613.200 338.850 623.400 ;
        RECT 337.050 611.400 339.450 613.200 ;
        RECT 351.000 612.600 352.800 623.400 ;
        RECT 351.000 611.400 354.600 612.600 ;
        RECT 356.100 611.400 357.900 624.000 ;
        RECT 369.000 612.600 370.800 623.400 ;
        RECT 369.000 611.400 372.600 612.600 ;
        RECT 374.100 611.400 375.900 624.000 ;
        RECT 386.100 612.300 387.900 623.400 ;
        RECT 389.100 613.200 390.900 624.000 ;
        RECT 392.100 612.300 393.900 623.400 ;
        RECT 386.100 611.400 393.900 612.300 ;
        RECT 395.100 611.400 396.900 623.400 ;
        RECT 399.150 613.200 400.950 623.400 ;
        RECT 398.550 611.400 400.950 613.200 ;
        RECT 402.150 611.400 403.950 624.000 ;
        RECT 407.550 614.400 409.350 623.400 ;
        RECT 412.350 617.400 414.150 624.000 ;
        RECT 415.350 616.500 417.150 623.400 ;
        RECT 418.350 617.400 420.150 624.000 ;
        RECT 422.850 617.400 424.650 623.400 ;
        RECT 411.450 615.450 418.050 616.500 ;
        RECT 411.450 614.700 413.250 615.450 ;
        RECT 416.250 614.700 418.050 615.450 ;
        RECT 422.550 615.300 424.650 617.400 ;
        RECT 407.250 613.500 409.350 614.400 ;
        RECT 419.850 613.800 421.650 614.400 ;
        RECT 407.250 612.300 415.050 613.500 ;
        RECT 413.250 611.700 415.050 612.300 ;
        RECT 415.950 612.900 421.650 613.800 ;
        RECT 321.150 610.500 329.550 610.800 ;
        RECT 338.550 610.500 339.450 611.400 ;
        RECT 321.150 609.900 339.450 610.500 ;
        RECT 327.750 609.300 339.450 609.900 ;
        RECT 327.750 609.000 329.550 609.300 ;
        RECT 325.800 602.400 327.900 604.050 ;
        RECT 325.800 601.200 333.900 602.400 ;
        RECT 334.950 601.950 337.050 604.050 ;
        RECT 332.100 600.600 333.900 601.200 ;
        RECT 329.100 599.400 330.900 600.000 ;
        RECT 335.250 599.400 337.050 601.950 ;
        RECT 329.100 598.200 337.050 599.400 ;
        RECT 318.150 597.000 330.150 598.200 ;
        RECT 318.150 596.400 319.950 597.000 ;
        RECT 329.100 595.200 330.150 597.000 ;
        RECT 257.850 593.550 259.650 594.300 ;
        RECT 257.850 592.500 262.800 593.550 ;
        RECT 251.850 591.600 255.750 592.200 ;
        RECT 261.750 591.600 262.800 592.500 ;
        RECT 269.250 591.600 271.650 593.700 ;
        RECT 252.150 590.700 255.750 591.600 ;
        RECT 253.950 588.600 255.750 590.700 ;
        RECT 258.450 588.000 260.250 591.600 ;
        RECT 261.750 588.600 263.550 591.600 ;
        RECT 264.750 588.000 266.550 591.600 ;
        RECT 269.250 588.600 271.050 591.600 ;
        RECT 274.350 588.000 276.150 594.600 ;
        RECT 277.650 588.600 279.450 594.600 ;
        RECT 290.700 588.000 292.500 594.600 ;
        RECT 295.200 588.600 297.000 594.600 ;
        RECT 299.700 588.000 301.500 594.600 ;
        RECT 305.550 588.600 307.350 594.600 ;
        RECT 308.850 588.000 310.650 594.600 ;
        RECT 313.350 591.600 315.750 593.700 ;
        RECT 325.350 593.550 327.150 594.300 ;
        RECT 322.200 592.500 327.150 593.550 ;
        RECT 328.350 593.400 330.150 595.200 ;
        RECT 338.550 594.600 339.450 609.300 ;
        RECT 350.100 604.050 351.900 605.850 ;
        RECT 353.700 604.050 354.600 611.400 ;
        RECT 355.950 604.050 357.750 605.850 ;
        RECT 368.100 604.050 369.900 605.850 ;
        RECT 371.700 604.050 372.600 611.400 ;
        RECT 373.950 609.450 376.050 610.050 ;
        RECT 391.950 609.450 394.050 610.050 ;
        RECT 373.950 608.550 394.050 609.450 ;
        RECT 373.950 607.950 376.050 608.550 ;
        RECT 391.950 607.950 394.050 608.550 ;
        RECT 373.950 604.050 375.750 605.850 ;
        RECT 389.250 604.050 391.050 605.850 ;
        RECT 395.700 604.050 396.600 611.400 ;
        RECT 398.550 610.500 399.450 611.400 ;
        RECT 415.950 610.800 416.850 612.900 ;
        RECT 419.850 612.600 421.650 612.900 ;
        RECT 422.550 612.600 425.550 614.400 ;
        RECT 422.550 611.700 423.750 612.600 ;
        RECT 408.450 610.500 416.850 610.800 ;
        RECT 398.550 609.900 416.850 610.500 ;
        RECT 418.950 610.800 423.750 611.700 ;
        RECT 427.650 611.400 429.450 624.000 ;
        RECT 430.650 611.400 432.450 623.400 ;
        RECT 443.700 617.400 445.500 624.000 ;
        RECT 444.000 614.100 445.800 615.900 ;
        RECT 446.700 612.900 448.500 623.400 ;
        RECT 398.550 609.300 410.250 609.900 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 352.950 601.950 355.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 322.200 591.600 323.250 592.500 ;
        RECT 331.050 592.200 333.150 593.700 ;
        RECT 329.250 591.600 333.150 592.200 ;
        RECT 313.950 588.600 315.750 591.600 ;
        RECT 318.450 588.000 320.250 591.600 ;
        RECT 321.450 588.600 323.250 591.600 ;
        RECT 324.750 588.000 326.550 591.600 ;
        RECT 329.250 590.700 332.850 591.600 ;
        RECT 329.250 588.600 331.050 590.700 ;
        RECT 334.050 588.000 335.850 594.600 ;
        RECT 337.050 592.800 339.450 594.600 ;
        RECT 337.050 588.600 338.850 592.800 ;
        RECT 353.700 591.600 354.600 601.950 ;
        RECT 371.700 591.600 372.600 601.950 ;
        RECT 386.100 600.150 387.900 601.950 ;
        RECT 392.250 600.150 394.050 601.950 ;
        RECT 395.700 594.600 396.600 601.950 ;
        RECT 350.100 588.000 351.900 591.600 ;
        RECT 353.100 588.600 354.900 591.600 ;
        RECT 356.100 588.000 357.900 591.600 ;
        RECT 368.100 588.000 369.900 591.600 ;
        RECT 371.100 588.600 372.900 591.600 ;
        RECT 374.100 588.000 375.900 591.600 ;
        RECT 387.000 588.000 388.800 594.600 ;
        RECT 391.500 593.400 396.600 594.600 ;
        RECT 398.550 594.600 399.450 609.300 ;
        RECT 408.450 609.000 410.250 609.300 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 410.100 602.400 412.200 604.050 ;
        RECT 400.950 599.400 402.750 601.950 ;
        RECT 404.100 601.200 412.200 602.400 ;
        RECT 404.100 600.600 405.900 601.200 ;
        RECT 407.100 599.400 408.900 600.000 ;
        RECT 400.950 598.200 408.900 599.400 ;
        RECT 418.950 598.200 419.850 610.800 ;
        RECT 422.550 608.100 424.650 608.700 ;
        RECT 428.550 608.100 430.350 608.550 ;
        RECT 422.550 606.900 430.350 608.100 ;
        RECT 422.550 606.600 424.650 606.900 ;
        RECT 428.550 606.750 430.350 606.900 ;
        RECT 431.250 604.050 432.450 611.400 ;
        RECT 446.100 611.400 448.500 612.900 ;
        RECT 451.800 611.400 453.600 624.000 ;
        RECT 464.100 617.400 465.900 624.000 ;
        RECT 467.100 617.400 468.900 623.400 ;
        RECT 470.100 618.000 471.900 624.000 ;
        RECT 467.400 617.100 468.900 617.400 ;
        RECT 473.100 617.400 474.900 623.400 ;
        RECT 473.100 617.100 474.000 617.400 ;
        RECT 467.400 616.200 474.000 617.100 ;
        RECT 446.100 604.050 447.300 611.400 ;
        RECT 459.000 606.450 463.050 607.050 ;
        RECT 452.100 604.050 453.900 605.850 ;
        RECT 458.550 604.950 463.050 606.450 ;
        RECT 427.950 603.750 432.450 604.050 ;
        RECT 426.150 601.950 432.450 603.750 ;
        RECT 442.950 601.950 445.050 604.050 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 407.850 597.000 419.850 598.200 ;
        RECT 407.850 595.200 408.900 597.000 ;
        RECT 418.050 596.400 419.850 597.000 ;
        RECT 391.500 588.600 393.300 593.400 ;
        RECT 398.550 592.800 400.950 594.600 ;
        RECT 394.500 588.000 396.300 591.600 ;
        RECT 399.150 588.600 400.950 592.800 ;
        RECT 402.150 588.000 403.950 594.600 ;
        RECT 404.850 592.200 406.950 593.700 ;
        RECT 407.850 593.400 409.650 595.200 ;
        RECT 431.250 594.600 432.450 601.950 ;
        RECT 443.100 600.150 444.900 601.950 ;
        RECT 446.100 597.600 447.300 601.950 ;
        RECT 449.100 600.150 450.900 601.950 ;
        RECT 458.550 601.050 459.450 604.950 ;
        RECT 467.100 604.050 468.900 605.850 ;
        RECT 473.100 604.050 474.000 616.200 ;
        RECT 485.400 611.400 487.200 624.000 ;
        RECT 490.500 612.900 492.300 623.400 ;
        RECT 493.500 617.400 495.300 624.000 ;
        RECT 506.100 617.400 507.900 624.000 ;
        RECT 509.100 617.400 510.900 623.400 ;
        RECT 512.100 617.400 513.900 624.000 ;
        RECT 524.100 617.400 525.900 623.400 ;
        RECT 493.200 614.100 495.000 615.900 ;
        RECT 490.500 611.400 492.900 612.900 ;
        RECT 485.100 604.050 486.900 605.850 ;
        RECT 491.700 604.050 492.900 611.400 ;
        RECT 493.950 609.450 496.050 610.050 ;
        RECT 502.950 609.450 505.050 610.050 ;
        RECT 493.950 608.550 505.050 609.450 ;
        RECT 493.950 607.950 496.050 608.550 ;
        RECT 502.950 607.950 505.050 608.550 ;
        RECT 509.100 604.050 510.300 617.400 ;
        RECT 524.100 610.500 525.300 617.400 ;
        RECT 527.100 613.200 528.900 624.000 ;
        RECT 530.100 611.400 531.900 623.400 ;
        RECT 511.950 609.450 514.050 610.050 ;
        RECT 520.950 609.450 523.050 609.900 ;
        RECT 524.100 609.600 529.800 610.500 ;
        RECT 511.950 608.550 523.050 609.450 ;
        RECT 511.950 607.950 514.050 608.550 ;
        RECT 520.950 607.800 523.050 608.550 ;
        RECT 528.000 608.700 529.800 609.600 ;
        RECT 524.400 604.050 526.200 605.850 ;
        RECT 463.950 601.950 466.050 604.050 ;
        RECT 466.950 601.950 469.050 604.050 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 484.950 601.950 487.050 604.050 ;
        RECT 487.950 601.950 490.050 604.050 ;
        RECT 490.950 601.950 493.050 604.050 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 505.950 601.950 508.050 604.050 ;
        RECT 508.950 601.950 511.050 604.050 ;
        RECT 511.950 601.950 514.050 604.050 ;
        RECT 524.400 601.950 526.500 604.050 ;
        RECT 458.550 599.550 463.050 601.050 ;
        RECT 464.100 600.150 465.900 601.950 ;
        RECT 470.100 600.150 471.900 601.950 ;
        RECT 459.000 598.950 463.050 599.550 ;
        RECT 473.100 598.200 474.000 601.950 ;
        RECT 488.100 600.150 489.900 601.950 ;
        RECT 443.700 596.700 447.300 597.600 ;
        RECT 443.700 594.600 444.900 596.700 ;
        RECT 410.850 593.550 412.650 594.300 ;
        RECT 410.850 592.500 415.800 593.550 ;
        RECT 404.850 591.600 408.750 592.200 ;
        RECT 414.750 591.600 415.800 592.500 ;
        RECT 422.250 591.600 424.650 593.700 ;
        RECT 405.150 590.700 408.750 591.600 ;
        RECT 406.950 588.600 408.750 590.700 ;
        RECT 411.450 588.000 413.250 591.600 ;
        RECT 414.750 588.600 416.550 591.600 ;
        RECT 417.750 588.000 419.550 591.600 ;
        RECT 422.250 588.600 424.050 591.600 ;
        RECT 427.350 588.000 429.150 594.600 ;
        RECT 430.650 588.600 432.450 594.600 ;
        RECT 443.100 588.600 444.900 594.600 ;
        RECT 446.100 593.700 453.900 595.050 ;
        RECT 446.100 588.600 447.900 593.700 ;
        RECT 449.100 588.000 450.900 592.800 ;
        RECT 452.100 588.600 453.900 593.700 ;
        RECT 464.100 588.000 465.900 597.600 ;
        RECT 470.700 597.000 474.000 598.200 ;
        RECT 491.700 597.600 492.900 601.950 ;
        RECT 494.100 600.150 495.900 601.950 ;
        RECT 506.250 600.150 508.050 601.950 ;
        RECT 470.700 588.600 472.500 597.000 ;
        RECT 491.700 596.700 495.300 597.600 ;
        RECT 485.100 593.700 492.900 595.050 ;
        RECT 485.100 588.600 486.900 593.700 ;
        RECT 488.100 588.000 489.900 592.800 ;
        RECT 491.100 588.600 492.900 593.700 ;
        RECT 494.100 594.600 495.300 596.700 ;
        RECT 509.100 596.700 510.300 601.950 ;
        RECT 512.100 600.150 513.900 601.950 ;
        RECT 528.000 597.300 528.900 608.700 ;
        RECT 530.700 604.050 531.900 611.400 ;
        RECT 542.100 617.400 543.900 623.400 ;
        RECT 542.100 610.500 543.300 617.400 ;
        RECT 545.100 613.200 546.900 624.000 ;
        RECT 548.100 611.400 549.900 623.400 ;
        RECT 560.100 612.300 561.900 623.400 ;
        RECT 563.100 613.200 564.900 624.000 ;
        RECT 566.100 612.300 567.900 623.400 ;
        RECT 560.100 611.400 567.900 612.300 ;
        RECT 569.100 611.400 570.900 623.400 ;
        RECT 582.000 612.600 583.800 623.400 ;
        RECT 582.000 611.400 585.600 612.600 ;
        RECT 587.100 611.400 588.900 624.000 ;
        RECT 599.100 617.400 600.900 624.000 ;
        RECT 602.100 617.400 603.900 623.400 ;
        RECT 605.100 617.400 606.900 624.000 ;
        RECT 542.100 609.600 547.800 610.500 ;
        RECT 546.000 608.700 547.800 609.600 ;
        RECT 529.800 601.950 531.900 604.050 ;
        RECT 542.400 604.050 544.200 605.850 ;
        RECT 542.400 601.950 544.500 604.050 ;
        RECT 509.100 595.800 513.300 596.700 ;
        RECT 528.000 596.400 529.800 597.300 ;
        RECT 494.100 588.600 495.900 594.600 ;
        RECT 506.400 588.000 508.200 594.600 ;
        RECT 511.500 588.600 513.300 595.800 ;
        RECT 524.100 595.500 529.800 596.400 ;
        RECT 524.100 591.600 525.300 595.500 ;
        RECT 530.700 594.600 531.900 601.950 ;
        RECT 546.000 597.300 546.900 608.700 ;
        RECT 548.700 604.050 549.900 611.400 ;
        RECT 563.250 604.050 565.050 605.850 ;
        RECT 569.700 604.050 570.600 611.400 ;
        RECT 581.100 604.050 582.900 605.850 ;
        RECT 584.700 604.050 585.600 611.400 ;
        RECT 586.950 609.450 589.050 610.050 ;
        RECT 598.950 609.450 601.050 610.050 ;
        RECT 586.950 608.550 601.050 609.450 ;
        RECT 586.950 607.950 589.050 608.550 ;
        RECT 598.950 607.950 601.050 608.550 ;
        RECT 589.950 606.450 594.000 607.050 ;
        RECT 586.950 604.050 588.750 605.850 ;
        RECT 589.950 604.950 594.450 606.450 ;
        RECT 547.800 601.950 549.900 604.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 580.950 601.950 583.050 604.050 ;
        RECT 583.950 601.950 586.050 604.050 ;
        RECT 586.950 601.950 589.050 604.050 ;
        RECT 546.000 596.400 547.800 597.300 ;
        RECT 524.100 588.600 525.900 591.600 ;
        RECT 527.100 588.000 528.900 594.600 ;
        RECT 530.100 588.600 531.900 594.600 ;
        RECT 542.100 595.500 547.800 596.400 ;
        RECT 542.100 591.600 543.300 595.500 ;
        RECT 548.700 594.600 549.900 601.950 ;
        RECT 560.100 600.150 561.900 601.950 ;
        RECT 566.250 600.150 568.050 601.950 ;
        RECT 569.700 594.600 570.600 601.950 ;
        RECT 542.100 588.600 543.900 591.600 ;
        RECT 545.100 588.000 546.900 594.600 ;
        RECT 548.100 588.600 549.900 594.600 ;
        RECT 561.000 588.000 562.800 594.600 ;
        RECT 565.500 593.400 570.600 594.600 ;
        RECT 565.500 588.600 567.300 593.400 ;
        RECT 584.700 591.600 585.600 601.950 ;
        RECT 593.550 601.050 594.450 604.950 ;
        RECT 602.700 604.050 603.900 617.400 ;
        RECT 609.150 613.200 610.950 623.400 ;
        RECT 608.550 611.400 610.950 613.200 ;
        RECT 612.150 611.400 613.950 624.000 ;
        RECT 617.550 614.400 619.350 623.400 ;
        RECT 622.350 617.400 624.150 624.000 ;
        RECT 625.350 616.500 627.150 623.400 ;
        RECT 628.350 617.400 630.150 624.000 ;
        RECT 632.850 617.400 634.650 623.400 ;
        RECT 621.450 615.450 628.050 616.500 ;
        RECT 621.450 614.700 623.250 615.450 ;
        RECT 626.250 614.700 628.050 615.450 ;
        RECT 632.550 615.300 634.650 617.400 ;
        RECT 617.250 613.500 619.350 614.400 ;
        RECT 629.850 613.800 631.650 614.400 ;
        RECT 617.250 612.300 625.050 613.500 ;
        RECT 623.250 611.700 625.050 612.300 ;
        RECT 625.950 612.900 631.650 613.800 ;
        RECT 608.550 610.500 609.450 611.400 ;
        RECT 625.950 610.800 626.850 612.900 ;
        RECT 629.850 612.600 631.650 612.900 ;
        RECT 632.550 612.600 635.550 614.400 ;
        RECT 632.550 611.700 633.750 612.600 ;
        RECT 618.450 610.500 626.850 610.800 ;
        RECT 608.550 609.900 626.850 610.500 ;
        RECT 628.950 610.800 633.750 611.700 ;
        RECT 637.650 611.400 639.450 624.000 ;
        RECT 640.650 611.400 642.450 623.400 ;
        RECT 653.100 617.400 654.900 624.000 ;
        RECT 656.100 617.400 657.900 623.400 ;
        RECT 659.100 617.400 660.900 624.000 ;
        RECT 671.100 617.400 672.900 624.000 ;
        RECT 674.100 617.400 675.900 623.400 ;
        RECT 677.100 617.400 678.900 624.000 ;
        RECT 689.700 617.400 691.500 624.000 ;
        RECT 608.550 609.300 620.250 609.900 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 589.950 599.550 594.450 601.050 ;
        RECT 599.100 600.150 600.900 601.950 ;
        RECT 589.950 598.950 594.000 599.550 ;
        RECT 602.700 596.700 603.900 601.950 ;
        RECT 604.950 600.150 606.750 601.950 ;
        RECT 599.700 595.800 603.900 596.700 ;
        RECT 586.950 594.450 589.050 595.050 ;
        RECT 595.950 594.450 598.050 595.050 ;
        RECT 586.950 593.550 598.050 594.450 ;
        RECT 586.950 592.950 589.050 593.550 ;
        RECT 595.950 592.950 598.050 593.550 ;
        RECT 568.500 588.000 570.300 591.600 ;
        RECT 581.100 588.000 582.900 591.600 ;
        RECT 584.100 588.600 585.900 591.600 ;
        RECT 587.100 588.000 588.900 591.600 ;
        RECT 599.700 588.600 601.500 595.800 ;
        RECT 608.550 594.600 609.450 609.300 ;
        RECT 618.450 609.000 620.250 609.300 ;
        RECT 610.950 601.950 613.050 604.050 ;
        RECT 620.100 602.400 622.200 604.050 ;
        RECT 610.950 599.400 612.750 601.950 ;
        RECT 614.100 601.200 622.200 602.400 ;
        RECT 614.100 600.600 615.900 601.200 ;
        RECT 617.100 599.400 618.900 600.000 ;
        RECT 610.950 598.200 618.900 599.400 ;
        RECT 628.950 598.200 629.850 610.800 ;
        RECT 632.550 608.100 634.650 608.700 ;
        RECT 638.550 608.100 640.350 608.550 ;
        RECT 632.550 606.900 640.350 608.100 ;
        RECT 632.550 606.600 634.650 606.900 ;
        RECT 638.550 606.750 640.350 606.900 ;
        RECT 641.250 604.050 642.450 611.400 ;
        RECT 656.700 604.050 657.900 617.400 ;
        RECT 674.700 604.050 675.900 617.400 ;
        RECT 690.000 614.100 691.800 615.900 ;
        RECT 692.700 612.900 694.500 623.400 ;
        RECT 692.100 611.400 694.500 612.900 ;
        RECT 697.800 611.400 699.600 624.000 ;
        RECT 702.150 613.200 703.950 623.400 ;
        RECT 701.550 611.400 703.950 613.200 ;
        RECT 705.150 611.400 706.950 624.000 ;
        RECT 710.550 614.400 712.350 623.400 ;
        RECT 715.350 617.400 717.150 624.000 ;
        RECT 718.350 616.500 720.150 623.400 ;
        RECT 721.350 617.400 723.150 624.000 ;
        RECT 725.850 617.400 727.650 623.400 ;
        RECT 714.450 615.450 721.050 616.500 ;
        RECT 714.450 614.700 716.250 615.450 ;
        RECT 719.250 614.700 721.050 615.450 ;
        RECT 725.550 615.300 727.650 617.400 ;
        RECT 710.250 613.500 712.350 614.400 ;
        RECT 722.850 613.800 724.650 614.400 ;
        RECT 710.250 612.300 718.050 613.500 ;
        RECT 716.250 611.700 718.050 612.300 ;
        RECT 718.950 612.900 724.650 613.800 ;
        RECT 692.100 604.050 693.300 611.400 ;
        RECT 701.550 610.500 702.450 611.400 ;
        RECT 718.950 610.800 719.850 612.900 ;
        RECT 722.850 612.600 724.650 612.900 ;
        RECT 725.550 612.600 728.550 614.400 ;
        RECT 725.550 611.700 726.750 612.600 ;
        RECT 711.450 610.500 719.850 610.800 ;
        RECT 701.550 609.900 719.850 610.500 ;
        RECT 721.950 610.800 726.750 611.700 ;
        RECT 730.650 611.400 732.450 624.000 ;
        RECT 733.650 611.400 735.450 623.400 ;
        RECT 746.400 611.400 748.200 624.000 ;
        RECT 751.500 612.900 753.300 623.400 ;
        RECT 754.500 617.400 756.300 624.000 ;
        RECT 754.200 614.100 756.000 615.900 ;
        RECT 751.500 611.400 753.900 612.900 ;
        RECT 767.100 612.600 768.900 623.400 ;
        RECT 770.100 613.500 771.900 624.000 ;
        RECT 773.100 622.500 780.900 623.400 ;
        RECT 773.100 612.600 774.900 622.500 ;
        RECT 767.100 611.700 774.900 612.600 ;
        RECT 701.550 609.300 713.250 609.900 ;
        RECT 698.100 604.050 699.900 605.850 ;
        RECT 637.950 603.750 642.450 604.050 ;
        RECT 636.150 601.950 642.450 603.750 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 673.950 601.950 676.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 691.950 601.950 694.050 604.050 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 697.950 601.950 700.050 604.050 ;
        RECT 617.850 597.000 629.850 598.200 ;
        RECT 617.850 595.200 618.900 597.000 ;
        RECT 628.050 596.400 629.850 597.000 ;
        RECT 604.800 588.000 606.600 594.600 ;
        RECT 608.550 592.800 610.950 594.600 ;
        RECT 609.150 588.600 610.950 592.800 ;
        RECT 612.150 588.000 613.950 594.600 ;
        RECT 614.850 592.200 616.950 593.700 ;
        RECT 617.850 593.400 619.650 595.200 ;
        RECT 641.250 594.600 642.450 601.950 ;
        RECT 653.100 600.150 654.900 601.950 ;
        RECT 656.700 596.700 657.900 601.950 ;
        RECT 658.950 600.150 660.750 601.950 ;
        RECT 671.100 600.150 672.900 601.950 ;
        RECT 674.700 596.700 675.900 601.950 ;
        RECT 676.950 600.150 678.750 601.950 ;
        RECT 689.100 600.150 690.900 601.950 ;
        RECT 692.100 597.600 693.300 601.950 ;
        RECT 695.100 600.150 696.900 601.950 ;
        RECT 620.850 593.550 622.650 594.300 ;
        RECT 620.850 592.500 625.800 593.550 ;
        RECT 614.850 591.600 618.750 592.200 ;
        RECT 624.750 591.600 625.800 592.500 ;
        RECT 632.250 591.600 634.650 593.700 ;
        RECT 615.150 590.700 618.750 591.600 ;
        RECT 616.950 588.600 618.750 590.700 ;
        RECT 621.450 588.000 623.250 591.600 ;
        RECT 624.750 588.600 626.550 591.600 ;
        RECT 627.750 588.000 629.550 591.600 ;
        RECT 632.250 588.600 634.050 591.600 ;
        RECT 637.350 588.000 639.150 594.600 ;
        RECT 640.650 588.600 642.450 594.600 ;
        RECT 653.700 595.800 657.900 596.700 ;
        RECT 671.700 595.800 675.900 596.700 ;
        RECT 689.700 596.700 693.300 597.600 ;
        RECT 653.700 588.600 655.500 595.800 ;
        RECT 658.800 588.000 660.600 594.600 ;
        RECT 671.700 588.600 673.500 595.800 ;
        RECT 689.700 594.600 690.900 596.700 ;
        RECT 676.800 588.000 678.600 594.600 ;
        RECT 689.100 588.600 690.900 594.600 ;
        RECT 692.100 593.700 699.900 595.050 ;
        RECT 692.100 588.600 693.900 593.700 ;
        RECT 695.100 588.000 696.900 592.800 ;
        RECT 698.100 588.600 699.900 593.700 ;
        RECT 701.550 594.600 702.450 609.300 ;
        RECT 711.450 609.000 713.250 609.300 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 713.100 602.400 715.200 604.050 ;
        RECT 703.950 599.400 705.750 601.950 ;
        RECT 707.100 601.200 715.200 602.400 ;
        RECT 707.100 600.600 708.900 601.200 ;
        RECT 710.100 599.400 711.900 600.000 ;
        RECT 703.950 598.200 711.900 599.400 ;
        RECT 721.950 598.200 722.850 610.800 ;
        RECT 725.550 608.100 727.650 608.700 ;
        RECT 731.550 608.100 733.350 608.550 ;
        RECT 725.550 606.900 733.350 608.100 ;
        RECT 725.550 606.600 727.650 606.900 ;
        RECT 731.550 606.750 733.350 606.900 ;
        RECT 734.250 604.050 735.450 611.400 ;
        RECT 746.100 604.050 747.900 605.850 ;
        RECT 752.700 604.050 753.900 611.400 ;
        RECT 776.100 610.500 777.900 621.600 ;
        RECT 779.100 611.400 780.900 622.500 ;
        RECT 791.700 617.400 793.500 624.000 ;
        RECT 792.000 614.100 793.800 615.900 ;
        RECT 794.700 612.900 796.500 623.400 ;
        RECT 794.100 611.400 796.500 612.900 ;
        RECT 799.800 611.400 801.600 624.000 ;
        RECT 812.100 617.400 813.900 623.400 ;
        RECT 815.100 617.400 816.900 624.000 ;
        RECT 760.950 609.450 763.050 610.050 ;
        RECT 766.950 609.450 769.050 610.050 ;
        RECT 760.950 608.550 769.050 609.450 ;
        RECT 760.950 607.950 763.050 608.550 ;
        RECT 766.950 607.950 769.050 608.550 ;
        RECT 773.100 609.600 777.900 610.500 ;
        RECT 770.250 604.050 772.050 605.850 ;
        RECT 773.100 604.050 774.000 609.600 ;
        RECT 778.950 609.450 781.050 610.050 ;
        RECT 784.950 609.450 787.050 610.050 ;
        RECT 778.950 608.550 787.050 609.450 ;
        RECT 778.950 607.950 781.050 608.550 ;
        RECT 784.950 607.950 787.050 608.550 ;
        RECT 776.100 604.050 777.900 605.850 ;
        RECT 794.100 604.050 795.300 611.400 ;
        RECT 802.950 606.450 807.000 607.050 ;
        RECT 800.100 604.050 801.900 605.850 ;
        RECT 802.950 604.950 807.450 606.450 ;
        RECT 730.950 603.750 735.450 604.050 ;
        RECT 729.150 601.950 735.450 603.750 ;
        RECT 745.950 601.950 748.050 604.050 ;
        RECT 748.950 601.950 751.050 604.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 766.950 601.950 769.050 604.050 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 710.850 597.000 722.850 598.200 ;
        RECT 710.850 595.200 711.900 597.000 ;
        RECT 721.050 596.400 722.850 597.000 ;
        RECT 701.550 592.800 703.950 594.600 ;
        RECT 702.150 588.600 703.950 592.800 ;
        RECT 705.150 588.000 706.950 594.600 ;
        RECT 707.850 592.200 709.950 593.700 ;
        RECT 710.850 593.400 712.650 595.200 ;
        RECT 734.250 594.600 735.450 601.950 ;
        RECT 749.100 600.150 750.900 601.950 ;
        RECT 752.700 597.600 753.900 601.950 ;
        RECT 755.100 600.150 756.900 601.950 ;
        RECT 767.250 600.150 769.050 601.950 ;
        RECT 752.700 596.700 756.300 597.600 ;
        RECT 713.850 593.550 715.650 594.300 ;
        RECT 713.850 592.500 718.800 593.550 ;
        RECT 707.850 591.600 711.750 592.200 ;
        RECT 717.750 591.600 718.800 592.500 ;
        RECT 725.250 591.600 727.650 593.700 ;
        RECT 708.150 590.700 711.750 591.600 ;
        RECT 709.950 588.600 711.750 590.700 ;
        RECT 714.450 588.000 716.250 591.600 ;
        RECT 717.750 588.600 719.550 591.600 ;
        RECT 720.750 588.000 722.550 591.600 ;
        RECT 725.250 588.600 727.050 591.600 ;
        RECT 730.350 588.000 732.150 594.600 ;
        RECT 733.650 588.600 735.450 594.600 ;
        RECT 746.100 593.700 753.900 595.050 ;
        RECT 746.100 588.600 747.900 593.700 ;
        RECT 749.100 588.000 750.900 592.800 ;
        RECT 752.100 588.600 753.900 593.700 ;
        RECT 755.100 594.600 756.300 596.700 ;
        RECT 773.100 594.600 774.300 601.950 ;
        RECT 779.100 600.150 780.900 601.950 ;
        RECT 791.100 600.150 792.900 601.950 ;
        RECT 794.100 597.600 795.300 601.950 ;
        RECT 797.100 600.150 798.900 601.950 ;
        RECT 806.550 601.050 807.450 604.950 ;
        RECT 812.700 604.050 813.900 617.400 ;
        RECT 819.150 613.200 820.950 623.400 ;
        RECT 818.550 611.400 820.950 613.200 ;
        RECT 822.150 611.400 823.950 624.000 ;
        RECT 827.550 614.400 829.350 623.400 ;
        RECT 832.350 617.400 834.150 624.000 ;
        RECT 835.350 616.500 837.150 623.400 ;
        RECT 838.350 617.400 840.150 624.000 ;
        RECT 842.850 617.400 844.650 623.400 ;
        RECT 831.450 615.450 838.050 616.500 ;
        RECT 831.450 614.700 833.250 615.450 ;
        RECT 836.250 614.700 838.050 615.450 ;
        RECT 842.550 615.300 844.650 617.400 ;
        RECT 827.250 613.500 829.350 614.400 ;
        RECT 839.850 613.800 841.650 614.400 ;
        RECT 827.250 612.300 835.050 613.500 ;
        RECT 833.250 611.700 835.050 612.300 ;
        RECT 835.950 612.900 841.650 613.800 ;
        RECT 818.550 610.500 819.450 611.400 ;
        RECT 835.950 610.800 836.850 612.900 ;
        RECT 839.850 612.600 841.650 612.900 ;
        RECT 842.550 612.600 845.550 614.400 ;
        RECT 842.550 611.700 843.750 612.600 ;
        RECT 828.450 610.500 836.850 610.800 ;
        RECT 818.550 609.900 836.850 610.500 ;
        RECT 838.950 610.800 843.750 611.700 ;
        RECT 847.650 611.400 849.450 624.000 ;
        RECT 850.650 611.400 852.450 623.400 ;
        RECT 863.100 617.400 864.900 624.000 ;
        RECT 866.100 617.400 867.900 623.400 ;
        RECT 818.550 609.300 830.250 609.900 ;
        RECT 815.100 604.050 816.900 605.850 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 601.950 817.050 604.050 ;
        RECT 802.950 599.550 807.450 601.050 ;
        RECT 802.950 598.950 807.000 599.550 ;
        RECT 791.700 596.700 795.300 597.600 ;
        RECT 791.700 594.600 792.900 596.700 ;
        RECT 755.100 588.600 756.900 594.600 ;
        RECT 767.700 588.000 769.500 594.600 ;
        RECT 772.200 588.600 774.000 594.600 ;
        RECT 776.700 588.000 778.500 594.600 ;
        RECT 791.100 588.600 792.900 594.600 ;
        RECT 794.100 593.700 801.900 595.050 ;
        RECT 794.100 588.600 795.900 593.700 ;
        RECT 797.100 588.000 798.900 592.800 ;
        RECT 800.100 588.600 801.900 593.700 ;
        RECT 812.700 591.600 813.900 601.950 ;
        RECT 818.550 594.600 819.450 609.300 ;
        RECT 828.450 609.000 830.250 609.300 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 830.100 602.400 832.200 604.050 ;
        RECT 820.950 599.400 822.750 601.950 ;
        RECT 824.100 601.200 832.200 602.400 ;
        RECT 824.100 600.600 825.900 601.200 ;
        RECT 827.100 599.400 828.900 600.000 ;
        RECT 820.950 598.200 828.900 599.400 ;
        RECT 838.950 598.200 839.850 610.800 ;
        RECT 842.550 608.100 844.650 608.700 ;
        RECT 848.550 608.100 850.350 608.550 ;
        RECT 842.550 606.900 850.350 608.100 ;
        RECT 842.550 606.600 844.650 606.900 ;
        RECT 848.550 606.750 850.350 606.900 ;
        RECT 851.250 604.050 852.450 611.400 ;
        RECT 861.000 609.450 865.050 610.050 ;
        RECT 860.550 607.950 865.050 609.450 ;
        RECT 860.550 606.450 861.450 607.950 ;
        RECT 847.950 603.750 852.450 604.050 ;
        RECT 846.150 601.950 852.450 603.750 ;
        RECT 827.850 597.000 839.850 598.200 ;
        RECT 827.850 595.200 828.900 597.000 ;
        RECT 838.050 596.400 839.850 597.000 ;
        RECT 818.550 592.800 820.950 594.600 ;
        RECT 812.100 588.600 813.900 591.600 ;
        RECT 815.100 588.000 816.900 591.600 ;
        RECT 819.150 588.600 820.950 592.800 ;
        RECT 822.150 588.000 823.950 594.600 ;
        RECT 824.850 592.200 826.950 593.700 ;
        RECT 827.850 593.400 829.650 595.200 ;
        RECT 851.250 594.600 852.450 601.950 ;
        RECT 857.550 605.550 861.450 606.450 ;
        RECT 857.550 601.050 858.450 605.550 ;
        RECT 863.100 604.050 864.900 605.850 ;
        RECT 866.100 604.050 867.300 617.400 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 857.550 599.550 862.050 601.050 ;
        RECT 858.000 598.950 862.050 599.550 ;
        RECT 830.850 593.550 832.650 594.300 ;
        RECT 830.850 592.500 835.800 593.550 ;
        RECT 824.850 591.600 828.750 592.200 ;
        RECT 834.750 591.600 835.800 592.500 ;
        RECT 842.250 591.600 844.650 593.700 ;
        RECT 825.150 590.700 828.750 591.600 ;
        RECT 826.950 588.600 828.750 590.700 ;
        RECT 831.450 588.000 833.250 591.600 ;
        RECT 834.750 588.600 836.550 591.600 ;
        RECT 837.750 588.000 839.550 591.600 ;
        RECT 842.250 588.600 844.050 591.600 ;
        RECT 847.350 588.000 849.150 594.600 ;
        RECT 850.650 588.600 852.450 594.600 ;
        RECT 866.100 591.600 867.300 601.950 ;
        RECT 863.100 588.000 864.900 591.600 ;
        RECT 866.100 588.600 867.900 591.600 ;
        RECT 11.700 577.200 13.500 584.400 ;
        RECT 16.800 578.400 18.600 585.000 ;
        RECT 29.100 579.300 30.900 584.400 ;
        RECT 32.100 580.200 33.900 585.000 ;
        RECT 35.100 579.300 36.900 584.400 ;
        RECT 29.100 577.950 36.900 579.300 ;
        RECT 38.100 578.400 39.900 584.400 ;
        RECT 53.100 581.400 54.900 585.000 ;
        RECT 56.100 581.400 57.900 584.400 ;
        RECT 11.700 576.300 15.900 577.200 ;
        RECT 38.100 576.300 39.300 578.400 ;
        RECT 11.100 571.050 12.900 572.850 ;
        RECT 14.700 571.050 15.900 576.300 ;
        RECT 35.700 575.400 39.300 576.300 ;
        RECT 16.950 571.050 18.750 572.850 ;
        RECT 32.100 571.050 33.900 572.850 ;
        RECT 35.700 571.050 36.900 575.400 ;
        RECT 38.100 571.050 39.900 572.850 ;
        RECT 56.100 571.050 57.300 581.400 ;
        RECT 68.100 579.300 69.900 584.400 ;
        RECT 71.100 580.200 72.900 585.000 ;
        RECT 74.100 579.300 75.900 584.400 ;
        RECT 68.100 577.950 75.900 579.300 ;
        RECT 77.100 578.400 78.900 584.400 ;
        RECT 89.100 578.400 90.900 584.400 ;
        RECT 77.100 576.300 78.300 578.400 ;
        RECT 74.700 575.400 78.300 576.300 ;
        RECT 89.700 576.300 90.900 578.400 ;
        RECT 92.100 579.300 93.900 584.400 ;
        RECT 95.100 580.200 96.900 585.000 ;
        RECT 98.100 579.300 99.900 584.400 ;
        RECT 92.100 577.950 99.900 579.300 ;
        RECT 110.100 579.300 111.900 584.400 ;
        RECT 113.100 580.200 114.900 585.000 ;
        RECT 116.100 579.300 117.900 584.400 ;
        RECT 110.100 577.950 117.900 579.300 ;
        RECT 119.100 578.400 120.900 584.400 ;
        RECT 119.100 576.300 120.300 578.400 ;
        RECT 131.700 577.200 133.500 584.400 ;
        RECT 136.800 578.400 138.600 585.000 ;
        RECT 149.100 578.400 150.900 584.400 ;
        RECT 131.700 576.300 135.900 577.200 ;
        RECT 89.700 575.400 93.300 576.300 ;
        RECT 71.100 571.050 72.900 572.850 ;
        RECT 74.700 571.050 75.900 575.400 ;
        RECT 79.950 573.450 84.000 574.050 ;
        RECT 77.100 571.050 78.900 572.850 ;
        RECT 79.950 571.950 84.450 573.450 ;
        RECT 10.950 568.950 13.050 571.050 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 568.950 34.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 67.950 568.950 70.050 571.050 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 14.700 555.600 15.900 568.950 ;
        RECT 29.100 567.150 30.900 568.950 ;
        RECT 35.700 561.600 36.900 568.950 ;
        RECT 53.100 567.150 54.900 568.950 ;
        RECT 11.100 549.000 12.900 555.600 ;
        RECT 14.100 549.600 15.900 555.600 ;
        RECT 17.100 549.000 18.900 555.600 ;
        RECT 29.400 549.000 31.200 561.600 ;
        RECT 34.500 560.100 36.900 561.600 ;
        RECT 34.500 549.600 36.300 560.100 ;
        RECT 37.200 557.100 39.000 558.900 ;
        RECT 56.100 555.600 57.300 568.950 ;
        RECT 68.100 567.150 69.900 568.950 ;
        RECT 74.700 561.600 75.900 568.950 ;
        RECT 83.550 568.050 84.450 571.950 ;
        RECT 89.100 571.050 90.900 572.850 ;
        RECT 92.100 571.050 93.300 575.400 ;
        RECT 116.700 575.400 120.300 576.300 ;
        RECT 105.000 573.450 109.050 574.050 ;
        RECT 95.100 571.050 96.900 572.850 ;
        RECT 104.550 571.950 109.050 573.450 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 91.950 568.950 94.050 571.050 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 79.950 566.550 84.450 568.050 ;
        RECT 79.950 565.950 84.000 566.550 ;
        RECT 37.500 549.000 39.300 555.600 ;
        RECT 53.100 549.000 54.900 555.600 ;
        RECT 56.100 549.600 57.900 555.600 ;
        RECT 68.400 549.000 70.200 561.600 ;
        RECT 73.500 560.100 75.900 561.600 ;
        RECT 92.100 561.600 93.300 568.950 ;
        RECT 98.100 567.150 99.900 568.950 ;
        RECT 104.550 568.050 105.450 571.950 ;
        RECT 113.100 571.050 114.900 572.850 ;
        RECT 116.700 571.050 117.900 575.400 ;
        RECT 121.950 573.450 126.000 574.050 ;
        RECT 119.100 571.050 120.900 572.850 ;
        RECT 121.950 571.950 126.450 573.450 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 112.950 568.950 115.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 104.550 566.550 109.050 568.050 ;
        RECT 110.100 567.150 111.900 568.950 ;
        RECT 105.000 565.950 109.050 566.550 ;
        RECT 94.950 564.450 97.050 565.050 ;
        RECT 112.950 564.450 115.050 565.050 ;
        RECT 94.950 563.550 115.050 564.450 ;
        RECT 94.950 562.950 97.050 563.550 ;
        RECT 112.950 562.950 115.050 563.550 ;
        RECT 116.700 561.600 117.900 568.950 ;
        RECT 125.550 568.050 126.450 571.950 ;
        RECT 131.100 571.050 132.900 572.850 ;
        RECT 134.700 571.050 135.900 576.300 ;
        RECT 149.700 576.300 150.900 578.400 ;
        RECT 152.100 579.300 153.900 584.400 ;
        RECT 155.100 580.200 156.900 585.000 ;
        RECT 158.100 579.300 159.900 584.400 ;
        RECT 162.150 580.200 163.950 584.400 ;
        RECT 152.100 577.950 159.900 579.300 ;
        RECT 161.550 578.400 163.950 580.200 ;
        RECT 165.150 578.400 166.950 585.000 ;
        RECT 169.950 582.300 171.750 584.400 ;
        RECT 168.150 581.400 171.750 582.300 ;
        RECT 174.450 581.400 176.250 585.000 ;
        RECT 177.750 581.400 179.550 584.400 ;
        RECT 180.750 581.400 182.550 585.000 ;
        RECT 185.250 581.400 187.050 584.400 ;
        RECT 167.850 580.800 171.750 581.400 ;
        RECT 167.850 579.300 169.950 580.800 ;
        RECT 177.750 580.500 178.800 581.400 ;
        RECT 149.700 575.400 153.300 576.300 ;
        RECT 136.950 571.050 138.750 572.850 ;
        RECT 149.100 571.050 150.900 572.850 ;
        RECT 152.100 571.050 153.300 575.400 ;
        RECT 155.100 571.050 156.900 572.850 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 136.950 568.950 139.050 571.050 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 125.550 566.550 130.050 568.050 ;
        RECT 126.000 565.950 130.050 566.550 ;
        RECT 92.100 560.100 94.500 561.600 ;
        RECT 73.500 549.600 75.300 560.100 ;
        RECT 76.200 557.100 78.000 558.900 ;
        RECT 90.000 557.100 91.800 558.900 ;
        RECT 76.500 549.000 78.300 555.600 ;
        RECT 89.700 549.000 91.500 555.600 ;
        RECT 92.700 549.600 94.500 560.100 ;
        RECT 97.800 549.000 99.600 561.600 ;
        RECT 110.400 549.000 112.200 561.600 ;
        RECT 115.500 560.100 117.900 561.600 ;
        RECT 115.500 549.600 117.300 560.100 ;
        RECT 118.200 557.100 120.000 558.900 ;
        RECT 134.700 555.600 135.900 568.950 ;
        RECT 152.100 561.600 153.300 568.950 ;
        RECT 158.100 567.150 159.900 568.950 ;
        RECT 161.550 563.700 162.450 578.400 ;
        RECT 170.850 577.800 172.650 579.600 ;
        RECT 173.850 579.450 178.800 580.500 ;
        RECT 173.850 578.700 175.650 579.450 ;
        RECT 185.250 579.300 187.650 581.400 ;
        RECT 190.350 578.400 192.150 585.000 ;
        RECT 193.650 578.400 195.450 584.400 ;
        RECT 170.850 576.000 171.900 577.800 ;
        RECT 181.050 576.000 182.850 576.600 ;
        RECT 170.850 574.800 182.850 576.000 ;
        RECT 163.950 573.600 171.900 574.800 ;
        RECT 163.950 571.050 165.750 573.600 ;
        RECT 170.100 573.000 171.900 573.600 ;
        RECT 167.100 571.800 168.900 572.400 ;
        RECT 163.950 568.950 166.050 571.050 ;
        RECT 167.100 570.600 175.200 571.800 ;
        RECT 173.100 568.950 175.200 570.600 ;
        RECT 171.450 563.700 173.250 564.000 ;
        RECT 161.550 563.100 173.250 563.700 ;
        RECT 161.550 562.500 179.850 563.100 ;
        RECT 161.550 561.600 162.450 562.500 ;
        RECT 171.450 562.200 179.850 562.500 ;
        RECT 152.100 560.100 154.500 561.600 ;
        RECT 150.000 557.100 151.800 558.900 ;
        RECT 118.500 549.000 120.300 555.600 ;
        RECT 131.100 549.000 132.900 555.600 ;
        RECT 134.100 549.600 135.900 555.600 ;
        RECT 137.100 549.000 138.900 555.600 ;
        RECT 149.700 549.000 151.500 555.600 ;
        RECT 152.700 549.600 154.500 560.100 ;
        RECT 157.800 549.000 159.600 561.600 ;
        RECT 161.550 559.800 163.950 561.600 ;
        RECT 162.150 549.600 163.950 559.800 ;
        RECT 165.150 549.000 166.950 561.600 ;
        RECT 176.250 560.700 178.050 561.300 ;
        RECT 170.250 559.500 178.050 560.700 ;
        RECT 178.950 560.100 179.850 562.200 ;
        RECT 181.950 562.200 182.850 574.800 ;
        RECT 194.250 571.050 195.450 578.400 ;
        RECT 206.100 579.300 207.900 584.400 ;
        RECT 209.100 580.200 210.900 585.000 ;
        RECT 212.100 579.300 213.900 584.400 ;
        RECT 206.100 577.950 213.900 579.300 ;
        RECT 215.100 578.400 216.900 584.400 ;
        RECT 215.100 576.300 216.300 578.400 ;
        RECT 227.700 577.200 229.500 584.400 ;
        RECT 232.800 578.400 234.600 585.000 ;
        RECT 248.100 578.400 249.900 584.400 ;
        RECT 251.100 578.400 252.900 585.000 ;
        RECT 254.100 581.400 255.900 584.400 ;
        RECT 227.700 576.300 231.900 577.200 ;
        RECT 212.700 575.400 216.300 576.300 ;
        RECT 196.950 573.450 199.050 574.050 ;
        RECT 202.950 573.450 205.050 574.050 ;
        RECT 196.950 572.550 205.050 573.450 ;
        RECT 196.950 571.950 199.050 572.550 ;
        RECT 202.950 571.950 205.050 572.550 ;
        RECT 209.100 571.050 210.900 572.850 ;
        RECT 212.700 571.050 213.900 575.400 ;
        RECT 217.950 573.450 222.000 574.050 ;
        RECT 215.100 571.050 216.900 572.850 ;
        RECT 217.950 571.950 222.450 573.450 ;
        RECT 189.150 569.250 195.450 571.050 ;
        RECT 190.950 568.950 195.450 569.250 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 185.550 566.100 187.650 566.400 ;
        RECT 191.550 566.100 193.350 566.250 ;
        RECT 185.550 564.900 193.350 566.100 ;
        RECT 185.550 564.300 187.650 564.900 ;
        RECT 191.550 564.450 193.350 564.900 ;
        RECT 181.950 561.300 186.750 562.200 ;
        RECT 194.250 561.600 195.450 568.950 ;
        RECT 206.100 567.150 207.900 568.950 ;
        RECT 212.700 561.600 213.900 568.950 ;
        RECT 221.550 568.050 222.450 571.950 ;
        RECT 227.100 571.050 228.900 572.850 ;
        RECT 230.700 571.050 231.900 576.300 ;
        RECT 232.950 576.450 235.050 577.050 ;
        RECT 244.950 576.450 247.050 577.050 ;
        RECT 232.950 575.550 247.050 576.450 ;
        RECT 232.950 574.950 235.050 575.550 ;
        RECT 244.950 574.950 247.050 575.550 ;
        RECT 232.950 571.050 234.750 572.850 ;
        RECT 248.100 571.050 249.300 578.400 ;
        RECT 254.700 577.500 255.900 581.400 ;
        RECT 266.100 579.300 267.900 584.400 ;
        RECT 269.100 580.200 270.900 585.000 ;
        RECT 272.100 579.300 273.900 584.400 ;
        RECT 266.100 577.950 273.900 579.300 ;
        RECT 275.100 578.400 276.900 584.400 ;
        RECT 289.500 578.400 291.300 585.000 ;
        RECT 294.000 578.400 295.800 584.400 ;
        RECT 298.500 578.400 300.300 585.000 ;
        RECT 311.400 578.400 313.200 585.000 ;
        RECT 250.200 576.600 255.900 577.500 ;
        RECT 250.200 575.700 252.000 576.600 ;
        RECT 275.100 576.300 276.300 578.400 ;
        RECT 226.950 568.950 229.050 571.050 ;
        RECT 229.950 568.950 232.050 571.050 ;
        RECT 232.950 568.950 235.050 571.050 ;
        RECT 248.100 568.950 250.200 571.050 ;
        RECT 217.950 566.550 222.450 568.050 ;
        RECT 217.950 565.950 222.000 566.550 ;
        RECT 185.550 560.400 186.750 561.300 ;
        RECT 182.850 560.100 184.650 560.400 ;
        RECT 170.250 558.600 172.350 559.500 ;
        RECT 178.950 559.200 184.650 560.100 ;
        RECT 182.850 558.600 184.650 559.200 ;
        RECT 185.550 558.600 188.550 560.400 ;
        RECT 170.550 549.600 172.350 558.600 ;
        RECT 174.450 557.550 176.250 558.300 ;
        RECT 179.250 557.550 181.050 558.300 ;
        RECT 174.450 556.500 181.050 557.550 ;
        RECT 175.350 549.000 177.150 555.600 ;
        RECT 178.350 549.600 180.150 556.500 ;
        RECT 185.550 555.600 187.650 557.700 ;
        RECT 181.350 549.000 183.150 555.600 ;
        RECT 185.850 549.600 187.650 555.600 ;
        RECT 190.650 549.000 192.450 561.600 ;
        RECT 193.650 549.600 195.450 561.600 ;
        RECT 206.400 549.000 208.200 561.600 ;
        RECT 211.500 560.100 213.900 561.600 ;
        RECT 211.500 549.600 213.300 560.100 ;
        RECT 214.200 557.100 216.000 558.900 ;
        RECT 230.700 555.600 231.900 568.950 ;
        RECT 248.100 561.600 249.300 568.950 ;
        RECT 251.100 564.300 252.000 575.700 ;
        RECT 272.700 575.400 276.300 576.300 ;
        RECT 269.100 571.050 270.900 572.850 ;
        RECT 272.700 571.050 273.900 575.400 ;
        RECT 277.950 573.450 282.000 574.050 ;
        RECT 275.100 571.050 276.900 572.850 ;
        RECT 277.950 571.950 282.450 573.450 ;
        RECT 253.500 568.950 255.600 571.050 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 253.800 567.150 255.600 568.950 ;
        RECT 266.100 567.150 267.900 568.950 ;
        RECT 250.200 563.400 252.000 564.300 ;
        RECT 250.200 562.500 255.900 563.400 ;
        RECT 214.500 549.000 216.300 555.600 ;
        RECT 227.100 549.000 228.900 555.600 ;
        RECT 230.100 549.600 231.900 555.600 ;
        RECT 233.100 549.000 234.900 555.600 ;
        RECT 248.100 549.600 249.900 561.600 ;
        RECT 251.100 549.000 252.900 559.800 ;
        RECT 254.700 555.600 255.900 562.500 ;
        RECT 272.700 561.600 273.900 568.950 ;
        RECT 281.550 568.050 282.450 571.950 ;
        RECT 287.100 571.050 288.900 572.850 ;
        RECT 293.700 571.050 294.900 578.400 ;
        RECT 316.500 577.200 318.300 584.400 ;
        RECT 329.100 579.300 330.900 584.400 ;
        RECT 332.100 580.200 333.900 585.000 ;
        RECT 335.100 579.300 336.900 584.400 ;
        RECT 329.100 577.950 336.900 579.300 ;
        RECT 338.100 578.400 339.900 584.400 ;
        RECT 350.400 578.400 352.200 585.000 ;
        RECT 314.100 576.300 318.300 577.200 ;
        RECT 338.100 576.300 339.300 578.400 ;
        RECT 355.500 577.200 357.300 584.400 ;
        RECT 306.000 573.450 310.050 574.050 ;
        RECT 298.950 571.050 300.750 572.850 ;
        RECT 305.550 571.950 310.050 573.450 ;
        RECT 286.950 568.950 289.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 292.950 568.950 295.050 571.050 ;
        RECT 295.950 568.950 298.050 571.050 ;
        RECT 298.950 568.950 301.050 571.050 ;
        RECT 281.550 566.550 286.050 568.050 ;
        RECT 290.100 567.150 291.900 568.950 ;
        RECT 282.000 565.950 286.050 566.550 ;
        RECT 294.000 563.400 294.900 568.950 ;
        RECT 295.950 567.150 297.750 568.950 ;
        RECT 305.550 567.450 306.450 571.950 ;
        RECT 311.250 571.050 313.050 572.850 ;
        RECT 314.100 571.050 315.300 576.300 ;
        RECT 335.700 575.400 339.300 576.300 ;
        RECT 340.950 576.450 343.050 577.050 ;
        RECT 349.950 576.450 352.050 577.050 ;
        RECT 340.950 575.550 352.050 576.450 ;
        RECT 317.100 571.050 318.900 572.850 ;
        RECT 332.100 571.050 333.900 572.850 ;
        RECT 335.700 571.050 336.900 575.400 ;
        RECT 340.950 574.950 343.050 575.550 ;
        RECT 349.950 574.950 352.050 575.550 ;
        RECT 353.100 576.300 357.300 577.200 ;
        RECT 368.100 581.400 369.900 584.400 ;
        RECT 368.100 577.500 369.300 581.400 ;
        RECT 371.100 578.400 372.900 585.000 ;
        RECT 374.100 578.400 375.900 584.400 ;
        RECT 368.100 576.600 373.800 577.500 ;
        RECT 338.100 571.050 339.900 572.850 ;
        RECT 350.250 571.050 352.050 572.850 ;
        RECT 353.100 571.050 354.300 576.300 ;
        RECT 372.000 575.700 373.800 576.600 ;
        RECT 356.100 571.050 357.900 572.850 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 349.950 568.950 352.050 571.050 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 355.950 568.950 358.050 571.050 ;
        RECT 368.400 568.950 370.500 571.050 ;
        RECT 302.550 567.000 306.450 567.450 ;
        RECT 290.100 562.500 294.900 563.400 ;
        RECT 301.950 566.550 306.450 567.000 ;
        RECT 301.950 562.950 304.050 566.550 ;
        RECT 254.100 549.600 255.900 555.600 ;
        RECT 266.400 549.000 268.200 561.600 ;
        RECT 271.500 560.100 273.900 561.600 ;
        RECT 271.500 549.600 273.300 560.100 ;
        RECT 274.200 557.100 276.000 558.900 ;
        RECT 274.500 549.000 276.300 555.600 ;
        RECT 287.100 550.500 288.900 561.600 ;
        RECT 290.100 551.400 291.900 562.500 ;
        RECT 293.100 560.400 300.900 561.300 ;
        RECT 293.100 550.500 294.900 560.400 ;
        RECT 287.100 549.600 294.900 550.500 ;
        RECT 296.100 549.000 297.900 559.500 ;
        RECT 299.100 549.600 300.900 560.400 ;
        RECT 314.100 555.600 315.300 568.950 ;
        RECT 329.100 567.150 330.900 568.950 ;
        RECT 335.700 561.600 336.900 568.950 ;
        RECT 311.100 549.000 312.900 555.600 ;
        RECT 314.100 549.600 315.900 555.600 ;
        RECT 317.100 549.000 318.900 555.600 ;
        RECT 329.400 549.000 331.200 561.600 ;
        RECT 334.500 560.100 336.900 561.600 ;
        RECT 334.500 549.600 336.300 560.100 ;
        RECT 337.200 557.100 339.000 558.900 ;
        RECT 353.100 555.600 354.300 568.950 ;
        RECT 368.400 567.150 370.200 568.950 ;
        RECT 372.000 564.300 372.900 575.700 ;
        RECT 374.700 571.050 375.900 578.400 ;
        RECT 373.800 568.950 375.900 571.050 ;
        RECT 372.000 563.400 373.800 564.300 ;
        RECT 368.100 562.500 373.800 563.400 ;
        RECT 368.100 555.600 369.300 562.500 ;
        RECT 374.700 561.600 375.900 568.950 ;
        RECT 337.500 549.000 339.300 555.600 ;
        RECT 350.100 549.000 351.900 555.600 ;
        RECT 353.100 549.600 354.900 555.600 ;
        RECT 356.100 549.000 357.900 555.600 ;
        RECT 368.100 549.600 369.900 555.600 ;
        RECT 371.100 549.000 372.900 559.800 ;
        RECT 374.100 549.600 375.900 561.600 ;
        RECT 377.550 578.400 379.350 584.400 ;
        RECT 380.850 578.400 382.650 585.000 ;
        RECT 385.950 581.400 387.750 584.400 ;
        RECT 390.450 581.400 392.250 585.000 ;
        RECT 393.450 581.400 395.250 584.400 ;
        RECT 396.750 581.400 398.550 585.000 ;
        RECT 401.250 582.300 403.050 584.400 ;
        RECT 401.250 581.400 404.850 582.300 ;
        RECT 385.350 579.300 387.750 581.400 ;
        RECT 394.200 580.500 395.250 581.400 ;
        RECT 401.250 580.800 405.150 581.400 ;
        RECT 394.200 579.450 399.150 580.500 ;
        RECT 397.350 578.700 399.150 579.450 ;
        RECT 377.550 571.050 378.750 578.400 ;
        RECT 400.350 577.800 402.150 579.600 ;
        RECT 403.050 579.300 405.150 580.800 ;
        RECT 406.050 578.400 407.850 585.000 ;
        RECT 409.050 580.200 410.850 584.400 ;
        RECT 414.150 580.200 415.950 584.400 ;
        RECT 409.050 578.400 411.450 580.200 ;
        RECT 390.150 576.000 391.950 576.600 ;
        RECT 401.100 576.000 402.150 577.800 ;
        RECT 390.150 574.800 402.150 576.000 ;
        RECT 377.550 569.250 383.850 571.050 ;
        RECT 377.550 568.950 382.050 569.250 ;
        RECT 377.550 561.600 378.750 568.950 ;
        RECT 379.650 566.100 381.450 566.250 ;
        RECT 385.350 566.100 387.450 566.400 ;
        RECT 379.650 564.900 387.450 566.100 ;
        RECT 379.650 564.450 381.450 564.900 ;
        RECT 385.350 564.300 387.450 564.900 ;
        RECT 390.150 562.200 391.050 574.800 ;
        RECT 401.100 573.600 409.050 574.800 ;
        RECT 401.100 573.000 402.900 573.600 ;
        RECT 404.100 571.800 405.900 572.400 ;
        RECT 397.800 570.600 405.900 571.800 ;
        RECT 407.250 571.050 409.050 573.600 ;
        RECT 397.800 568.950 399.900 570.600 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 399.750 563.700 401.550 564.000 ;
        RECT 410.550 563.700 411.450 578.400 ;
        RECT 399.750 563.100 411.450 563.700 ;
        RECT 377.550 549.600 379.350 561.600 ;
        RECT 380.550 549.000 382.350 561.600 ;
        RECT 386.250 561.300 391.050 562.200 ;
        RECT 393.150 562.500 411.450 563.100 ;
        RECT 393.150 562.200 401.550 562.500 ;
        RECT 386.250 560.400 387.450 561.300 ;
        RECT 384.450 558.600 387.450 560.400 ;
        RECT 388.350 560.100 390.150 560.400 ;
        RECT 393.150 560.100 394.050 562.200 ;
        RECT 410.550 561.600 411.450 562.500 ;
        RECT 388.350 559.200 394.050 560.100 ;
        RECT 394.950 560.700 396.750 561.300 ;
        RECT 394.950 559.500 402.750 560.700 ;
        RECT 388.350 558.600 390.150 559.200 ;
        RECT 400.650 558.600 402.750 559.500 ;
        RECT 385.350 555.600 387.450 557.700 ;
        RECT 391.950 557.550 393.750 558.300 ;
        RECT 396.750 557.550 398.550 558.300 ;
        RECT 391.950 556.500 398.550 557.550 ;
        RECT 385.350 549.600 387.150 555.600 ;
        RECT 389.850 549.000 391.650 555.600 ;
        RECT 392.850 549.600 394.650 556.500 ;
        RECT 395.850 549.000 397.650 555.600 ;
        RECT 400.650 549.600 402.450 558.600 ;
        RECT 406.050 549.000 407.850 561.600 ;
        RECT 409.050 559.800 411.450 561.600 ;
        RECT 413.550 578.400 415.950 580.200 ;
        RECT 417.150 578.400 418.950 585.000 ;
        RECT 421.950 582.300 423.750 584.400 ;
        RECT 420.150 581.400 423.750 582.300 ;
        RECT 426.450 581.400 428.250 585.000 ;
        RECT 429.750 581.400 431.550 584.400 ;
        RECT 432.750 581.400 434.550 585.000 ;
        RECT 437.250 581.400 439.050 584.400 ;
        RECT 419.850 580.800 423.750 581.400 ;
        RECT 419.850 579.300 421.950 580.800 ;
        RECT 429.750 580.500 430.800 581.400 ;
        RECT 413.550 563.700 414.450 578.400 ;
        RECT 422.850 577.800 424.650 579.600 ;
        RECT 425.850 579.450 430.800 580.500 ;
        RECT 425.850 578.700 427.650 579.450 ;
        RECT 437.250 579.300 439.650 581.400 ;
        RECT 442.350 578.400 444.150 585.000 ;
        RECT 445.650 578.400 447.450 584.400 ;
        RECT 422.850 576.000 423.900 577.800 ;
        RECT 433.050 576.000 434.850 576.600 ;
        RECT 422.850 574.800 434.850 576.000 ;
        RECT 415.950 573.600 423.900 574.800 ;
        RECT 415.950 571.050 417.750 573.600 ;
        RECT 422.100 573.000 423.900 573.600 ;
        RECT 419.100 571.800 420.900 572.400 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 419.100 570.600 427.200 571.800 ;
        RECT 425.100 568.950 427.200 570.600 ;
        RECT 423.450 563.700 425.250 564.000 ;
        RECT 413.550 563.100 425.250 563.700 ;
        RECT 413.550 562.500 431.850 563.100 ;
        RECT 413.550 561.600 414.450 562.500 ;
        RECT 423.450 562.200 431.850 562.500 ;
        RECT 413.550 559.800 415.950 561.600 ;
        RECT 409.050 549.600 410.850 559.800 ;
        RECT 414.150 549.600 415.950 559.800 ;
        RECT 417.150 549.000 418.950 561.600 ;
        RECT 428.250 560.700 430.050 561.300 ;
        RECT 422.250 559.500 430.050 560.700 ;
        RECT 430.950 560.100 431.850 562.200 ;
        RECT 433.950 562.200 434.850 574.800 ;
        RECT 446.250 571.050 447.450 578.400 ;
        RECT 441.150 569.250 447.450 571.050 ;
        RECT 442.950 568.950 447.450 569.250 ;
        RECT 437.550 566.100 439.650 566.400 ;
        RECT 443.550 566.100 445.350 566.250 ;
        RECT 437.550 564.900 445.350 566.100 ;
        RECT 437.550 564.300 439.650 564.900 ;
        RECT 443.550 564.450 445.350 564.900 ;
        RECT 433.950 561.300 438.750 562.200 ;
        RECT 446.250 561.600 447.450 568.950 ;
        RECT 437.550 560.400 438.750 561.300 ;
        RECT 434.850 560.100 436.650 560.400 ;
        RECT 422.250 558.600 424.350 559.500 ;
        RECT 430.950 559.200 436.650 560.100 ;
        RECT 434.850 558.600 436.650 559.200 ;
        RECT 437.550 558.600 440.550 560.400 ;
        RECT 422.550 549.600 424.350 558.600 ;
        RECT 426.450 557.550 428.250 558.300 ;
        RECT 431.250 557.550 433.050 558.300 ;
        RECT 426.450 556.500 433.050 557.550 ;
        RECT 427.350 549.000 429.150 555.600 ;
        RECT 430.350 549.600 432.150 556.500 ;
        RECT 437.550 555.600 439.650 557.700 ;
        RECT 433.350 549.000 435.150 555.600 ;
        RECT 437.850 549.600 439.650 555.600 ;
        RECT 442.650 549.000 444.450 561.600 ;
        RECT 445.650 549.600 447.450 561.600 ;
        RECT 449.550 578.400 451.350 584.400 ;
        RECT 452.850 578.400 454.650 585.000 ;
        RECT 457.950 581.400 459.750 584.400 ;
        RECT 462.450 581.400 464.250 585.000 ;
        RECT 465.450 581.400 467.250 584.400 ;
        RECT 468.750 581.400 470.550 585.000 ;
        RECT 473.250 582.300 475.050 584.400 ;
        RECT 473.250 581.400 476.850 582.300 ;
        RECT 457.350 579.300 459.750 581.400 ;
        RECT 466.200 580.500 467.250 581.400 ;
        RECT 473.250 580.800 477.150 581.400 ;
        RECT 466.200 579.450 471.150 580.500 ;
        RECT 469.350 578.700 471.150 579.450 ;
        RECT 449.550 571.050 450.750 578.400 ;
        RECT 472.350 577.800 474.150 579.600 ;
        RECT 475.050 579.300 477.150 580.800 ;
        RECT 478.050 578.400 479.850 585.000 ;
        RECT 481.050 580.200 482.850 584.400 ;
        RECT 494.100 581.400 495.900 584.400 ;
        RECT 481.050 578.400 483.450 580.200 ;
        RECT 462.150 576.000 463.950 576.600 ;
        RECT 473.100 576.000 474.150 577.800 ;
        RECT 462.150 574.800 474.150 576.000 ;
        RECT 449.550 569.250 455.850 571.050 ;
        RECT 449.550 568.950 454.050 569.250 ;
        RECT 449.550 561.600 450.750 568.950 ;
        RECT 451.650 566.100 453.450 566.250 ;
        RECT 457.350 566.100 459.450 566.400 ;
        RECT 451.650 564.900 459.450 566.100 ;
        RECT 451.650 564.450 453.450 564.900 ;
        RECT 457.350 564.300 459.450 564.900 ;
        RECT 462.150 562.200 463.050 574.800 ;
        RECT 473.100 573.600 481.050 574.800 ;
        RECT 473.100 573.000 474.900 573.600 ;
        RECT 476.100 571.800 477.900 572.400 ;
        RECT 469.800 570.600 477.900 571.800 ;
        RECT 479.250 571.050 481.050 573.600 ;
        RECT 469.800 568.950 471.900 570.600 ;
        RECT 478.950 568.950 481.050 571.050 ;
        RECT 471.750 563.700 473.550 564.000 ;
        RECT 482.550 563.700 483.450 578.400 ;
        RECT 494.100 577.500 495.300 581.400 ;
        RECT 497.100 578.400 498.900 585.000 ;
        RECT 500.100 578.400 501.900 584.400 ;
        RECT 494.100 576.600 499.800 577.500 ;
        RECT 498.000 575.700 499.800 576.600 ;
        RECT 494.400 568.950 496.500 571.050 ;
        RECT 494.400 567.150 496.200 568.950 ;
        RECT 471.750 563.100 483.450 563.700 ;
        RECT 498.000 564.300 498.900 575.700 ;
        RECT 500.700 571.050 501.900 578.400 ;
        RECT 512.700 577.200 514.500 584.400 ;
        RECT 517.800 578.400 519.600 585.000 ;
        RECT 521.550 578.400 523.350 584.400 ;
        RECT 524.850 578.400 526.650 585.000 ;
        RECT 529.950 581.400 531.750 584.400 ;
        RECT 534.450 581.400 536.250 585.000 ;
        RECT 537.450 581.400 539.250 584.400 ;
        RECT 540.750 581.400 542.550 585.000 ;
        RECT 545.250 582.300 547.050 584.400 ;
        RECT 545.250 581.400 548.850 582.300 ;
        RECT 529.350 579.300 531.750 581.400 ;
        RECT 538.200 580.500 539.250 581.400 ;
        RECT 545.250 580.800 549.150 581.400 ;
        RECT 538.200 579.450 543.150 580.500 ;
        RECT 541.350 578.700 543.150 579.450 ;
        RECT 512.700 576.300 516.900 577.200 ;
        RECT 512.100 571.050 513.900 572.850 ;
        RECT 515.700 571.050 516.900 576.300 ;
        RECT 517.950 571.050 519.750 572.850 ;
        RECT 521.550 571.050 522.750 578.400 ;
        RECT 544.350 577.800 546.150 579.600 ;
        RECT 547.050 579.300 549.150 580.800 ;
        RECT 550.050 578.400 551.850 585.000 ;
        RECT 553.050 580.200 554.850 584.400 ;
        RECT 553.050 578.400 555.450 580.200 ;
        RECT 566.100 578.400 567.900 584.400 ;
        RECT 534.150 576.000 535.950 576.600 ;
        RECT 545.100 576.000 546.150 577.800 ;
        RECT 534.150 574.800 546.150 576.000 ;
        RECT 499.800 568.950 501.900 571.050 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 517.950 568.950 520.050 571.050 ;
        RECT 521.550 569.250 527.850 571.050 ;
        RECT 521.550 568.950 526.050 569.250 ;
        RECT 498.000 563.400 499.800 564.300 ;
        RECT 449.550 549.600 451.350 561.600 ;
        RECT 452.550 549.000 454.350 561.600 ;
        RECT 458.250 561.300 463.050 562.200 ;
        RECT 465.150 562.500 483.450 563.100 ;
        RECT 465.150 562.200 473.550 562.500 ;
        RECT 458.250 560.400 459.450 561.300 ;
        RECT 456.450 558.600 459.450 560.400 ;
        RECT 460.350 560.100 462.150 560.400 ;
        RECT 465.150 560.100 466.050 562.200 ;
        RECT 482.550 561.600 483.450 562.500 ;
        RECT 460.350 559.200 466.050 560.100 ;
        RECT 466.950 560.700 468.750 561.300 ;
        RECT 466.950 559.500 474.750 560.700 ;
        RECT 460.350 558.600 462.150 559.200 ;
        RECT 472.650 558.600 474.750 559.500 ;
        RECT 457.350 555.600 459.450 557.700 ;
        RECT 463.950 557.550 465.750 558.300 ;
        RECT 468.750 557.550 470.550 558.300 ;
        RECT 463.950 556.500 470.550 557.550 ;
        RECT 457.350 549.600 459.150 555.600 ;
        RECT 461.850 549.000 463.650 555.600 ;
        RECT 464.850 549.600 466.650 556.500 ;
        RECT 467.850 549.000 469.650 555.600 ;
        RECT 472.650 549.600 474.450 558.600 ;
        RECT 478.050 549.000 479.850 561.600 ;
        RECT 481.050 559.800 483.450 561.600 ;
        RECT 494.100 562.500 499.800 563.400 ;
        RECT 481.050 549.600 482.850 559.800 ;
        RECT 494.100 555.600 495.300 562.500 ;
        RECT 500.700 561.600 501.900 568.950 ;
        RECT 494.100 549.600 495.900 555.600 ;
        RECT 497.100 549.000 498.900 559.800 ;
        RECT 500.100 549.600 501.900 561.600 ;
        RECT 515.700 555.600 516.900 568.950 ;
        RECT 521.550 561.600 522.750 568.950 ;
        RECT 523.650 566.100 525.450 566.250 ;
        RECT 529.350 566.100 531.450 566.400 ;
        RECT 523.650 564.900 531.450 566.100 ;
        RECT 523.650 564.450 525.450 564.900 ;
        RECT 529.350 564.300 531.450 564.900 ;
        RECT 534.150 562.200 535.050 574.800 ;
        RECT 545.100 573.600 553.050 574.800 ;
        RECT 545.100 573.000 546.900 573.600 ;
        RECT 548.100 571.800 549.900 572.400 ;
        RECT 541.800 570.600 549.900 571.800 ;
        RECT 551.250 571.050 553.050 573.600 ;
        RECT 541.800 568.950 543.900 570.600 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 543.750 563.700 545.550 564.000 ;
        RECT 554.550 563.700 555.450 578.400 ;
        RECT 566.700 576.300 567.900 578.400 ;
        RECT 569.100 579.300 570.900 584.400 ;
        RECT 572.100 580.200 573.900 585.000 ;
        RECT 575.100 579.300 576.900 584.400 ;
        RECT 569.100 577.950 576.900 579.300 ;
        RECT 587.100 579.300 588.900 584.400 ;
        RECT 590.100 580.200 591.900 585.000 ;
        RECT 593.100 579.300 594.900 584.400 ;
        RECT 587.100 577.950 594.900 579.300 ;
        RECT 596.100 578.400 597.900 584.400 ;
        RECT 599.550 578.400 601.350 584.400 ;
        RECT 602.850 578.400 604.650 585.000 ;
        RECT 607.950 581.400 609.750 584.400 ;
        RECT 612.450 581.400 614.250 585.000 ;
        RECT 615.450 581.400 617.250 584.400 ;
        RECT 618.750 581.400 620.550 585.000 ;
        RECT 623.250 582.300 625.050 584.400 ;
        RECT 623.250 581.400 626.850 582.300 ;
        RECT 607.350 579.300 609.750 581.400 ;
        RECT 616.200 580.500 617.250 581.400 ;
        RECT 623.250 580.800 627.150 581.400 ;
        RECT 616.200 579.450 621.150 580.500 ;
        RECT 619.350 578.700 621.150 579.450 ;
        RECT 596.100 576.300 597.300 578.400 ;
        RECT 566.700 575.400 570.300 576.300 ;
        RECT 566.100 571.050 567.900 572.850 ;
        RECT 569.100 571.050 570.300 575.400 ;
        RECT 593.700 575.400 597.300 576.300 ;
        RECT 582.000 573.450 586.050 574.050 ;
        RECT 572.100 571.050 573.900 572.850 ;
        RECT 581.550 571.950 586.050 573.450 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 543.750 563.100 555.450 563.700 ;
        RECT 512.100 549.000 513.900 555.600 ;
        RECT 515.100 549.600 516.900 555.600 ;
        RECT 518.100 549.000 519.900 555.600 ;
        RECT 521.550 549.600 523.350 561.600 ;
        RECT 524.550 549.000 526.350 561.600 ;
        RECT 530.250 561.300 535.050 562.200 ;
        RECT 537.150 562.500 555.450 563.100 ;
        RECT 537.150 562.200 545.550 562.500 ;
        RECT 530.250 560.400 531.450 561.300 ;
        RECT 528.450 558.600 531.450 560.400 ;
        RECT 532.350 560.100 534.150 560.400 ;
        RECT 537.150 560.100 538.050 562.200 ;
        RECT 554.550 561.600 555.450 562.500 ;
        RECT 532.350 559.200 538.050 560.100 ;
        RECT 538.950 560.700 540.750 561.300 ;
        RECT 538.950 559.500 546.750 560.700 ;
        RECT 532.350 558.600 534.150 559.200 ;
        RECT 544.650 558.600 546.750 559.500 ;
        RECT 529.350 555.600 531.450 557.700 ;
        RECT 535.950 557.550 537.750 558.300 ;
        RECT 540.750 557.550 542.550 558.300 ;
        RECT 535.950 556.500 542.550 557.550 ;
        RECT 529.350 549.600 531.150 555.600 ;
        RECT 533.850 549.000 535.650 555.600 ;
        RECT 536.850 549.600 538.650 556.500 ;
        RECT 539.850 549.000 541.650 555.600 ;
        RECT 544.650 549.600 546.450 558.600 ;
        RECT 550.050 549.000 551.850 561.600 ;
        RECT 553.050 559.800 555.450 561.600 ;
        RECT 569.100 561.600 570.300 568.950 ;
        RECT 575.100 567.150 576.900 568.950 ;
        RECT 581.550 568.050 582.450 571.950 ;
        RECT 590.100 571.050 591.900 572.850 ;
        RECT 593.700 571.050 594.900 575.400 ;
        RECT 596.100 571.050 597.900 572.850 ;
        RECT 599.550 571.050 600.750 578.400 ;
        RECT 622.350 577.800 624.150 579.600 ;
        RECT 625.050 579.300 627.150 580.800 ;
        RECT 628.050 578.400 629.850 585.000 ;
        RECT 631.050 580.200 632.850 584.400 ;
        RECT 631.050 578.400 633.450 580.200 ;
        RECT 644.100 578.400 645.900 585.000 ;
        RECT 612.150 576.000 613.950 576.600 ;
        RECT 623.100 576.000 624.150 577.800 ;
        RECT 612.150 574.800 624.150 576.000 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 595.950 568.950 598.050 571.050 ;
        RECT 599.550 569.250 605.850 571.050 ;
        RECT 599.550 568.950 604.050 569.250 ;
        RECT 581.550 566.550 586.050 568.050 ;
        RECT 587.100 567.150 588.900 568.950 ;
        RECT 582.000 565.950 586.050 566.550 ;
        RECT 593.700 561.600 594.900 568.950 ;
        RECT 569.100 560.100 571.500 561.600 ;
        RECT 553.050 549.600 554.850 559.800 ;
        RECT 567.000 557.100 568.800 558.900 ;
        RECT 566.700 549.000 568.500 555.600 ;
        RECT 569.700 549.600 571.500 560.100 ;
        RECT 574.800 549.000 576.600 561.600 ;
        RECT 587.400 549.000 589.200 561.600 ;
        RECT 592.500 560.100 594.900 561.600 ;
        RECT 599.550 561.600 600.750 568.950 ;
        RECT 601.650 566.100 603.450 566.250 ;
        RECT 607.350 566.100 609.450 566.400 ;
        RECT 601.650 564.900 609.450 566.100 ;
        RECT 601.650 564.450 603.450 564.900 ;
        RECT 607.350 564.300 609.450 564.900 ;
        RECT 612.150 562.200 613.050 574.800 ;
        RECT 623.100 573.600 631.050 574.800 ;
        RECT 623.100 573.000 624.900 573.600 ;
        RECT 626.100 571.800 627.900 572.400 ;
        RECT 619.800 570.600 627.900 571.800 ;
        RECT 629.250 571.050 631.050 573.600 ;
        RECT 619.800 568.950 621.900 570.600 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 621.750 563.700 623.550 564.000 ;
        RECT 632.550 563.700 633.450 578.400 ;
        RECT 647.100 577.500 648.900 584.400 ;
        RECT 650.100 578.400 651.900 585.000 ;
        RECT 653.100 577.500 654.900 584.400 ;
        RECT 656.100 578.400 657.900 585.000 ;
        RECT 659.100 577.500 660.900 584.400 ;
        RECT 662.100 578.400 663.900 585.000 ;
        RECT 665.100 577.500 666.900 584.400 ;
        RECT 668.100 578.400 669.900 585.000 ;
        RECT 680.100 581.400 681.900 584.400 ;
        RECT 680.100 577.500 681.300 581.400 ;
        RECT 683.100 578.400 684.900 585.000 ;
        RECT 686.100 578.400 687.900 584.400 ;
        RECT 647.100 576.300 651.000 577.500 ;
        RECT 653.100 576.300 657.000 577.500 ;
        RECT 659.100 576.300 663.000 577.500 ;
        RECT 665.100 576.300 667.950 577.500 ;
        RECT 680.100 576.600 685.800 577.500 ;
        RECT 649.800 575.400 651.000 576.300 ;
        RECT 655.800 575.400 657.000 576.300 ;
        RECT 661.800 575.400 663.000 576.300 ;
        RECT 649.800 574.200 654.000 575.400 ;
        RECT 646.800 571.050 648.600 572.850 ;
        RECT 646.800 568.950 648.900 571.050 ;
        RECT 649.800 563.700 651.000 574.200 ;
        RECT 652.200 573.600 654.000 574.200 ;
        RECT 655.800 574.200 660.000 575.400 ;
        RECT 655.800 563.700 657.000 574.200 ;
        RECT 658.200 573.600 660.000 574.200 ;
        RECT 661.800 574.200 666.000 575.400 ;
        RECT 661.800 563.700 663.000 574.200 ;
        RECT 664.200 573.600 666.000 574.200 ;
        RECT 666.900 571.050 667.950 576.300 ;
        RECT 684.000 575.700 685.800 576.600 ;
        RECT 664.800 568.950 667.950 571.050 ;
        RECT 666.900 563.700 667.950 568.950 ;
        RECT 680.400 568.950 682.500 571.050 ;
        RECT 680.400 567.150 682.200 568.950 ;
        RECT 621.750 563.100 633.450 563.700 ;
        RECT 592.500 549.600 594.300 560.100 ;
        RECT 595.200 557.100 597.000 558.900 ;
        RECT 595.500 549.000 597.300 555.600 ;
        RECT 599.550 549.600 601.350 561.600 ;
        RECT 602.550 549.000 604.350 561.600 ;
        RECT 608.250 561.300 613.050 562.200 ;
        RECT 615.150 562.500 633.450 563.100 ;
        RECT 615.150 562.200 623.550 562.500 ;
        RECT 608.250 560.400 609.450 561.300 ;
        RECT 606.450 558.600 609.450 560.400 ;
        RECT 610.350 560.100 612.150 560.400 ;
        RECT 615.150 560.100 616.050 562.200 ;
        RECT 632.550 561.600 633.450 562.500 ;
        RECT 647.100 562.500 651.000 563.700 ;
        RECT 653.100 562.500 657.000 563.700 ;
        RECT 659.100 562.500 663.000 563.700 ;
        RECT 665.100 562.500 667.950 563.700 ;
        RECT 684.000 564.300 684.900 575.700 ;
        RECT 686.700 571.050 687.900 578.400 ;
        RECT 698.100 579.300 699.900 584.400 ;
        RECT 701.100 580.200 702.900 585.000 ;
        RECT 704.100 579.300 705.900 584.400 ;
        RECT 698.100 577.950 705.900 579.300 ;
        RECT 707.100 578.400 708.900 584.400 ;
        RECT 707.100 576.300 708.300 578.400 ;
        RECT 719.700 577.200 721.500 584.400 ;
        RECT 724.800 578.400 726.600 585.000 ;
        RECT 729.150 580.200 730.950 584.400 ;
        RECT 728.550 578.400 730.950 580.200 ;
        RECT 732.150 578.400 733.950 585.000 ;
        RECT 736.950 582.300 738.750 584.400 ;
        RECT 735.150 581.400 738.750 582.300 ;
        RECT 741.450 581.400 743.250 585.000 ;
        RECT 744.750 581.400 746.550 584.400 ;
        RECT 747.750 581.400 749.550 585.000 ;
        RECT 752.250 581.400 754.050 584.400 ;
        RECT 734.850 580.800 738.750 581.400 ;
        RECT 734.850 579.300 736.950 580.800 ;
        RECT 744.750 580.500 745.800 581.400 ;
        RECT 719.700 576.300 723.900 577.200 ;
        RECT 704.700 575.400 708.300 576.300 ;
        RECT 701.100 571.050 702.900 572.850 ;
        RECT 704.700 571.050 705.900 575.400 ;
        RECT 707.100 571.050 708.900 572.850 ;
        RECT 719.100 571.050 720.900 572.850 ;
        RECT 722.700 571.050 723.900 576.300 ;
        RECT 724.950 571.050 726.750 572.850 ;
        RECT 685.800 568.950 687.900 571.050 ;
        RECT 684.000 563.400 685.800 564.300 ;
        RECT 680.100 562.500 685.800 563.400 ;
        RECT 610.350 559.200 616.050 560.100 ;
        RECT 616.950 560.700 618.750 561.300 ;
        RECT 616.950 559.500 624.750 560.700 ;
        RECT 610.350 558.600 612.150 559.200 ;
        RECT 622.650 558.600 624.750 559.500 ;
        RECT 607.350 555.600 609.450 557.700 ;
        RECT 613.950 557.550 615.750 558.300 ;
        RECT 618.750 557.550 620.550 558.300 ;
        RECT 613.950 556.500 620.550 557.550 ;
        RECT 607.350 549.600 609.150 555.600 ;
        RECT 611.850 549.000 613.650 555.600 ;
        RECT 614.850 549.600 616.650 556.500 ;
        RECT 617.850 549.000 619.650 555.600 ;
        RECT 622.650 549.600 624.450 558.600 ;
        RECT 628.050 549.000 629.850 561.600 ;
        RECT 631.050 559.800 633.450 561.600 ;
        RECT 631.050 549.600 632.850 559.800 ;
        RECT 644.100 549.000 645.900 561.600 ;
        RECT 647.100 549.600 648.900 562.500 ;
        RECT 650.100 549.000 651.900 561.600 ;
        RECT 653.100 549.600 654.900 562.500 ;
        RECT 656.100 549.000 657.900 561.600 ;
        RECT 659.100 549.600 660.900 562.500 ;
        RECT 662.100 549.000 663.900 561.600 ;
        RECT 665.100 549.600 666.900 562.500 ;
        RECT 668.100 549.000 669.900 561.600 ;
        RECT 680.100 555.600 681.300 562.500 ;
        RECT 686.700 561.600 687.900 568.950 ;
        RECT 691.950 568.050 694.050 571.050 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 718.950 568.950 721.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 691.950 567.000 697.050 568.050 ;
        RECT 698.100 567.150 699.900 568.950 ;
        RECT 692.550 566.550 697.050 567.000 ;
        RECT 693.000 565.950 697.050 566.550 ;
        RECT 704.700 561.600 705.900 568.950 ;
        RECT 680.100 549.600 681.900 555.600 ;
        RECT 683.100 549.000 684.900 559.800 ;
        RECT 686.100 549.600 687.900 561.600 ;
        RECT 698.400 549.000 700.200 561.600 ;
        RECT 703.500 560.100 705.900 561.600 ;
        RECT 703.500 549.600 705.300 560.100 ;
        RECT 706.200 557.100 708.000 558.900 ;
        RECT 722.700 555.600 723.900 568.950 ;
        RECT 728.550 563.700 729.450 578.400 ;
        RECT 737.850 577.800 739.650 579.600 ;
        RECT 740.850 579.450 745.800 580.500 ;
        RECT 740.850 578.700 742.650 579.450 ;
        RECT 752.250 579.300 754.650 581.400 ;
        RECT 757.350 578.400 759.150 585.000 ;
        RECT 760.650 578.400 762.450 584.400 ;
        RECT 737.850 576.000 738.900 577.800 ;
        RECT 748.050 576.000 749.850 576.600 ;
        RECT 737.850 574.800 749.850 576.000 ;
        RECT 730.950 573.600 738.900 574.800 ;
        RECT 730.950 571.050 732.750 573.600 ;
        RECT 737.100 573.000 738.900 573.600 ;
        RECT 734.100 571.800 735.900 572.400 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 734.100 570.600 742.200 571.800 ;
        RECT 740.100 568.950 742.200 570.600 ;
        RECT 738.450 563.700 740.250 564.000 ;
        RECT 728.550 563.100 740.250 563.700 ;
        RECT 728.550 562.500 746.850 563.100 ;
        RECT 728.550 561.600 729.450 562.500 ;
        RECT 738.450 562.200 746.850 562.500 ;
        RECT 728.550 559.800 730.950 561.600 ;
        RECT 706.500 549.000 708.300 555.600 ;
        RECT 719.100 549.000 720.900 555.600 ;
        RECT 722.100 549.600 723.900 555.600 ;
        RECT 725.100 549.000 726.900 555.600 ;
        RECT 729.150 549.600 730.950 559.800 ;
        RECT 732.150 549.000 733.950 561.600 ;
        RECT 743.250 560.700 745.050 561.300 ;
        RECT 737.250 559.500 745.050 560.700 ;
        RECT 745.950 560.100 746.850 562.200 ;
        RECT 748.950 562.200 749.850 574.800 ;
        RECT 761.250 571.050 762.450 578.400 ;
        RECT 773.100 576.600 774.900 584.400 ;
        RECT 777.600 578.400 779.400 585.000 ;
        RECT 780.600 580.200 782.400 584.400 ;
        RECT 780.600 578.400 783.300 580.200 ;
        RECT 795.000 578.400 796.800 585.000 ;
        RECT 799.500 579.600 801.300 584.400 ;
        RECT 802.500 581.400 804.300 585.000 ;
        RECT 815.100 581.400 816.900 585.000 ;
        RECT 818.100 581.400 819.900 584.400 ;
        RECT 821.100 581.400 822.900 585.000 ;
        RECT 799.500 578.400 804.600 579.600 ;
        RECT 779.700 576.600 781.500 577.500 ;
        RECT 773.100 575.700 781.500 576.600 ;
        RECT 773.250 571.050 775.050 572.850 ;
        RECT 756.150 569.250 762.450 571.050 ;
        RECT 757.950 568.950 762.450 569.250 ;
        RECT 773.100 568.950 775.200 571.050 ;
        RECT 752.550 566.100 754.650 566.400 ;
        RECT 758.550 566.100 760.350 566.250 ;
        RECT 752.550 564.900 760.350 566.100 ;
        RECT 752.550 564.300 754.650 564.900 ;
        RECT 758.550 564.450 760.350 564.900 ;
        RECT 748.950 561.300 753.750 562.200 ;
        RECT 761.250 561.600 762.450 568.950 ;
        RECT 752.550 560.400 753.750 561.300 ;
        RECT 749.850 560.100 751.650 560.400 ;
        RECT 737.250 558.600 739.350 559.500 ;
        RECT 745.950 559.200 751.650 560.100 ;
        RECT 749.850 558.600 751.650 559.200 ;
        RECT 752.550 558.600 755.550 560.400 ;
        RECT 737.550 549.600 739.350 558.600 ;
        RECT 741.450 557.550 743.250 558.300 ;
        RECT 746.250 557.550 748.050 558.300 ;
        RECT 741.450 556.500 748.050 557.550 ;
        RECT 742.350 549.000 744.150 555.600 ;
        RECT 745.350 549.600 747.150 556.500 ;
        RECT 752.550 555.600 754.650 557.700 ;
        RECT 748.350 549.000 750.150 555.600 ;
        RECT 752.850 549.600 754.650 555.600 ;
        RECT 757.650 549.000 759.450 561.600 ;
        RECT 760.650 549.600 762.450 561.600 ;
        RECT 776.100 555.600 777.000 575.700 ;
        RECT 782.400 571.050 783.300 578.400 ;
        RECT 794.100 571.050 795.900 572.850 ;
        RECT 800.250 571.050 802.050 572.850 ;
        RECT 803.700 571.050 804.600 578.400 ;
        RECT 811.950 573.450 814.050 577.050 ;
        RECT 809.550 573.000 814.050 573.450 ;
        RECT 809.550 572.550 813.450 573.000 ;
        RECT 778.500 568.950 780.600 571.050 ;
        RECT 781.800 568.950 783.900 571.050 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 778.200 567.150 780.000 568.950 ;
        RECT 782.400 561.600 783.300 568.950 ;
        RECT 797.250 567.150 799.050 568.950 ;
        RECT 803.700 561.600 804.600 568.950 ;
        RECT 809.550 568.050 810.450 572.550 ;
        RECT 818.700 571.050 819.600 581.400 ;
        RECT 836.700 577.200 838.500 584.400 ;
        RECT 841.800 578.400 843.600 585.000 ;
        RECT 836.700 576.300 840.900 577.200 ;
        RECT 836.100 571.050 837.900 572.850 ;
        RECT 839.700 571.050 840.900 576.300 ;
        RECT 854.100 575.400 855.900 585.000 ;
        RECT 860.700 576.000 862.500 584.400 ;
        RECT 860.700 574.800 864.000 576.000 ;
        RECT 841.950 571.050 843.750 572.850 ;
        RECT 854.100 571.050 855.900 572.850 ;
        RECT 860.100 571.050 861.900 572.850 ;
        RECT 863.100 571.050 864.000 574.800 ;
        RECT 865.950 573.450 870.000 574.050 ;
        RECT 865.950 571.950 870.450 573.450 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 856.950 568.950 859.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 805.950 566.550 810.450 568.050 ;
        RECT 815.100 567.150 816.900 568.950 ;
        RECT 805.950 565.950 810.000 566.550 ;
        RECT 818.700 561.600 819.600 568.950 ;
        RECT 820.950 567.150 822.750 568.950 ;
        RECT 773.100 549.000 774.900 555.600 ;
        RECT 776.100 549.600 777.900 555.600 ;
        RECT 779.100 549.000 780.900 561.000 ;
        RECT 782.100 549.600 783.900 561.600 ;
        RECT 794.100 560.700 801.900 561.600 ;
        RECT 794.100 549.600 795.900 560.700 ;
        RECT 797.100 549.000 798.900 559.800 ;
        RECT 800.100 549.600 801.900 560.700 ;
        RECT 803.100 549.600 804.900 561.600 ;
        RECT 816.000 560.400 819.600 561.600 ;
        RECT 816.000 549.600 817.800 560.400 ;
        RECT 821.100 549.000 822.900 561.600 ;
        RECT 839.700 555.600 840.900 568.950 ;
        RECT 857.100 567.150 858.900 568.950 ;
        RECT 863.100 556.800 864.000 568.950 ;
        RECT 869.550 568.050 870.450 571.950 ;
        RECT 865.950 566.550 870.450 568.050 ;
        RECT 865.950 565.950 870.000 566.550 ;
        RECT 857.400 555.900 864.000 556.800 ;
        RECT 857.400 555.600 858.900 555.900 ;
        RECT 836.100 549.000 837.900 555.600 ;
        RECT 839.100 549.600 840.900 555.600 ;
        RECT 842.100 549.000 843.900 555.600 ;
        RECT 854.100 549.000 855.900 555.600 ;
        RECT 857.100 549.600 858.900 555.600 ;
        RECT 863.100 555.600 864.000 555.900 ;
        RECT 860.100 549.000 861.900 555.000 ;
        RECT 863.100 549.600 864.900 555.600 ;
        RECT 11.100 539.400 12.900 546.000 ;
        RECT 14.100 539.400 15.900 545.400 ;
        RECT 11.100 526.050 12.900 527.850 ;
        RECT 14.100 526.050 15.300 539.400 ;
        RECT 17.550 533.400 19.350 545.400 ;
        RECT 20.550 533.400 22.350 546.000 ;
        RECT 25.350 539.400 27.150 545.400 ;
        RECT 29.850 539.400 31.650 546.000 ;
        RECT 25.350 537.300 27.450 539.400 ;
        RECT 32.850 538.500 34.650 545.400 ;
        RECT 35.850 539.400 37.650 546.000 ;
        RECT 31.950 537.450 38.550 538.500 ;
        RECT 31.950 536.700 33.750 537.450 ;
        RECT 36.750 536.700 38.550 537.450 ;
        RECT 40.650 536.400 42.450 545.400 ;
        RECT 24.450 534.600 27.450 536.400 ;
        RECT 28.350 535.800 30.150 536.400 ;
        RECT 28.350 534.900 34.050 535.800 ;
        RECT 40.650 535.500 42.750 536.400 ;
        RECT 28.350 534.600 30.150 534.900 ;
        RECT 26.250 533.700 27.450 534.600 ;
        RECT 17.550 526.050 18.750 533.400 ;
        RECT 26.250 532.800 31.050 533.700 ;
        RECT 19.650 530.100 21.450 530.550 ;
        RECT 25.350 530.100 27.450 530.700 ;
        RECT 19.650 528.900 27.450 530.100 ;
        RECT 19.650 528.750 21.450 528.900 ;
        RECT 25.350 528.600 27.450 528.900 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 17.550 525.750 22.050 526.050 ;
        RECT 17.550 523.950 23.850 525.750 ;
        RECT 14.100 513.600 15.300 523.950 ;
        RECT 17.550 516.600 18.750 523.950 ;
        RECT 30.150 520.200 31.050 532.800 ;
        RECT 33.150 532.800 34.050 534.900 ;
        RECT 34.950 534.300 42.750 535.500 ;
        RECT 34.950 533.700 36.750 534.300 ;
        RECT 46.050 533.400 47.850 546.000 ;
        RECT 49.050 535.200 50.850 545.400 ;
        RECT 62.100 539.400 63.900 546.000 ;
        RECT 65.100 539.400 66.900 545.400 ;
        RECT 49.050 533.400 51.450 535.200 ;
        RECT 33.150 532.500 41.550 532.800 ;
        RECT 50.550 532.500 51.450 533.400 ;
        RECT 33.150 531.900 51.450 532.500 ;
        RECT 39.750 531.300 51.450 531.900 ;
        RECT 39.750 531.000 41.550 531.300 ;
        RECT 37.800 524.400 39.900 526.050 ;
        RECT 37.800 523.200 45.900 524.400 ;
        RECT 46.950 523.950 49.050 526.050 ;
        RECT 44.100 522.600 45.900 523.200 ;
        RECT 41.100 521.400 42.900 522.000 ;
        RECT 47.250 521.400 49.050 523.950 ;
        RECT 41.100 520.200 49.050 521.400 ;
        RECT 30.150 519.000 42.150 520.200 ;
        RECT 30.150 518.400 31.950 519.000 ;
        RECT 41.100 517.200 42.150 519.000 ;
        RECT 11.100 510.000 12.900 513.600 ;
        RECT 14.100 510.600 15.900 513.600 ;
        RECT 17.550 510.600 19.350 516.600 ;
        RECT 20.850 510.000 22.650 516.600 ;
        RECT 25.350 513.600 27.750 515.700 ;
        RECT 37.350 515.550 39.150 516.300 ;
        RECT 34.200 514.500 39.150 515.550 ;
        RECT 40.350 515.400 42.150 517.200 ;
        RECT 50.550 516.600 51.450 531.300 ;
        RECT 62.100 526.050 63.900 527.850 ;
        RECT 65.100 526.050 66.300 539.400 ;
        RECT 68.550 533.400 70.350 545.400 ;
        RECT 71.550 533.400 73.350 546.000 ;
        RECT 76.350 539.400 78.150 545.400 ;
        RECT 80.850 539.400 82.650 546.000 ;
        RECT 76.350 537.300 78.450 539.400 ;
        RECT 83.850 538.500 85.650 545.400 ;
        RECT 86.850 539.400 88.650 546.000 ;
        RECT 82.950 537.450 89.550 538.500 ;
        RECT 82.950 536.700 84.750 537.450 ;
        RECT 87.750 536.700 89.550 537.450 ;
        RECT 91.650 536.400 93.450 545.400 ;
        RECT 75.450 534.600 78.450 536.400 ;
        RECT 79.350 535.800 81.150 536.400 ;
        RECT 79.350 534.900 85.050 535.800 ;
        RECT 91.650 535.500 93.750 536.400 ;
        RECT 79.350 534.600 81.150 534.900 ;
        RECT 77.250 533.700 78.450 534.600 ;
        RECT 68.550 526.050 69.750 533.400 ;
        RECT 77.250 532.800 82.050 533.700 ;
        RECT 70.650 530.100 72.450 530.550 ;
        RECT 76.350 530.100 78.450 530.700 ;
        RECT 70.650 528.900 78.450 530.100 ;
        RECT 70.650 528.750 72.450 528.900 ;
        RECT 76.350 528.600 78.450 528.900 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 64.950 523.950 67.050 526.050 ;
        RECT 68.550 525.750 73.050 526.050 ;
        RECT 68.550 523.950 74.850 525.750 ;
        RECT 34.200 513.600 35.250 514.500 ;
        RECT 43.050 514.200 45.150 515.700 ;
        RECT 41.250 513.600 45.150 514.200 ;
        RECT 25.950 510.600 27.750 513.600 ;
        RECT 30.450 510.000 32.250 513.600 ;
        RECT 33.450 510.600 35.250 513.600 ;
        RECT 36.750 510.000 38.550 513.600 ;
        RECT 41.250 512.700 44.850 513.600 ;
        RECT 41.250 510.600 43.050 512.700 ;
        RECT 46.050 510.000 47.850 516.600 ;
        RECT 49.050 514.800 51.450 516.600 ;
        RECT 49.050 510.600 50.850 514.800 ;
        RECT 65.100 513.600 66.300 523.950 ;
        RECT 68.550 516.600 69.750 523.950 ;
        RECT 81.150 520.200 82.050 532.800 ;
        RECT 84.150 532.800 85.050 534.900 ;
        RECT 85.950 534.300 93.750 535.500 ;
        RECT 85.950 533.700 87.750 534.300 ;
        RECT 97.050 533.400 98.850 546.000 ;
        RECT 100.050 535.200 101.850 545.400 ;
        RECT 100.050 533.400 102.450 535.200 ;
        RECT 113.400 533.400 115.200 546.000 ;
        RECT 118.500 534.900 120.300 545.400 ;
        RECT 121.500 539.400 123.300 546.000 ;
        RECT 134.100 539.400 135.900 546.000 ;
        RECT 137.100 539.400 138.900 545.400 ;
        RECT 140.100 540.000 141.900 546.000 ;
        RECT 137.400 539.100 138.900 539.400 ;
        RECT 143.100 539.400 144.900 545.400 ;
        RECT 143.100 539.100 144.000 539.400 ;
        RECT 137.400 538.200 144.000 539.100 ;
        RECT 121.200 536.100 123.000 537.900 ;
        RECT 118.500 533.400 120.900 534.900 ;
        RECT 84.150 532.500 92.550 532.800 ;
        RECT 101.550 532.500 102.450 533.400 ;
        RECT 84.150 531.900 102.450 532.500 ;
        RECT 90.750 531.300 102.450 531.900 ;
        RECT 90.750 531.000 92.550 531.300 ;
        RECT 88.800 524.400 90.900 526.050 ;
        RECT 88.800 523.200 96.900 524.400 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 95.100 522.600 96.900 523.200 ;
        RECT 92.100 521.400 93.900 522.000 ;
        RECT 98.250 521.400 100.050 523.950 ;
        RECT 92.100 520.200 100.050 521.400 ;
        RECT 81.150 519.000 93.150 520.200 ;
        RECT 81.150 518.400 82.950 519.000 ;
        RECT 92.100 517.200 93.150 519.000 ;
        RECT 62.100 510.000 63.900 513.600 ;
        RECT 65.100 510.600 66.900 513.600 ;
        RECT 68.550 510.600 70.350 516.600 ;
        RECT 71.850 510.000 73.650 516.600 ;
        RECT 76.350 513.600 78.750 515.700 ;
        RECT 88.350 515.550 90.150 516.300 ;
        RECT 85.200 514.500 90.150 515.550 ;
        RECT 91.350 515.400 93.150 517.200 ;
        RECT 101.550 516.600 102.450 531.300 ;
        RECT 113.100 526.050 114.900 527.850 ;
        RECT 119.700 526.050 120.900 533.400 ;
        RECT 137.100 526.050 138.900 527.850 ;
        RECT 143.100 526.050 144.000 538.200 ;
        RECT 155.100 534.300 156.900 545.400 ;
        RECT 158.100 535.200 159.900 546.000 ;
        RECT 161.100 534.300 162.900 545.400 ;
        RECT 155.100 533.400 162.900 534.300 ;
        RECT 164.100 533.400 165.900 545.400 ;
        RECT 176.100 539.400 177.900 546.000 ;
        RECT 179.100 539.400 180.900 545.400 ;
        RECT 182.100 539.400 183.900 546.000 ;
        RECT 158.250 526.050 160.050 527.850 ;
        RECT 164.700 526.050 165.600 533.400 ;
        RECT 179.100 526.050 180.300 539.400 ;
        RECT 194.100 533.400 195.900 546.000 ;
        RECT 197.100 532.500 198.900 545.400 ;
        RECT 200.100 533.400 201.900 546.000 ;
        RECT 203.100 532.500 204.900 545.400 ;
        RECT 206.100 533.400 207.900 546.000 ;
        RECT 209.100 532.500 210.900 545.400 ;
        RECT 212.100 533.400 213.900 546.000 ;
        RECT 215.100 532.500 216.900 545.400 ;
        RECT 218.100 533.400 219.900 546.000 ;
        RECT 230.100 539.400 231.900 546.000 ;
        RECT 233.100 539.400 234.900 545.400 ;
        RECT 236.100 539.400 237.900 546.000 ;
        RECT 196.050 531.300 198.900 532.500 ;
        RECT 201.000 531.300 204.900 532.500 ;
        RECT 207.000 531.300 210.900 532.500 ;
        RECT 213.000 531.300 216.900 532.500 ;
        RECT 196.050 526.050 197.100 531.300 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 121.950 523.950 124.050 526.050 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 196.050 523.950 199.200 526.050 ;
        RECT 116.100 522.150 117.900 523.950 ;
        RECT 119.700 519.600 120.900 523.950 ;
        RECT 122.100 522.150 123.900 523.950 ;
        RECT 134.100 522.150 135.900 523.950 ;
        RECT 140.100 522.150 141.900 523.950 ;
        RECT 143.100 520.200 144.000 523.950 ;
        RECT 155.100 522.150 156.900 523.950 ;
        RECT 161.250 522.150 163.050 523.950 ;
        RECT 119.700 518.700 123.300 519.600 ;
        RECT 85.200 513.600 86.250 514.500 ;
        RECT 94.050 514.200 96.150 515.700 ;
        RECT 92.250 513.600 96.150 514.200 ;
        RECT 76.950 510.600 78.750 513.600 ;
        RECT 81.450 510.000 83.250 513.600 ;
        RECT 84.450 510.600 86.250 513.600 ;
        RECT 87.750 510.000 89.550 513.600 ;
        RECT 92.250 512.700 95.850 513.600 ;
        RECT 92.250 510.600 94.050 512.700 ;
        RECT 97.050 510.000 98.850 516.600 ;
        RECT 100.050 514.800 102.450 516.600 ;
        RECT 113.100 515.700 120.900 517.050 ;
        RECT 100.050 510.600 101.850 514.800 ;
        RECT 113.100 510.600 114.900 515.700 ;
        RECT 116.100 510.000 117.900 514.800 ;
        RECT 119.100 510.600 120.900 515.700 ;
        RECT 122.100 516.600 123.300 518.700 ;
        RECT 122.100 510.600 123.900 516.600 ;
        RECT 134.100 510.000 135.900 519.600 ;
        RECT 140.700 519.000 144.000 520.200 ;
        RECT 140.700 510.600 142.500 519.000 ;
        RECT 164.700 516.600 165.600 523.950 ;
        RECT 176.250 522.150 178.050 523.950 ;
        RECT 179.100 518.700 180.300 523.950 ;
        RECT 182.100 522.150 183.900 523.950 ;
        RECT 196.050 518.700 197.100 523.950 ;
        RECT 198.000 520.800 199.800 521.400 ;
        RECT 201.000 520.800 202.200 531.300 ;
        RECT 198.000 519.600 202.200 520.800 ;
        RECT 204.000 520.800 205.800 521.400 ;
        RECT 207.000 520.800 208.200 531.300 ;
        RECT 204.000 519.600 208.200 520.800 ;
        RECT 210.000 520.800 211.800 521.400 ;
        RECT 213.000 520.800 214.200 531.300 ;
        RECT 233.700 526.050 234.900 539.400 ;
        RECT 248.100 534.300 249.900 545.400 ;
        RECT 251.100 535.500 252.900 546.000 ;
        RECT 255.600 534.300 257.400 545.400 ;
        RECT 259.800 535.500 261.900 546.000 ;
        RECT 263.100 534.600 264.900 545.400 ;
        RECT 248.100 533.100 252.900 534.300 ;
        RECT 255.600 533.400 258.900 534.300 ;
        RECT 250.800 532.200 252.900 533.100 ;
        RECT 235.950 531.450 238.050 532.050 ;
        RECT 235.950 530.550 243.450 531.450 ;
        RECT 250.800 531.300 256.200 532.200 ;
        RECT 235.950 529.950 238.050 530.550 ;
        RECT 215.100 523.950 217.200 526.050 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 215.400 522.150 217.200 523.950 ;
        RECT 230.100 522.150 231.900 523.950 ;
        RECT 210.000 519.600 214.200 520.800 ;
        RECT 201.000 518.700 202.200 519.600 ;
        RECT 207.000 518.700 208.200 519.600 ;
        RECT 213.000 518.700 214.200 519.600 ;
        RECT 233.700 518.700 234.900 523.950 ;
        RECT 235.950 522.150 237.750 523.950 ;
        RECT 242.550 523.050 243.450 530.550 ;
        RECT 254.400 529.500 256.200 531.300 ;
        RECT 257.700 529.050 258.900 533.400 ;
        RECT 259.800 533.400 264.900 534.600 ;
        RECT 275.100 534.300 276.900 545.400 ;
        RECT 278.100 535.200 279.900 546.000 ;
        RECT 281.100 534.300 282.900 545.400 ;
        RECT 275.100 533.400 282.900 534.300 ;
        RECT 284.100 533.400 285.900 545.400 ;
        RECT 297.000 534.600 298.800 545.400 ;
        RECT 297.000 533.400 300.600 534.600 ;
        RECT 302.100 533.400 303.900 546.000 ;
        RECT 317.100 539.400 318.900 546.000 ;
        RECT 320.100 539.400 321.900 545.400 ;
        RECT 259.800 532.500 261.900 533.400 ;
        RECT 257.100 528.300 259.200 529.050 ;
        RECT 252.900 526.200 254.700 528.000 ;
        RECT 256.200 526.950 259.200 528.300 ;
        RECT 248.100 523.800 250.200 526.050 ;
        RECT 252.900 524.100 255.000 526.200 ;
        RECT 238.950 521.550 243.450 523.050 ;
        RECT 248.400 523.200 250.200 523.800 ;
        RECT 248.400 522.000 255.000 523.200 ;
        RECT 238.950 520.950 243.000 521.550 ;
        RECT 252.900 521.100 255.000 522.000 ;
        RECT 250.500 519.000 252.600 519.600 ;
        RECT 253.500 519.300 255.300 521.100 ;
        RECT 256.200 520.200 257.100 526.950 ;
        RECT 262.800 526.050 264.600 527.850 ;
        RECT 278.250 526.050 280.050 527.850 ;
        RECT 284.700 526.050 285.600 533.400 ;
        RECT 296.100 526.050 297.900 527.850 ;
        RECT 299.700 526.050 300.600 533.400 ;
        RECT 301.950 526.050 303.750 527.850 ;
        RECT 317.100 526.050 318.900 527.850 ;
        RECT 320.100 526.050 321.300 539.400 ;
        RECT 332.400 533.400 334.200 546.000 ;
        RECT 337.500 534.900 339.300 545.400 ;
        RECT 340.500 539.400 342.300 546.000 ;
        RECT 353.100 539.400 354.900 545.400 ;
        RECT 340.200 536.100 342.000 537.900 ;
        RECT 337.500 533.400 339.900 534.900 ;
        RECT 332.100 526.050 333.900 527.850 ;
        RECT 338.700 526.050 339.900 533.400 ;
        RECT 353.100 532.500 354.300 539.400 ;
        RECT 356.100 535.200 357.900 546.000 ;
        RECT 359.100 533.400 360.900 545.400 ;
        RECT 371.100 539.400 372.900 546.000 ;
        RECT 374.100 539.400 375.900 545.400 ;
        RECT 377.100 539.400 378.900 546.000 ;
        RECT 389.100 539.400 390.900 546.000 ;
        RECT 392.100 539.400 393.900 545.400 ;
        RECT 395.100 539.400 396.900 546.000 ;
        RECT 407.100 539.400 408.900 546.000 ;
        RECT 410.100 539.400 411.900 545.400 ;
        RECT 413.100 539.400 414.900 546.000 ;
        RECT 353.100 531.600 358.800 532.500 ;
        RECT 357.000 530.700 358.800 531.600 ;
        RECT 353.400 526.050 355.200 527.850 ;
        RECT 258.000 524.100 259.800 525.900 ;
        RECT 258.000 522.000 260.100 524.100 ;
        RECT 262.800 523.950 264.900 526.050 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 334.950 523.950 337.050 526.050 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 353.400 523.950 355.500 526.050 ;
        RECT 275.100 522.150 276.900 523.950 ;
        RECT 281.250 522.150 283.050 523.950 ;
        RECT 179.100 517.800 183.300 518.700 ;
        RECT 156.000 510.000 157.800 516.600 ;
        RECT 160.500 515.400 165.600 516.600 ;
        RECT 160.500 510.600 162.300 515.400 ;
        RECT 163.500 510.000 165.300 513.600 ;
        RECT 176.400 510.000 178.200 516.600 ;
        RECT 181.500 510.600 183.300 517.800 ;
        RECT 196.050 517.500 198.900 518.700 ;
        RECT 201.000 517.500 204.900 518.700 ;
        RECT 207.000 517.500 210.900 518.700 ;
        RECT 213.000 517.500 216.900 518.700 ;
        RECT 194.100 510.000 195.900 516.600 ;
        RECT 197.100 510.600 198.900 517.500 ;
        RECT 200.100 510.000 201.900 516.600 ;
        RECT 203.100 510.600 204.900 517.500 ;
        RECT 206.100 510.000 207.900 516.600 ;
        RECT 209.100 510.600 210.900 517.500 ;
        RECT 212.100 510.000 213.900 516.600 ;
        RECT 215.100 510.600 216.900 517.500 ;
        RECT 230.700 517.800 234.900 518.700 ;
        RECT 218.100 510.000 219.900 516.600 ;
        RECT 230.700 510.600 232.500 517.800 ;
        RECT 248.100 517.500 252.600 519.000 ;
        RECT 256.200 518.100 259.200 520.200 ;
        RECT 248.100 516.600 249.600 517.500 ;
        RECT 235.800 510.000 237.600 516.600 ;
        RECT 248.100 510.600 249.900 516.600 ;
        RECT 256.200 516.000 257.100 518.100 ;
        RECT 260.400 517.500 262.500 519.900 ;
        RECT 260.400 516.600 264.900 517.500 ;
        RECT 284.700 516.600 285.600 523.950 ;
        RECT 251.100 510.000 252.900 515.700 ;
        RECT 255.300 510.600 257.100 516.000 ;
        RECT 259.800 510.000 261.600 515.700 ;
        RECT 263.100 510.600 264.900 516.600 ;
        RECT 276.000 510.000 277.800 516.600 ;
        RECT 280.500 515.400 285.600 516.600 ;
        RECT 280.500 510.600 282.300 515.400 ;
        RECT 299.700 513.600 300.600 523.950 ;
        RECT 307.950 522.450 310.050 523.050 ;
        RECT 313.950 522.450 316.050 523.050 ;
        RECT 307.950 521.550 316.050 522.450 ;
        RECT 307.950 520.950 310.050 521.550 ;
        RECT 313.950 520.950 316.050 521.550 ;
        RECT 320.100 513.600 321.300 523.950 ;
        RECT 335.100 522.150 336.900 523.950 ;
        RECT 338.700 519.600 339.900 523.950 ;
        RECT 341.100 522.150 342.900 523.950 ;
        RECT 338.700 518.700 342.300 519.600 ;
        RECT 332.100 515.700 339.900 517.050 ;
        RECT 283.500 510.000 285.300 513.600 ;
        RECT 296.100 510.000 297.900 513.600 ;
        RECT 299.100 510.600 300.900 513.600 ;
        RECT 302.100 510.000 303.900 513.600 ;
        RECT 317.100 510.000 318.900 513.600 ;
        RECT 320.100 510.600 321.900 513.600 ;
        RECT 332.100 510.600 333.900 515.700 ;
        RECT 335.100 510.000 336.900 514.800 ;
        RECT 338.100 510.600 339.900 515.700 ;
        RECT 341.100 516.600 342.300 518.700 ;
        RECT 357.000 519.300 357.900 530.700 ;
        RECT 359.700 526.050 360.900 533.400 ;
        RECT 374.100 526.050 375.300 539.400 ;
        RECT 392.100 526.050 393.300 539.400 ;
        RECT 410.700 526.050 411.900 539.400 ;
        RECT 417.150 535.200 418.950 545.400 ;
        RECT 416.550 533.400 418.950 535.200 ;
        RECT 420.150 533.400 421.950 546.000 ;
        RECT 425.550 536.400 427.350 545.400 ;
        RECT 430.350 539.400 432.150 546.000 ;
        RECT 433.350 538.500 435.150 545.400 ;
        RECT 436.350 539.400 438.150 546.000 ;
        RECT 440.850 539.400 442.650 545.400 ;
        RECT 429.450 537.450 436.050 538.500 ;
        RECT 429.450 536.700 431.250 537.450 ;
        RECT 434.250 536.700 436.050 537.450 ;
        RECT 440.550 537.300 442.650 539.400 ;
        RECT 425.250 535.500 427.350 536.400 ;
        RECT 437.850 535.800 439.650 536.400 ;
        RECT 425.250 534.300 433.050 535.500 ;
        RECT 431.250 533.700 433.050 534.300 ;
        RECT 433.950 534.900 439.650 535.800 ;
        RECT 416.550 532.500 417.450 533.400 ;
        RECT 433.950 532.800 434.850 534.900 ;
        RECT 437.850 534.600 439.650 534.900 ;
        RECT 440.550 534.600 443.550 536.400 ;
        RECT 440.550 533.700 441.750 534.600 ;
        RECT 426.450 532.500 434.850 532.800 ;
        RECT 416.550 531.900 434.850 532.500 ;
        RECT 436.950 532.800 441.750 533.700 ;
        RECT 445.650 533.400 447.450 546.000 ;
        RECT 448.650 533.400 450.450 545.400 ;
        RECT 464.100 533.400 465.900 546.000 ;
        RECT 467.100 533.400 468.900 545.400 ;
        RECT 479.100 533.400 480.900 546.000 ;
        RECT 484.200 534.600 486.000 545.400 ;
        RECT 482.400 533.400 486.000 534.600 ;
        RECT 488.550 533.400 490.350 545.400 ;
        RECT 491.550 533.400 493.350 546.000 ;
        RECT 496.350 539.400 498.150 545.400 ;
        RECT 500.850 539.400 502.650 546.000 ;
        RECT 496.350 537.300 498.450 539.400 ;
        RECT 503.850 538.500 505.650 545.400 ;
        RECT 506.850 539.400 508.650 546.000 ;
        RECT 502.950 537.450 509.550 538.500 ;
        RECT 502.950 536.700 504.750 537.450 ;
        RECT 507.750 536.700 509.550 537.450 ;
        RECT 511.650 536.400 513.450 545.400 ;
        RECT 495.450 534.600 498.450 536.400 ;
        RECT 499.350 535.800 501.150 536.400 ;
        RECT 499.350 534.900 505.050 535.800 ;
        RECT 511.650 535.500 513.750 536.400 ;
        RECT 499.350 534.600 501.150 534.900 ;
        RECT 497.250 533.700 498.450 534.600 ;
        RECT 416.550 531.300 428.250 531.900 ;
        RECT 358.800 523.950 360.900 526.050 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 357.000 518.400 358.800 519.300 ;
        RECT 353.100 517.500 358.800 518.400 ;
        RECT 341.100 510.600 342.900 516.600 ;
        RECT 353.100 513.600 354.300 517.500 ;
        RECT 359.700 516.600 360.900 523.950 ;
        RECT 371.250 522.150 373.050 523.950 ;
        RECT 374.100 518.700 375.300 523.950 ;
        RECT 377.100 522.150 378.900 523.950 ;
        RECT 389.250 522.150 391.050 523.950 ;
        RECT 392.100 518.700 393.300 523.950 ;
        RECT 395.100 522.150 396.900 523.950 ;
        RECT 407.100 522.150 408.900 523.950 ;
        RECT 410.700 518.700 411.900 523.950 ;
        RECT 412.950 522.150 414.750 523.950 ;
        RECT 374.100 517.800 378.300 518.700 ;
        RECT 392.100 517.800 396.300 518.700 ;
        RECT 353.100 510.600 354.900 513.600 ;
        RECT 356.100 510.000 357.900 516.600 ;
        RECT 359.100 510.600 360.900 516.600 ;
        RECT 371.400 510.000 373.200 516.600 ;
        RECT 376.500 510.600 378.300 517.800 ;
        RECT 389.400 510.000 391.200 516.600 ;
        RECT 394.500 510.600 396.300 517.800 ;
        RECT 407.700 517.800 411.900 518.700 ;
        RECT 407.700 510.600 409.500 517.800 ;
        RECT 416.550 516.600 417.450 531.300 ;
        RECT 426.450 531.000 428.250 531.300 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 428.100 524.400 430.200 526.050 ;
        RECT 418.950 521.400 420.750 523.950 ;
        RECT 422.100 523.200 430.200 524.400 ;
        RECT 422.100 522.600 423.900 523.200 ;
        RECT 425.100 521.400 426.900 522.000 ;
        RECT 418.950 520.200 426.900 521.400 ;
        RECT 436.950 520.200 437.850 532.800 ;
        RECT 440.550 530.100 442.650 530.700 ;
        RECT 446.550 530.100 448.350 530.550 ;
        RECT 440.550 528.900 448.350 530.100 ;
        RECT 440.550 528.600 442.650 528.900 ;
        RECT 446.550 528.750 448.350 528.900 ;
        RECT 449.250 526.050 450.450 533.400 ;
        RECT 467.100 526.050 468.300 533.400 ;
        RECT 479.250 526.050 481.050 527.850 ;
        RECT 482.400 526.050 483.300 533.400 ;
        RECT 485.100 526.050 486.900 527.850 ;
        RECT 488.550 526.050 489.750 533.400 ;
        RECT 497.250 532.800 502.050 533.700 ;
        RECT 490.650 530.100 492.450 530.550 ;
        RECT 496.350 530.100 498.450 530.700 ;
        RECT 490.650 528.900 498.450 530.100 ;
        RECT 490.650 528.750 492.450 528.900 ;
        RECT 496.350 528.600 498.450 528.900 ;
        RECT 445.950 525.750 450.450 526.050 ;
        RECT 444.150 523.950 450.450 525.750 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 478.950 523.950 481.050 526.050 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 488.550 525.750 493.050 526.050 ;
        RECT 488.550 523.950 494.850 525.750 ;
        RECT 425.850 519.000 437.850 520.200 ;
        RECT 425.850 517.200 426.900 519.000 ;
        RECT 436.050 518.400 437.850 519.000 ;
        RECT 412.800 510.000 414.600 516.600 ;
        RECT 416.550 514.800 418.950 516.600 ;
        RECT 417.150 510.600 418.950 514.800 ;
        RECT 420.150 510.000 421.950 516.600 ;
        RECT 422.850 514.200 424.950 515.700 ;
        RECT 425.850 515.400 427.650 517.200 ;
        RECT 449.250 516.600 450.450 523.950 ;
        RECT 464.100 522.150 465.900 523.950 ;
        RECT 467.100 516.600 468.300 523.950 ;
        RECT 428.850 515.550 430.650 516.300 ;
        RECT 428.850 514.500 433.800 515.550 ;
        RECT 422.850 513.600 426.750 514.200 ;
        RECT 432.750 513.600 433.800 514.500 ;
        RECT 440.250 513.600 442.650 515.700 ;
        RECT 423.150 512.700 426.750 513.600 ;
        RECT 424.950 510.600 426.750 512.700 ;
        RECT 429.450 510.000 431.250 513.600 ;
        RECT 432.750 510.600 434.550 513.600 ;
        RECT 435.750 510.000 437.550 513.600 ;
        RECT 440.250 510.600 442.050 513.600 ;
        RECT 445.350 510.000 447.150 516.600 ;
        RECT 448.650 510.600 450.450 516.600 ;
        RECT 464.100 510.000 465.900 516.600 ;
        RECT 467.100 510.600 468.900 516.600 ;
        RECT 482.400 513.600 483.300 523.950 ;
        RECT 488.550 516.600 489.750 523.950 ;
        RECT 501.150 520.200 502.050 532.800 ;
        RECT 504.150 532.800 505.050 534.900 ;
        RECT 505.950 534.300 513.750 535.500 ;
        RECT 505.950 533.700 507.750 534.300 ;
        RECT 517.050 533.400 518.850 546.000 ;
        RECT 520.050 535.200 521.850 545.400 ;
        RECT 520.050 533.400 522.450 535.200 ;
        RECT 533.100 533.400 534.900 545.400 ;
        RECT 536.100 534.300 537.900 545.400 ;
        RECT 539.100 535.200 540.900 546.000 ;
        RECT 542.100 534.300 543.900 545.400 ;
        RECT 536.100 533.400 543.900 534.300 ;
        RECT 555.000 534.600 556.800 545.400 ;
        RECT 555.000 533.400 558.600 534.600 ;
        RECT 560.100 533.400 561.900 546.000 ;
        RECT 573.000 534.600 574.800 545.400 ;
        RECT 573.000 533.400 576.600 534.600 ;
        RECT 578.100 533.400 579.900 546.000 ;
        RECT 590.100 533.400 591.900 545.400 ;
        RECT 593.100 534.300 594.900 545.400 ;
        RECT 596.100 535.200 597.900 546.000 ;
        RECT 599.100 534.300 600.900 545.400 ;
        RECT 593.100 533.400 600.900 534.300 ;
        RECT 611.400 533.400 613.200 546.000 ;
        RECT 616.500 534.900 618.300 545.400 ;
        RECT 619.500 539.400 621.300 546.000 ;
        RECT 619.200 536.100 621.000 537.900 ;
        RECT 624.150 535.200 625.950 545.400 ;
        RECT 616.500 533.400 618.900 534.900 ;
        RECT 504.150 532.500 512.550 532.800 ;
        RECT 521.550 532.500 522.450 533.400 ;
        RECT 504.150 531.900 522.450 532.500 ;
        RECT 510.750 531.300 522.450 531.900 ;
        RECT 510.750 531.000 512.550 531.300 ;
        RECT 508.800 524.400 510.900 526.050 ;
        RECT 508.800 523.200 516.900 524.400 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 515.100 522.600 516.900 523.200 ;
        RECT 512.100 521.400 513.900 522.000 ;
        RECT 518.250 521.400 520.050 523.950 ;
        RECT 512.100 520.200 520.050 521.400 ;
        RECT 501.150 519.000 513.150 520.200 ;
        RECT 501.150 518.400 502.950 519.000 ;
        RECT 512.100 517.200 513.150 519.000 ;
        RECT 479.100 510.000 480.900 513.600 ;
        RECT 482.100 510.600 483.900 513.600 ;
        RECT 485.100 510.000 486.900 513.600 ;
        RECT 488.550 510.600 490.350 516.600 ;
        RECT 491.850 510.000 493.650 516.600 ;
        RECT 496.350 513.600 498.750 515.700 ;
        RECT 508.350 515.550 510.150 516.300 ;
        RECT 505.200 514.500 510.150 515.550 ;
        RECT 511.350 515.400 513.150 517.200 ;
        RECT 521.550 516.600 522.450 531.300 ;
        RECT 533.400 526.050 534.300 533.400 ;
        RECT 538.950 526.050 540.750 527.850 ;
        RECT 554.100 526.050 555.900 527.850 ;
        RECT 557.700 526.050 558.600 533.400 ;
        RECT 559.950 526.050 561.750 527.850 ;
        RECT 572.100 526.050 573.900 527.850 ;
        RECT 575.700 526.050 576.600 533.400 ;
        RECT 577.950 526.050 579.750 527.850 ;
        RECT 590.400 526.050 591.300 533.400 ;
        RECT 595.950 526.050 597.750 527.850 ;
        RECT 611.100 526.050 612.900 527.850 ;
        RECT 617.700 526.050 618.900 533.400 ;
        RECT 623.550 533.400 625.950 535.200 ;
        RECT 627.150 533.400 628.950 546.000 ;
        RECT 632.550 536.400 634.350 545.400 ;
        RECT 637.350 539.400 639.150 546.000 ;
        RECT 640.350 538.500 642.150 545.400 ;
        RECT 643.350 539.400 645.150 546.000 ;
        RECT 647.850 539.400 649.650 545.400 ;
        RECT 636.450 537.450 643.050 538.500 ;
        RECT 636.450 536.700 638.250 537.450 ;
        RECT 641.250 536.700 643.050 537.450 ;
        RECT 647.550 537.300 649.650 539.400 ;
        RECT 632.250 535.500 634.350 536.400 ;
        RECT 644.850 535.800 646.650 536.400 ;
        RECT 632.250 534.300 640.050 535.500 ;
        RECT 638.250 533.700 640.050 534.300 ;
        RECT 640.950 534.900 646.650 535.800 ;
        RECT 623.550 532.500 624.450 533.400 ;
        RECT 640.950 532.800 641.850 534.900 ;
        RECT 644.850 534.600 646.650 534.900 ;
        RECT 647.550 534.600 650.550 536.400 ;
        RECT 647.550 533.700 648.750 534.600 ;
        RECT 633.450 532.500 641.850 532.800 ;
        RECT 623.550 531.900 641.850 532.500 ;
        RECT 643.950 532.800 648.750 533.700 ;
        RECT 652.650 533.400 654.450 546.000 ;
        RECT 655.650 533.400 657.450 545.400 ;
        RECT 668.100 539.400 669.900 546.000 ;
        RECT 671.100 539.400 672.900 545.400 ;
        RECT 674.100 539.400 675.900 546.000 ;
        RECT 686.100 539.400 687.900 546.000 ;
        RECT 689.100 539.400 690.900 545.400 ;
        RECT 692.100 539.400 693.900 546.000 ;
        RECT 704.100 539.400 705.900 545.400 ;
        RECT 623.550 531.300 635.250 531.900 ;
        RECT 532.950 523.950 535.050 526.050 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 541.950 523.950 544.050 526.050 ;
        RECT 553.950 523.950 556.050 526.050 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 577.950 523.950 580.050 526.050 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 595.950 523.950 598.050 526.050 ;
        RECT 598.950 523.950 601.050 526.050 ;
        RECT 610.950 523.950 613.050 526.050 ;
        RECT 613.950 523.950 616.050 526.050 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 505.200 513.600 506.250 514.500 ;
        RECT 514.050 514.200 516.150 515.700 ;
        RECT 512.250 513.600 516.150 514.200 ;
        RECT 496.950 510.600 498.750 513.600 ;
        RECT 501.450 510.000 503.250 513.600 ;
        RECT 504.450 510.600 506.250 513.600 ;
        RECT 507.750 510.000 509.550 513.600 ;
        RECT 512.250 512.700 515.850 513.600 ;
        RECT 512.250 510.600 514.050 512.700 ;
        RECT 517.050 510.000 518.850 516.600 ;
        RECT 520.050 514.800 522.450 516.600 ;
        RECT 533.400 516.600 534.300 523.950 ;
        RECT 535.950 522.150 537.750 523.950 ;
        RECT 542.100 522.150 543.900 523.950 ;
        RECT 533.400 515.400 538.500 516.600 ;
        RECT 520.050 510.600 521.850 514.800 ;
        RECT 533.700 510.000 535.500 513.600 ;
        RECT 536.700 510.600 538.500 515.400 ;
        RECT 541.200 510.000 543.000 516.600 ;
        RECT 557.700 513.600 558.600 523.950 ;
        RECT 575.700 513.600 576.600 523.950 ;
        RECT 590.400 516.600 591.300 523.950 ;
        RECT 592.950 522.150 594.750 523.950 ;
        RECT 599.100 522.150 600.900 523.950 ;
        RECT 614.100 522.150 615.900 523.950 ;
        RECT 595.950 519.450 598.050 520.050 ;
        RECT 604.950 519.450 607.050 520.050 ;
        RECT 595.950 518.550 607.050 519.450 ;
        RECT 617.700 519.600 618.900 523.950 ;
        RECT 620.100 522.150 621.900 523.950 ;
        RECT 617.700 518.700 621.300 519.600 ;
        RECT 595.950 517.950 598.050 518.550 ;
        RECT 604.950 517.950 607.050 518.550 ;
        RECT 590.400 515.400 595.500 516.600 ;
        RECT 554.100 510.000 555.900 513.600 ;
        RECT 557.100 510.600 558.900 513.600 ;
        RECT 560.100 510.000 561.900 513.600 ;
        RECT 572.100 510.000 573.900 513.600 ;
        RECT 575.100 510.600 576.900 513.600 ;
        RECT 578.100 510.000 579.900 513.600 ;
        RECT 590.700 510.000 592.500 513.600 ;
        RECT 593.700 510.600 595.500 515.400 ;
        RECT 598.200 510.000 600.000 516.600 ;
        RECT 611.100 515.700 618.900 517.050 ;
        RECT 611.100 510.600 612.900 515.700 ;
        RECT 614.100 510.000 615.900 514.800 ;
        RECT 617.100 510.600 618.900 515.700 ;
        RECT 620.100 516.600 621.300 518.700 ;
        RECT 623.550 516.600 624.450 531.300 ;
        RECT 633.450 531.000 635.250 531.300 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 635.100 524.400 637.200 526.050 ;
        RECT 625.950 521.400 627.750 523.950 ;
        RECT 629.100 523.200 637.200 524.400 ;
        RECT 629.100 522.600 630.900 523.200 ;
        RECT 632.100 521.400 633.900 522.000 ;
        RECT 625.950 520.200 633.900 521.400 ;
        RECT 643.950 520.200 644.850 532.800 ;
        RECT 647.550 530.100 649.650 530.700 ;
        RECT 653.550 530.100 655.350 530.550 ;
        RECT 647.550 528.900 655.350 530.100 ;
        RECT 647.550 528.600 649.650 528.900 ;
        RECT 653.550 528.750 655.350 528.900 ;
        RECT 656.250 526.050 657.450 533.400 ;
        RECT 671.700 526.050 672.900 539.400 ;
        RECT 689.100 526.050 690.300 539.400 ;
        RECT 704.100 532.500 705.300 539.400 ;
        RECT 707.100 535.200 708.900 546.000 ;
        RECT 710.100 533.400 711.900 545.400 ;
        RECT 722.400 533.400 724.200 546.000 ;
        RECT 727.500 534.900 729.300 545.400 ;
        RECT 730.500 539.400 732.300 546.000 ;
        RECT 743.100 539.400 744.900 545.400 ;
        RECT 746.100 539.400 747.900 546.000 ;
        RECT 758.100 539.400 759.900 545.400 ;
        RECT 761.100 540.000 762.900 546.000 ;
        RECT 730.200 536.100 732.000 537.900 ;
        RECT 727.500 533.400 729.900 534.900 ;
        RECT 704.100 531.600 709.800 532.500 ;
        RECT 708.000 530.700 709.800 531.600 ;
        RECT 704.400 526.050 706.200 527.850 ;
        RECT 652.950 525.750 657.450 526.050 ;
        RECT 651.150 523.950 657.450 525.750 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 704.400 523.950 706.500 526.050 ;
        RECT 632.850 519.000 644.850 520.200 ;
        RECT 632.850 517.200 633.900 519.000 ;
        RECT 643.050 518.400 644.850 519.000 ;
        RECT 620.100 510.600 621.900 516.600 ;
        RECT 623.550 514.800 625.950 516.600 ;
        RECT 624.150 510.600 625.950 514.800 ;
        RECT 627.150 510.000 628.950 516.600 ;
        RECT 629.850 514.200 631.950 515.700 ;
        RECT 632.850 515.400 634.650 517.200 ;
        RECT 656.250 516.600 657.450 523.950 ;
        RECT 668.100 522.150 669.900 523.950 ;
        RECT 671.700 518.700 672.900 523.950 ;
        RECT 673.950 522.150 675.750 523.950 ;
        RECT 686.250 522.150 688.050 523.950 ;
        RECT 635.850 515.550 637.650 516.300 ;
        RECT 635.850 514.500 640.800 515.550 ;
        RECT 629.850 513.600 633.750 514.200 ;
        RECT 639.750 513.600 640.800 514.500 ;
        RECT 647.250 513.600 649.650 515.700 ;
        RECT 630.150 512.700 633.750 513.600 ;
        RECT 631.950 510.600 633.750 512.700 ;
        RECT 636.450 510.000 638.250 513.600 ;
        RECT 639.750 510.600 641.550 513.600 ;
        RECT 642.750 510.000 644.550 513.600 ;
        RECT 647.250 510.600 649.050 513.600 ;
        RECT 652.350 510.000 654.150 516.600 ;
        RECT 655.650 510.600 657.450 516.600 ;
        RECT 668.700 517.800 672.900 518.700 ;
        RECT 689.100 518.700 690.300 523.950 ;
        RECT 692.100 522.150 693.900 523.950 ;
        RECT 708.000 519.300 708.900 530.700 ;
        RECT 710.700 526.050 711.900 533.400 ;
        RECT 722.100 526.050 723.900 527.850 ;
        RECT 728.700 526.050 729.900 533.400 ;
        RECT 743.700 526.050 744.900 539.400 ;
        RECT 759.000 539.100 759.900 539.400 ;
        RECT 764.100 539.400 765.900 545.400 ;
        RECT 767.100 539.400 768.900 546.000 ;
        RECT 779.100 539.400 780.900 546.000 ;
        RECT 782.100 539.400 783.900 545.400 ;
        RECT 785.100 539.400 786.900 546.000 ;
        RECT 797.700 539.400 799.500 546.000 ;
        RECT 764.100 539.100 765.600 539.400 ;
        RECT 759.000 538.200 765.600 539.100 ;
        RECT 746.100 526.050 747.900 527.850 ;
        RECT 759.000 526.050 759.900 538.200 ;
        RECT 763.950 531.450 766.050 532.050 ;
        RECT 763.950 530.550 771.450 531.450 ;
        RECT 763.950 529.950 766.050 530.550 ;
        RECT 770.550 528.450 771.450 530.550 ;
        RECT 764.100 526.050 765.900 527.850 ;
        RECT 770.550 527.550 774.450 528.450 ;
        RECT 709.800 523.950 711.900 526.050 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 727.950 523.950 730.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 757.950 523.950 760.050 526.050 ;
        RECT 760.950 523.950 763.050 526.050 ;
        RECT 763.950 523.950 766.050 526.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 689.100 517.800 693.300 518.700 ;
        RECT 708.000 518.400 709.800 519.300 ;
        RECT 668.700 510.600 670.500 517.800 ;
        RECT 673.800 510.000 675.600 516.600 ;
        RECT 686.400 510.000 688.200 516.600 ;
        RECT 691.500 510.600 693.300 517.800 ;
        RECT 704.100 517.500 709.800 518.400 ;
        RECT 704.100 513.600 705.300 517.500 ;
        RECT 710.700 516.600 711.900 523.950 ;
        RECT 725.100 522.150 726.900 523.950 ;
        RECT 728.700 519.600 729.900 523.950 ;
        RECT 731.100 522.150 732.900 523.950 ;
        RECT 728.700 518.700 732.300 519.600 ;
        RECT 704.100 510.600 705.900 513.600 ;
        RECT 707.100 510.000 708.900 516.600 ;
        RECT 710.100 510.600 711.900 516.600 ;
        RECT 722.100 515.700 729.900 517.050 ;
        RECT 722.100 510.600 723.900 515.700 ;
        RECT 725.100 510.000 726.900 514.800 ;
        RECT 728.100 510.600 729.900 515.700 ;
        RECT 731.100 516.600 732.300 518.700 ;
        RECT 731.100 510.600 732.900 516.600 ;
        RECT 743.700 513.600 744.900 523.950 ;
        RECT 759.000 520.200 759.900 523.950 ;
        RECT 761.100 522.150 762.900 523.950 ;
        RECT 767.100 522.150 768.900 523.950 ;
        RECT 773.550 523.050 774.450 527.550 ;
        RECT 782.700 526.050 783.900 539.400 ;
        RECT 798.000 536.100 799.800 537.900 ;
        RECT 800.700 534.900 802.500 545.400 ;
        RECT 800.100 533.400 802.500 534.900 ;
        RECT 805.800 533.400 807.600 546.000 ;
        RECT 821.100 539.400 822.900 545.400 ;
        RECT 824.100 539.400 825.900 546.000 ;
        RECT 800.100 526.050 801.300 533.400 ;
        RECT 817.950 528.450 820.050 529.050 ;
        RECT 806.100 526.050 807.900 527.850 ;
        RECT 812.550 527.550 820.050 528.450 ;
        RECT 778.950 523.950 781.050 526.050 ;
        RECT 781.950 523.950 784.050 526.050 ;
        RECT 784.950 523.950 787.050 526.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 805.950 523.950 808.050 526.050 ;
        RECT 769.950 521.550 774.450 523.050 ;
        RECT 779.100 522.150 780.900 523.950 ;
        RECT 769.950 520.950 774.000 521.550 ;
        RECT 759.000 519.000 762.300 520.200 ;
        RECT 743.100 510.600 744.900 513.600 ;
        RECT 746.100 510.000 747.900 513.600 ;
        RECT 760.500 510.600 762.300 519.000 ;
        RECT 767.100 510.000 768.900 519.600 ;
        RECT 782.700 518.700 783.900 523.950 ;
        RECT 784.950 522.150 786.750 523.950 ;
        RECT 797.100 522.150 798.900 523.950 ;
        RECT 800.100 519.600 801.300 523.950 ;
        RECT 803.100 522.150 804.900 523.950 ;
        RECT 812.550 523.050 813.450 527.550 ;
        RECT 817.950 526.950 820.050 527.550 ;
        RECT 821.700 526.050 822.900 539.400 ;
        RECT 836.400 533.400 838.200 546.000 ;
        RECT 841.500 534.900 843.300 545.400 ;
        RECT 844.500 539.400 846.300 546.000 ;
        RECT 857.100 539.400 858.900 546.000 ;
        RECT 860.100 539.400 861.900 545.400 ;
        RECT 863.100 539.400 864.900 546.000 ;
        RECT 844.200 536.100 846.000 537.900 ;
        RECT 841.500 533.400 843.900 534.900 ;
        RECT 824.100 526.050 825.900 527.850 ;
        RECT 836.100 526.050 837.900 527.850 ;
        RECT 842.700 526.050 843.900 533.400 ;
        RECT 844.950 534.450 847.050 535.050 ;
        RECT 856.950 534.450 859.050 535.050 ;
        RECT 844.950 533.550 859.050 534.450 ;
        RECT 844.950 532.950 847.050 533.550 ;
        RECT 856.950 532.950 859.050 533.550 ;
        RECT 850.950 529.950 853.050 532.050 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 835.950 523.950 838.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 808.950 521.550 813.450 523.050 ;
        RECT 808.950 520.950 813.000 521.550 ;
        RECT 779.700 517.800 783.900 518.700 ;
        RECT 797.700 518.700 801.300 519.600 ;
        RECT 779.700 510.600 781.500 517.800 ;
        RECT 797.700 516.600 798.900 518.700 ;
        RECT 784.800 510.000 786.600 516.600 ;
        RECT 797.100 510.600 798.900 516.600 ;
        RECT 800.100 515.700 807.900 517.050 ;
        RECT 800.100 510.600 801.900 515.700 ;
        RECT 803.100 510.000 804.900 514.800 ;
        RECT 806.100 510.600 807.900 515.700 ;
        RECT 821.700 513.600 822.900 523.950 ;
        RECT 839.100 522.150 840.900 523.950 ;
        RECT 842.700 519.600 843.900 523.950 ;
        RECT 845.100 522.150 846.900 523.950 ;
        RECT 851.550 523.050 852.450 529.950 ;
        RECT 860.700 526.050 861.900 539.400 ;
        RECT 865.950 528.450 868.050 529.050 ;
        RECT 871.950 528.450 874.050 529.050 ;
        RECT 865.950 527.550 874.050 528.450 ;
        RECT 865.950 526.950 868.050 527.550 ;
        RECT 871.950 526.950 874.050 527.550 ;
        RECT 856.950 523.950 859.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 851.550 521.550 856.050 523.050 ;
        RECT 857.100 522.150 858.900 523.950 ;
        RECT 852.000 520.950 856.050 521.550 ;
        RECT 842.700 518.700 846.300 519.600 ;
        RECT 860.700 518.700 861.900 523.950 ;
        RECT 862.950 522.150 864.750 523.950 ;
        RECT 836.100 515.700 843.900 517.050 ;
        RECT 821.100 510.600 822.900 513.600 ;
        RECT 824.100 510.000 825.900 513.600 ;
        RECT 836.100 510.600 837.900 515.700 ;
        RECT 839.100 510.000 840.900 514.800 ;
        RECT 842.100 510.600 843.900 515.700 ;
        RECT 845.100 516.600 846.300 518.700 ;
        RECT 857.700 517.800 861.900 518.700 ;
        RECT 845.100 510.600 846.900 516.600 ;
        RECT 857.700 510.600 859.500 517.800 ;
        RECT 862.800 510.000 864.600 516.600 ;
        RECT 11.400 500.400 13.200 507.000 ;
        RECT 16.500 499.200 18.300 506.400 ;
        RECT 32.100 501.300 33.900 506.400 ;
        RECT 35.100 502.200 36.900 507.000 ;
        RECT 38.100 501.300 39.900 506.400 ;
        RECT 32.100 499.950 39.900 501.300 ;
        RECT 41.100 500.400 42.900 506.400 ;
        RECT 53.400 500.400 55.200 507.000 ;
        RECT 14.100 498.300 18.300 499.200 ;
        RECT 41.100 498.300 42.300 500.400 ;
        RECT 58.500 499.200 60.300 506.400 ;
        RECT 71.100 501.300 72.900 506.400 ;
        RECT 74.100 502.200 75.900 507.000 ;
        RECT 77.100 501.300 78.900 506.400 ;
        RECT 71.100 499.950 78.900 501.300 ;
        RECT 80.100 500.400 81.900 506.400 ;
        RECT 92.100 503.400 93.900 506.400 ;
        RECT 95.100 503.400 96.900 507.000 ;
        RECT 107.100 503.400 108.900 507.000 ;
        RECT 110.100 503.400 111.900 506.400 ;
        RECT 113.100 503.400 114.900 507.000 ;
        RECT 11.250 493.050 13.050 494.850 ;
        RECT 14.100 493.050 15.300 498.300 ;
        RECT 38.700 497.400 42.300 498.300 ;
        RECT 56.100 498.300 60.300 499.200 ;
        RECT 80.100 498.300 81.300 500.400 ;
        RECT 22.950 495.450 25.050 496.050 ;
        RECT 28.950 495.450 31.050 496.050 ;
        RECT 17.100 493.050 18.900 494.850 ;
        RECT 22.950 494.550 31.050 495.450 ;
        RECT 22.950 493.950 25.050 494.550 ;
        RECT 28.950 493.950 31.050 494.550 ;
        RECT 35.100 493.050 36.900 494.850 ;
        RECT 38.700 493.050 39.900 497.400 ;
        RECT 41.100 493.050 42.900 494.850 ;
        RECT 53.250 493.050 55.050 494.850 ;
        RECT 56.100 493.050 57.300 498.300 ;
        RECT 77.700 497.400 81.300 498.300 ;
        RECT 59.100 493.050 60.900 494.850 ;
        RECT 74.100 493.050 75.900 494.850 ;
        RECT 77.700 493.050 78.900 497.400 ;
        RECT 80.100 493.050 81.900 494.850 ;
        RECT 92.700 493.050 93.900 503.400 ;
        RECT 94.950 498.450 97.050 499.050 ;
        RECT 100.950 498.450 103.050 499.050 ;
        RECT 94.950 497.550 103.050 498.450 ;
        RECT 94.950 496.950 97.050 497.550 ;
        RECT 100.950 496.950 103.050 497.550 ;
        RECT 110.400 493.050 111.300 503.400 ;
        RECT 125.100 500.400 126.900 506.400 ;
        RECT 128.100 501.300 129.900 507.000 ;
        RECT 132.600 500.400 134.400 506.400 ;
        RECT 137.100 501.300 138.900 507.000 ;
        RECT 140.100 500.400 141.900 506.400 ;
        RECT 152.100 503.400 153.900 507.000 ;
        RECT 155.100 503.400 156.900 506.400 ;
        RECT 158.100 503.400 159.900 507.000 ;
        RECT 125.100 499.500 129.900 500.400 ;
        RECT 127.800 498.300 129.900 499.500 ;
        RECT 132.900 498.900 134.100 500.400 ;
        RECT 131.100 496.800 134.100 498.900 ;
        RECT 140.100 498.600 141.300 500.400 ;
        RECT 129.900 493.800 132.000 495.900 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 31.950 490.950 34.050 493.050 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 55.950 490.950 58.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 70.950 490.950 73.050 493.050 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 94.950 490.950 97.050 493.050 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 112.950 490.950 115.050 493.050 ;
        RECT 125.100 490.950 127.200 493.050 ;
        RECT 129.900 492.000 131.700 493.800 ;
        RECT 132.900 491.100 134.100 496.800 ;
        RECT 135.000 497.700 141.300 498.600 ;
        RECT 135.000 495.600 137.100 497.700 ;
        RECT 135.000 493.800 136.800 495.600 ;
        RECT 148.950 495.450 151.050 496.050 ;
        RECT 139.800 493.050 141.600 494.850 ;
        RECT 143.550 494.550 151.050 495.450 ;
        RECT 139.800 492.300 141.900 493.050 ;
        RECT 14.100 477.600 15.300 490.950 ;
        RECT 32.100 489.150 33.900 490.950 ;
        RECT 38.700 483.600 39.900 490.950 ;
        RECT 40.950 486.450 43.050 487.050 ;
        RECT 46.950 486.450 49.050 487.050 ;
        RECT 40.950 485.550 49.050 486.450 ;
        RECT 40.950 484.950 43.050 485.550 ;
        RECT 46.950 484.950 49.050 485.550 ;
        RECT 11.100 471.000 12.900 477.600 ;
        RECT 14.100 471.600 15.900 477.600 ;
        RECT 17.100 471.000 18.900 477.600 ;
        RECT 32.400 471.000 34.200 483.600 ;
        RECT 37.500 482.100 39.900 483.600 ;
        RECT 37.500 471.600 39.300 482.100 ;
        RECT 40.200 479.100 42.000 480.900 ;
        RECT 56.100 477.600 57.300 490.950 ;
        RECT 71.100 489.150 72.900 490.950 ;
        RECT 77.700 483.600 78.900 490.950 ;
        RECT 40.500 471.000 42.300 477.600 ;
        RECT 53.100 471.000 54.900 477.600 ;
        RECT 56.100 471.600 57.900 477.600 ;
        RECT 59.100 471.000 60.900 477.600 ;
        RECT 71.400 471.000 73.200 483.600 ;
        RECT 76.500 482.100 78.900 483.600 ;
        RECT 76.500 471.600 78.300 482.100 ;
        RECT 79.200 479.100 81.000 480.900 ;
        RECT 92.700 477.600 93.900 490.950 ;
        RECT 95.100 489.150 96.900 490.950 ;
        RECT 107.250 489.150 109.050 490.950 ;
        RECT 110.400 483.600 111.300 490.950 ;
        RECT 113.100 489.150 114.900 490.950 ;
        RECT 125.400 489.150 127.200 490.950 ;
        RECT 131.700 490.200 134.100 491.100 ;
        RECT 135.000 490.950 141.900 492.300 ;
        RECT 135.000 490.500 136.800 490.950 ;
        RECT 131.700 490.050 133.200 490.200 ;
        RECT 131.100 487.950 133.200 490.050 ;
        RECT 132.300 486.000 133.200 487.950 ;
        RECT 134.100 487.500 138.000 489.300 ;
        RECT 134.100 487.200 136.200 487.500 ;
        RECT 143.550 487.050 144.450 494.550 ;
        RECT 148.950 493.950 151.050 494.550 ;
        RECT 155.700 493.050 156.600 503.400 ;
        RECT 174.600 502.200 176.400 506.400 ;
        RECT 157.950 501.450 160.050 502.050 ;
        RECT 169.950 501.450 172.050 502.050 ;
        RECT 157.950 500.550 172.050 501.450 ;
        RECT 157.950 499.950 160.050 500.550 ;
        RECT 169.950 499.950 172.050 500.550 ;
        RECT 173.700 500.400 176.400 502.200 ;
        RECT 177.600 500.400 179.400 507.000 ;
        RECT 173.700 493.050 174.600 500.400 ;
        RECT 175.500 498.600 177.300 499.500 ;
        RECT 182.100 498.600 183.900 506.400 ;
        RECT 184.950 504.450 187.050 505.050 ;
        RECT 190.950 504.450 193.050 505.050 ;
        RECT 184.950 503.550 193.050 504.450 ;
        RECT 184.950 502.950 187.050 503.550 ;
        RECT 190.950 502.950 193.050 503.550 ;
        RECT 194.100 501.300 195.900 506.400 ;
        RECT 197.100 502.200 198.900 507.000 ;
        RECT 200.100 501.300 201.900 506.400 ;
        RECT 194.100 499.950 201.900 501.300 ;
        RECT 203.100 500.400 204.900 506.400 ;
        RECT 207.150 502.200 208.950 506.400 ;
        RECT 206.550 500.400 208.950 502.200 ;
        RECT 210.150 500.400 211.950 507.000 ;
        RECT 214.950 504.300 216.750 506.400 ;
        RECT 213.150 503.400 216.750 504.300 ;
        RECT 219.450 503.400 221.250 507.000 ;
        RECT 222.750 503.400 224.550 506.400 ;
        RECT 225.750 503.400 227.550 507.000 ;
        RECT 230.250 503.400 232.050 506.400 ;
        RECT 212.850 502.800 216.750 503.400 ;
        RECT 212.850 501.300 214.950 502.800 ;
        RECT 222.750 502.500 223.800 503.400 ;
        RECT 175.500 497.700 183.900 498.600 ;
        RECT 203.100 498.300 204.300 500.400 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 157.950 490.950 160.050 493.050 ;
        RECT 173.100 490.950 175.200 493.050 ;
        RECT 176.400 490.950 178.500 493.050 ;
        RECT 152.100 489.150 153.900 490.950 ;
        RECT 132.300 484.950 133.800 486.000 ;
        RECT 127.800 483.600 129.900 484.500 ;
        RECT 79.500 471.000 81.300 477.600 ;
        RECT 92.100 471.600 93.900 477.600 ;
        RECT 95.100 471.000 96.900 477.600 ;
        RECT 107.100 471.000 108.900 483.600 ;
        RECT 110.400 482.400 114.000 483.600 ;
        RECT 112.200 471.600 114.000 482.400 ;
        RECT 125.100 482.400 129.900 483.600 ;
        RECT 132.600 483.600 133.800 484.950 ;
        RECT 137.400 483.600 139.500 485.700 ;
        RECT 142.950 484.950 145.050 487.050 ;
        RECT 155.700 483.600 156.600 490.950 ;
        RECT 157.950 489.150 159.750 490.950 ;
        RECT 173.700 483.600 174.600 490.950 ;
        RECT 177.000 489.150 178.800 490.950 ;
        RECT 125.100 471.600 126.900 482.400 ;
        RECT 128.100 471.000 129.900 481.500 ;
        RECT 132.600 471.600 134.400 483.600 ;
        RECT 137.400 482.700 141.900 483.600 ;
        RECT 137.100 471.000 138.900 481.500 ;
        RECT 140.100 471.600 141.900 482.700 ;
        RECT 153.000 482.400 156.600 483.600 ;
        RECT 153.000 471.600 154.800 482.400 ;
        RECT 158.100 471.000 159.900 483.600 ;
        RECT 173.100 471.600 174.900 483.600 ;
        RECT 176.100 471.000 177.900 483.000 ;
        RECT 180.000 477.600 180.900 497.700 ;
        RECT 200.700 497.400 204.300 498.300 ;
        RECT 181.950 493.050 183.750 494.850 ;
        RECT 197.100 493.050 198.900 494.850 ;
        RECT 200.700 493.050 201.900 497.400 ;
        RECT 203.100 493.050 204.900 494.850 ;
        RECT 181.800 490.950 183.900 493.050 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 199.950 490.950 202.050 493.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 194.100 489.150 195.900 490.950 ;
        RECT 200.700 483.600 201.900 490.950 ;
        RECT 179.100 471.600 180.900 477.600 ;
        RECT 182.100 471.000 183.900 477.600 ;
        RECT 194.400 471.000 196.200 483.600 ;
        RECT 199.500 482.100 201.900 483.600 ;
        RECT 206.550 485.700 207.450 500.400 ;
        RECT 215.850 499.800 217.650 501.600 ;
        RECT 218.850 501.450 223.800 502.500 ;
        RECT 218.850 500.700 220.650 501.450 ;
        RECT 230.250 501.300 232.650 503.400 ;
        RECT 235.350 500.400 237.150 507.000 ;
        RECT 238.650 500.400 240.450 506.400 ;
        RECT 215.850 498.000 216.900 499.800 ;
        RECT 226.050 498.000 227.850 498.600 ;
        RECT 215.850 496.800 227.850 498.000 ;
        RECT 208.950 495.600 216.900 496.800 ;
        RECT 208.950 493.050 210.750 495.600 ;
        RECT 215.100 495.000 216.900 495.600 ;
        RECT 212.100 493.800 213.900 494.400 ;
        RECT 208.950 490.950 211.050 493.050 ;
        RECT 212.100 492.600 220.200 493.800 ;
        RECT 218.100 490.950 220.200 492.600 ;
        RECT 216.450 485.700 218.250 486.000 ;
        RECT 206.550 485.100 218.250 485.700 ;
        RECT 206.550 484.500 224.850 485.100 ;
        RECT 206.550 483.600 207.450 484.500 ;
        RECT 216.450 484.200 224.850 484.500 ;
        RECT 199.500 471.600 201.300 482.100 ;
        RECT 206.550 481.800 208.950 483.600 ;
        RECT 202.200 479.100 204.000 480.900 ;
        RECT 202.500 471.000 204.300 477.600 ;
        RECT 207.150 471.600 208.950 481.800 ;
        RECT 210.150 471.000 211.950 483.600 ;
        RECT 221.250 482.700 223.050 483.300 ;
        RECT 215.250 481.500 223.050 482.700 ;
        RECT 223.950 482.100 224.850 484.200 ;
        RECT 226.950 484.200 227.850 496.800 ;
        RECT 239.250 493.050 240.450 500.400 ;
        RECT 251.100 500.400 252.900 506.400 ;
        RECT 254.100 501.300 255.900 507.000 ;
        RECT 258.300 501.000 260.100 506.400 ;
        RECT 262.800 501.300 264.600 507.000 ;
        RECT 251.100 499.500 252.600 500.400 ;
        RECT 251.100 498.000 255.600 499.500 ;
        RECT 253.500 497.400 255.600 498.000 ;
        RECT 259.200 498.900 260.100 501.000 ;
        RECT 266.100 500.400 267.900 506.400 ;
        RECT 263.400 499.500 267.900 500.400 ;
        RECT 281.100 500.400 282.900 506.400 ;
        RECT 284.100 501.300 285.900 507.000 ;
        RECT 288.600 500.400 290.400 506.400 ;
        RECT 293.100 501.300 294.900 507.000 ;
        RECT 296.100 500.400 297.900 506.400 ;
        RECT 299.550 500.400 301.350 506.400 ;
        RECT 302.850 500.400 304.650 507.000 ;
        RECT 307.950 503.400 309.750 506.400 ;
        RECT 312.450 503.400 314.250 507.000 ;
        RECT 315.450 503.400 317.250 506.400 ;
        RECT 318.750 503.400 320.550 507.000 ;
        RECT 323.250 504.300 325.050 506.400 ;
        RECT 323.250 503.400 326.850 504.300 ;
        RECT 307.350 501.300 309.750 503.400 ;
        RECT 316.200 502.500 317.250 503.400 ;
        RECT 323.250 502.800 327.150 503.400 ;
        RECT 316.200 501.450 321.150 502.500 ;
        RECT 319.350 500.700 321.150 501.450 ;
        RECT 281.100 499.500 285.900 500.400 ;
        RECT 256.500 495.900 258.300 497.700 ;
        RECT 259.200 496.800 262.200 498.900 ;
        RECT 263.400 497.100 265.500 499.500 ;
        RECT 283.800 498.300 285.900 499.500 ;
        RECT 288.900 498.900 290.100 500.400 ;
        RECT 287.100 496.800 290.100 498.900 ;
        RECT 296.100 498.600 297.300 500.400 ;
        RECT 255.900 495.000 258.000 495.900 ;
        RECT 251.400 493.800 258.000 495.000 ;
        RECT 251.400 493.200 253.200 493.800 ;
        RECT 234.150 491.250 240.450 493.050 ;
        RECT 235.950 490.950 240.450 491.250 ;
        RECT 251.100 490.950 253.200 493.200 ;
        RECT 230.550 488.100 232.650 488.400 ;
        RECT 236.550 488.100 238.350 488.250 ;
        RECT 230.550 486.900 238.350 488.100 ;
        RECT 230.550 486.300 232.650 486.900 ;
        RECT 236.550 486.450 238.350 486.900 ;
        RECT 226.950 483.300 231.750 484.200 ;
        RECT 239.250 483.600 240.450 490.950 ;
        RECT 255.900 490.800 258.000 492.900 ;
        RECT 255.900 489.000 257.700 490.800 ;
        RECT 259.200 490.050 260.100 496.800 ;
        RECT 261.000 492.900 263.100 495.000 ;
        RECT 285.900 493.800 288.000 495.900 ;
        RECT 261.000 491.100 262.800 492.900 ;
        RECT 265.800 490.950 267.900 493.050 ;
        RECT 281.100 490.950 283.200 493.050 ;
        RECT 285.900 492.000 287.700 493.800 ;
        RECT 288.900 491.100 290.100 496.800 ;
        RECT 291.000 497.700 297.300 498.600 ;
        RECT 291.000 495.600 293.100 497.700 ;
        RECT 291.000 493.800 292.800 495.600 ;
        RECT 295.800 493.050 297.600 494.850 ;
        RECT 299.550 493.050 300.750 500.400 ;
        RECT 322.350 499.800 324.150 501.600 ;
        RECT 325.050 501.300 327.150 502.800 ;
        RECT 328.050 500.400 329.850 507.000 ;
        RECT 331.050 502.200 332.850 506.400 ;
        RECT 331.050 500.400 333.450 502.200 ;
        RECT 344.100 500.400 345.900 507.000 ;
        RECT 312.150 498.000 313.950 498.600 ;
        RECT 323.100 498.000 324.150 499.800 ;
        RECT 312.150 496.800 324.150 498.000 ;
        RECT 295.800 492.300 297.900 493.050 ;
        RECT 259.200 488.700 262.200 490.050 ;
        RECT 265.800 489.150 267.600 490.950 ;
        RECT 281.400 489.150 283.200 490.950 ;
        RECT 287.700 490.200 290.100 491.100 ;
        RECT 291.000 490.950 297.900 492.300 ;
        RECT 299.550 491.250 305.850 493.050 ;
        RECT 299.550 490.950 304.050 491.250 ;
        RECT 291.000 490.500 292.800 490.950 ;
        RECT 287.700 490.050 289.200 490.200 ;
        RECT 260.100 487.950 262.200 488.700 ;
        RECT 287.100 487.950 289.200 490.050 ;
        RECT 257.400 485.700 259.200 487.500 ;
        RECT 253.800 484.800 259.200 485.700 ;
        RECT 253.800 483.900 255.900 484.800 ;
        RECT 230.550 482.400 231.750 483.300 ;
        RECT 227.850 482.100 229.650 482.400 ;
        RECT 215.250 480.600 217.350 481.500 ;
        RECT 223.950 481.200 229.650 482.100 ;
        RECT 227.850 480.600 229.650 481.200 ;
        RECT 230.550 480.600 233.550 482.400 ;
        RECT 215.550 471.600 217.350 480.600 ;
        RECT 219.450 479.550 221.250 480.300 ;
        RECT 224.250 479.550 226.050 480.300 ;
        RECT 219.450 478.500 226.050 479.550 ;
        RECT 220.350 471.000 222.150 477.600 ;
        RECT 223.350 471.600 225.150 478.500 ;
        RECT 230.550 477.600 232.650 479.700 ;
        RECT 226.350 471.000 228.150 477.600 ;
        RECT 230.850 471.600 232.650 477.600 ;
        RECT 235.650 471.000 237.450 483.600 ;
        RECT 238.650 471.600 240.450 483.600 ;
        RECT 251.100 482.700 255.900 483.900 ;
        RECT 260.700 483.600 261.900 487.950 ;
        RECT 288.300 486.000 289.200 487.950 ;
        RECT 290.100 487.500 294.000 489.300 ;
        RECT 290.100 487.200 292.200 487.500 ;
        RECT 288.300 484.950 289.800 486.000 ;
        RECT 258.600 482.700 261.900 483.600 ;
        RECT 262.800 483.600 264.900 484.500 ;
        RECT 283.800 483.600 285.900 484.500 ;
        RECT 251.100 471.600 252.900 482.700 ;
        RECT 254.100 471.000 255.900 481.500 ;
        RECT 258.600 471.600 260.400 482.700 ;
        RECT 262.800 482.400 267.900 483.600 ;
        RECT 262.800 471.000 264.900 481.500 ;
        RECT 266.100 471.600 267.900 482.400 ;
        RECT 281.100 482.400 285.900 483.600 ;
        RECT 288.600 483.600 289.800 484.950 ;
        RECT 293.400 483.600 295.500 485.700 ;
        RECT 299.550 483.600 300.750 490.950 ;
        RECT 301.650 488.100 303.450 488.250 ;
        RECT 307.350 488.100 309.450 488.400 ;
        RECT 301.650 486.900 309.450 488.100 ;
        RECT 301.650 486.450 303.450 486.900 ;
        RECT 307.350 486.300 309.450 486.900 ;
        RECT 312.150 484.200 313.050 496.800 ;
        RECT 323.100 495.600 331.050 496.800 ;
        RECT 323.100 495.000 324.900 495.600 ;
        RECT 326.100 493.800 327.900 494.400 ;
        RECT 319.800 492.600 327.900 493.800 ;
        RECT 329.250 493.050 331.050 495.600 ;
        RECT 319.800 490.950 321.900 492.600 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 321.750 485.700 323.550 486.000 ;
        RECT 332.550 485.700 333.450 500.400 ;
        RECT 347.100 499.500 348.900 506.400 ;
        RECT 350.100 500.400 351.900 507.000 ;
        RECT 353.100 499.500 354.900 506.400 ;
        RECT 356.100 500.400 357.900 507.000 ;
        RECT 359.100 499.500 360.900 506.400 ;
        RECT 362.100 500.400 363.900 507.000 ;
        RECT 365.100 499.500 366.900 506.400 ;
        RECT 368.100 500.400 369.900 507.000 ;
        RECT 371.550 500.400 373.350 506.400 ;
        RECT 374.850 500.400 376.650 507.000 ;
        RECT 379.950 503.400 381.750 506.400 ;
        RECT 384.450 503.400 386.250 507.000 ;
        RECT 387.450 503.400 389.250 506.400 ;
        RECT 390.750 503.400 392.550 507.000 ;
        RECT 395.250 504.300 397.050 506.400 ;
        RECT 395.250 503.400 398.850 504.300 ;
        RECT 379.350 501.300 381.750 503.400 ;
        RECT 388.200 502.500 389.250 503.400 ;
        RECT 395.250 502.800 399.150 503.400 ;
        RECT 388.200 501.450 393.150 502.500 ;
        RECT 391.350 500.700 393.150 501.450 ;
        RECT 347.100 498.300 351.000 499.500 ;
        RECT 353.100 498.300 357.000 499.500 ;
        RECT 359.100 498.300 363.000 499.500 ;
        RECT 365.100 498.300 367.950 499.500 ;
        RECT 349.800 497.400 351.000 498.300 ;
        RECT 355.800 497.400 357.000 498.300 ;
        RECT 361.800 497.400 363.000 498.300 ;
        RECT 349.800 496.200 354.000 497.400 ;
        RECT 346.800 493.050 348.600 494.850 ;
        RECT 346.800 490.950 348.900 493.050 ;
        RECT 349.800 485.700 351.000 496.200 ;
        RECT 352.200 495.600 354.000 496.200 ;
        RECT 355.800 496.200 360.000 497.400 ;
        RECT 355.800 485.700 357.000 496.200 ;
        RECT 358.200 495.600 360.000 496.200 ;
        RECT 361.800 496.200 366.000 497.400 ;
        RECT 361.800 485.700 363.000 496.200 ;
        RECT 364.200 495.600 366.000 496.200 ;
        RECT 366.900 493.050 367.950 498.300 ;
        RECT 364.800 490.950 367.950 493.050 ;
        RECT 366.900 485.700 367.950 490.950 ;
        RECT 321.750 485.100 333.450 485.700 ;
        RECT 281.100 471.600 282.900 482.400 ;
        RECT 284.100 471.000 285.900 481.500 ;
        RECT 288.600 471.600 290.400 483.600 ;
        RECT 293.400 482.700 297.900 483.600 ;
        RECT 293.100 471.000 294.900 481.500 ;
        RECT 296.100 471.600 297.900 482.700 ;
        RECT 299.550 471.600 301.350 483.600 ;
        RECT 302.550 471.000 304.350 483.600 ;
        RECT 308.250 483.300 313.050 484.200 ;
        RECT 315.150 484.500 333.450 485.100 ;
        RECT 315.150 484.200 323.550 484.500 ;
        RECT 308.250 482.400 309.450 483.300 ;
        RECT 306.450 480.600 309.450 482.400 ;
        RECT 310.350 482.100 312.150 482.400 ;
        RECT 315.150 482.100 316.050 484.200 ;
        RECT 332.550 483.600 333.450 484.500 ;
        RECT 347.100 484.500 351.000 485.700 ;
        RECT 353.100 484.500 357.000 485.700 ;
        RECT 359.100 484.500 363.000 485.700 ;
        RECT 365.100 484.500 367.950 485.700 ;
        RECT 371.550 493.050 372.750 500.400 ;
        RECT 394.350 499.800 396.150 501.600 ;
        RECT 397.050 501.300 399.150 502.800 ;
        RECT 400.050 500.400 401.850 507.000 ;
        RECT 403.050 502.200 404.850 506.400 ;
        RECT 403.050 500.400 405.450 502.200 ;
        RECT 416.100 500.400 417.900 506.400 ;
        RECT 384.150 498.000 385.950 498.600 ;
        RECT 395.100 498.000 396.150 499.800 ;
        RECT 384.150 496.800 396.150 498.000 ;
        RECT 371.550 491.250 377.850 493.050 ;
        RECT 371.550 490.950 376.050 491.250 ;
        RECT 310.350 481.200 316.050 482.100 ;
        RECT 316.950 482.700 318.750 483.300 ;
        RECT 316.950 481.500 324.750 482.700 ;
        RECT 310.350 480.600 312.150 481.200 ;
        RECT 322.650 480.600 324.750 481.500 ;
        RECT 307.350 477.600 309.450 479.700 ;
        RECT 313.950 479.550 315.750 480.300 ;
        RECT 318.750 479.550 320.550 480.300 ;
        RECT 313.950 478.500 320.550 479.550 ;
        RECT 307.350 471.600 309.150 477.600 ;
        RECT 311.850 471.000 313.650 477.600 ;
        RECT 314.850 471.600 316.650 478.500 ;
        RECT 317.850 471.000 319.650 477.600 ;
        RECT 322.650 471.600 324.450 480.600 ;
        RECT 328.050 471.000 329.850 483.600 ;
        RECT 331.050 481.800 333.450 483.600 ;
        RECT 331.050 471.600 332.850 481.800 ;
        RECT 344.100 471.000 345.900 483.600 ;
        RECT 347.100 471.600 348.900 484.500 ;
        RECT 350.100 471.000 351.900 483.600 ;
        RECT 353.100 471.600 354.900 484.500 ;
        RECT 356.100 471.000 357.900 483.600 ;
        RECT 359.100 471.600 360.900 484.500 ;
        RECT 362.100 471.000 363.900 483.600 ;
        RECT 365.100 471.600 366.900 484.500 ;
        RECT 371.550 483.600 372.750 490.950 ;
        RECT 373.650 488.100 375.450 488.250 ;
        RECT 379.350 488.100 381.450 488.400 ;
        RECT 373.650 486.900 381.450 488.100 ;
        RECT 373.650 486.450 375.450 486.900 ;
        RECT 379.350 486.300 381.450 486.900 ;
        RECT 384.150 484.200 385.050 496.800 ;
        RECT 395.100 495.600 403.050 496.800 ;
        RECT 395.100 495.000 396.900 495.600 ;
        RECT 398.100 493.800 399.900 494.400 ;
        RECT 391.800 492.600 399.900 493.800 ;
        RECT 401.250 493.050 403.050 495.600 ;
        RECT 391.800 490.950 393.900 492.600 ;
        RECT 400.950 490.950 403.050 493.050 ;
        RECT 393.750 485.700 395.550 486.000 ;
        RECT 404.550 485.700 405.450 500.400 ;
        RECT 416.700 498.300 417.900 500.400 ;
        RECT 419.100 501.300 420.900 506.400 ;
        RECT 422.100 502.200 423.900 507.000 ;
        RECT 425.100 501.300 426.900 506.400 ;
        RECT 419.100 499.950 426.900 501.300 ;
        RECT 437.100 500.400 438.900 506.400 ;
        RECT 437.700 498.300 438.900 500.400 ;
        RECT 440.100 501.300 441.900 506.400 ;
        RECT 443.100 502.200 444.900 507.000 ;
        RECT 446.100 501.300 447.900 506.400 ;
        RECT 440.100 499.950 447.900 501.300 ;
        RECT 449.550 500.400 451.350 506.400 ;
        RECT 452.850 500.400 454.650 507.000 ;
        RECT 457.950 503.400 459.750 506.400 ;
        RECT 462.450 503.400 464.250 507.000 ;
        RECT 465.450 503.400 467.250 506.400 ;
        RECT 468.750 503.400 470.550 507.000 ;
        RECT 473.250 504.300 475.050 506.400 ;
        RECT 473.250 503.400 476.850 504.300 ;
        RECT 457.350 501.300 459.750 503.400 ;
        RECT 466.200 502.500 467.250 503.400 ;
        RECT 473.250 502.800 477.150 503.400 ;
        RECT 466.200 501.450 471.150 502.500 ;
        RECT 469.350 500.700 471.150 501.450 ;
        RECT 416.700 497.400 420.300 498.300 ;
        RECT 437.700 497.400 441.300 498.300 ;
        RECT 416.100 493.050 417.900 494.850 ;
        RECT 419.100 493.050 420.300 497.400 ;
        RECT 422.100 493.050 423.900 494.850 ;
        RECT 437.100 493.050 438.900 494.850 ;
        RECT 440.100 493.050 441.300 497.400 ;
        RECT 443.100 493.050 444.900 494.850 ;
        RECT 449.550 493.050 450.750 500.400 ;
        RECT 472.350 499.800 474.150 501.600 ;
        RECT 475.050 501.300 477.150 502.800 ;
        RECT 478.050 500.400 479.850 507.000 ;
        RECT 481.050 502.200 482.850 506.400 ;
        RECT 481.050 500.400 483.450 502.200 ;
        RECT 462.150 498.000 463.950 498.600 ;
        RECT 473.100 498.000 474.150 499.800 ;
        RECT 462.150 496.800 474.150 498.000 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 445.950 490.950 448.050 493.050 ;
        RECT 449.550 491.250 455.850 493.050 ;
        RECT 449.550 490.950 454.050 491.250 ;
        RECT 393.750 485.100 405.450 485.700 ;
        RECT 368.100 471.000 369.900 483.600 ;
        RECT 371.550 471.600 373.350 483.600 ;
        RECT 374.550 471.000 376.350 483.600 ;
        RECT 380.250 483.300 385.050 484.200 ;
        RECT 387.150 484.500 405.450 485.100 ;
        RECT 387.150 484.200 395.550 484.500 ;
        RECT 380.250 482.400 381.450 483.300 ;
        RECT 378.450 480.600 381.450 482.400 ;
        RECT 382.350 482.100 384.150 482.400 ;
        RECT 387.150 482.100 388.050 484.200 ;
        RECT 404.550 483.600 405.450 484.500 ;
        RECT 382.350 481.200 388.050 482.100 ;
        RECT 388.950 482.700 390.750 483.300 ;
        RECT 388.950 481.500 396.750 482.700 ;
        RECT 382.350 480.600 384.150 481.200 ;
        RECT 394.650 480.600 396.750 481.500 ;
        RECT 379.350 477.600 381.450 479.700 ;
        RECT 385.950 479.550 387.750 480.300 ;
        RECT 390.750 479.550 392.550 480.300 ;
        RECT 385.950 478.500 392.550 479.550 ;
        RECT 379.350 471.600 381.150 477.600 ;
        RECT 383.850 471.000 385.650 477.600 ;
        RECT 386.850 471.600 388.650 478.500 ;
        RECT 389.850 471.000 391.650 477.600 ;
        RECT 394.650 471.600 396.450 480.600 ;
        RECT 400.050 471.000 401.850 483.600 ;
        RECT 403.050 481.800 405.450 483.600 ;
        RECT 419.100 483.600 420.300 490.950 ;
        RECT 425.100 489.150 426.900 490.950 ;
        RECT 440.100 483.600 441.300 490.950 ;
        RECT 446.100 489.150 447.900 490.950 ;
        RECT 449.550 483.600 450.750 490.950 ;
        RECT 451.650 488.100 453.450 488.250 ;
        RECT 457.350 488.100 459.450 488.400 ;
        RECT 451.650 486.900 459.450 488.100 ;
        RECT 451.650 486.450 453.450 486.900 ;
        RECT 457.350 486.300 459.450 486.900 ;
        RECT 462.150 484.200 463.050 496.800 ;
        RECT 473.100 495.600 481.050 496.800 ;
        RECT 473.100 495.000 474.900 495.600 ;
        RECT 476.100 493.800 477.900 494.400 ;
        RECT 469.800 492.600 477.900 493.800 ;
        RECT 479.250 493.050 481.050 495.600 ;
        RECT 469.800 490.950 471.900 492.600 ;
        RECT 478.950 490.950 481.050 493.050 ;
        RECT 471.750 485.700 473.550 486.000 ;
        RECT 482.550 485.700 483.450 500.400 ;
        RECT 494.100 501.300 495.900 506.400 ;
        RECT 497.100 502.200 498.900 507.000 ;
        RECT 500.100 501.300 501.900 506.400 ;
        RECT 494.100 499.950 501.900 501.300 ;
        RECT 503.100 500.400 504.900 506.400 ;
        RECT 515.100 500.400 516.900 506.400 ;
        RECT 503.100 498.300 504.300 500.400 ;
        RECT 500.700 497.400 504.300 498.300 ;
        RECT 515.700 498.300 516.900 500.400 ;
        RECT 518.100 501.300 519.900 506.400 ;
        RECT 521.100 502.200 522.900 507.000 ;
        RECT 524.100 501.300 525.900 506.400 ;
        RECT 518.100 499.950 525.900 501.300 ;
        RECT 536.100 500.400 537.900 507.000 ;
        RECT 539.100 499.500 540.900 506.400 ;
        RECT 542.100 500.400 543.900 507.000 ;
        RECT 545.100 499.500 546.900 506.400 ;
        RECT 548.100 500.400 549.900 507.000 ;
        RECT 551.100 499.500 552.900 506.400 ;
        RECT 554.100 500.400 555.900 507.000 ;
        RECT 557.100 499.500 558.900 506.400 ;
        RECT 560.100 500.400 561.900 507.000 ;
        RECT 563.550 500.400 565.350 506.400 ;
        RECT 566.850 500.400 568.650 507.000 ;
        RECT 571.950 503.400 573.750 506.400 ;
        RECT 576.450 503.400 578.250 507.000 ;
        RECT 579.450 503.400 581.250 506.400 ;
        RECT 582.750 503.400 584.550 507.000 ;
        RECT 587.250 504.300 589.050 506.400 ;
        RECT 587.250 503.400 590.850 504.300 ;
        RECT 571.350 501.300 573.750 503.400 ;
        RECT 580.200 502.500 581.250 503.400 ;
        RECT 587.250 502.800 591.150 503.400 ;
        RECT 580.200 501.450 585.150 502.500 ;
        RECT 583.350 500.700 585.150 501.450 ;
        RECT 538.050 498.300 540.900 499.500 ;
        RECT 543.000 498.300 546.900 499.500 ;
        RECT 549.000 498.300 552.900 499.500 ;
        RECT 555.000 498.300 558.900 499.500 ;
        RECT 515.700 497.400 519.300 498.300 ;
        RECT 497.100 493.050 498.900 494.850 ;
        RECT 500.700 493.050 501.900 497.400 ;
        RECT 503.100 493.050 504.900 494.850 ;
        RECT 515.100 493.050 516.900 494.850 ;
        RECT 518.100 493.050 519.300 497.400 ;
        RECT 521.100 493.050 522.900 494.850 ;
        RECT 538.050 493.050 539.100 498.300 ;
        RECT 543.000 497.400 544.200 498.300 ;
        RECT 549.000 497.400 550.200 498.300 ;
        RECT 555.000 497.400 556.200 498.300 ;
        RECT 540.000 496.200 544.200 497.400 ;
        RECT 540.000 495.600 541.800 496.200 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 499.950 490.950 502.050 493.050 ;
        RECT 502.950 490.950 505.050 493.050 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 520.950 490.950 523.050 493.050 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 538.050 490.950 541.200 493.050 ;
        RECT 494.100 489.150 495.900 490.950 ;
        RECT 471.750 485.100 483.450 485.700 ;
        RECT 419.100 482.100 421.500 483.600 ;
        RECT 403.050 471.600 404.850 481.800 ;
        RECT 417.000 479.100 418.800 480.900 ;
        RECT 416.700 471.000 418.500 477.600 ;
        RECT 419.700 471.600 421.500 482.100 ;
        RECT 424.800 471.000 426.600 483.600 ;
        RECT 440.100 482.100 442.500 483.600 ;
        RECT 438.000 479.100 439.800 480.900 ;
        RECT 437.700 471.000 439.500 477.600 ;
        RECT 440.700 471.600 442.500 482.100 ;
        RECT 445.800 471.000 447.600 483.600 ;
        RECT 449.550 471.600 451.350 483.600 ;
        RECT 452.550 471.000 454.350 483.600 ;
        RECT 458.250 483.300 463.050 484.200 ;
        RECT 465.150 484.500 483.450 485.100 ;
        RECT 484.950 486.450 487.050 487.050 ;
        RECT 496.950 486.450 499.050 487.050 ;
        RECT 484.950 485.550 499.050 486.450 ;
        RECT 484.950 484.950 487.050 485.550 ;
        RECT 496.950 484.950 499.050 485.550 ;
        RECT 465.150 484.200 473.550 484.500 ;
        RECT 458.250 482.400 459.450 483.300 ;
        RECT 456.450 480.600 459.450 482.400 ;
        RECT 460.350 482.100 462.150 482.400 ;
        RECT 465.150 482.100 466.050 484.200 ;
        RECT 482.550 483.600 483.450 484.500 ;
        RECT 500.700 483.600 501.900 490.950 ;
        RECT 460.350 481.200 466.050 482.100 ;
        RECT 466.950 482.700 468.750 483.300 ;
        RECT 466.950 481.500 474.750 482.700 ;
        RECT 460.350 480.600 462.150 481.200 ;
        RECT 472.650 480.600 474.750 481.500 ;
        RECT 457.350 477.600 459.450 479.700 ;
        RECT 463.950 479.550 465.750 480.300 ;
        RECT 468.750 479.550 470.550 480.300 ;
        RECT 463.950 478.500 470.550 479.550 ;
        RECT 457.350 471.600 459.150 477.600 ;
        RECT 461.850 471.000 463.650 477.600 ;
        RECT 464.850 471.600 466.650 478.500 ;
        RECT 467.850 471.000 469.650 477.600 ;
        RECT 472.650 471.600 474.450 480.600 ;
        RECT 478.050 471.000 479.850 483.600 ;
        RECT 481.050 481.800 483.450 483.600 ;
        RECT 481.050 471.600 482.850 481.800 ;
        RECT 494.400 471.000 496.200 483.600 ;
        RECT 499.500 482.100 501.900 483.600 ;
        RECT 518.100 483.600 519.300 490.950 ;
        RECT 524.100 489.150 525.900 490.950 ;
        RECT 538.050 485.700 539.100 490.950 ;
        RECT 543.000 485.700 544.200 496.200 ;
        RECT 546.000 496.200 550.200 497.400 ;
        RECT 546.000 495.600 547.800 496.200 ;
        RECT 549.000 485.700 550.200 496.200 ;
        RECT 552.000 496.200 556.200 497.400 ;
        RECT 552.000 495.600 553.800 496.200 ;
        RECT 555.000 485.700 556.200 496.200 ;
        RECT 557.400 493.050 559.200 494.850 ;
        RECT 557.100 490.950 559.200 493.050 ;
        RECT 563.550 493.050 564.750 500.400 ;
        RECT 586.350 499.800 588.150 501.600 ;
        RECT 589.050 501.300 591.150 502.800 ;
        RECT 592.050 500.400 593.850 507.000 ;
        RECT 595.050 502.200 596.850 506.400 ;
        RECT 595.050 500.400 597.450 502.200 ;
        RECT 576.150 498.000 577.950 498.600 ;
        RECT 587.100 498.000 588.150 499.800 ;
        RECT 576.150 496.800 588.150 498.000 ;
        RECT 563.550 491.250 569.850 493.050 ;
        RECT 563.550 490.950 568.050 491.250 ;
        RECT 538.050 484.500 540.900 485.700 ;
        RECT 543.000 484.500 546.900 485.700 ;
        RECT 549.000 484.500 552.900 485.700 ;
        RECT 555.000 484.500 558.900 485.700 ;
        RECT 518.100 482.100 520.500 483.600 ;
        RECT 499.500 471.600 501.300 482.100 ;
        RECT 502.200 479.100 504.000 480.900 ;
        RECT 516.000 479.100 517.800 480.900 ;
        RECT 502.500 471.000 504.300 477.600 ;
        RECT 515.700 471.000 517.500 477.600 ;
        RECT 518.700 471.600 520.500 482.100 ;
        RECT 523.800 471.000 525.600 483.600 ;
        RECT 536.100 471.000 537.900 483.600 ;
        RECT 539.100 471.600 540.900 484.500 ;
        RECT 542.100 471.000 543.900 483.600 ;
        RECT 545.100 471.600 546.900 484.500 ;
        RECT 548.100 471.000 549.900 483.600 ;
        RECT 551.100 471.600 552.900 484.500 ;
        RECT 554.100 471.000 555.900 483.600 ;
        RECT 557.100 471.600 558.900 484.500 ;
        RECT 563.550 483.600 564.750 490.950 ;
        RECT 565.650 488.100 567.450 488.250 ;
        RECT 571.350 488.100 573.450 488.400 ;
        RECT 565.650 486.900 573.450 488.100 ;
        RECT 565.650 486.450 567.450 486.900 ;
        RECT 571.350 486.300 573.450 486.900 ;
        RECT 576.150 484.200 577.050 496.800 ;
        RECT 587.100 495.600 595.050 496.800 ;
        RECT 587.100 495.000 588.900 495.600 ;
        RECT 590.100 493.800 591.900 494.400 ;
        RECT 583.800 492.600 591.900 493.800 ;
        RECT 593.250 493.050 595.050 495.600 ;
        RECT 583.800 490.950 585.900 492.600 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 585.750 485.700 587.550 486.000 ;
        RECT 596.550 485.700 597.450 500.400 ;
        RECT 608.100 500.400 609.900 506.400 ;
        RECT 611.100 501.300 612.900 507.000 ;
        RECT 615.600 500.400 617.400 506.400 ;
        RECT 620.100 501.300 621.900 507.000 ;
        RECT 623.100 500.400 624.900 506.400 ;
        RECT 635.100 500.400 636.900 506.400 ;
        RECT 638.100 501.300 639.900 507.000 ;
        RECT 642.600 500.400 644.400 506.400 ;
        RECT 647.100 501.300 648.900 507.000 ;
        RECT 650.100 500.400 651.900 506.400 ;
        RECT 663.000 500.400 664.800 507.000 ;
        RECT 667.500 501.600 669.300 506.400 ;
        RECT 670.500 503.400 672.300 507.000 ;
        RECT 683.100 503.400 684.900 506.400 ;
        RECT 686.100 503.400 687.900 507.000 ;
        RECT 698.100 503.400 699.900 506.400 ;
        RECT 701.100 503.400 702.900 507.000 ;
        RECT 667.500 500.400 672.600 501.600 ;
        RECT 608.100 499.500 612.900 500.400 ;
        RECT 610.800 498.300 612.900 499.500 ;
        RECT 615.900 498.900 617.100 500.400 ;
        RECT 614.100 496.800 617.100 498.900 ;
        RECT 623.100 498.600 624.300 500.400 ;
        RECT 612.900 493.800 615.000 495.900 ;
        RECT 608.100 490.950 610.200 493.050 ;
        RECT 612.900 492.000 614.700 493.800 ;
        RECT 615.900 491.100 617.100 496.800 ;
        RECT 618.000 497.700 624.300 498.600 ;
        RECT 635.700 498.600 636.900 500.400 ;
        RECT 642.900 498.900 644.100 500.400 ;
        RECT 647.100 499.500 651.900 500.400 ;
        RECT 635.700 497.700 642.000 498.600 ;
        RECT 618.000 495.600 620.100 497.700 ;
        RECT 639.900 495.600 642.000 497.700 ;
        RECT 618.000 493.800 619.800 495.600 ;
        RECT 622.800 493.050 624.600 494.850 ;
        RECT 635.400 493.050 637.200 494.850 ;
        RECT 640.200 493.800 642.000 495.600 ;
        RECT 642.900 496.800 645.900 498.900 ;
        RECT 647.100 498.300 649.200 499.500 ;
        RECT 622.800 492.300 624.900 493.050 ;
        RECT 608.400 489.150 610.200 490.950 ;
        RECT 614.700 490.200 617.100 491.100 ;
        RECT 618.000 490.950 624.900 492.300 ;
        RECT 635.100 492.300 637.200 493.050 ;
        RECT 635.100 490.950 642.000 492.300 ;
        RECT 618.000 490.500 619.800 490.950 ;
        RECT 640.200 490.500 642.000 490.950 ;
        RECT 642.900 491.100 644.100 496.800 ;
        RECT 645.000 493.800 647.100 495.900 ;
        RECT 645.300 492.000 647.100 493.800 ;
        RECT 662.100 493.050 663.900 494.850 ;
        RECT 668.250 493.050 670.050 494.850 ;
        RECT 671.700 493.050 672.600 500.400 ;
        RECT 683.700 493.050 684.900 503.400 ;
        RECT 698.700 493.050 699.900 503.400 ;
        RECT 714.000 500.400 715.800 507.000 ;
        RECT 718.500 501.600 720.300 506.400 ;
        RECT 721.500 503.400 723.300 507.000 ;
        RECT 718.500 500.400 723.600 501.600 ;
        RECT 715.950 498.450 718.050 499.050 ;
        RECT 710.550 497.550 718.050 498.450 ;
        RECT 710.550 495.450 711.450 497.550 ;
        RECT 715.950 496.950 718.050 497.550 ;
        RECT 707.550 494.550 711.450 495.450 ;
        RECT 642.900 490.200 645.300 491.100 ;
        RECT 614.700 490.050 616.200 490.200 ;
        RECT 614.100 487.950 616.200 490.050 ;
        RECT 643.800 490.050 645.300 490.200 ;
        RECT 649.800 490.950 651.900 493.050 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 585.750 485.100 597.450 485.700 ;
        RECT 560.100 471.000 561.900 483.600 ;
        RECT 563.550 471.600 565.350 483.600 ;
        RECT 566.550 471.000 568.350 483.600 ;
        RECT 572.250 483.300 577.050 484.200 ;
        RECT 579.150 484.500 597.450 485.100 ;
        RECT 615.300 486.000 616.200 487.950 ;
        RECT 617.100 487.500 621.000 489.300 ;
        RECT 639.000 487.500 642.900 489.300 ;
        RECT 617.100 487.200 619.200 487.500 ;
        RECT 640.800 487.200 642.900 487.500 ;
        RECT 643.800 487.950 645.900 490.050 ;
        RECT 649.800 489.150 651.600 490.950 ;
        RECT 665.250 489.150 667.050 490.950 ;
        RECT 643.800 486.000 644.700 487.950 ;
        RECT 615.300 484.950 616.800 486.000 ;
        RECT 579.150 484.200 587.550 484.500 ;
        RECT 572.250 482.400 573.450 483.300 ;
        RECT 570.450 480.600 573.450 482.400 ;
        RECT 574.350 482.100 576.150 482.400 ;
        RECT 579.150 482.100 580.050 484.200 ;
        RECT 596.550 483.600 597.450 484.500 ;
        RECT 610.800 483.600 612.900 484.500 ;
        RECT 574.350 481.200 580.050 482.100 ;
        RECT 580.950 482.700 582.750 483.300 ;
        RECT 580.950 481.500 588.750 482.700 ;
        RECT 574.350 480.600 576.150 481.200 ;
        RECT 586.650 480.600 588.750 481.500 ;
        RECT 571.350 477.600 573.450 479.700 ;
        RECT 577.950 479.550 579.750 480.300 ;
        RECT 582.750 479.550 584.550 480.300 ;
        RECT 577.950 478.500 584.550 479.550 ;
        RECT 571.350 471.600 573.150 477.600 ;
        RECT 575.850 471.000 577.650 477.600 ;
        RECT 578.850 471.600 580.650 478.500 ;
        RECT 581.850 471.000 583.650 477.600 ;
        RECT 586.650 471.600 588.450 480.600 ;
        RECT 592.050 471.000 593.850 483.600 ;
        RECT 595.050 481.800 597.450 483.600 ;
        RECT 608.100 482.400 612.900 483.600 ;
        RECT 615.600 483.600 616.800 484.950 ;
        RECT 620.400 483.600 622.500 485.700 ;
        RECT 637.500 483.600 639.600 485.700 ;
        RECT 643.200 484.950 644.700 486.000 ;
        RECT 643.200 483.600 644.400 484.950 ;
        RECT 595.050 471.600 596.850 481.800 ;
        RECT 608.100 471.600 609.900 482.400 ;
        RECT 611.100 471.000 612.900 481.500 ;
        RECT 615.600 471.600 617.400 483.600 ;
        RECT 620.400 482.700 624.900 483.600 ;
        RECT 620.100 471.000 621.900 481.500 ;
        RECT 623.100 471.600 624.900 482.700 ;
        RECT 635.100 482.700 639.600 483.600 ;
        RECT 635.100 471.600 636.900 482.700 ;
        RECT 638.100 471.000 639.900 481.500 ;
        RECT 642.600 471.600 644.400 483.600 ;
        RECT 647.100 483.600 649.200 484.500 ;
        RECT 671.700 483.600 672.600 490.950 ;
        RECT 647.100 482.400 651.900 483.600 ;
        RECT 647.100 471.000 648.900 481.500 ;
        RECT 650.100 471.600 651.900 482.400 ;
        RECT 662.100 482.700 669.900 483.600 ;
        RECT 662.100 471.600 663.900 482.700 ;
        RECT 665.100 471.000 666.900 481.800 ;
        RECT 668.100 471.600 669.900 482.700 ;
        RECT 671.100 471.600 672.900 483.600 ;
        RECT 683.700 477.600 684.900 490.950 ;
        RECT 686.100 489.150 687.900 490.950 ;
        RECT 698.700 477.600 699.900 490.950 ;
        RECT 701.100 489.150 702.900 490.950 ;
        RECT 707.550 490.050 708.450 494.550 ;
        RECT 713.100 493.050 714.900 494.850 ;
        RECT 719.250 493.050 721.050 494.850 ;
        RECT 722.700 493.050 723.600 500.400 ;
        RECT 734.100 501.300 735.900 506.400 ;
        RECT 737.100 502.200 738.900 507.000 ;
        RECT 740.100 501.300 741.900 506.400 ;
        RECT 734.100 499.950 741.900 501.300 ;
        RECT 743.100 500.400 744.900 506.400 ;
        RECT 743.100 498.300 744.300 500.400 ;
        RECT 740.700 497.400 744.300 498.300 ;
        RECT 755.100 498.600 756.900 506.400 ;
        RECT 759.600 500.400 761.400 507.000 ;
        RECT 762.600 502.200 764.400 506.400 ;
        RECT 762.600 500.400 765.300 502.200 ;
        RECT 776.100 500.400 777.900 506.400 ;
        RECT 761.700 498.600 763.500 499.500 ;
        RECT 755.100 497.700 763.500 498.600 ;
        RECT 729.000 495.450 733.050 496.050 ;
        RECT 728.550 493.950 733.050 495.450 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 715.950 490.950 718.050 493.050 ;
        RECT 718.950 490.950 721.050 493.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 703.950 488.550 708.450 490.050 ;
        RECT 716.250 489.150 718.050 490.950 ;
        RECT 703.950 487.950 708.000 488.550 ;
        RECT 722.700 483.600 723.600 490.950 ;
        RECT 728.550 489.450 729.450 493.950 ;
        RECT 737.100 493.050 738.900 494.850 ;
        RECT 740.700 493.050 741.900 497.400 ;
        RECT 743.100 493.050 744.900 494.850 ;
        RECT 755.250 493.050 757.050 494.850 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 755.100 490.950 757.200 493.050 ;
        RECT 725.550 489.000 729.450 489.450 ;
        RECT 734.100 489.150 735.900 490.950 ;
        RECT 724.950 488.550 729.450 489.000 ;
        RECT 724.950 484.950 727.050 488.550 ;
        RECT 740.700 483.600 741.900 490.950 ;
        RECT 713.100 482.700 720.900 483.600 ;
        RECT 683.100 471.600 684.900 477.600 ;
        RECT 686.100 471.000 687.900 477.600 ;
        RECT 698.100 471.600 699.900 477.600 ;
        RECT 701.100 471.000 702.900 477.600 ;
        RECT 713.100 471.600 714.900 482.700 ;
        RECT 716.100 471.000 717.900 481.800 ;
        RECT 719.100 471.600 720.900 482.700 ;
        RECT 722.100 471.600 723.900 483.600 ;
        RECT 734.400 471.000 736.200 483.600 ;
        RECT 739.500 482.100 741.900 483.600 ;
        RECT 739.500 471.600 741.300 482.100 ;
        RECT 742.200 479.100 744.000 480.900 ;
        RECT 758.100 477.600 759.000 497.700 ;
        RECT 764.400 493.050 765.300 500.400 ;
        RECT 776.700 498.300 777.900 500.400 ;
        RECT 779.100 501.300 780.900 506.400 ;
        RECT 782.100 502.200 783.900 507.000 ;
        RECT 785.100 501.300 786.900 506.400 ;
        RECT 779.100 499.950 786.900 501.300 ;
        RECT 776.700 497.400 780.300 498.300 ;
        RECT 799.500 498.000 801.300 506.400 ;
        RECT 776.100 493.050 777.900 494.850 ;
        RECT 779.100 493.050 780.300 497.400 ;
        RECT 798.000 496.800 801.300 498.000 ;
        RECT 806.100 497.400 807.900 507.000 ;
        RECT 818.700 499.200 820.500 506.400 ;
        RECT 823.800 500.400 825.600 507.000 ;
        RECT 839.100 500.400 840.900 506.400 ;
        RECT 842.100 501.300 843.900 507.000 ;
        RECT 846.600 500.400 848.400 506.400 ;
        RECT 851.100 501.300 852.900 507.000 ;
        RECT 854.100 500.400 855.900 506.400 ;
        RECT 818.700 498.300 822.900 499.200 ;
        RECT 782.100 493.050 783.900 494.850 ;
        RECT 798.000 493.050 798.900 496.800 ;
        RECT 800.100 493.050 801.900 494.850 ;
        RECT 806.100 493.050 807.900 494.850 ;
        RECT 818.100 493.050 819.900 494.850 ;
        RECT 821.700 493.050 822.900 498.300 ;
        RECT 839.700 498.600 840.900 500.400 ;
        RECT 846.900 498.900 848.100 500.400 ;
        RECT 851.100 499.500 855.900 500.400 ;
        RECT 839.700 497.700 846.000 498.600 ;
        RECT 843.900 495.600 846.000 497.700 ;
        RECT 823.950 493.050 825.750 494.850 ;
        RECT 839.400 493.050 841.200 494.850 ;
        RECT 844.200 493.800 846.000 495.600 ;
        RECT 846.900 496.800 849.900 498.900 ;
        RECT 851.100 498.300 853.200 499.500 ;
        RECT 760.500 490.950 762.600 493.050 ;
        RECT 763.800 490.950 765.900 493.050 ;
        RECT 775.950 490.950 778.050 493.050 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 799.950 490.950 802.050 493.050 ;
        RECT 802.950 490.950 805.050 493.050 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 823.950 490.950 826.050 493.050 ;
        RECT 839.100 492.300 841.200 493.050 ;
        RECT 839.100 490.950 846.000 492.300 ;
        RECT 760.200 489.150 762.000 490.950 ;
        RECT 764.400 483.600 765.300 490.950 ;
        RECT 779.100 483.600 780.300 490.950 ;
        RECT 785.100 489.150 786.900 490.950 ;
        RECT 742.500 471.000 744.300 477.600 ;
        RECT 755.100 471.000 756.900 477.600 ;
        RECT 758.100 471.600 759.900 477.600 ;
        RECT 761.100 471.000 762.900 483.000 ;
        RECT 764.100 471.600 765.900 483.600 ;
        RECT 779.100 482.100 781.500 483.600 ;
        RECT 777.000 479.100 778.800 480.900 ;
        RECT 776.700 471.000 778.500 477.600 ;
        RECT 779.700 471.600 781.500 482.100 ;
        RECT 784.800 471.000 786.600 483.600 ;
        RECT 798.000 478.800 798.900 490.950 ;
        RECT 803.100 489.150 804.900 490.950 ;
        RECT 799.950 486.450 802.050 487.050 ;
        RECT 817.950 486.450 820.050 487.050 ;
        RECT 799.950 485.550 820.050 486.450 ;
        RECT 799.950 484.950 802.050 485.550 ;
        RECT 817.950 484.950 820.050 485.550 ;
        RECT 798.000 477.900 804.600 478.800 ;
        RECT 798.000 477.600 798.900 477.900 ;
        RECT 797.100 471.600 798.900 477.600 ;
        RECT 803.100 477.600 804.600 477.900 ;
        RECT 821.700 477.600 822.900 490.950 ;
        RECT 844.200 490.500 846.000 490.950 ;
        RECT 846.900 491.100 848.100 496.800 ;
        RECT 849.000 493.800 851.100 495.900 ;
        RECT 849.300 492.000 851.100 493.800 ;
        RECT 846.900 490.200 849.300 491.100 ;
        RECT 847.800 490.050 849.300 490.200 ;
        RECT 853.800 490.950 855.900 493.050 ;
        RECT 843.000 487.500 846.900 489.300 ;
        RECT 844.800 487.200 846.900 487.500 ;
        RECT 847.800 487.950 849.900 490.050 ;
        RECT 853.800 489.150 855.600 490.950 ;
        RECT 847.800 486.000 848.700 487.950 ;
        RECT 841.500 483.600 843.600 485.700 ;
        RECT 847.200 484.950 848.700 486.000 ;
        RECT 847.200 483.600 848.400 484.950 ;
        RECT 839.100 482.700 843.600 483.600 ;
        RECT 800.100 471.000 801.900 477.000 ;
        RECT 803.100 471.600 804.900 477.600 ;
        RECT 806.100 471.000 807.900 477.600 ;
        RECT 818.100 471.000 819.900 477.600 ;
        RECT 821.100 471.600 822.900 477.600 ;
        RECT 824.100 471.000 825.900 477.600 ;
        RECT 839.100 471.600 840.900 482.700 ;
        RECT 842.100 471.000 843.900 481.500 ;
        RECT 846.600 471.600 848.400 483.600 ;
        RECT 851.100 483.600 853.200 484.500 ;
        RECT 851.100 482.400 855.900 483.600 ;
        RECT 851.100 471.000 852.900 481.500 ;
        RECT 854.100 471.600 855.900 482.400 ;
        RECT 11.100 455.400 12.900 467.400 ;
        RECT 14.100 457.200 15.900 468.000 ;
        RECT 17.100 461.400 18.900 467.400 ;
        RECT 11.100 448.050 12.300 455.400 ;
        RECT 17.700 454.500 18.900 461.400 ;
        RECT 21.150 457.200 22.950 467.400 ;
        RECT 13.200 453.600 18.900 454.500 ;
        RECT 20.550 455.400 22.950 457.200 ;
        RECT 24.150 455.400 25.950 468.000 ;
        RECT 29.550 458.400 31.350 467.400 ;
        RECT 34.350 461.400 36.150 468.000 ;
        RECT 37.350 460.500 39.150 467.400 ;
        RECT 40.350 461.400 42.150 468.000 ;
        RECT 44.850 461.400 46.650 467.400 ;
        RECT 33.450 459.450 40.050 460.500 ;
        RECT 33.450 458.700 35.250 459.450 ;
        RECT 38.250 458.700 40.050 459.450 ;
        RECT 44.550 459.300 46.650 461.400 ;
        RECT 29.250 457.500 31.350 458.400 ;
        RECT 41.850 457.800 43.650 458.400 ;
        RECT 29.250 456.300 37.050 457.500 ;
        RECT 35.250 455.700 37.050 456.300 ;
        RECT 37.950 456.900 43.650 457.800 ;
        RECT 20.550 454.500 21.450 455.400 ;
        RECT 37.950 454.800 38.850 456.900 ;
        RECT 41.850 456.600 43.650 456.900 ;
        RECT 44.550 456.600 47.550 458.400 ;
        RECT 44.550 455.700 45.750 456.600 ;
        RECT 30.450 454.500 38.850 454.800 ;
        RECT 20.550 453.900 38.850 454.500 ;
        RECT 40.950 454.800 45.750 455.700 ;
        RECT 49.650 455.400 51.450 468.000 ;
        RECT 52.650 455.400 54.450 467.400 ;
        RECT 65.100 461.400 66.900 468.000 ;
        RECT 68.100 461.400 69.900 467.400 ;
        RECT 13.200 452.700 15.000 453.600 ;
        RECT 11.100 445.950 13.200 448.050 ;
        RECT 11.100 438.600 12.300 445.950 ;
        RECT 14.100 441.300 15.000 452.700 ;
        RECT 20.550 453.300 32.250 453.900 ;
        RECT 16.800 448.050 18.600 449.850 ;
        RECT 16.500 445.950 18.600 448.050 ;
        RECT 13.200 440.400 15.000 441.300 ;
        RECT 13.200 439.500 18.900 440.400 ;
        RECT 11.100 432.600 12.900 438.600 ;
        RECT 14.100 432.000 15.900 438.600 ;
        RECT 17.700 435.600 18.900 439.500 ;
        RECT 20.550 438.600 21.450 453.300 ;
        RECT 30.450 453.000 32.250 453.300 ;
        RECT 22.950 445.950 25.050 448.050 ;
        RECT 32.100 446.400 34.200 448.050 ;
        RECT 22.950 443.400 24.750 445.950 ;
        RECT 26.100 445.200 34.200 446.400 ;
        RECT 26.100 444.600 27.900 445.200 ;
        RECT 29.100 443.400 30.900 444.000 ;
        RECT 22.950 442.200 30.900 443.400 ;
        RECT 40.950 442.200 41.850 454.800 ;
        RECT 44.550 452.100 46.650 452.700 ;
        RECT 50.550 452.100 52.350 452.550 ;
        RECT 44.550 450.900 52.350 452.100 ;
        RECT 44.550 450.600 46.650 450.900 ;
        RECT 50.550 450.750 52.350 450.900 ;
        RECT 53.250 448.050 54.450 455.400 ;
        RECT 65.100 448.050 66.900 449.850 ;
        RECT 68.100 448.050 69.300 461.400 ;
        RECT 84.000 456.600 85.800 467.400 ;
        RECT 84.000 455.400 87.600 456.600 ;
        RECT 89.100 455.400 90.900 468.000 ;
        RECT 101.400 455.400 103.200 468.000 ;
        RECT 106.500 456.900 108.300 467.400 ;
        RECT 109.500 461.400 111.300 468.000 ;
        RECT 122.100 461.400 123.900 467.400 ;
        RECT 109.200 458.100 111.000 459.900 ;
        RECT 106.500 455.400 108.900 456.900 ;
        RECT 83.100 448.050 84.900 449.850 ;
        RECT 86.700 448.050 87.600 455.400 ;
        RECT 88.950 448.050 90.750 449.850 ;
        RECT 101.100 448.050 102.900 449.850 ;
        RECT 107.700 448.050 108.900 455.400 ;
        RECT 122.100 454.500 123.300 461.400 ;
        RECT 125.100 457.200 126.900 468.000 ;
        RECT 128.100 455.400 129.900 467.400 ;
        RECT 143.100 461.400 144.900 468.000 ;
        RECT 146.100 461.400 147.900 467.400 ;
        RECT 149.100 461.400 150.900 468.000 ;
        RECT 161.100 461.400 162.900 468.000 ;
        RECT 164.100 461.400 165.900 467.400 ;
        RECT 167.100 461.400 168.900 468.000 ;
        RECT 179.700 461.400 181.500 468.000 ;
        RECT 122.100 453.600 127.800 454.500 ;
        RECT 126.000 452.700 127.800 453.600 ;
        RECT 122.400 448.050 124.200 449.850 ;
        RECT 49.950 447.750 54.450 448.050 ;
        RECT 48.150 445.950 54.450 447.750 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 67.950 445.950 70.050 448.050 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 122.400 445.950 124.500 448.050 ;
        RECT 29.850 441.000 41.850 442.200 ;
        RECT 29.850 439.200 30.900 441.000 ;
        RECT 40.050 440.400 41.850 441.000 ;
        RECT 20.550 436.800 22.950 438.600 ;
        RECT 17.100 432.600 18.900 435.600 ;
        RECT 21.150 432.600 22.950 436.800 ;
        RECT 24.150 432.000 25.950 438.600 ;
        RECT 26.850 436.200 28.950 437.700 ;
        RECT 29.850 437.400 31.650 439.200 ;
        RECT 53.250 438.600 54.450 445.950 ;
        RECT 32.850 437.550 34.650 438.300 ;
        RECT 32.850 436.500 37.800 437.550 ;
        RECT 26.850 435.600 30.750 436.200 ;
        RECT 36.750 435.600 37.800 436.500 ;
        RECT 44.250 435.600 46.650 437.700 ;
        RECT 27.150 434.700 30.750 435.600 ;
        RECT 28.950 432.600 30.750 434.700 ;
        RECT 33.450 432.000 35.250 435.600 ;
        RECT 36.750 432.600 38.550 435.600 ;
        RECT 39.750 432.000 41.550 435.600 ;
        RECT 44.250 432.600 46.050 435.600 ;
        RECT 49.350 432.000 51.150 438.600 ;
        RECT 52.650 432.600 54.450 438.600 ;
        RECT 68.100 435.600 69.300 445.950 ;
        RECT 86.700 435.600 87.600 445.950 ;
        RECT 104.100 444.150 105.900 445.950 ;
        RECT 107.700 441.600 108.900 445.950 ;
        RECT 110.100 444.150 111.900 445.950 ;
        RECT 107.700 440.700 111.300 441.600 ;
        RECT 101.100 437.700 108.900 439.050 ;
        RECT 65.100 432.000 66.900 435.600 ;
        RECT 68.100 432.600 69.900 435.600 ;
        RECT 83.100 432.000 84.900 435.600 ;
        RECT 86.100 432.600 87.900 435.600 ;
        RECT 89.100 432.000 90.900 435.600 ;
        RECT 101.100 432.600 102.900 437.700 ;
        RECT 104.100 432.000 105.900 436.800 ;
        RECT 107.100 432.600 108.900 437.700 ;
        RECT 110.100 438.600 111.300 440.700 ;
        RECT 126.000 441.300 126.900 452.700 ;
        RECT 128.700 448.050 129.900 455.400 ;
        RECT 146.700 448.050 147.900 461.400 ;
        RECT 164.100 448.050 165.300 461.400 ;
        RECT 180.000 458.100 181.800 459.900 ;
        RECT 182.700 456.900 184.500 467.400 ;
        RECT 182.100 455.400 184.500 456.900 ;
        RECT 187.800 455.400 189.600 468.000 ;
        RECT 200.100 461.400 201.900 467.400 ;
        RECT 203.100 461.400 204.900 468.000 ;
        RECT 182.100 448.050 183.300 455.400 ;
        RECT 190.950 450.450 195.000 451.050 ;
        RECT 188.100 448.050 189.900 449.850 ;
        RECT 190.950 448.950 195.450 450.450 ;
        RECT 127.800 445.950 129.900 448.050 ;
        RECT 142.950 445.950 145.050 448.050 ;
        RECT 145.950 445.950 148.050 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 166.950 445.950 169.050 448.050 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 187.950 445.950 190.050 448.050 ;
        RECT 126.000 440.400 127.800 441.300 ;
        RECT 122.100 439.500 127.800 440.400 ;
        RECT 110.100 432.600 111.900 438.600 ;
        RECT 122.100 435.600 123.300 439.500 ;
        RECT 128.700 438.600 129.900 445.950 ;
        RECT 143.100 444.150 144.900 445.950 ;
        RECT 146.700 440.700 147.900 445.950 ;
        RECT 148.950 444.150 150.750 445.950 ;
        RECT 161.250 444.150 163.050 445.950 ;
        RECT 122.100 432.600 123.900 435.600 ;
        RECT 125.100 432.000 126.900 438.600 ;
        RECT 128.100 432.600 129.900 438.600 ;
        RECT 143.700 439.800 147.900 440.700 ;
        RECT 164.100 440.700 165.300 445.950 ;
        RECT 167.100 444.150 168.900 445.950 ;
        RECT 179.100 444.150 180.900 445.950 ;
        RECT 182.100 441.600 183.300 445.950 ;
        RECT 185.100 444.150 186.900 445.950 ;
        RECT 194.550 445.050 195.450 448.950 ;
        RECT 200.700 448.050 201.900 461.400 ;
        RECT 206.550 455.400 208.350 467.400 ;
        RECT 209.550 455.400 211.350 468.000 ;
        RECT 214.350 461.400 216.150 467.400 ;
        RECT 218.850 461.400 220.650 468.000 ;
        RECT 214.350 459.300 216.450 461.400 ;
        RECT 221.850 460.500 223.650 467.400 ;
        RECT 224.850 461.400 226.650 468.000 ;
        RECT 220.950 459.450 227.550 460.500 ;
        RECT 220.950 458.700 222.750 459.450 ;
        RECT 225.750 458.700 227.550 459.450 ;
        RECT 229.650 458.400 231.450 467.400 ;
        RECT 213.450 456.600 216.450 458.400 ;
        RECT 217.350 457.800 219.150 458.400 ;
        RECT 217.350 456.900 223.050 457.800 ;
        RECT 229.650 457.500 231.750 458.400 ;
        RECT 217.350 456.600 219.150 456.900 ;
        RECT 215.250 455.700 216.450 456.600 ;
        RECT 203.100 448.050 204.900 449.850 ;
        RECT 206.550 448.050 207.750 455.400 ;
        RECT 215.250 454.800 220.050 455.700 ;
        RECT 208.650 452.100 210.450 452.550 ;
        RECT 214.350 452.100 216.450 452.700 ;
        RECT 208.650 450.900 216.450 452.100 ;
        RECT 208.650 450.750 210.450 450.900 ;
        RECT 214.350 450.600 216.450 450.900 ;
        RECT 199.950 445.950 202.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 206.550 447.750 211.050 448.050 ;
        RECT 206.550 445.950 212.850 447.750 ;
        RECT 190.950 443.550 195.450 445.050 ;
        RECT 190.950 442.950 195.000 443.550 ;
        RECT 179.700 440.700 183.300 441.600 ;
        RECT 164.100 439.800 168.300 440.700 ;
        RECT 143.700 432.600 145.500 439.800 ;
        RECT 148.800 432.000 150.600 438.600 ;
        RECT 161.400 432.000 163.200 438.600 ;
        RECT 166.500 432.600 168.300 439.800 ;
        RECT 179.700 438.600 180.900 440.700 ;
        RECT 179.100 432.600 180.900 438.600 ;
        RECT 182.100 437.700 189.900 439.050 ;
        RECT 182.100 432.600 183.900 437.700 ;
        RECT 185.100 432.000 186.900 436.800 ;
        RECT 188.100 432.600 189.900 437.700 ;
        RECT 200.700 435.600 201.900 445.950 ;
        RECT 206.550 438.600 207.750 445.950 ;
        RECT 219.150 442.200 220.050 454.800 ;
        RECT 222.150 454.800 223.050 456.900 ;
        RECT 223.950 456.300 231.750 457.500 ;
        RECT 223.950 455.700 225.750 456.300 ;
        RECT 235.050 455.400 236.850 468.000 ;
        RECT 238.050 457.200 239.850 467.400 ;
        RECT 238.050 455.400 240.450 457.200 ;
        RECT 251.400 455.400 253.200 468.000 ;
        RECT 256.500 456.900 258.300 467.400 ;
        RECT 259.500 461.400 261.300 468.000 ;
        RECT 272.100 461.400 273.900 468.000 ;
        RECT 275.100 461.400 276.900 467.400 ;
        RECT 278.100 461.400 279.900 468.000 ;
        RECT 290.100 461.400 291.900 468.000 ;
        RECT 293.100 461.400 294.900 467.400 ;
        RECT 259.200 458.100 261.000 459.900 ;
        RECT 256.500 455.400 258.900 456.900 ;
        RECT 222.150 454.500 230.550 454.800 ;
        RECT 239.550 454.500 240.450 455.400 ;
        RECT 222.150 453.900 240.450 454.500 ;
        RECT 228.750 453.300 240.450 453.900 ;
        RECT 228.750 453.000 230.550 453.300 ;
        RECT 226.800 446.400 228.900 448.050 ;
        RECT 226.800 445.200 234.900 446.400 ;
        RECT 235.950 445.950 238.050 448.050 ;
        RECT 233.100 444.600 234.900 445.200 ;
        RECT 230.100 443.400 231.900 444.000 ;
        RECT 236.250 443.400 238.050 445.950 ;
        RECT 230.100 442.200 238.050 443.400 ;
        RECT 219.150 441.000 231.150 442.200 ;
        RECT 219.150 440.400 220.950 441.000 ;
        RECT 230.100 439.200 231.150 441.000 ;
        RECT 200.100 432.600 201.900 435.600 ;
        RECT 203.100 432.000 204.900 435.600 ;
        RECT 206.550 432.600 208.350 438.600 ;
        RECT 209.850 432.000 211.650 438.600 ;
        RECT 214.350 435.600 216.750 437.700 ;
        RECT 226.350 437.550 228.150 438.300 ;
        RECT 223.200 436.500 228.150 437.550 ;
        RECT 229.350 437.400 231.150 439.200 ;
        RECT 239.550 438.600 240.450 453.300 ;
        RECT 251.100 448.050 252.900 449.850 ;
        RECT 257.700 448.050 258.900 455.400 ;
        RECT 275.700 448.050 276.900 461.400 ;
        RECT 290.100 448.050 291.900 449.850 ;
        RECT 293.100 448.050 294.300 461.400 ;
        RECT 305.100 455.400 306.900 467.400 ;
        RECT 308.100 457.200 309.900 468.000 ;
        RECT 311.100 461.400 312.900 467.400 ;
        RECT 323.100 461.400 324.900 468.000 ;
        RECT 326.100 461.400 327.900 467.400 ;
        RECT 329.100 461.400 330.900 468.000 ;
        RECT 341.100 461.400 342.900 468.000 ;
        RECT 344.100 461.400 345.900 467.400 ;
        RECT 347.100 461.400 348.900 468.000 ;
        RECT 305.100 448.050 306.300 455.400 ;
        RECT 311.700 454.500 312.900 461.400 ;
        RECT 307.200 453.600 312.900 454.500 ;
        RECT 307.200 452.700 309.000 453.600 ;
        RECT 250.950 445.950 253.050 448.050 ;
        RECT 253.950 445.950 256.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 277.950 445.950 280.050 448.050 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 292.950 445.950 295.050 448.050 ;
        RECT 305.100 445.950 307.200 448.050 ;
        RECT 254.100 444.150 255.900 445.950 ;
        RECT 257.700 441.600 258.900 445.950 ;
        RECT 260.100 444.150 261.900 445.950 ;
        RECT 272.100 444.150 273.900 445.950 ;
        RECT 257.700 440.700 261.300 441.600 ;
        RECT 275.700 440.700 276.900 445.950 ;
        RECT 277.950 444.150 279.750 445.950 ;
        RECT 223.200 435.600 224.250 436.500 ;
        RECT 232.050 436.200 234.150 437.700 ;
        RECT 230.250 435.600 234.150 436.200 ;
        RECT 214.950 432.600 216.750 435.600 ;
        RECT 219.450 432.000 221.250 435.600 ;
        RECT 222.450 432.600 224.250 435.600 ;
        RECT 225.750 432.000 227.550 435.600 ;
        RECT 230.250 434.700 233.850 435.600 ;
        RECT 230.250 432.600 232.050 434.700 ;
        RECT 235.050 432.000 236.850 438.600 ;
        RECT 238.050 436.800 240.450 438.600 ;
        RECT 251.100 437.700 258.900 439.050 ;
        RECT 238.050 432.600 239.850 436.800 ;
        RECT 251.100 432.600 252.900 437.700 ;
        RECT 254.100 432.000 255.900 436.800 ;
        RECT 257.100 432.600 258.900 437.700 ;
        RECT 260.100 438.600 261.300 440.700 ;
        RECT 272.700 439.800 276.900 440.700 ;
        RECT 260.100 432.600 261.900 438.600 ;
        RECT 272.700 432.600 274.500 439.800 ;
        RECT 277.800 432.000 279.600 438.600 ;
        RECT 293.100 435.600 294.300 445.950 ;
        RECT 305.100 438.600 306.300 445.950 ;
        RECT 308.100 441.300 309.000 452.700 ;
        RECT 310.800 448.050 312.600 449.850 ;
        RECT 326.100 448.050 327.300 461.400 ;
        RECT 344.100 448.050 345.300 461.400 ;
        RECT 350.550 455.400 352.350 467.400 ;
        RECT 353.550 455.400 355.350 468.000 ;
        RECT 358.350 461.400 360.150 467.400 ;
        RECT 362.850 461.400 364.650 468.000 ;
        RECT 358.350 459.300 360.450 461.400 ;
        RECT 365.850 460.500 367.650 467.400 ;
        RECT 368.850 461.400 370.650 468.000 ;
        RECT 364.950 459.450 371.550 460.500 ;
        RECT 364.950 458.700 366.750 459.450 ;
        RECT 369.750 458.700 371.550 459.450 ;
        RECT 373.650 458.400 375.450 467.400 ;
        RECT 357.450 456.600 360.450 458.400 ;
        RECT 361.350 457.800 363.150 458.400 ;
        RECT 361.350 456.900 367.050 457.800 ;
        RECT 373.650 457.500 375.750 458.400 ;
        RECT 361.350 456.600 363.150 456.900 ;
        RECT 359.250 455.700 360.450 456.600 ;
        RECT 350.550 448.050 351.750 455.400 ;
        RECT 359.250 454.800 364.050 455.700 ;
        RECT 352.650 452.100 354.450 452.550 ;
        RECT 358.350 452.100 360.450 452.700 ;
        RECT 352.650 450.900 360.450 452.100 ;
        RECT 352.650 450.750 354.450 450.900 ;
        RECT 358.350 450.600 360.450 450.900 ;
        RECT 310.500 445.950 312.600 448.050 ;
        RECT 322.950 445.950 325.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 350.550 447.750 355.050 448.050 ;
        RECT 350.550 445.950 356.850 447.750 ;
        RECT 323.250 444.150 325.050 445.950 ;
        RECT 307.200 440.400 309.000 441.300 ;
        RECT 326.100 440.700 327.300 445.950 ;
        RECT 329.100 444.150 330.900 445.950 ;
        RECT 341.250 444.150 343.050 445.950 ;
        RECT 344.100 440.700 345.300 445.950 ;
        RECT 347.100 444.150 348.900 445.950 ;
        RECT 307.200 439.500 312.900 440.400 ;
        RECT 326.100 439.800 330.300 440.700 ;
        RECT 344.100 439.800 348.300 440.700 ;
        RECT 290.100 432.000 291.900 435.600 ;
        RECT 293.100 432.600 294.900 435.600 ;
        RECT 305.100 432.600 306.900 438.600 ;
        RECT 308.100 432.000 309.900 438.600 ;
        RECT 311.700 435.600 312.900 439.500 ;
        RECT 311.100 432.600 312.900 435.600 ;
        RECT 323.400 432.000 325.200 438.600 ;
        RECT 328.500 432.600 330.300 439.800 ;
        RECT 341.400 432.000 343.200 438.600 ;
        RECT 346.500 432.600 348.300 439.800 ;
        RECT 350.550 438.600 351.750 445.950 ;
        RECT 363.150 442.200 364.050 454.800 ;
        RECT 366.150 454.800 367.050 456.900 ;
        RECT 367.950 456.300 375.750 457.500 ;
        RECT 367.950 455.700 369.750 456.300 ;
        RECT 379.050 455.400 380.850 468.000 ;
        RECT 382.050 457.200 383.850 467.400 ;
        RECT 395.700 461.400 397.500 468.000 ;
        RECT 396.000 458.100 397.800 459.900 ;
        RECT 382.050 455.400 384.450 457.200 ;
        RECT 398.700 456.900 400.500 467.400 ;
        RECT 366.150 454.500 374.550 454.800 ;
        RECT 383.550 454.500 384.450 455.400 ;
        RECT 366.150 453.900 384.450 454.500 ;
        RECT 372.750 453.300 384.450 453.900 ;
        RECT 372.750 453.000 374.550 453.300 ;
        RECT 370.800 446.400 372.900 448.050 ;
        RECT 370.800 445.200 378.900 446.400 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 377.100 444.600 378.900 445.200 ;
        RECT 374.100 443.400 375.900 444.000 ;
        RECT 380.250 443.400 382.050 445.950 ;
        RECT 374.100 442.200 382.050 443.400 ;
        RECT 363.150 441.000 375.150 442.200 ;
        RECT 363.150 440.400 364.950 441.000 ;
        RECT 374.100 439.200 375.150 441.000 ;
        RECT 350.550 432.600 352.350 438.600 ;
        RECT 353.850 432.000 355.650 438.600 ;
        RECT 358.350 435.600 360.750 437.700 ;
        RECT 370.350 437.550 372.150 438.300 ;
        RECT 367.200 436.500 372.150 437.550 ;
        RECT 373.350 437.400 375.150 439.200 ;
        RECT 383.550 438.600 384.450 453.300 ;
        RECT 398.100 455.400 400.500 456.900 ;
        RECT 403.800 455.400 405.600 468.000 ;
        RECT 416.700 461.400 418.500 468.000 ;
        RECT 417.000 458.100 418.800 459.900 ;
        RECT 419.700 456.900 421.500 467.400 ;
        RECT 419.100 455.400 421.500 456.900 ;
        RECT 424.800 455.400 426.600 468.000 ;
        RECT 440.100 461.400 441.900 467.400 ;
        RECT 443.100 461.400 444.900 468.000 ;
        RECT 455.700 461.400 457.500 468.000 ;
        RECT 398.100 448.050 399.300 455.400 ;
        RECT 404.100 448.050 405.900 449.850 ;
        RECT 419.100 448.050 420.300 455.400 ;
        RECT 425.100 448.050 426.900 449.850 ;
        RECT 440.700 448.050 441.900 461.400 ;
        RECT 456.000 458.100 457.800 459.900 ;
        RECT 458.700 456.900 460.500 467.400 ;
        RECT 458.100 455.400 460.500 456.900 ;
        RECT 463.800 455.400 465.600 468.000 ;
        RECT 479.700 461.400 481.500 468.000 ;
        RECT 480.000 458.100 481.800 459.900 ;
        RECT 482.700 456.900 484.500 467.400 ;
        RECT 482.100 455.400 484.500 456.900 ;
        RECT 487.800 455.400 489.600 468.000 ;
        RECT 504.000 456.600 505.800 467.400 ;
        RECT 504.000 455.400 507.600 456.600 ;
        RECT 509.100 455.400 510.900 468.000 ;
        RECT 521.100 456.300 522.900 467.400 ;
        RECT 524.100 457.200 525.900 468.000 ;
        RECT 527.100 456.300 528.900 467.400 ;
        RECT 521.100 455.400 528.900 456.300 ;
        RECT 530.100 455.400 531.900 467.400 ;
        RECT 545.100 455.400 546.900 467.400 ;
        RECT 548.100 457.200 549.900 468.000 ;
        RECT 551.100 461.400 552.900 467.400 ;
        RECT 443.100 448.050 444.900 449.850 ;
        RECT 458.100 448.050 459.300 455.400 ;
        RECT 464.100 448.050 465.900 449.850 ;
        RECT 482.100 448.050 483.300 455.400 ;
        RECT 488.100 448.050 489.900 449.850 ;
        RECT 503.100 448.050 504.900 449.850 ;
        RECT 506.700 448.050 507.600 455.400 ;
        RECT 508.950 453.450 511.050 453.900 ;
        RECT 526.950 453.450 529.050 454.050 ;
        RECT 508.950 452.550 529.050 453.450 ;
        RECT 508.950 451.800 511.050 452.550 ;
        RECT 526.950 451.950 529.050 452.550 ;
        RECT 508.950 448.050 510.750 449.850 ;
        RECT 524.250 448.050 526.050 449.850 ;
        RECT 530.700 448.050 531.600 455.400 ;
        RECT 545.100 448.050 546.300 455.400 ;
        RECT 551.700 454.500 552.900 461.400 ;
        RECT 566.100 456.300 567.900 467.400 ;
        RECT 569.100 457.200 570.900 468.000 ;
        RECT 572.100 456.300 573.900 467.400 ;
        RECT 566.100 455.400 573.900 456.300 ;
        RECT 575.100 455.400 576.900 467.400 ;
        RECT 587.100 461.400 588.900 467.400 ;
        RECT 590.100 462.000 591.900 468.000 ;
        RECT 588.000 461.100 588.900 461.400 ;
        RECT 593.100 461.400 594.900 467.400 ;
        RECT 596.100 461.400 597.900 468.000 ;
        RECT 608.100 461.400 609.900 468.000 ;
        RECT 611.100 461.400 612.900 467.400 ;
        RECT 593.100 461.100 594.600 461.400 ;
        RECT 588.000 460.200 594.600 461.100 ;
        RECT 547.200 453.600 552.900 454.500 ;
        RECT 547.200 452.700 549.000 453.600 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 400.950 445.950 403.050 448.050 ;
        RECT 403.950 445.950 406.050 448.050 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 424.950 445.950 427.050 448.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 463.950 445.950 466.050 448.050 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 520.950 445.950 523.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 445.950 532.050 448.050 ;
        RECT 545.100 445.950 547.200 448.050 ;
        RECT 395.100 444.150 396.900 445.950 ;
        RECT 398.100 441.600 399.300 445.950 ;
        RECT 401.100 444.150 402.900 445.950 ;
        RECT 416.100 444.150 417.900 445.950 ;
        RECT 419.100 441.600 420.300 445.950 ;
        RECT 422.100 444.150 423.900 445.950 ;
        RECT 395.700 440.700 399.300 441.600 ;
        RECT 416.700 440.700 420.300 441.600 ;
        RECT 395.700 438.600 396.900 440.700 ;
        RECT 367.200 435.600 368.250 436.500 ;
        RECT 376.050 436.200 378.150 437.700 ;
        RECT 374.250 435.600 378.150 436.200 ;
        RECT 358.950 432.600 360.750 435.600 ;
        RECT 363.450 432.000 365.250 435.600 ;
        RECT 366.450 432.600 368.250 435.600 ;
        RECT 369.750 432.000 371.550 435.600 ;
        RECT 374.250 434.700 377.850 435.600 ;
        RECT 374.250 432.600 376.050 434.700 ;
        RECT 379.050 432.000 380.850 438.600 ;
        RECT 382.050 436.800 384.450 438.600 ;
        RECT 382.050 432.600 383.850 436.800 ;
        RECT 395.100 432.600 396.900 438.600 ;
        RECT 398.100 437.700 405.900 439.050 ;
        RECT 416.700 438.600 417.900 440.700 ;
        RECT 398.100 432.600 399.900 437.700 ;
        RECT 401.100 432.000 402.900 436.800 ;
        RECT 404.100 432.600 405.900 437.700 ;
        RECT 416.100 432.600 417.900 438.600 ;
        RECT 419.100 437.700 426.900 439.050 ;
        RECT 419.100 432.600 420.900 437.700 ;
        RECT 422.100 432.000 423.900 436.800 ;
        RECT 425.100 432.600 426.900 437.700 ;
        RECT 440.700 435.600 441.900 445.950 ;
        RECT 455.100 444.150 456.900 445.950 ;
        RECT 458.100 441.600 459.300 445.950 ;
        RECT 461.100 444.150 462.900 445.950 ;
        RECT 479.100 444.150 480.900 445.950 ;
        RECT 482.100 441.600 483.300 445.950 ;
        RECT 485.100 444.150 486.900 445.950 ;
        RECT 455.700 440.700 459.300 441.600 ;
        RECT 479.700 440.700 483.300 441.600 ;
        RECT 455.700 438.600 456.900 440.700 ;
        RECT 440.100 432.600 441.900 435.600 ;
        RECT 443.100 432.000 444.900 435.600 ;
        RECT 455.100 432.600 456.900 438.600 ;
        RECT 458.100 437.700 465.900 439.050 ;
        RECT 479.700 438.600 480.900 440.700 ;
        RECT 458.100 432.600 459.900 437.700 ;
        RECT 461.100 432.000 462.900 436.800 ;
        RECT 464.100 432.600 465.900 437.700 ;
        RECT 479.100 432.600 480.900 438.600 ;
        RECT 482.100 437.700 489.900 439.050 ;
        RECT 482.100 432.600 483.900 437.700 ;
        RECT 485.100 432.000 486.900 436.800 ;
        RECT 488.100 432.600 489.900 437.700 ;
        RECT 506.700 435.600 507.600 445.950 ;
        RECT 521.100 444.150 522.900 445.950 ;
        RECT 527.250 444.150 529.050 445.950 ;
        RECT 530.700 438.600 531.600 445.950 ;
        RECT 503.100 432.000 504.900 435.600 ;
        RECT 506.100 432.600 507.900 435.600 ;
        RECT 509.100 432.000 510.900 435.600 ;
        RECT 522.000 432.000 523.800 438.600 ;
        RECT 526.500 437.400 531.600 438.600 ;
        RECT 545.100 438.600 546.300 445.950 ;
        RECT 548.100 441.300 549.000 452.700 ;
        RECT 550.800 448.050 552.600 449.850 ;
        RECT 569.250 448.050 571.050 449.850 ;
        RECT 575.700 448.050 576.600 455.400 ;
        RECT 588.000 448.050 588.900 460.200 ;
        RECT 593.100 448.050 594.900 449.850 ;
        RECT 608.100 448.050 609.900 449.850 ;
        RECT 611.100 448.050 612.300 461.400 ;
        RECT 623.100 455.400 624.900 467.400 ;
        RECT 626.100 456.300 627.900 467.400 ;
        RECT 629.100 457.200 630.900 468.000 ;
        RECT 632.100 456.300 633.900 467.400 ;
        RECT 644.100 461.400 645.900 468.000 ;
        RECT 647.100 461.400 648.900 467.400 ;
        RECT 650.100 461.400 651.900 468.000 ;
        RECT 626.100 455.400 633.900 456.300 ;
        RECT 623.400 448.050 624.300 455.400 ;
        RECT 628.950 448.050 630.750 449.850 ;
        RECT 647.700 448.050 648.900 461.400 ;
        RECT 663.000 456.600 664.800 467.400 ;
        RECT 663.000 455.400 666.600 456.600 ;
        RECT 668.100 455.400 669.900 468.000 ;
        RECT 680.100 455.400 681.900 467.400 ;
        RECT 683.100 456.000 684.900 468.000 ;
        RECT 686.100 461.400 687.900 467.400 ;
        RECT 689.100 461.400 690.900 468.000 ;
        RECT 701.100 461.400 702.900 468.000 ;
        RECT 704.100 461.400 705.900 467.400 ;
        RECT 707.100 461.400 708.900 468.000 ;
        RECT 719.100 461.400 720.900 468.000 ;
        RECT 722.100 461.400 723.900 467.400 ;
        RECT 725.100 461.400 726.900 468.000 ;
        RECT 737.100 461.400 738.900 468.000 ;
        RECT 740.100 461.400 741.900 467.400 ;
        RECT 743.100 461.400 744.900 468.000 ;
        RECT 755.700 461.400 757.500 468.000 ;
        RECT 662.100 448.050 663.900 449.850 ;
        RECT 665.700 448.050 666.600 455.400 ;
        RECT 667.950 448.050 669.750 449.850 ;
        RECT 680.700 448.050 681.600 455.400 ;
        RECT 684.000 448.050 685.800 449.850 ;
        RECT 550.500 445.950 552.600 448.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 622.950 445.950 625.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 628.950 445.950 631.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 680.100 445.950 682.200 448.050 ;
        RECT 683.400 445.950 685.500 448.050 ;
        RECT 566.100 444.150 567.900 445.950 ;
        RECT 572.250 444.150 574.050 445.950 ;
        RECT 547.200 440.400 549.000 441.300 ;
        RECT 547.200 439.500 552.900 440.400 ;
        RECT 526.500 432.600 528.300 437.400 ;
        RECT 529.500 432.000 531.300 435.600 ;
        RECT 545.100 432.600 546.900 438.600 ;
        RECT 548.100 432.000 549.900 438.600 ;
        RECT 551.700 435.600 552.900 439.500 ;
        RECT 575.700 438.600 576.600 445.950 ;
        RECT 588.000 442.200 588.900 445.950 ;
        RECT 590.100 444.150 591.900 445.950 ;
        RECT 596.100 444.150 597.900 445.950 ;
        RECT 588.000 441.000 591.300 442.200 ;
        RECT 551.100 432.600 552.900 435.600 ;
        RECT 567.000 432.000 568.800 438.600 ;
        RECT 571.500 437.400 576.600 438.600 ;
        RECT 571.500 432.600 573.300 437.400 ;
        RECT 574.500 432.000 576.300 435.600 ;
        RECT 589.500 432.600 591.300 441.000 ;
        RECT 596.100 432.000 597.900 441.600 ;
        RECT 611.100 435.600 612.300 445.950 ;
        RECT 623.400 438.600 624.300 445.950 ;
        RECT 625.950 444.150 627.750 445.950 ;
        RECT 632.100 444.150 633.900 445.950 ;
        RECT 644.100 444.150 645.900 445.950 ;
        RECT 647.700 440.700 648.900 445.950 ;
        RECT 649.950 444.150 651.750 445.950 ;
        RECT 644.700 439.800 648.900 440.700 ;
        RECT 623.400 437.400 628.500 438.600 ;
        RECT 608.100 432.000 609.900 435.600 ;
        RECT 611.100 432.600 612.900 435.600 ;
        RECT 623.700 432.000 625.500 435.600 ;
        RECT 626.700 432.600 628.500 437.400 ;
        RECT 631.200 432.000 633.000 438.600 ;
        RECT 644.700 432.600 646.500 439.800 ;
        RECT 649.800 432.000 651.600 438.600 ;
        RECT 665.700 435.600 666.600 445.950 ;
        RECT 680.700 438.600 681.600 445.950 ;
        RECT 687.000 441.300 687.900 461.400 ;
        RECT 704.100 448.050 705.300 461.400 ;
        RECT 722.100 448.050 723.300 461.400 ;
        RECT 740.700 448.050 741.900 461.400 ;
        RECT 756.000 458.100 757.800 459.900 ;
        RECT 758.700 456.900 760.500 467.400 ;
        RECT 758.100 455.400 760.500 456.900 ;
        RECT 763.800 455.400 765.600 468.000 ;
        RECT 779.100 461.400 780.900 468.000 ;
        RECT 782.100 461.400 783.900 467.400 ;
        RECT 758.100 448.050 759.300 455.400 ;
        RECT 764.100 448.050 765.900 449.850 ;
        RECT 779.100 448.050 780.900 449.850 ;
        RECT 782.100 448.050 783.300 461.400 ;
        RECT 794.100 455.400 795.900 467.400 ;
        RECT 797.100 456.300 798.900 467.400 ;
        RECT 800.100 457.200 801.900 468.000 ;
        RECT 803.100 456.300 804.900 467.400 ;
        RECT 797.100 455.400 804.900 456.300 ;
        RECT 819.000 456.600 820.800 467.400 ;
        RECT 819.000 455.400 822.600 456.600 ;
        RECT 824.100 455.400 825.900 468.000 ;
        RECT 837.600 456.900 839.400 467.400 ;
        RECT 837.000 455.400 839.400 456.900 ;
        RECT 840.600 455.400 842.400 468.000 ;
        RECT 845.100 455.400 846.900 467.400 ;
        RECT 860.100 461.400 861.900 468.000 ;
        RECT 863.100 461.400 864.900 467.400 ;
        RECT 866.100 461.400 867.900 468.000 ;
        RECT 794.400 448.050 795.300 455.400 ;
        RECT 799.950 448.050 801.750 449.850 ;
        RECT 818.100 448.050 819.900 449.850 ;
        RECT 821.700 448.050 822.600 455.400 ;
        RECT 823.950 448.050 825.750 449.850 ;
        RECT 837.000 448.050 838.200 455.400 ;
        RECT 845.700 453.900 846.900 455.400 ;
        RECT 839.100 452.700 846.900 453.900 ;
        RECT 839.100 452.100 840.900 452.700 ;
        RECT 688.800 445.950 690.900 448.050 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 736.950 445.950 739.050 448.050 ;
        RECT 739.950 445.950 742.050 448.050 ;
        RECT 742.950 445.950 745.050 448.050 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 757.950 445.950 760.050 448.050 ;
        RECT 760.950 445.950 763.050 448.050 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 793.950 445.950 796.050 448.050 ;
        RECT 796.950 445.950 799.050 448.050 ;
        RECT 799.950 445.950 802.050 448.050 ;
        RECT 802.950 445.950 805.050 448.050 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 823.950 445.950 826.050 448.050 ;
        RECT 836.100 445.950 838.200 448.050 ;
        RECT 688.950 444.150 690.750 445.950 ;
        RECT 701.250 444.150 703.050 445.950 ;
        RECT 682.500 440.400 690.900 441.300 ;
        RECT 682.500 439.500 684.300 440.400 ;
        RECT 680.700 436.800 683.400 438.600 ;
        RECT 662.100 432.000 663.900 435.600 ;
        RECT 665.100 432.600 666.900 435.600 ;
        RECT 668.100 432.000 669.900 435.600 ;
        RECT 681.600 432.600 683.400 436.800 ;
        RECT 684.600 432.000 686.400 438.600 ;
        RECT 689.100 432.600 690.900 440.400 ;
        RECT 704.100 440.700 705.300 445.950 ;
        RECT 707.100 444.150 708.900 445.950 ;
        RECT 719.250 444.150 721.050 445.950 ;
        RECT 722.100 440.700 723.300 445.950 ;
        RECT 725.100 444.150 726.900 445.950 ;
        RECT 737.100 444.150 738.900 445.950 ;
        RECT 740.700 440.700 741.900 445.950 ;
        RECT 742.950 444.150 744.750 445.950 ;
        RECT 755.100 444.150 756.900 445.950 ;
        RECT 758.100 441.600 759.300 445.950 ;
        RECT 761.100 444.150 762.900 445.950 ;
        RECT 704.100 439.800 708.300 440.700 ;
        RECT 722.100 439.800 726.300 440.700 ;
        RECT 701.400 432.000 703.200 438.600 ;
        RECT 706.500 432.600 708.300 439.800 ;
        RECT 719.400 432.000 721.200 438.600 ;
        RECT 724.500 432.600 726.300 439.800 ;
        RECT 737.700 439.800 741.900 440.700 ;
        RECT 755.700 440.700 759.300 441.600 ;
        RECT 737.700 432.600 739.500 439.800 ;
        RECT 755.700 438.600 756.900 440.700 ;
        RECT 742.800 432.000 744.600 438.600 ;
        RECT 755.100 432.600 756.900 438.600 ;
        RECT 758.100 437.700 765.900 439.050 ;
        RECT 758.100 432.600 759.900 437.700 ;
        RECT 761.100 432.000 762.900 436.800 ;
        RECT 764.100 432.600 765.900 437.700 ;
        RECT 782.100 435.600 783.300 445.950 ;
        RECT 794.400 438.600 795.300 445.950 ;
        RECT 796.950 444.150 798.750 445.950 ;
        RECT 803.100 444.150 804.900 445.950 ;
        RECT 799.950 441.450 802.050 442.050 ;
        RECT 808.950 441.450 811.050 442.050 ;
        RECT 817.950 441.450 820.050 442.050 ;
        RECT 799.950 440.550 820.050 441.450 ;
        RECT 799.950 439.950 802.050 440.550 ;
        RECT 808.950 439.950 811.050 440.550 ;
        RECT 817.950 439.950 820.050 440.550 ;
        RECT 794.400 437.400 799.500 438.600 ;
        RECT 779.100 432.000 780.900 435.600 ;
        RECT 782.100 432.600 783.900 435.600 ;
        RECT 794.700 432.000 796.500 435.600 ;
        RECT 797.700 432.600 799.500 437.400 ;
        RECT 802.200 432.000 804.000 438.600 ;
        RECT 821.700 435.600 822.600 445.950 ;
        RECT 836.100 438.600 837.000 445.950 ;
        RECT 839.400 441.600 840.300 452.100 ;
        RECT 841.200 448.050 843.000 449.850 ;
        RECT 863.100 448.050 864.300 461.400 ;
        RECT 841.500 445.950 843.600 448.050 ;
        RECT 844.800 445.950 846.900 448.050 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 865.950 445.950 868.050 448.050 ;
        RECT 844.800 444.150 846.600 445.950 ;
        RECT 860.250 444.150 862.050 445.950 ;
        RECT 838.200 440.700 840.300 441.600 ;
        RECT 863.100 440.700 864.300 445.950 ;
        RECT 866.100 444.150 867.900 445.950 ;
        RECT 838.200 439.800 843.600 440.700 ;
        RECT 863.100 439.800 867.300 440.700 ;
        RECT 818.100 432.000 819.900 435.600 ;
        RECT 821.100 432.600 822.900 435.600 ;
        RECT 824.100 432.000 825.900 435.600 ;
        RECT 836.100 432.600 837.900 438.600 ;
        RECT 839.100 432.000 840.900 438.000 ;
        RECT 842.700 435.600 843.600 439.800 ;
        RECT 842.100 432.600 843.900 435.600 ;
        RECT 845.100 432.600 846.900 435.600 ;
        RECT 845.700 432.000 846.900 432.600 ;
        RECT 860.400 432.000 862.200 438.600 ;
        RECT 865.500 432.600 867.300 439.800 ;
        RECT 3.150 424.200 4.950 428.400 ;
        RECT 2.550 422.400 4.950 424.200 ;
        RECT 6.150 422.400 7.950 429.000 ;
        RECT 10.950 426.300 12.750 428.400 ;
        RECT 9.150 425.400 12.750 426.300 ;
        RECT 15.450 425.400 17.250 429.000 ;
        RECT 18.750 425.400 20.550 428.400 ;
        RECT 21.750 425.400 23.550 429.000 ;
        RECT 26.250 425.400 28.050 428.400 ;
        RECT 8.850 424.800 12.750 425.400 ;
        RECT 8.850 423.300 10.950 424.800 ;
        RECT 18.750 424.500 19.800 425.400 ;
        RECT 2.550 407.700 3.450 422.400 ;
        RECT 11.850 421.800 13.650 423.600 ;
        RECT 14.850 423.450 19.800 424.500 ;
        RECT 14.850 422.700 16.650 423.450 ;
        RECT 26.250 423.300 28.650 425.400 ;
        RECT 31.350 422.400 33.150 429.000 ;
        RECT 34.650 422.400 36.450 428.400 ;
        RECT 47.100 425.400 48.900 429.000 ;
        RECT 50.100 425.400 51.900 428.400 ;
        RECT 53.100 425.400 54.900 429.000 ;
        RECT 65.100 425.400 66.900 429.000 ;
        RECT 68.100 425.400 69.900 428.400 ;
        RECT 11.850 420.000 12.900 421.800 ;
        RECT 22.050 420.000 23.850 420.600 ;
        RECT 11.850 418.800 23.850 420.000 ;
        RECT 4.950 417.600 12.900 418.800 ;
        RECT 4.950 415.050 6.750 417.600 ;
        RECT 11.100 417.000 12.900 417.600 ;
        RECT 8.100 415.800 9.900 416.400 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 8.100 414.600 16.200 415.800 ;
        RECT 14.100 412.950 16.200 414.600 ;
        RECT 12.450 407.700 14.250 408.000 ;
        RECT 2.550 407.100 14.250 407.700 ;
        RECT 2.550 406.500 20.850 407.100 ;
        RECT 2.550 405.600 3.450 406.500 ;
        RECT 12.450 406.200 20.850 406.500 ;
        RECT 2.550 403.800 4.950 405.600 ;
        RECT 3.150 393.600 4.950 403.800 ;
        RECT 6.150 393.000 7.950 405.600 ;
        RECT 17.250 404.700 19.050 405.300 ;
        RECT 11.250 403.500 19.050 404.700 ;
        RECT 19.950 404.100 20.850 406.200 ;
        RECT 22.950 406.200 23.850 418.800 ;
        RECT 35.250 415.050 36.450 422.400 ;
        RECT 50.400 415.050 51.300 425.400 ;
        RECT 68.100 415.050 69.300 425.400 ;
        RECT 71.550 422.400 73.350 428.400 ;
        RECT 74.850 422.400 76.650 429.000 ;
        RECT 79.950 425.400 81.750 428.400 ;
        RECT 84.450 425.400 86.250 429.000 ;
        RECT 87.450 425.400 89.250 428.400 ;
        RECT 90.750 425.400 92.550 429.000 ;
        RECT 95.250 426.300 97.050 428.400 ;
        RECT 95.250 425.400 98.850 426.300 ;
        RECT 79.350 423.300 81.750 425.400 ;
        RECT 88.200 424.500 89.250 425.400 ;
        RECT 95.250 424.800 99.150 425.400 ;
        RECT 88.200 423.450 93.150 424.500 ;
        RECT 91.350 422.700 93.150 423.450 ;
        RECT 71.550 415.050 72.750 422.400 ;
        RECT 94.350 421.800 96.150 423.600 ;
        RECT 97.050 423.300 99.150 424.800 ;
        RECT 100.050 422.400 101.850 429.000 ;
        RECT 103.050 424.200 104.850 428.400 ;
        RECT 103.050 422.400 105.450 424.200 ;
        RECT 84.150 420.000 85.950 420.600 ;
        RECT 95.100 420.000 96.150 421.800 ;
        RECT 84.150 418.800 96.150 420.000 ;
        RECT 30.150 413.250 36.450 415.050 ;
        RECT 31.950 412.950 36.450 413.250 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 64.950 412.950 67.050 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 71.550 413.250 77.850 415.050 ;
        RECT 71.550 412.950 76.050 413.250 ;
        RECT 26.550 410.100 28.650 410.400 ;
        RECT 32.550 410.100 34.350 410.250 ;
        RECT 26.550 408.900 34.350 410.100 ;
        RECT 26.550 408.300 28.650 408.900 ;
        RECT 32.550 408.450 34.350 408.900 ;
        RECT 22.950 405.300 27.750 406.200 ;
        RECT 35.250 405.600 36.450 412.950 ;
        RECT 47.250 411.150 49.050 412.950 ;
        RECT 50.400 405.600 51.300 412.950 ;
        RECT 53.100 411.150 54.900 412.950 ;
        RECT 65.100 411.150 66.900 412.950 ;
        RECT 26.550 404.400 27.750 405.300 ;
        RECT 23.850 404.100 25.650 404.400 ;
        RECT 11.250 402.600 13.350 403.500 ;
        RECT 19.950 403.200 25.650 404.100 ;
        RECT 23.850 402.600 25.650 403.200 ;
        RECT 26.550 402.600 29.550 404.400 ;
        RECT 11.550 393.600 13.350 402.600 ;
        RECT 15.450 401.550 17.250 402.300 ;
        RECT 20.250 401.550 22.050 402.300 ;
        RECT 15.450 400.500 22.050 401.550 ;
        RECT 16.350 393.000 18.150 399.600 ;
        RECT 19.350 393.600 21.150 400.500 ;
        RECT 26.550 399.600 28.650 401.700 ;
        RECT 22.350 393.000 24.150 399.600 ;
        RECT 26.850 393.600 28.650 399.600 ;
        RECT 31.650 393.000 33.450 405.600 ;
        RECT 34.650 393.600 36.450 405.600 ;
        RECT 47.100 393.000 48.900 405.600 ;
        RECT 50.400 404.400 54.000 405.600 ;
        RECT 52.200 393.600 54.000 404.400 ;
        RECT 68.100 399.600 69.300 412.950 ;
        RECT 71.550 405.600 72.750 412.950 ;
        RECT 73.650 410.100 75.450 410.250 ;
        RECT 79.350 410.100 81.450 410.400 ;
        RECT 73.650 408.900 81.450 410.100 ;
        RECT 73.650 408.450 75.450 408.900 ;
        RECT 79.350 408.300 81.450 408.900 ;
        RECT 84.150 406.200 85.050 418.800 ;
        RECT 95.100 417.600 103.050 418.800 ;
        RECT 95.100 417.000 96.900 417.600 ;
        RECT 98.100 415.800 99.900 416.400 ;
        RECT 91.800 414.600 99.900 415.800 ;
        RECT 101.250 415.050 103.050 417.600 ;
        RECT 91.800 412.950 93.900 414.600 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 93.750 407.700 95.550 408.000 ;
        RECT 104.550 407.700 105.450 422.400 ;
        RECT 93.750 407.100 105.450 407.700 ;
        RECT 65.100 393.000 66.900 399.600 ;
        RECT 68.100 393.600 69.900 399.600 ;
        RECT 71.550 393.600 73.350 405.600 ;
        RECT 74.550 393.000 76.350 405.600 ;
        RECT 80.250 405.300 85.050 406.200 ;
        RECT 87.150 406.500 105.450 407.100 ;
        RECT 87.150 406.200 95.550 406.500 ;
        RECT 80.250 404.400 81.450 405.300 ;
        RECT 78.450 402.600 81.450 404.400 ;
        RECT 82.350 404.100 84.150 404.400 ;
        RECT 87.150 404.100 88.050 406.200 ;
        RECT 104.550 405.600 105.450 406.500 ;
        RECT 82.350 403.200 88.050 404.100 ;
        RECT 88.950 404.700 90.750 405.300 ;
        RECT 88.950 403.500 96.750 404.700 ;
        RECT 82.350 402.600 84.150 403.200 ;
        RECT 94.650 402.600 96.750 403.500 ;
        RECT 79.350 399.600 81.450 401.700 ;
        RECT 85.950 401.550 87.750 402.300 ;
        RECT 90.750 401.550 92.550 402.300 ;
        RECT 85.950 400.500 92.550 401.550 ;
        RECT 79.350 393.600 81.150 399.600 ;
        RECT 83.850 393.000 85.650 399.600 ;
        RECT 86.850 393.600 88.650 400.500 ;
        RECT 89.850 393.000 91.650 399.600 ;
        RECT 94.650 393.600 96.450 402.600 ;
        RECT 100.050 393.000 101.850 405.600 ;
        RECT 103.050 403.800 105.450 405.600 ;
        RECT 116.100 422.400 117.900 428.400 ;
        RECT 119.100 422.400 120.900 429.000 ;
        RECT 122.100 425.400 123.900 428.400 ;
        RECT 116.100 415.050 117.300 422.400 ;
        RECT 122.700 421.500 123.900 425.400 ;
        RECT 134.100 422.400 135.900 428.400 ;
        RECT 137.100 423.300 138.900 429.000 ;
        RECT 141.600 422.400 143.400 428.400 ;
        RECT 146.100 423.300 147.900 429.000 ;
        RECT 149.100 422.400 150.900 428.400 ;
        RECT 118.200 420.600 123.900 421.500 ;
        RECT 134.700 420.600 135.900 422.400 ;
        RECT 141.900 420.900 143.100 422.400 ;
        RECT 146.100 421.500 150.900 422.400 ;
        RECT 118.200 419.700 120.000 420.600 ;
        RECT 134.700 419.700 141.000 420.600 ;
        RECT 116.100 412.950 118.200 415.050 ;
        RECT 116.100 405.600 117.300 412.950 ;
        RECT 119.100 408.300 120.000 419.700 ;
        RECT 138.900 417.600 141.000 419.700 ;
        RECT 134.400 415.050 136.200 416.850 ;
        RECT 139.200 415.800 141.000 417.600 ;
        RECT 141.900 418.800 144.900 420.900 ;
        RECT 146.100 420.300 148.200 421.500 ;
        RECT 161.700 421.200 163.500 428.400 ;
        RECT 166.800 422.400 168.600 429.000 ;
        RECT 179.100 423.300 180.900 428.400 ;
        RECT 182.100 424.200 183.900 429.000 ;
        RECT 185.100 423.300 186.900 428.400 ;
        RECT 179.100 421.950 186.900 423.300 ;
        RECT 188.100 422.400 189.900 428.400 ;
        RECT 200.100 425.400 201.900 429.000 ;
        RECT 203.100 425.400 204.900 428.400 ;
        RECT 218.100 425.400 219.900 429.000 ;
        RECT 221.100 425.400 222.900 428.400 ;
        RECT 224.100 425.400 225.900 429.000 ;
        RECT 161.700 420.300 165.900 421.200 ;
        RECT 188.100 420.300 189.300 422.400 ;
        RECT 121.500 412.950 123.600 415.050 ;
        RECT 134.100 414.300 136.200 415.050 ;
        RECT 134.100 412.950 141.000 414.300 ;
        RECT 121.800 411.150 123.600 412.950 ;
        RECT 139.200 412.500 141.000 412.950 ;
        RECT 141.900 413.100 143.100 418.800 ;
        RECT 144.000 415.800 146.100 417.900 ;
        RECT 144.300 414.000 146.100 415.800 ;
        RECT 161.100 415.050 162.900 416.850 ;
        RECT 164.700 415.050 165.900 420.300 ;
        RECT 185.700 419.400 189.300 420.300 ;
        RECT 166.950 415.050 168.750 416.850 ;
        RECT 182.100 415.050 183.900 416.850 ;
        RECT 185.700 415.050 186.900 419.400 ;
        RECT 188.100 415.050 189.900 416.850 ;
        RECT 203.100 415.050 204.300 425.400 ;
        RECT 213.000 417.450 217.050 418.050 ;
        RECT 212.550 415.950 217.050 417.450 ;
        RECT 141.900 412.200 144.300 413.100 ;
        RECT 142.800 412.050 144.300 412.200 ;
        RECT 148.800 412.950 150.900 415.050 ;
        RECT 160.950 412.950 163.050 415.050 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 138.000 409.500 141.900 411.300 ;
        RECT 139.800 409.200 141.900 409.500 ;
        RECT 142.800 409.950 144.900 412.050 ;
        RECT 148.800 411.150 150.600 412.950 ;
        RECT 118.200 407.400 120.000 408.300 ;
        RECT 142.800 408.000 143.700 409.950 ;
        RECT 118.200 406.500 123.900 407.400 ;
        RECT 103.050 393.600 104.850 403.800 ;
        RECT 116.100 393.600 117.900 405.600 ;
        RECT 119.100 393.000 120.900 403.800 ;
        RECT 122.700 399.600 123.900 406.500 ;
        RECT 136.500 405.600 138.600 407.700 ;
        RECT 142.200 406.950 143.700 408.000 ;
        RECT 142.200 405.600 143.400 406.950 ;
        RECT 122.100 393.600 123.900 399.600 ;
        RECT 134.100 404.700 138.600 405.600 ;
        RECT 134.100 393.600 135.900 404.700 ;
        RECT 137.100 393.000 138.900 403.500 ;
        RECT 141.600 393.600 143.400 405.600 ;
        RECT 146.100 405.600 148.200 406.500 ;
        RECT 146.100 404.400 150.900 405.600 ;
        RECT 146.100 393.000 147.900 403.500 ;
        RECT 149.100 393.600 150.900 404.400 ;
        RECT 164.700 399.600 165.900 412.950 ;
        RECT 179.100 411.150 180.900 412.950 ;
        RECT 185.700 405.600 186.900 412.950 ;
        RECT 200.100 411.150 201.900 412.950 ;
        RECT 161.100 393.000 162.900 399.600 ;
        RECT 164.100 393.600 165.900 399.600 ;
        RECT 167.100 393.000 168.900 399.600 ;
        RECT 179.400 393.000 181.200 405.600 ;
        RECT 184.500 404.100 186.900 405.600 ;
        RECT 184.500 393.600 186.300 404.100 ;
        RECT 187.200 401.100 189.000 402.900 ;
        RECT 203.100 399.600 204.300 412.950 ;
        RECT 205.950 411.450 208.050 412.050 ;
        RECT 212.550 411.450 213.450 415.950 ;
        RECT 221.700 415.050 222.600 425.400 ;
        RECT 236.700 421.200 238.500 428.400 ;
        RECT 241.800 422.400 243.600 429.000 ;
        RECT 254.100 425.400 255.900 429.000 ;
        RECT 257.100 425.400 258.900 428.400 ;
        RECT 260.100 425.400 261.900 429.000 ;
        RECT 236.700 420.300 240.900 421.200 ;
        RECT 236.100 415.050 237.900 416.850 ;
        RECT 239.700 415.050 240.900 420.300 ;
        RECT 244.950 417.450 249.000 418.050 ;
        RECT 241.950 415.050 243.750 416.850 ;
        RECT 244.950 415.950 249.450 417.450 ;
        RECT 217.950 412.950 220.050 415.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 235.950 412.950 238.050 415.050 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 205.950 410.550 213.450 411.450 ;
        RECT 218.100 411.150 219.900 412.950 ;
        RECT 205.950 409.950 208.050 410.550 ;
        RECT 221.700 405.600 222.600 412.950 ;
        RECT 223.950 411.150 225.750 412.950 ;
        RECT 219.000 404.400 222.600 405.600 ;
        RECT 187.500 393.000 189.300 399.600 ;
        RECT 200.100 393.000 201.900 399.600 ;
        RECT 203.100 393.600 204.900 399.600 ;
        RECT 219.000 393.600 220.800 404.400 ;
        RECT 224.100 393.000 225.900 405.600 ;
        RECT 239.700 399.600 240.900 412.950 ;
        RECT 248.550 412.050 249.450 415.950 ;
        RECT 257.400 415.050 258.300 425.400 ;
        RECT 263.550 422.400 265.350 428.400 ;
        RECT 266.850 422.400 268.650 429.000 ;
        RECT 271.950 425.400 273.750 428.400 ;
        RECT 276.450 425.400 278.250 429.000 ;
        RECT 279.450 425.400 281.250 428.400 ;
        RECT 282.750 425.400 284.550 429.000 ;
        RECT 287.250 426.300 289.050 428.400 ;
        RECT 287.250 425.400 290.850 426.300 ;
        RECT 271.350 423.300 273.750 425.400 ;
        RECT 280.200 424.500 281.250 425.400 ;
        RECT 287.250 424.800 291.150 425.400 ;
        RECT 280.200 423.450 285.150 424.500 ;
        RECT 283.350 422.700 285.150 423.450 ;
        RECT 263.550 415.050 264.750 422.400 ;
        RECT 286.350 421.800 288.150 423.600 ;
        RECT 289.050 423.300 291.150 424.800 ;
        RECT 292.050 422.400 293.850 429.000 ;
        RECT 295.050 424.200 296.850 428.400 ;
        RECT 295.050 422.400 297.450 424.200 ;
        RECT 276.150 420.000 277.950 420.600 ;
        RECT 287.100 420.000 288.150 421.800 ;
        RECT 276.150 418.800 288.150 420.000 ;
        RECT 253.950 412.950 256.050 415.050 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 259.950 412.950 262.050 415.050 ;
        RECT 263.550 413.250 269.850 415.050 ;
        RECT 263.550 412.950 268.050 413.250 ;
        RECT 248.550 410.550 253.050 412.050 ;
        RECT 254.250 411.150 256.050 412.950 ;
        RECT 249.000 409.950 253.050 410.550 ;
        RECT 257.400 405.600 258.300 412.950 ;
        RECT 260.100 411.150 261.900 412.950 ;
        RECT 263.550 405.600 264.750 412.950 ;
        RECT 265.650 410.100 267.450 410.250 ;
        RECT 271.350 410.100 273.450 410.400 ;
        RECT 265.650 408.900 273.450 410.100 ;
        RECT 265.650 408.450 267.450 408.900 ;
        RECT 271.350 408.300 273.450 408.900 ;
        RECT 276.150 406.200 277.050 418.800 ;
        RECT 287.100 417.600 295.050 418.800 ;
        RECT 287.100 417.000 288.900 417.600 ;
        RECT 290.100 415.800 291.900 416.400 ;
        RECT 283.800 414.600 291.900 415.800 ;
        RECT 293.250 415.050 295.050 417.600 ;
        RECT 283.800 412.950 285.900 414.600 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 285.750 407.700 287.550 408.000 ;
        RECT 296.550 407.700 297.450 422.400 ;
        RECT 308.100 423.300 309.900 428.400 ;
        RECT 311.100 424.200 312.900 429.000 ;
        RECT 314.100 423.300 315.900 428.400 ;
        RECT 308.100 421.950 315.900 423.300 ;
        RECT 317.100 422.400 318.900 428.400 ;
        RECT 329.400 422.400 331.200 429.000 ;
        RECT 317.100 420.300 318.300 422.400 ;
        RECT 334.500 421.200 336.300 428.400 ;
        RECT 347.100 425.400 348.900 429.000 ;
        RECT 350.100 425.400 351.900 428.400 ;
        RECT 314.700 419.400 318.300 420.300 ;
        RECT 311.100 415.050 312.900 416.850 ;
        RECT 314.700 415.050 315.900 419.400 ;
        RECT 325.950 417.450 328.050 421.050 ;
        RECT 323.550 417.000 328.050 417.450 ;
        RECT 332.100 420.300 336.300 421.200 ;
        RECT 317.100 415.050 318.900 416.850 ;
        RECT 323.550 416.550 327.450 417.000 ;
        RECT 307.950 412.950 310.050 415.050 ;
        RECT 310.950 412.950 313.050 415.050 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 308.100 411.150 309.900 412.950 ;
        RECT 285.750 407.100 297.450 407.700 ;
        RECT 236.100 393.000 237.900 399.600 ;
        RECT 239.100 393.600 240.900 399.600 ;
        RECT 242.100 393.000 243.900 399.600 ;
        RECT 254.100 393.000 255.900 405.600 ;
        RECT 257.400 404.400 261.000 405.600 ;
        RECT 259.200 393.600 261.000 404.400 ;
        RECT 263.550 393.600 265.350 405.600 ;
        RECT 266.550 393.000 268.350 405.600 ;
        RECT 272.250 405.300 277.050 406.200 ;
        RECT 279.150 406.500 297.450 407.100 ;
        RECT 279.150 406.200 287.550 406.500 ;
        RECT 272.250 404.400 273.450 405.300 ;
        RECT 270.450 402.600 273.450 404.400 ;
        RECT 274.350 404.100 276.150 404.400 ;
        RECT 279.150 404.100 280.050 406.200 ;
        RECT 296.550 405.600 297.450 406.500 ;
        RECT 314.700 405.600 315.900 412.950 ;
        RECT 323.550 412.050 324.450 416.550 ;
        RECT 329.250 415.050 331.050 416.850 ;
        RECT 332.100 415.050 333.300 420.300 ;
        RECT 335.100 415.050 336.900 416.850 ;
        RECT 350.100 415.050 351.300 425.400 ;
        RECT 353.550 422.400 355.350 428.400 ;
        RECT 356.850 422.400 358.650 429.000 ;
        RECT 361.950 425.400 363.750 428.400 ;
        RECT 366.450 425.400 368.250 429.000 ;
        RECT 369.450 425.400 371.250 428.400 ;
        RECT 372.750 425.400 374.550 429.000 ;
        RECT 377.250 426.300 379.050 428.400 ;
        RECT 377.250 425.400 380.850 426.300 ;
        RECT 361.350 423.300 363.750 425.400 ;
        RECT 370.200 424.500 371.250 425.400 ;
        RECT 377.250 424.800 381.150 425.400 ;
        RECT 370.200 423.450 375.150 424.500 ;
        RECT 373.350 422.700 375.150 423.450 ;
        RECT 353.550 415.050 354.750 422.400 ;
        RECT 376.350 421.800 378.150 423.600 ;
        RECT 379.050 423.300 381.150 424.800 ;
        RECT 382.050 422.400 383.850 429.000 ;
        RECT 385.050 424.200 386.850 428.400 ;
        RECT 385.050 422.400 387.450 424.200 ;
        RECT 366.150 420.000 367.950 420.600 ;
        RECT 377.100 420.000 378.150 421.800 ;
        RECT 366.150 418.800 378.150 420.000 ;
        RECT 328.950 412.950 331.050 415.050 ;
        RECT 331.950 412.950 334.050 415.050 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 353.550 413.250 359.850 415.050 ;
        RECT 353.550 412.950 358.050 413.250 ;
        RECT 319.950 410.550 324.450 412.050 ;
        RECT 319.950 409.950 324.000 410.550 ;
        RECT 274.350 403.200 280.050 404.100 ;
        RECT 280.950 404.700 282.750 405.300 ;
        RECT 280.950 403.500 288.750 404.700 ;
        RECT 274.350 402.600 276.150 403.200 ;
        RECT 286.650 402.600 288.750 403.500 ;
        RECT 271.350 399.600 273.450 401.700 ;
        RECT 277.950 401.550 279.750 402.300 ;
        RECT 282.750 401.550 284.550 402.300 ;
        RECT 277.950 400.500 284.550 401.550 ;
        RECT 271.350 393.600 273.150 399.600 ;
        RECT 275.850 393.000 277.650 399.600 ;
        RECT 278.850 393.600 280.650 400.500 ;
        RECT 281.850 393.000 283.650 399.600 ;
        RECT 286.650 393.600 288.450 402.600 ;
        RECT 292.050 393.000 293.850 405.600 ;
        RECT 295.050 403.800 297.450 405.600 ;
        RECT 295.050 393.600 296.850 403.800 ;
        RECT 308.400 393.000 310.200 405.600 ;
        RECT 313.500 404.100 315.900 405.600 ;
        RECT 313.500 393.600 315.300 404.100 ;
        RECT 316.200 401.100 318.000 402.900 ;
        RECT 332.100 399.600 333.300 412.950 ;
        RECT 347.100 411.150 348.900 412.950 ;
        RECT 350.100 399.600 351.300 412.950 ;
        RECT 353.550 405.600 354.750 412.950 ;
        RECT 355.650 410.100 357.450 410.250 ;
        RECT 361.350 410.100 363.450 410.400 ;
        RECT 355.650 408.900 363.450 410.100 ;
        RECT 355.650 408.450 357.450 408.900 ;
        RECT 361.350 408.300 363.450 408.900 ;
        RECT 366.150 406.200 367.050 418.800 ;
        RECT 377.100 417.600 385.050 418.800 ;
        RECT 377.100 417.000 378.900 417.600 ;
        RECT 380.100 415.800 381.900 416.400 ;
        RECT 373.800 414.600 381.900 415.800 ;
        RECT 383.250 415.050 385.050 417.600 ;
        RECT 373.800 412.950 375.900 414.600 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 375.750 407.700 377.550 408.000 ;
        RECT 386.550 407.700 387.450 422.400 ;
        RECT 398.100 423.300 399.900 428.400 ;
        RECT 401.100 424.200 402.900 429.000 ;
        RECT 404.100 423.300 405.900 428.400 ;
        RECT 398.100 421.950 405.900 423.300 ;
        RECT 407.100 422.400 408.900 428.400 ;
        RECT 422.400 422.400 424.200 429.000 ;
        RECT 388.950 420.450 391.050 421.050 ;
        RECT 394.950 420.450 397.050 421.050 ;
        RECT 388.950 419.550 397.050 420.450 ;
        RECT 407.100 420.300 408.300 422.400 ;
        RECT 427.500 421.200 429.300 428.400 ;
        RECT 388.950 418.950 391.050 419.550 ;
        RECT 394.950 418.950 397.050 419.550 ;
        RECT 404.700 419.400 408.300 420.300 ;
        RECT 425.100 420.300 429.300 421.200 ;
        RECT 440.100 422.400 441.900 428.400 ;
        RECT 443.100 422.400 444.900 429.000 ;
        RECT 446.100 425.400 447.900 428.400 ;
        RECT 401.100 415.050 402.900 416.850 ;
        RECT 404.700 415.050 405.900 419.400 ;
        RECT 407.100 415.050 408.900 416.850 ;
        RECT 422.250 415.050 424.050 416.850 ;
        RECT 425.100 415.050 426.300 420.300 ;
        RECT 428.100 415.050 429.900 416.850 ;
        RECT 440.100 415.050 441.300 422.400 ;
        RECT 446.700 421.500 447.900 425.400 ;
        RECT 442.200 420.600 447.900 421.500 ;
        RECT 449.550 422.400 451.350 428.400 ;
        RECT 452.850 422.400 454.650 429.000 ;
        RECT 457.950 425.400 459.750 428.400 ;
        RECT 462.450 425.400 464.250 429.000 ;
        RECT 465.450 425.400 467.250 428.400 ;
        RECT 468.750 425.400 470.550 429.000 ;
        RECT 473.250 426.300 475.050 428.400 ;
        RECT 473.250 425.400 476.850 426.300 ;
        RECT 457.350 423.300 459.750 425.400 ;
        RECT 466.200 424.500 467.250 425.400 ;
        RECT 473.250 424.800 477.150 425.400 ;
        RECT 466.200 423.450 471.150 424.500 ;
        RECT 469.350 422.700 471.150 423.450 ;
        RECT 442.200 419.700 444.000 420.600 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 440.100 412.950 442.200 415.050 ;
        RECT 398.100 411.150 399.900 412.950 ;
        RECT 375.750 407.100 387.450 407.700 ;
        RECT 316.500 393.000 318.300 399.600 ;
        RECT 329.100 393.000 330.900 399.600 ;
        RECT 332.100 393.600 333.900 399.600 ;
        RECT 335.100 393.000 336.900 399.600 ;
        RECT 347.100 393.000 348.900 399.600 ;
        RECT 350.100 393.600 351.900 399.600 ;
        RECT 353.550 393.600 355.350 405.600 ;
        RECT 356.550 393.000 358.350 405.600 ;
        RECT 362.250 405.300 367.050 406.200 ;
        RECT 369.150 406.500 387.450 407.100 ;
        RECT 369.150 406.200 377.550 406.500 ;
        RECT 362.250 404.400 363.450 405.300 ;
        RECT 360.450 402.600 363.450 404.400 ;
        RECT 364.350 404.100 366.150 404.400 ;
        RECT 369.150 404.100 370.050 406.200 ;
        RECT 386.550 405.600 387.450 406.500 ;
        RECT 404.700 405.600 405.900 412.950 ;
        RECT 364.350 403.200 370.050 404.100 ;
        RECT 370.950 404.700 372.750 405.300 ;
        RECT 370.950 403.500 378.750 404.700 ;
        RECT 364.350 402.600 366.150 403.200 ;
        RECT 376.650 402.600 378.750 403.500 ;
        RECT 361.350 399.600 363.450 401.700 ;
        RECT 367.950 401.550 369.750 402.300 ;
        RECT 372.750 401.550 374.550 402.300 ;
        RECT 367.950 400.500 374.550 401.550 ;
        RECT 361.350 393.600 363.150 399.600 ;
        RECT 365.850 393.000 367.650 399.600 ;
        RECT 368.850 393.600 370.650 400.500 ;
        RECT 371.850 393.000 373.650 399.600 ;
        RECT 376.650 393.600 378.450 402.600 ;
        RECT 382.050 393.000 383.850 405.600 ;
        RECT 385.050 403.800 387.450 405.600 ;
        RECT 385.050 393.600 386.850 403.800 ;
        RECT 398.400 393.000 400.200 405.600 ;
        RECT 403.500 404.100 405.900 405.600 ;
        RECT 403.500 393.600 405.300 404.100 ;
        RECT 406.200 401.100 408.000 402.900 ;
        RECT 425.100 399.600 426.300 412.950 ;
        RECT 440.100 405.600 441.300 412.950 ;
        RECT 443.100 408.300 444.000 419.700 ;
        RECT 449.550 415.050 450.750 422.400 ;
        RECT 472.350 421.800 474.150 423.600 ;
        RECT 475.050 423.300 477.150 424.800 ;
        RECT 478.050 422.400 479.850 429.000 ;
        RECT 481.050 424.200 482.850 428.400 ;
        RECT 481.050 422.400 483.450 424.200 ;
        RECT 462.150 420.000 463.950 420.600 ;
        RECT 473.100 420.000 474.150 421.800 ;
        RECT 462.150 418.800 474.150 420.000 ;
        RECT 445.500 412.950 447.600 415.050 ;
        RECT 445.800 411.150 447.600 412.950 ;
        RECT 449.550 413.250 455.850 415.050 ;
        RECT 449.550 412.950 454.050 413.250 ;
        RECT 442.200 407.400 444.000 408.300 ;
        RECT 442.200 406.500 447.900 407.400 ;
        RECT 406.500 393.000 408.300 399.600 ;
        RECT 422.100 393.000 423.900 399.600 ;
        RECT 425.100 393.600 426.900 399.600 ;
        RECT 428.100 393.000 429.900 399.600 ;
        RECT 440.100 393.600 441.900 405.600 ;
        RECT 443.100 393.000 444.900 403.800 ;
        RECT 446.700 399.600 447.900 406.500 ;
        RECT 446.100 393.600 447.900 399.600 ;
        RECT 449.550 405.600 450.750 412.950 ;
        RECT 451.650 410.100 453.450 410.250 ;
        RECT 457.350 410.100 459.450 410.400 ;
        RECT 451.650 408.900 459.450 410.100 ;
        RECT 451.650 408.450 453.450 408.900 ;
        RECT 457.350 408.300 459.450 408.900 ;
        RECT 462.150 406.200 463.050 418.800 ;
        RECT 473.100 417.600 481.050 418.800 ;
        RECT 473.100 417.000 474.900 417.600 ;
        RECT 476.100 415.800 477.900 416.400 ;
        RECT 469.800 414.600 477.900 415.800 ;
        RECT 479.250 415.050 481.050 417.600 ;
        RECT 469.800 412.950 471.900 414.600 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 471.750 407.700 473.550 408.000 ;
        RECT 482.550 407.700 483.450 422.400 ;
        RECT 471.750 407.100 483.450 407.700 ;
        RECT 449.550 393.600 451.350 405.600 ;
        RECT 452.550 393.000 454.350 405.600 ;
        RECT 458.250 405.300 463.050 406.200 ;
        RECT 465.150 406.500 483.450 407.100 ;
        RECT 465.150 406.200 473.550 406.500 ;
        RECT 458.250 404.400 459.450 405.300 ;
        RECT 456.450 402.600 459.450 404.400 ;
        RECT 460.350 404.100 462.150 404.400 ;
        RECT 465.150 404.100 466.050 406.200 ;
        RECT 482.550 405.600 483.450 406.500 ;
        RECT 460.350 403.200 466.050 404.100 ;
        RECT 466.950 404.700 468.750 405.300 ;
        RECT 466.950 403.500 474.750 404.700 ;
        RECT 460.350 402.600 462.150 403.200 ;
        RECT 472.650 402.600 474.750 403.500 ;
        RECT 457.350 399.600 459.450 401.700 ;
        RECT 463.950 401.550 465.750 402.300 ;
        RECT 468.750 401.550 470.550 402.300 ;
        RECT 463.950 400.500 470.550 401.550 ;
        RECT 457.350 393.600 459.150 399.600 ;
        RECT 461.850 393.000 463.650 399.600 ;
        RECT 464.850 393.600 466.650 400.500 ;
        RECT 467.850 393.000 469.650 399.600 ;
        RECT 472.650 393.600 474.450 402.600 ;
        RECT 478.050 393.000 479.850 405.600 ;
        RECT 481.050 403.800 483.450 405.600 ;
        RECT 494.100 422.400 495.900 428.400 ;
        RECT 497.100 422.400 498.900 429.000 ;
        RECT 500.100 425.400 501.900 428.400 ;
        RECT 494.100 415.050 495.300 422.400 ;
        RECT 500.700 421.500 501.900 425.400 ;
        RECT 496.200 420.600 501.900 421.500 ;
        RECT 503.550 422.400 505.350 428.400 ;
        RECT 506.850 422.400 508.650 429.000 ;
        RECT 511.950 425.400 513.750 428.400 ;
        RECT 516.450 425.400 518.250 429.000 ;
        RECT 519.450 425.400 521.250 428.400 ;
        RECT 522.750 425.400 524.550 429.000 ;
        RECT 527.250 426.300 529.050 428.400 ;
        RECT 527.250 425.400 530.850 426.300 ;
        RECT 511.350 423.300 513.750 425.400 ;
        RECT 520.200 424.500 521.250 425.400 ;
        RECT 527.250 424.800 531.150 425.400 ;
        RECT 520.200 423.450 525.150 424.500 ;
        RECT 523.350 422.700 525.150 423.450 ;
        RECT 496.200 419.700 498.000 420.600 ;
        RECT 494.100 412.950 496.200 415.050 ;
        RECT 494.100 405.600 495.300 412.950 ;
        RECT 497.100 408.300 498.000 419.700 ;
        RECT 503.550 415.050 504.750 422.400 ;
        RECT 526.350 421.800 528.150 423.600 ;
        RECT 529.050 423.300 531.150 424.800 ;
        RECT 532.050 422.400 533.850 429.000 ;
        RECT 535.050 424.200 536.850 428.400 ;
        RECT 535.050 422.400 537.450 424.200 ;
        RECT 516.150 420.000 517.950 420.600 ;
        RECT 527.100 420.000 528.150 421.800 ;
        RECT 516.150 418.800 528.150 420.000 ;
        RECT 499.500 412.950 501.600 415.050 ;
        RECT 499.800 411.150 501.600 412.950 ;
        RECT 503.550 413.250 509.850 415.050 ;
        RECT 503.550 412.950 508.050 413.250 ;
        RECT 496.200 407.400 498.000 408.300 ;
        RECT 496.200 406.500 501.900 407.400 ;
        RECT 481.050 393.600 482.850 403.800 ;
        RECT 494.100 393.600 495.900 405.600 ;
        RECT 497.100 393.000 498.900 403.800 ;
        RECT 500.700 399.600 501.900 406.500 ;
        RECT 500.100 393.600 501.900 399.600 ;
        RECT 503.550 405.600 504.750 412.950 ;
        RECT 505.650 410.100 507.450 410.250 ;
        RECT 511.350 410.100 513.450 410.400 ;
        RECT 505.650 408.900 513.450 410.100 ;
        RECT 505.650 408.450 507.450 408.900 ;
        RECT 511.350 408.300 513.450 408.900 ;
        RECT 516.150 406.200 517.050 418.800 ;
        RECT 527.100 417.600 535.050 418.800 ;
        RECT 527.100 417.000 528.900 417.600 ;
        RECT 530.100 415.800 531.900 416.400 ;
        RECT 523.800 414.600 531.900 415.800 ;
        RECT 533.250 415.050 535.050 417.600 ;
        RECT 523.800 412.950 525.900 414.600 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 525.750 407.700 527.550 408.000 ;
        RECT 536.550 407.700 537.450 422.400 ;
        RECT 525.750 407.100 537.450 407.700 ;
        RECT 503.550 393.600 505.350 405.600 ;
        RECT 506.550 393.000 508.350 405.600 ;
        RECT 512.250 405.300 517.050 406.200 ;
        RECT 519.150 406.500 537.450 407.100 ;
        RECT 519.150 406.200 527.550 406.500 ;
        RECT 512.250 404.400 513.450 405.300 ;
        RECT 510.450 402.600 513.450 404.400 ;
        RECT 514.350 404.100 516.150 404.400 ;
        RECT 519.150 404.100 520.050 406.200 ;
        RECT 536.550 405.600 537.450 406.500 ;
        RECT 514.350 403.200 520.050 404.100 ;
        RECT 520.950 404.700 522.750 405.300 ;
        RECT 520.950 403.500 528.750 404.700 ;
        RECT 514.350 402.600 516.150 403.200 ;
        RECT 526.650 402.600 528.750 403.500 ;
        RECT 511.350 399.600 513.450 401.700 ;
        RECT 517.950 401.550 519.750 402.300 ;
        RECT 522.750 401.550 524.550 402.300 ;
        RECT 517.950 400.500 524.550 401.550 ;
        RECT 511.350 393.600 513.150 399.600 ;
        RECT 515.850 393.000 517.650 399.600 ;
        RECT 518.850 393.600 520.650 400.500 ;
        RECT 521.850 393.000 523.650 399.600 ;
        RECT 526.650 393.600 528.450 402.600 ;
        RECT 532.050 393.000 533.850 405.600 ;
        RECT 535.050 403.800 537.450 405.600 ;
        RECT 548.100 422.400 549.900 428.400 ;
        RECT 551.100 422.400 552.900 429.000 ;
        RECT 554.100 425.400 555.900 428.400 ;
        RECT 548.100 415.050 549.300 422.400 ;
        RECT 554.700 421.500 555.900 425.400 ;
        RECT 550.200 420.600 555.900 421.500 ;
        RECT 557.550 422.400 559.350 428.400 ;
        RECT 560.850 422.400 562.650 429.000 ;
        RECT 565.950 425.400 567.750 428.400 ;
        RECT 570.450 425.400 572.250 429.000 ;
        RECT 573.450 425.400 575.250 428.400 ;
        RECT 576.750 425.400 578.550 429.000 ;
        RECT 581.250 426.300 583.050 428.400 ;
        RECT 581.250 425.400 584.850 426.300 ;
        RECT 565.350 423.300 567.750 425.400 ;
        RECT 574.200 424.500 575.250 425.400 ;
        RECT 581.250 424.800 585.150 425.400 ;
        RECT 574.200 423.450 579.150 424.500 ;
        RECT 577.350 422.700 579.150 423.450 ;
        RECT 550.200 419.700 552.000 420.600 ;
        RECT 548.100 412.950 550.200 415.050 ;
        RECT 548.100 405.600 549.300 412.950 ;
        RECT 551.100 408.300 552.000 419.700 ;
        RECT 557.550 415.050 558.750 422.400 ;
        RECT 580.350 421.800 582.150 423.600 ;
        RECT 583.050 423.300 585.150 424.800 ;
        RECT 586.050 422.400 587.850 429.000 ;
        RECT 589.050 424.200 590.850 428.400 ;
        RECT 589.050 422.400 591.450 424.200 ;
        RECT 570.150 420.000 571.950 420.600 ;
        RECT 581.100 420.000 582.150 421.800 ;
        RECT 570.150 418.800 582.150 420.000 ;
        RECT 553.500 412.950 555.600 415.050 ;
        RECT 553.800 411.150 555.600 412.950 ;
        RECT 557.550 413.250 563.850 415.050 ;
        RECT 557.550 412.950 562.050 413.250 ;
        RECT 550.200 407.400 552.000 408.300 ;
        RECT 550.200 406.500 555.900 407.400 ;
        RECT 535.050 393.600 536.850 403.800 ;
        RECT 548.100 393.600 549.900 405.600 ;
        RECT 551.100 393.000 552.900 403.800 ;
        RECT 554.700 399.600 555.900 406.500 ;
        RECT 554.100 393.600 555.900 399.600 ;
        RECT 557.550 405.600 558.750 412.950 ;
        RECT 559.650 410.100 561.450 410.250 ;
        RECT 565.350 410.100 567.450 410.400 ;
        RECT 559.650 408.900 567.450 410.100 ;
        RECT 559.650 408.450 561.450 408.900 ;
        RECT 565.350 408.300 567.450 408.900 ;
        RECT 570.150 406.200 571.050 418.800 ;
        RECT 581.100 417.600 589.050 418.800 ;
        RECT 581.100 417.000 582.900 417.600 ;
        RECT 584.100 415.800 585.900 416.400 ;
        RECT 577.800 414.600 585.900 415.800 ;
        RECT 587.250 415.050 589.050 417.600 ;
        RECT 577.800 412.950 579.900 414.600 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 579.750 407.700 581.550 408.000 ;
        RECT 590.550 407.700 591.450 422.400 ;
        RECT 602.100 423.300 603.900 428.400 ;
        RECT 605.100 424.200 606.900 429.000 ;
        RECT 608.100 423.300 609.900 428.400 ;
        RECT 602.100 421.950 609.900 423.300 ;
        RECT 611.100 422.400 612.900 428.400 ;
        RECT 611.100 420.300 612.300 422.400 ;
        RECT 623.700 421.200 625.500 428.400 ;
        RECT 628.800 422.400 630.600 429.000 ;
        RECT 641.100 422.400 642.900 429.000 ;
        RECT 644.100 422.400 645.900 428.400 ;
        RECT 656.100 422.400 657.900 428.400 ;
        RECT 659.100 422.400 660.900 429.000 ;
        RECT 623.700 420.300 627.900 421.200 ;
        RECT 608.700 419.400 612.300 420.300 ;
        RECT 605.100 415.050 606.900 416.850 ;
        RECT 608.700 415.050 609.900 419.400 ;
        RECT 611.100 415.050 612.900 416.850 ;
        RECT 623.100 415.050 624.900 416.850 ;
        RECT 626.700 415.050 627.900 420.300 ;
        RECT 628.950 415.050 630.750 416.850 ;
        RECT 641.100 415.050 642.900 416.850 ;
        RECT 644.100 415.050 645.300 422.400 ;
        RECT 656.700 415.050 657.900 422.400 ;
        RECT 671.700 421.200 673.500 428.400 ;
        RECT 676.800 422.400 678.600 429.000 ;
        RECT 689.100 423.300 690.900 428.400 ;
        RECT 692.100 424.200 693.900 429.000 ;
        RECT 695.100 423.300 696.900 428.400 ;
        RECT 689.100 421.950 696.900 423.300 ;
        RECT 698.100 422.400 699.900 428.400 ;
        RECT 710.100 423.300 711.900 428.400 ;
        RECT 713.100 424.200 714.900 429.000 ;
        RECT 716.100 423.300 717.900 428.400 ;
        RECT 671.700 420.300 675.900 421.200 ;
        RECT 698.100 420.300 699.300 422.400 ;
        RECT 710.100 421.950 717.900 423.300 ;
        RECT 719.100 422.400 720.900 428.400 ;
        RECT 731.100 425.400 732.900 429.000 ;
        RECT 746.100 428.400 747.300 429.000 ;
        RECT 734.100 425.400 735.900 428.400 ;
        RECT 719.100 420.300 720.300 422.400 ;
        RECT 659.100 415.050 660.900 416.850 ;
        RECT 671.100 415.050 672.900 416.850 ;
        RECT 674.700 415.050 675.900 420.300 ;
        RECT 695.700 419.400 699.300 420.300 ;
        RECT 716.700 419.400 720.300 420.300 ;
        RECT 676.950 415.050 678.750 416.850 ;
        RECT 692.100 415.050 693.900 416.850 ;
        RECT 695.700 415.050 696.900 419.400 ;
        RECT 698.100 415.050 699.900 416.850 ;
        RECT 713.100 415.050 714.900 416.850 ;
        RECT 716.700 415.050 717.900 419.400 ;
        RECT 719.100 415.050 720.900 416.850 ;
        RECT 734.100 415.050 735.300 425.400 ;
        RECT 736.950 423.450 739.050 427.050 ;
        RECT 746.100 425.400 747.900 428.400 ;
        RECT 749.100 425.400 750.900 428.400 ;
        RECT 745.950 423.450 748.050 424.050 ;
        RECT 736.950 423.000 748.050 423.450 ;
        RECT 737.550 422.550 748.050 423.000 ;
        RECT 745.950 421.950 748.050 422.550 ;
        RECT 749.400 421.200 750.300 425.400 ;
        RECT 752.100 423.000 753.900 429.000 ;
        RECT 767.100 428.400 768.300 429.000 ;
        RECT 755.100 422.400 756.900 428.400 ;
        RECT 767.100 425.400 768.900 428.400 ;
        RECT 770.100 425.400 771.900 428.400 ;
        RECT 749.400 420.300 754.800 421.200 ;
        RECT 752.700 419.400 754.800 420.300 ;
        RECT 746.400 415.050 748.200 416.850 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 746.100 412.950 748.200 415.050 ;
        RECT 749.400 412.950 751.500 415.050 ;
        RECT 602.100 411.150 603.900 412.950 ;
        RECT 579.750 407.100 591.450 407.700 ;
        RECT 557.550 393.600 559.350 405.600 ;
        RECT 560.550 393.000 562.350 405.600 ;
        RECT 566.250 405.300 571.050 406.200 ;
        RECT 573.150 406.500 591.450 407.100 ;
        RECT 573.150 406.200 581.550 406.500 ;
        RECT 566.250 404.400 567.450 405.300 ;
        RECT 564.450 402.600 567.450 404.400 ;
        RECT 568.350 404.100 570.150 404.400 ;
        RECT 573.150 404.100 574.050 406.200 ;
        RECT 590.550 405.600 591.450 406.500 ;
        RECT 608.700 405.600 609.900 412.950 ;
        RECT 610.950 408.450 613.050 409.050 ;
        RECT 616.950 408.450 619.050 409.050 ;
        RECT 610.950 407.550 619.050 408.450 ;
        RECT 610.950 406.950 613.050 407.550 ;
        RECT 616.950 406.950 619.050 407.550 ;
        RECT 568.350 403.200 574.050 404.100 ;
        RECT 574.950 404.700 576.750 405.300 ;
        RECT 574.950 403.500 582.750 404.700 ;
        RECT 568.350 402.600 570.150 403.200 ;
        RECT 580.650 402.600 582.750 403.500 ;
        RECT 565.350 399.600 567.450 401.700 ;
        RECT 571.950 401.550 573.750 402.300 ;
        RECT 576.750 401.550 578.550 402.300 ;
        RECT 571.950 400.500 578.550 401.550 ;
        RECT 565.350 393.600 567.150 399.600 ;
        RECT 569.850 393.000 571.650 399.600 ;
        RECT 572.850 393.600 574.650 400.500 ;
        RECT 575.850 393.000 577.650 399.600 ;
        RECT 580.650 393.600 582.450 402.600 ;
        RECT 586.050 393.000 587.850 405.600 ;
        RECT 589.050 403.800 591.450 405.600 ;
        RECT 589.050 393.600 590.850 403.800 ;
        RECT 602.400 393.000 604.200 405.600 ;
        RECT 607.500 404.100 609.900 405.600 ;
        RECT 607.500 393.600 609.300 404.100 ;
        RECT 610.200 401.100 612.000 402.900 ;
        RECT 626.700 399.600 627.900 412.950 ;
        RECT 644.100 405.600 645.300 412.950 ;
        RECT 656.700 405.600 657.900 412.950 ;
        RECT 610.500 393.000 612.300 399.600 ;
        RECT 623.100 393.000 624.900 399.600 ;
        RECT 626.100 393.600 627.900 399.600 ;
        RECT 629.100 393.000 630.900 399.600 ;
        RECT 641.100 393.000 642.900 405.600 ;
        RECT 644.100 393.600 645.900 405.600 ;
        RECT 656.100 393.600 657.900 405.600 ;
        RECT 659.100 393.000 660.900 405.600 ;
        RECT 674.700 399.600 675.900 412.950 ;
        RECT 689.100 411.150 690.900 412.950 ;
        RECT 695.700 405.600 696.900 412.950 ;
        RECT 710.100 411.150 711.900 412.950 ;
        RECT 716.700 405.600 717.900 412.950 ;
        RECT 731.100 411.150 732.900 412.950 ;
        RECT 671.100 393.000 672.900 399.600 ;
        RECT 674.100 393.600 675.900 399.600 ;
        RECT 677.100 393.000 678.900 399.600 ;
        RECT 689.400 393.000 691.200 405.600 ;
        RECT 694.500 404.100 696.900 405.600 ;
        RECT 694.500 393.600 696.300 404.100 ;
        RECT 697.200 401.100 699.000 402.900 ;
        RECT 697.500 393.000 699.300 399.600 ;
        RECT 710.400 393.000 712.200 405.600 ;
        RECT 715.500 404.100 717.900 405.600 ;
        RECT 715.500 393.600 717.300 404.100 ;
        RECT 718.200 401.100 720.000 402.900 ;
        RECT 734.100 399.600 735.300 412.950 ;
        RECT 750.000 411.150 751.800 412.950 ;
        RECT 752.700 408.900 753.600 419.400 ;
        RECT 756.000 415.050 756.900 422.400 ;
        RECT 770.400 421.200 771.300 425.400 ;
        RECT 773.100 423.000 774.900 429.000 ;
        RECT 776.100 422.400 777.900 428.400 ;
        RECT 770.400 420.300 775.800 421.200 ;
        RECT 773.700 419.400 775.800 420.300 ;
        RECT 767.400 415.050 769.200 416.850 ;
        RECT 754.800 412.950 756.900 415.050 ;
        RECT 767.100 412.950 769.200 415.050 ;
        RECT 770.400 412.950 772.500 415.050 ;
        RECT 752.100 408.300 753.900 408.900 ;
        RECT 746.100 407.100 753.900 408.300 ;
        RECT 746.100 405.600 747.300 407.100 ;
        RECT 754.800 405.600 756.000 412.950 ;
        RECT 771.000 411.150 772.800 412.950 ;
        RECT 773.700 408.900 774.600 419.400 ;
        RECT 777.000 415.050 777.900 422.400 ;
        RECT 788.100 420.600 789.900 428.400 ;
        RECT 792.600 422.400 794.400 429.000 ;
        RECT 795.600 424.200 797.400 428.400 ;
        RECT 795.600 422.400 798.300 424.200 ;
        RECT 809.400 422.400 811.200 429.000 ;
        RECT 794.700 420.600 796.500 421.500 ;
        RECT 788.100 419.700 796.500 420.600 ;
        RECT 788.250 415.050 790.050 416.850 ;
        RECT 775.800 412.950 777.900 415.050 ;
        RECT 788.100 412.950 790.200 415.050 ;
        RECT 773.100 408.300 774.900 408.900 ;
        RECT 718.500 393.000 720.300 399.600 ;
        RECT 731.100 393.000 732.900 399.600 ;
        RECT 734.100 393.600 735.900 399.600 ;
        RECT 746.100 393.600 747.900 405.600 ;
        RECT 750.600 393.000 752.400 405.600 ;
        RECT 753.600 404.100 756.000 405.600 ;
        RECT 767.100 407.100 774.900 408.300 ;
        RECT 767.100 405.600 768.300 407.100 ;
        RECT 775.800 405.600 777.000 412.950 ;
        RECT 753.600 393.600 755.400 404.100 ;
        RECT 767.100 393.600 768.900 405.600 ;
        RECT 771.600 393.000 773.400 405.600 ;
        RECT 774.600 404.100 777.000 405.600 ;
        RECT 774.600 393.600 776.400 404.100 ;
        RECT 791.100 399.600 792.000 419.700 ;
        RECT 797.400 415.050 798.300 422.400 ;
        RECT 814.500 421.200 816.300 428.400 ;
        RECT 827.100 422.400 828.900 428.400 ;
        RECT 830.400 423.300 832.200 429.000 ;
        RECT 834.900 423.000 836.700 428.400 ;
        RECT 839.100 423.300 840.900 429.000 ;
        RECT 827.100 421.500 831.600 422.400 ;
        RECT 812.100 420.300 816.300 421.200 ;
        RECT 809.250 415.050 811.050 416.850 ;
        RECT 812.100 415.050 813.300 420.300 ;
        RECT 829.500 419.100 831.600 421.500 ;
        RECT 834.900 420.900 835.800 423.000 ;
        RECT 842.100 422.400 843.900 428.400 ;
        RECT 854.700 425.400 856.500 429.000 ;
        RECT 857.700 423.600 859.500 428.400 ;
        RECT 842.400 421.500 843.900 422.400 ;
        RECT 832.800 418.800 835.800 420.900 ;
        RECT 839.400 420.000 843.900 421.500 ;
        RECT 854.400 422.400 859.500 423.600 ;
        RECT 862.200 422.400 864.000 429.000 ;
        RECT 815.100 415.050 816.900 416.850 ;
        RECT 793.500 412.950 795.600 415.050 ;
        RECT 796.800 412.950 798.900 415.050 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 827.100 412.950 829.200 415.050 ;
        RECT 831.900 414.900 834.000 417.000 ;
        RECT 832.200 413.100 834.000 414.900 ;
        RECT 793.200 411.150 795.000 412.950 ;
        RECT 797.400 405.600 798.300 412.950 ;
        RECT 788.100 393.000 789.900 399.600 ;
        RECT 791.100 393.600 792.900 399.600 ;
        RECT 794.100 393.000 795.900 405.000 ;
        RECT 797.100 393.600 798.900 405.600 ;
        RECT 812.100 399.600 813.300 412.950 ;
        RECT 827.400 411.150 829.200 412.950 ;
        RECT 834.900 412.050 835.800 418.800 ;
        RECT 836.700 417.900 838.500 419.700 ;
        RECT 839.400 419.400 841.500 420.000 ;
        RECT 837.000 417.000 839.100 417.900 ;
        RECT 837.000 415.800 843.600 417.000 ;
        RECT 841.800 415.200 843.600 415.800 ;
        RECT 837.000 412.800 839.100 414.900 ;
        RECT 841.800 412.950 843.900 415.200 ;
        RECT 854.400 415.050 855.300 422.400 ;
        RECT 856.950 415.050 858.750 416.850 ;
        RECT 863.100 415.050 864.900 416.850 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 832.800 410.700 835.800 412.050 ;
        RECT 837.300 411.000 839.100 412.800 ;
        RECT 832.800 409.950 834.900 410.700 ;
        RECT 830.100 405.600 832.200 406.500 ;
        RECT 827.100 404.400 832.200 405.600 ;
        RECT 833.100 405.600 834.300 409.950 ;
        RECT 835.800 407.700 837.600 409.500 ;
        RECT 835.800 406.800 841.200 407.700 ;
        RECT 839.100 405.900 841.200 406.800 ;
        RECT 833.100 404.700 836.400 405.600 ;
        RECT 839.100 404.700 843.900 405.900 ;
        RECT 854.400 405.600 855.300 412.950 ;
        RECT 859.950 411.150 861.750 412.950 ;
        RECT 865.950 411.450 868.050 412.050 ;
        RECT 871.950 411.450 874.050 412.050 ;
        RECT 865.950 410.550 874.050 411.450 ;
        RECT 865.950 409.950 868.050 410.550 ;
        RECT 871.950 409.950 874.050 410.550 ;
        RECT 809.100 393.000 810.900 399.600 ;
        RECT 812.100 393.600 813.900 399.600 ;
        RECT 815.100 393.000 816.900 399.600 ;
        RECT 827.100 393.600 828.900 404.400 ;
        RECT 830.100 393.000 832.200 403.500 ;
        RECT 834.600 393.600 836.400 404.700 ;
        RECT 839.100 393.000 840.900 403.500 ;
        RECT 842.100 393.600 843.900 404.700 ;
        RECT 854.100 393.600 855.900 405.600 ;
        RECT 857.100 404.700 864.900 405.600 ;
        RECT 857.100 393.600 858.900 404.700 ;
        RECT 860.100 393.000 861.900 403.800 ;
        RECT 863.100 393.600 864.900 404.700 ;
        RECT 11.100 383.400 12.900 389.400 ;
        RECT 14.100 383.400 15.900 390.000 ;
        RECT 11.700 370.050 12.900 383.400 ;
        RECT 17.550 377.400 19.350 389.400 ;
        RECT 20.550 377.400 22.350 390.000 ;
        RECT 25.350 383.400 27.150 389.400 ;
        RECT 29.850 383.400 31.650 390.000 ;
        RECT 25.350 381.300 27.450 383.400 ;
        RECT 32.850 382.500 34.650 389.400 ;
        RECT 35.850 383.400 37.650 390.000 ;
        RECT 31.950 381.450 38.550 382.500 ;
        RECT 31.950 380.700 33.750 381.450 ;
        RECT 36.750 380.700 38.550 381.450 ;
        RECT 40.650 380.400 42.450 389.400 ;
        RECT 24.450 378.600 27.450 380.400 ;
        RECT 28.350 379.800 30.150 380.400 ;
        RECT 28.350 378.900 34.050 379.800 ;
        RECT 40.650 379.500 42.750 380.400 ;
        RECT 28.350 378.600 30.150 378.900 ;
        RECT 26.250 377.700 27.450 378.600 ;
        RECT 14.100 370.050 15.900 371.850 ;
        RECT 17.550 370.050 18.750 377.400 ;
        RECT 26.250 376.800 31.050 377.700 ;
        RECT 19.650 374.100 21.450 374.550 ;
        RECT 25.350 374.100 27.450 374.700 ;
        RECT 19.650 372.900 27.450 374.100 ;
        RECT 19.650 372.750 21.450 372.900 ;
        RECT 25.350 372.600 27.450 372.900 ;
        RECT 10.950 367.950 13.050 370.050 ;
        RECT 13.950 367.950 16.050 370.050 ;
        RECT 17.550 369.750 22.050 370.050 ;
        RECT 17.550 367.950 23.850 369.750 ;
        RECT 11.700 357.600 12.900 367.950 ;
        RECT 17.550 360.600 18.750 367.950 ;
        RECT 30.150 364.200 31.050 376.800 ;
        RECT 33.150 376.800 34.050 378.900 ;
        RECT 34.950 378.300 42.750 379.500 ;
        RECT 34.950 377.700 36.750 378.300 ;
        RECT 46.050 377.400 47.850 390.000 ;
        RECT 49.050 379.200 50.850 389.400 ;
        RECT 54.150 379.200 55.950 389.400 ;
        RECT 49.050 377.400 51.450 379.200 ;
        RECT 33.150 376.500 41.550 376.800 ;
        RECT 50.550 376.500 51.450 377.400 ;
        RECT 33.150 375.900 51.450 376.500 ;
        RECT 39.750 375.300 51.450 375.900 ;
        RECT 39.750 375.000 41.550 375.300 ;
        RECT 37.800 368.400 39.900 370.050 ;
        RECT 37.800 367.200 45.900 368.400 ;
        RECT 46.950 367.950 49.050 370.050 ;
        RECT 44.100 366.600 45.900 367.200 ;
        RECT 41.100 365.400 42.900 366.000 ;
        RECT 47.250 365.400 49.050 367.950 ;
        RECT 41.100 364.200 49.050 365.400 ;
        RECT 30.150 363.000 42.150 364.200 ;
        RECT 30.150 362.400 31.950 363.000 ;
        RECT 41.100 361.200 42.150 363.000 ;
        RECT 11.100 354.600 12.900 357.600 ;
        RECT 14.100 354.000 15.900 357.600 ;
        RECT 17.550 354.600 19.350 360.600 ;
        RECT 20.850 354.000 22.650 360.600 ;
        RECT 25.350 357.600 27.750 359.700 ;
        RECT 37.350 359.550 39.150 360.300 ;
        RECT 34.200 358.500 39.150 359.550 ;
        RECT 40.350 359.400 42.150 361.200 ;
        RECT 50.550 360.600 51.450 375.300 ;
        RECT 34.200 357.600 35.250 358.500 ;
        RECT 43.050 358.200 45.150 359.700 ;
        RECT 41.250 357.600 45.150 358.200 ;
        RECT 25.950 354.600 27.750 357.600 ;
        RECT 30.450 354.000 32.250 357.600 ;
        RECT 33.450 354.600 35.250 357.600 ;
        RECT 36.750 354.000 38.550 357.600 ;
        RECT 41.250 356.700 44.850 357.600 ;
        RECT 41.250 354.600 43.050 356.700 ;
        RECT 46.050 354.000 47.850 360.600 ;
        RECT 49.050 358.800 51.450 360.600 ;
        RECT 53.550 377.400 55.950 379.200 ;
        RECT 57.150 377.400 58.950 390.000 ;
        RECT 62.550 380.400 64.350 389.400 ;
        RECT 67.350 383.400 69.150 390.000 ;
        RECT 70.350 382.500 72.150 389.400 ;
        RECT 73.350 383.400 75.150 390.000 ;
        RECT 77.850 383.400 79.650 389.400 ;
        RECT 66.450 381.450 73.050 382.500 ;
        RECT 66.450 380.700 68.250 381.450 ;
        RECT 71.250 380.700 73.050 381.450 ;
        RECT 77.550 381.300 79.650 383.400 ;
        RECT 62.250 379.500 64.350 380.400 ;
        RECT 74.850 379.800 76.650 380.400 ;
        RECT 62.250 378.300 70.050 379.500 ;
        RECT 68.250 377.700 70.050 378.300 ;
        RECT 70.950 378.900 76.650 379.800 ;
        RECT 53.550 376.500 54.450 377.400 ;
        RECT 70.950 376.800 71.850 378.900 ;
        RECT 74.850 378.600 76.650 378.900 ;
        RECT 77.550 378.600 80.550 380.400 ;
        RECT 77.550 377.700 78.750 378.600 ;
        RECT 63.450 376.500 71.850 376.800 ;
        RECT 53.550 375.900 71.850 376.500 ;
        RECT 73.950 376.800 78.750 377.700 ;
        RECT 82.650 377.400 84.450 390.000 ;
        RECT 85.650 377.400 87.450 389.400 ;
        RECT 98.100 383.400 99.900 390.000 ;
        RECT 101.100 383.400 102.900 389.400 ;
        RECT 53.550 375.300 65.250 375.900 ;
        RECT 53.550 360.600 54.450 375.300 ;
        RECT 63.450 375.000 65.250 375.300 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 65.100 368.400 67.200 370.050 ;
        RECT 55.950 365.400 57.750 367.950 ;
        RECT 59.100 367.200 67.200 368.400 ;
        RECT 59.100 366.600 60.900 367.200 ;
        RECT 62.100 365.400 63.900 366.000 ;
        RECT 55.950 364.200 63.900 365.400 ;
        RECT 73.950 364.200 74.850 376.800 ;
        RECT 77.550 374.100 79.650 374.700 ;
        RECT 83.550 374.100 85.350 374.550 ;
        RECT 77.550 372.900 85.350 374.100 ;
        RECT 77.550 372.600 79.650 372.900 ;
        RECT 83.550 372.750 85.350 372.900 ;
        RECT 86.250 370.050 87.450 377.400 ;
        RECT 98.100 370.050 99.900 371.850 ;
        RECT 101.100 370.050 102.300 383.400 ;
        RECT 113.400 377.400 115.200 390.000 ;
        RECT 118.500 378.900 120.300 389.400 ;
        RECT 121.500 383.400 123.300 390.000 ;
        RECT 121.200 380.100 123.000 381.900 ;
        RECT 126.150 379.200 127.950 389.400 ;
        RECT 118.500 377.400 120.900 378.900 ;
        RECT 113.100 370.050 114.900 371.850 ;
        RECT 119.700 370.050 120.900 377.400 ;
        RECT 125.550 377.400 127.950 379.200 ;
        RECT 129.150 377.400 130.950 390.000 ;
        RECT 134.550 380.400 136.350 389.400 ;
        RECT 139.350 383.400 141.150 390.000 ;
        RECT 142.350 382.500 144.150 389.400 ;
        RECT 145.350 383.400 147.150 390.000 ;
        RECT 149.850 383.400 151.650 389.400 ;
        RECT 138.450 381.450 145.050 382.500 ;
        RECT 138.450 380.700 140.250 381.450 ;
        RECT 143.250 380.700 145.050 381.450 ;
        RECT 149.550 381.300 151.650 383.400 ;
        RECT 134.250 379.500 136.350 380.400 ;
        RECT 146.850 379.800 148.650 380.400 ;
        RECT 134.250 378.300 142.050 379.500 ;
        RECT 140.250 377.700 142.050 378.300 ;
        RECT 142.950 378.900 148.650 379.800 ;
        RECT 125.550 376.500 126.450 377.400 ;
        RECT 142.950 376.800 143.850 378.900 ;
        RECT 146.850 378.600 148.650 378.900 ;
        RECT 149.550 378.600 152.550 380.400 ;
        RECT 149.550 377.700 150.750 378.600 ;
        RECT 135.450 376.500 143.850 376.800 ;
        RECT 125.550 375.900 143.850 376.500 ;
        RECT 145.950 376.800 150.750 377.700 ;
        RECT 154.650 377.400 156.450 390.000 ;
        RECT 157.650 377.400 159.450 389.400 ;
        RECT 170.100 383.400 171.900 390.000 ;
        RECT 173.100 383.400 174.900 389.400 ;
        RECT 125.550 375.300 137.250 375.900 ;
        RECT 82.950 369.750 87.450 370.050 ;
        RECT 81.150 367.950 87.450 369.750 ;
        RECT 97.950 367.950 100.050 370.050 ;
        RECT 100.950 367.950 103.050 370.050 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 62.850 363.000 74.850 364.200 ;
        RECT 62.850 361.200 63.900 363.000 ;
        RECT 73.050 362.400 74.850 363.000 ;
        RECT 53.550 358.800 55.950 360.600 ;
        RECT 49.050 354.600 50.850 358.800 ;
        RECT 54.150 354.600 55.950 358.800 ;
        RECT 57.150 354.000 58.950 360.600 ;
        RECT 59.850 358.200 61.950 359.700 ;
        RECT 62.850 359.400 64.650 361.200 ;
        RECT 86.250 360.600 87.450 367.950 ;
        RECT 65.850 359.550 67.650 360.300 ;
        RECT 65.850 358.500 70.800 359.550 ;
        RECT 59.850 357.600 63.750 358.200 ;
        RECT 69.750 357.600 70.800 358.500 ;
        RECT 77.250 357.600 79.650 359.700 ;
        RECT 60.150 356.700 63.750 357.600 ;
        RECT 61.950 354.600 63.750 356.700 ;
        RECT 66.450 354.000 68.250 357.600 ;
        RECT 69.750 354.600 71.550 357.600 ;
        RECT 72.750 354.000 74.550 357.600 ;
        RECT 77.250 354.600 79.050 357.600 ;
        RECT 82.350 354.000 84.150 360.600 ;
        RECT 85.650 354.600 87.450 360.600 ;
        RECT 101.100 357.600 102.300 367.950 ;
        RECT 116.100 366.150 117.900 367.950 ;
        RECT 119.700 363.600 120.900 367.950 ;
        RECT 122.100 366.150 123.900 367.950 ;
        RECT 119.700 362.700 123.300 363.600 ;
        RECT 113.100 359.700 120.900 361.050 ;
        RECT 98.100 354.000 99.900 357.600 ;
        RECT 101.100 354.600 102.900 357.600 ;
        RECT 113.100 354.600 114.900 359.700 ;
        RECT 116.100 354.000 117.900 358.800 ;
        RECT 119.100 354.600 120.900 359.700 ;
        RECT 122.100 360.600 123.300 362.700 ;
        RECT 125.550 360.600 126.450 375.300 ;
        RECT 135.450 375.000 137.250 375.300 ;
        RECT 127.950 367.950 130.050 370.050 ;
        RECT 137.100 368.400 139.200 370.050 ;
        RECT 127.950 365.400 129.750 367.950 ;
        RECT 131.100 367.200 139.200 368.400 ;
        RECT 131.100 366.600 132.900 367.200 ;
        RECT 134.100 365.400 135.900 366.000 ;
        RECT 127.950 364.200 135.900 365.400 ;
        RECT 145.950 364.200 146.850 376.800 ;
        RECT 149.550 374.100 151.650 374.700 ;
        RECT 155.550 374.100 157.350 374.550 ;
        RECT 149.550 372.900 157.350 374.100 ;
        RECT 149.550 372.600 151.650 372.900 ;
        RECT 155.550 372.750 157.350 372.900 ;
        RECT 158.250 370.050 159.450 377.400 ;
        RECT 170.100 370.050 171.900 371.850 ;
        RECT 173.100 370.050 174.300 383.400 ;
        RECT 185.100 377.400 186.900 390.000 ;
        RECT 189.600 377.400 192.900 389.400 ;
        RECT 195.600 377.400 197.400 390.000 ;
        RECT 209.100 383.400 210.900 390.000 ;
        RECT 212.100 383.400 213.900 389.400 ;
        RECT 215.100 383.400 216.900 390.000 ;
        RECT 185.100 370.050 186.900 371.850 ;
        RECT 190.950 370.050 192.000 377.400 ;
        RECT 196.950 370.050 198.750 371.850 ;
        RECT 212.100 370.050 213.300 383.400 ;
        RECT 227.100 378.300 228.900 389.400 ;
        RECT 230.100 379.500 231.900 390.000 ;
        RECT 234.600 378.300 236.400 389.400 ;
        RECT 238.800 379.500 240.900 390.000 ;
        RECT 242.100 378.600 243.900 389.400 ;
        RECT 254.100 383.400 255.900 390.000 ;
        RECT 257.100 383.400 258.900 389.400 ;
        RECT 227.100 377.100 231.900 378.300 ;
        RECT 234.600 377.400 237.900 378.300 ;
        RECT 229.800 376.200 231.900 377.100 ;
        RECT 229.800 375.300 235.200 376.200 ;
        RECT 233.400 373.500 235.200 375.300 ;
        RECT 236.700 373.050 237.900 377.400 ;
        RECT 238.800 377.400 243.900 378.600 ;
        RECT 238.800 376.500 240.900 377.400 ;
        RECT 236.100 372.300 238.200 373.050 ;
        RECT 231.900 370.200 233.700 372.000 ;
        RECT 235.200 370.950 238.200 372.300 ;
        RECT 154.950 369.750 159.450 370.050 ;
        RECT 153.150 367.950 159.450 369.750 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 184.950 367.950 187.050 370.050 ;
        RECT 187.950 367.950 190.050 370.050 ;
        RECT 134.850 363.000 146.850 364.200 ;
        RECT 134.850 361.200 135.900 363.000 ;
        RECT 145.050 362.400 146.850 363.000 ;
        RECT 122.100 354.600 123.900 360.600 ;
        RECT 125.550 358.800 127.950 360.600 ;
        RECT 126.150 354.600 127.950 358.800 ;
        RECT 129.150 354.000 130.950 360.600 ;
        RECT 131.850 358.200 133.950 359.700 ;
        RECT 134.850 359.400 136.650 361.200 ;
        RECT 158.250 360.600 159.450 367.950 ;
        RECT 137.850 359.550 139.650 360.300 ;
        RECT 137.850 358.500 142.800 359.550 ;
        RECT 131.850 357.600 135.750 358.200 ;
        RECT 141.750 357.600 142.800 358.500 ;
        RECT 149.250 357.600 151.650 359.700 ;
        RECT 132.150 356.700 135.750 357.600 ;
        RECT 133.950 354.600 135.750 356.700 ;
        RECT 138.450 354.000 140.250 357.600 ;
        RECT 141.750 354.600 143.550 357.600 ;
        RECT 144.750 354.000 146.550 357.600 ;
        RECT 149.250 354.600 151.050 357.600 ;
        RECT 154.350 354.000 156.150 360.600 ;
        RECT 157.650 354.600 159.450 360.600 ;
        RECT 173.100 357.600 174.300 367.950 ;
        RECT 188.250 366.150 190.050 367.950 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 208.950 367.950 211.050 370.050 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 190.950 363.300 192.000 367.950 ;
        RECT 193.950 366.150 195.750 367.950 ;
        RECT 209.250 366.150 211.050 367.950 ;
        RECT 190.950 362.100 195.300 363.300 ;
        RECT 185.100 360.000 192.900 360.900 ;
        RECT 194.400 360.600 195.300 362.100 ;
        RECT 212.100 362.700 213.300 367.950 ;
        RECT 215.100 366.150 216.900 367.950 ;
        RECT 227.100 367.800 229.200 370.050 ;
        RECT 231.900 368.100 234.000 370.200 ;
        RECT 227.400 367.200 229.200 367.800 ;
        RECT 227.400 366.000 234.000 367.200 ;
        RECT 231.900 365.100 234.000 366.000 ;
        RECT 229.500 363.000 231.600 363.600 ;
        RECT 232.500 363.300 234.300 365.100 ;
        RECT 235.200 364.200 236.100 370.950 ;
        RECT 241.800 370.050 243.600 371.850 ;
        RECT 237.000 368.100 238.800 369.900 ;
        RECT 237.000 366.000 239.100 368.100 ;
        RECT 241.800 367.950 243.900 370.050 ;
        RECT 254.100 367.950 256.200 370.050 ;
        RECT 254.250 366.150 256.050 367.950 ;
        RECT 212.100 361.800 216.300 362.700 ;
        RECT 170.100 354.000 171.900 357.600 ;
        RECT 173.100 354.600 174.900 357.600 ;
        RECT 185.100 354.600 186.900 360.000 ;
        RECT 188.100 354.000 189.900 359.100 ;
        RECT 191.100 355.500 192.900 360.000 ;
        RECT 194.100 356.400 195.900 360.600 ;
        RECT 197.100 355.500 198.900 360.600 ;
        RECT 191.100 354.600 198.900 355.500 ;
        RECT 209.400 354.000 211.200 360.600 ;
        RECT 214.500 354.600 216.300 361.800 ;
        RECT 227.100 361.500 231.600 363.000 ;
        RECT 235.200 362.100 238.200 364.200 ;
        RECT 227.100 360.600 228.600 361.500 ;
        RECT 227.100 354.600 228.900 360.600 ;
        RECT 235.200 360.000 236.100 362.100 ;
        RECT 239.400 361.500 241.500 363.900 ;
        RECT 257.100 363.300 258.000 383.400 ;
        RECT 260.100 378.000 261.900 390.000 ;
        RECT 263.100 377.400 264.900 389.400 ;
        RECT 267.150 379.200 268.950 389.400 ;
        RECT 266.550 377.400 268.950 379.200 ;
        RECT 270.150 377.400 271.950 390.000 ;
        RECT 275.550 380.400 277.350 389.400 ;
        RECT 280.350 383.400 282.150 390.000 ;
        RECT 283.350 382.500 285.150 389.400 ;
        RECT 286.350 383.400 288.150 390.000 ;
        RECT 290.850 383.400 292.650 389.400 ;
        RECT 279.450 381.450 286.050 382.500 ;
        RECT 279.450 380.700 281.250 381.450 ;
        RECT 284.250 380.700 286.050 381.450 ;
        RECT 290.550 381.300 292.650 383.400 ;
        RECT 275.250 379.500 277.350 380.400 ;
        RECT 287.850 379.800 289.650 380.400 ;
        RECT 275.250 378.300 283.050 379.500 ;
        RECT 281.250 377.700 283.050 378.300 ;
        RECT 283.950 378.900 289.650 379.800 ;
        RECT 259.200 370.050 261.000 371.850 ;
        RECT 263.400 370.050 264.300 377.400 ;
        RECT 266.550 376.500 267.450 377.400 ;
        RECT 283.950 376.800 284.850 378.900 ;
        RECT 287.850 378.600 289.650 378.900 ;
        RECT 290.550 378.600 293.550 380.400 ;
        RECT 290.550 377.700 291.750 378.600 ;
        RECT 276.450 376.500 284.850 376.800 ;
        RECT 266.550 375.900 284.850 376.500 ;
        RECT 286.950 376.800 291.750 377.700 ;
        RECT 295.650 377.400 297.450 390.000 ;
        RECT 298.650 377.400 300.450 389.400 ;
        RECT 311.100 383.400 312.900 389.400 ;
        RECT 314.100 384.000 315.900 390.000 ;
        RECT 266.550 375.300 278.250 375.900 ;
        RECT 259.500 367.950 261.600 370.050 ;
        RECT 262.800 367.950 264.900 370.050 ;
        RECT 254.100 362.400 262.500 363.300 ;
        RECT 239.400 360.600 243.900 361.500 ;
        RECT 230.100 354.000 231.900 359.700 ;
        RECT 234.300 354.600 236.100 360.000 ;
        RECT 238.800 354.000 240.600 359.700 ;
        RECT 242.100 354.600 243.900 360.600 ;
        RECT 254.100 354.600 255.900 362.400 ;
        RECT 260.700 361.500 262.500 362.400 ;
        RECT 263.400 360.600 264.300 367.950 ;
        RECT 258.600 354.000 260.400 360.600 ;
        RECT 261.600 358.800 264.300 360.600 ;
        RECT 266.550 360.600 267.450 375.300 ;
        RECT 276.450 375.000 278.250 375.300 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 278.100 368.400 280.200 370.050 ;
        RECT 268.950 365.400 270.750 367.950 ;
        RECT 272.100 367.200 280.200 368.400 ;
        RECT 272.100 366.600 273.900 367.200 ;
        RECT 275.100 365.400 276.900 366.000 ;
        RECT 268.950 364.200 276.900 365.400 ;
        RECT 286.950 364.200 287.850 376.800 ;
        RECT 290.550 374.100 292.650 374.700 ;
        RECT 296.550 374.100 298.350 374.550 ;
        RECT 290.550 372.900 298.350 374.100 ;
        RECT 290.550 372.600 292.650 372.900 ;
        RECT 296.550 372.750 298.350 372.900 ;
        RECT 299.250 370.050 300.450 377.400 ;
        RECT 312.000 383.100 312.900 383.400 ;
        RECT 317.100 383.400 318.900 389.400 ;
        RECT 320.100 383.400 321.900 390.000 ;
        RECT 332.100 383.400 333.900 390.000 ;
        RECT 335.100 383.400 336.900 389.400 ;
        RECT 317.100 383.100 318.600 383.400 ;
        RECT 312.000 382.200 318.600 383.100 ;
        RECT 312.000 370.050 312.900 382.200 ;
        RECT 317.100 370.050 318.900 371.850 ;
        RECT 332.100 370.050 333.900 371.850 ;
        RECT 335.100 370.050 336.300 383.400 ;
        RECT 338.550 377.400 340.350 389.400 ;
        RECT 341.550 377.400 343.350 390.000 ;
        RECT 346.350 383.400 348.150 389.400 ;
        RECT 350.850 383.400 352.650 390.000 ;
        RECT 346.350 381.300 348.450 383.400 ;
        RECT 353.850 382.500 355.650 389.400 ;
        RECT 356.850 383.400 358.650 390.000 ;
        RECT 352.950 381.450 359.550 382.500 ;
        RECT 352.950 380.700 354.750 381.450 ;
        RECT 357.750 380.700 359.550 381.450 ;
        RECT 361.650 380.400 363.450 389.400 ;
        RECT 345.450 378.600 348.450 380.400 ;
        RECT 349.350 379.800 351.150 380.400 ;
        RECT 349.350 378.900 355.050 379.800 ;
        RECT 361.650 379.500 363.750 380.400 ;
        RECT 349.350 378.600 351.150 378.900 ;
        RECT 347.250 377.700 348.450 378.600 ;
        RECT 338.550 370.050 339.750 377.400 ;
        RECT 347.250 376.800 352.050 377.700 ;
        RECT 340.650 374.100 342.450 374.550 ;
        RECT 346.350 374.100 348.450 374.700 ;
        RECT 340.650 372.900 348.450 374.100 ;
        RECT 340.650 372.750 342.450 372.900 ;
        RECT 346.350 372.600 348.450 372.900 ;
        RECT 295.950 369.750 300.450 370.050 ;
        RECT 294.150 367.950 300.450 369.750 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 338.550 369.750 343.050 370.050 ;
        RECT 338.550 367.950 344.850 369.750 ;
        RECT 275.850 363.000 287.850 364.200 ;
        RECT 275.850 361.200 276.900 363.000 ;
        RECT 286.050 362.400 287.850 363.000 ;
        RECT 266.550 358.800 268.950 360.600 ;
        RECT 261.600 354.600 263.400 358.800 ;
        RECT 267.150 354.600 268.950 358.800 ;
        RECT 270.150 354.000 271.950 360.600 ;
        RECT 272.850 358.200 274.950 359.700 ;
        RECT 275.850 359.400 277.650 361.200 ;
        RECT 299.250 360.600 300.450 367.950 ;
        RECT 312.000 364.200 312.900 367.950 ;
        RECT 314.100 366.150 315.900 367.950 ;
        RECT 320.100 366.150 321.900 367.950 ;
        RECT 312.000 363.000 315.300 364.200 ;
        RECT 278.850 359.550 280.650 360.300 ;
        RECT 278.850 358.500 283.800 359.550 ;
        RECT 272.850 357.600 276.750 358.200 ;
        RECT 282.750 357.600 283.800 358.500 ;
        RECT 290.250 357.600 292.650 359.700 ;
        RECT 273.150 356.700 276.750 357.600 ;
        RECT 274.950 354.600 276.750 356.700 ;
        RECT 279.450 354.000 281.250 357.600 ;
        RECT 282.750 354.600 284.550 357.600 ;
        RECT 285.750 354.000 287.550 357.600 ;
        RECT 290.250 354.600 292.050 357.600 ;
        RECT 295.350 354.000 297.150 360.600 ;
        RECT 298.650 354.600 300.450 360.600 ;
        RECT 313.500 354.600 315.300 363.000 ;
        RECT 320.100 354.000 321.900 363.600 ;
        RECT 335.100 357.600 336.300 367.950 ;
        RECT 338.550 360.600 339.750 367.950 ;
        RECT 351.150 364.200 352.050 376.800 ;
        RECT 354.150 376.800 355.050 378.900 ;
        RECT 355.950 378.300 363.750 379.500 ;
        RECT 355.950 377.700 357.750 378.300 ;
        RECT 367.050 377.400 368.850 390.000 ;
        RECT 370.050 379.200 371.850 389.400 ;
        RECT 383.700 383.400 385.500 390.000 ;
        RECT 384.000 380.100 385.800 381.900 ;
        RECT 370.050 377.400 372.450 379.200 ;
        RECT 386.700 378.900 388.500 389.400 ;
        RECT 354.150 376.500 362.550 376.800 ;
        RECT 371.550 376.500 372.450 377.400 ;
        RECT 354.150 375.900 372.450 376.500 ;
        RECT 360.750 375.300 372.450 375.900 ;
        RECT 360.750 375.000 362.550 375.300 ;
        RECT 358.800 368.400 360.900 370.050 ;
        RECT 358.800 367.200 366.900 368.400 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 365.100 366.600 366.900 367.200 ;
        RECT 362.100 365.400 363.900 366.000 ;
        RECT 368.250 365.400 370.050 367.950 ;
        RECT 362.100 364.200 370.050 365.400 ;
        RECT 351.150 363.000 363.150 364.200 ;
        RECT 351.150 362.400 352.950 363.000 ;
        RECT 362.100 361.200 363.150 363.000 ;
        RECT 332.100 354.000 333.900 357.600 ;
        RECT 335.100 354.600 336.900 357.600 ;
        RECT 338.550 354.600 340.350 360.600 ;
        RECT 341.850 354.000 343.650 360.600 ;
        RECT 346.350 357.600 348.750 359.700 ;
        RECT 358.350 359.550 360.150 360.300 ;
        RECT 355.200 358.500 360.150 359.550 ;
        RECT 361.350 359.400 363.150 361.200 ;
        RECT 371.550 360.600 372.450 375.300 ;
        RECT 386.100 377.400 388.500 378.900 ;
        RECT 391.800 377.400 393.600 390.000 ;
        RECT 404.100 383.400 405.900 390.000 ;
        RECT 407.100 383.400 408.900 389.400 ;
        RECT 410.100 383.400 411.900 390.000 ;
        RECT 422.100 383.400 423.900 390.000 ;
        RECT 425.100 383.400 426.900 389.400 ;
        RECT 428.100 383.400 429.900 390.000 ;
        RECT 440.700 383.400 442.500 390.000 ;
        RECT 386.100 370.050 387.300 377.400 ;
        RECT 392.100 370.050 393.900 371.850 ;
        RECT 407.100 370.050 408.300 383.400 ;
        RECT 425.100 370.050 426.300 383.400 ;
        RECT 441.000 380.100 442.800 381.900 ;
        RECT 427.950 378.450 430.050 379.050 ;
        RECT 436.950 378.450 439.050 379.050 ;
        RECT 443.700 378.900 445.500 389.400 ;
        RECT 427.950 377.550 439.050 378.450 ;
        RECT 427.950 376.950 430.050 377.550 ;
        RECT 436.950 376.950 439.050 377.550 ;
        RECT 443.100 377.400 445.500 378.900 ;
        RECT 448.800 377.400 450.600 390.000 ;
        RECT 453.150 379.200 454.950 389.400 ;
        RECT 452.550 377.400 454.950 379.200 ;
        RECT 456.150 377.400 457.950 390.000 ;
        RECT 461.550 380.400 463.350 389.400 ;
        RECT 466.350 383.400 468.150 390.000 ;
        RECT 469.350 382.500 471.150 389.400 ;
        RECT 472.350 383.400 474.150 390.000 ;
        RECT 476.850 383.400 478.650 389.400 ;
        RECT 465.450 381.450 472.050 382.500 ;
        RECT 465.450 380.700 467.250 381.450 ;
        RECT 470.250 380.700 472.050 381.450 ;
        RECT 476.550 381.300 478.650 383.400 ;
        RECT 461.250 379.500 463.350 380.400 ;
        RECT 473.850 379.800 475.650 380.400 ;
        RECT 461.250 378.300 469.050 379.500 ;
        RECT 467.250 377.700 469.050 378.300 ;
        RECT 469.950 378.900 475.650 379.800 ;
        RECT 443.100 370.050 444.300 377.400 ;
        RECT 452.550 376.500 453.450 377.400 ;
        RECT 469.950 376.800 470.850 378.900 ;
        RECT 473.850 378.600 475.650 378.900 ;
        RECT 476.550 378.600 479.550 380.400 ;
        RECT 476.550 377.700 477.750 378.600 ;
        RECT 462.450 376.500 470.850 376.800 ;
        RECT 452.550 375.900 470.850 376.500 ;
        RECT 472.950 376.800 477.750 377.700 ;
        RECT 481.650 377.400 483.450 390.000 ;
        RECT 484.650 377.400 486.450 389.400 ;
        RECT 497.100 383.400 498.900 390.000 ;
        RECT 500.100 383.400 501.900 389.400 ;
        RECT 503.100 383.400 504.900 390.000 ;
        RECT 515.700 383.400 517.500 390.000 ;
        RECT 452.550 375.300 464.250 375.900 ;
        RECT 449.100 370.050 450.900 371.850 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 406.950 367.950 409.050 370.050 ;
        RECT 409.950 367.950 412.050 370.050 ;
        RECT 421.950 367.950 424.050 370.050 ;
        RECT 424.950 367.950 427.050 370.050 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 442.950 367.950 445.050 370.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 383.100 366.150 384.900 367.950 ;
        RECT 386.100 363.600 387.300 367.950 ;
        RECT 389.100 366.150 390.900 367.950 ;
        RECT 404.250 366.150 406.050 367.950 ;
        RECT 383.700 362.700 387.300 363.600 ;
        RECT 407.100 362.700 408.300 367.950 ;
        RECT 410.100 366.150 411.900 367.950 ;
        RECT 422.250 366.150 424.050 367.950 ;
        RECT 425.100 362.700 426.300 367.950 ;
        RECT 428.100 366.150 429.900 367.950 ;
        RECT 440.100 366.150 441.900 367.950 ;
        RECT 443.100 363.600 444.300 367.950 ;
        RECT 446.100 366.150 447.900 367.950 ;
        RECT 440.700 362.700 444.300 363.600 ;
        RECT 383.700 360.600 384.900 362.700 ;
        RECT 407.100 361.800 411.300 362.700 ;
        RECT 425.100 361.800 429.300 362.700 ;
        RECT 355.200 357.600 356.250 358.500 ;
        RECT 364.050 358.200 366.150 359.700 ;
        RECT 362.250 357.600 366.150 358.200 ;
        RECT 346.950 354.600 348.750 357.600 ;
        RECT 351.450 354.000 353.250 357.600 ;
        RECT 354.450 354.600 356.250 357.600 ;
        RECT 357.750 354.000 359.550 357.600 ;
        RECT 362.250 356.700 365.850 357.600 ;
        RECT 362.250 354.600 364.050 356.700 ;
        RECT 367.050 354.000 368.850 360.600 ;
        RECT 370.050 358.800 372.450 360.600 ;
        RECT 370.050 354.600 371.850 358.800 ;
        RECT 383.100 354.600 384.900 360.600 ;
        RECT 386.100 359.700 393.900 361.050 ;
        RECT 386.100 354.600 387.900 359.700 ;
        RECT 389.100 354.000 390.900 358.800 ;
        RECT 392.100 354.600 393.900 359.700 ;
        RECT 404.400 354.000 406.200 360.600 ;
        RECT 409.500 354.600 411.300 361.800 ;
        RECT 422.400 354.000 424.200 360.600 ;
        RECT 427.500 354.600 429.300 361.800 ;
        RECT 440.700 360.600 441.900 362.700 ;
        RECT 440.100 354.600 441.900 360.600 ;
        RECT 443.100 359.700 450.900 361.050 ;
        RECT 443.100 354.600 444.900 359.700 ;
        RECT 446.100 354.000 447.900 358.800 ;
        RECT 449.100 354.600 450.900 359.700 ;
        RECT 452.550 360.600 453.450 375.300 ;
        RECT 462.450 375.000 464.250 375.300 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 464.100 368.400 466.200 370.050 ;
        RECT 454.950 365.400 456.750 367.950 ;
        RECT 458.100 367.200 466.200 368.400 ;
        RECT 458.100 366.600 459.900 367.200 ;
        RECT 461.100 365.400 462.900 366.000 ;
        RECT 454.950 364.200 462.900 365.400 ;
        RECT 472.950 364.200 473.850 376.800 ;
        RECT 476.550 374.100 478.650 374.700 ;
        RECT 482.550 374.100 484.350 374.550 ;
        RECT 476.550 372.900 484.350 374.100 ;
        RECT 476.550 372.600 478.650 372.900 ;
        RECT 482.550 372.750 484.350 372.900 ;
        RECT 485.250 370.050 486.450 377.400 ;
        RECT 500.100 370.050 501.300 383.400 ;
        RECT 516.000 380.100 517.800 381.900 ;
        RECT 518.700 378.900 520.500 389.400 ;
        RECT 518.100 377.400 520.500 378.900 ;
        RECT 523.800 377.400 525.600 390.000 ;
        RECT 539.100 383.400 540.900 390.000 ;
        RECT 542.100 383.400 543.900 389.400 ;
        RECT 545.100 383.400 546.900 390.000 ;
        RECT 557.100 383.400 558.900 390.000 ;
        RECT 560.100 383.400 561.900 389.400 ;
        RECT 563.100 383.400 564.900 390.000 ;
        RECT 578.700 383.400 580.500 390.000 ;
        RECT 518.100 370.050 519.300 377.400 ;
        RECT 534.000 372.450 538.050 373.050 ;
        RECT 524.100 370.050 525.900 371.850 ;
        RECT 533.550 370.950 538.050 372.450 ;
        RECT 481.950 369.750 486.450 370.050 ;
        RECT 480.150 367.950 486.450 369.750 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 514.950 367.950 517.050 370.050 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 461.850 363.000 473.850 364.200 ;
        RECT 461.850 361.200 462.900 363.000 ;
        RECT 472.050 362.400 473.850 363.000 ;
        RECT 452.550 358.800 454.950 360.600 ;
        RECT 453.150 354.600 454.950 358.800 ;
        RECT 456.150 354.000 457.950 360.600 ;
        RECT 458.850 358.200 460.950 359.700 ;
        RECT 461.850 359.400 463.650 361.200 ;
        RECT 485.250 360.600 486.450 367.950 ;
        RECT 497.250 366.150 499.050 367.950 ;
        RECT 500.100 362.700 501.300 367.950 ;
        RECT 503.100 366.150 504.900 367.950 ;
        RECT 515.100 366.150 516.900 367.950 ;
        RECT 518.100 363.600 519.300 367.950 ;
        RECT 521.100 366.150 522.900 367.950 ;
        RECT 526.950 366.450 529.050 367.050 ;
        RECT 533.550 366.450 534.450 370.950 ;
        RECT 542.100 370.050 543.300 383.400 ;
        RECT 560.100 370.050 561.300 383.400 ;
        RECT 579.000 380.100 580.800 381.900 ;
        RECT 581.700 378.900 583.500 389.400 ;
        RECT 581.100 377.400 583.500 378.900 ;
        RECT 586.800 377.400 588.600 390.000 ;
        RECT 591.150 379.200 592.950 389.400 ;
        RECT 590.550 377.400 592.950 379.200 ;
        RECT 594.150 377.400 595.950 390.000 ;
        RECT 599.550 380.400 601.350 389.400 ;
        RECT 604.350 383.400 606.150 390.000 ;
        RECT 607.350 382.500 609.150 389.400 ;
        RECT 610.350 383.400 612.150 390.000 ;
        RECT 614.850 383.400 616.650 389.400 ;
        RECT 603.450 381.450 610.050 382.500 ;
        RECT 603.450 380.700 605.250 381.450 ;
        RECT 608.250 380.700 610.050 381.450 ;
        RECT 614.550 381.300 616.650 383.400 ;
        RECT 599.250 379.500 601.350 380.400 ;
        RECT 611.850 379.800 613.650 380.400 ;
        RECT 599.250 378.300 607.050 379.500 ;
        RECT 605.250 377.700 607.050 378.300 ;
        RECT 607.950 378.900 613.650 379.800 ;
        RECT 581.100 370.050 582.300 377.400 ;
        RECT 590.550 376.500 591.450 377.400 ;
        RECT 607.950 376.800 608.850 378.900 ;
        RECT 611.850 378.600 613.650 378.900 ;
        RECT 614.550 378.600 617.550 380.400 ;
        RECT 614.550 377.700 615.750 378.600 ;
        RECT 600.450 376.500 608.850 376.800 ;
        RECT 590.550 375.900 608.850 376.500 ;
        RECT 610.950 376.800 615.750 377.700 ;
        RECT 619.650 377.400 621.450 390.000 ;
        RECT 622.650 377.400 624.450 389.400 ;
        RECT 635.400 377.400 637.200 390.000 ;
        RECT 640.500 378.900 642.300 389.400 ;
        RECT 643.500 383.400 645.300 390.000 ;
        RECT 643.200 380.100 645.000 381.900 ;
        RECT 640.500 377.400 642.900 378.900 ;
        RECT 656.400 377.400 658.200 390.000 ;
        RECT 661.500 378.900 663.300 389.400 ;
        RECT 664.500 383.400 666.300 390.000 ;
        RECT 664.200 380.100 666.000 381.900 ;
        RECT 661.500 377.400 663.900 378.900 ;
        RECT 677.100 377.400 678.900 390.000 ;
        RECT 682.200 378.600 684.000 389.400 ;
        RECT 680.400 377.400 684.000 378.600 ;
        RECT 696.000 378.600 697.800 389.400 ;
        RECT 696.000 377.400 699.600 378.600 ;
        RECT 701.100 377.400 702.900 390.000 ;
        RECT 713.100 383.400 714.900 390.000 ;
        RECT 716.100 383.400 717.900 389.400 ;
        RECT 719.100 383.400 720.900 390.000 ;
        RECT 731.700 383.400 733.500 390.000 ;
        RECT 590.550 375.300 602.250 375.900 ;
        RECT 587.100 370.050 588.900 371.850 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 544.950 367.950 547.050 370.050 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 559.950 367.950 562.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 580.950 367.950 583.050 370.050 ;
        RECT 583.950 367.950 586.050 370.050 ;
        RECT 586.950 367.950 589.050 370.050 ;
        RECT 526.950 365.550 534.450 366.450 ;
        RECT 539.250 366.150 541.050 367.950 ;
        RECT 526.950 364.950 529.050 365.550 ;
        RECT 515.700 362.700 519.300 363.600 ;
        RECT 542.100 362.700 543.300 367.950 ;
        RECT 545.100 366.150 546.900 367.950 ;
        RECT 557.250 366.150 559.050 367.950 ;
        RECT 560.100 362.700 561.300 367.950 ;
        RECT 563.100 366.150 564.900 367.950 ;
        RECT 578.100 366.150 579.900 367.950 ;
        RECT 581.100 363.600 582.300 367.950 ;
        RECT 584.100 366.150 585.900 367.950 ;
        RECT 578.700 362.700 582.300 363.600 ;
        RECT 500.100 361.800 504.300 362.700 ;
        RECT 464.850 359.550 466.650 360.300 ;
        RECT 464.850 358.500 469.800 359.550 ;
        RECT 458.850 357.600 462.750 358.200 ;
        RECT 468.750 357.600 469.800 358.500 ;
        RECT 476.250 357.600 478.650 359.700 ;
        RECT 459.150 356.700 462.750 357.600 ;
        RECT 460.950 354.600 462.750 356.700 ;
        RECT 465.450 354.000 467.250 357.600 ;
        RECT 468.750 354.600 470.550 357.600 ;
        RECT 471.750 354.000 473.550 357.600 ;
        RECT 476.250 354.600 478.050 357.600 ;
        RECT 481.350 354.000 483.150 360.600 ;
        RECT 484.650 354.600 486.450 360.600 ;
        RECT 497.400 354.000 499.200 360.600 ;
        RECT 502.500 354.600 504.300 361.800 ;
        RECT 515.700 360.600 516.900 362.700 ;
        RECT 542.100 361.800 546.300 362.700 ;
        RECT 560.100 361.800 564.300 362.700 ;
        RECT 515.100 354.600 516.900 360.600 ;
        RECT 518.100 359.700 525.900 361.050 ;
        RECT 518.100 354.600 519.900 359.700 ;
        RECT 521.100 354.000 522.900 358.800 ;
        RECT 524.100 354.600 525.900 359.700 ;
        RECT 539.400 354.000 541.200 360.600 ;
        RECT 544.500 354.600 546.300 361.800 ;
        RECT 557.400 354.000 559.200 360.600 ;
        RECT 562.500 354.600 564.300 361.800 ;
        RECT 578.700 360.600 579.900 362.700 ;
        RECT 578.100 354.600 579.900 360.600 ;
        RECT 581.100 359.700 588.900 361.050 ;
        RECT 581.100 354.600 582.900 359.700 ;
        RECT 584.100 354.000 585.900 358.800 ;
        RECT 587.100 354.600 588.900 359.700 ;
        RECT 590.550 360.600 591.450 375.300 ;
        RECT 600.450 375.000 602.250 375.300 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 602.100 368.400 604.200 370.050 ;
        RECT 592.950 365.400 594.750 367.950 ;
        RECT 596.100 367.200 604.200 368.400 ;
        RECT 596.100 366.600 597.900 367.200 ;
        RECT 599.100 365.400 600.900 366.000 ;
        RECT 592.950 364.200 600.900 365.400 ;
        RECT 610.950 364.200 611.850 376.800 ;
        RECT 614.550 374.100 616.650 374.700 ;
        RECT 620.550 374.100 622.350 374.550 ;
        RECT 614.550 372.900 622.350 374.100 ;
        RECT 614.550 372.600 616.650 372.900 ;
        RECT 620.550 372.750 622.350 372.900 ;
        RECT 623.250 370.050 624.450 377.400 ;
        RECT 635.100 370.050 636.900 371.850 ;
        RECT 641.700 370.050 642.900 377.400 ;
        RECT 656.100 370.050 657.900 371.850 ;
        RECT 662.700 370.050 663.900 377.400 ;
        RECT 677.250 370.050 679.050 371.850 ;
        RECT 680.400 370.050 681.300 377.400 ;
        RECT 685.950 372.450 690.000 373.050 ;
        RECT 683.100 370.050 684.900 371.850 ;
        RECT 685.950 370.950 690.450 372.450 ;
        RECT 619.950 369.750 624.450 370.050 ;
        RECT 618.150 367.950 624.450 369.750 ;
        RECT 634.950 367.950 637.050 370.050 ;
        RECT 637.950 367.950 640.050 370.050 ;
        RECT 640.950 367.950 643.050 370.050 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 658.950 367.950 661.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 599.850 363.000 611.850 364.200 ;
        RECT 599.850 361.200 600.900 363.000 ;
        RECT 610.050 362.400 611.850 363.000 ;
        RECT 590.550 358.800 592.950 360.600 ;
        RECT 591.150 354.600 592.950 358.800 ;
        RECT 594.150 354.000 595.950 360.600 ;
        RECT 596.850 358.200 598.950 359.700 ;
        RECT 599.850 359.400 601.650 361.200 ;
        RECT 623.250 360.600 624.450 367.950 ;
        RECT 638.100 366.150 639.900 367.950 ;
        RECT 641.700 363.600 642.900 367.950 ;
        RECT 644.100 366.150 645.900 367.950 ;
        RECT 659.100 366.150 660.900 367.950 ;
        RECT 662.700 363.600 663.900 367.950 ;
        RECT 665.100 366.150 666.900 367.950 ;
        RECT 641.700 362.700 645.300 363.600 ;
        RECT 662.700 362.700 666.300 363.600 ;
        RECT 602.850 359.550 604.650 360.300 ;
        RECT 602.850 358.500 607.800 359.550 ;
        RECT 596.850 357.600 600.750 358.200 ;
        RECT 606.750 357.600 607.800 358.500 ;
        RECT 614.250 357.600 616.650 359.700 ;
        RECT 597.150 356.700 600.750 357.600 ;
        RECT 598.950 354.600 600.750 356.700 ;
        RECT 603.450 354.000 605.250 357.600 ;
        RECT 606.750 354.600 608.550 357.600 ;
        RECT 609.750 354.000 611.550 357.600 ;
        RECT 614.250 354.600 616.050 357.600 ;
        RECT 619.350 354.000 621.150 360.600 ;
        RECT 622.650 354.600 624.450 360.600 ;
        RECT 635.100 359.700 642.900 361.050 ;
        RECT 635.100 354.600 636.900 359.700 ;
        RECT 638.100 354.000 639.900 358.800 ;
        RECT 641.100 354.600 642.900 359.700 ;
        RECT 644.100 360.600 645.300 362.700 ;
        RECT 644.100 354.600 645.900 360.600 ;
        RECT 656.100 359.700 663.900 361.050 ;
        RECT 656.100 354.600 657.900 359.700 ;
        RECT 659.100 354.000 660.900 358.800 ;
        RECT 662.100 354.600 663.900 359.700 ;
        RECT 665.100 360.600 666.300 362.700 ;
        RECT 665.100 354.600 666.900 360.600 ;
        RECT 680.400 357.600 681.300 367.950 ;
        RECT 689.550 367.050 690.450 370.950 ;
        RECT 695.100 370.050 696.900 371.850 ;
        RECT 698.700 370.050 699.600 377.400 ;
        RECT 708.000 372.450 712.050 373.050 ;
        RECT 700.950 370.050 702.750 371.850 ;
        RECT 707.550 370.950 712.050 372.450 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 697.950 367.950 700.050 370.050 ;
        RECT 700.950 367.950 703.050 370.050 ;
        RECT 685.950 365.550 690.450 367.050 ;
        RECT 685.950 364.950 690.000 365.550 ;
        RECT 698.700 357.600 699.600 367.950 ;
        RECT 707.550 367.050 708.450 370.950 ;
        RECT 716.100 370.050 717.300 383.400 ;
        RECT 732.000 380.100 733.800 381.900 ;
        RECT 734.700 378.900 736.500 389.400 ;
        RECT 734.100 377.400 736.500 378.900 ;
        RECT 739.800 377.400 741.600 390.000 ;
        RECT 755.100 377.400 756.900 390.000 ;
        RECT 759.600 377.400 762.900 389.400 ;
        RECT 765.600 377.400 767.400 390.000 ;
        RECT 779.100 383.400 780.900 390.000 ;
        RECT 782.100 383.400 783.900 389.400 ;
        RECT 721.950 372.450 726.000 373.050 ;
        RECT 721.950 370.950 726.450 372.450 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 715.950 367.950 718.050 370.050 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 703.950 365.550 708.450 367.050 ;
        RECT 713.250 366.150 715.050 367.950 ;
        RECT 703.950 364.950 708.000 365.550 ;
        RECT 716.100 362.700 717.300 367.950 ;
        RECT 719.100 366.150 720.900 367.950 ;
        RECT 725.550 367.050 726.450 370.950 ;
        RECT 734.100 370.050 735.300 377.400 ;
        RECT 742.950 372.450 747.000 373.050 ;
        RECT 740.100 370.050 741.900 371.850 ;
        RECT 742.950 370.950 747.450 372.450 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 739.950 367.950 742.050 370.050 ;
        RECT 725.550 365.550 730.050 367.050 ;
        RECT 731.100 366.150 732.900 367.950 ;
        RECT 726.000 364.950 730.050 365.550 ;
        RECT 734.100 363.600 735.300 367.950 ;
        RECT 737.100 366.150 738.900 367.950 ;
        RECT 746.550 366.450 747.450 370.950 ;
        RECT 755.100 370.050 756.900 371.850 ;
        RECT 760.950 370.050 762.000 377.400 ;
        RECT 763.950 375.450 766.050 376.050 ;
        RECT 763.950 374.550 771.450 375.450 ;
        RECT 763.950 373.950 766.050 374.550 ;
        RECT 770.550 372.450 771.450 374.550 ;
        RECT 766.950 370.050 768.750 371.850 ;
        RECT 770.550 371.550 774.450 372.450 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 751.950 366.450 754.050 367.050 ;
        RECT 746.550 365.550 754.050 366.450 ;
        RECT 758.250 366.150 760.050 367.950 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 751.950 364.950 754.050 365.550 ;
        RECT 731.700 362.700 735.300 363.600 ;
        RECT 760.950 363.300 762.000 367.950 ;
        RECT 763.950 366.150 765.750 367.950 ;
        RECT 773.550 367.050 774.450 371.550 ;
        RECT 779.100 370.050 780.900 371.850 ;
        RECT 782.100 370.050 783.300 383.400 ;
        RECT 797.100 378.300 798.900 389.400 ;
        RECT 800.100 379.500 801.900 390.000 ;
        RECT 797.100 377.400 801.600 378.300 ;
        RECT 804.600 377.400 806.400 389.400 ;
        RECT 809.100 379.500 810.900 390.000 ;
        RECT 812.100 378.600 813.900 389.400 ;
        RECT 824.100 383.400 825.900 390.000 ;
        RECT 827.100 383.400 828.900 389.400 ;
        RECT 839.700 383.400 841.500 390.000 ;
        RECT 799.500 375.300 801.600 377.400 ;
        RECT 805.200 376.050 806.400 377.400 ;
        RECT 809.100 377.400 813.900 378.600 ;
        RECT 809.100 376.500 811.200 377.400 ;
        RECT 805.200 375.000 806.700 376.050 ;
        RECT 802.800 373.500 804.900 373.800 ;
        RECT 801.000 371.700 804.900 373.500 ;
        RECT 805.800 373.050 806.700 375.000 ;
        RECT 805.800 370.950 807.900 373.050 ;
        RECT 805.800 370.800 807.300 370.950 ;
        RECT 802.200 370.050 804.000 370.500 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 797.100 368.700 804.000 370.050 ;
        RECT 804.900 369.900 807.300 370.800 ;
        RECT 811.800 370.050 813.600 371.850 ;
        RECT 824.100 370.050 825.900 371.850 ;
        RECT 827.100 370.050 828.300 383.400 ;
        RECT 840.000 380.100 841.800 381.900 ;
        RECT 842.700 378.900 844.500 389.400 ;
        RECT 842.100 377.400 844.500 378.900 ;
        RECT 847.800 377.400 849.600 390.000 ;
        RECT 860.100 383.400 861.900 389.400 ;
        RECT 863.100 383.400 864.900 390.000 ;
        RECT 842.100 370.050 843.300 377.400 ;
        RECT 848.100 370.050 849.900 371.850 ;
        RECT 860.700 370.050 861.900 383.400 ;
        RECT 862.950 375.450 865.050 376.050 ;
        RECT 862.950 374.550 870.450 375.450 ;
        RECT 862.950 373.950 865.050 374.550 ;
        RECT 863.100 370.050 864.900 371.850 ;
        RECT 797.100 367.950 799.200 368.700 ;
        RECT 769.950 365.550 774.450 367.050 ;
        RECT 769.950 364.950 774.000 365.550 ;
        RECT 716.100 361.800 720.300 362.700 ;
        RECT 677.100 354.000 678.900 357.600 ;
        RECT 680.100 354.600 681.900 357.600 ;
        RECT 683.100 354.000 684.900 357.600 ;
        RECT 695.100 354.000 696.900 357.600 ;
        RECT 698.100 354.600 699.900 357.600 ;
        RECT 701.100 354.000 702.900 357.600 ;
        RECT 713.400 354.000 715.200 360.600 ;
        RECT 718.500 354.600 720.300 361.800 ;
        RECT 731.700 360.600 732.900 362.700 ;
        RECT 760.950 362.100 765.300 363.300 ;
        RECT 731.100 354.600 732.900 360.600 ;
        RECT 734.100 359.700 741.900 361.050 ;
        RECT 734.100 354.600 735.900 359.700 ;
        RECT 737.100 354.000 738.900 358.800 ;
        RECT 740.100 354.600 741.900 359.700 ;
        RECT 755.100 360.000 762.900 360.900 ;
        RECT 764.400 360.600 765.300 362.100 ;
        RECT 755.100 354.600 756.900 360.000 ;
        RECT 758.100 354.000 759.900 359.100 ;
        RECT 761.100 355.500 762.900 360.000 ;
        RECT 764.100 356.400 765.900 360.600 ;
        RECT 767.100 355.500 768.900 360.600 ;
        RECT 782.100 357.600 783.300 367.950 ;
        RECT 797.400 366.150 799.200 367.950 ;
        RECT 802.200 365.400 804.000 367.200 ;
        RECT 801.900 363.300 804.000 365.400 ;
        RECT 797.700 362.400 804.000 363.300 ;
        RECT 804.900 364.200 806.100 369.900 ;
        RECT 807.300 367.200 809.100 369.000 ;
        RECT 811.800 367.950 813.900 370.050 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 807.000 365.100 809.100 367.200 ;
        RECT 797.700 360.600 798.900 362.400 ;
        RECT 804.900 362.100 807.900 364.200 ;
        RECT 804.900 360.600 806.100 362.100 ;
        RECT 809.100 361.500 811.200 362.700 ;
        RECT 809.100 360.600 813.900 361.500 ;
        RECT 761.100 354.600 768.900 355.500 ;
        RECT 779.100 354.000 780.900 357.600 ;
        RECT 782.100 354.600 783.900 357.600 ;
        RECT 797.100 354.600 798.900 360.600 ;
        RECT 800.100 354.000 801.900 359.700 ;
        RECT 804.600 354.600 806.400 360.600 ;
        RECT 809.100 354.000 810.900 359.700 ;
        RECT 812.100 354.600 813.900 360.600 ;
        RECT 827.100 357.600 828.300 367.950 ;
        RECT 832.950 367.050 835.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 829.950 366.000 835.050 367.050 ;
        RECT 839.100 366.150 840.900 367.950 ;
        RECT 829.950 365.550 834.450 366.000 ;
        RECT 829.950 364.950 834.000 365.550 ;
        RECT 842.100 363.600 843.300 367.950 ;
        RECT 845.100 366.150 846.900 367.950 ;
        RECT 839.700 362.700 843.300 363.600 ;
        RECT 839.700 360.600 840.900 362.700 ;
        RECT 824.100 354.000 825.900 357.600 ;
        RECT 827.100 354.600 828.900 357.600 ;
        RECT 839.100 354.600 840.900 360.600 ;
        RECT 842.100 359.700 849.900 361.050 ;
        RECT 842.100 354.600 843.900 359.700 ;
        RECT 845.100 354.000 846.900 358.800 ;
        RECT 848.100 354.600 849.900 359.700 ;
        RECT 860.700 357.600 861.900 367.950 ;
        RECT 869.550 367.050 870.450 374.550 ;
        RECT 865.950 365.550 870.450 367.050 ;
        RECT 865.950 364.950 870.000 365.550 ;
        RECT 860.100 354.600 861.900 357.600 ;
        RECT 863.100 354.000 864.900 357.600 ;
        RECT 11.100 345.000 12.900 350.400 ;
        RECT 14.100 345.900 15.900 351.000 ;
        RECT 17.100 349.500 24.900 350.400 ;
        RECT 17.100 345.000 18.900 349.500 ;
        RECT 11.100 344.100 18.900 345.000 ;
        RECT 20.100 344.400 21.900 348.600 ;
        RECT 23.100 344.400 24.900 349.500 ;
        RECT 38.400 344.400 40.200 351.000 ;
        RECT 20.400 342.900 21.300 344.400 ;
        RECT 43.500 343.200 45.300 350.400 ;
        RECT 56.400 344.400 58.200 351.000 ;
        RECT 61.500 343.200 63.300 350.400 ;
        RECT 74.100 345.000 75.900 350.400 ;
        RECT 77.100 345.900 78.900 351.000 ;
        RECT 80.100 349.500 87.900 350.400 ;
        RECT 80.100 345.000 81.900 349.500 ;
        RECT 74.100 344.100 81.900 345.000 ;
        RECT 83.100 344.400 84.900 348.600 ;
        RECT 86.100 344.400 87.900 349.500 ;
        RECT 98.700 347.400 100.500 351.000 ;
        RECT 101.700 345.600 103.500 350.400 ;
        RECT 98.400 344.400 103.500 345.600 ;
        RECT 106.200 344.400 108.000 351.000 ;
        RECT 16.950 341.700 21.300 342.900 ;
        RECT 41.100 342.300 45.300 343.200 ;
        RECT 59.100 342.300 63.300 343.200 ;
        RECT 83.400 342.900 84.300 344.400 ;
        RECT 14.250 337.050 16.050 338.850 ;
        RECT 10.950 334.950 13.050 337.050 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 16.950 337.050 18.000 341.700 ;
        RECT 19.950 337.050 21.750 338.850 ;
        RECT 38.250 337.050 40.050 338.850 ;
        RECT 41.100 337.050 42.300 342.300 ;
        RECT 44.100 337.050 45.900 338.850 ;
        RECT 56.250 337.050 58.050 338.850 ;
        RECT 59.100 337.050 60.300 342.300 ;
        RECT 79.950 341.700 84.300 342.900 ;
        RECT 62.100 337.050 63.900 338.850 ;
        RECT 77.250 337.050 79.050 338.850 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 19.950 334.950 22.050 337.050 ;
        RECT 22.950 334.950 25.050 337.050 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 337.050 81.000 341.700 ;
        RECT 82.950 337.050 84.750 338.850 ;
        RECT 98.400 337.050 99.300 344.400 ;
        RECT 121.500 342.000 123.300 350.400 ;
        RECT 120.000 340.800 123.300 342.000 ;
        RECT 128.100 341.400 129.900 351.000 ;
        RECT 140.100 347.400 141.900 350.400 ;
        RECT 143.100 347.400 144.900 351.000 ;
        RECT 100.950 337.050 102.750 338.850 ;
        RECT 107.100 337.050 108.900 338.850 ;
        RECT 120.000 337.050 120.900 340.800 ;
        RECT 122.100 337.050 123.900 338.850 ;
        RECT 128.100 337.050 129.900 338.850 ;
        RECT 140.700 337.050 141.900 347.400 ;
        RECT 158.100 344.400 159.900 350.400 ;
        RECT 158.700 342.300 159.900 344.400 ;
        RECT 161.100 345.300 162.900 350.400 ;
        RECT 164.100 346.200 165.900 351.000 ;
        RECT 167.100 345.300 168.900 350.400 ;
        RECT 179.700 347.400 181.500 351.000 ;
        RECT 182.700 345.600 184.500 350.400 ;
        RECT 161.100 343.950 168.900 345.300 ;
        RECT 179.400 344.400 184.500 345.600 ;
        RECT 187.200 344.400 189.000 351.000 ;
        RECT 158.700 341.400 162.300 342.300 ;
        RECT 158.100 337.050 159.900 338.850 ;
        RECT 161.100 337.050 162.300 341.400 ;
        RECT 164.100 337.050 165.900 338.850 ;
        RECT 179.400 337.050 180.300 344.400 ;
        RECT 181.950 342.450 184.050 343.200 ;
        RECT 196.950 342.450 199.050 343.050 ;
        RECT 181.950 341.550 199.050 342.450 ;
        RECT 202.500 342.000 204.300 350.400 ;
        RECT 181.950 341.100 184.050 341.550 ;
        RECT 196.950 340.950 199.050 341.550 ;
        RECT 201.000 340.800 204.300 342.000 ;
        RECT 209.100 341.400 210.900 351.000 ;
        RECT 221.100 347.400 222.900 351.000 ;
        RECT 224.100 347.400 225.900 350.400 ;
        RECT 227.100 347.400 228.900 351.000 ;
        RECT 181.950 337.050 183.750 338.850 ;
        RECT 188.100 337.050 189.900 338.850 ;
        RECT 201.000 337.050 201.900 340.800 ;
        RECT 203.100 337.050 204.900 338.850 ;
        RECT 209.100 337.050 210.900 338.850 ;
        RECT 224.700 337.050 225.600 347.400 ;
        RECT 242.400 344.400 244.200 351.000 ;
        RECT 247.500 343.200 249.300 350.400 ;
        RECT 245.100 342.300 249.300 343.200 ;
        RECT 260.700 343.200 262.500 350.400 ;
        RECT 265.800 344.400 267.600 351.000 ;
        RECT 281.100 347.400 282.900 351.000 ;
        RECT 284.100 347.400 285.900 350.400 ;
        RECT 260.700 342.300 264.900 343.200 ;
        RECT 242.250 337.050 244.050 338.850 ;
        RECT 245.100 337.050 246.300 342.300 ;
        RECT 248.100 337.050 249.900 338.850 ;
        RECT 260.100 337.050 261.900 338.850 ;
        RECT 263.700 337.050 264.900 342.300 ;
        RECT 265.950 337.050 267.750 338.850 ;
        RECT 284.100 337.050 285.300 347.400 ;
        RECT 296.700 343.200 298.500 350.400 ;
        RECT 301.800 344.400 303.600 351.000 ;
        RECT 314.700 343.200 316.500 350.400 ;
        RECT 319.800 344.400 321.600 351.000 ;
        RECT 335.100 345.300 336.900 350.400 ;
        RECT 338.100 346.200 339.900 351.000 ;
        RECT 341.100 345.300 342.900 350.400 ;
        RECT 335.100 343.950 342.900 345.300 ;
        RECT 344.100 344.400 345.900 350.400 ;
        RECT 356.100 345.300 357.900 350.400 ;
        RECT 359.100 346.200 360.900 351.000 ;
        RECT 362.100 345.300 363.900 350.400 ;
        RECT 296.700 342.300 300.900 343.200 ;
        RECT 314.700 342.300 318.900 343.200 ;
        RECT 344.100 342.300 345.300 344.400 ;
        RECT 356.100 343.950 363.900 345.300 ;
        RECT 365.100 344.400 366.900 350.400 ;
        RECT 377.400 344.400 379.200 351.000 ;
        RECT 365.100 342.300 366.300 344.400 ;
        RECT 382.500 343.200 384.300 350.400 ;
        RECT 296.100 337.050 297.900 338.850 ;
        RECT 299.700 337.050 300.900 342.300 ;
        RECT 309.000 339.450 313.050 340.050 ;
        RECT 301.950 337.050 303.750 338.850 ;
        RECT 308.550 337.950 313.050 339.450 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 100.950 334.950 103.050 337.050 ;
        RECT 103.950 334.950 106.050 337.050 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 121.950 334.950 124.050 337.050 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 127.950 334.950 130.050 337.050 ;
        RECT 139.950 334.950 142.050 337.050 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 265.950 334.950 268.050 337.050 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 283.950 334.950 286.050 337.050 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 11.100 333.150 12.900 334.950 ;
        RECT 16.950 327.600 18.000 334.950 ;
        RECT 22.950 333.150 24.750 334.950 ;
        RECT 11.100 315.000 12.900 327.600 ;
        RECT 15.600 315.600 18.900 327.600 ;
        RECT 21.600 315.000 23.400 327.600 ;
        RECT 41.100 321.600 42.300 334.950 ;
        RECT 59.100 321.600 60.300 334.950 ;
        RECT 74.100 333.150 75.900 334.950 ;
        RECT 79.950 327.600 81.000 334.950 ;
        RECT 85.950 333.150 87.750 334.950 ;
        RECT 98.400 327.600 99.300 334.950 ;
        RECT 103.950 333.150 105.750 334.950 ;
        RECT 38.100 315.000 39.900 321.600 ;
        RECT 41.100 315.600 42.900 321.600 ;
        RECT 44.100 315.000 45.900 321.600 ;
        RECT 56.100 315.000 57.900 321.600 ;
        RECT 59.100 315.600 60.900 321.600 ;
        RECT 62.100 315.000 63.900 321.600 ;
        RECT 74.100 315.000 75.900 327.600 ;
        RECT 78.600 315.600 81.900 327.600 ;
        RECT 84.600 315.000 86.400 327.600 ;
        RECT 98.100 315.600 99.900 327.600 ;
        RECT 101.100 326.700 108.900 327.600 ;
        RECT 101.100 315.600 102.900 326.700 ;
        RECT 104.100 315.000 105.900 325.800 ;
        RECT 107.100 315.600 108.900 326.700 ;
        RECT 120.000 322.800 120.900 334.950 ;
        RECT 125.100 333.150 126.900 334.950 ;
        RECT 120.000 321.900 126.600 322.800 ;
        RECT 120.000 321.600 120.900 321.900 ;
        RECT 119.100 315.600 120.900 321.600 ;
        RECT 125.100 321.600 126.600 321.900 ;
        RECT 140.700 321.600 141.900 334.950 ;
        RECT 143.100 333.150 144.900 334.950 ;
        RECT 161.100 327.600 162.300 334.950 ;
        RECT 167.100 333.150 168.900 334.950 ;
        RECT 179.400 327.600 180.300 334.950 ;
        RECT 184.950 333.150 186.750 334.950 ;
        RECT 161.100 326.100 163.500 327.600 ;
        RECT 159.000 323.100 160.800 324.900 ;
        RECT 122.100 315.000 123.900 321.000 ;
        RECT 125.100 315.600 126.900 321.600 ;
        RECT 128.100 315.000 129.900 321.600 ;
        RECT 140.100 315.600 141.900 321.600 ;
        RECT 143.100 315.000 144.900 321.600 ;
        RECT 158.700 315.000 160.500 321.600 ;
        RECT 161.700 315.600 163.500 326.100 ;
        RECT 166.800 315.000 168.600 327.600 ;
        RECT 179.100 315.600 180.900 327.600 ;
        RECT 182.100 326.700 189.900 327.600 ;
        RECT 182.100 315.600 183.900 326.700 ;
        RECT 185.100 315.000 186.900 325.800 ;
        RECT 188.100 315.600 189.900 326.700 ;
        RECT 201.000 322.800 201.900 334.950 ;
        RECT 206.100 333.150 207.900 334.950 ;
        RECT 221.100 333.150 222.900 334.950 ;
        RECT 224.700 327.600 225.600 334.950 ;
        RECT 226.950 333.150 228.750 334.950 ;
        RECT 222.000 326.400 225.600 327.600 ;
        RECT 201.000 321.900 207.600 322.800 ;
        RECT 201.000 321.600 201.900 321.900 ;
        RECT 200.100 315.600 201.900 321.600 ;
        RECT 206.100 321.600 207.600 321.900 ;
        RECT 203.100 315.000 204.900 321.000 ;
        RECT 206.100 315.600 207.900 321.600 ;
        RECT 209.100 315.000 210.900 321.600 ;
        RECT 222.000 315.600 223.800 326.400 ;
        RECT 227.100 315.000 228.900 327.600 ;
        RECT 245.100 321.600 246.300 334.950 ;
        RECT 263.700 321.600 264.900 334.950 ;
        RECT 281.100 333.150 282.900 334.950 ;
        RECT 284.100 321.600 285.300 334.950 ;
        RECT 299.700 321.600 300.900 334.950 ;
        RECT 308.550 333.450 309.450 337.950 ;
        RECT 314.100 337.050 315.900 338.850 ;
        RECT 317.700 337.050 318.900 342.300 ;
        RECT 341.700 341.400 345.300 342.300 ;
        RECT 362.700 341.400 366.300 342.300 ;
        RECT 380.100 342.300 384.300 343.200 ;
        RECT 386.550 344.400 388.350 350.400 ;
        RECT 389.850 344.400 391.650 351.000 ;
        RECT 394.950 347.400 396.750 350.400 ;
        RECT 399.450 347.400 401.250 351.000 ;
        RECT 402.450 347.400 404.250 350.400 ;
        RECT 405.750 347.400 407.550 351.000 ;
        RECT 410.250 348.300 412.050 350.400 ;
        RECT 410.250 347.400 413.850 348.300 ;
        RECT 394.350 345.300 396.750 347.400 ;
        RECT 403.200 346.500 404.250 347.400 ;
        RECT 410.250 346.800 414.150 347.400 ;
        RECT 403.200 345.450 408.150 346.500 ;
        RECT 406.350 344.700 408.150 345.450 ;
        RECT 319.950 337.050 321.750 338.850 ;
        RECT 338.100 337.050 339.900 338.850 ;
        RECT 341.700 337.050 342.900 341.400 ;
        RECT 344.100 337.050 345.900 338.850 ;
        RECT 359.100 337.050 360.900 338.850 ;
        RECT 362.700 337.050 363.900 341.400 ;
        RECT 365.100 337.050 366.900 338.850 ;
        RECT 377.250 337.050 379.050 338.850 ;
        RECT 380.100 337.050 381.300 342.300 ;
        RECT 383.100 337.050 384.900 338.850 ;
        RECT 386.550 337.050 387.750 344.400 ;
        RECT 409.350 343.800 411.150 345.600 ;
        RECT 412.050 345.300 414.150 346.800 ;
        RECT 415.050 344.400 416.850 351.000 ;
        RECT 418.050 346.200 419.850 350.400 ;
        RECT 418.050 344.400 420.450 346.200 ;
        RECT 431.100 344.400 432.900 350.400 ;
        RECT 434.100 344.400 435.900 351.000 ;
        RECT 437.550 344.400 439.350 350.400 ;
        RECT 440.850 344.400 442.650 351.000 ;
        RECT 445.950 347.400 447.750 350.400 ;
        RECT 450.450 347.400 452.250 351.000 ;
        RECT 453.450 347.400 455.250 350.400 ;
        RECT 456.750 347.400 458.550 351.000 ;
        RECT 461.250 348.300 463.050 350.400 ;
        RECT 461.250 347.400 464.850 348.300 ;
        RECT 445.350 345.300 447.750 347.400 ;
        RECT 454.200 346.500 455.250 347.400 ;
        RECT 461.250 346.800 465.150 347.400 ;
        RECT 454.200 345.450 459.150 346.500 ;
        RECT 457.350 344.700 459.150 345.450 ;
        RECT 399.150 342.000 400.950 342.600 ;
        RECT 410.100 342.000 411.150 343.800 ;
        RECT 399.150 340.800 411.150 342.000 ;
        RECT 313.950 334.950 316.050 337.050 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 305.550 332.550 309.450 333.450 ;
        RECT 305.550 331.050 306.450 332.550 ;
        RECT 301.950 329.550 306.450 331.050 ;
        RECT 301.950 328.950 306.000 329.550 ;
        RECT 317.700 321.600 318.900 334.950 ;
        RECT 335.100 333.150 336.900 334.950 ;
        RECT 341.700 327.600 342.900 334.950 ;
        RECT 349.950 334.050 352.050 337.050 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 358.950 334.950 361.050 337.050 ;
        RECT 361.950 334.950 364.050 337.050 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 382.950 334.950 385.050 337.050 ;
        RECT 386.550 335.250 392.850 337.050 ;
        RECT 386.550 334.950 391.050 335.250 ;
        RECT 349.950 333.000 355.050 334.050 ;
        RECT 356.100 333.150 357.900 334.950 ;
        RECT 350.550 332.550 355.050 333.000 ;
        RECT 351.000 331.950 355.050 332.550 ;
        RECT 362.700 327.600 363.900 334.950 ;
        RECT 242.100 315.000 243.900 321.600 ;
        RECT 245.100 315.600 246.900 321.600 ;
        RECT 248.100 315.000 249.900 321.600 ;
        RECT 260.100 315.000 261.900 321.600 ;
        RECT 263.100 315.600 264.900 321.600 ;
        RECT 266.100 315.000 267.900 321.600 ;
        RECT 281.100 315.000 282.900 321.600 ;
        RECT 284.100 315.600 285.900 321.600 ;
        RECT 296.100 315.000 297.900 321.600 ;
        RECT 299.100 315.600 300.900 321.600 ;
        RECT 302.100 315.000 303.900 321.600 ;
        RECT 314.100 315.000 315.900 321.600 ;
        RECT 317.100 315.600 318.900 321.600 ;
        RECT 320.100 315.000 321.900 321.600 ;
        RECT 335.400 315.000 337.200 327.600 ;
        RECT 340.500 326.100 342.900 327.600 ;
        RECT 340.500 315.600 342.300 326.100 ;
        RECT 343.200 323.100 345.000 324.900 ;
        RECT 343.500 315.000 345.300 321.600 ;
        RECT 356.400 315.000 358.200 327.600 ;
        RECT 361.500 326.100 363.900 327.600 ;
        RECT 361.500 315.600 363.300 326.100 ;
        RECT 364.200 323.100 366.000 324.900 ;
        RECT 380.100 321.600 381.300 334.950 ;
        RECT 386.550 327.600 387.750 334.950 ;
        RECT 388.650 332.100 390.450 332.250 ;
        RECT 394.350 332.100 396.450 332.400 ;
        RECT 388.650 330.900 396.450 332.100 ;
        RECT 388.650 330.450 390.450 330.900 ;
        RECT 394.350 330.300 396.450 330.900 ;
        RECT 399.150 328.200 400.050 340.800 ;
        RECT 410.100 339.600 418.050 340.800 ;
        RECT 410.100 339.000 411.900 339.600 ;
        RECT 413.100 337.800 414.900 338.400 ;
        RECT 406.800 336.600 414.900 337.800 ;
        RECT 416.250 337.050 418.050 339.600 ;
        RECT 406.800 334.950 408.900 336.600 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 408.750 329.700 410.550 330.000 ;
        RECT 419.550 329.700 420.450 344.400 ;
        RECT 431.700 337.050 432.900 344.400 ;
        RECT 434.100 337.050 435.900 338.850 ;
        RECT 437.550 337.050 438.750 344.400 ;
        RECT 460.350 343.800 462.150 345.600 ;
        RECT 463.050 345.300 465.150 346.800 ;
        RECT 466.050 344.400 467.850 351.000 ;
        RECT 469.050 346.200 470.850 350.400 ;
        RECT 469.050 344.400 471.450 346.200 ;
        RECT 450.150 342.000 451.950 342.600 ;
        RECT 461.100 342.000 462.150 343.800 ;
        RECT 450.150 340.800 462.150 342.000 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 437.550 335.250 443.850 337.050 ;
        RECT 437.550 334.950 442.050 335.250 ;
        RECT 408.750 329.100 420.450 329.700 ;
        RECT 364.500 315.000 366.300 321.600 ;
        RECT 377.100 315.000 378.900 321.600 ;
        RECT 380.100 315.600 381.900 321.600 ;
        RECT 383.100 315.000 384.900 321.600 ;
        RECT 386.550 315.600 388.350 327.600 ;
        RECT 389.550 315.000 391.350 327.600 ;
        RECT 395.250 327.300 400.050 328.200 ;
        RECT 402.150 328.500 420.450 329.100 ;
        RECT 402.150 328.200 410.550 328.500 ;
        RECT 395.250 326.400 396.450 327.300 ;
        RECT 393.450 324.600 396.450 326.400 ;
        RECT 397.350 326.100 399.150 326.400 ;
        RECT 402.150 326.100 403.050 328.200 ;
        RECT 419.550 327.600 420.450 328.500 ;
        RECT 431.700 327.600 432.900 334.950 ;
        RECT 437.550 327.600 438.750 334.950 ;
        RECT 439.650 332.100 441.450 332.250 ;
        RECT 445.350 332.100 447.450 332.400 ;
        RECT 439.650 330.900 447.450 332.100 ;
        RECT 439.650 330.450 441.450 330.900 ;
        RECT 445.350 330.300 447.450 330.900 ;
        RECT 450.150 328.200 451.050 340.800 ;
        RECT 461.100 339.600 469.050 340.800 ;
        RECT 461.100 339.000 462.900 339.600 ;
        RECT 464.100 337.800 465.900 338.400 ;
        RECT 457.800 336.600 465.900 337.800 ;
        RECT 467.250 337.050 469.050 339.600 ;
        RECT 457.800 334.950 459.900 336.600 ;
        RECT 466.950 334.950 469.050 337.050 ;
        RECT 459.750 329.700 461.550 330.000 ;
        RECT 470.550 329.700 471.450 344.400 ;
        RECT 459.750 329.100 471.450 329.700 ;
        RECT 397.350 325.200 403.050 326.100 ;
        RECT 403.950 326.700 405.750 327.300 ;
        RECT 403.950 325.500 411.750 326.700 ;
        RECT 397.350 324.600 399.150 325.200 ;
        RECT 409.650 324.600 411.750 325.500 ;
        RECT 394.350 321.600 396.450 323.700 ;
        RECT 400.950 323.550 402.750 324.300 ;
        RECT 405.750 323.550 407.550 324.300 ;
        RECT 400.950 322.500 407.550 323.550 ;
        RECT 394.350 315.600 396.150 321.600 ;
        RECT 398.850 315.000 400.650 321.600 ;
        RECT 401.850 315.600 403.650 322.500 ;
        RECT 404.850 315.000 406.650 321.600 ;
        RECT 409.650 315.600 411.450 324.600 ;
        RECT 415.050 315.000 416.850 327.600 ;
        RECT 418.050 325.800 420.450 327.600 ;
        RECT 418.050 315.600 419.850 325.800 ;
        RECT 431.100 315.600 432.900 327.600 ;
        RECT 434.100 315.000 435.900 327.600 ;
        RECT 437.550 315.600 439.350 327.600 ;
        RECT 440.550 315.000 442.350 327.600 ;
        RECT 446.250 327.300 451.050 328.200 ;
        RECT 453.150 328.500 471.450 329.100 ;
        RECT 453.150 328.200 461.550 328.500 ;
        RECT 446.250 326.400 447.450 327.300 ;
        RECT 444.450 324.600 447.450 326.400 ;
        RECT 448.350 326.100 450.150 326.400 ;
        RECT 453.150 326.100 454.050 328.200 ;
        RECT 470.550 327.600 471.450 328.500 ;
        RECT 448.350 325.200 454.050 326.100 ;
        RECT 454.950 326.700 456.750 327.300 ;
        RECT 454.950 325.500 462.750 326.700 ;
        RECT 448.350 324.600 450.150 325.200 ;
        RECT 460.650 324.600 462.750 325.500 ;
        RECT 445.350 321.600 447.450 323.700 ;
        RECT 451.950 323.550 453.750 324.300 ;
        RECT 456.750 323.550 458.550 324.300 ;
        RECT 451.950 322.500 458.550 323.550 ;
        RECT 445.350 315.600 447.150 321.600 ;
        RECT 449.850 315.000 451.650 321.600 ;
        RECT 452.850 315.600 454.650 322.500 ;
        RECT 455.850 315.000 457.650 321.600 ;
        RECT 460.650 315.600 462.450 324.600 ;
        RECT 466.050 315.000 467.850 327.600 ;
        RECT 469.050 325.800 471.450 327.600 ;
        RECT 473.550 344.400 475.350 350.400 ;
        RECT 476.850 344.400 478.650 351.000 ;
        RECT 481.950 347.400 483.750 350.400 ;
        RECT 486.450 347.400 488.250 351.000 ;
        RECT 489.450 347.400 491.250 350.400 ;
        RECT 492.750 347.400 494.550 351.000 ;
        RECT 497.250 348.300 499.050 350.400 ;
        RECT 497.250 347.400 500.850 348.300 ;
        RECT 481.350 345.300 483.750 347.400 ;
        RECT 490.200 346.500 491.250 347.400 ;
        RECT 497.250 346.800 501.150 347.400 ;
        RECT 490.200 345.450 495.150 346.500 ;
        RECT 493.350 344.700 495.150 345.450 ;
        RECT 473.550 337.050 474.750 344.400 ;
        RECT 496.350 343.800 498.150 345.600 ;
        RECT 499.050 345.300 501.150 346.800 ;
        RECT 502.050 344.400 503.850 351.000 ;
        RECT 505.050 346.200 506.850 350.400 ;
        RECT 505.050 344.400 507.450 346.200 ;
        RECT 486.150 342.000 487.950 342.600 ;
        RECT 497.100 342.000 498.150 343.800 ;
        RECT 486.150 340.800 498.150 342.000 ;
        RECT 473.550 335.250 479.850 337.050 ;
        RECT 473.550 334.950 478.050 335.250 ;
        RECT 473.550 327.600 474.750 334.950 ;
        RECT 475.650 332.100 477.450 332.250 ;
        RECT 481.350 332.100 483.450 332.400 ;
        RECT 475.650 330.900 483.450 332.100 ;
        RECT 475.650 330.450 477.450 330.900 ;
        RECT 481.350 330.300 483.450 330.900 ;
        RECT 486.150 328.200 487.050 340.800 ;
        RECT 497.100 339.600 505.050 340.800 ;
        RECT 497.100 339.000 498.900 339.600 ;
        RECT 500.100 337.800 501.900 338.400 ;
        RECT 493.800 336.600 501.900 337.800 ;
        RECT 503.250 337.050 505.050 339.600 ;
        RECT 493.800 334.950 495.900 336.600 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 495.750 329.700 497.550 330.000 ;
        RECT 506.550 329.700 507.450 344.400 ;
        RECT 518.100 345.300 519.900 350.400 ;
        RECT 521.100 346.200 522.900 351.000 ;
        RECT 524.100 345.300 525.900 350.400 ;
        RECT 518.100 343.950 525.900 345.300 ;
        RECT 527.100 344.400 528.900 350.400 ;
        RECT 539.100 344.400 540.900 350.400 ;
        RECT 527.100 342.300 528.300 344.400 ;
        RECT 524.700 341.400 528.300 342.300 ;
        RECT 539.700 342.300 540.900 344.400 ;
        RECT 542.100 345.300 543.900 350.400 ;
        RECT 545.100 346.200 546.900 351.000 ;
        RECT 548.100 345.300 549.900 350.400 ;
        RECT 542.100 343.950 549.900 345.300 ;
        RECT 560.400 344.400 562.200 351.000 ;
        RECT 565.500 343.200 567.300 350.400 ;
        RECT 563.100 342.300 567.300 343.200 ;
        RECT 578.700 343.200 580.500 350.400 ;
        RECT 583.800 344.400 585.600 351.000 ;
        RECT 599.100 344.400 600.900 350.400 ;
        RECT 578.700 342.300 582.900 343.200 ;
        RECT 539.700 341.400 543.300 342.300 ;
        RECT 521.100 337.050 522.900 338.850 ;
        RECT 524.700 337.050 525.900 341.400 ;
        RECT 527.100 337.050 528.900 338.850 ;
        RECT 539.100 337.050 540.900 338.850 ;
        RECT 542.100 337.050 543.300 341.400 ;
        RECT 545.100 337.050 546.900 338.850 ;
        RECT 560.250 337.050 562.050 338.850 ;
        RECT 563.100 337.050 564.300 342.300 ;
        RECT 573.000 339.450 577.050 340.050 ;
        RECT 566.100 337.050 567.900 338.850 ;
        RECT 572.550 337.950 577.050 339.450 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 526.950 334.950 529.050 337.050 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 518.100 333.150 519.900 334.950 ;
        RECT 495.750 329.100 507.450 329.700 ;
        RECT 469.050 315.600 470.850 325.800 ;
        RECT 473.550 315.600 475.350 327.600 ;
        RECT 476.550 315.000 478.350 327.600 ;
        RECT 482.250 327.300 487.050 328.200 ;
        RECT 489.150 328.500 507.450 329.100 ;
        RECT 508.950 330.450 511.050 331.050 ;
        RECT 520.950 330.450 523.050 331.050 ;
        RECT 508.950 329.550 523.050 330.450 ;
        RECT 508.950 328.950 511.050 329.550 ;
        RECT 520.950 328.950 523.050 329.550 ;
        RECT 489.150 328.200 497.550 328.500 ;
        RECT 482.250 326.400 483.450 327.300 ;
        RECT 480.450 324.600 483.450 326.400 ;
        RECT 484.350 326.100 486.150 326.400 ;
        RECT 489.150 326.100 490.050 328.200 ;
        RECT 506.550 327.600 507.450 328.500 ;
        RECT 524.700 327.600 525.900 334.950 ;
        RECT 484.350 325.200 490.050 326.100 ;
        RECT 490.950 326.700 492.750 327.300 ;
        RECT 490.950 325.500 498.750 326.700 ;
        RECT 484.350 324.600 486.150 325.200 ;
        RECT 496.650 324.600 498.750 325.500 ;
        RECT 481.350 321.600 483.450 323.700 ;
        RECT 487.950 323.550 489.750 324.300 ;
        RECT 492.750 323.550 494.550 324.300 ;
        RECT 487.950 322.500 494.550 323.550 ;
        RECT 481.350 315.600 483.150 321.600 ;
        RECT 485.850 315.000 487.650 321.600 ;
        RECT 488.850 315.600 490.650 322.500 ;
        RECT 491.850 315.000 493.650 321.600 ;
        RECT 496.650 315.600 498.450 324.600 ;
        RECT 502.050 315.000 503.850 327.600 ;
        RECT 505.050 325.800 507.450 327.600 ;
        RECT 505.050 315.600 506.850 325.800 ;
        RECT 518.400 315.000 520.200 327.600 ;
        RECT 523.500 326.100 525.900 327.600 ;
        RECT 542.100 327.600 543.300 334.950 ;
        RECT 548.100 333.150 549.900 334.950 ;
        RECT 544.950 330.450 547.050 331.050 ;
        RECT 544.950 329.550 552.450 330.450 ;
        RECT 544.950 328.950 547.050 329.550 ;
        RECT 542.100 326.100 544.500 327.600 ;
        RECT 523.500 315.600 525.300 326.100 ;
        RECT 526.200 323.100 528.000 324.900 ;
        RECT 540.000 323.100 541.800 324.900 ;
        RECT 526.500 315.000 528.300 321.600 ;
        RECT 539.700 315.000 541.500 321.600 ;
        RECT 542.700 315.600 544.500 326.100 ;
        RECT 547.800 315.000 549.600 327.600 ;
        RECT 551.550 327.450 552.450 329.550 ;
        RECT 559.950 327.450 562.050 328.050 ;
        RECT 551.550 326.550 562.050 327.450 ;
        RECT 559.950 325.950 562.050 326.550 ;
        RECT 563.100 321.600 564.300 334.950 ;
        RECT 572.550 334.050 573.450 337.950 ;
        RECT 578.100 337.050 579.900 338.850 ;
        RECT 581.700 337.050 582.900 342.300 ;
        RECT 583.950 342.450 586.050 343.050 ;
        RECT 592.950 342.450 595.050 343.050 ;
        RECT 583.950 341.550 595.050 342.450 ;
        RECT 583.950 340.950 586.050 341.550 ;
        RECT 592.950 340.950 595.050 341.550 ;
        RECT 599.700 342.300 600.900 344.400 ;
        RECT 602.100 345.300 603.900 350.400 ;
        RECT 605.100 346.200 606.900 351.000 ;
        RECT 608.100 345.300 609.900 350.400 ;
        RECT 602.100 343.950 609.900 345.300 ;
        RECT 620.700 343.200 622.500 350.400 ;
        RECT 625.800 344.400 627.600 351.000 ;
        RECT 638.100 345.300 639.900 350.400 ;
        RECT 641.100 346.200 642.900 351.000 ;
        RECT 644.100 345.300 645.900 350.400 ;
        RECT 638.100 343.950 645.900 345.300 ;
        RECT 647.100 344.400 648.900 350.400 ;
        RECT 659.100 347.400 660.900 351.000 ;
        RECT 662.100 347.400 663.900 350.400 ;
        RECT 665.100 347.400 666.900 351.000 ;
        RECT 620.700 342.300 624.900 343.200 ;
        RECT 647.100 342.300 648.300 344.400 ;
        RECT 599.700 341.400 603.300 342.300 ;
        RECT 583.950 337.050 585.750 338.850 ;
        RECT 599.100 337.050 600.900 338.850 ;
        RECT 602.100 337.050 603.300 341.400 ;
        RECT 605.100 337.050 606.900 338.850 ;
        RECT 620.100 337.050 621.900 338.850 ;
        RECT 623.700 337.050 624.900 342.300 ;
        RECT 644.700 341.400 648.300 342.300 ;
        RECT 633.000 339.450 637.050 340.050 ;
        RECT 625.950 337.050 627.750 338.850 ;
        RECT 632.550 337.950 637.050 339.450 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 568.950 332.550 573.450 334.050 ;
        RECT 568.950 331.950 573.000 332.550 ;
        RECT 565.950 330.450 568.050 330.750 ;
        RECT 577.950 330.450 580.050 331.050 ;
        RECT 565.950 329.550 580.050 330.450 ;
        RECT 565.950 328.650 568.050 329.550 ;
        RECT 577.950 328.950 580.050 329.550 ;
        RECT 581.700 321.600 582.900 334.950 ;
        RECT 602.100 327.600 603.300 334.950 ;
        RECT 608.100 333.150 609.900 334.950 ;
        RECT 602.100 326.100 604.500 327.600 ;
        RECT 600.000 323.100 601.800 324.900 ;
        RECT 560.100 315.000 561.900 321.600 ;
        RECT 563.100 315.600 564.900 321.600 ;
        RECT 566.100 315.000 567.900 321.600 ;
        RECT 578.100 315.000 579.900 321.600 ;
        RECT 581.100 315.600 582.900 321.600 ;
        RECT 584.100 315.000 585.900 321.600 ;
        RECT 599.700 315.000 601.500 321.600 ;
        RECT 602.700 315.600 604.500 326.100 ;
        RECT 607.800 315.000 609.600 327.600 ;
        RECT 623.700 321.600 624.900 334.950 ;
        RECT 632.550 334.050 633.450 337.950 ;
        RECT 641.100 337.050 642.900 338.850 ;
        RECT 644.700 337.050 645.900 341.400 ;
        RECT 649.950 339.450 654.000 340.050 ;
        RECT 647.100 337.050 648.900 338.850 ;
        RECT 649.950 337.950 654.450 339.450 ;
        RECT 637.950 334.950 640.050 337.050 ;
        RECT 640.950 334.950 643.050 337.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 632.550 332.550 637.050 334.050 ;
        RECT 638.100 333.150 639.900 334.950 ;
        RECT 633.000 331.950 637.050 332.550 ;
        RECT 644.700 327.600 645.900 334.950 ;
        RECT 653.550 334.050 654.450 337.950 ;
        RECT 662.400 337.050 663.300 347.400 ;
        RECT 680.400 344.400 682.200 351.000 ;
        RECT 698.100 350.400 699.300 351.000 ;
        RECT 685.500 343.200 687.300 350.400 ;
        RECT 698.100 347.400 699.900 350.400 ;
        RECT 701.100 347.400 702.900 350.400 ;
        RECT 688.950 343.950 691.050 346.050 ;
        RECT 664.950 342.450 667.050 343.050 ;
        RECT 670.950 342.450 673.050 343.050 ;
        RECT 679.950 342.450 682.050 343.050 ;
        RECT 664.950 341.550 682.050 342.450 ;
        RECT 664.950 340.950 667.050 341.550 ;
        RECT 670.950 340.950 673.050 341.550 ;
        RECT 679.950 340.950 682.050 341.550 ;
        RECT 683.100 342.300 687.300 343.200 ;
        RECT 680.250 337.050 682.050 338.850 ;
        RECT 683.100 337.050 684.300 342.300 ;
        RECT 689.550 339.450 690.450 343.950 ;
        RECT 701.400 343.200 702.300 347.400 ;
        RECT 704.100 345.000 705.900 351.000 ;
        RECT 707.100 344.400 708.900 350.400 ;
        RECT 701.400 342.300 706.800 343.200 ;
        RECT 704.700 341.400 706.800 342.300 ;
        RECT 686.100 337.050 687.900 338.850 ;
        RECT 689.550 338.550 693.450 339.450 ;
        RECT 658.950 334.950 661.050 337.050 ;
        RECT 661.950 334.950 664.050 337.050 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 679.950 334.950 682.050 337.050 ;
        RECT 682.950 334.950 685.050 337.050 ;
        RECT 685.950 334.950 688.050 337.050 ;
        RECT 653.550 332.550 658.050 334.050 ;
        RECT 659.250 333.150 661.050 334.950 ;
        RECT 654.000 331.950 658.050 332.550 ;
        RECT 662.400 327.600 663.300 334.950 ;
        RECT 665.100 333.150 666.900 334.950 ;
        RECT 664.950 330.450 667.050 331.050 ;
        RECT 670.950 330.450 673.050 331.050 ;
        RECT 664.950 329.550 673.050 330.450 ;
        RECT 664.950 328.950 667.050 329.550 ;
        RECT 670.950 328.950 673.050 329.550 ;
        RECT 620.100 315.000 621.900 321.600 ;
        RECT 623.100 315.600 624.900 321.600 ;
        RECT 626.100 315.000 627.900 321.600 ;
        RECT 638.400 315.000 640.200 327.600 ;
        RECT 643.500 326.100 645.900 327.600 ;
        RECT 643.500 315.600 645.300 326.100 ;
        RECT 646.200 323.100 648.000 324.900 ;
        RECT 646.500 315.000 648.300 321.600 ;
        RECT 659.100 315.000 660.900 327.600 ;
        RECT 662.400 326.400 666.000 327.600 ;
        RECT 664.200 315.600 666.000 326.400 ;
        RECT 683.100 321.600 684.300 334.950 ;
        RECT 692.550 334.050 693.450 338.550 ;
        RECT 698.400 337.050 700.200 338.850 ;
        RECT 698.100 334.950 700.200 337.050 ;
        RECT 701.400 334.950 703.500 337.050 ;
        RECT 688.950 332.550 693.450 334.050 ;
        RECT 702.000 333.150 703.800 334.950 ;
        RECT 688.950 331.950 693.000 332.550 ;
        RECT 704.700 330.900 705.600 341.400 ;
        RECT 708.000 337.050 708.900 344.400 ;
        RECT 719.100 341.400 720.900 351.000 ;
        RECT 725.700 342.000 727.500 350.400 ;
        RECT 740.100 344.400 741.900 350.400 ;
        RECT 740.700 342.300 741.900 344.400 ;
        RECT 743.100 345.300 744.900 350.400 ;
        RECT 746.100 346.200 747.900 351.000 ;
        RECT 749.100 345.300 750.900 350.400 ;
        RECT 743.100 343.950 750.900 345.300 ;
        RECT 764.100 344.400 765.900 350.400 ;
        RECT 764.700 342.300 765.900 344.400 ;
        RECT 767.100 345.300 768.900 350.400 ;
        RECT 770.100 346.200 771.900 351.000 ;
        RECT 773.100 345.300 774.900 350.400 ;
        RECT 767.100 343.950 774.900 345.300 ;
        RECT 785.700 343.200 787.500 350.400 ;
        RECT 790.800 344.400 792.600 351.000 ;
        RECT 785.700 342.300 789.900 343.200 ;
        RECT 725.700 340.800 729.000 342.000 ;
        RECT 740.700 341.400 744.300 342.300 ;
        RECT 764.700 341.400 768.300 342.300 ;
        RECT 719.100 337.050 720.900 338.850 ;
        RECT 725.100 337.050 726.900 338.850 ;
        RECT 728.100 337.050 729.000 340.800 ;
        RECT 730.950 339.450 735.000 340.050 ;
        RECT 730.950 337.950 735.450 339.450 ;
        RECT 706.800 334.950 708.900 337.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 727.950 334.950 730.050 337.050 ;
        RECT 704.100 330.300 705.900 330.900 ;
        RECT 698.100 329.100 705.900 330.300 ;
        RECT 698.100 327.600 699.300 329.100 ;
        RECT 706.800 327.600 708.000 334.950 ;
        RECT 722.100 333.150 723.900 334.950 ;
        RECT 685.950 324.450 688.050 324.900 ;
        RECT 694.950 324.450 697.050 325.050 ;
        RECT 685.950 323.550 697.050 324.450 ;
        RECT 685.950 322.800 688.050 323.550 ;
        RECT 694.950 322.950 697.050 323.550 ;
        RECT 680.100 315.000 681.900 321.600 ;
        RECT 683.100 315.600 684.900 321.600 ;
        RECT 686.100 315.000 687.900 321.600 ;
        RECT 698.100 315.600 699.900 327.600 ;
        RECT 702.600 315.000 704.400 327.600 ;
        RECT 705.600 326.100 708.000 327.600 ;
        RECT 705.600 315.600 707.400 326.100 ;
        RECT 728.100 322.800 729.000 334.950 ;
        RECT 734.550 334.050 735.450 337.950 ;
        RECT 740.100 337.050 741.900 338.850 ;
        RECT 743.100 337.050 744.300 341.400 ;
        RECT 751.950 339.450 756.000 340.050 ;
        RECT 746.100 337.050 747.900 338.850 ;
        RECT 751.950 337.950 756.450 339.450 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 734.550 332.550 739.050 334.050 ;
        RECT 735.000 331.950 739.050 332.550 ;
        RECT 743.100 327.600 744.300 334.950 ;
        RECT 749.100 333.150 750.900 334.950 ;
        RECT 755.550 334.050 756.450 337.950 ;
        RECT 764.100 337.050 765.900 338.850 ;
        RECT 767.100 337.050 768.300 341.400 ;
        RECT 770.100 337.050 771.900 338.850 ;
        RECT 785.100 337.050 786.900 338.850 ;
        RECT 788.700 337.050 789.900 342.300 ;
        RECT 803.100 341.400 804.900 351.000 ;
        RECT 809.700 342.000 811.500 350.400 ;
        RECT 825.000 344.400 826.800 351.000 ;
        RECT 829.500 345.600 831.300 350.400 ;
        RECT 832.500 347.400 834.300 351.000 ;
        RECT 845.100 347.400 846.900 350.400 ;
        RECT 829.500 344.400 834.600 345.600 ;
        RECT 817.950 342.450 820.050 343.050 ;
        RECT 826.950 342.450 829.050 342.900 ;
        RECT 809.700 340.800 813.000 342.000 ;
        RECT 817.950 341.550 829.050 342.450 ;
        RECT 817.950 340.950 820.050 341.550 ;
        RECT 826.950 340.800 829.050 341.550 ;
        RECT 790.950 337.050 792.750 338.850 ;
        RECT 803.100 337.050 804.900 338.850 ;
        RECT 809.100 337.050 810.900 338.850 ;
        RECT 812.100 337.050 813.000 340.800 ;
        RECT 814.950 339.450 819.000 340.050 ;
        RECT 814.950 337.950 819.450 339.450 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 751.950 332.550 756.450 334.050 ;
        RECT 751.950 331.950 756.000 332.550 ;
        RECT 767.100 327.600 768.300 334.950 ;
        RECT 773.100 333.150 774.900 334.950 ;
        RECT 743.100 326.100 745.500 327.600 ;
        RECT 741.000 323.100 742.800 324.900 ;
        RECT 722.400 321.900 729.000 322.800 ;
        RECT 722.400 321.600 723.900 321.900 ;
        RECT 719.100 315.000 720.900 321.600 ;
        RECT 722.100 315.600 723.900 321.600 ;
        RECT 728.100 321.600 729.000 321.900 ;
        RECT 725.100 315.000 726.900 321.000 ;
        RECT 728.100 315.600 729.900 321.600 ;
        RECT 740.700 315.000 742.500 321.600 ;
        RECT 743.700 315.600 745.500 326.100 ;
        RECT 748.800 315.000 750.600 327.600 ;
        RECT 767.100 326.100 769.500 327.600 ;
        RECT 765.000 323.100 766.800 324.900 ;
        RECT 764.700 315.000 766.500 321.600 ;
        RECT 767.700 315.600 769.500 326.100 ;
        RECT 772.800 315.000 774.600 327.600 ;
        RECT 788.700 321.600 789.900 334.950 ;
        RECT 806.100 333.150 807.900 334.950 ;
        RECT 812.100 322.800 813.000 334.950 ;
        RECT 818.550 333.450 819.450 337.950 ;
        RECT 824.100 337.050 825.900 338.850 ;
        RECT 830.250 337.050 832.050 338.850 ;
        RECT 833.700 337.050 834.600 344.400 ;
        RECT 845.100 343.500 846.300 347.400 ;
        RECT 848.100 344.400 849.900 351.000 ;
        RECT 851.100 344.400 852.900 350.400 ;
        RECT 845.100 342.600 850.800 343.500 ;
        RECT 849.000 341.700 850.800 342.600 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 818.550 332.550 822.450 333.450 ;
        RECT 827.250 333.150 829.050 334.950 ;
        RECT 821.550 330.450 822.450 332.550 ;
        RECT 829.950 330.450 832.050 330.750 ;
        RECT 821.550 329.550 832.050 330.450 ;
        RECT 829.950 328.650 832.050 329.550 ;
        RECT 833.700 327.600 834.600 334.950 ;
        RECT 835.950 333.450 838.050 334.050 ;
        RECT 841.950 333.450 844.050 337.050 ;
        RECT 835.950 333.000 844.050 333.450 ;
        RECT 845.400 334.950 847.500 337.050 ;
        RECT 845.400 333.150 847.200 334.950 ;
        RECT 835.950 332.550 843.450 333.000 ;
        RECT 835.950 331.950 838.050 332.550 ;
        RECT 849.000 330.300 849.900 341.700 ;
        RECT 851.700 337.050 852.900 344.400 ;
        RECT 863.100 347.400 864.900 350.400 ;
        RECT 863.100 343.500 864.300 347.400 ;
        RECT 866.100 344.400 867.900 351.000 ;
        RECT 869.100 344.400 870.900 350.400 ;
        RECT 863.100 342.600 868.800 343.500 ;
        RECT 867.000 341.700 868.800 342.600 ;
        RECT 850.800 334.950 852.900 337.050 ;
        RECT 849.000 329.400 850.800 330.300 ;
        RECT 845.100 328.500 850.800 329.400 ;
        RECT 806.400 321.900 813.000 322.800 ;
        RECT 806.400 321.600 807.900 321.900 ;
        RECT 785.100 315.000 786.900 321.600 ;
        RECT 788.100 315.600 789.900 321.600 ;
        RECT 791.100 315.000 792.900 321.600 ;
        RECT 803.100 315.000 804.900 321.600 ;
        RECT 806.100 315.600 807.900 321.600 ;
        RECT 812.100 321.600 813.000 321.900 ;
        RECT 824.100 326.700 831.900 327.600 ;
        RECT 809.100 315.000 810.900 321.000 ;
        RECT 812.100 315.600 813.900 321.600 ;
        RECT 824.100 315.600 825.900 326.700 ;
        RECT 827.100 315.000 828.900 325.800 ;
        RECT 830.100 315.600 831.900 326.700 ;
        RECT 833.100 315.600 834.900 327.600 ;
        RECT 845.100 321.600 846.300 328.500 ;
        RECT 851.700 327.600 852.900 334.950 ;
        RECT 863.400 334.950 865.500 337.050 ;
        RECT 863.400 333.150 865.200 334.950 ;
        RECT 853.950 328.950 856.050 331.050 ;
        RECT 867.000 330.300 867.900 341.700 ;
        RECT 869.700 337.050 870.900 344.400 ;
        RECT 868.800 334.950 870.900 337.050 ;
        RECT 867.000 329.400 868.800 330.300 ;
        RECT 845.100 315.600 846.900 321.600 ;
        RECT 848.100 315.000 849.900 325.800 ;
        RECT 851.100 315.600 852.900 327.600 ;
        RECT 854.550 325.050 855.450 328.950 ;
        RECT 863.100 328.500 868.800 329.400 ;
        RECT 853.950 322.950 856.050 325.050 ;
        RECT 863.100 321.600 864.300 328.500 ;
        RECT 869.700 327.600 870.900 334.950 ;
        RECT 863.100 315.600 864.900 321.600 ;
        RECT 866.100 315.000 867.900 325.800 ;
        RECT 869.100 315.600 870.900 327.600 ;
        RECT 11.100 300.300 12.900 311.400 ;
        RECT 14.100 301.200 15.900 312.000 ;
        RECT 17.100 300.300 18.900 311.400 ;
        RECT 11.100 299.400 18.900 300.300 ;
        RECT 20.100 299.400 21.900 311.400 ;
        RECT 32.100 305.400 33.900 312.000 ;
        RECT 35.100 305.400 36.900 311.400 ;
        RECT 38.100 306.000 39.900 312.000 ;
        RECT 35.400 305.100 36.900 305.400 ;
        RECT 41.100 305.400 42.900 311.400 ;
        RECT 56.100 305.400 57.900 311.400 ;
        RECT 59.100 305.400 60.900 312.000 ;
        RECT 71.100 305.400 72.900 311.400 ;
        RECT 74.100 305.400 75.900 312.000 ;
        RECT 86.100 305.400 87.900 312.000 ;
        RECT 89.100 305.400 90.900 311.400 ;
        RECT 92.100 306.000 93.900 312.000 ;
        RECT 41.100 305.100 42.000 305.400 ;
        RECT 35.400 304.200 42.000 305.100 ;
        RECT 14.250 292.050 16.050 293.850 ;
        RECT 20.700 292.050 21.600 299.400 ;
        RECT 25.950 297.450 28.050 298.050 ;
        RECT 37.950 297.450 40.050 298.050 ;
        RECT 25.950 296.550 40.050 297.450 ;
        RECT 25.950 295.950 28.050 296.550 ;
        RECT 37.950 295.950 40.050 296.550 ;
        RECT 35.100 292.050 36.900 293.850 ;
        RECT 41.100 292.050 42.000 304.200 ;
        RECT 56.700 292.050 57.900 305.400 ;
        RECT 59.100 292.050 60.900 293.850 ;
        RECT 71.700 292.050 72.900 305.400 ;
        RECT 89.400 305.100 90.900 305.400 ;
        RECT 95.100 305.400 96.900 311.400 ;
        RECT 107.100 305.400 108.900 312.000 ;
        RECT 110.100 305.400 111.900 311.400 ;
        RECT 113.100 306.000 114.900 312.000 ;
        RECT 95.100 305.100 96.000 305.400 ;
        RECT 89.400 304.200 96.000 305.100 ;
        RECT 110.400 305.100 111.900 305.400 ;
        RECT 116.100 305.400 117.900 311.400 ;
        RECT 128.100 305.400 129.900 312.000 ;
        RECT 131.100 305.400 132.900 311.400 ;
        RECT 134.100 306.000 135.900 312.000 ;
        RECT 116.100 305.100 117.000 305.400 ;
        RECT 110.400 304.200 117.000 305.100 ;
        RECT 131.400 305.100 132.900 305.400 ;
        RECT 137.100 305.400 138.900 311.400 ;
        RECT 137.100 305.100 138.000 305.400 ;
        RECT 131.400 304.200 138.000 305.100 ;
        RECT 74.100 292.050 75.900 293.850 ;
        RECT 89.100 292.050 90.900 293.850 ;
        RECT 95.100 292.050 96.000 304.200 ;
        RECT 102.000 294.450 106.050 295.050 ;
        RECT 101.550 292.950 106.050 294.450 ;
        RECT 10.950 289.950 13.050 292.050 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 31.950 289.950 34.050 292.050 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 70.950 289.950 73.050 292.050 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 88.950 289.950 91.050 292.050 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 94.950 289.950 97.050 292.050 ;
        RECT 11.100 288.150 12.900 289.950 ;
        RECT 17.250 288.150 19.050 289.950 ;
        RECT 20.700 282.600 21.600 289.950 ;
        RECT 32.100 288.150 33.900 289.950 ;
        RECT 38.100 288.150 39.900 289.950 ;
        RECT 41.100 286.200 42.000 289.950 ;
        RECT 12.000 276.000 13.800 282.600 ;
        RECT 16.500 281.400 21.600 282.600 ;
        RECT 16.500 276.600 18.300 281.400 ;
        RECT 19.500 276.000 21.300 279.600 ;
        RECT 32.100 276.000 33.900 285.600 ;
        RECT 38.700 285.000 42.000 286.200 ;
        RECT 38.700 276.600 40.500 285.000 ;
        RECT 56.700 279.600 57.900 289.950 ;
        RECT 71.700 279.600 72.900 289.950 ;
        RECT 86.100 288.150 87.900 289.950 ;
        RECT 92.100 288.150 93.900 289.950 ;
        RECT 95.100 286.200 96.000 289.950 ;
        RECT 101.550 289.050 102.450 292.950 ;
        RECT 110.100 292.050 111.900 293.850 ;
        RECT 116.100 292.050 117.000 304.200 ;
        RECT 131.100 292.050 132.900 293.850 ;
        RECT 137.100 292.050 138.000 304.200 ;
        RECT 149.100 299.400 150.900 311.400 ;
        RECT 152.100 300.300 153.900 311.400 ;
        RECT 155.100 301.200 156.900 312.000 ;
        RECT 158.100 300.300 159.900 311.400 ;
        RECT 152.100 299.400 159.900 300.300 ;
        RECT 171.000 300.600 172.800 311.400 ;
        RECT 171.000 299.400 174.600 300.600 ;
        RECT 176.100 299.400 177.900 312.000 ;
        RECT 188.400 299.400 190.200 312.000 ;
        RECT 193.500 300.900 195.300 311.400 ;
        RECT 196.500 305.400 198.300 312.000 ;
        RECT 209.100 305.400 210.900 311.400 ;
        RECT 212.100 306.000 213.900 312.000 ;
        RECT 210.000 305.100 210.900 305.400 ;
        RECT 215.100 305.400 216.900 311.400 ;
        RECT 218.100 305.400 219.900 312.000 ;
        RECT 230.100 305.400 231.900 312.000 ;
        RECT 233.100 305.400 234.900 311.400 ;
        RECT 236.100 305.400 237.900 312.000 ;
        RECT 215.100 305.100 216.600 305.400 ;
        RECT 210.000 304.200 216.600 305.100 ;
        RECT 196.200 302.100 198.000 303.900 ;
        RECT 193.500 299.400 195.900 300.900 ;
        RECT 149.400 292.050 150.300 299.400 ;
        RECT 160.950 294.450 165.000 295.050 ;
        RECT 154.950 292.050 156.750 293.850 ;
        RECT 160.950 292.950 165.450 294.450 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 112.950 289.950 115.050 292.050 ;
        RECT 115.950 289.950 118.050 292.050 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 136.950 289.950 139.050 292.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 157.950 289.950 160.050 292.050 ;
        RECT 97.950 287.550 102.450 289.050 ;
        RECT 107.100 288.150 108.900 289.950 ;
        RECT 113.100 288.150 114.900 289.950 ;
        RECT 97.950 286.950 102.000 287.550 ;
        RECT 116.100 286.200 117.000 289.950 ;
        RECT 128.100 288.150 129.900 289.950 ;
        RECT 134.100 288.150 135.900 289.950 ;
        RECT 137.100 286.200 138.000 289.950 ;
        RECT 56.100 276.600 57.900 279.600 ;
        RECT 59.100 276.000 60.900 279.600 ;
        RECT 71.100 276.600 72.900 279.600 ;
        RECT 74.100 276.000 75.900 279.600 ;
        RECT 86.100 276.000 87.900 285.600 ;
        RECT 92.700 285.000 96.000 286.200 ;
        RECT 92.700 276.600 94.500 285.000 ;
        RECT 107.100 276.000 108.900 285.600 ;
        RECT 113.700 285.000 117.000 286.200 ;
        RECT 113.700 276.600 115.500 285.000 ;
        RECT 128.100 276.000 129.900 285.600 ;
        RECT 134.700 285.000 138.000 286.200 ;
        RECT 134.700 276.600 136.500 285.000 ;
        RECT 149.400 282.600 150.300 289.950 ;
        RECT 151.950 288.150 153.750 289.950 ;
        RECT 158.100 288.150 159.900 289.950 ;
        RECT 164.550 289.050 165.450 292.950 ;
        RECT 170.100 292.050 171.900 293.850 ;
        RECT 173.700 292.050 174.600 299.400 ;
        RECT 175.950 292.050 177.750 293.850 ;
        RECT 188.100 292.050 189.900 293.850 ;
        RECT 194.700 292.050 195.900 299.400 ;
        RECT 199.950 294.450 204.000 295.050 ;
        RECT 199.950 292.950 204.450 294.450 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 164.550 287.550 169.050 289.050 ;
        RECT 165.000 286.950 169.050 287.550 ;
        RECT 149.400 281.400 154.500 282.600 ;
        RECT 149.700 276.000 151.500 279.600 ;
        RECT 152.700 276.600 154.500 281.400 ;
        RECT 157.200 276.000 159.000 282.600 ;
        RECT 173.700 279.600 174.600 289.950 ;
        RECT 191.100 288.150 192.900 289.950 ;
        RECT 194.700 285.600 195.900 289.950 ;
        RECT 197.100 288.150 198.900 289.950 ;
        RECT 203.550 289.050 204.450 292.950 ;
        RECT 210.000 292.050 210.900 304.200 ;
        RECT 214.950 297.450 217.050 298.050 ;
        RECT 214.950 296.550 222.450 297.450 ;
        RECT 214.950 295.950 217.050 296.550 ;
        RECT 221.550 294.450 222.450 296.550 ;
        RECT 215.100 292.050 216.900 293.850 ;
        RECT 221.550 293.550 225.450 294.450 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 203.550 287.550 208.050 289.050 ;
        RECT 204.000 286.950 208.050 287.550 ;
        RECT 210.000 286.200 210.900 289.950 ;
        RECT 212.100 288.150 213.900 289.950 ;
        RECT 218.100 288.150 219.900 289.950 ;
        RECT 224.550 289.050 225.450 293.550 ;
        RECT 233.100 292.050 234.300 305.400 ;
        RECT 248.100 300.600 249.900 311.400 ;
        RECT 251.100 301.500 252.900 312.000 ;
        RECT 254.100 310.500 261.900 311.400 ;
        RECT 254.100 300.600 255.900 310.500 ;
        RECT 248.100 299.700 255.900 300.600 ;
        RECT 257.100 298.500 258.900 309.600 ;
        RECT 260.100 299.400 261.900 310.500 ;
        RECT 272.100 305.400 273.900 312.000 ;
        RECT 275.100 305.400 276.900 311.400 ;
        RECT 254.100 297.600 258.900 298.500 ;
        RECT 243.000 294.450 247.050 295.050 ;
        RECT 242.550 292.950 247.050 294.450 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 220.950 287.550 225.450 289.050 ;
        RECT 230.250 288.150 232.050 289.950 ;
        RECT 220.950 286.950 225.000 287.550 ;
        RECT 194.700 284.700 198.300 285.600 ;
        RECT 210.000 285.000 213.300 286.200 ;
        RECT 188.100 281.700 195.900 283.050 ;
        RECT 170.100 276.000 171.900 279.600 ;
        RECT 173.100 276.600 174.900 279.600 ;
        RECT 176.100 276.000 177.900 279.600 ;
        RECT 188.100 276.600 189.900 281.700 ;
        RECT 191.100 276.000 192.900 280.800 ;
        RECT 194.100 276.600 195.900 281.700 ;
        RECT 197.100 282.600 198.300 284.700 ;
        RECT 197.100 276.600 198.900 282.600 ;
        RECT 211.500 276.600 213.300 285.000 ;
        RECT 218.100 276.000 219.900 285.600 ;
        RECT 233.100 284.700 234.300 289.950 ;
        RECT 236.100 288.150 237.900 289.950 ;
        RECT 242.550 289.050 243.450 292.950 ;
        RECT 251.250 292.050 253.050 293.850 ;
        RECT 254.100 292.050 255.000 297.600 ;
        RECT 262.950 294.450 267.000 295.050 ;
        RECT 257.100 292.050 258.900 293.850 ;
        RECT 262.950 292.950 267.450 294.450 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 250.950 289.950 253.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 242.550 287.550 247.050 289.050 ;
        RECT 248.250 288.150 250.050 289.950 ;
        RECT 243.000 286.950 247.050 287.550 ;
        RECT 233.100 283.800 237.300 284.700 ;
        RECT 230.400 276.000 232.200 282.600 ;
        RECT 235.500 276.600 237.300 283.800 ;
        RECT 254.100 282.600 255.300 289.950 ;
        RECT 260.100 288.150 261.900 289.950 ;
        RECT 266.550 285.450 267.450 292.950 ;
        RECT 272.100 292.050 273.900 293.850 ;
        RECT 275.100 292.050 276.300 305.400 ;
        RECT 287.400 299.400 289.200 312.000 ;
        RECT 292.500 300.900 294.300 311.400 ;
        RECT 295.500 305.400 297.300 312.000 ;
        RECT 295.200 302.100 297.000 303.900 ;
        RECT 292.500 299.400 294.900 300.900 ;
        RECT 280.950 297.450 283.050 298.050 ;
        RECT 289.950 297.450 292.050 298.050 ;
        RECT 280.950 296.550 292.050 297.450 ;
        RECT 280.950 295.950 283.050 296.550 ;
        RECT 289.950 295.950 292.050 296.550 ;
        RECT 282.000 294.450 286.050 295.050 ;
        RECT 281.550 292.950 286.050 294.450 ;
        RECT 271.950 289.950 274.050 292.050 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 271.950 285.450 274.050 285.750 ;
        RECT 266.550 284.550 274.050 285.450 ;
        RECT 271.950 283.650 274.050 284.550 ;
        RECT 248.700 276.000 250.500 282.600 ;
        RECT 253.200 276.600 255.000 282.600 ;
        RECT 257.700 276.000 259.500 282.600 ;
        RECT 275.100 279.600 276.300 289.950 ;
        RECT 281.550 289.050 282.450 292.950 ;
        RECT 287.100 292.050 288.900 293.850 ;
        RECT 293.700 292.050 294.900 299.400 ;
        RECT 311.100 299.400 312.900 311.400 ;
        RECT 314.100 301.200 315.900 312.000 ;
        RECT 317.100 305.400 318.900 311.400 ;
        RECT 329.100 305.400 330.900 312.000 ;
        RECT 332.100 305.400 333.900 311.400 ;
        RECT 335.100 305.400 336.900 312.000 ;
        RECT 347.700 305.400 349.500 312.000 ;
        RECT 311.100 292.050 312.300 299.400 ;
        RECT 317.700 298.500 318.900 305.400 ;
        RECT 313.200 297.600 318.900 298.500 ;
        RECT 313.200 296.700 315.000 297.600 ;
        RECT 286.950 289.950 289.050 292.050 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 311.100 289.950 313.200 292.050 ;
        RECT 281.550 287.550 286.050 289.050 ;
        RECT 290.100 288.150 291.900 289.950 ;
        RECT 282.000 286.950 286.050 287.550 ;
        RECT 293.700 285.600 294.900 289.950 ;
        RECT 296.100 288.150 297.900 289.950 ;
        RECT 293.700 284.700 297.300 285.600 ;
        RECT 287.100 281.700 294.900 283.050 ;
        RECT 272.100 276.000 273.900 279.600 ;
        RECT 275.100 276.600 276.900 279.600 ;
        RECT 287.100 276.600 288.900 281.700 ;
        RECT 290.100 276.000 291.900 280.800 ;
        RECT 293.100 276.600 294.900 281.700 ;
        RECT 296.100 282.600 297.300 284.700 ;
        RECT 311.100 282.600 312.300 289.950 ;
        RECT 314.100 285.300 315.000 296.700 ;
        RECT 316.800 292.050 318.600 293.850 ;
        RECT 332.700 292.050 333.900 305.400 ;
        RECT 348.000 302.100 349.800 303.900 ;
        RECT 350.700 300.900 352.500 311.400 ;
        RECT 350.100 299.400 352.500 300.900 ;
        RECT 355.800 299.400 357.600 312.000 ;
        RECT 368.100 305.400 369.900 312.000 ;
        RECT 371.100 305.400 372.900 311.400 ;
        RECT 374.100 305.400 375.900 312.000 ;
        RECT 350.100 292.050 351.300 299.400 ;
        RECT 356.100 292.050 357.900 293.850 ;
        RECT 371.100 292.050 372.300 305.400 ;
        RECT 386.400 299.400 388.200 312.000 ;
        RECT 391.500 300.900 393.300 311.400 ;
        RECT 394.500 305.400 396.300 312.000 ;
        RECT 410.100 305.400 411.900 312.000 ;
        RECT 413.100 305.400 414.900 311.400 ;
        RECT 416.100 305.400 417.900 312.000 ;
        RECT 394.200 302.100 396.000 303.900 ;
        RECT 391.500 299.400 393.900 300.900 ;
        RECT 386.100 292.050 387.900 293.850 ;
        RECT 392.700 292.050 393.900 299.400 ;
        RECT 413.100 292.050 414.300 305.400 ;
        RECT 431.100 299.400 432.900 311.400 ;
        RECT 434.100 299.400 435.900 312.000 ;
        RECT 449.100 305.400 450.900 312.000 ;
        RECT 452.100 305.400 453.900 311.400 ;
        RECT 455.100 305.400 456.900 312.000 ;
        RECT 431.700 292.050 432.900 299.400 ;
        RECT 452.100 292.050 453.300 305.400 ;
        RECT 467.400 299.400 469.200 312.000 ;
        RECT 472.500 300.900 474.300 311.400 ;
        RECT 475.500 305.400 477.300 312.000 ;
        RECT 475.200 302.100 477.000 303.900 ;
        RECT 480.150 301.200 481.950 311.400 ;
        RECT 472.500 299.400 474.900 300.900 ;
        RECT 467.100 292.050 468.900 293.850 ;
        RECT 473.700 292.050 474.900 299.400 ;
        RECT 479.550 299.400 481.950 301.200 ;
        RECT 483.150 299.400 484.950 312.000 ;
        RECT 488.550 302.400 490.350 311.400 ;
        RECT 493.350 305.400 495.150 312.000 ;
        RECT 496.350 304.500 498.150 311.400 ;
        RECT 499.350 305.400 501.150 312.000 ;
        RECT 503.850 305.400 505.650 311.400 ;
        RECT 492.450 303.450 499.050 304.500 ;
        RECT 492.450 302.700 494.250 303.450 ;
        RECT 497.250 302.700 499.050 303.450 ;
        RECT 503.550 303.300 505.650 305.400 ;
        RECT 488.250 301.500 490.350 302.400 ;
        RECT 500.850 301.800 502.650 302.400 ;
        RECT 488.250 300.300 496.050 301.500 ;
        RECT 494.250 299.700 496.050 300.300 ;
        RECT 496.950 300.900 502.650 301.800 ;
        RECT 479.550 298.500 480.450 299.400 ;
        RECT 496.950 298.800 497.850 300.900 ;
        RECT 500.850 300.600 502.650 300.900 ;
        RECT 503.550 300.600 506.550 302.400 ;
        RECT 503.550 299.700 504.750 300.600 ;
        RECT 489.450 298.500 497.850 298.800 ;
        RECT 479.550 297.900 497.850 298.500 ;
        RECT 499.950 298.800 504.750 299.700 ;
        RECT 508.650 299.400 510.450 312.000 ;
        RECT 511.650 299.400 513.450 311.400 ;
        RECT 524.100 305.400 525.900 312.000 ;
        RECT 527.100 305.400 528.900 311.400 ;
        RECT 479.550 297.300 491.250 297.900 ;
        RECT 316.500 289.950 318.600 292.050 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 346.950 289.950 349.050 292.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 352.950 289.950 355.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 367.950 289.950 370.050 292.050 ;
        RECT 370.950 289.950 373.050 292.050 ;
        RECT 373.950 289.950 376.050 292.050 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 388.950 289.950 391.050 292.050 ;
        RECT 391.950 289.950 394.050 292.050 ;
        RECT 394.950 289.950 397.050 292.050 ;
        RECT 409.950 289.950 412.050 292.050 ;
        RECT 412.950 289.950 415.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 430.950 289.950 433.050 292.050 ;
        RECT 433.950 289.950 436.050 292.050 ;
        RECT 448.950 289.950 451.050 292.050 ;
        RECT 451.950 289.950 454.050 292.050 ;
        RECT 454.950 289.950 457.050 292.050 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 472.950 289.950 475.050 292.050 ;
        RECT 475.950 289.950 478.050 292.050 ;
        RECT 329.100 288.150 330.900 289.950 ;
        RECT 313.200 284.400 315.000 285.300 ;
        RECT 332.700 284.700 333.900 289.950 ;
        RECT 334.950 288.150 336.750 289.950 ;
        RECT 347.100 288.150 348.900 289.950 ;
        RECT 350.100 285.600 351.300 289.950 ;
        RECT 353.100 288.150 354.900 289.950 ;
        RECT 368.250 288.150 370.050 289.950 ;
        RECT 313.200 283.500 318.900 284.400 ;
        RECT 296.100 276.600 297.900 282.600 ;
        RECT 311.100 276.600 312.900 282.600 ;
        RECT 314.100 276.000 315.900 282.600 ;
        RECT 317.700 279.600 318.900 283.500 ;
        RECT 317.100 276.600 318.900 279.600 ;
        RECT 329.700 283.800 333.900 284.700 ;
        RECT 347.700 284.700 351.300 285.600 ;
        RECT 371.100 284.700 372.300 289.950 ;
        RECT 374.100 288.150 375.900 289.950 ;
        RECT 389.100 288.150 390.900 289.950 ;
        RECT 392.700 285.600 393.900 289.950 ;
        RECT 395.100 288.150 396.900 289.950 ;
        RECT 410.250 288.150 412.050 289.950 ;
        RECT 392.700 284.700 396.300 285.600 ;
        RECT 329.700 276.600 331.500 283.800 ;
        RECT 347.700 282.600 348.900 284.700 ;
        RECT 371.100 283.800 375.300 284.700 ;
        RECT 334.800 276.000 336.600 282.600 ;
        RECT 347.100 276.600 348.900 282.600 ;
        RECT 350.100 281.700 357.900 283.050 ;
        RECT 350.100 276.600 351.900 281.700 ;
        RECT 353.100 276.000 354.900 280.800 ;
        RECT 356.100 276.600 357.900 281.700 ;
        RECT 368.400 276.000 370.200 282.600 ;
        RECT 373.500 276.600 375.300 283.800 ;
        RECT 386.100 281.700 393.900 283.050 ;
        RECT 386.100 276.600 387.900 281.700 ;
        RECT 389.100 276.000 390.900 280.800 ;
        RECT 392.100 276.600 393.900 281.700 ;
        RECT 395.100 282.600 396.300 284.700 ;
        RECT 413.100 284.700 414.300 289.950 ;
        RECT 416.100 288.150 417.900 289.950 ;
        RECT 413.100 283.800 417.300 284.700 ;
        RECT 395.100 276.600 396.900 282.600 ;
        RECT 410.400 276.000 412.200 282.600 ;
        RECT 415.500 276.600 417.300 283.800 ;
        RECT 431.700 282.600 432.900 289.950 ;
        RECT 434.100 288.150 435.900 289.950 ;
        RECT 449.250 288.150 451.050 289.950 ;
        RECT 452.100 284.700 453.300 289.950 ;
        RECT 455.100 288.150 456.900 289.950 ;
        RECT 470.100 288.150 471.900 289.950 ;
        RECT 473.700 285.600 474.900 289.950 ;
        RECT 476.100 288.150 477.900 289.950 ;
        RECT 473.700 284.700 477.300 285.600 ;
        RECT 452.100 283.800 456.300 284.700 ;
        RECT 431.100 276.600 432.900 282.600 ;
        RECT 434.100 276.000 435.900 282.600 ;
        RECT 449.400 276.000 451.200 282.600 ;
        RECT 454.500 276.600 456.300 283.800 ;
        RECT 467.100 281.700 474.900 283.050 ;
        RECT 467.100 276.600 468.900 281.700 ;
        RECT 470.100 276.000 471.900 280.800 ;
        RECT 473.100 276.600 474.900 281.700 ;
        RECT 476.100 282.600 477.300 284.700 ;
        RECT 479.550 282.600 480.450 297.300 ;
        RECT 489.450 297.000 491.250 297.300 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 491.100 290.400 493.200 292.050 ;
        RECT 481.950 287.400 483.750 289.950 ;
        RECT 485.100 289.200 493.200 290.400 ;
        RECT 485.100 288.600 486.900 289.200 ;
        RECT 488.100 287.400 489.900 288.000 ;
        RECT 481.950 286.200 489.900 287.400 ;
        RECT 499.950 286.200 500.850 298.800 ;
        RECT 503.550 296.100 505.650 296.700 ;
        RECT 509.550 296.100 511.350 296.550 ;
        RECT 503.550 294.900 511.350 296.100 ;
        RECT 503.550 294.600 505.650 294.900 ;
        RECT 509.550 294.750 511.350 294.900 ;
        RECT 512.250 292.050 513.450 299.400 ;
        RECT 508.950 291.750 513.450 292.050 ;
        RECT 507.150 289.950 513.450 291.750 ;
        RECT 524.100 289.950 526.200 292.050 ;
        RECT 488.850 285.000 500.850 286.200 ;
        RECT 488.850 283.200 489.900 285.000 ;
        RECT 499.050 284.400 500.850 285.000 ;
        RECT 476.100 276.600 477.900 282.600 ;
        RECT 479.550 280.800 481.950 282.600 ;
        RECT 480.150 276.600 481.950 280.800 ;
        RECT 483.150 276.000 484.950 282.600 ;
        RECT 485.850 280.200 487.950 281.700 ;
        RECT 488.850 281.400 490.650 283.200 ;
        RECT 512.250 282.600 513.450 289.950 ;
        RECT 524.250 288.150 526.050 289.950 ;
        RECT 527.100 285.300 528.000 305.400 ;
        RECT 530.100 300.000 531.900 312.000 ;
        RECT 533.100 299.400 534.900 311.400 ;
        RECT 545.400 299.400 547.200 312.000 ;
        RECT 550.500 300.900 552.300 311.400 ;
        RECT 553.500 305.400 555.300 312.000 ;
        RECT 566.100 305.400 567.900 312.000 ;
        RECT 569.100 305.400 570.900 311.400 ;
        RECT 553.200 302.100 555.000 303.900 ;
        RECT 550.500 299.400 552.900 300.900 ;
        RECT 529.200 292.050 531.000 293.850 ;
        RECT 533.400 292.050 534.300 299.400 ;
        RECT 544.950 297.450 547.050 298.050 ;
        RECT 536.550 296.550 547.050 297.450 ;
        RECT 529.500 289.950 531.600 292.050 ;
        RECT 532.800 289.950 534.900 292.050 ;
        RECT 491.850 281.550 493.650 282.300 ;
        RECT 491.850 280.500 496.800 281.550 ;
        RECT 485.850 279.600 489.750 280.200 ;
        RECT 495.750 279.600 496.800 280.500 ;
        RECT 503.250 279.600 505.650 281.700 ;
        RECT 486.150 278.700 489.750 279.600 ;
        RECT 487.950 276.600 489.750 278.700 ;
        RECT 492.450 276.000 494.250 279.600 ;
        RECT 495.750 276.600 497.550 279.600 ;
        RECT 498.750 276.000 500.550 279.600 ;
        RECT 503.250 276.600 505.050 279.600 ;
        RECT 508.350 276.000 510.150 282.600 ;
        RECT 511.650 276.600 513.450 282.600 ;
        RECT 524.100 284.400 532.500 285.300 ;
        RECT 524.100 276.600 525.900 284.400 ;
        RECT 530.700 283.500 532.500 284.400 ;
        RECT 533.400 282.600 534.300 289.950 ;
        RECT 528.600 276.000 530.400 282.600 ;
        RECT 531.600 280.800 534.300 282.600 ;
        RECT 531.600 276.600 533.400 280.800 ;
        RECT 536.550 280.050 537.450 296.550 ;
        RECT 544.950 295.950 547.050 296.550 ;
        RECT 540.000 294.450 544.050 295.050 ;
        RECT 539.550 292.950 544.050 294.450 ;
        RECT 539.550 283.050 540.450 292.950 ;
        RECT 545.100 292.050 546.900 293.850 ;
        RECT 551.700 292.050 552.900 299.400 ;
        RECT 556.950 294.450 561.000 295.050 ;
        RECT 556.950 292.950 561.450 294.450 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 548.100 288.150 549.900 289.950 ;
        RECT 551.700 285.600 552.900 289.950 ;
        RECT 554.100 288.150 555.900 289.950 ;
        RECT 560.550 289.050 561.450 292.950 ;
        RECT 566.100 289.950 568.200 292.050 ;
        RECT 556.950 287.550 561.450 289.050 ;
        RECT 566.250 288.150 568.050 289.950 ;
        RECT 556.950 286.950 561.000 287.550 ;
        RECT 551.700 284.700 555.300 285.600 ;
        RECT 569.100 285.300 570.000 305.400 ;
        RECT 572.100 300.000 573.900 312.000 ;
        RECT 575.100 299.400 576.900 311.400 ;
        RECT 587.100 305.400 588.900 312.000 ;
        RECT 590.100 305.400 591.900 311.400 ;
        RECT 593.100 305.400 594.900 312.000 ;
        RECT 608.100 305.400 609.900 312.000 ;
        RECT 611.100 305.400 612.900 311.400 ;
        RECT 614.100 305.400 615.900 312.000 ;
        RECT 626.100 305.400 627.900 312.000 ;
        RECT 629.100 305.400 630.900 311.400 ;
        RECT 632.100 305.400 633.900 312.000 ;
        RECT 571.200 292.050 573.000 293.850 ;
        RECT 575.400 292.050 576.300 299.400 ;
        RECT 582.000 294.450 586.050 295.050 ;
        RECT 581.550 292.950 586.050 294.450 ;
        RECT 571.500 289.950 573.600 292.050 ;
        RECT 574.800 289.950 576.900 292.050 ;
        RECT 538.950 280.950 541.050 283.050 ;
        RECT 545.100 281.700 552.900 283.050 ;
        RECT 535.950 277.950 538.050 280.050 ;
        RECT 545.100 276.600 546.900 281.700 ;
        RECT 548.100 276.000 549.900 280.800 ;
        RECT 551.100 276.600 552.900 281.700 ;
        RECT 554.100 282.600 555.300 284.700 ;
        RECT 566.100 284.400 574.500 285.300 ;
        RECT 554.100 276.600 555.900 282.600 ;
        RECT 566.100 276.600 567.900 284.400 ;
        RECT 572.700 283.500 574.500 284.400 ;
        RECT 575.400 282.600 576.300 289.950 ;
        RECT 570.600 276.000 572.400 282.600 ;
        RECT 573.600 280.800 576.300 282.600 ;
        RECT 581.550 283.050 582.450 292.950 ;
        RECT 590.100 292.050 591.300 305.400 ;
        RECT 611.100 292.050 612.300 305.400 ;
        RECT 621.000 294.450 625.050 295.050 ;
        RECT 620.550 292.950 625.050 294.450 ;
        RECT 586.950 289.950 589.050 292.050 ;
        RECT 589.950 289.950 592.050 292.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 610.950 289.950 613.050 292.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 587.250 288.150 589.050 289.950 ;
        RECT 590.100 284.700 591.300 289.950 ;
        RECT 593.100 288.150 594.900 289.950 ;
        RECT 608.250 288.150 610.050 289.950 ;
        RECT 611.100 284.700 612.300 289.950 ;
        RECT 614.100 288.150 615.900 289.950 ;
        RECT 620.550 285.450 621.450 292.950 ;
        RECT 629.100 292.050 630.300 305.400 ;
        RECT 644.100 299.400 645.900 312.000 ;
        RECT 647.100 299.400 648.900 311.400 ;
        RECT 662.400 299.400 664.200 312.000 ;
        RECT 667.500 300.900 669.300 311.400 ;
        RECT 670.500 305.400 672.300 312.000 ;
        RECT 683.100 305.400 684.900 312.000 ;
        RECT 686.100 305.400 687.900 311.400 ;
        RECT 689.100 305.400 690.900 312.000 ;
        RECT 670.200 302.100 672.000 303.900 ;
        RECT 667.500 299.400 669.900 300.900 ;
        RECT 639.000 294.450 643.050 295.050 ;
        RECT 638.550 292.950 643.050 294.450 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 626.250 288.150 628.050 289.950 ;
        RECT 625.950 285.450 628.050 286.050 ;
        RECT 590.100 283.800 594.300 284.700 ;
        RECT 611.100 283.800 615.300 284.700 ;
        RECT 620.550 284.550 628.050 285.450 ;
        RECT 625.950 283.950 628.050 284.550 ;
        RECT 629.100 284.700 630.300 289.950 ;
        RECT 632.100 288.150 633.900 289.950 ;
        RECT 638.550 289.050 639.450 292.950 ;
        RECT 647.100 292.050 648.300 299.400 ;
        RECT 662.100 292.050 663.900 293.850 ;
        RECT 668.700 292.050 669.900 299.400 ;
        RECT 686.700 292.050 687.900 305.400 ;
        RECT 688.950 303.450 691.050 304.050 ;
        RECT 694.950 303.450 697.050 304.050 ;
        RECT 688.950 302.550 697.050 303.450 ;
        RECT 688.950 301.950 691.050 302.550 ;
        RECT 694.950 301.950 697.050 302.550 ;
        RECT 701.100 300.300 702.900 311.400 ;
        RECT 704.100 301.200 705.900 312.000 ;
        RECT 707.100 300.300 708.900 311.400 ;
        RECT 701.100 299.400 708.900 300.300 ;
        RECT 710.100 299.400 711.900 311.400 ;
        RECT 722.100 305.400 723.900 312.000 ;
        RECT 725.100 305.400 726.900 311.400 ;
        RECT 728.100 306.000 729.900 312.000 ;
        RECT 725.400 305.100 726.900 305.400 ;
        RECT 731.100 305.400 732.900 311.400 ;
        RECT 746.100 305.400 747.900 312.000 ;
        RECT 749.100 305.400 750.900 311.400 ;
        RECT 731.100 305.100 732.000 305.400 ;
        RECT 725.400 304.200 732.000 305.100 ;
        RECT 688.950 297.450 691.050 298.050 ;
        RECT 703.950 297.450 706.050 298.050 ;
        RECT 688.950 296.550 706.050 297.450 ;
        RECT 688.950 295.950 691.050 296.550 ;
        RECT 703.950 295.950 706.050 296.550 ;
        RECT 704.250 292.050 706.050 293.850 ;
        RECT 710.700 292.050 711.600 299.400 ;
        RECT 712.950 294.450 717.000 295.050 ;
        RECT 712.950 292.950 717.450 294.450 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 646.950 289.950 649.050 292.050 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 667.950 289.950 670.050 292.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 703.950 289.950 706.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 634.950 287.550 639.450 289.050 ;
        RECT 644.100 288.150 645.900 289.950 ;
        RECT 634.950 286.950 639.000 287.550 ;
        RECT 629.100 283.800 633.300 284.700 ;
        RECT 581.550 281.550 586.050 283.050 ;
        RECT 582.000 280.950 586.050 281.550 ;
        RECT 573.600 276.600 575.400 280.800 ;
        RECT 587.400 276.000 589.200 282.600 ;
        RECT 592.500 276.600 594.300 283.800 ;
        RECT 608.400 276.000 610.200 282.600 ;
        RECT 613.500 276.600 615.300 283.800 ;
        RECT 626.400 276.000 628.200 282.600 ;
        RECT 631.500 276.600 633.300 283.800 ;
        RECT 647.100 282.600 648.300 289.950 ;
        RECT 665.100 288.150 666.900 289.950 ;
        RECT 668.700 285.600 669.900 289.950 ;
        RECT 671.100 288.150 672.900 289.950 ;
        RECT 683.100 288.150 684.900 289.950 ;
        RECT 668.700 284.700 672.300 285.600 ;
        RECT 686.700 284.700 687.900 289.950 ;
        RECT 688.950 288.150 690.750 289.950 ;
        RECT 701.100 288.150 702.900 289.950 ;
        RECT 707.250 288.150 709.050 289.950 ;
        RECT 644.100 276.000 645.900 282.600 ;
        RECT 647.100 276.600 648.900 282.600 ;
        RECT 662.100 281.700 669.900 283.050 ;
        RECT 662.100 276.600 663.900 281.700 ;
        RECT 665.100 276.000 666.900 280.800 ;
        RECT 668.100 276.600 669.900 281.700 ;
        RECT 671.100 282.600 672.300 284.700 ;
        RECT 683.700 283.800 687.900 284.700 ;
        RECT 671.100 276.600 672.900 282.600 ;
        RECT 683.700 276.600 685.500 283.800 ;
        RECT 710.700 282.600 711.600 289.950 ;
        RECT 716.550 289.050 717.450 292.950 ;
        RECT 725.100 292.050 726.900 293.850 ;
        RECT 731.100 292.050 732.000 304.200 ;
        RECT 746.100 292.050 747.900 293.850 ;
        RECT 749.100 292.050 750.300 305.400 ;
        RECT 761.400 299.400 763.200 312.000 ;
        RECT 766.500 300.900 768.300 311.400 ;
        RECT 769.500 305.400 771.300 312.000 ;
        RECT 769.200 302.100 771.000 303.900 ;
        RECT 766.500 299.400 768.900 300.900 ;
        RECT 782.400 299.400 784.200 312.000 ;
        RECT 787.500 300.900 789.300 311.400 ;
        RECT 790.500 305.400 792.300 312.000 ;
        RECT 803.100 305.400 804.900 312.000 ;
        RECT 806.100 305.400 807.900 311.400 ;
        RECT 809.100 306.000 810.900 312.000 ;
        RECT 806.400 305.100 807.900 305.400 ;
        RECT 812.100 305.400 813.900 311.400 ;
        RECT 824.100 305.400 825.900 311.400 ;
        RECT 827.100 306.000 828.900 312.000 ;
        RECT 812.100 305.100 813.000 305.400 ;
        RECT 806.400 304.200 813.000 305.100 ;
        RECT 790.200 302.100 792.000 303.900 ;
        RECT 787.500 299.400 789.900 300.900 ;
        RECT 751.950 294.450 756.000 295.050 ;
        RECT 751.950 292.950 756.450 294.450 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 727.950 289.950 730.050 292.050 ;
        RECT 730.950 289.950 733.050 292.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 748.950 289.950 751.050 292.050 ;
        RECT 716.550 287.550 721.050 289.050 ;
        RECT 722.100 288.150 723.900 289.950 ;
        RECT 728.100 288.150 729.900 289.950 ;
        RECT 717.000 286.950 721.050 287.550 ;
        RECT 731.100 286.200 732.000 289.950 ;
        RECT 688.800 276.000 690.600 282.600 ;
        RECT 702.000 276.000 703.800 282.600 ;
        RECT 706.500 281.400 711.600 282.600 ;
        RECT 706.500 276.600 708.300 281.400 ;
        RECT 709.500 276.000 711.300 279.600 ;
        RECT 722.100 276.000 723.900 285.600 ;
        RECT 728.700 285.000 732.000 286.200 ;
        RECT 728.700 276.600 730.500 285.000 ;
        RECT 739.950 282.450 742.050 283.050 ;
        RECT 745.950 282.450 748.050 283.050 ;
        RECT 739.950 281.550 748.050 282.450 ;
        RECT 739.950 280.950 742.050 281.550 ;
        RECT 745.950 280.950 748.050 281.550 ;
        RECT 749.100 279.600 750.300 289.950 ;
        RECT 755.550 289.050 756.450 292.950 ;
        RECT 761.100 292.050 762.900 293.850 ;
        RECT 767.700 292.050 768.900 299.400 ;
        RECT 782.100 292.050 783.900 293.850 ;
        RECT 788.700 292.050 789.900 299.400 ;
        RECT 796.950 297.450 799.050 298.050 ;
        RECT 808.950 297.450 811.050 298.050 ;
        RECT 796.950 296.550 811.050 297.450 ;
        RECT 796.950 295.950 799.050 296.550 ;
        RECT 808.950 295.950 811.050 296.550 ;
        RECT 793.950 294.450 798.000 295.050 ;
        RECT 793.950 292.950 798.450 294.450 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 769.950 289.950 772.050 292.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 790.950 289.950 793.050 292.050 ;
        RECT 755.550 287.550 760.050 289.050 ;
        RECT 764.100 288.150 765.900 289.950 ;
        RECT 756.000 286.950 760.050 287.550 ;
        RECT 767.700 285.600 768.900 289.950 ;
        RECT 770.100 288.150 771.900 289.950 ;
        RECT 785.100 288.150 786.900 289.950 ;
        RECT 788.700 285.600 789.900 289.950 ;
        RECT 791.100 288.150 792.900 289.950 ;
        RECT 797.550 289.050 798.450 292.950 ;
        RECT 806.100 292.050 807.900 293.850 ;
        RECT 812.100 292.050 813.000 304.200 ;
        RECT 825.000 305.100 825.900 305.400 ;
        RECT 830.100 305.400 831.900 311.400 ;
        RECT 833.100 305.400 834.900 312.000 ;
        RECT 830.100 305.100 831.600 305.400 ;
        RECT 825.000 304.200 831.600 305.100 ;
        RECT 825.000 292.050 825.900 304.200 ;
        RECT 845.100 299.400 846.900 311.400 ;
        RECT 848.100 300.000 849.900 312.000 ;
        RECT 851.100 305.400 852.900 311.400 ;
        RECT 854.100 305.400 855.900 312.000 ;
        RECT 830.100 292.050 831.900 293.850 ;
        RECT 845.700 292.050 846.600 299.400 ;
        RECT 849.000 292.050 850.800 293.850 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 805.950 289.950 808.050 292.050 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 823.950 289.950 826.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 845.100 289.950 847.200 292.050 ;
        RECT 848.400 289.950 850.500 292.050 ;
        RECT 793.950 287.550 798.450 289.050 ;
        RECT 803.100 288.150 804.900 289.950 ;
        RECT 809.100 288.150 810.900 289.950 ;
        RECT 793.950 286.950 798.000 287.550 ;
        RECT 812.100 286.200 813.000 289.950 ;
        RECT 767.700 284.700 771.300 285.600 ;
        RECT 788.700 284.700 792.300 285.600 ;
        RECT 761.100 281.700 768.900 283.050 ;
        RECT 746.100 276.000 747.900 279.600 ;
        RECT 749.100 276.600 750.900 279.600 ;
        RECT 761.100 276.600 762.900 281.700 ;
        RECT 764.100 276.000 765.900 280.800 ;
        RECT 767.100 276.600 768.900 281.700 ;
        RECT 770.100 282.600 771.300 284.700 ;
        RECT 770.100 276.600 771.900 282.600 ;
        RECT 782.100 281.700 789.900 283.050 ;
        RECT 782.100 276.600 783.900 281.700 ;
        RECT 785.100 276.000 786.900 280.800 ;
        RECT 788.100 276.600 789.900 281.700 ;
        RECT 791.100 282.600 792.300 284.700 ;
        RECT 791.100 276.600 792.900 282.600 ;
        RECT 803.100 276.000 804.900 285.600 ;
        RECT 809.700 285.000 813.000 286.200 ;
        RECT 825.000 286.200 825.900 289.950 ;
        RECT 827.100 288.150 828.900 289.950 ;
        RECT 833.100 288.150 834.900 289.950 ;
        RECT 825.000 285.000 828.300 286.200 ;
        RECT 809.700 276.600 811.500 285.000 ;
        RECT 826.500 276.600 828.300 285.000 ;
        RECT 833.100 276.000 834.900 285.600 ;
        RECT 845.700 282.600 846.600 289.950 ;
        RECT 852.000 285.300 852.900 305.400 ;
        RECT 862.950 297.450 865.050 298.050 ;
        RECT 871.950 297.450 874.050 298.050 ;
        RECT 862.950 296.550 874.050 297.450 ;
        RECT 862.950 295.950 865.050 296.550 ;
        RECT 871.950 295.950 874.050 296.550 ;
        RECT 853.800 289.950 855.900 292.050 ;
        RECT 853.950 288.150 855.750 289.950 ;
        RECT 847.500 284.400 855.900 285.300 ;
        RECT 847.500 283.500 849.300 284.400 ;
        RECT 845.700 280.800 848.400 282.600 ;
        RECT 846.600 276.600 848.400 280.800 ;
        RECT 849.600 276.000 851.400 282.600 ;
        RECT 854.100 276.600 855.900 284.400 ;
        RECT 11.100 266.400 12.900 272.400 ;
        RECT 14.100 267.300 15.900 273.000 ;
        RECT 18.300 267.000 20.100 272.400 ;
        RECT 22.800 267.300 24.600 273.000 ;
        RECT 11.100 265.500 12.600 266.400 ;
        RECT 11.100 264.000 15.600 265.500 ;
        RECT 13.500 263.400 15.600 264.000 ;
        RECT 19.200 264.900 20.100 267.000 ;
        RECT 26.100 266.400 27.900 272.400 ;
        RECT 38.700 269.400 40.500 273.000 ;
        RECT 41.700 267.600 43.500 272.400 ;
        RECT 23.400 265.500 27.900 266.400 ;
        RECT 38.400 266.400 43.500 267.600 ;
        RECT 46.200 266.400 48.000 273.000 ;
        RECT 62.100 269.400 63.900 273.000 ;
        RECT 65.100 269.400 66.900 272.400 ;
        RECT 77.700 269.400 79.500 273.000 ;
        RECT 16.500 261.900 18.300 263.700 ;
        RECT 19.200 262.800 22.200 264.900 ;
        RECT 23.400 263.100 25.500 265.500 ;
        RECT 15.900 261.000 18.000 261.900 ;
        RECT 11.400 259.800 18.000 261.000 ;
        RECT 11.400 259.200 13.200 259.800 ;
        RECT 11.100 256.950 13.200 259.200 ;
        RECT 15.900 256.800 18.000 258.900 ;
        RECT 15.900 255.000 17.700 256.800 ;
        RECT 19.200 256.050 20.100 262.800 ;
        RECT 21.000 258.900 23.100 261.000 ;
        RECT 38.400 259.050 39.300 266.400 ;
        RECT 40.950 259.050 42.750 260.850 ;
        RECT 47.100 259.050 48.900 260.850 ;
        RECT 65.100 259.050 66.300 269.400 ;
        RECT 80.700 267.600 82.500 272.400 ;
        RECT 77.400 266.400 82.500 267.600 ;
        RECT 85.200 266.400 87.000 273.000 ;
        RECT 77.400 259.050 78.300 266.400 ;
        RECT 100.500 264.000 102.300 272.400 ;
        RECT 99.000 262.800 102.300 264.000 ;
        RECT 107.100 263.400 108.900 273.000 ;
        RECT 119.400 266.400 121.200 273.000 ;
        RECT 124.500 265.200 126.300 272.400 ;
        RECT 140.100 266.400 141.900 272.400 ;
        RECT 122.100 264.300 126.300 265.200 ;
        RECT 140.700 264.300 141.900 266.400 ;
        RECT 143.100 267.300 144.900 272.400 ;
        RECT 146.100 268.200 147.900 273.000 ;
        RECT 149.100 267.300 150.900 272.400 ;
        RECT 143.100 265.950 150.900 267.300 ;
        RECT 161.100 267.300 162.900 272.400 ;
        RECT 164.100 268.200 165.900 273.000 ;
        RECT 167.100 267.300 168.900 272.400 ;
        RECT 161.100 265.950 168.900 267.300 ;
        RECT 170.100 266.400 171.900 272.400 ;
        RECT 182.100 266.400 183.900 272.400 ;
        RECT 170.100 264.300 171.300 266.400 ;
        RECT 79.950 259.050 81.750 260.850 ;
        RECT 86.100 259.050 87.900 260.850 ;
        RECT 99.000 259.050 99.900 262.800 ;
        RECT 101.100 259.050 102.900 260.850 ;
        RECT 107.100 259.050 108.900 260.850 ;
        RECT 119.250 259.050 121.050 260.850 ;
        RECT 122.100 259.050 123.300 264.300 ;
        RECT 140.700 263.400 144.300 264.300 ;
        RECT 125.100 259.050 126.900 260.850 ;
        RECT 140.100 259.050 141.900 260.850 ;
        RECT 143.100 259.050 144.300 263.400 ;
        RECT 167.700 263.400 171.300 264.300 ;
        RECT 182.700 264.300 183.900 266.400 ;
        RECT 185.100 267.300 186.900 272.400 ;
        RECT 188.100 268.200 189.900 273.000 ;
        RECT 191.100 267.300 192.900 272.400 ;
        RECT 203.100 269.400 204.900 273.000 ;
        RECT 206.100 269.400 207.900 272.400 ;
        RECT 185.100 265.950 192.900 267.300 ;
        RECT 182.700 263.400 186.300 264.300 ;
        RECT 146.100 259.050 147.900 260.850 ;
        RECT 164.100 259.050 165.900 260.850 ;
        RECT 167.700 259.050 168.900 263.400 ;
        RECT 170.100 259.050 171.900 260.850 ;
        RECT 182.100 259.050 183.900 260.850 ;
        RECT 185.100 259.050 186.300 263.400 ;
        RECT 188.100 259.050 189.900 260.850 ;
        RECT 206.100 259.050 207.300 269.400 ;
        RECT 218.700 265.200 220.500 272.400 ;
        RECT 223.800 266.400 225.600 273.000 ;
        RECT 237.600 268.200 239.400 272.400 ;
        RECT 236.700 266.400 239.400 268.200 ;
        RECT 240.600 266.400 242.400 273.000 ;
        RECT 218.700 264.300 222.900 265.200 ;
        RECT 218.100 259.050 219.900 260.850 ;
        RECT 221.700 259.050 222.900 264.300 ;
        RECT 223.950 259.050 225.750 260.850 ;
        RECT 236.700 259.050 237.600 266.400 ;
        RECT 238.500 264.600 240.300 265.500 ;
        RECT 245.100 264.600 246.900 272.400 ;
        RECT 238.500 263.700 246.900 264.600 ;
        RECT 257.100 264.600 258.900 272.400 ;
        RECT 261.600 266.400 263.400 273.000 ;
        RECT 264.600 268.200 266.400 272.400 ;
        RECT 278.100 269.400 279.900 272.400 ;
        RECT 264.600 266.400 267.300 268.200 ;
        RECT 263.700 264.600 265.500 265.500 ;
        RECT 257.100 263.700 265.500 264.600 ;
        RECT 21.000 257.100 22.800 258.900 ;
        RECT 25.800 256.950 27.900 259.050 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 46.950 256.950 49.050 259.050 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 76.950 256.950 79.050 259.050 ;
        RECT 79.950 256.950 82.050 259.050 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 139.950 256.950 142.050 259.050 ;
        RECT 142.950 256.950 145.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 160.950 256.950 163.050 259.050 ;
        RECT 163.950 256.950 166.050 259.050 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 217.950 256.950 220.050 259.050 ;
        RECT 220.950 256.950 223.050 259.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 236.100 256.950 238.200 259.050 ;
        RECT 239.400 256.950 241.500 259.050 ;
        RECT 19.200 254.700 22.200 256.050 ;
        RECT 25.800 255.150 27.600 256.950 ;
        RECT 20.100 253.950 22.200 254.700 ;
        RECT 17.400 251.700 19.200 253.500 ;
        RECT 13.800 250.800 19.200 251.700 ;
        RECT 13.800 249.900 15.900 250.800 ;
        RECT 11.100 248.700 15.900 249.900 ;
        RECT 20.700 249.600 21.900 253.950 ;
        RECT 18.600 248.700 21.900 249.600 ;
        RECT 22.800 249.600 24.900 250.500 ;
        RECT 38.400 249.600 39.300 256.950 ;
        RECT 43.950 255.150 45.750 256.950 ;
        RECT 62.100 255.150 63.900 256.950 ;
        RECT 40.950 252.450 43.050 253.050 ;
        RECT 61.950 252.450 64.050 253.050 ;
        RECT 40.950 251.550 64.050 252.450 ;
        RECT 40.950 250.950 43.050 251.550 ;
        RECT 61.950 250.950 64.050 251.550 ;
        RECT 11.100 237.600 12.900 248.700 ;
        RECT 14.100 237.000 15.900 247.500 ;
        RECT 18.600 237.600 20.400 248.700 ;
        RECT 22.800 248.400 27.900 249.600 ;
        RECT 22.800 237.000 24.900 247.500 ;
        RECT 26.100 237.600 27.900 248.400 ;
        RECT 38.100 237.600 39.900 249.600 ;
        RECT 41.100 248.700 48.900 249.600 ;
        RECT 41.100 237.600 42.900 248.700 ;
        RECT 44.100 237.000 45.900 247.800 ;
        RECT 47.100 237.600 48.900 248.700 ;
        RECT 65.100 243.600 66.300 256.950 ;
        RECT 77.400 249.600 78.300 256.950 ;
        RECT 82.950 255.150 84.750 256.950 ;
        RECT 62.100 237.000 63.900 243.600 ;
        RECT 65.100 237.600 66.900 243.600 ;
        RECT 77.100 237.600 78.900 249.600 ;
        RECT 80.100 248.700 87.900 249.600 ;
        RECT 80.100 237.600 81.900 248.700 ;
        RECT 83.100 237.000 84.900 247.800 ;
        RECT 86.100 237.600 87.900 248.700 ;
        RECT 99.000 244.800 99.900 256.950 ;
        RECT 104.100 255.150 105.900 256.950 ;
        RECT 99.000 243.900 105.600 244.800 ;
        RECT 99.000 243.600 99.900 243.900 ;
        RECT 98.100 237.600 99.900 243.600 ;
        RECT 104.100 243.600 105.600 243.900 ;
        RECT 122.100 243.600 123.300 256.950 ;
        RECT 143.100 249.600 144.300 256.950 ;
        RECT 149.100 255.150 150.900 256.950 ;
        RECT 161.100 255.150 162.900 256.950 ;
        RECT 167.700 249.600 168.900 256.950 ;
        RECT 143.100 248.100 145.500 249.600 ;
        RECT 141.000 245.100 142.800 246.900 ;
        RECT 101.100 237.000 102.900 243.000 ;
        RECT 104.100 237.600 105.900 243.600 ;
        RECT 107.100 237.000 108.900 243.600 ;
        RECT 119.100 237.000 120.900 243.600 ;
        RECT 122.100 237.600 123.900 243.600 ;
        RECT 125.100 237.000 126.900 243.600 ;
        RECT 140.700 237.000 142.500 243.600 ;
        RECT 143.700 237.600 145.500 248.100 ;
        RECT 148.800 237.000 150.600 249.600 ;
        RECT 161.400 237.000 163.200 249.600 ;
        RECT 166.500 248.100 168.900 249.600 ;
        RECT 185.100 249.600 186.300 256.950 ;
        RECT 191.100 255.150 192.900 256.950 ;
        RECT 203.100 255.150 204.900 256.950 ;
        RECT 185.100 248.100 187.500 249.600 ;
        RECT 166.500 237.600 168.300 248.100 ;
        RECT 169.200 245.100 171.000 246.900 ;
        RECT 183.000 245.100 184.800 246.900 ;
        RECT 169.500 237.000 171.300 243.600 ;
        RECT 182.700 237.000 184.500 243.600 ;
        RECT 185.700 237.600 187.500 248.100 ;
        RECT 190.800 237.000 192.600 249.600 ;
        RECT 206.100 243.600 207.300 256.950 ;
        RECT 221.700 243.600 222.900 256.950 ;
        RECT 236.700 249.600 237.600 256.950 ;
        RECT 240.000 255.150 241.800 256.950 ;
        RECT 203.100 237.000 204.900 243.600 ;
        RECT 206.100 237.600 207.900 243.600 ;
        RECT 218.100 237.000 219.900 243.600 ;
        RECT 221.100 237.600 222.900 243.600 ;
        RECT 224.100 237.000 225.900 243.600 ;
        RECT 236.100 237.600 237.900 249.600 ;
        RECT 239.100 237.000 240.900 249.000 ;
        RECT 243.000 243.600 243.900 263.700 ;
        RECT 244.950 259.050 246.750 260.850 ;
        RECT 257.250 259.050 259.050 260.850 ;
        RECT 244.800 256.950 246.900 259.050 ;
        RECT 257.100 256.950 259.200 259.050 ;
        RECT 260.100 243.600 261.000 263.700 ;
        RECT 266.400 259.050 267.300 266.400 ;
        RECT 278.100 265.500 279.300 269.400 ;
        RECT 281.100 266.400 282.900 273.000 ;
        RECT 284.100 266.400 285.900 272.400 ;
        RECT 296.100 266.400 297.900 273.000 ;
        RECT 299.100 266.400 300.900 272.400 ;
        RECT 278.100 264.600 283.800 265.500 ;
        RECT 282.000 263.700 283.800 264.600 ;
        RECT 262.500 256.950 264.600 259.050 ;
        RECT 265.800 256.950 267.900 259.050 ;
        RECT 278.400 256.950 280.500 259.050 ;
        RECT 262.200 255.150 264.000 256.950 ;
        RECT 266.400 249.600 267.300 256.950 ;
        RECT 278.400 255.150 280.200 256.950 ;
        RECT 282.000 252.300 282.900 263.700 ;
        RECT 284.700 259.050 285.900 266.400 ;
        RECT 296.100 259.050 297.900 260.850 ;
        RECT 299.100 259.050 300.300 266.400 ;
        RECT 311.100 264.600 312.900 272.400 ;
        RECT 315.600 266.400 317.400 273.000 ;
        RECT 318.600 268.200 320.400 272.400 ;
        RECT 318.600 266.400 321.300 268.200 ;
        RECT 317.700 264.600 319.500 265.500 ;
        RECT 311.100 263.700 319.500 264.600 ;
        RECT 301.950 261.450 306.000 262.050 ;
        RECT 301.950 259.950 306.450 261.450 ;
        RECT 283.800 256.950 285.900 259.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 282.000 251.400 283.800 252.300 ;
        RECT 278.100 250.500 283.800 251.400 ;
        RECT 242.100 237.600 243.900 243.600 ;
        RECT 245.100 237.000 246.900 243.600 ;
        RECT 257.100 237.000 258.900 243.600 ;
        RECT 260.100 237.600 261.900 243.600 ;
        RECT 263.100 237.000 264.900 249.000 ;
        RECT 266.100 237.600 267.900 249.600 ;
        RECT 278.100 243.600 279.300 250.500 ;
        RECT 284.700 249.600 285.900 256.950 ;
        RECT 299.100 249.600 300.300 256.950 ;
        RECT 305.550 256.050 306.450 259.950 ;
        RECT 311.250 259.050 313.050 260.850 ;
        RECT 311.100 256.950 313.200 259.050 ;
        RECT 301.950 254.550 306.450 256.050 ;
        RECT 301.950 253.950 306.000 254.550 ;
        RECT 278.100 237.600 279.900 243.600 ;
        RECT 281.100 237.000 282.900 247.800 ;
        RECT 284.100 237.600 285.900 249.600 ;
        RECT 296.100 237.000 297.900 249.600 ;
        RECT 299.100 237.600 300.900 249.600 ;
        RECT 314.100 243.600 315.000 263.700 ;
        RECT 320.400 259.050 321.300 266.400 ;
        RECT 335.100 267.300 336.900 272.400 ;
        RECT 338.100 268.200 339.900 273.000 ;
        RECT 341.100 267.300 342.900 272.400 ;
        RECT 335.100 265.950 342.900 267.300 ;
        RECT 344.100 266.400 345.900 272.400 ;
        RECT 356.400 266.400 358.200 273.000 ;
        RECT 344.100 264.300 345.300 266.400 ;
        RECT 361.500 265.200 363.300 272.400 ;
        RECT 374.100 269.400 375.900 272.400 ;
        RECT 377.100 269.400 378.900 273.000 ;
        RECT 341.700 263.400 345.300 264.300 ;
        RECT 359.100 264.300 363.300 265.200 ;
        RECT 338.100 259.050 339.900 260.850 ;
        RECT 341.700 259.050 342.900 263.400 ;
        RECT 346.950 261.450 351.000 262.050 ;
        RECT 344.100 259.050 345.900 260.850 ;
        RECT 346.950 259.950 351.450 261.450 ;
        RECT 316.500 256.950 318.600 259.050 ;
        RECT 319.800 256.950 321.900 259.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 316.200 255.150 318.000 256.950 ;
        RECT 320.400 249.600 321.300 256.950 ;
        RECT 335.100 255.150 336.900 256.950 ;
        RECT 341.700 249.600 342.900 256.950 ;
        RECT 343.950 252.450 346.050 252.750 ;
        RECT 350.550 252.450 351.450 259.950 ;
        RECT 356.250 259.050 358.050 260.850 ;
        RECT 359.100 259.050 360.300 264.300 ;
        RECT 364.950 261.450 369.000 262.050 ;
        RECT 362.100 259.050 363.900 260.850 ;
        RECT 364.950 259.950 369.450 261.450 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 343.950 251.550 351.450 252.450 ;
        RECT 343.950 250.650 346.050 251.550 ;
        RECT 311.100 237.000 312.900 243.600 ;
        RECT 314.100 237.600 315.900 243.600 ;
        RECT 317.100 237.000 318.900 249.000 ;
        RECT 320.100 237.600 321.900 249.600 ;
        RECT 335.400 237.000 337.200 249.600 ;
        RECT 340.500 248.100 342.900 249.600 ;
        RECT 340.500 237.600 342.300 248.100 ;
        RECT 343.200 245.100 345.000 246.900 ;
        RECT 359.100 243.600 360.300 256.950 ;
        RECT 368.550 256.050 369.450 259.950 ;
        RECT 374.700 259.050 375.900 269.400 ;
        RECT 389.100 263.400 390.900 273.000 ;
        RECT 395.700 264.000 397.500 272.400 ;
        RECT 410.100 266.400 411.900 272.400 ;
        RECT 410.700 264.300 411.900 266.400 ;
        RECT 413.100 267.300 414.900 272.400 ;
        RECT 416.100 268.200 417.900 273.000 ;
        RECT 419.100 267.300 420.900 272.400 ;
        RECT 413.100 265.950 420.900 267.300 ;
        RECT 395.700 262.800 399.000 264.000 ;
        RECT 410.700 263.400 414.300 264.300 ;
        RECT 384.000 261.450 388.050 262.050 ;
        RECT 383.550 259.950 388.050 261.450 ;
        RECT 373.950 256.950 376.050 259.050 ;
        RECT 376.950 256.950 379.050 259.050 ;
        RECT 364.950 254.550 369.450 256.050 ;
        RECT 364.950 253.950 369.000 254.550 ;
        RECT 374.700 243.600 375.900 256.950 ;
        RECT 377.100 255.150 378.900 256.950 ;
        RECT 383.550 256.050 384.450 259.950 ;
        RECT 389.100 259.050 390.900 260.850 ;
        RECT 395.100 259.050 396.900 260.850 ;
        RECT 398.100 259.050 399.000 262.800 ;
        RECT 410.100 259.050 411.900 260.850 ;
        RECT 413.100 259.050 414.300 263.400 ;
        RECT 427.950 262.950 430.050 265.050 ;
        RECT 431.100 264.600 432.900 272.400 ;
        RECT 435.600 266.400 437.400 273.000 ;
        RECT 438.600 268.200 440.400 272.400 ;
        RECT 452.100 269.400 453.900 272.400 ;
        RECT 455.100 269.400 456.900 273.000 ;
        RECT 438.600 266.400 441.300 268.200 ;
        RECT 437.700 264.600 439.500 265.500 ;
        RECT 431.100 263.700 439.500 264.600 ;
        RECT 421.950 261.450 426.000 262.050 ;
        RECT 416.100 259.050 417.900 260.850 ;
        RECT 421.950 259.950 426.450 261.450 ;
        RECT 388.950 256.950 391.050 259.050 ;
        RECT 391.950 256.950 394.050 259.050 ;
        RECT 394.950 256.950 397.050 259.050 ;
        RECT 397.950 256.950 400.050 259.050 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 412.950 256.950 415.050 259.050 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 418.950 256.950 421.050 259.050 ;
        RECT 383.550 254.550 388.050 256.050 ;
        RECT 392.100 255.150 393.900 256.950 ;
        RECT 384.000 253.950 388.050 254.550 ;
        RECT 398.100 244.800 399.000 256.950 ;
        RECT 413.100 249.600 414.300 256.950 ;
        RECT 419.100 255.150 420.900 256.950 ;
        RECT 425.550 255.450 426.450 259.950 ;
        RECT 422.550 254.550 426.450 255.450 ;
        RECT 422.550 253.050 423.450 254.550 ;
        RECT 418.950 251.550 423.450 253.050 ;
        RECT 428.550 253.050 429.450 262.950 ;
        RECT 431.250 259.050 433.050 260.850 ;
        RECT 431.100 256.950 433.200 259.050 ;
        RECT 428.550 251.550 433.050 253.050 ;
        RECT 418.950 250.950 423.000 251.550 ;
        RECT 429.000 250.950 433.050 251.550 ;
        RECT 413.100 248.100 415.500 249.600 ;
        RECT 411.000 245.100 412.800 246.900 ;
        RECT 392.400 243.900 399.000 244.800 ;
        RECT 392.400 243.600 393.900 243.900 ;
        RECT 343.500 237.000 345.300 243.600 ;
        RECT 356.100 237.000 357.900 243.600 ;
        RECT 359.100 237.600 360.900 243.600 ;
        RECT 362.100 237.000 363.900 243.600 ;
        RECT 374.100 237.600 375.900 243.600 ;
        RECT 377.100 237.000 378.900 243.600 ;
        RECT 389.100 237.000 390.900 243.600 ;
        RECT 392.100 237.600 393.900 243.600 ;
        RECT 398.100 243.600 399.000 243.900 ;
        RECT 395.100 237.000 396.900 243.000 ;
        RECT 398.100 237.600 399.900 243.600 ;
        RECT 410.700 237.000 412.500 243.600 ;
        RECT 413.700 237.600 415.500 248.100 ;
        RECT 418.800 237.000 420.600 249.600 ;
        RECT 434.100 243.600 435.000 263.700 ;
        RECT 440.400 259.050 441.300 266.400 ;
        RECT 452.700 259.050 453.900 269.400 ;
        RECT 469.500 264.000 471.300 272.400 ;
        RECT 468.000 262.800 471.300 264.000 ;
        RECT 476.100 263.400 477.900 273.000 ;
        RECT 488.100 267.300 489.900 272.400 ;
        RECT 491.100 268.200 492.900 273.000 ;
        RECT 494.100 267.300 495.900 272.400 ;
        RECT 488.100 265.950 495.900 267.300 ;
        RECT 497.100 266.400 498.900 272.400 ;
        RECT 510.600 268.200 512.400 272.400 ;
        RECT 509.700 266.400 512.400 268.200 ;
        RECT 513.600 266.400 515.400 273.000 ;
        RECT 497.100 264.300 498.300 266.400 ;
        RECT 494.700 263.400 498.300 264.300 ;
        RECT 468.000 259.050 468.900 262.800 ;
        RECT 483.000 261.450 487.050 262.050 ;
        RECT 470.100 259.050 471.900 260.850 ;
        RECT 476.100 259.050 477.900 260.850 ;
        RECT 482.550 259.950 487.050 261.450 ;
        RECT 436.500 256.950 438.600 259.050 ;
        RECT 439.800 256.950 441.900 259.050 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 466.950 256.950 469.050 259.050 ;
        RECT 469.950 256.950 472.050 259.050 ;
        RECT 472.950 256.950 475.050 259.050 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 436.200 255.150 438.000 256.950 ;
        RECT 440.400 249.600 441.300 256.950 ;
        RECT 431.100 237.000 432.900 243.600 ;
        RECT 434.100 237.600 435.900 243.600 ;
        RECT 437.100 237.000 438.900 249.000 ;
        RECT 440.100 237.600 441.900 249.600 ;
        RECT 452.700 243.600 453.900 256.950 ;
        RECT 455.100 255.150 456.900 256.950 ;
        RECT 468.000 244.800 468.900 256.950 ;
        RECT 473.100 255.150 474.900 256.950 ;
        RECT 482.550 256.050 483.450 259.950 ;
        RECT 491.100 259.050 492.900 260.850 ;
        RECT 494.700 259.050 495.900 263.400 ;
        RECT 499.950 261.450 504.000 262.050 ;
        RECT 497.100 259.050 498.900 260.850 ;
        RECT 499.950 259.950 504.450 261.450 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 490.950 256.950 493.050 259.050 ;
        RECT 493.950 256.950 496.050 259.050 ;
        RECT 496.950 256.950 499.050 259.050 ;
        RECT 482.550 254.550 487.050 256.050 ;
        RECT 488.100 255.150 489.900 256.950 ;
        RECT 483.000 253.950 487.050 254.550 ;
        RECT 469.950 252.450 472.050 252.750 ;
        RECT 475.950 252.450 478.050 253.050 ;
        RECT 469.950 251.550 478.050 252.450 ;
        RECT 469.950 250.650 472.050 251.550 ;
        RECT 475.950 250.950 478.050 251.550 ;
        RECT 494.700 249.600 495.900 256.950 ;
        RECT 503.550 256.050 504.450 259.950 ;
        RECT 509.700 259.050 510.600 266.400 ;
        RECT 511.500 264.600 513.300 265.500 ;
        RECT 518.100 264.600 519.900 272.400 ;
        RECT 530.100 266.400 531.900 272.400 ;
        RECT 511.500 263.700 519.900 264.600 ;
        RECT 530.700 264.300 531.900 266.400 ;
        RECT 533.100 267.300 534.900 272.400 ;
        RECT 536.100 268.200 537.900 273.000 ;
        RECT 539.100 267.300 540.900 272.400 ;
        RECT 533.100 265.950 540.900 267.300 ;
        RECT 554.700 265.200 556.500 272.400 ;
        RECT 559.800 266.400 561.600 273.000 ;
        RECT 572.100 266.400 573.900 272.400 ;
        RECT 554.700 264.300 558.900 265.200 ;
        RECT 509.100 256.950 511.200 259.050 ;
        RECT 512.400 256.950 514.500 259.050 ;
        RECT 499.950 254.550 504.450 256.050 ;
        RECT 499.950 253.950 504.000 254.550 ;
        RECT 509.700 249.600 510.600 256.950 ;
        RECT 513.000 255.150 514.800 256.950 ;
        RECT 468.000 243.900 474.600 244.800 ;
        RECT 468.000 243.600 468.900 243.900 ;
        RECT 452.100 237.600 453.900 243.600 ;
        RECT 455.100 237.000 456.900 243.600 ;
        RECT 467.100 237.600 468.900 243.600 ;
        RECT 473.100 243.600 474.600 243.900 ;
        RECT 470.100 237.000 471.900 243.000 ;
        RECT 473.100 237.600 474.900 243.600 ;
        RECT 476.100 237.000 477.900 243.600 ;
        RECT 488.400 237.000 490.200 249.600 ;
        RECT 493.500 248.100 495.900 249.600 ;
        RECT 493.500 237.600 495.300 248.100 ;
        RECT 496.200 245.100 498.000 246.900 ;
        RECT 496.500 237.000 498.300 243.600 ;
        RECT 509.100 237.600 510.900 249.600 ;
        RECT 512.100 237.000 513.900 249.000 ;
        RECT 516.000 243.600 516.900 263.700 ;
        RECT 530.700 263.400 534.300 264.300 ;
        RECT 517.950 259.050 519.750 260.850 ;
        RECT 530.100 259.050 531.900 260.850 ;
        RECT 533.100 259.050 534.300 263.400 ;
        RECT 536.100 259.050 537.900 260.850 ;
        RECT 554.100 259.050 555.900 260.850 ;
        RECT 557.700 259.050 558.900 264.300 ;
        RECT 572.700 264.300 573.900 266.400 ;
        RECT 575.100 267.300 576.900 272.400 ;
        RECT 578.100 268.200 579.900 273.000 ;
        RECT 581.100 267.300 582.900 272.400 ;
        RECT 575.100 265.950 582.900 267.300 ;
        RECT 572.700 263.400 576.300 264.300 ;
        RECT 595.500 264.000 597.300 272.400 ;
        RECT 567.000 261.450 571.050 262.050 ;
        RECT 559.950 259.050 561.750 260.850 ;
        RECT 566.550 259.950 571.050 261.450 ;
        RECT 517.800 256.950 519.900 259.050 ;
        RECT 529.950 256.950 532.050 259.050 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 538.950 256.950 541.050 259.050 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 533.100 249.600 534.300 256.950 ;
        RECT 539.100 255.150 540.900 256.950 ;
        RECT 533.100 248.100 535.500 249.600 ;
        RECT 531.000 245.100 532.800 246.900 ;
        RECT 515.100 237.600 516.900 243.600 ;
        RECT 518.100 237.000 519.900 243.600 ;
        RECT 530.700 237.000 532.500 243.600 ;
        RECT 533.700 237.600 535.500 248.100 ;
        RECT 538.800 237.000 540.600 249.600 ;
        RECT 557.700 243.600 558.900 256.950 ;
        RECT 566.550 256.050 567.450 259.950 ;
        RECT 572.100 259.050 573.900 260.850 ;
        RECT 575.100 259.050 576.300 263.400 ;
        RECT 594.000 262.800 597.300 264.000 ;
        RECT 602.100 263.400 603.900 273.000 ;
        RECT 614.100 269.400 615.900 272.400 ;
        RECT 617.100 269.400 618.900 273.000 ;
        RECT 588.000 261.900 591.000 262.050 ;
        RECT 588.000 261.450 592.050 261.900 ;
        RECT 578.100 259.050 579.900 260.850 ;
        RECT 587.550 259.950 592.050 261.450 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 562.950 254.550 567.450 256.050 ;
        RECT 562.950 253.950 567.000 254.550 ;
        RECT 575.100 249.600 576.300 256.950 ;
        RECT 581.100 255.150 582.900 256.950 ;
        RECT 587.550 256.050 588.450 259.950 ;
        RECT 589.950 259.800 592.050 259.950 ;
        RECT 594.000 259.050 594.900 262.800 ;
        RECT 604.950 261.450 609.000 262.050 ;
        RECT 596.100 259.050 597.900 260.850 ;
        RECT 602.100 259.050 603.900 260.850 ;
        RECT 604.950 259.950 609.450 261.450 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 595.950 256.950 598.050 259.050 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 583.950 254.550 588.450 256.050 ;
        RECT 583.950 253.950 588.000 254.550 ;
        RECT 577.950 252.450 580.050 253.050 ;
        RECT 589.950 252.450 592.050 253.050 ;
        RECT 577.950 251.550 592.050 252.450 ;
        RECT 577.950 250.950 580.050 251.550 ;
        RECT 589.950 250.950 592.050 251.550 ;
        RECT 575.100 248.100 577.500 249.600 ;
        RECT 573.000 245.100 574.800 246.900 ;
        RECT 554.100 237.000 555.900 243.600 ;
        RECT 557.100 237.600 558.900 243.600 ;
        RECT 560.100 237.000 561.900 243.600 ;
        RECT 572.700 237.000 574.500 243.600 ;
        RECT 575.700 237.600 577.500 248.100 ;
        RECT 580.800 237.000 582.600 249.600 ;
        RECT 594.000 244.800 594.900 256.950 ;
        RECT 599.100 255.150 600.900 256.950 ;
        RECT 608.550 256.050 609.450 259.950 ;
        RECT 614.700 259.050 615.900 269.400 ;
        RECT 629.100 263.400 630.900 273.000 ;
        RECT 635.700 264.000 637.500 272.400 ;
        RECT 650.100 266.400 651.900 272.400 ;
        RECT 635.700 262.800 639.000 264.000 ;
        RECT 619.950 261.450 624.000 262.050 ;
        RECT 619.950 259.950 624.450 261.450 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 608.550 254.550 613.050 256.050 ;
        RECT 609.000 253.950 613.050 254.550 ;
        RECT 594.000 243.900 600.600 244.800 ;
        RECT 594.000 243.600 594.900 243.900 ;
        RECT 593.100 237.600 594.900 243.600 ;
        RECT 599.100 243.600 600.600 243.900 ;
        RECT 614.700 243.600 615.900 256.950 ;
        RECT 617.100 255.150 618.900 256.950 ;
        RECT 623.550 256.050 624.450 259.950 ;
        RECT 629.100 259.050 630.900 260.850 ;
        RECT 635.100 259.050 636.900 260.850 ;
        RECT 638.100 259.050 639.000 262.800 ;
        RECT 640.950 261.450 643.050 264.900 ;
        RECT 650.700 264.300 651.900 266.400 ;
        RECT 653.100 267.300 654.900 272.400 ;
        RECT 656.100 268.200 657.900 273.000 ;
        RECT 659.100 267.300 660.900 272.400 ;
        RECT 671.100 269.400 672.900 273.000 ;
        RECT 674.100 269.400 675.900 272.400 ;
        RECT 677.100 269.400 678.900 273.000 ;
        RECT 653.100 265.950 660.900 267.300 ;
        RECT 650.700 263.400 654.300 264.300 ;
        RECT 646.950 261.450 649.050 262.050 ;
        RECT 640.950 261.000 649.050 261.450 ;
        RECT 641.550 260.550 649.050 261.000 ;
        RECT 646.950 259.950 649.050 260.550 ;
        RECT 650.100 259.050 651.900 260.850 ;
        RECT 653.100 259.050 654.300 263.400 ;
        RECT 661.950 261.450 666.000 262.050 ;
        RECT 656.100 259.050 657.900 260.850 ;
        RECT 661.950 259.950 666.450 261.450 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 637.950 256.950 640.050 259.050 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 619.950 254.550 624.450 256.050 ;
        RECT 632.100 255.150 633.900 256.950 ;
        RECT 619.950 253.950 624.000 254.550 ;
        RECT 616.950 249.450 619.050 250.050 ;
        RECT 631.950 249.450 634.050 250.050 ;
        RECT 616.950 248.550 634.050 249.450 ;
        RECT 616.950 247.950 619.050 248.550 ;
        RECT 631.950 247.950 634.050 248.550 ;
        RECT 638.100 244.800 639.000 256.950 ;
        RECT 653.100 249.600 654.300 256.950 ;
        RECT 659.100 255.150 660.900 256.950 ;
        RECT 665.550 255.450 666.450 259.950 ;
        RECT 674.700 259.050 675.600 269.400 ;
        RECT 689.400 266.400 691.200 273.000 ;
        RECT 694.500 265.200 696.300 272.400 ;
        RECT 707.100 269.400 708.900 273.000 ;
        RECT 710.100 269.400 711.900 272.400 ;
        RECT 713.100 269.400 714.900 273.000 ;
        RECT 692.100 264.300 696.300 265.200 ;
        RECT 684.000 261.450 688.050 262.050 ;
        RECT 683.550 259.950 688.050 261.450 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 665.550 254.550 669.450 255.450 ;
        RECT 671.100 255.150 672.900 256.950 ;
        RECT 668.550 253.050 669.450 254.550 ;
        RECT 668.550 251.550 673.050 253.050 ;
        RECT 669.000 250.950 673.050 251.550 ;
        RECT 674.700 249.600 675.600 256.950 ;
        RECT 676.950 255.150 678.750 256.950 ;
        RECT 683.550 256.050 684.450 259.950 ;
        RECT 689.250 259.050 691.050 260.850 ;
        RECT 692.100 259.050 693.300 264.300 ;
        RECT 695.100 259.050 696.900 260.850 ;
        RECT 710.400 259.050 711.300 269.400 ;
        RECT 725.100 267.300 726.900 272.400 ;
        RECT 728.100 268.200 729.900 273.000 ;
        RECT 731.100 267.300 732.900 272.400 ;
        RECT 725.100 265.950 732.900 267.300 ;
        RECT 734.100 266.400 735.900 272.400 ;
        RECT 734.100 264.300 735.300 266.400 ;
        RECT 731.700 263.400 735.300 264.300 ;
        RECT 751.500 264.000 753.300 272.400 ;
        RECT 720.000 261.450 724.050 262.050 ;
        RECT 719.550 259.950 724.050 261.450 ;
        RECT 688.950 256.950 691.050 259.050 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 709.950 256.950 712.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 683.550 254.550 688.050 256.050 ;
        RECT 684.000 253.950 688.050 254.550 ;
        RECT 653.100 248.100 655.500 249.600 ;
        RECT 651.000 245.100 652.800 246.900 ;
        RECT 632.400 243.900 639.000 244.800 ;
        RECT 632.400 243.600 633.900 243.900 ;
        RECT 596.100 237.000 597.900 243.000 ;
        RECT 599.100 237.600 600.900 243.600 ;
        RECT 602.100 237.000 603.900 243.600 ;
        RECT 614.100 237.600 615.900 243.600 ;
        RECT 617.100 237.000 618.900 243.600 ;
        RECT 629.100 237.000 630.900 243.600 ;
        RECT 632.100 237.600 633.900 243.600 ;
        RECT 638.100 243.600 639.000 243.900 ;
        RECT 635.100 237.000 636.900 243.000 ;
        RECT 638.100 237.600 639.900 243.600 ;
        RECT 650.700 237.000 652.500 243.600 ;
        RECT 653.700 237.600 655.500 248.100 ;
        RECT 658.800 237.000 660.600 249.600 ;
        RECT 672.000 248.400 675.600 249.600 ;
        RECT 672.000 237.600 673.800 248.400 ;
        RECT 677.100 237.000 678.900 249.600 ;
        RECT 692.100 243.600 693.300 256.950 ;
        RECT 707.250 255.150 709.050 256.950 ;
        RECT 710.400 249.600 711.300 256.950 ;
        RECT 713.100 255.150 714.900 256.950 ;
        RECT 712.950 252.450 715.050 253.050 ;
        RECT 719.550 252.450 720.450 259.950 ;
        RECT 728.100 259.050 729.900 260.850 ;
        RECT 731.700 259.050 732.900 263.400 ;
        RECT 750.000 262.800 753.300 264.000 ;
        RECT 758.100 263.400 759.900 273.000 ;
        RECT 770.400 266.400 772.200 273.000 ;
        RECT 775.500 265.200 777.300 272.400 ;
        RECT 773.100 264.300 777.300 265.200 ;
        RECT 734.100 259.050 735.900 260.850 ;
        RECT 750.000 259.050 750.900 262.800 ;
        RECT 765.000 261.450 769.050 262.050 ;
        RECT 752.100 259.050 753.900 260.850 ;
        RECT 758.100 259.050 759.900 260.850 ;
        RECT 764.550 259.950 769.050 261.450 ;
        RECT 724.950 256.950 727.050 259.050 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 730.950 256.950 733.050 259.050 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 748.950 256.950 751.050 259.050 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 725.100 255.150 726.900 256.950 ;
        RECT 712.950 251.550 720.450 252.450 ;
        RECT 712.950 250.950 715.050 251.550 ;
        RECT 731.700 249.600 732.900 256.950 ;
        RECT 689.100 237.000 690.900 243.600 ;
        RECT 692.100 237.600 693.900 243.600 ;
        RECT 695.100 237.000 696.900 243.600 ;
        RECT 707.100 237.000 708.900 249.600 ;
        RECT 710.400 248.400 714.000 249.600 ;
        RECT 712.200 237.600 714.000 248.400 ;
        RECT 725.400 237.000 727.200 249.600 ;
        RECT 730.500 248.100 732.900 249.600 ;
        RECT 730.500 237.600 732.300 248.100 ;
        RECT 733.200 245.100 735.000 246.900 ;
        RECT 750.000 244.800 750.900 256.950 ;
        RECT 755.100 255.150 756.900 256.950 ;
        RECT 764.550 256.050 765.450 259.950 ;
        RECT 770.250 259.050 772.050 260.850 ;
        RECT 773.100 259.050 774.300 264.300 ;
        RECT 790.500 264.000 792.300 272.400 ;
        RECT 789.000 262.800 792.300 264.000 ;
        RECT 797.100 263.400 798.900 273.000 ;
        RECT 809.100 263.400 810.900 273.000 ;
        RECT 815.700 264.000 817.500 272.400 ;
        RECT 832.500 264.000 834.300 272.400 ;
        RECT 815.700 262.800 819.000 264.000 ;
        RECT 783.000 261.450 787.050 262.050 ;
        RECT 776.100 259.050 777.900 260.850 ;
        RECT 782.550 259.950 787.050 261.450 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 760.950 254.550 765.450 256.050 ;
        RECT 760.950 253.950 765.000 254.550 ;
        RECT 750.000 243.900 756.600 244.800 ;
        RECT 750.000 243.600 750.900 243.900 ;
        RECT 733.500 237.000 735.300 243.600 ;
        RECT 749.100 237.600 750.900 243.600 ;
        RECT 755.100 243.600 756.600 243.900 ;
        RECT 773.100 243.600 774.300 256.950 ;
        RECT 782.550 256.050 783.450 259.950 ;
        RECT 789.000 259.050 789.900 262.800 ;
        RECT 791.100 259.050 792.900 260.850 ;
        RECT 797.100 259.050 798.900 260.850 ;
        RECT 809.100 259.050 810.900 260.850 ;
        RECT 815.100 259.050 816.900 260.850 ;
        RECT 818.100 259.050 819.000 262.800 ;
        RECT 831.000 262.800 834.300 264.000 ;
        RECT 839.100 263.400 840.900 273.000 ;
        RECT 851.100 269.400 852.900 273.000 ;
        RECT 854.100 269.400 855.900 272.400 ;
        RECT 831.000 259.050 831.900 262.800 ;
        RECT 846.000 261.450 850.050 262.050 ;
        RECT 833.100 259.050 834.900 260.850 ;
        RECT 839.100 259.050 840.900 260.850 ;
        RECT 845.550 259.950 850.050 261.450 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 835.950 256.950 838.050 259.050 ;
        RECT 838.950 256.950 841.050 259.050 ;
        RECT 782.550 254.550 787.050 256.050 ;
        RECT 783.000 253.950 787.050 254.550 ;
        RECT 789.000 244.800 789.900 256.950 ;
        RECT 794.100 255.150 795.900 256.950 ;
        RECT 812.100 255.150 813.900 256.950 ;
        RECT 818.100 244.800 819.000 256.950 ;
        RECT 789.000 243.900 795.600 244.800 ;
        RECT 789.000 243.600 789.900 243.900 ;
        RECT 752.100 237.000 753.900 243.000 ;
        RECT 755.100 237.600 756.900 243.600 ;
        RECT 758.100 237.000 759.900 243.600 ;
        RECT 770.100 237.000 771.900 243.600 ;
        RECT 773.100 237.600 774.900 243.600 ;
        RECT 776.100 237.000 777.900 243.600 ;
        RECT 788.100 237.600 789.900 243.600 ;
        RECT 794.100 243.600 795.600 243.900 ;
        RECT 812.400 243.900 819.000 244.800 ;
        RECT 812.400 243.600 813.900 243.900 ;
        RECT 791.100 237.000 792.900 243.000 ;
        RECT 794.100 237.600 795.900 243.600 ;
        RECT 797.100 237.000 798.900 243.600 ;
        RECT 809.100 237.000 810.900 243.600 ;
        RECT 812.100 237.600 813.900 243.600 ;
        RECT 818.100 243.600 819.000 243.900 ;
        RECT 831.000 244.800 831.900 256.950 ;
        RECT 836.100 255.150 837.900 256.950 ;
        RECT 845.550 256.050 846.450 259.950 ;
        RECT 854.100 259.050 855.300 269.400 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 845.550 254.550 850.050 256.050 ;
        RECT 851.100 255.150 852.900 256.950 ;
        RECT 846.000 253.950 850.050 254.550 ;
        RECT 831.000 243.900 837.600 244.800 ;
        RECT 831.000 243.600 831.900 243.900 ;
        RECT 815.100 237.000 816.900 243.000 ;
        RECT 818.100 237.600 819.900 243.600 ;
        RECT 830.100 237.600 831.900 243.600 ;
        RECT 836.100 243.600 837.600 243.900 ;
        RECT 854.100 243.600 855.300 256.950 ;
        RECT 833.100 237.000 834.900 243.000 ;
        RECT 836.100 237.600 837.900 243.600 ;
        RECT 839.100 237.000 840.900 243.600 ;
        RECT 851.100 237.000 852.900 243.600 ;
        RECT 854.100 237.600 855.900 243.600 ;
        RECT 11.100 227.400 12.900 234.000 ;
        RECT 14.100 227.400 15.900 233.400 ;
        RECT 17.100 227.400 18.900 234.000 ;
        RECT 14.100 214.050 15.300 227.400 ;
        RECT 29.400 221.400 31.200 234.000 ;
        RECT 34.500 222.900 36.300 233.400 ;
        RECT 37.500 227.400 39.300 234.000 ;
        RECT 50.100 227.400 51.900 233.400 ;
        RECT 53.100 227.400 54.900 234.000 ;
        RECT 65.700 227.400 67.500 234.000 ;
        RECT 37.200 224.100 39.000 225.900 ;
        RECT 34.500 221.400 36.900 222.900 ;
        RECT 16.950 219.450 19.050 220.050 ;
        RECT 28.950 219.450 31.050 220.050 ;
        RECT 16.950 218.550 31.050 219.450 ;
        RECT 16.950 217.950 19.050 218.550 ;
        RECT 28.950 217.950 31.050 218.550 ;
        RECT 29.100 214.050 30.900 215.850 ;
        RECT 35.700 214.050 36.900 221.400 ;
        RECT 50.700 214.050 51.900 227.400 ;
        RECT 66.000 224.100 67.800 225.900 ;
        RECT 68.700 222.900 70.500 233.400 ;
        RECT 68.100 221.400 70.500 222.900 ;
        RECT 73.800 221.400 75.600 234.000 ;
        RECT 86.100 227.400 87.900 233.400 ;
        RECT 89.100 228.000 90.900 234.000 ;
        RECT 87.000 227.100 87.900 227.400 ;
        RECT 92.100 227.400 93.900 233.400 ;
        RECT 95.100 227.400 96.900 234.000 ;
        RECT 107.700 227.400 109.500 234.000 ;
        RECT 92.100 227.100 93.600 227.400 ;
        RECT 87.000 226.200 93.600 227.100 ;
        RECT 53.100 214.050 54.900 215.850 ;
        RECT 68.100 214.050 69.300 221.400 ;
        RECT 74.100 214.050 75.900 215.850 ;
        RECT 87.000 214.050 87.900 226.200 ;
        RECT 108.000 224.100 109.800 225.900 ;
        RECT 110.700 222.900 112.500 233.400 ;
        RECT 110.100 221.400 112.500 222.900 ;
        RECT 115.800 221.400 117.600 234.000 ;
        RECT 128.100 221.400 129.900 233.400 ;
        RECT 131.100 222.300 132.900 233.400 ;
        RECT 134.100 223.200 135.900 234.000 ;
        RECT 137.100 222.300 138.900 233.400 ;
        RECT 131.100 221.400 138.900 222.300 ;
        RECT 150.000 222.600 151.800 233.400 ;
        RECT 150.000 221.400 153.600 222.600 ;
        RECT 155.100 221.400 156.900 234.000 ;
        RECT 167.100 227.400 168.900 234.000 ;
        RECT 170.100 227.400 171.900 233.400 ;
        RECT 173.100 227.400 174.900 234.000 ;
        RECT 185.100 227.400 186.900 234.000 ;
        RECT 188.100 227.400 189.900 233.400 ;
        RECT 191.100 227.400 192.900 234.000 ;
        RECT 206.100 227.400 207.900 234.000 ;
        RECT 209.100 227.400 210.900 233.400 ;
        RECT 212.100 227.400 213.900 234.000 ;
        RECT 227.100 227.400 228.900 234.000 ;
        RECT 230.100 227.400 231.900 233.400 ;
        RECT 233.100 227.400 234.900 234.000 ;
        RECT 92.100 214.050 93.900 215.850 ;
        RECT 110.100 214.050 111.300 221.400 ;
        RECT 116.100 214.050 117.900 215.850 ;
        RECT 128.400 214.050 129.300 221.400 ;
        RECT 133.950 214.050 135.750 215.850 ;
        RECT 149.100 214.050 150.900 215.850 ;
        RECT 152.700 214.050 153.600 221.400 ;
        RECT 154.950 214.050 156.750 215.850 ;
        RECT 170.100 214.050 171.300 227.400 ;
        RECT 188.700 214.050 189.900 227.400 ;
        RECT 201.000 216.450 205.050 217.050 ;
        RECT 200.550 214.950 205.050 216.450 ;
        RECT 10.950 211.950 13.050 214.050 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 28.950 211.950 31.050 214.050 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 109.950 211.950 112.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 127.950 211.950 130.050 214.050 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 148.950 211.950 151.050 214.050 ;
        RECT 151.950 211.950 154.050 214.050 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 184.950 211.950 187.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 11.250 210.150 13.050 211.950 ;
        RECT 14.100 206.700 15.300 211.950 ;
        RECT 17.100 210.150 18.900 211.950 ;
        RECT 32.100 210.150 33.900 211.950 ;
        RECT 35.700 207.600 36.900 211.950 ;
        RECT 38.100 210.150 39.900 211.950 ;
        RECT 35.700 206.700 39.300 207.600 ;
        RECT 14.100 205.800 18.300 206.700 ;
        RECT 11.400 198.000 13.200 204.600 ;
        RECT 16.500 198.600 18.300 205.800 ;
        RECT 29.100 203.700 36.900 205.050 ;
        RECT 29.100 198.600 30.900 203.700 ;
        RECT 32.100 198.000 33.900 202.800 ;
        RECT 35.100 198.600 36.900 203.700 ;
        RECT 38.100 204.600 39.300 206.700 ;
        RECT 38.100 198.600 39.900 204.600 ;
        RECT 50.700 201.600 51.900 211.950 ;
        RECT 65.100 210.150 66.900 211.950 ;
        RECT 68.100 207.600 69.300 211.950 ;
        RECT 71.100 210.150 72.900 211.950 ;
        RECT 65.700 206.700 69.300 207.600 ;
        RECT 87.000 208.200 87.900 211.950 ;
        RECT 89.100 210.150 90.900 211.950 ;
        RECT 95.100 210.150 96.900 211.950 ;
        RECT 107.100 210.150 108.900 211.950 ;
        RECT 87.000 207.000 90.300 208.200 ;
        RECT 110.100 207.600 111.300 211.950 ;
        RECT 113.100 210.150 114.900 211.950 ;
        RECT 65.700 204.600 66.900 206.700 ;
        RECT 50.100 198.600 51.900 201.600 ;
        RECT 53.100 198.000 54.900 201.600 ;
        RECT 65.100 198.600 66.900 204.600 ;
        RECT 68.100 203.700 75.900 205.050 ;
        RECT 68.100 198.600 69.900 203.700 ;
        RECT 71.100 198.000 72.900 202.800 ;
        RECT 74.100 198.600 75.900 203.700 ;
        RECT 88.500 198.600 90.300 207.000 ;
        RECT 95.100 198.000 96.900 207.600 ;
        RECT 107.700 206.700 111.300 207.600 ;
        RECT 107.700 204.600 108.900 206.700 ;
        RECT 107.100 198.600 108.900 204.600 ;
        RECT 110.100 203.700 117.900 205.050 ;
        RECT 110.100 198.600 111.900 203.700 ;
        RECT 113.100 198.000 114.900 202.800 ;
        RECT 116.100 198.600 117.900 203.700 ;
        RECT 128.400 204.600 129.300 211.950 ;
        RECT 130.950 210.150 132.750 211.950 ;
        RECT 137.100 210.150 138.900 211.950 ;
        RECT 128.400 203.400 133.500 204.600 ;
        RECT 128.700 198.000 130.500 201.600 ;
        RECT 131.700 198.600 133.500 203.400 ;
        RECT 136.200 198.000 138.000 204.600 ;
        RECT 152.700 201.600 153.600 211.950 ;
        RECT 167.250 210.150 169.050 211.950 ;
        RECT 170.100 206.700 171.300 211.950 ;
        RECT 173.100 210.150 174.900 211.950 ;
        RECT 185.100 210.150 186.900 211.950 ;
        RECT 188.700 206.700 189.900 211.950 ;
        RECT 190.950 210.150 192.750 211.950 ;
        RECT 200.550 211.050 201.450 214.950 ;
        RECT 209.100 214.050 210.300 227.400 ;
        RECT 230.700 214.050 231.900 227.400 ;
        RECT 245.100 221.400 246.900 233.400 ;
        RECT 248.100 222.300 249.900 233.400 ;
        RECT 251.100 223.200 252.900 234.000 ;
        RECT 254.100 222.300 255.900 233.400 ;
        RECT 266.700 227.400 268.500 234.000 ;
        RECT 267.000 224.100 268.800 225.900 ;
        RECT 269.700 222.900 271.500 233.400 ;
        RECT 248.100 221.400 255.900 222.300 ;
        RECT 269.100 221.400 271.500 222.900 ;
        RECT 274.800 221.400 276.600 234.000 ;
        RECT 287.100 221.400 288.900 233.400 ;
        RECT 290.100 223.200 291.900 234.000 ;
        RECT 293.100 227.400 294.900 233.400 ;
        RECT 305.700 227.400 307.500 234.000 ;
        RECT 235.950 216.450 240.000 217.050 ;
        RECT 235.950 214.950 240.450 216.450 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 229.950 211.950 232.050 214.050 ;
        RECT 232.950 211.950 235.050 214.050 ;
        RECT 200.550 209.550 205.050 211.050 ;
        RECT 206.250 210.150 208.050 211.950 ;
        RECT 201.000 208.950 205.050 209.550 ;
        RECT 170.100 205.800 174.300 206.700 ;
        RECT 149.100 198.000 150.900 201.600 ;
        RECT 152.100 198.600 153.900 201.600 ;
        RECT 155.100 198.000 156.900 201.600 ;
        RECT 167.400 198.000 169.200 204.600 ;
        RECT 172.500 198.600 174.300 205.800 ;
        RECT 185.700 205.800 189.900 206.700 ;
        RECT 209.100 206.700 210.300 211.950 ;
        RECT 212.100 210.150 213.900 211.950 ;
        RECT 227.100 210.150 228.900 211.950 ;
        RECT 230.700 206.700 231.900 211.950 ;
        RECT 232.950 210.150 234.750 211.950 ;
        RECT 239.550 211.050 240.450 214.950 ;
        RECT 245.400 214.050 246.300 221.400 ;
        RECT 250.950 214.050 252.750 215.850 ;
        RECT 269.100 214.050 270.300 221.400 ;
        RECT 275.100 214.050 276.900 215.850 ;
        RECT 287.100 214.050 288.300 221.400 ;
        RECT 293.700 220.500 294.900 227.400 ;
        RECT 306.000 224.100 307.800 225.900 ;
        RECT 308.700 222.900 310.500 233.400 ;
        RECT 289.200 219.600 294.900 220.500 ;
        RECT 308.100 221.400 310.500 222.900 ;
        RECT 313.800 221.400 315.600 234.000 ;
        RECT 326.700 227.400 328.500 234.000 ;
        RECT 327.000 224.100 328.800 225.900 ;
        RECT 329.700 222.900 331.500 233.400 ;
        RECT 329.100 221.400 331.500 222.900 ;
        RECT 334.800 221.400 336.600 234.000 ;
        RECT 347.100 227.400 348.900 234.000 ;
        RECT 350.100 227.400 351.900 233.400 ;
        RECT 353.100 227.400 354.900 234.000 ;
        RECT 368.100 227.400 369.900 233.400 ;
        RECT 371.100 228.000 372.900 234.000 ;
        RECT 289.200 218.700 291.000 219.600 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 211.950 256.050 214.050 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 287.100 211.950 289.200 214.050 ;
        RECT 239.550 209.550 244.050 211.050 ;
        RECT 240.000 208.950 244.050 209.550 ;
        RECT 209.100 205.800 213.300 206.700 ;
        RECT 185.700 198.600 187.500 205.800 ;
        RECT 190.800 198.000 192.600 204.600 ;
        RECT 206.400 198.000 208.200 204.600 ;
        RECT 211.500 198.600 213.300 205.800 ;
        RECT 227.700 205.800 231.900 206.700 ;
        RECT 227.700 198.600 229.500 205.800 ;
        RECT 245.400 204.600 246.300 211.950 ;
        RECT 247.950 210.150 249.750 211.950 ;
        RECT 254.100 210.150 255.900 211.950 ;
        RECT 266.100 210.150 267.900 211.950 ;
        RECT 269.100 207.600 270.300 211.950 ;
        RECT 272.100 210.150 273.900 211.950 ;
        RECT 266.700 206.700 270.300 207.600 ;
        RECT 266.700 204.600 267.900 206.700 ;
        RECT 232.800 198.000 234.600 204.600 ;
        RECT 245.400 203.400 250.500 204.600 ;
        RECT 245.700 198.000 247.500 201.600 ;
        RECT 248.700 198.600 250.500 203.400 ;
        RECT 253.200 198.000 255.000 204.600 ;
        RECT 266.100 198.600 267.900 204.600 ;
        RECT 269.100 203.700 276.900 205.050 ;
        RECT 269.100 198.600 270.900 203.700 ;
        RECT 272.100 198.000 273.900 202.800 ;
        RECT 275.100 198.600 276.900 203.700 ;
        RECT 287.100 204.600 288.300 211.950 ;
        RECT 290.100 207.300 291.000 218.700 ;
        RECT 292.800 214.050 294.600 215.850 ;
        RECT 308.100 214.050 309.300 221.400 ;
        RECT 316.950 216.450 321.000 217.050 ;
        RECT 314.100 214.050 315.900 215.850 ;
        RECT 316.950 214.950 321.450 216.450 ;
        RECT 292.500 211.950 294.600 214.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 307.950 211.950 310.050 214.050 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 305.100 210.150 306.900 211.950 ;
        RECT 308.100 207.600 309.300 211.950 ;
        RECT 311.100 210.150 312.900 211.950 ;
        RECT 320.550 211.050 321.450 214.950 ;
        RECT 329.100 214.050 330.300 221.400 ;
        RECT 335.100 214.050 336.900 215.850 ;
        RECT 350.700 214.050 351.900 227.400 ;
        RECT 369.000 227.100 369.900 227.400 ;
        RECT 374.100 227.400 375.900 233.400 ;
        RECT 377.100 227.400 378.900 234.000 ;
        RECT 389.700 227.400 391.500 234.000 ;
        RECT 374.100 227.100 375.600 227.400 ;
        RECT 369.000 226.200 375.600 227.100 ;
        RECT 369.000 214.050 369.900 226.200 ;
        RECT 390.000 224.100 391.800 225.900 ;
        RECT 392.700 222.900 394.500 233.400 ;
        RECT 392.100 221.400 394.500 222.900 ;
        RECT 397.800 221.400 399.600 234.000 ;
        RECT 410.100 227.400 411.900 234.000 ;
        RECT 413.100 227.400 414.900 233.400 ;
        RECT 416.100 227.400 417.900 234.000 ;
        RECT 428.100 227.400 429.900 234.000 ;
        RECT 431.100 227.400 432.900 233.400 ;
        RECT 434.100 227.400 435.900 234.000 ;
        RECT 446.700 227.400 448.500 234.000 ;
        RECT 384.000 216.450 388.050 217.050 ;
        RECT 374.100 214.050 375.900 215.850 ;
        RECT 383.550 214.950 388.050 216.450 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 328.950 211.950 331.050 214.050 ;
        RECT 331.950 211.950 334.050 214.050 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 346.950 211.950 349.050 214.050 ;
        RECT 349.950 211.950 352.050 214.050 ;
        RECT 352.950 211.950 355.050 214.050 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 373.950 211.950 376.050 214.050 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 320.550 209.550 325.050 211.050 ;
        RECT 326.100 210.150 327.900 211.950 ;
        RECT 321.000 208.950 325.050 209.550 ;
        RECT 329.100 207.600 330.300 211.950 ;
        RECT 332.100 210.150 333.900 211.950 ;
        RECT 347.100 210.150 348.900 211.950 ;
        RECT 289.200 206.400 291.000 207.300 ;
        RECT 305.700 206.700 309.300 207.600 ;
        RECT 326.700 206.700 330.300 207.600 ;
        RECT 350.700 206.700 351.900 211.950 ;
        RECT 352.950 210.150 354.750 211.950 ;
        RECT 369.000 208.200 369.900 211.950 ;
        RECT 371.100 210.150 372.900 211.950 ;
        RECT 377.100 210.150 378.900 211.950 ;
        RECT 383.550 211.050 384.450 214.950 ;
        RECT 392.100 214.050 393.300 221.400 ;
        RECT 397.950 219.450 400.050 220.050 ;
        RECT 409.950 219.450 412.050 220.050 ;
        RECT 397.950 218.550 412.050 219.450 ;
        RECT 397.950 217.950 400.050 218.550 ;
        RECT 409.950 217.950 412.050 218.550 ;
        RECT 398.100 214.050 399.900 215.850 ;
        RECT 413.100 214.050 414.300 227.400 ;
        RECT 431.100 214.050 432.300 227.400 ;
        RECT 447.000 224.100 448.800 225.900 ;
        RECT 449.700 222.900 451.500 233.400 ;
        RECT 449.100 221.400 451.500 222.900 ;
        RECT 454.800 221.400 456.600 234.000 ;
        RECT 467.100 227.400 468.900 234.000 ;
        RECT 470.100 227.400 471.900 233.400 ;
        RECT 473.100 228.000 474.900 234.000 ;
        RECT 470.400 227.100 471.900 227.400 ;
        RECT 476.100 227.400 477.900 233.400 ;
        RECT 488.100 227.400 489.900 234.000 ;
        RECT 491.100 227.400 492.900 233.400 ;
        RECT 494.100 227.400 495.900 234.000 ;
        RECT 509.100 227.400 510.900 234.000 ;
        RECT 512.100 227.400 513.900 233.400 ;
        RECT 515.100 227.400 516.900 234.000 ;
        RECT 476.100 227.100 477.000 227.400 ;
        RECT 470.400 226.200 477.000 227.100 ;
        RECT 449.100 214.050 450.300 221.400 ;
        RECT 455.100 214.050 456.900 215.850 ;
        RECT 470.100 214.050 471.900 215.850 ;
        RECT 476.100 214.050 477.000 226.200 ;
        RECT 491.700 214.050 492.900 227.400 ;
        RECT 512.700 214.050 513.900 227.400 ;
        RECT 527.100 221.400 528.900 233.400 ;
        RECT 530.100 222.000 531.900 234.000 ;
        RECT 533.100 227.400 534.900 233.400 ;
        RECT 536.100 227.400 537.900 234.000 ;
        RECT 548.100 227.400 549.900 233.400 ;
        RECT 527.700 214.050 528.600 221.400 ;
        RECT 531.000 214.050 532.800 215.850 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 391.950 211.950 394.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 412.950 211.950 415.050 214.050 ;
        RECT 415.950 211.950 418.050 214.050 ;
        RECT 427.950 211.950 430.050 214.050 ;
        RECT 430.950 211.950 433.050 214.050 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 448.950 211.950 451.050 214.050 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 454.950 211.950 457.050 214.050 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 469.950 211.950 472.050 214.050 ;
        RECT 472.950 211.950 475.050 214.050 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 508.950 211.950 511.050 214.050 ;
        RECT 511.950 211.950 514.050 214.050 ;
        RECT 514.950 211.950 517.050 214.050 ;
        RECT 527.100 211.950 529.200 214.050 ;
        RECT 530.400 211.950 532.500 214.050 ;
        RECT 383.550 209.550 388.050 211.050 ;
        RECT 389.100 210.150 390.900 211.950 ;
        RECT 384.000 208.950 388.050 209.550 ;
        RECT 369.000 207.000 372.300 208.200 ;
        RECT 392.100 207.600 393.300 211.950 ;
        RECT 395.100 210.150 396.900 211.950 ;
        RECT 410.250 210.150 412.050 211.950 ;
        RECT 289.200 205.500 294.900 206.400 ;
        RECT 287.100 198.600 288.900 204.600 ;
        RECT 290.100 198.000 291.900 204.600 ;
        RECT 293.700 201.600 294.900 205.500 ;
        RECT 305.700 204.600 306.900 206.700 ;
        RECT 293.100 198.600 294.900 201.600 ;
        RECT 305.100 198.600 306.900 204.600 ;
        RECT 308.100 203.700 315.900 205.050 ;
        RECT 326.700 204.600 327.900 206.700 ;
        RECT 347.700 205.800 351.900 206.700 ;
        RECT 308.100 198.600 309.900 203.700 ;
        RECT 311.100 198.000 312.900 202.800 ;
        RECT 314.100 198.600 315.900 203.700 ;
        RECT 326.100 198.600 327.900 204.600 ;
        RECT 329.100 203.700 336.900 205.050 ;
        RECT 329.100 198.600 330.900 203.700 ;
        RECT 332.100 198.000 333.900 202.800 ;
        RECT 335.100 198.600 336.900 203.700 ;
        RECT 347.700 198.600 349.500 205.800 ;
        RECT 352.800 198.000 354.600 204.600 ;
        RECT 370.500 198.600 372.300 207.000 ;
        RECT 377.100 198.000 378.900 207.600 ;
        RECT 389.700 206.700 393.300 207.600 ;
        RECT 413.100 206.700 414.300 211.950 ;
        RECT 416.100 210.150 417.900 211.950 ;
        RECT 428.250 210.150 430.050 211.950 ;
        RECT 431.100 206.700 432.300 211.950 ;
        RECT 434.100 210.150 435.900 211.950 ;
        RECT 446.100 210.150 447.900 211.950 ;
        RECT 449.100 207.600 450.300 211.950 ;
        RECT 452.100 210.150 453.900 211.950 ;
        RECT 467.100 210.150 468.900 211.950 ;
        RECT 473.100 210.150 474.900 211.950 ;
        RECT 476.100 208.200 477.000 211.950 ;
        RECT 488.100 210.150 489.900 211.950 ;
        RECT 446.700 206.700 450.300 207.600 ;
        RECT 389.700 204.600 390.900 206.700 ;
        RECT 413.100 205.800 417.300 206.700 ;
        RECT 431.100 205.800 435.300 206.700 ;
        RECT 389.100 198.600 390.900 204.600 ;
        RECT 392.100 203.700 399.900 205.050 ;
        RECT 392.100 198.600 393.900 203.700 ;
        RECT 395.100 198.000 396.900 202.800 ;
        RECT 398.100 198.600 399.900 203.700 ;
        RECT 410.400 198.000 412.200 204.600 ;
        RECT 415.500 198.600 417.300 205.800 ;
        RECT 428.400 198.000 430.200 204.600 ;
        RECT 433.500 198.600 435.300 205.800 ;
        RECT 446.700 204.600 447.900 206.700 ;
        RECT 446.100 198.600 447.900 204.600 ;
        RECT 449.100 203.700 456.900 205.050 ;
        RECT 449.100 198.600 450.900 203.700 ;
        RECT 452.100 198.000 453.900 202.800 ;
        RECT 455.100 198.600 456.900 203.700 ;
        RECT 467.100 198.000 468.900 207.600 ;
        RECT 473.700 207.000 477.000 208.200 ;
        RECT 473.700 198.600 475.500 207.000 ;
        RECT 491.700 206.700 492.900 211.950 ;
        RECT 493.950 210.150 495.750 211.950 ;
        RECT 509.100 210.150 510.900 211.950 ;
        RECT 512.700 206.700 513.900 211.950 ;
        RECT 514.950 210.150 516.750 211.950 ;
        RECT 488.700 205.800 492.900 206.700 ;
        RECT 509.700 205.800 513.900 206.700 ;
        RECT 488.700 198.600 490.500 205.800 ;
        RECT 493.800 198.000 495.600 204.600 ;
        RECT 509.700 198.600 511.500 205.800 ;
        RECT 527.700 204.600 528.600 211.950 ;
        RECT 534.000 207.300 534.900 227.400 ;
        RECT 548.100 220.500 549.300 227.400 ;
        RECT 551.100 223.200 552.900 234.000 ;
        RECT 554.100 221.400 555.900 233.400 ;
        RECT 566.100 221.400 567.900 233.400 ;
        RECT 569.100 222.000 570.900 234.000 ;
        RECT 572.100 227.400 573.900 233.400 ;
        RECT 575.100 227.400 576.900 234.000 ;
        RECT 577.950 231.450 580.050 232.050 ;
        RECT 583.950 231.450 586.050 232.050 ;
        RECT 577.950 230.550 586.050 231.450 ;
        RECT 577.950 229.950 580.050 230.550 ;
        RECT 583.950 229.950 586.050 230.550 ;
        RECT 548.100 219.600 553.800 220.500 ;
        RECT 552.000 218.700 553.800 219.600 ;
        RECT 548.400 214.050 550.200 215.850 ;
        RECT 535.800 211.950 537.900 214.050 ;
        RECT 548.400 211.950 550.500 214.050 ;
        RECT 535.950 210.150 537.750 211.950 ;
        RECT 552.000 207.300 552.900 218.700 ;
        RECT 554.700 214.050 555.900 221.400 ;
        RECT 566.700 214.050 567.600 221.400 ;
        RECT 570.000 214.050 571.800 215.850 ;
        RECT 553.800 211.950 555.900 214.050 ;
        RECT 566.100 211.950 568.200 214.050 ;
        RECT 569.400 211.950 571.500 214.050 ;
        RECT 529.500 206.400 537.900 207.300 ;
        RECT 552.000 206.400 553.800 207.300 ;
        RECT 529.500 205.500 531.300 206.400 ;
        RECT 514.800 198.000 516.600 204.600 ;
        RECT 527.700 202.800 530.400 204.600 ;
        RECT 528.600 198.600 530.400 202.800 ;
        RECT 531.600 198.000 533.400 204.600 ;
        RECT 536.100 198.600 537.900 206.400 ;
        RECT 548.100 205.500 553.800 206.400 ;
        RECT 548.100 201.600 549.300 205.500 ;
        RECT 554.700 204.600 555.900 211.950 ;
        RECT 548.100 198.600 549.900 201.600 ;
        RECT 551.100 198.000 552.900 204.600 ;
        RECT 554.100 198.600 555.900 204.600 ;
        RECT 566.700 204.600 567.600 211.950 ;
        RECT 573.000 207.300 573.900 227.400 ;
        RECT 587.100 221.400 588.900 234.000 ;
        RECT 590.100 221.400 591.900 233.400 ;
        RECT 602.400 221.400 604.200 234.000 ;
        RECT 607.500 222.900 609.300 233.400 ;
        RECT 610.500 227.400 612.300 234.000 ;
        RECT 610.200 224.100 612.000 225.900 ;
        RECT 607.500 221.400 609.900 222.900 ;
        RECT 623.100 221.400 624.900 233.400 ;
        RECT 626.100 221.400 627.900 234.000 ;
        RECT 641.400 221.400 643.200 234.000 ;
        RECT 646.500 222.900 648.300 233.400 ;
        RECT 649.500 227.400 651.300 234.000 ;
        RECT 662.100 227.400 663.900 234.000 ;
        RECT 665.100 227.400 666.900 233.400 ;
        RECT 668.100 227.400 669.900 234.000 ;
        RECT 680.100 227.400 681.900 234.000 ;
        RECT 683.100 227.400 684.900 233.400 ;
        RECT 686.100 227.400 687.900 234.000 ;
        RECT 649.200 224.100 651.000 225.900 ;
        RECT 646.500 221.400 648.900 222.900 ;
        RECT 590.100 214.050 591.300 221.400 ;
        RECT 602.100 214.050 603.900 215.850 ;
        RECT 608.700 214.050 609.900 221.400 ;
        RECT 610.950 219.450 615.000 220.050 ;
        RECT 610.950 217.950 615.450 219.450 ;
        RECT 614.550 216.450 615.450 217.950 ;
        RECT 614.550 215.550 618.450 216.450 ;
        RECT 574.800 211.950 576.900 214.050 ;
        RECT 586.950 211.950 589.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 574.950 210.150 576.750 211.950 ;
        RECT 587.100 210.150 588.900 211.950 ;
        RECT 568.500 206.400 576.900 207.300 ;
        RECT 568.500 205.500 570.300 206.400 ;
        RECT 566.700 202.800 569.400 204.600 ;
        RECT 567.600 198.600 569.400 202.800 ;
        RECT 570.600 198.000 572.400 204.600 ;
        RECT 575.100 198.600 576.900 206.400 ;
        RECT 590.100 204.600 591.300 211.950 ;
        RECT 605.100 210.150 606.900 211.950 ;
        RECT 608.700 207.600 609.900 211.950 ;
        RECT 611.100 210.150 612.900 211.950 ;
        RECT 617.550 211.050 618.450 215.550 ;
        RECT 623.700 214.050 624.900 221.400 ;
        RECT 641.100 214.050 642.900 215.850 ;
        RECT 647.700 214.050 648.900 221.400 ;
        RECT 649.950 222.450 652.050 223.050 ;
        RECT 661.950 222.450 664.050 223.050 ;
        RECT 649.950 221.550 664.050 222.450 ;
        RECT 649.950 220.950 652.050 221.550 ;
        RECT 661.950 220.950 664.050 221.550 ;
        RECT 665.100 214.050 666.300 227.400 ;
        RECT 683.100 214.050 684.300 227.400 ;
        RECT 698.400 221.400 700.200 234.000 ;
        RECT 703.500 222.900 705.300 233.400 ;
        RECT 706.500 227.400 708.300 234.000 ;
        RECT 706.200 224.100 708.000 225.900 ;
        RECT 703.500 221.400 705.900 222.900 ;
        RECT 719.100 222.600 720.900 233.400 ;
        RECT 722.100 223.500 723.900 234.000 ;
        RECT 719.100 221.400 723.900 222.600 ;
        RECT 698.100 214.050 699.900 215.850 ;
        RECT 704.700 214.050 705.900 221.400 ;
        RECT 721.800 220.500 723.900 221.400 ;
        RECT 726.600 221.400 728.400 233.400 ;
        RECT 731.100 223.500 732.900 234.000 ;
        RECT 734.100 222.300 735.900 233.400 ;
        RECT 731.400 221.400 735.900 222.300 ;
        RECT 746.100 221.400 747.900 233.400 ;
        RECT 750.600 221.400 752.400 234.000 ;
        RECT 753.600 222.900 755.400 233.400 ;
        RECT 753.600 221.400 756.000 222.900 ;
        RECT 767.100 222.600 768.900 233.400 ;
        RECT 770.100 223.500 771.900 234.000 ;
        RECT 773.100 232.500 780.900 233.400 ;
        RECT 773.100 222.600 774.900 232.500 ;
        RECT 767.100 221.700 774.900 222.600 ;
        RECT 726.600 220.050 727.800 221.400 ;
        RECT 726.300 219.000 727.800 220.050 ;
        RECT 731.400 219.300 733.500 221.400 ;
        RECT 746.100 219.900 747.300 221.400 ;
        RECT 726.300 217.050 727.200 219.000 ;
        RECT 746.100 218.700 753.900 219.900 ;
        RECT 752.100 218.100 753.900 218.700 ;
        RECT 719.400 214.050 721.200 215.850 ;
        RECT 725.100 214.950 727.200 217.050 ;
        RECT 728.100 217.500 730.200 217.800 ;
        RECT 728.100 215.700 732.000 217.500 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 625.950 211.950 628.050 214.050 ;
        RECT 640.950 211.950 643.050 214.050 ;
        RECT 643.950 211.950 646.050 214.050 ;
        RECT 646.950 211.950 649.050 214.050 ;
        RECT 649.950 211.950 652.050 214.050 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 697.950 211.950 700.050 214.050 ;
        RECT 700.950 211.950 703.050 214.050 ;
        RECT 703.950 211.950 706.050 214.050 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 719.100 211.950 721.200 214.050 ;
        RECT 725.700 214.800 727.200 214.950 ;
        RECT 725.700 213.900 728.100 214.800 ;
        RECT 617.550 209.550 622.050 211.050 ;
        RECT 618.000 208.950 622.050 209.550 ;
        RECT 608.700 206.700 612.300 207.600 ;
        RECT 587.100 198.000 588.900 204.600 ;
        RECT 590.100 198.600 591.900 204.600 ;
        RECT 602.100 203.700 609.900 205.050 ;
        RECT 602.100 198.600 603.900 203.700 ;
        RECT 605.100 198.000 606.900 202.800 ;
        RECT 608.100 198.600 609.900 203.700 ;
        RECT 611.100 204.600 612.300 206.700 ;
        RECT 623.700 204.600 624.900 211.950 ;
        RECT 626.100 210.150 627.900 211.950 ;
        RECT 644.100 210.150 645.900 211.950 ;
        RECT 647.700 207.600 648.900 211.950 ;
        RECT 650.100 210.150 651.900 211.950 ;
        RECT 662.250 210.150 664.050 211.950 ;
        RECT 647.700 206.700 651.300 207.600 ;
        RECT 611.100 198.600 612.900 204.600 ;
        RECT 623.100 198.600 624.900 204.600 ;
        RECT 626.100 198.000 627.900 204.600 ;
        RECT 628.950 201.450 631.050 202.050 ;
        RECT 637.950 201.450 640.050 205.050 ;
        RECT 628.950 201.000 640.050 201.450 ;
        RECT 641.100 203.700 648.900 205.050 ;
        RECT 628.950 200.550 639.450 201.000 ;
        RECT 628.950 199.950 631.050 200.550 ;
        RECT 641.100 198.600 642.900 203.700 ;
        RECT 644.100 198.000 645.900 202.800 ;
        RECT 647.100 198.600 648.900 203.700 ;
        RECT 650.100 204.600 651.300 206.700 ;
        RECT 665.100 206.700 666.300 211.950 ;
        RECT 668.100 210.150 669.900 211.950 ;
        RECT 680.250 210.150 682.050 211.950 ;
        RECT 683.100 206.700 684.300 211.950 ;
        RECT 686.100 210.150 687.900 211.950 ;
        RECT 701.100 210.150 702.900 211.950 ;
        RECT 704.700 207.600 705.900 211.950 ;
        RECT 707.100 210.150 708.900 211.950 ;
        RECT 723.900 211.200 725.700 213.000 ;
        RECT 723.900 209.100 726.000 211.200 ;
        RECT 726.900 208.200 728.100 213.900 ;
        RECT 729.000 214.050 730.800 214.500 ;
        RECT 750.000 214.050 751.800 215.850 ;
        RECT 729.000 212.700 735.900 214.050 ;
        RECT 733.800 211.950 735.900 212.700 ;
        RECT 746.100 211.950 748.200 214.050 ;
        RECT 749.400 211.950 751.500 214.050 ;
        RECT 704.700 206.700 708.300 207.600 ;
        RECT 665.100 205.800 669.300 206.700 ;
        RECT 683.100 205.800 687.300 206.700 ;
        RECT 650.100 198.600 651.900 204.600 ;
        RECT 662.400 198.000 664.200 204.600 ;
        RECT 667.500 198.600 669.300 205.800 ;
        RECT 680.400 198.000 682.200 204.600 ;
        RECT 685.500 198.600 687.300 205.800 ;
        RECT 698.100 203.700 705.900 205.050 ;
        RECT 698.100 198.600 699.900 203.700 ;
        RECT 701.100 198.000 702.900 202.800 ;
        RECT 704.100 198.600 705.900 203.700 ;
        RECT 707.100 204.600 708.300 206.700 ;
        RECT 721.800 205.500 723.900 206.700 ;
        RECT 725.100 206.100 728.100 208.200 ;
        RECT 729.000 209.400 730.800 211.200 ;
        RECT 733.800 210.150 735.600 211.950 ;
        RECT 746.400 210.150 748.200 211.950 ;
        RECT 729.000 207.300 731.100 209.400 ;
        RECT 752.700 207.600 753.600 218.100 ;
        RECT 754.800 214.050 756.000 221.400 ;
        RECT 776.100 220.500 777.900 231.600 ;
        RECT 779.100 221.400 780.900 232.500 ;
        RECT 794.100 227.400 795.900 234.000 ;
        RECT 797.100 227.400 798.900 233.400 ;
        RECT 773.100 219.600 777.900 220.500 ;
        RECT 762.000 216.450 766.050 217.050 ;
        RECT 761.550 214.950 766.050 216.450 ;
        RECT 754.800 211.950 756.900 214.050 ;
        RECT 729.000 206.400 735.300 207.300 ;
        RECT 752.700 206.700 754.800 207.600 ;
        RECT 719.100 204.600 723.900 205.500 ;
        RECT 726.900 204.600 728.100 206.100 ;
        RECT 734.100 204.600 735.300 206.400 ;
        RECT 749.400 205.800 754.800 206.700 ;
        RECT 707.100 198.600 708.900 204.600 ;
        RECT 719.100 198.600 720.900 204.600 ;
        RECT 722.100 198.000 723.900 203.700 ;
        RECT 726.600 198.600 728.400 204.600 ;
        RECT 731.100 198.000 732.900 203.700 ;
        RECT 734.100 198.600 735.900 204.600 ;
        RECT 749.400 201.600 750.300 205.800 ;
        RECT 756.000 204.600 756.900 211.950 ;
        RECT 761.550 211.050 762.450 214.950 ;
        RECT 770.250 214.050 772.050 215.850 ;
        RECT 773.100 214.050 774.000 219.600 ;
        RECT 776.100 214.050 777.900 215.850 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 772.950 211.950 775.050 214.050 ;
        RECT 775.950 211.950 778.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 794.100 211.950 796.200 214.050 ;
        RECT 761.550 209.550 766.050 211.050 ;
        RECT 767.250 210.150 769.050 211.950 ;
        RECT 762.000 208.950 766.050 209.550 ;
        RECT 773.100 204.600 774.300 211.950 ;
        RECT 779.100 210.150 780.900 211.950 ;
        RECT 794.250 210.150 796.050 211.950 ;
        RECT 778.950 207.450 781.050 208.050 ;
        RECT 784.950 207.450 787.050 208.050 ;
        RECT 778.950 206.550 787.050 207.450 ;
        RECT 797.100 207.300 798.000 227.400 ;
        RECT 800.100 222.000 801.900 234.000 ;
        RECT 803.100 221.400 804.900 233.400 ;
        RECT 815.100 222.300 816.900 233.400 ;
        RECT 818.100 223.200 819.900 234.000 ;
        RECT 821.100 222.300 822.900 233.400 ;
        RECT 815.100 221.400 822.900 222.300 ;
        RECT 824.100 221.400 825.900 233.400 ;
        RECT 836.100 222.600 837.900 233.400 ;
        RECT 839.100 223.500 840.900 234.000 ;
        RECT 842.100 232.500 849.900 233.400 ;
        RECT 842.100 222.600 843.900 232.500 ;
        RECT 836.100 221.700 843.900 222.600 ;
        RECT 799.200 214.050 801.000 215.850 ;
        RECT 803.400 214.050 804.300 221.400 ;
        RECT 818.250 214.050 820.050 215.850 ;
        RECT 824.700 214.050 825.600 221.400 ;
        RECT 845.100 220.500 846.900 231.600 ;
        RECT 848.100 221.400 849.900 232.500 ;
        RECT 860.100 227.400 861.900 234.000 ;
        RECT 863.100 227.400 864.900 233.400 ;
        RECT 866.100 228.000 867.900 234.000 ;
        RECT 863.400 227.100 864.900 227.400 ;
        RECT 869.100 227.400 870.900 233.400 ;
        RECT 869.100 227.100 870.000 227.400 ;
        RECT 863.400 226.200 870.000 227.100 ;
        RECT 853.950 222.450 856.050 223.050 ;
        RECT 865.950 222.450 868.050 223.050 ;
        RECT 853.950 221.550 868.050 222.450 ;
        RECT 853.950 220.950 856.050 221.550 ;
        RECT 865.950 220.950 868.050 221.550 ;
        RECT 842.100 219.600 846.900 220.500 ;
        RECT 831.000 216.450 835.050 217.050 ;
        RECT 830.550 214.950 835.050 216.450 ;
        RECT 799.500 211.950 801.600 214.050 ;
        RECT 802.800 211.950 804.900 214.050 ;
        RECT 814.950 211.950 817.050 214.050 ;
        RECT 817.950 211.950 820.050 214.050 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 778.950 205.950 781.050 206.550 ;
        RECT 784.950 205.950 787.050 206.550 ;
        RECT 794.100 206.400 802.500 207.300 ;
        RECT 746.100 198.600 747.900 201.600 ;
        RECT 749.100 198.600 750.900 201.600 ;
        RECT 746.100 198.000 747.300 198.600 ;
        RECT 752.100 198.000 753.900 204.000 ;
        RECT 755.100 198.600 756.900 204.600 ;
        RECT 767.700 198.000 769.500 204.600 ;
        RECT 772.200 198.600 774.000 204.600 ;
        RECT 776.700 198.000 778.500 204.600 ;
        RECT 794.100 198.600 795.900 206.400 ;
        RECT 800.700 205.500 802.500 206.400 ;
        RECT 803.400 204.600 804.300 211.950 ;
        RECT 815.100 210.150 816.900 211.950 ;
        RECT 821.250 210.150 823.050 211.950 ;
        RECT 808.950 207.450 811.050 208.050 ;
        RECT 817.950 207.450 820.050 207.750 ;
        RECT 808.950 206.550 820.050 207.450 ;
        RECT 808.950 205.950 811.050 206.550 ;
        RECT 817.950 205.650 820.050 206.550 ;
        RECT 824.700 204.600 825.600 211.950 ;
        RECT 830.550 211.050 831.450 214.950 ;
        RECT 839.250 214.050 841.050 215.850 ;
        RECT 842.100 214.050 843.000 219.600 ;
        RECT 862.950 219.450 865.050 220.050 ;
        RECT 854.550 218.550 865.050 219.450 ;
        RECT 845.100 214.050 846.900 215.850 ;
        RECT 835.950 211.950 838.050 214.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 826.950 209.550 831.450 211.050 ;
        RECT 836.250 210.150 838.050 211.950 ;
        RECT 826.950 208.950 831.000 209.550 ;
        RECT 842.100 204.600 843.300 211.950 ;
        RECT 848.100 210.150 849.900 211.950 ;
        RECT 854.550 211.050 855.450 218.550 ;
        RECT 862.950 217.950 865.050 218.550 ;
        RECT 863.100 214.050 864.900 215.850 ;
        RECT 869.100 214.050 870.000 226.200 ;
        RECT 859.950 211.950 862.050 214.050 ;
        RECT 862.950 211.950 865.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 854.550 209.550 859.050 211.050 ;
        RECT 860.100 210.150 861.900 211.950 ;
        RECT 866.100 210.150 867.900 211.950 ;
        RECT 855.000 208.950 859.050 209.550 ;
        RECT 869.100 208.200 870.000 211.950 ;
        RECT 798.600 198.000 800.400 204.600 ;
        RECT 801.600 202.800 804.300 204.600 ;
        RECT 801.600 198.600 803.400 202.800 ;
        RECT 816.000 198.000 817.800 204.600 ;
        RECT 820.500 203.400 825.600 204.600 ;
        RECT 820.500 198.600 822.300 203.400 ;
        RECT 823.500 198.000 825.300 201.600 ;
        RECT 836.700 198.000 838.500 204.600 ;
        RECT 841.200 198.600 843.000 204.600 ;
        RECT 845.700 198.000 847.500 204.600 ;
        RECT 860.100 198.000 861.900 207.600 ;
        RECT 866.700 207.000 870.000 208.200 ;
        RECT 866.700 198.600 868.500 207.000 ;
        RECT 11.700 187.200 13.500 194.400 ;
        RECT 16.800 188.400 18.600 195.000 ;
        RECT 32.700 188.400 34.500 195.000 ;
        RECT 37.200 188.400 39.000 194.400 ;
        RECT 41.700 188.400 43.500 195.000 ;
        RECT 11.700 186.300 15.900 187.200 ;
        RECT 11.100 181.050 12.900 182.850 ;
        RECT 14.700 181.050 15.900 186.300 ;
        RECT 22.950 186.450 25.050 187.050 ;
        RECT 34.950 186.450 37.050 187.050 ;
        RECT 22.950 185.550 37.050 186.450 ;
        RECT 22.950 184.950 25.050 185.550 ;
        RECT 34.950 184.950 37.050 185.550 ;
        RECT 16.950 181.050 18.750 182.850 ;
        RECT 32.250 181.050 34.050 182.850 ;
        RECT 38.100 181.050 39.300 188.400 ;
        RECT 58.500 186.000 60.300 194.400 ;
        RECT 57.000 184.800 60.300 186.000 ;
        RECT 65.100 185.400 66.900 195.000 ;
        RECT 80.100 191.400 81.900 195.000 ;
        RECT 83.100 191.400 84.900 194.400 ;
        RECT 44.100 181.050 45.900 182.850 ;
        RECT 57.000 181.050 57.900 184.800 ;
        RECT 59.100 181.050 60.900 182.850 ;
        RECT 65.100 181.050 66.900 182.850 ;
        RECT 83.100 181.050 84.300 191.400 ;
        RECT 95.100 188.400 96.900 194.400 ;
        RECT 95.700 186.300 96.900 188.400 ;
        RECT 98.100 189.300 99.900 194.400 ;
        RECT 101.100 190.200 102.900 195.000 ;
        RECT 104.100 189.300 105.900 194.400 ;
        RECT 116.700 191.400 118.500 195.000 ;
        RECT 119.700 189.600 121.500 194.400 ;
        RECT 98.100 187.950 105.900 189.300 ;
        RECT 116.400 188.400 121.500 189.600 ;
        RECT 124.200 188.400 126.000 195.000 ;
        RECT 137.100 191.400 138.900 194.400 ;
        RECT 140.100 191.400 141.900 195.000 ;
        RECT 152.100 191.400 153.900 194.400 ;
        RECT 155.100 191.400 156.900 195.000 ;
        RECT 95.700 185.400 99.300 186.300 ;
        RECT 95.100 181.050 96.900 182.850 ;
        RECT 98.100 181.050 99.300 185.400 ;
        RECT 101.100 181.050 102.900 182.850 ;
        RECT 116.400 181.050 117.300 188.400 ;
        RECT 124.950 186.450 127.050 187.050 ;
        RECT 130.950 186.450 133.050 187.050 ;
        RECT 124.950 185.550 133.050 186.450 ;
        RECT 124.950 184.950 127.050 185.550 ;
        RECT 130.950 184.950 133.050 185.550 ;
        RECT 118.950 181.050 120.750 182.850 ;
        RECT 125.100 181.050 126.900 182.850 ;
        RECT 137.700 181.050 138.900 191.400 ;
        RECT 152.700 181.050 153.900 191.400 ;
        RECT 167.100 186.600 168.900 194.400 ;
        RECT 171.600 188.400 173.400 195.000 ;
        RECT 174.600 190.200 176.400 194.400 ;
        RECT 174.600 188.400 177.300 190.200 ;
        RECT 190.500 188.400 192.300 195.000 ;
        RECT 195.000 188.400 196.800 194.400 ;
        RECT 199.500 188.400 201.300 195.000 ;
        RECT 212.700 188.400 214.500 195.000 ;
        RECT 217.200 188.400 219.000 194.400 ;
        RECT 221.700 188.400 223.500 195.000 ;
        RECT 236.400 188.400 238.200 195.000 ;
        RECT 173.700 186.600 175.500 187.500 ;
        RECT 167.100 185.700 175.500 186.600 ;
        RECT 167.250 181.050 169.050 182.850 ;
        RECT 10.950 178.950 13.050 181.050 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 31.950 178.950 34.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 167.100 178.950 169.200 181.050 ;
        RECT 14.700 165.600 15.900 178.950 ;
        RECT 35.250 177.150 37.050 178.950 ;
        RECT 38.100 173.400 39.000 178.950 ;
        RECT 41.100 177.150 42.900 178.950 ;
        RECT 38.100 172.500 42.900 173.400 ;
        RECT 32.100 170.400 39.900 171.300 ;
        RECT 11.100 159.000 12.900 165.600 ;
        RECT 14.100 159.600 15.900 165.600 ;
        RECT 17.100 159.000 18.900 165.600 ;
        RECT 32.100 159.600 33.900 170.400 ;
        RECT 35.100 159.000 36.900 169.500 ;
        RECT 38.100 160.500 39.900 170.400 ;
        RECT 41.100 161.400 42.900 172.500 ;
        RECT 44.100 160.500 45.900 171.600 ;
        RECT 57.000 166.800 57.900 178.950 ;
        RECT 62.100 177.150 63.900 178.950 ;
        RECT 80.100 177.150 81.900 178.950 ;
        RECT 58.950 171.450 61.050 172.050 ;
        RECT 64.950 171.450 67.050 171.900 ;
        RECT 58.950 170.550 67.050 171.450 ;
        RECT 58.950 169.950 61.050 170.550 ;
        RECT 64.950 169.800 67.050 170.550 ;
        RECT 57.000 165.900 63.600 166.800 ;
        RECT 57.000 165.600 57.900 165.900 ;
        RECT 38.100 159.600 45.900 160.500 ;
        RECT 56.100 159.600 57.900 165.600 ;
        RECT 62.100 165.600 63.600 165.900 ;
        RECT 83.100 165.600 84.300 178.950 ;
        RECT 98.100 171.600 99.300 178.950 ;
        RECT 104.100 177.150 105.900 178.950 ;
        RECT 116.400 171.600 117.300 178.950 ;
        RECT 121.950 177.150 123.750 178.950 ;
        RECT 118.950 174.450 121.050 175.050 ;
        RECT 130.950 174.450 133.050 175.050 ;
        RECT 118.950 173.550 133.050 174.450 ;
        RECT 118.950 172.950 121.050 173.550 ;
        RECT 130.950 172.950 133.050 173.550 ;
        RECT 98.100 170.100 100.500 171.600 ;
        RECT 96.000 167.100 97.800 168.900 ;
        RECT 59.100 159.000 60.900 165.000 ;
        RECT 62.100 159.600 63.900 165.600 ;
        RECT 65.100 159.000 66.900 165.600 ;
        RECT 80.100 159.000 81.900 165.600 ;
        RECT 83.100 159.600 84.900 165.600 ;
        RECT 95.700 159.000 97.500 165.600 ;
        RECT 98.700 159.600 100.500 170.100 ;
        RECT 103.800 159.000 105.600 171.600 ;
        RECT 116.100 159.600 117.900 171.600 ;
        RECT 119.100 170.700 126.900 171.600 ;
        RECT 119.100 159.600 120.900 170.700 ;
        RECT 122.100 159.000 123.900 169.800 ;
        RECT 125.100 159.600 126.900 170.700 ;
        RECT 137.700 165.600 138.900 178.950 ;
        RECT 140.100 177.150 141.900 178.950 ;
        RECT 152.700 165.600 153.900 178.950 ;
        RECT 155.100 177.150 156.900 178.950 ;
        RECT 170.100 165.600 171.000 185.700 ;
        RECT 176.400 181.050 177.300 188.400 ;
        RECT 188.100 181.050 189.900 182.850 ;
        RECT 194.700 181.050 195.900 188.400 ;
        RECT 196.950 186.450 199.050 187.050 ;
        RECT 208.950 186.450 211.050 187.050 ;
        RECT 196.950 185.550 211.050 186.450 ;
        RECT 196.950 184.950 199.050 185.550 ;
        RECT 208.950 184.950 211.050 185.550 ;
        RECT 199.950 181.050 201.750 182.850 ;
        RECT 212.250 181.050 214.050 182.850 ;
        RECT 218.100 181.050 219.300 188.400 ;
        RECT 241.500 187.200 243.300 194.400 ;
        RECT 220.950 186.450 223.050 186.900 ;
        RECT 229.950 186.450 232.050 187.050 ;
        RECT 220.950 185.550 232.050 186.450 ;
        RECT 220.950 184.800 223.050 185.550 ;
        RECT 229.950 184.950 232.050 185.550 ;
        RECT 239.100 186.300 243.300 187.200 ;
        RECT 257.100 188.400 258.900 194.400 ;
        RECT 260.100 188.400 261.900 195.000 ;
        RECT 263.100 191.400 264.900 194.400 ;
        RECT 224.100 181.050 225.900 182.850 ;
        RECT 236.250 181.050 238.050 182.850 ;
        RECT 239.100 181.050 240.300 186.300 ;
        RECT 242.100 181.050 243.900 182.850 ;
        RECT 257.100 181.050 258.300 188.400 ;
        RECT 263.700 187.500 264.900 191.400 ;
        RECT 278.100 188.400 279.900 194.400 ;
        RECT 281.100 189.300 282.900 195.000 ;
        RECT 285.600 188.400 287.400 194.400 ;
        RECT 290.100 189.300 291.900 195.000 ;
        RECT 293.100 188.400 294.900 194.400 ;
        RECT 306.600 190.200 308.400 194.400 ;
        RECT 259.200 186.600 264.900 187.500 ;
        RECT 278.700 186.600 279.900 188.400 ;
        RECT 285.900 186.900 287.100 188.400 ;
        RECT 290.100 187.500 294.900 188.400 ;
        RECT 305.700 188.400 308.400 190.200 ;
        RECT 309.600 188.400 311.400 195.000 ;
        RECT 259.200 185.700 261.000 186.600 ;
        RECT 278.700 185.700 285.000 186.600 ;
        RECT 172.500 178.950 174.600 181.050 ;
        RECT 175.800 178.950 177.900 181.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 257.100 178.950 259.200 181.050 ;
        RECT 172.200 177.150 174.000 178.950 ;
        RECT 176.400 171.600 177.300 178.950 ;
        RECT 191.100 177.150 192.900 178.950 ;
        RECT 195.000 173.400 195.900 178.950 ;
        RECT 196.950 177.150 198.750 178.950 ;
        RECT 215.250 177.150 217.050 178.950 ;
        RECT 191.100 172.500 195.900 173.400 ;
        RECT 218.100 173.400 219.000 178.950 ;
        RECT 221.100 177.150 222.900 178.950 ;
        RECT 223.950 174.450 226.050 175.050 ;
        RECT 235.950 174.450 238.050 175.050 ;
        RECT 223.950 173.550 238.050 174.450 ;
        RECT 218.100 172.500 222.900 173.400 ;
        RECT 223.950 172.950 226.050 173.550 ;
        RECT 235.950 172.950 238.050 173.550 ;
        RECT 137.100 159.600 138.900 165.600 ;
        RECT 140.100 159.000 141.900 165.600 ;
        RECT 152.100 159.600 153.900 165.600 ;
        RECT 155.100 159.000 156.900 165.600 ;
        RECT 167.100 159.000 168.900 165.600 ;
        RECT 170.100 159.600 171.900 165.600 ;
        RECT 173.100 159.000 174.900 171.000 ;
        RECT 176.100 159.600 177.900 171.600 ;
        RECT 188.100 160.500 189.900 171.600 ;
        RECT 191.100 161.400 192.900 172.500 ;
        RECT 194.100 170.400 201.900 171.300 ;
        RECT 194.100 160.500 195.900 170.400 ;
        RECT 188.100 159.600 195.900 160.500 ;
        RECT 197.100 159.000 198.900 169.500 ;
        RECT 200.100 159.600 201.900 170.400 ;
        RECT 212.100 170.400 219.900 171.300 ;
        RECT 212.100 159.600 213.900 170.400 ;
        RECT 215.100 159.000 216.900 169.500 ;
        RECT 218.100 160.500 219.900 170.400 ;
        RECT 221.100 161.400 222.900 172.500 ;
        RECT 224.100 160.500 225.900 171.600 ;
        RECT 239.100 165.600 240.300 178.950 ;
        RECT 257.100 171.600 258.300 178.950 ;
        RECT 260.100 174.300 261.000 185.700 ;
        RECT 282.900 183.600 285.000 185.700 ;
        RECT 278.400 181.050 280.200 182.850 ;
        RECT 283.200 181.800 285.000 183.600 ;
        RECT 285.900 184.800 288.900 186.900 ;
        RECT 290.100 186.300 292.200 187.500 ;
        RECT 262.500 178.950 264.600 181.050 ;
        RECT 278.100 180.300 280.200 181.050 ;
        RECT 278.100 178.950 285.000 180.300 ;
        RECT 262.800 177.150 264.600 178.950 ;
        RECT 283.200 178.500 285.000 178.950 ;
        RECT 285.900 179.100 287.100 184.800 ;
        RECT 288.000 181.800 290.100 183.900 ;
        RECT 288.300 180.000 290.100 181.800 ;
        RECT 305.700 181.050 306.600 188.400 ;
        RECT 307.500 186.600 309.300 187.500 ;
        RECT 314.100 186.600 315.900 194.400 ;
        RECT 307.500 185.700 315.900 186.600 ;
        RECT 326.700 187.200 328.500 194.400 ;
        RECT 331.800 188.400 333.600 195.000 ;
        RECT 344.100 189.300 345.900 194.400 ;
        RECT 347.100 190.200 348.900 195.000 ;
        RECT 350.100 189.300 351.900 194.400 ;
        RECT 344.100 187.950 351.900 189.300 ;
        RECT 353.100 188.400 354.900 194.400 ;
        RECT 365.100 191.400 366.900 194.400 ;
        RECT 326.700 186.300 330.900 187.200 ;
        RECT 285.900 178.200 288.300 179.100 ;
        RECT 286.800 178.050 288.300 178.200 ;
        RECT 292.800 178.950 294.900 181.050 ;
        RECT 305.100 178.950 307.200 181.050 ;
        RECT 308.400 178.950 310.500 181.050 ;
        RECT 282.000 175.500 285.900 177.300 ;
        RECT 283.800 175.200 285.900 175.500 ;
        RECT 286.800 175.950 288.900 178.050 ;
        RECT 292.800 177.150 294.600 178.950 ;
        RECT 259.200 173.400 261.000 174.300 ;
        RECT 286.800 174.000 287.700 175.950 ;
        RECT 259.200 172.500 264.900 173.400 ;
        RECT 218.100 159.600 225.900 160.500 ;
        RECT 236.100 159.000 237.900 165.600 ;
        RECT 239.100 159.600 240.900 165.600 ;
        RECT 242.100 159.000 243.900 165.600 ;
        RECT 257.100 159.600 258.900 171.600 ;
        RECT 260.100 159.000 261.900 169.800 ;
        RECT 263.700 165.600 264.900 172.500 ;
        RECT 280.500 171.600 282.600 173.700 ;
        RECT 286.200 172.950 287.700 174.000 ;
        RECT 286.200 171.600 287.400 172.950 ;
        RECT 263.100 159.600 264.900 165.600 ;
        RECT 278.100 170.700 282.600 171.600 ;
        RECT 278.100 159.600 279.900 170.700 ;
        RECT 281.100 159.000 282.900 169.500 ;
        RECT 285.600 159.600 287.400 171.600 ;
        RECT 290.100 171.600 292.200 172.500 ;
        RECT 305.700 171.600 306.600 178.950 ;
        RECT 309.000 177.150 310.800 178.950 ;
        RECT 290.100 170.400 294.900 171.600 ;
        RECT 290.100 159.000 291.900 169.500 ;
        RECT 293.100 159.600 294.900 170.400 ;
        RECT 305.100 159.600 306.900 171.600 ;
        RECT 308.100 159.000 309.900 171.000 ;
        RECT 312.000 165.600 312.900 185.700 ;
        RECT 321.000 183.450 325.050 184.050 ;
        RECT 313.950 181.050 315.750 182.850 ;
        RECT 320.550 181.950 325.050 183.450 ;
        RECT 313.800 178.950 315.900 181.050 ;
        RECT 320.550 177.450 321.450 181.950 ;
        RECT 326.100 181.050 327.900 182.850 ;
        RECT 329.700 181.050 330.900 186.300 ;
        RECT 340.950 183.450 343.050 187.050 ;
        RECT 353.100 186.300 354.300 188.400 ;
        RECT 365.100 187.500 366.300 191.400 ;
        RECT 368.100 188.400 369.900 195.000 ;
        RECT 371.100 188.400 372.900 194.400 ;
        RECT 365.100 186.600 370.800 187.500 ;
        RECT 338.550 183.000 343.050 183.450 ;
        RECT 350.700 185.400 354.300 186.300 ;
        RECT 369.000 185.700 370.800 186.600 ;
        RECT 331.950 181.050 333.750 182.850 ;
        RECT 338.550 182.550 342.450 183.000 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 320.550 176.550 324.450 177.450 ;
        RECT 323.550 175.050 324.450 176.550 ;
        RECT 313.950 174.450 316.050 175.050 ;
        RECT 323.550 174.450 328.050 175.050 ;
        RECT 313.950 173.550 328.050 174.450 ;
        RECT 313.950 172.950 316.050 173.550 ;
        RECT 324.000 172.950 328.050 173.550 ;
        RECT 329.700 165.600 330.900 178.950 ;
        RECT 338.550 178.050 339.450 182.550 ;
        RECT 347.100 181.050 348.900 182.850 ;
        RECT 350.700 181.050 351.900 185.400 ;
        RECT 353.100 181.050 354.900 182.850 ;
        RECT 343.950 178.950 346.050 181.050 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 365.400 178.950 367.500 181.050 ;
        RECT 334.950 176.550 339.450 178.050 ;
        RECT 344.100 177.150 345.900 178.950 ;
        RECT 334.950 175.950 339.000 176.550 ;
        RECT 350.700 171.600 351.900 178.950 ;
        RECT 365.400 177.150 367.200 178.950 ;
        RECT 352.950 174.450 355.050 175.050 ;
        RECT 361.950 174.450 364.050 175.050 ;
        RECT 352.950 173.550 364.050 174.450 ;
        RECT 352.950 172.950 355.050 173.550 ;
        RECT 361.950 172.950 364.050 173.550 ;
        RECT 369.000 174.300 369.900 185.700 ;
        RECT 371.700 181.050 372.900 188.400 ;
        RECT 370.800 178.950 372.900 181.050 ;
        RECT 369.000 173.400 370.800 174.300 ;
        RECT 311.100 159.600 312.900 165.600 ;
        RECT 314.100 159.000 315.900 165.600 ;
        RECT 326.100 159.000 327.900 165.600 ;
        RECT 329.100 159.600 330.900 165.600 ;
        RECT 332.100 159.000 333.900 165.600 ;
        RECT 344.400 159.000 346.200 171.600 ;
        RECT 349.500 170.100 351.900 171.600 ;
        RECT 365.100 172.500 370.800 173.400 ;
        RECT 349.500 159.600 351.300 170.100 ;
        RECT 352.200 167.100 354.000 168.900 ;
        RECT 365.100 165.600 366.300 172.500 ;
        RECT 371.700 171.600 372.900 178.950 ;
        RECT 352.500 159.000 354.300 165.600 ;
        RECT 365.100 159.600 366.900 165.600 ;
        RECT 368.100 159.000 369.900 169.800 ;
        RECT 371.100 159.600 372.900 171.600 ;
        RECT 383.100 188.400 384.900 194.400 ;
        RECT 386.100 188.400 387.900 195.000 ;
        RECT 389.100 191.400 390.900 194.400 ;
        RECT 383.100 181.050 384.300 188.400 ;
        RECT 389.700 187.500 390.900 191.400 ;
        RECT 385.200 186.600 390.900 187.500 ;
        RECT 401.100 191.400 402.900 194.400 ;
        RECT 401.100 187.500 402.300 191.400 ;
        RECT 404.100 188.400 405.900 195.000 ;
        RECT 407.100 188.400 408.900 194.400 ;
        RECT 401.100 186.600 406.800 187.500 ;
        RECT 385.200 185.700 387.000 186.600 ;
        RECT 383.100 178.950 385.200 181.050 ;
        RECT 383.100 171.600 384.300 178.950 ;
        RECT 386.100 174.300 387.000 185.700 ;
        RECT 405.000 185.700 406.800 186.600 ;
        RECT 388.500 178.950 390.600 181.050 ;
        RECT 388.800 177.150 390.600 178.950 ;
        RECT 401.400 178.950 403.500 181.050 ;
        RECT 401.400 177.150 403.200 178.950 ;
        RECT 385.200 173.400 387.000 174.300 ;
        RECT 405.000 174.300 405.900 185.700 ;
        RECT 407.700 181.050 408.900 188.400 ;
        RECT 419.100 191.400 420.900 194.400 ;
        RECT 419.100 187.500 420.300 191.400 ;
        RECT 422.100 188.400 423.900 195.000 ;
        RECT 425.100 188.400 426.900 194.400 ;
        RECT 419.100 186.600 424.800 187.500 ;
        RECT 423.000 185.700 424.800 186.600 ;
        RECT 406.800 178.950 408.900 181.050 ;
        RECT 405.000 173.400 406.800 174.300 ;
        RECT 385.200 172.500 390.900 173.400 ;
        RECT 383.100 159.600 384.900 171.600 ;
        RECT 386.100 159.000 387.900 169.800 ;
        RECT 389.700 165.600 390.900 172.500 ;
        RECT 389.100 159.600 390.900 165.600 ;
        RECT 401.100 172.500 406.800 173.400 ;
        RECT 401.100 165.600 402.300 172.500 ;
        RECT 407.700 171.600 408.900 178.950 ;
        RECT 419.400 178.950 421.500 181.050 ;
        RECT 419.400 177.150 421.200 178.950 ;
        RECT 423.000 174.300 423.900 185.700 ;
        RECT 425.700 181.050 426.900 188.400 ;
        RECT 437.700 187.200 439.500 194.400 ;
        RECT 442.800 188.400 444.600 195.000 ;
        RECT 437.700 186.300 441.900 187.200 ;
        RECT 437.100 181.050 438.900 182.850 ;
        RECT 440.700 181.050 441.900 186.300 ;
        RECT 455.100 186.600 456.900 194.400 ;
        RECT 459.600 188.400 461.400 195.000 ;
        RECT 462.600 190.200 464.400 194.400 ;
        RECT 462.600 188.400 465.300 190.200 ;
        RECT 461.700 186.600 463.500 187.500 ;
        RECT 455.100 185.700 463.500 186.600 ;
        RECT 442.950 181.050 444.750 182.850 ;
        RECT 455.250 181.050 457.050 182.850 ;
        RECT 424.800 178.950 426.900 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 439.950 178.950 442.050 181.050 ;
        RECT 442.950 178.950 445.050 181.050 ;
        RECT 455.100 178.950 457.200 181.050 ;
        RECT 423.000 173.400 424.800 174.300 ;
        RECT 401.100 159.600 402.900 165.600 ;
        RECT 404.100 159.000 405.900 169.800 ;
        RECT 407.100 159.600 408.900 171.600 ;
        RECT 419.100 172.500 424.800 173.400 ;
        RECT 419.100 165.600 420.300 172.500 ;
        RECT 425.700 171.600 426.900 178.950 ;
        RECT 419.100 159.600 420.900 165.600 ;
        RECT 422.100 159.000 423.900 169.800 ;
        RECT 425.100 159.600 426.900 171.600 ;
        RECT 440.700 165.600 441.900 178.950 ;
        RECT 458.100 165.600 459.000 185.700 ;
        RECT 464.400 181.050 465.300 188.400 ;
        RECT 476.700 187.200 478.500 194.400 ;
        RECT 481.800 188.400 483.600 195.000 ;
        RECT 497.100 188.400 498.900 194.400 ;
        RECT 476.700 186.300 480.900 187.200 ;
        RECT 476.100 181.050 477.900 182.850 ;
        RECT 479.700 181.050 480.900 186.300 ;
        RECT 497.700 186.300 498.900 188.400 ;
        RECT 500.100 189.300 501.900 194.400 ;
        RECT 503.100 190.200 504.900 195.000 ;
        RECT 506.100 189.300 507.900 194.400 ;
        RECT 500.100 187.950 507.900 189.300 ;
        RECT 497.700 185.400 501.300 186.300 ;
        RECT 523.500 186.000 525.300 194.400 ;
        RECT 481.950 181.050 483.750 182.850 ;
        RECT 497.100 181.050 498.900 182.850 ;
        RECT 500.100 181.050 501.300 185.400 ;
        RECT 522.000 184.800 525.300 186.000 ;
        RECT 530.100 185.400 531.900 195.000 ;
        RECT 544.500 188.400 546.300 195.000 ;
        RECT 549.000 188.400 550.800 194.400 ;
        RECT 553.500 188.400 555.300 195.000 ;
        RECT 503.100 181.050 504.900 182.850 ;
        RECT 522.000 181.050 522.900 184.800 ;
        RECT 524.100 181.050 525.900 182.850 ;
        RECT 530.100 181.050 531.900 182.850 ;
        RECT 542.100 181.050 543.900 182.850 ;
        RECT 548.700 181.050 549.900 188.400 ;
        RECT 566.700 187.200 568.500 194.400 ;
        RECT 571.800 188.400 573.600 195.000 ;
        RECT 584.100 189.300 585.900 194.400 ;
        RECT 587.100 190.200 588.900 195.000 ;
        RECT 590.100 189.300 591.900 194.400 ;
        RECT 584.100 187.950 591.900 189.300 ;
        RECT 593.100 188.400 594.900 194.400 ;
        RECT 606.000 188.400 607.800 195.000 ;
        RECT 610.500 189.600 612.300 194.400 ;
        RECT 613.500 191.400 615.300 195.000 ;
        RECT 627.600 190.200 629.400 194.400 ;
        RECT 610.500 188.400 615.600 189.600 ;
        RECT 566.700 186.300 570.900 187.200 ;
        RECT 593.100 186.300 594.300 188.400 ;
        RECT 607.950 186.450 610.050 187.200 ;
        RECT 553.950 181.050 555.750 182.850 ;
        RECT 566.100 181.050 567.900 182.850 ;
        RECT 569.700 181.050 570.900 186.300 ;
        RECT 590.700 185.400 594.300 186.300 ;
        RECT 599.550 185.550 610.050 186.450 ;
        RECT 571.950 181.050 573.750 182.850 ;
        RECT 587.100 181.050 588.900 182.850 ;
        RECT 590.700 181.050 591.900 185.400 ;
        RECT 593.100 181.050 594.900 182.850 ;
        RECT 460.500 178.950 462.600 181.050 ;
        RECT 463.800 178.950 465.900 181.050 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 478.950 178.950 481.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 505.950 178.950 508.050 181.050 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 529.950 178.950 532.050 181.050 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 460.200 177.150 462.000 178.950 ;
        RECT 464.400 171.600 465.300 178.950 ;
        RECT 437.100 159.000 438.900 165.600 ;
        RECT 440.100 159.600 441.900 165.600 ;
        RECT 443.100 159.000 444.900 165.600 ;
        RECT 455.100 159.000 456.900 165.600 ;
        RECT 458.100 159.600 459.900 165.600 ;
        RECT 461.100 159.000 462.900 171.000 ;
        RECT 464.100 159.600 465.900 171.600 ;
        RECT 479.700 165.600 480.900 178.950 ;
        RECT 484.950 171.450 487.050 172.050 ;
        RECT 496.950 171.450 499.050 172.050 ;
        RECT 484.950 170.550 499.050 171.450 ;
        RECT 484.950 169.950 487.050 170.550 ;
        RECT 496.950 169.950 499.050 170.550 ;
        RECT 500.100 171.600 501.300 178.950 ;
        RECT 506.100 177.150 507.900 178.950 ;
        RECT 500.100 170.100 502.500 171.600 ;
        RECT 498.000 167.100 499.800 168.900 ;
        RECT 476.100 159.000 477.900 165.600 ;
        RECT 479.100 159.600 480.900 165.600 ;
        RECT 482.100 159.000 483.900 165.600 ;
        RECT 497.700 159.000 499.500 165.600 ;
        RECT 500.700 159.600 502.500 170.100 ;
        RECT 505.800 159.000 507.600 171.600 ;
        RECT 522.000 166.800 522.900 178.950 ;
        RECT 527.100 177.150 528.900 178.950 ;
        RECT 545.100 177.150 546.900 178.950 ;
        RECT 526.950 174.450 529.050 175.050 ;
        RECT 535.950 174.450 538.050 175.050 ;
        RECT 526.950 173.550 538.050 174.450 ;
        RECT 526.950 172.950 529.050 173.550 ;
        RECT 535.950 172.950 538.050 173.550 ;
        RECT 549.000 173.400 549.900 178.950 ;
        RECT 550.950 177.150 552.750 178.950 ;
        RECT 559.950 178.050 562.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 559.950 177.000 565.050 178.050 ;
        RECT 560.550 176.550 565.050 177.000 ;
        RECT 561.000 175.950 565.050 176.550 ;
        RECT 545.100 172.500 549.900 173.400 ;
        RECT 522.000 165.900 528.600 166.800 ;
        RECT 522.000 165.600 522.900 165.900 ;
        RECT 521.100 159.600 522.900 165.600 ;
        RECT 527.100 165.600 528.600 165.900 ;
        RECT 524.100 159.000 525.900 165.000 ;
        RECT 527.100 159.600 528.900 165.600 ;
        RECT 530.100 159.000 531.900 165.600 ;
        RECT 542.100 160.500 543.900 171.600 ;
        RECT 545.100 161.400 546.900 172.500 ;
        RECT 548.100 170.400 555.900 171.300 ;
        RECT 548.100 160.500 549.900 170.400 ;
        RECT 542.100 159.600 549.900 160.500 ;
        RECT 551.100 159.000 552.900 169.500 ;
        RECT 554.100 159.600 555.900 170.400 ;
        RECT 569.700 165.600 570.900 178.950 ;
        RECT 584.100 177.150 585.900 178.950 ;
        RECT 574.950 174.450 577.050 175.050 ;
        RECT 586.950 174.450 589.050 175.050 ;
        RECT 574.950 173.550 589.050 174.450 ;
        RECT 574.950 172.950 577.050 173.550 ;
        RECT 586.950 172.950 589.050 173.550 ;
        RECT 590.700 171.600 591.900 178.950 ;
        RECT 599.550 178.050 600.450 185.550 ;
        RECT 607.950 185.100 610.050 185.550 ;
        RECT 605.100 181.050 606.900 182.850 ;
        RECT 611.250 181.050 613.050 182.850 ;
        RECT 614.700 181.050 615.600 188.400 ;
        RECT 626.700 188.400 629.400 190.200 ;
        RECT 630.600 188.400 632.400 195.000 ;
        RECT 626.700 181.050 627.600 188.400 ;
        RECT 628.500 186.600 630.300 187.500 ;
        RECT 635.100 186.600 636.900 194.400 ;
        RECT 628.500 185.700 636.900 186.600 ;
        RECT 647.700 187.200 649.500 194.400 ;
        RECT 652.800 188.400 654.600 195.000 ;
        RECT 667.500 188.400 669.300 195.000 ;
        RECT 672.000 188.400 673.800 194.400 ;
        RECT 676.500 188.400 678.300 195.000 ;
        RECT 689.100 189.300 690.900 194.400 ;
        RECT 692.100 190.200 693.900 195.000 ;
        RECT 695.100 189.300 696.900 194.400 ;
        RECT 647.700 186.300 651.900 187.200 ;
        RECT 604.950 178.950 607.050 181.050 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 626.100 178.950 628.200 181.050 ;
        RECT 629.400 178.950 631.500 181.050 ;
        RECT 599.550 176.550 604.050 178.050 ;
        RECT 608.250 177.150 610.050 178.950 ;
        RECT 600.000 175.950 604.050 176.550 ;
        RECT 614.700 171.600 615.600 178.950 ;
        RECT 626.700 171.600 627.600 178.950 ;
        RECT 630.000 177.150 631.800 178.950 ;
        RECT 566.100 159.000 567.900 165.600 ;
        RECT 569.100 159.600 570.900 165.600 ;
        RECT 572.100 159.000 573.900 165.600 ;
        RECT 584.400 159.000 586.200 171.600 ;
        RECT 589.500 170.100 591.900 171.600 ;
        RECT 605.100 170.700 612.900 171.600 ;
        RECT 589.500 159.600 591.300 170.100 ;
        RECT 592.200 167.100 594.000 168.900 ;
        RECT 592.500 159.000 594.300 165.600 ;
        RECT 605.100 159.600 606.900 170.700 ;
        RECT 608.100 159.000 609.900 169.800 ;
        RECT 611.100 159.600 612.900 170.700 ;
        RECT 614.100 159.600 615.900 171.600 ;
        RECT 626.100 159.600 627.900 171.600 ;
        RECT 629.100 159.000 630.900 171.000 ;
        RECT 633.000 165.600 633.900 185.700 ;
        RECT 643.950 183.450 646.050 184.050 ;
        RECT 634.950 181.050 636.750 182.850 ;
        RECT 638.550 182.550 646.050 183.450 ;
        RECT 634.800 178.950 636.900 181.050 ;
        RECT 638.550 175.050 639.450 182.550 ;
        RECT 643.950 181.950 646.050 182.550 ;
        RECT 647.100 181.050 648.900 182.850 ;
        RECT 650.700 181.050 651.900 186.300 ;
        RECT 652.950 181.050 654.750 182.850 ;
        RECT 665.100 181.050 666.900 182.850 ;
        RECT 671.700 181.050 672.900 188.400 ;
        RECT 689.100 187.950 696.900 189.300 ;
        RECT 698.100 188.400 699.900 194.400 ;
        RECT 710.100 191.400 711.900 194.400 ;
        RECT 713.100 191.400 714.900 195.000 ;
        RECT 698.100 186.300 699.300 188.400 ;
        RECT 695.700 185.400 699.300 186.300 ;
        RECT 676.950 181.050 678.750 182.850 ;
        RECT 692.100 181.050 693.900 182.850 ;
        RECT 695.700 181.050 696.900 185.400 ;
        RECT 700.950 183.450 705.000 184.050 ;
        RECT 698.100 181.050 699.900 182.850 ;
        RECT 700.950 181.950 705.450 183.450 ;
        RECT 646.950 178.950 649.050 181.050 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 667.950 178.950 670.050 181.050 ;
        RECT 670.950 178.950 673.050 181.050 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 691.950 178.950 694.050 181.050 ;
        RECT 694.950 178.950 697.050 181.050 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 634.950 173.550 639.450 175.050 ;
        RECT 634.950 172.950 639.000 173.550 ;
        RECT 650.700 165.600 651.900 178.950 ;
        RECT 668.100 177.150 669.900 178.950 ;
        RECT 672.000 173.400 672.900 178.950 ;
        RECT 673.950 177.150 675.750 178.950 ;
        RECT 689.100 177.150 690.900 178.950 ;
        RECT 668.100 172.500 672.900 173.400 ;
        RECT 632.100 159.600 633.900 165.600 ;
        RECT 635.100 159.000 636.900 165.600 ;
        RECT 647.100 159.000 648.900 165.600 ;
        RECT 650.100 159.600 651.900 165.600 ;
        RECT 653.100 159.000 654.900 165.600 ;
        RECT 665.100 160.500 666.900 171.600 ;
        RECT 668.100 161.400 669.900 172.500 ;
        RECT 695.700 171.600 696.900 178.950 ;
        RECT 704.550 178.050 705.450 181.950 ;
        RECT 710.700 181.050 711.900 191.400 ;
        RECT 725.400 188.400 727.200 195.000 ;
        RECT 730.500 187.200 732.300 194.400 ;
        RECT 746.100 191.400 747.900 195.000 ;
        RECT 749.100 191.400 750.900 194.400 ;
        RECT 752.100 191.400 753.900 195.000 ;
        RECT 712.950 186.450 715.050 187.200 ;
        RECT 718.950 186.450 721.050 187.050 ;
        RECT 712.950 185.550 721.050 186.450 ;
        RECT 712.950 185.100 715.050 185.550 ;
        RECT 718.950 184.950 721.050 185.550 ;
        RECT 728.100 186.300 732.300 187.200 ;
        RECT 725.250 181.050 727.050 182.850 ;
        RECT 728.100 181.050 729.300 186.300 ;
        RECT 733.950 183.450 738.000 184.050 ;
        RECT 731.100 181.050 732.900 182.850 ;
        RECT 733.950 181.950 738.450 183.450 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 712.950 178.950 715.050 181.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 700.950 176.550 705.450 178.050 ;
        RECT 700.950 175.950 705.000 176.550 ;
        RECT 671.100 170.400 678.900 171.300 ;
        RECT 671.100 160.500 672.900 170.400 ;
        RECT 665.100 159.600 672.900 160.500 ;
        RECT 674.100 159.000 675.900 169.500 ;
        RECT 677.100 159.600 678.900 170.400 ;
        RECT 689.400 159.000 691.200 171.600 ;
        RECT 694.500 170.100 696.900 171.600 ;
        RECT 694.500 159.600 696.300 170.100 ;
        RECT 697.200 167.100 699.000 168.900 ;
        RECT 710.700 165.600 711.900 178.950 ;
        RECT 713.100 177.150 714.900 178.950 ;
        RECT 728.100 165.600 729.300 178.950 ;
        RECT 737.550 177.450 738.450 181.950 ;
        RECT 749.400 181.050 750.300 191.400 ;
        RECT 764.100 189.300 765.900 194.400 ;
        RECT 767.100 190.200 768.900 195.000 ;
        RECT 770.100 189.300 771.900 194.400 ;
        RECT 764.100 187.950 771.900 189.300 ;
        RECT 773.100 188.400 774.900 194.400 ;
        RECT 785.100 191.400 786.900 195.000 ;
        RECT 788.100 191.400 789.900 194.400 ;
        RECT 791.100 191.400 792.900 195.000 ;
        RECT 757.950 184.950 760.050 187.050 ;
        RECT 773.100 186.300 774.300 188.400 ;
        RECT 770.700 185.400 774.300 186.300 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 748.950 178.950 751.050 181.050 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 742.950 177.450 745.050 178.050 ;
        RECT 737.550 176.550 745.050 177.450 ;
        RECT 746.250 177.150 748.050 178.950 ;
        RECT 742.950 175.950 745.050 176.550 ;
        RECT 749.400 171.600 750.300 178.950 ;
        RECT 752.100 177.150 753.900 178.950 ;
        RECT 758.550 178.050 759.450 184.950 ;
        RECT 767.100 181.050 768.900 182.850 ;
        RECT 770.700 181.050 771.900 185.400 ;
        RECT 773.100 181.050 774.900 182.850 ;
        RECT 788.700 181.050 789.600 191.400 ;
        RECT 803.100 188.400 804.900 194.400 ;
        RECT 803.700 186.300 804.900 188.400 ;
        RECT 806.100 189.300 807.900 194.400 ;
        RECT 809.100 190.200 810.900 195.000 ;
        RECT 812.100 189.300 813.900 194.400 ;
        RECT 806.100 187.950 813.900 189.300 ;
        RECT 827.100 188.400 828.900 194.400 ;
        RECT 830.100 189.300 831.900 195.000 ;
        RECT 834.600 188.400 836.400 194.400 ;
        RECT 839.100 189.300 840.900 195.000 ;
        RECT 842.100 188.400 843.900 194.400 ;
        RECT 854.100 188.400 855.900 194.400 ;
        RECT 857.400 189.300 859.200 195.000 ;
        RECT 861.900 189.000 863.700 194.400 ;
        RECT 866.100 189.300 867.900 195.000 ;
        RECT 827.100 187.500 831.900 188.400 ;
        RECT 829.800 186.300 831.900 187.500 ;
        RECT 834.900 186.900 836.100 188.400 ;
        RECT 803.700 185.400 807.300 186.300 ;
        RECT 803.100 181.050 804.900 182.850 ;
        RECT 806.100 181.050 807.300 185.400 ;
        RECT 833.100 184.800 836.100 186.900 ;
        RECT 842.100 186.600 843.300 188.400 ;
        RECT 854.100 187.500 858.600 188.400 ;
        RECT 814.950 183.450 817.050 184.050 ;
        RECT 814.950 183.000 825.450 183.450 ;
        RECT 809.100 181.050 810.900 182.850 ;
        RECT 814.950 182.550 826.050 183.000 ;
        RECT 814.950 181.950 817.050 182.550 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 769.950 178.950 772.050 181.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 823.950 178.950 826.050 182.550 ;
        RECT 831.900 181.800 834.000 183.900 ;
        RECT 827.100 178.950 829.200 181.050 ;
        RECT 831.900 180.000 833.700 181.800 ;
        RECT 834.900 179.100 836.100 184.800 ;
        RECT 837.000 185.700 843.300 186.600 ;
        RECT 837.000 183.600 839.100 185.700 ;
        RECT 856.500 185.100 858.600 187.500 ;
        RECT 861.900 186.900 862.800 189.000 ;
        RECT 869.100 188.400 870.900 194.400 ;
        RECT 869.400 187.500 870.900 188.400 ;
        RECT 859.800 184.800 862.800 186.900 ;
        RECT 866.400 186.000 870.900 187.500 ;
        RECT 837.000 181.800 838.800 183.600 ;
        RECT 841.800 181.050 843.600 182.850 ;
        RECT 841.800 180.300 843.900 181.050 ;
        RECT 758.550 176.550 763.050 178.050 ;
        RECT 764.100 177.150 765.900 178.950 ;
        RECT 759.000 175.950 763.050 176.550 ;
        RECT 770.700 171.600 771.900 178.950 ;
        RECT 785.100 177.150 786.900 178.950 ;
        RECT 788.700 171.600 789.600 178.950 ;
        RECT 790.950 177.150 792.750 178.950 ;
        RECT 806.100 171.600 807.300 178.950 ;
        RECT 812.100 177.150 813.900 178.950 ;
        RECT 827.400 177.150 829.200 178.950 ;
        RECT 833.700 178.200 836.100 179.100 ;
        RECT 837.000 178.950 843.900 180.300 ;
        RECT 854.100 178.950 856.200 181.050 ;
        RECT 858.900 180.900 861.000 183.000 ;
        RECT 859.200 179.100 861.000 180.900 ;
        RECT 837.000 178.500 838.800 178.950 ;
        RECT 833.700 178.050 835.200 178.200 ;
        RECT 833.100 175.950 835.200 178.050 ;
        RECT 834.300 174.000 835.200 175.950 ;
        RECT 836.100 175.500 840.000 177.300 ;
        RECT 854.400 177.150 856.200 178.950 ;
        RECT 861.900 178.050 862.800 184.800 ;
        RECT 863.700 183.900 865.500 185.700 ;
        RECT 866.400 185.400 868.500 186.000 ;
        RECT 864.000 183.000 866.100 183.900 ;
        RECT 864.000 181.800 870.600 183.000 ;
        RECT 868.800 181.200 870.600 181.800 ;
        RECT 864.000 178.800 866.100 180.900 ;
        RECT 868.800 178.950 870.900 181.200 ;
        RECT 859.800 176.700 862.800 178.050 ;
        RECT 864.300 177.000 866.100 178.800 ;
        RECT 859.800 175.950 861.900 176.700 ;
        RECT 836.100 175.200 838.200 175.500 ;
        RECT 834.300 172.950 835.800 174.000 ;
        RECT 829.800 171.600 831.900 172.500 ;
        RECT 697.500 159.000 699.300 165.600 ;
        RECT 710.100 159.600 711.900 165.600 ;
        RECT 713.100 159.000 714.900 165.600 ;
        RECT 725.100 159.000 726.900 165.600 ;
        RECT 728.100 159.600 729.900 165.600 ;
        RECT 731.100 159.000 732.900 165.600 ;
        RECT 746.100 159.000 747.900 171.600 ;
        RECT 749.400 170.400 753.000 171.600 ;
        RECT 751.200 159.600 753.000 170.400 ;
        RECT 764.400 159.000 766.200 171.600 ;
        RECT 769.500 170.100 771.900 171.600 ;
        RECT 786.000 170.400 789.600 171.600 ;
        RECT 769.500 159.600 771.300 170.100 ;
        RECT 772.200 167.100 774.000 168.900 ;
        RECT 772.500 159.000 774.300 165.600 ;
        RECT 786.000 159.600 787.800 170.400 ;
        RECT 791.100 159.000 792.900 171.600 ;
        RECT 806.100 170.100 808.500 171.600 ;
        RECT 804.000 167.100 805.800 168.900 ;
        RECT 803.700 159.000 805.500 165.600 ;
        RECT 806.700 159.600 808.500 170.100 ;
        RECT 811.800 159.000 813.600 171.600 ;
        RECT 827.100 170.400 831.900 171.600 ;
        RECT 834.600 171.600 835.800 172.950 ;
        RECT 839.400 171.600 841.500 173.700 ;
        RECT 857.100 171.600 859.200 172.500 ;
        RECT 827.100 159.600 828.900 170.400 ;
        RECT 830.100 159.000 831.900 169.500 ;
        RECT 834.600 159.600 836.400 171.600 ;
        RECT 839.400 170.700 843.900 171.600 ;
        RECT 839.100 159.000 840.900 169.500 ;
        RECT 842.100 159.600 843.900 170.700 ;
        RECT 854.100 170.400 859.200 171.600 ;
        RECT 860.100 171.600 861.300 175.950 ;
        RECT 862.800 173.700 864.600 175.500 ;
        RECT 862.800 172.800 868.200 173.700 ;
        RECT 866.100 171.900 868.200 172.800 ;
        RECT 860.100 170.700 863.400 171.600 ;
        RECT 866.100 170.700 870.900 171.900 ;
        RECT 854.100 159.600 855.900 170.400 ;
        RECT 857.100 159.000 859.200 169.500 ;
        RECT 861.600 159.600 863.400 170.700 ;
        RECT 866.100 159.000 867.900 169.500 ;
        RECT 869.100 159.600 870.900 170.700 ;
        RECT 11.100 143.400 12.900 155.400 ;
        RECT 14.100 144.300 15.900 155.400 ;
        RECT 17.100 145.200 18.900 156.000 ;
        RECT 20.100 144.300 21.900 155.400 ;
        RECT 32.100 149.400 33.900 156.000 ;
        RECT 35.100 149.400 36.900 155.400 ;
        RECT 38.100 150.000 39.900 156.000 ;
        RECT 35.400 149.100 36.900 149.400 ;
        RECT 41.100 149.400 42.900 155.400 ;
        RECT 41.100 149.100 42.000 149.400 ;
        RECT 35.400 148.200 42.000 149.100 ;
        RECT 14.100 143.400 21.900 144.300 ;
        RECT 11.400 136.050 12.300 143.400 ;
        RECT 13.950 141.450 16.050 142.050 ;
        RECT 31.950 141.450 34.050 142.050 ;
        RECT 13.950 140.550 34.050 141.450 ;
        RECT 13.950 139.950 16.050 140.550 ;
        RECT 31.950 139.950 34.050 140.550 ;
        RECT 16.950 136.050 18.750 137.850 ;
        RECT 35.100 136.050 36.900 137.850 ;
        RECT 41.100 136.050 42.000 148.200 ;
        RECT 53.400 143.400 55.200 156.000 ;
        RECT 58.500 144.900 60.300 155.400 ;
        RECT 61.500 149.400 63.300 156.000 ;
        RECT 74.100 149.400 75.900 155.400 ;
        RECT 77.100 150.000 78.900 156.000 ;
        RECT 75.000 149.100 75.900 149.400 ;
        RECT 80.100 149.400 81.900 155.400 ;
        RECT 83.100 149.400 84.900 156.000 ;
        RECT 80.100 149.100 81.600 149.400 ;
        RECT 75.000 148.200 81.600 149.100 ;
        RECT 61.200 146.100 63.000 147.900 ;
        RECT 58.500 143.400 60.900 144.900 ;
        RECT 48.000 138.450 52.050 139.050 ;
        RECT 47.550 136.950 52.050 138.450 ;
        RECT 10.950 133.950 13.050 136.050 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 11.400 126.600 12.300 133.950 ;
        RECT 13.950 132.150 15.750 133.950 ;
        RECT 20.100 132.150 21.900 133.950 ;
        RECT 25.950 133.050 28.050 136.050 ;
        RECT 31.950 133.950 34.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 25.950 132.000 31.050 133.050 ;
        RECT 32.100 132.150 33.900 133.950 ;
        RECT 38.100 132.150 39.900 133.950 ;
        RECT 26.550 131.550 31.050 132.000 ;
        RECT 27.000 130.950 31.050 131.550 ;
        RECT 41.100 130.200 42.000 133.950 ;
        RECT 47.550 133.050 48.450 136.950 ;
        RECT 53.100 136.050 54.900 137.850 ;
        RECT 59.700 136.050 60.900 143.400 ;
        RECT 75.000 136.050 75.900 148.200 ;
        RECT 82.950 144.450 85.050 145.050 ;
        RECT 88.950 144.450 91.050 145.050 ;
        RECT 82.950 143.550 91.050 144.450 ;
        RECT 82.950 142.950 85.050 143.550 ;
        RECT 88.950 142.950 91.050 143.550 ;
        RECT 95.100 143.400 96.900 155.400 ;
        RECT 98.100 144.300 99.900 155.400 ;
        RECT 101.100 145.200 102.900 156.000 ;
        RECT 104.100 144.300 105.900 155.400 ;
        RECT 98.100 143.400 105.900 144.300 ;
        RECT 116.400 143.400 118.200 156.000 ;
        RECT 121.500 144.900 123.300 155.400 ;
        RECT 124.500 149.400 126.300 156.000 ;
        RECT 137.100 149.400 138.900 155.400 ;
        RECT 140.100 150.000 141.900 156.000 ;
        RECT 138.000 149.100 138.900 149.400 ;
        RECT 143.100 149.400 144.900 155.400 ;
        RECT 146.100 149.400 147.900 156.000 ;
        RECT 161.100 149.400 162.900 155.400 ;
        RECT 164.100 150.000 165.900 156.000 ;
        RECT 143.100 149.100 144.600 149.400 ;
        RECT 138.000 148.200 144.600 149.100 ;
        RECT 162.000 149.100 162.900 149.400 ;
        RECT 167.100 149.400 168.900 155.400 ;
        RECT 170.100 149.400 171.900 156.000 ;
        RECT 182.100 149.400 183.900 156.000 ;
        RECT 185.100 149.400 186.900 155.400 ;
        RECT 188.100 149.400 189.900 156.000 ;
        RECT 203.100 149.400 204.900 156.000 ;
        RECT 206.100 149.400 207.900 155.400 ;
        RECT 209.100 149.400 210.900 156.000 ;
        RECT 221.100 149.400 222.900 155.400 ;
        RECT 224.100 150.000 225.900 156.000 ;
        RECT 167.100 149.100 168.600 149.400 ;
        RECT 162.000 148.200 168.600 149.100 ;
        RECT 124.200 146.100 126.000 147.900 ;
        RECT 121.500 143.400 123.900 144.900 ;
        RECT 80.100 136.050 81.900 137.850 ;
        RECT 95.400 136.050 96.300 143.400 ;
        RECT 100.950 136.050 102.750 137.850 ;
        RECT 116.100 136.050 117.900 137.850 ;
        RECT 122.700 136.050 123.900 143.400 ;
        RECT 138.000 136.050 138.900 148.200 ;
        RECT 145.950 147.450 148.050 148.050 ;
        RECT 154.950 147.450 157.050 148.050 ;
        RECT 145.950 146.550 157.050 147.450 ;
        RECT 145.950 145.950 148.050 146.550 ;
        RECT 154.950 145.950 157.050 146.550 ;
        RECT 143.100 136.050 144.900 137.850 ;
        RECT 162.000 136.050 162.900 148.200 ;
        RECT 175.950 147.450 178.050 148.050 ;
        RECT 181.950 147.450 184.050 148.050 ;
        RECT 175.950 146.550 184.050 147.450 ;
        RECT 175.950 145.950 178.050 146.550 ;
        RECT 181.950 145.950 184.050 146.550 ;
        RECT 163.950 141.450 166.050 142.200 ;
        RECT 175.950 141.450 178.050 142.050 ;
        RECT 163.950 140.550 178.050 141.450 ;
        RECT 163.950 140.100 166.050 140.550 ;
        RECT 175.950 139.950 178.050 140.550 ;
        RECT 167.100 136.050 168.900 137.850 ;
        RECT 185.100 136.050 186.300 149.400 ;
        RECT 206.100 136.050 207.300 149.400 ;
        RECT 222.000 149.100 222.900 149.400 ;
        RECT 227.100 149.400 228.900 155.400 ;
        RECT 230.100 149.400 231.900 156.000 ;
        RECT 242.100 149.400 243.900 156.000 ;
        RECT 245.100 149.400 246.900 155.400 ;
        RECT 227.100 149.100 228.600 149.400 ;
        RECT 222.000 148.200 228.600 149.100 ;
        RECT 222.000 136.050 222.900 148.200 ;
        RECT 229.950 141.450 232.050 142.050 ;
        RECT 241.950 141.450 244.050 141.900 ;
        RECT 229.950 140.550 244.050 141.450 ;
        RECT 229.950 139.950 232.050 140.550 ;
        RECT 241.950 139.800 244.050 140.550 ;
        RECT 227.100 136.050 228.900 137.850 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 94.950 133.950 97.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 115.950 133.950 118.050 136.050 ;
        RECT 118.950 133.950 121.050 136.050 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 136.950 133.950 139.050 136.050 ;
        RECT 139.950 133.950 142.050 136.050 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 160.950 133.950 163.050 136.050 ;
        RECT 163.950 133.950 166.050 136.050 ;
        RECT 166.950 133.950 169.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 184.950 133.950 187.050 136.050 ;
        RECT 187.950 133.950 190.050 136.050 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 205.950 133.950 208.050 136.050 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 242.100 133.950 244.200 136.050 ;
        RECT 43.950 131.550 48.450 133.050 ;
        RECT 56.100 132.150 57.900 133.950 ;
        RECT 43.950 130.950 48.000 131.550 ;
        RECT 16.950 129.450 19.050 130.050 ;
        RECT 25.950 129.450 28.050 130.050 ;
        RECT 16.950 128.550 28.050 129.450 ;
        RECT 16.950 127.950 19.050 128.550 ;
        RECT 25.950 127.950 28.050 128.550 ;
        RECT 11.400 125.400 16.500 126.600 ;
        RECT 11.700 120.000 13.500 123.600 ;
        RECT 14.700 120.600 16.500 125.400 ;
        RECT 19.200 120.000 21.000 126.600 ;
        RECT 32.100 120.000 33.900 129.600 ;
        RECT 38.700 129.000 42.000 130.200 ;
        RECT 59.700 129.600 60.900 133.950 ;
        RECT 62.100 132.150 63.900 133.950 ;
        RECT 75.000 130.200 75.900 133.950 ;
        RECT 77.100 132.150 78.900 133.950 ;
        RECT 83.100 132.150 84.900 133.950 ;
        RECT 38.700 120.600 40.500 129.000 ;
        RECT 59.700 128.700 63.300 129.600 ;
        RECT 75.000 129.000 78.300 130.200 ;
        RECT 53.100 125.700 60.900 127.050 ;
        RECT 53.100 120.600 54.900 125.700 ;
        RECT 56.100 120.000 57.900 124.800 ;
        RECT 59.100 120.600 60.900 125.700 ;
        RECT 62.100 126.600 63.300 128.700 ;
        RECT 62.100 120.600 63.900 126.600 ;
        RECT 76.500 120.600 78.300 129.000 ;
        RECT 83.100 120.000 84.900 129.600 ;
        RECT 95.400 126.600 96.300 133.950 ;
        RECT 97.950 132.150 99.750 133.950 ;
        RECT 104.100 132.150 105.900 133.950 ;
        RECT 119.100 132.150 120.900 133.950 ;
        RECT 122.700 129.600 123.900 133.950 ;
        RECT 125.100 132.150 126.900 133.950 ;
        RECT 138.000 130.200 138.900 133.950 ;
        RECT 140.100 132.150 141.900 133.950 ;
        RECT 146.100 132.150 147.900 133.950 ;
        RECT 162.000 130.200 162.900 133.950 ;
        RECT 164.100 132.150 165.900 133.950 ;
        RECT 170.100 132.150 171.900 133.950 ;
        RECT 182.250 132.150 184.050 133.950 ;
        RECT 122.700 128.700 126.300 129.600 ;
        RECT 138.000 129.000 141.300 130.200 ;
        RECT 95.400 125.400 100.500 126.600 ;
        RECT 95.700 120.000 97.500 123.600 ;
        RECT 98.700 120.600 100.500 125.400 ;
        RECT 103.200 120.000 105.000 126.600 ;
        RECT 116.100 125.700 123.900 127.050 ;
        RECT 116.100 120.600 117.900 125.700 ;
        RECT 119.100 120.000 120.900 124.800 ;
        RECT 122.100 120.600 123.900 125.700 ;
        RECT 125.100 126.600 126.300 128.700 ;
        RECT 125.100 120.600 126.900 126.600 ;
        RECT 139.500 120.600 141.300 129.000 ;
        RECT 146.100 120.000 147.900 129.600 ;
        RECT 162.000 129.000 165.300 130.200 ;
        RECT 163.500 120.600 165.300 129.000 ;
        RECT 170.100 120.000 171.900 129.600 ;
        RECT 185.100 128.700 186.300 133.950 ;
        RECT 188.100 132.150 189.900 133.950 ;
        RECT 203.250 132.150 205.050 133.950 ;
        RECT 206.100 128.700 207.300 133.950 ;
        RECT 209.100 132.150 210.900 133.950 ;
        RECT 222.000 130.200 222.900 133.950 ;
        RECT 224.100 132.150 225.900 133.950 ;
        RECT 230.100 132.150 231.900 133.950 ;
        RECT 242.250 132.150 244.050 133.950 ;
        RECT 222.000 129.000 225.300 130.200 ;
        RECT 185.100 127.800 189.300 128.700 ;
        RECT 206.100 127.800 210.300 128.700 ;
        RECT 182.400 120.000 184.200 126.600 ;
        RECT 187.500 120.600 189.300 127.800 ;
        RECT 203.400 120.000 205.200 126.600 ;
        RECT 208.500 120.600 210.300 127.800 ;
        RECT 223.500 120.600 225.300 129.000 ;
        RECT 230.100 120.000 231.900 129.600 ;
        RECT 245.100 129.300 246.000 149.400 ;
        RECT 248.100 144.000 249.900 156.000 ;
        RECT 251.100 143.400 252.900 155.400 ;
        RECT 263.100 149.400 264.900 155.400 ;
        RECT 266.100 149.400 267.900 156.000 ;
        RECT 278.100 149.400 279.900 156.000 ;
        RECT 281.100 149.400 282.900 155.400 ;
        RECT 284.100 149.400 285.900 156.000 ;
        RECT 247.200 136.050 249.000 137.850 ;
        RECT 251.400 136.050 252.300 143.400 ;
        RECT 263.700 136.050 264.900 149.400 ;
        RECT 266.100 136.050 267.900 137.850 ;
        RECT 281.100 136.050 282.300 149.400 ;
        RECT 296.100 144.300 297.900 155.400 ;
        RECT 299.100 145.200 300.900 156.000 ;
        RECT 302.100 144.300 303.900 155.400 ;
        RECT 296.100 143.400 303.900 144.300 ;
        RECT 305.100 143.400 306.900 155.400 ;
        RECT 318.000 144.600 319.800 155.400 ;
        RECT 318.000 143.400 321.600 144.600 ;
        RECT 323.100 143.400 324.900 156.000 ;
        RECT 335.100 149.400 336.900 156.000 ;
        RECT 338.100 149.400 339.900 155.400 ;
        RECT 341.100 149.400 342.900 156.000 ;
        RECT 353.100 149.400 354.900 156.000 ;
        RECT 356.100 149.400 357.900 155.400 ;
        RECT 359.100 149.400 360.900 156.000 ;
        RECT 371.700 149.400 373.500 156.000 ;
        RECT 299.250 136.050 301.050 137.850 ;
        RECT 305.700 136.050 306.600 143.400 ;
        RECT 317.100 136.050 318.900 137.850 ;
        RECT 320.700 136.050 321.600 143.400 ;
        RECT 322.950 136.050 324.750 137.850 ;
        RECT 338.700 136.050 339.900 149.400 ;
        RECT 343.950 138.450 348.000 139.050 ;
        RECT 343.950 136.950 348.450 138.450 ;
        RECT 247.500 133.950 249.600 136.050 ;
        RECT 250.800 133.950 252.900 136.050 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 304.950 133.950 307.050 136.050 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 242.100 128.400 250.500 129.300 ;
        RECT 242.100 120.600 243.900 128.400 ;
        RECT 248.700 127.500 250.500 128.400 ;
        RECT 251.400 126.600 252.300 133.950 ;
        RECT 246.600 120.000 248.400 126.600 ;
        RECT 249.600 124.800 252.300 126.600 ;
        RECT 249.600 120.600 251.400 124.800 ;
        RECT 263.700 123.600 264.900 133.950 ;
        RECT 278.250 132.150 280.050 133.950 ;
        RECT 281.100 128.700 282.300 133.950 ;
        RECT 284.100 132.150 285.900 133.950 ;
        RECT 296.100 132.150 297.900 133.950 ;
        RECT 302.250 132.150 304.050 133.950 ;
        RECT 281.100 127.800 285.300 128.700 ;
        RECT 263.100 120.600 264.900 123.600 ;
        RECT 266.100 120.000 267.900 123.600 ;
        RECT 278.400 120.000 280.200 126.600 ;
        RECT 283.500 120.600 285.300 127.800 ;
        RECT 305.700 126.600 306.600 133.950 ;
        RECT 297.000 120.000 298.800 126.600 ;
        RECT 301.500 125.400 306.600 126.600 ;
        RECT 301.500 120.600 303.300 125.400 ;
        RECT 320.700 123.600 321.600 133.950 ;
        RECT 335.100 132.150 336.900 133.950 ;
        RECT 338.700 128.700 339.900 133.950 ;
        RECT 340.950 132.150 342.750 133.950 ;
        RECT 335.700 127.800 339.900 128.700 ;
        RECT 340.950 129.450 343.050 130.050 ;
        RECT 347.550 129.450 348.450 136.950 ;
        RECT 356.700 136.050 357.900 149.400 ;
        RECT 358.950 144.450 361.050 148.050 ;
        RECT 372.000 146.100 373.800 147.900 ;
        RECT 370.950 144.450 373.050 145.050 ;
        RECT 374.700 144.900 376.500 155.400 ;
        RECT 358.950 144.000 373.050 144.450 ;
        RECT 359.550 143.550 373.050 144.000 ;
        RECT 370.950 142.950 373.050 143.550 ;
        RECT 374.100 143.400 376.500 144.900 ;
        RECT 379.800 143.400 381.600 156.000 ;
        RECT 392.100 143.400 393.900 155.400 ;
        RECT 395.100 145.200 396.900 156.000 ;
        RECT 398.100 149.400 399.900 155.400 ;
        RECT 410.100 149.400 411.900 155.400 ;
        RECT 413.100 149.400 414.900 156.000 ;
        RECT 361.950 138.450 366.000 139.050 ;
        RECT 361.950 136.950 366.450 138.450 ;
        RECT 352.950 133.950 355.050 136.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 353.100 132.150 354.900 133.950 ;
        RECT 340.950 128.550 348.450 129.450 ;
        RECT 356.700 128.700 357.900 133.950 ;
        RECT 358.950 132.150 360.750 133.950 ;
        RECT 365.550 132.900 366.450 136.950 ;
        RECT 374.100 136.050 375.300 143.400 ;
        RECT 380.100 136.050 381.900 137.850 ;
        RECT 392.100 136.050 393.300 143.400 ;
        RECT 398.700 142.500 399.900 149.400 ;
        RECT 394.200 141.600 399.900 142.500 ;
        RECT 394.200 140.700 396.000 141.600 ;
        RECT 370.950 133.950 373.050 136.050 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 392.100 133.950 394.200 136.050 ;
        RECT 364.950 130.800 367.050 132.900 ;
        RECT 371.100 132.150 372.900 133.950 ;
        RECT 374.100 129.600 375.300 133.950 ;
        RECT 377.100 132.150 378.900 133.950 ;
        RECT 340.950 127.950 343.050 128.550 ;
        RECT 353.700 127.800 357.900 128.700 ;
        RECT 371.700 128.700 375.300 129.600 ;
        RECT 304.500 120.000 306.300 123.600 ;
        RECT 317.100 120.000 318.900 123.600 ;
        RECT 320.100 120.600 321.900 123.600 ;
        RECT 323.100 120.000 324.900 123.600 ;
        RECT 335.700 120.600 337.500 127.800 ;
        RECT 340.800 120.000 342.600 126.600 ;
        RECT 353.700 120.600 355.500 127.800 ;
        RECT 371.700 126.600 372.900 128.700 ;
        RECT 358.800 120.000 360.600 126.600 ;
        RECT 371.100 120.600 372.900 126.600 ;
        RECT 374.100 125.700 381.900 127.050 ;
        RECT 374.100 120.600 375.900 125.700 ;
        RECT 377.100 120.000 378.900 124.800 ;
        RECT 380.100 120.600 381.900 125.700 ;
        RECT 392.100 126.600 393.300 133.950 ;
        RECT 395.100 129.300 396.000 140.700 ;
        RECT 397.800 136.050 399.600 137.850 ;
        RECT 410.700 136.050 411.900 149.400 ;
        RECT 425.100 143.400 426.900 155.400 ;
        RECT 428.100 144.000 429.900 156.000 ;
        RECT 431.100 149.400 432.900 155.400 ;
        RECT 434.100 149.400 435.900 156.000 ;
        RECT 446.700 149.400 448.500 156.000 ;
        RECT 413.100 136.050 414.900 137.850 ;
        RECT 425.700 136.050 426.600 143.400 ;
        RECT 429.000 136.050 430.800 137.850 ;
        RECT 397.500 133.950 399.600 136.050 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 425.100 133.950 427.200 136.050 ;
        RECT 428.400 133.950 430.500 136.050 ;
        RECT 394.200 128.400 396.000 129.300 ;
        RECT 394.200 127.500 399.900 128.400 ;
        RECT 392.100 120.600 393.900 126.600 ;
        RECT 395.100 120.000 396.900 126.600 ;
        RECT 398.700 123.600 399.900 127.500 ;
        RECT 410.700 123.600 411.900 133.950 ;
        RECT 425.700 126.600 426.600 133.950 ;
        RECT 432.000 129.300 432.900 149.400 ;
        RECT 447.000 146.100 448.800 147.900 ;
        RECT 449.700 144.900 451.500 155.400 ;
        RECT 449.100 143.400 451.500 144.900 ;
        RECT 454.800 143.400 456.600 156.000 ;
        RECT 467.700 149.400 469.500 156.000 ;
        RECT 468.000 146.100 469.800 147.900 ;
        RECT 470.700 144.900 472.500 155.400 ;
        RECT 470.100 143.400 472.500 144.900 ;
        RECT 475.800 143.400 477.600 156.000 ;
        RECT 488.100 144.600 489.900 155.400 ;
        RECT 491.100 145.500 492.900 156.000 ;
        RECT 494.100 154.500 501.900 155.400 ;
        RECT 494.100 144.600 495.900 154.500 ;
        RECT 488.100 143.700 495.900 144.600 ;
        RECT 449.100 136.050 450.300 143.400 ;
        RECT 462.000 138.450 466.050 139.050 ;
        RECT 455.100 136.050 456.900 137.850 ;
        RECT 461.550 136.950 466.050 138.450 ;
        RECT 433.800 133.950 435.900 136.050 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 433.950 132.150 435.750 133.950 ;
        RECT 446.100 132.150 447.900 133.950 ;
        RECT 449.100 129.600 450.300 133.950 ;
        RECT 452.100 132.150 453.900 133.950 ;
        RECT 461.550 133.050 462.450 136.950 ;
        RECT 470.100 136.050 471.300 143.400 ;
        RECT 497.100 142.500 498.900 153.600 ;
        RECT 500.100 143.400 501.900 154.500 ;
        RECT 512.100 143.400 513.900 155.400 ;
        RECT 515.100 144.300 516.900 155.400 ;
        RECT 518.100 145.200 519.900 156.000 ;
        RECT 521.100 144.300 522.900 155.400 ;
        RECT 533.100 149.400 534.900 155.400 ;
        RECT 536.100 150.000 537.900 156.000 ;
        RECT 515.100 143.400 522.900 144.300 ;
        RECT 534.000 149.100 534.900 149.400 ;
        RECT 539.100 149.400 540.900 155.400 ;
        RECT 542.100 149.400 543.900 156.000 ;
        RECT 554.700 149.400 556.500 156.000 ;
        RECT 539.100 149.100 540.600 149.400 ;
        RECT 534.000 148.200 540.600 149.100 ;
        RECT 494.100 141.600 498.900 142.500 ;
        RECT 476.100 136.050 477.900 137.850 ;
        RECT 491.250 136.050 493.050 137.850 ;
        RECT 494.100 136.050 495.000 141.600 ;
        RECT 502.950 138.450 507.000 139.050 ;
        RECT 497.100 136.050 498.900 137.850 ;
        RECT 502.950 136.950 507.450 138.450 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 499.950 133.950 502.050 136.050 ;
        RECT 457.950 131.550 462.450 133.050 ;
        RECT 467.100 132.150 468.900 133.950 ;
        RECT 457.950 130.950 462.000 131.550 ;
        RECT 470.100 129.600 471.300 133.950 ;
        RECT 473.100 132.150 474.900 133.950 ;
        RECT 488.250 132.150 490.050 133.950 ;
        RECT 427.500 128.400 435.900 129.300 ;
        RECT 427.500 127.500 429.300 128.400 ;
        RECT 425.700 124.800 428.400 126.600 ;
        RECT 398.100 120.600 399.900 123.600 ;
        RECT 410.100 120.600 411.900 123.600 ;
        RECT 413.100 120.000 414.900 123.600 ;
        RECT 426.600 120.600 428.400 124.800 ;
        RECT 429.600 120.000 431.400 126.600 ;
        RECT 434.100 120.600 435.900 128.400 ;
        RECT 446.700 128.700 450.300 129.600 ;
        RECT 467.700 128.700 471.300 129.600 ;
        RECT 446.700 126.600 447.900 128.700 ;
        RECT 446.100 120.600 447.900 126.600 ;
        RECT 449.100 125.700 456.900 127.050 ;
        RECT 467.700 126.600 468.900 128.700 ;
        RECT 449.100 120.600 450.900 125.700 ;
        RECT 452.100 120.000 453.900 124.800 ;
        RECT 455.100 120.600 456.900 125.700 ;
        RECT 467.100 120.600 468.900 126.600 ;
        RECT 470.100 125.700 477.900 127.050 ;
        RECT 494.100 126.600 495.300 133.950 ;
        RECT 500.100 132.150 501.900 133.950 ;
        RECT 506.550 133.050 507.450 136.950 ;
        RECT 512.400 136.050 513.300 143.400 ;
        RECT 529.950 138.450 532.050 142.050 ;
        RECT 527.550 138.000 532.050 138.450 ;
        RECT 517.950 136.050 519.750 137.850 ;
        RECT 527.550 137.550 531.450 138.000 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 514.950 133.950 517.050 136.050 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 506.550 131.550 511.050 133.050 ;
        RECT 507.000 130.950 511.050 131.550 ;
        RECT 512.400 126.600 513.300 133.950 ;
        RECT 514.950 132.150 516.750 133.950 ;
        RECT 521.100 132.150 522.900 133.950 ;
        RECT 517.950 129.450 520.050 130.050 ;
        RECT 527.550 129.450 528.450 137.550 ;
        RECT 534.000 136.050 534.900 148.200 ;
        RECT 555.000 146.100 556.800 147.900 ;
        RECT 557.700 144.900 559.500 155.400 ;
        RECT 557.100 143.400 559.500 144.900 ;
        RECT 562.800 143.400 564.600 156.000 ;
        RECT 575.100 149.400 576.900 155.400 ;
        RECT 578.100 150.000 579.900 156.000 ;
        RECT 576.000 149.100 576.900 149.400 ;
        RECT 581.100 149.400 582.900 155.400 ;
        RECT 584.100 149.400 585.900 156.000 ;
        RECT 596.100 149.400 597.900 156.000 ;
        RECT 599.100 149.400 600.900 155.400 ;
        RECT 602.100 149.400 603.900 156.000 ;
        RECT 614.100 149.400 615.900 156.000 ;
        RECT 617.100 149.400 618.900 155.400 ;
        RECT 581.100 149.100 582.600 149.400 ;
        RECT 576.000 148.200 582.600 149.100 ;
        RECT 535.950 141.450 538.050 142.050 ;
        RECT 547.950 141.450 550.050 141.900 ;
        RECT 535.950 140.550 550.050 141.450 ;
        RECT 535.950 139.950 538.050 140.550 ;
        RECT 547.950 139.800 550.050 140.550 ;
        RECT 539.100 136.050 540.900 137.850 ;
        RECT 557.100 136.050 558.300 143.400 ;
        RECT 563.100 136.050 564.900 137.850 ;
        RECT 576.000 136.050 576.900 148.200 ;
        RECT 581.100 136.050 582.900 137.850 ;
        RECT 599.100 136.050 600.300 149.400 ;
        RECT 614.100 136.050 615.900 137.850 ;
        RECT 617.100 136.050 618.300 149.400 ;
        RECT 629.100 143.400 630.900 155.400 ;
        RECT 632.100 144.300 633.900 155.400 ;
        RECT 635.100 145.200 636.900 156.000 ;
        RECT 638.100 144.300 639.900 155.400 ;
        RECT 650.100 149.400 651.900 156.000 ;
        RECT 653.100 149.400 654.900 155.400 ;
        RECT 656.100 150.000 657.900 156.000 ;
        RECT 653.400 149.100 654.900 149.400 ;
        RECT 659.100 149.400 660.900 155.400 ;
        RECT 671.700 149.400 673.500 156.000 ;
        RECT 659.100 149.100 660.000 149.400 ;
        RECT 653.400 148.200 660.000 149.100 ;
        RECT 632.100 143.400 639.900 144.300 ;
        RECT 629.400 136.050 630.300 143.400 ;
        RECT 637.950 141.450 640.050 142.050 ;
        RECT 655.950 141.450 658.050 142.050 ;
        RECT 637.950 140.550 658.050 141.450 ;
        RECT 637.950 139.950 640.050 140.550 ;
        RECT 655.950 139.950 658.050 140.550 ;
        RECT 634.950 136.050 636.750 137.850 ;
        RECT 653.100 136.050 654.900 137.850 ;
        RECT 659.100 136.050 660.000 148.200 ;
        RECT 672.000 146.100 673.800 147.900 ;
        RECT 674.700 144.900 676.500 155.400 ;
        RECT 674.100 143.400 676.500 144.900 ;
        RECT 679.800 143.400 681.600 156.000 ;
        RECT 692.100 149.400 693.900 156.000 ;
        RECT 695.100 149.400 696.900 155.400 ;
        RECT 674.100 136.050 675.300 143.400 ;
        RECT 680.100 136.050 681.900 137.850 ;
        RECT 692.100 136.050 693.900 137.850 ;
        RECT 695.100 136.050 696.300 149.400 ;
        RECT 707.100 144.300 708.900 155.400 ;
        RECT 710.100 145.200 711.900 156.000 ;
        RECT 713.100 144.300 714.900 155.400 ;
        RECT 707.100 143.400 714.900 144.300 ;
        RECT 716.100 143.400 717.900 155.400 ;
        RECT 731.100 149.400 732.900 156.000 ;
        RECT 734.100 149.400 735.900 155.400 ;
        RECT 737.100 149.400 738.900 156.000 ;
        RECT 700.950 139.950 703.050 142.050 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 535.950 133.950 538.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 541.950 133.950 544.050 136.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 556.950 133.950 559.050 136.050 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 577.950 133.950 580.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 631.950 133.950 634.050 136.050 ;
        RECT 634.950 133.950 637.050 136.050 ;
        RECT 637.950 133.950 640.050 136.050 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 655.950 133.950 658.050 136.050 ;
        RECT 658.950 133.950 661.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 701.550 135.900 702.450 139.950 ;
        RECT 710.250 136.050 712.050 137.850 ;
        RECT 716.700 136.050 717.600 143.400 ;
        RECT 734.700 136.050 735.900 149.400 ;
        RECT 749.400 143.400 751.200 156.000 ;
        RECT 754.500 144.900 756.300 155.400 ;
        RECT 757.500 149.400 759.300 156.000 ;
        RECT 757.200 146.100 759.000 147.900 ;
        RECT 754.500 143.400 756.900 144.900 ;
        RECT 770.100 144.300 771.900 155.400 ;
        RECT 773.100 145.200 774.900 156.000 ;
        RECT 776.100 144.300 777.900 155.400 ;
        RECT 770.100 143.400 777.900 144.300 ;
        RECT 779.100 143.400 780.900 155.400 ;
        RECT 791.100 149.400 792.900 156.000 ;
        RECT 794.100 149.400 795.900 155.400 ;
        RECT 797.100 149.400 798.900 156.000 ;
        RECT 749.100 136.050 750.900 137.850 ;
        RECT 755.700 136.050 756.900 143.400 ;
        RECT 760.950 138.450 765.000 139.050 ;
        RECT 760.950 136.950 765.450 138.450 ;
        RECT 517.950 128.550 528.450 129.450 ;
        RECT 534.000 130.200 534.900 133.950 ;
        RECT 536.100 132.150 537.900 133.950 ;
        RECT 542.100 132.150 543.900 133.950 ;
        RECT 554.100 132.150 555.900 133.950 ;
        RECT 534.000 129.000 537.300 130.200 ;
        RECT 557.100 129.600 558.300 133.950 ;
        RECT 560.100 132.150 561.900 133.950 ;
        RECT 517.950 127.950 520.050 128.550 ;
        RECT 470.100 120.600 471.900 125.700 ;
        RECT 473.100 120.000 474.900 124.800 ;
        RECT 476.100 120.600 477.900 125.700 ;
        RECT 488.700 120.000 490.500 126.600 ;
        RECT 493.200 120.600 495.000 126.600 ;
        RECT 497.700 120.000 499.500 126.600 ;
        RECT 512.400 125.400 517.500 126.600 ;
        RECT 512.700 120.000 514.500 123.600 ;
        RECT 515.700 120.600 517.500 125.400 ;
        RECT 520.200 120.000 522.000 126.600 ;
        RECT 535.500 120.600 537.300 129.000 ;
        RECT 542.100 120.000 543.900 129.600 ;
        RECT 554.700 128.700 558.300 129.600 ;
        RECT 576.000 130.200 576.900 133.950 ;
        RECT 578.100 132.150 579.900 133.950 ;
        RECT 584.100 132.150 585.900 133.950 ;
        RECT 596.250 132.150 598.050 133.950 ;
        RECT 576.000 129.000 579.300 130.200 ;
        RECT 554.700 126.600 555.900 128.700 ;
        RECT 554.100 120.600 555.900 126.600 ;
        RECT 557.100 125.700 564.900 127.050 ;
        RECT 557.100 120.600 558.900 125.700 ;
        RECT 560.100 120.000 561.900 124.800 ;
        RECT 563.100 120.600 564.900 125.700 ;
        RECT 577.500 120.600 579.300 129.000 ;
        RECT 584.100 120.000 585.900 129.600 ;
        RECT 599.100 128.700 600.300 133.950 ;
        RECT 602.100 132.150 603.900 133.950 ;
        RECT 599.100 127.800 603.300 128.700 ;
        RECT 596.400 120.000 598.200 126.600 ;
        RECT 601.500 120.600 603.300 127.800 ;
        RECT 617.100 123.600 618.300 133.950 ;
        RECT 629.400 126.600 630.300 133.950 ;
        RECT 631.950 132.150 633.750 133.950 ;
        RECT 638.100 132.150 639.900 133.950 ;
        RECT 650.100 132.150 651.900 133.950 ;
        RECT 656.100 132.150 657.900 133.950 ;
        RECT 659.100 130.200 660.000 133.950 ;
        RECT 671.100 132.150 672.900 133.950 ;
        RECT 629.400 125.400 634.500 126.600 ;
        RECT 614.100 120.000 615.900 123.600 ;
        RECT 617.100 120.600 618.900 123.600 ;
        RECT 629.700 120.000 631.500 123.600 ;
        RECT 632.700 120.600 634.500 125.400 ;
        RECT 637.200 120.000 639.000 126.600 ;
        RECT 650.100 120.000 651.900 129.600 ;
        RECT 656.700 129.000 660.000 130.200 ;
        RECT 674.100 129.600 675.300 133.950 ;
        RECT 677.100 132.150 678.900 133.950 ;
        RECT 656.700 120.600 658.500 129.000 ;
        RECT 671.700 128.700 675.300 129.600 ;
        RECT 671.700 126.600 672.900 128.700 ;
        RECT 671.100 120.600 672.900 126.600 ;
        RECT 674.100 125.700 681.900 127.050 ;
        RECT 674.100 120.600 675.900 125.700 ;
        RECT 677.100 120.000 678.900 124.800 ;
        RECT 680.100 120.600 681.900 125.700 ;
        RECT 695.100 123.600 696.300 133.950 ;
        RECT 700.950 133.800 703.050 135.900 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 709.950 133.950 712.050 136.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 707.100 132.150 708.900 133.950 ;
        RECT 713.250 132.150 715.050 133.950 ;
        RECT 716.700 126.600 717.600 133.950 ;
        RECT 731.100 132.150 732.900 133.950 ;
        RECT 734.700 128.700 735.900 133.950 ;
        RECT 736.950 132.150 738.750 133.950 ;
        RECT 752.100 132.150 753.900 133.950 ;
        RECT 755.700 129.600 756.900 133.950 ;
        RECT 758.100 132.150 759.900 133.950 ;
        RECT 764.550 133.050 765.450 136.950 ;
        RECT 773.250 136.050 775.050 137.850 ;
        RECT 779.700 136.050 780.600 143.400 ;
        RECT 786.000 138.450 790.050 139.050 ;
        RECT 785.550 136.950 790.050 138.450 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 764.550 131.550 769.050 133.050 ;
        RECT 770.100 132.150 771.900 133.950 ;
        RECT 776.250 132.150 778.050 133.950 ;
        RECT 765.000 130.950 769.050 131.550 ;
        RECT 755.700 128.700 759.300 129.600 ;
        RECT 692.100 120.000 693.900 123.600 ;
        RECT 695.100 120.600 696.900 123.600 ;
        RECT 708.000 120.000 709.800 126.600 ;
        RECT 712.500 125.400 717.600 126.600 ;
        RECT 731.700 127.800 735.900 128.700 ;
        RECT 712.500 120.600 714.300 125.400 ;
        RECT 715.500 120.000 717.300 123.600 ;
        RECT 731.700 120.600 733.500 127.800 ;
        RECT 736.800 120.000 738.600 126.600 ;
        RECT 749.100 125.700 756.900 127.050 ;
        RECT 749.100 120.600 750.900 125.700 ;
        RECT 752.100 120.000 753.900 124.800 ;
        RECT 755.100 120.600 756.900 125.700 ;
        RECT 758.100 126.600 759.300 128.700 ;
        RECT 779.700 126.600 780.600 133.950 ;
        RECT 785.550 133.050 786.450 136.950 ;
        RECT 794.700 136.050 795.900 149.400 ;
        RECT 810.000 144.600 811.800 155.400 ;
        RECT 810.000 143.400 813.600 144.600 ;
        RECT 815.100 143.400 816.900 156.000 ;
        RECT 827.100 143.400 828.900 155.400 ;
        RECT 830.100 144.300 831.900 155.400 ;
        RECT 833.100 145.200 834.900 156.000 ;
        RECT 836.100 144.300 837.900 155.400 ;
        RECT 830.100 143.400 837.900 144.300 ;
        RECT 848.400 143.400 850.200 156.000 ;
        RECT 853.500 144.900 855.300 155.400 ;
        RECT 856.500 149.400 858.300 156.000 ;
        RECT 856.200 146.100 858.000 147.900 ;
        RECT 853.500 143.400 855.900 144.900 ;
        RECT 804.000 138.450 808.050 139.050 ;
        RECT 803.550 136.950 808.050 138.450 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 785.550 131.550 790.050 133.050 ;
        RECT 791.100 132.150 792.900 133.950 ;
        RECT 786.000 130.950 790.050 131.550 ;
        RECT 794.700 128.700 795.900 133.950 ;
        RECT 796.950 132.150 798.750 133.950 ;
        RECT 803.550 133.050 804.450 136.950 ;
        RECT 809.100 136.050 810.900 137.850 ;
        RECT 812.700 136.050 813.600 143.400 ;
        RECT 814.950 141.450 817.050 142.050 ;
        RECT 823.950 141.450 826.050 142.050 ;
        RECT 814.950 140.550 826.050 141.450 ;
        RECT 814.950 139.950 817.050 140.550 ;
        RECT 823.950 139.950 826.050 140.550 ;
        RECT 814.950 136.050 816.750 137.850 ;
        RECT 827.400 136.050 828.300 143.400 ;
        RECT 829.950 141.450 832.050 142.050 ;
        RECT 850.950 141.450 853.050 141.900 ;
        RECT 829.950 140.550 853.050 141.450 ;
        RECT 829.950 139.950 832.050 140.550 ;
        RECT 850.950 139.800 853.050 140.550 ;
        RECT 832.950 136.050 834.750 137.850 ;
        RECT 848.100 136.050 849.900 137.850 ;
        RECT 854.700 136.050 855.900 143.400 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 826.950 133.950 829.050 136.050 ;
        RECT 829.950 133.950 832.050 136.050 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 847.950 133.950 850.050 136.050 ;
        RECT 850.950 133.950 853.050 136.050 ;
        RECT 853.950 133.950 856.050 136.050 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 799.950 131.550 804.450 133.050 ;
        RECT 799.950 130.950 804.000 131.550 ;
        RECT 758.100 120.600 759.900 126.600 ;
        RECT 771.000 120.000 772.800 126.600 ;
        RECT 775.500 125.400 780.600 126.600 ;
        RECT 791.700 127.800 795.900 128.700 ;
        RECT 775.500 120.600 777.300 125.400 ;
        RECT 778.500 120.000 780.300 123.600 ;
        RECT 791.700 120.600 793.500 127.800 ;
        RECT 796.800 120.000 798.600 126.600 ;
        RECT 812.700 123.600 813.600 133.950 ;
        RECT 827.400 126.600 828.300 133.950 ;
        RECT 829.950 132.150 831.750 133.950 ;
        RECT 836.100 132.150 837.900 133.950 ;
        RECT 851.100 132.150 852.900 133.950 ;
        RECT 854.700 129.600 855.900 133.950 ;
        RECT 857.100 132.150 858.900 133.950 ;
        RECT 854.700 128.700 858.300 129.600 ;
        RECT 827.400 125.400 832.500 126.600 ;
        RECT 809.100 120.000 810.900 123.600 ;
        RECT 812.100 120.600 813.900 123.600 ;
        RECT 815.100 120.000 816.900 123.600 ;
        RECT 827.700 120.000 829.500 123.600 ;
        RECT 830.700 120.600 832.500 125.400 ;
        RECT 835.200 120.000 837.000 126.600 ;
        RECT 848.100 125.700 855.900 127.050 ;
        RECT 848.100 120.600 849.900 125.700 ;
        RECT 851.100 120.000 852.900 124.800 ;
        RECT 854.100 120.600 855.900 125.700 ;
        RECT 857.100 126.600 858.300 128.700 ;
        RECT 857.100 120.600 858.900 126.600 ;
        RECT 11.100 113.400 12.900 117.000 ;
        RECT 14.100 113.400 15.900 116.400 ;
        RECT 14.100 103.050 15.300 113.400 ;
        RECT 16.950 109.950 19.050 112.050 ;
        RECT 27.000 110.400 28.800 117.000 ;
        RECT 31.500 111.600 33.300 116.400 ;
        RECT 34.500 113.400 36.300 117.000 ;
        RECT 31.500 110.400 36.600 111.600 ;
        RECT 47.100 110.400 48.900 116.400 ;
        RECT 17.550 105.450 18.450 109.950 ;
        RECT 19.950 108.450 22.050 109.050 ;
        RECT 28.950 108.450 31.050 109.050 ;
        RECT 19.950 107.550 31.050 108.450 ;
        RECT 19.950 106.950 22.050 107.550 ;
        RECT 28.950 106.950 31.050 107.550 ;
        RECT 17.550 104.550 21.450 105.450 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 11.100 99.150 12.900 100.950 ;
        RECT 14.100 87.600 15.300 100.950 ;
        RECT 20.550 100.050 21.450 104.550 ;
        RECT 26.100 103.050 27.900 104.850 ;
        RECT 32.250 103.050 34.050 104.850 ;
        RECT 35.700 103.050 36.600 110.400 ;
        RECT 47.700 108.300 48.900 110.400 ;
        RECT 50.100 111.300 51.900 116.400 ;
        RECT 53.100 112.200 54.900 117.000 ;
        RECT 56.100 111.300 57.900 116.400 ;
        RECT 68.700 113.400 70.500 117.000 ;
        RECT 71.700 111.600 73.500 116.400 ;
        RECT 50.100 109.950 57.900 111.300 ;
        RECT 68.400 110.400 73.500 111.600 ;
        RECT 76.200 110.400 78.000 117.000 ;
        RECT 47.700 107.400 51.300 108.300 ;
        RECT 47.100 103.050 48.900 104.850 ;
        RECT 50.100 103.050 51.300 107.400 ;
        RECT 58.950 105.450 63.000 106.050 ;
        RECT 53.100 103.050 54.900 104.850 ;
        RECT 58.950 103.950 63.450 105.450 ;
        RECT 25.950 100.950 28.050 103.050 ;
        RECT 28.950 100.950 31.050 103.050 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 20.550 98.550 25.050 100.050 ;
        RECT 29.250 99.150 31.050 100.950 ;
        RECT 21.000 97.950 25.050 98.550 ;
        RECT 35.700 93.600 36.600 100.950 ;
        RECT 50.100 93.600 51.300 100.950 ;
        RECT 56.100 99.150 57.900 100.950 ;
        RECT 62.550 99.450 63.450 103.950 ;
        RECT 68.400 103.050 69.300 110.400 ;
        RECT 91.500 108.000 93.300 116.400 ;
        RECT 90.000 106.800 93.300 108.000 ;
        RECT 98.100 107.400 99.900 117.000 ;
        RECT 110.100 110.400 111.900 116.400 ;
        RECT 70.950 103.050 72.750 104.850 ;
        RECT 77.100 103.050 78.900 104.850 ;
        RECT 90.000 103.050 90.900 106.800 ;
        RECT 100.950 105.450 103.050 109.050 ;
        RECT 106.950 105.450 109.050 109.050 ;
        RECT 110.700 108.300 111.900 110.400 ;
        RECT 113.100 111.300 114.900 116.400 ;
        RECT 116.100 112.200 117.900 117.000 ;
        RECT 119.100 111.300 120.900 116.400 ;
        RECT 131.100 113.400 132.900 116.400 ;
        RECT 134.100 113.400 135.900 117.000 ;
        RECT 146.100 113.400 147.900 117.000 ;
        RECT 149.100 113.400 150.900 116.400 ;
        RECT 152.100 113.400 153.900 117.000 ;
        RECT 113.100 109.950 120.900 111.300 ;
        RECT 110.700 107.400 114.300 108.300 ;
        RECT 100.950 105.000 109.050 105.450 ;
        RECT 92.100 103.050 93.900 104.850 ;
        RECT 98.100 103.050 99.900 104.850 ;
        RECT 101.550 104.550 108.450 105.000 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 76.950 100.950 79.050 103.050 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 94.950 100.950 97.050 103.050 ;
        RECT 97.950 100.950 100.050 103.050 ;
        RECT 59.550 98.550 63.450 99.450 ;
        RECT 52.950 96.450 55.050 97.050 ;
        RECT 59.550 96.450 60.450 98.550 ;
        RECT 52.950 95.550 60.450 96.450 ;
        RECT 52.950 94.950 55.050 95.550 ;
        RECT 68.400 93.600 69.300 100.950 ;
        RECT 73.950 99.150 75.750 100.950 ;
        RECT 70.950 96.450 73.050 97.050 ;
        RECT 82.950 96.450 85.050 97.050 ;
        RECT 70.950 95.550 85.050 96.450 ;
        RECT 70.950 94.950 73.050 95.550 ;
        RECT 82.950 94.950 85.050 95.550 ;
        RECT 26.100 92.700 33.900 93.600 ;
        RECT 11.100 81.000 12.900 87.600 ;
        RECT 14.100 81.600 15.900 87.600 ;
        RECT 26.100 81.600 27.900 92.700 ;
        RECT 29.100 81.000 30.900 91.800 ;
        RECT 32.100 81.600 33.900 92.700 ;
        RECT 35.100 81.600 36.900 93.600 ;
        RECT 50.100 92.100 52.500 93.600 ;
        RECT 48.000 89.100 49.800 90.900 ;
        RECT 47.700 81.000 49.500 87.600 ;
        RECT 50.700 81.600 52.500 92.100 ;
        RECT 55.800 81.000 57.600 93.600 ;
        RECT 68.100 81.600 69.900 93.600 ;
        RECT 71.100 92.700 78.900 93.600 ;
        RECT 71.100 81.600 72.900 92.700 ;
        RECT 74.100 81.000 75.900 91.800 ;
        RECT 77.100 81.600 78.900 92.700 ;
        RECT 90.000 88.800 90.900 100.950 ;
        RECT 95.100 99.150 96.900 100.950 ;
        RECT 104.550 100.050 105.450 104.550 ;
        RECT 110.100 103.050 111.900 104.850 ;
        RECT 113.100 103.050 114.300 107.400 ;
        RECT 121.950 105.450 126.000 106.050 ;
        RECT 116.100 103.050 117.900 104.850 ;
        RECT 121.950 103.950 126.450 105.450 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 100.950 98.550 105.450 100.050 ;
        RECT 100.950 97.950 105.000 98.550 ;
        RECT 113.100 93.600 114.300 100.950 ;
        RECT 119.100 99.150 120.900 100.950 ;
        RECT 125.550 100.050 126.450 103.950 ;
        RECT 131.700 103.050 132.900 113.400 ;
        RECT 149.400 103.050 150.300 113.400 ;
        RECT 164.100 111.000 165.900 116.400 ;
        RECT 167.100 111.900 168.900 117.000 ;
        RECT 170.100 115.500 177.900 116.400 ;
        RECT 170.100 111.000 171.900 115.500 ;
        RECT 164.100 110.100 171.900 111.000 ;
        RECT 173.100 110.400 174.900 114.600 ;
        RECT 176.100 110.400 177.900 115.500 ;
        RECT 191.700 113.400 193.500 117.000 ;
        RECT 194.700 111.600 196.500 116.400 ;
        RECT 191.400 110.400 196.500 111.600 ;
        RECT 199.200 110.400 201.000 117.000 ;
        RECT 173.400 108.900 174.300 110.400 ;
        RECT 169.950 107.700 174.300 108.900 ;
        RECT 167.250 103.050 169.050 104.850 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 151.950 100.950 154.050 103.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 169.950 103.050 171.000 107.700 ;
        RECT 172.950 103.050 174.750 104.850 ;
        RECT 191.400 103.050 192.300 110.400 ;
        RECT 217.500 108.000 219.300 116.400 ;
        RECT 216.000 106.800 219.300 108.000 ;
        RECT 224.100 107.400 225.900 117.000 ;
        RECT 238.500 108.000 240.300 116.400 ;
        RECT 237.000 106.800 240.300 108.000 ;
        RECT 245.100 107.400 246.900 117.000 ;
        RECT 257.700 113.400 259.500 117.000 ;
        RECT 260.700 111.600 262.500 116.400 ;
        RECT 257.400 110.400 262.500 111.600 ;
        RECT 265.200 110.400 267.000 117.000 ;
        RECT 281.100 111.300 282.900 116.400 ;
        RECT 284.100 112.200 285.900 117.000 ;
        RECT 287.100 111.300 288.900 116.400 ;
        RECT 210.000 105.450 214.050 106.050 ;
        RECT 193.950 103.050 195.750 104.850 ;
        RECT 200.100 103.050 201.900 104.850 ;
        RECT 209.550 103.950 214.050 105.450 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 175.950 100.950 178.050 103.050 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 121.950 98.550 126.450 100.050 ;
        RECT 121.950 97.950 126.000 98.550 ;
        RECT 113.100 92.100 115.500 93.600 ;
        RECT 111.000 89.100 112.800 90.900 ;
        RECT 90.000 87.900 96.600 88.800 ;
        RECT 90.000 87.600 90.900 87.900 ;
        RECT 89.100 81.600 90.900 87.600 ;
        RECT 95.100 87.600 96.600 87.900 ;
        RECT 92.100 81.000 93.900 87.000 ;
        RECT 95.100 81.600 96.900 87.600 ;
        RECT 98.100 81.000 99.900 87.600 ;
        RECT 110.700 81.000 112.500 87.600 ;
        RECT 113.700 81.600 115.500 92.100 ;
        RECT 118.800 81.000 120.600 93.600 ;
        RECT 131.700 87.600 132.900 100.950 ;
        RECT 134.100 99.150 135.900 100.950 ;
        RECT 146.250 99.150 148.050 100.950 ;
        RECT 149.400 93.600 150.300 100.950 ;
        RECT 152.100 99.150 153.900 100.950 ;
        RECT 164.100 99.150 165.900 100.950 ;
        RECT 169.950 93.600 171.000 100.950 ;
        RECT 175.950 99.150 177.750 100.950 ;
        RECT 191.400 93.600 192.300 100.950 ;
        RECT 196.950 99.150 198.750 100.950 ;
        RECT 199.950 96.450 202.050 97.050 ;
        RECT 209.550 96.450 210.450 103.950 ;
        RECT 216.000 103.050 216.900 106.800 ;
        RECT 218.100 103.050 219.900 104.850 ;
        RECT 224.100 103.050 225.900 104.850 ;
        RECT 237.000 103.050 237.900 106.800 ;
        RECT 252.000 105.450 256.050 106.050 ;
        RECT 239.100 103.050 240.900 104.850 ;
        RECT 245.100 103.050 246.900 104.850 ;
        RECT 251.550 103.950 256.050 105.450 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 220.950 100.950 223.050 103.050 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 199.950 95.550 210.450 96.450 ;
        RECT 199.950 94.950 202.050 95.550 ;
        RECT 131.100 81.600 132.900 87.600 ;
        RECT 134.100 81.000 135.900 87.600 ;
        RECT 146.100 81.000 147.900 93.600 ;
        RECT 149.400 92.400 153.000 93.600 ;
        RECT 151.200 81.600 153.000 92.400 ;
        RECT 164.100 81.000 165.900 93.600 ;
        RECT 168.600 81.600 171.900 93.600 ;
        RECT 174.600 81.000 176.400 93.600 ;
        RECT 191.100 81.600 192.900 93.600 ;
        RECT 194.100 92.700 201.900 93.600 ;
        RECT 194.100 81.600 195.900 92.700 ;
        RECT 197.100 81.000 198.900 91.800 ;
        RECT 200.100 81.600 201.900 92.700 ;
        RECT 216.000 88.800 216.900 100.950 ;
        RECT 221.100 99.150 222.900 100.950 ;
        RECT 237.000 88.800 237.900 100.950 ;
        RECT 242.100 99.150 243.900 100.950 ;
        RECT 251.550 100.050 252.450 103.950 ;
        RECT 257.400 103.050 258.300 110.400 ;
        RECT 281.100 109.950 288.900 111.300 ;
        RECT 290.100 110.400 291.900 116.400 ;
        RECT 290.100 108.300 291.300 110.400 ;
        RECT 287.700 107.400 291.300 108.300 ;
        RECT 304.500 108.000 306.300 116.400 ;
        RECT 276.000 105.450 280.050 106.050 ;
        RECT 259.950 103.050 261.750 104.850 ;
        RECT 266.100 103.050 267.900 104.850 ;
        RECT 275.550 103.950 280.050 105.450 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 275.550 102.450 276.450 103.950 ;
        RECT 284.100 103.050 285.900 104.850 ;
        RECT 287.700 103.050 288.900 107.400 ;
        RECT 303.000 106.800 306.300 108.000 ;
        RECT 311.100 107.400 312.900 117.000 ;
        RECT 325.500 110.400 327.300 117.000 ;
        RECT 330.000 110.400 331.800 116.400 ;
        RECT 334.500 110.400 336.300 117.000 ;
        RECT 347.100 113.400 348.900 117.000 ;
        RECT 350.100 113.400 351.900 116.400 ;
        RECT 362.700 113.400 364.500 117.000 ;
        RECT 297.000 105.450 301.050 106.050 ;
        RECT 290.100 103.050 291.900 104.850 ;
        RECT 296.550 103.950 301.050 105.450 ;
        RECT 272.550 101.550 276.450 102.450 ;
        RECT 247.950 98.550 252.450 100.050 ;
        RECT 247.950 97.950 252.000 98.550 ;
        RECT 257.400 93.600 258.300 100.950 ;
        RECT 262.950 99.150 264.750 100.950 ;
        RECT 272.550 100.050 273.450 101.550 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 268.950 98.550 273.450 100.050 ;
        RECT 281.100 99.150 282.900 100.950 ;
        RECT 268.950 97.950 273.000 98.550 ;
        RECT 262.950 96.450 265.050 97.050 ;
        RECT 274.950 96.450 277.050 97.050 ;
        RECT 262.950 95.550 277.050 96.450 ;
        RECT 262.950 94.950 265.050 95.550 ;
        RECT 274.950 94.950 277.050 95.550 ;
        RECT 287.700 93.600 288.900 100.950 ;
        RECT 296.550 100.050 297.450 103.950 ;
        RECT 303.000 103.050 303.900 106.800 ;
        RECT 318.000 105.450 322.050 106.050 ;
        RECT 305.100 103.050 306.900 104.850 ;
        RECT 311.100 103.050 312.900 104.850 ;
        RECT 317.550 103.950 322.050 105.450 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 292.950 98.550 297.450 100.050 ;
        RECT 292.950 97.950 297.000 98.550 ;
        RECT 216.000 87.900 222.600 88.800 ;
        RECT 216.000 87.600 216.900 87.900 ;
        RECT 215.100 81.600 216.900 87.600 ;
        RECT 221.100 87.600 222.600 87.900 ;
        RECT 237.000 87.900 243.600 88.800 ;
        RECT 237.000 87.600 237.900 87.900 ;
        RECT 218.100 81.000 219.900 87.000 ;
        RECT 221.100 81.600 222.900 87.600 ;
        RECT 224.100 81.000 225.900 87.600 ;
        RECT 236.100 81.600 237.900 87.600 ;
        RECT 242.100 87.600 243.600 87.900 ;
        RECT 239.100 81.000 240.900 87.000 ;
        RECT 242.100 81.600 243.900 87.600 ;
        RECT 245.100 81.000 246.900 87.600 ;
        RECT 257.100 81.600 258.900 93.600 ;
        RECT 260.100 92.700 267.900 93.600 ;
        RECT 260.100 81.600 261.900 92.700 ;
        RECT 263.100 81.000 264.900 91.800 ;
        RECT 266.100 81.600 267.900 92.700 ;
        RECT 281.400 81.000 283.200 93.600 ;
        RECT 286.500 92.100 288.900 93.600 ;
        RECT 286.500 81.600 288.300 92.100 ;
        RECT 289.200 89.100 291.000 90.900 ;
        RECT 303.000 88.800 303.900 100.950 ;
        RECT 308.100 99.150 309.900 100.950 ;
        RECT 317.550 100.050 318.450 103.950 ;
        RECT 323.100 103.050 324.900 104.850 ;
        RECT 329.700 103.050 330.900 110.400 ;
        RECT 334.950 103.050 336.750 104.850 ;
        RECT 350.100 103.050 351.300 113.400 ;
        RECT 365.700 111.600 367.500 116.400 ;
        RECT 362.400 110.400 367.500 111.600 ;
        RECT 370.200 110.400 372.000 117.000 ;
        RECT 362.400 103.050 363.300 110.400 ;
        RECT 383.100 107.400 384.900 117.000 ;
        RECT 389.700 108.000 391.500 116.400 ;
        RECT 406.500 108.000 408.300 116.400 ;
        RECT 389.700 106.800 393.000 108.000 ;
        RECT 373.950 105.450 378.000 106.050 ;
        RECT 364.950 103.050 366.750 104.850 ;
        RECT 371.100 103.050 372.900 104.850 ;
        RECT 373.950 103.950 378.450 105.450 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 328.950 100.950 331.050 103.050 ;
        RECT 331.950 100.950 334.050 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 317.550 98.550 322.050 100.050 ;
        RECT 326.100 99.150 327.900 100.950 ;
        RECT 318.000 97.950 322.050 98.550 ;
        RECT 310.950 96.450 313.050 97.050 ;
        RECT 322.950 96.450 325.050 97.050 ;
        RECT 310.950 95.550 325.050 96.450 ;
        RECT 310.950 94.950 313.050 95.550 ;
        RECT 322.950 94.950 325.050 95.550 ;
        RECT 330.000 95.400 330.900 100.950 ;
        RECT 331.950 99.150 333.750 100.950 ;
        RECT 347.100 99.150 348.900 100.950 ;
        RECT 326.100 94.500 330.900 95.400 ;
        RECT 331.950 96.450 334.050 97.050 ;
        RECT 340.950 96.450 343.050 97.050 ;
        RECT 331.950 95.550 343.050 96.450 ;
        RECT 331.950 94.950 334.050 95.550 ;
        RECT 340.950 94.950 343.050 95.550 ;
        RECT 303.000 87.900 309.600 88.800 ;
        RECT 303.000 87.600 303.900 87.900 ;
        RECT 289.500 81.000 291.300 87.600 ;
        RECT 302.100 81.600 303.900 87.600 ;
        RECT 308.100 87.600 309.600 87.900 ;
        RECT 305.100 81.000 306.900 87.000 ;
        RECT 308.100 81.600 309.900 87.600 ;
        RECT 311.100 81.000 312.900 87.600 ;
        RECT 323.100 82.500 324.900 93.600 ;
        RECT 326.100 83.400 327.900 94.500 ;
        RECT 329.100 92.400 336.900 93.300 ;
        RECT 329.100 82.500 330.900 92.400 ;
        RECT 323.100 81.600 330.900 82.500 ;
        RECT 332.100 81.000 333.900 91.500 ;
        RECT 335.100 81.600 336.900 92.400 ;
        RECT 350.100 87.600 351.300 100.950 ;
        RECT 362.400 93.600 363.300 100.950 ;
        RECT 367.950 99.150 369.750 100.950 ;
        RECT 377.550 100.050 378.450 103.950 ;
        RECT 383.100 103.050 384.900 104.850 ;
        RECT 389.100 103.050 390.900 104.850 ;
        RECT 392.100 103.050 393.000 106.800 ;
        RECT 405.000 106.800 408.300 108.000 ;
        RECT 413.100 107.400 414.900 117.000 ;
        RECT 426.000 110.400 427.800 117.000 ;
        RECT 430.500 111.600 432.300 116.400 ;
        RECT 433.500 113.400 435.300 117.000 ;
        RECT 430.500 110.400 435.600 111.600 ;
        RECT 405.000 103.050 405.900 106.800 ;
        RECT 407.100 103.050 408.900 104.850 ;
        RECT 413.100 103.050 414.900 104.850 ;
        RECT 425.100 103.050 426.900 104.850 ;
        RECT 431.250 103.050 433.050 104.850 ;
        RECT 434.700 103.050 435.600 110.400 ;
        RECT 446.100 107.400 447.900 117.000 ;
        RECT 452.700 108.000 454.500 116.400 ;
        RECT 470.100 111.300 471.900 116.400 ;
        RECT 473.100 112.200 474.900 117.000 ;
        RECT 476.100 111.300 477.900 116.400 ;
        RECT 470.100 109.950 477.900 111.300 ;
        RECT 479.100 110.400 480.900 116.400 ;
        RECT 479.100 108.300 480.300 110.400 ;
        RECT 452.700 106.800 456.000 108.000 ;
        RECT 436.950 105.450 441.000 106.050 ;
        RECT 436.950 103.950 441.450 105.450 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 403.950 100.950 406.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 377.550 98.550 382.050 100.050 ;
        RECT 386.100 99.150 387.900 100.950 ;
        RECT 378.000 97.950 382.050 98.550 ;
        RECT 370.950 96.450 373.050 97.050 ;
        RECT 388.950 96.450 391.050 97.050 ;
        RECT 370.950 95.550 391.050 96.450 ;
        RECT 370.950 94.950 373.050 95.550 ;
        RECT 388.950 94.950 391.050 95.550 ;
        RECT 347.100 81.000 348.900 87.600 ;
        RECT 350.100 81.600 351.900 87.600 ;
        RECT 362.100 81.600 363.900 93.600 ;
        RECT 365.100 92.700 372.900 93.600 ;
        RECT 365.100 81.600 366.900 92.700 ;
        RECT 368.100 81.000 369.900 91.800 ;
        RECT 371.100 81.600 372.900 92.700 ;
        RECT 392.100 88.800 393.000 100.950 ;
        RECT 386.400 87.900 393.000 88.800 ;
        RECT 386.400 87.600 387.900 87.900 ;
        RECT 383.100 81.000 384.900 87.600 ;
        RECT 386.100 81.600 387.900 87.600 ;
        RECT 392.100 87.600 393.000 87.900 ;
        RECT 405.000 88.800 405.900 100.950 ;
        RECT 410.100 99.150 411.900 100.950 ;
        RECT 428.250 99.150 430.050 100.950 ;
        RECT 434.700 93.600 435.600 100.950 ;
        RECT 440.550 99.450 441.450 103.950 ;
        RECT 446.100 103.050 447.900 104.850 ;
        RECT 452.100 103.050 453.900 104.850 ;
        RECT 455.100 103.050 456.000 106.800 ;
        RECT 476.700 107.400 480.300 108.300 ;
        RECT 493.500 108.000 495.300 116.400 ;
        RECT 457.950 105.450 462.000 106.050 ;
        RECT 457.950 103.950 462.450 105.450 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 448.950 100.950 451.050 103.050 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 440.550 98.550 444.450 99.450 ;
        RECT 449.100 99.150 450.900 100.950 ;
        RECT 443.550 96.450 444.450 98.550 ;
        RECT 451.950 96.450 454.050 96.750 ;
        RECT 443.550 95.550 454.050 96.450 ;
        RECT 451.950 94.650 454.050 95.550 ;
        RECT 425.100 92.700 432.900 93.600 ;
        RECT 405.000 87.900 411.600 88.800 ;
        RECT 405.000 87.600 405.900 87.900 ;
        RECT 389.100 81.000 390.900 87.000 ;
        RECT 392.100 81.600 393.900 87.600 ;
        RECT 404.100 81.600 405.900 87.600 ;
        RECT 410.100 87.600 411.600 87.900 ;
        RECT 407.100 81.000 408.900 87.000 ;
        RECT 410.100 81.600 411.900 87.600 ;
        RECT 413.100 81.000 414.900 87.600 ;
        RECT 425.100 81.600 426.900 92.700 ;
        RECT 428.100 81.000 429.900 91.800 ;
        RECT 431.100 81.600 432.900 92.700 ;
        RECT 434.100 81.600 435.900 93.600 ;
        RECT 455.100 88.800 456.000 100.950 ;
        RECT 461.550 100.050 462.450 103.950 ;
        RECT 473.100 103.050 474.900 104.850 ;
        RECT 476.700 103.050 477.900 107.400 ;
        RECT 492.000 106.800 495.300 108.000 ;
        RECT 500.100 107.400 501.900 117.000 ;
        RECT 512.100 113.400 513.900 116.400 ;
        RECT 515.100 113.400 516.900 117.000 ;
        RECT 481.950 105.450 486.000 106.050 ;
        RECT 479.100 103.050 480.900 104.850 ;
        RECT 481.950 103.950 486.450 105.450 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 457.950 98.550 462.450 100.050 ;
        RECT 470.100 99.150 471.900 100.950 ;
        RECT 457.950 97.950 462.000 98.550 ;
        RECT 476.700 93.600 477.900 100.950 ;
        RECT 485.550 100.050 486.450 103.950 ;
        RECT 492.000 103.050 492.900 106.800 ;
        RECT 507.000 105.450 511.050 106.050 ;
        RECT 494.100 103.050 495.900 104.850 ;
        RECT 500.100 103.050 501.900 104.850 ;
        RECT 506.550 103.950 511.050 105.450 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 496.950 100.950 499.050 103.050 ;
        RECT 499.950 100.950 502.050 103.050 ;
        RECT 481.950 98.550 486.450 100.050 ;
        RECT 481.950 97.950 486.000 98.550 ;
        RECT 449.400 87.900 456.000 88.800 ;
        RECT 449.400 87.600 450.900 87.900 ;
        RECT 446.100 81.000 447.900 87.600 ;
        RECT 449.100 81.600 450.900 87.600 ;
        RECT 455.100 87.600 456.000 87.900 ;
        RECT 452.100 81.000 453.900 87.000 ;
        RECT 455.100 81.600 456.900 87.600 ;
        RECT 470.400 81.000 472.200 93.600 ;
        RECT 475.500 92.100 477.900 93.600 ;
        RECT 475.500 81.600 477.300 92.100 ;
        RECT 478.200 89.100 480.000 90.900 ;
        RECT 492.000 88.800 492.900 100.950 ;
        RECT 497.100 99.150 498.900 100.950 ;
        RECT 506.550 100.050 507.450 103.950 ;
        RECT 512.700 103.050 513.900 113.400 ;
        RECT 529.500 110.400 531.300 117.000 ;
        RECT 534.000 110.400 535.800 116.400 ;
        RECT 538.500 110.400 540.300 117.000 ;
        RECT 551.400 110.400 553.200 117.000 ;
        RECT 517.950 105.450 522.000 106.050 ;
        RECT 517.950 103.950 522.450 105.450 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 502.950 98.550 507.450 100.050 ;
        RECT 502.950 97.950 507.000 98.550 ;
        RECT 492.000 87.900 498.600 88.800 ;
        RECT 492.000 87.600 492.900 87.900 ;
        RECT 478.500 81.000 480.300 87.600 ;
        RECT 491.100 81.600 492.900 87.600 ;
        RECT 497.100 87.600 498.600 87.900 ;
        RECT 512.700 87.600 513.900 100.950 ;
        RECT 515.100 99.150 516.900 100.950 ;
        RECT 521.550 100.050 522.450 103.950 ;
        RECT 527.100 103.050 528.900 104.850 ;
        RECT 533.700 103.050 534.900 110.400 ;
        RECT 556.500 109.200 558.300 116.400 ;
        RECT 569.400 110.400 571.200 117.000 ;
        RECT 574.500 109.200 576.300 116.400 ;
        RECT 587.400 110.400 589.200 117.000 ;
        RECT 592.500 109.200 594.300 116.400 ;
        RECT 608.100 110.400 609.900 116.400 ;
        RECT 554.100 108.300 558.300 109.200 ;
        RECT 572.100 108.300 576.300 109.200 ;
        RECT 590.100 108.300 594.300 109.200 ;
        RECT 608.700 108.300 609.900 110.400 ;
        RECT 611.100 111.300 612.900 116.400 ;
        RECT 614.100 112.200 615.900 117.000 ;
        RECT 617.100 111.300 618.900 116.400 ;
        RECT 611.100 109.950 618.900 111.300 ;
        RECT 629.100 111.300 630.900 116.400 ;
        RECT 632.100 112.200 633.900 117.000 ;
        RECT 635.100 111.300 636.900 116.400 ;
        RECT 629.100 109.950 636.900 111.300 ;
        RECT 638.100 110.400 639.900 116.400 ;
        RECT 650.700 113.400 652.500 117.000 ;
        RECT 653.700 111.600 655.500 116.400 ;
        RECT 650.400 110.400 655.500 111.600 ;
        RECT 658.200 110.400 660.000 117.000 ;
        RECT 638.100 108.300 639.300 110.400 ;
        RECT 538.950 103.050 540.750 104.850 ;
        RECT 551.250 103.050 553.050 104.850 ;
        RECT 554.100 103.050 555.300 108.300 ;
        RECT 557.100 103.050 558.900 104.850 ;
        RECT 569.250 103.050 571.050 104.850 ;
        RECT 572.100 103.050 573.300 108.300 ;
        RECT 575.100 103.050 576.900 104.850 ;
        RECT 587.250 103.050 589.050 104.850 ;
        RECT 590.100 103.050 591.300 108.300 ;
        RECT 608.700 107.400 612.300 108.300 ;
        RECT 593.100 103.050 594.900 104.850 ;
        RECT 608.100 103.050 609.900 104.850 ;
        RECT 611.100 103.050 612.300 107.400 ;
        RECT 635.700 107.400 639.300 108.300 ;
        RECT 614.100 103.050 615.900 104.850 ;
        RECT 632.100 103.050 633.900 104.850 ;
        RECT 635.700 103.050 636.900 107.400 ;
        RECT 638.100 103.050 639.900 104.850 ;
        RECT 650.400 103.050 651.300 110.400 ;
        RECT 671.100 107.400 672.900 117.000 ;
        RECT 677.700 108.000 679.500 116.400 ;
        RECT 692.100 110.400 693.900 116.400 ;
        RECT 692.700 108.300 693.900 110.400 ;
        RECT 695.100 111.300 696.900 116.400 ;
        RECT 698.100 112.200 699.900 117.000 ;
        RECT 701.100 111.300 702.900 116.400 ;
        RECT 713.700 113.400 715.500 117.000 ;
        RECT 716.700 111.600 718.500 116.400 ;
        RECT 695.100 109.950 702.900 111.300 ;
        RECT 713.400 110.400 718.500 111.600 ;
        RECT 721.200 110.400 723.000 117.000 ;
        RECT 677.700 106.800 681.000 108.000 ;
        RECT 692.700 107.400 696.300 108.300 ;
        RECT 666.000 105.450 670.050 106.050 ;
        RECT 652.950 103.050 654.750 104.850 ;
        RECT 659.100 103.050 660.900 104.850 ;
        RECT 665.550 103.950 670.050 105.450 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 568.950 100.950 571.050 103.050 ;
        RECT 571.950 100.950 574.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 586.950 100.950 589.050 103.050 ;
        RECT 589.950 100.950 592.050 103.050 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 610.950 100.950 613.050 103.050 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 631.950 100.950 634.050 103.050 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 517.950 98.550 522.450 100.050 ;
        RECT 530.100 99.150 531.900 100.950 ;
        RECT 517.950 97.950 522.000 98.550 ;
        RECT 534.000 95.400 534.900 100.950 ;
        RECT 535.950 99.150 537.750 100.950 ;
        RECT 530.100 94.500 534.900 95.400 ;
        RECT 494.100 81.000 495.900 87.000 ;
        RECT 497.100 81.600 498.900 87.600 ;
        RECT 500.100 81.000 501.900 87.600 ;
        RECT 512.100 81.600 513.900 87.600 ;
        RECT 515.100 81.000 516.900 87.600 ;
        RECT 527.100 82.500 528.900 93.600 ;
        RECT 530.100 83.400 531.900 94.500 ;
        RECT 533.100 92.400 540.900 93.300 ;
        RECT 533.100 82.500 534.900 92.400 ;
        RECT 527.100 81.600 534.900 82.500 ;
        RECT 536.100 81.000 537.900 91.500 ;
        RECT 539.100 81.600 540.900 92.400 ;
        RECT 554.100 87.600 555.300 100.950 ;
        RECT 572.100 87.600 573.300 100.950 ;
        RECT 590.100 87.600 591.300 100.950 ;
        RECT 592.950 96.450 595.050 97.050 ;
        RECT 598.950 96.450 601.050 97.050 ;
        RECT 592.950 95.550 601.050 96.450 ;
        RECT 592.950 94.950 595.050 95.550 ;
        RECT 598.950 94.950 601.050 95.550 ;
        RECT 611.100 93.600 612.300 100.950 ;
        RECT 617.100 99.150 618.900 100.950 ;
        RECT 629.100 99.150 630.900 100.950 ;
        RECT 613.950 96.450 616.050 97.050 ;
        RECT 622.950 96.450 625.050 97.050 ;
        RECT 631.950 96.450 634.050 97.050 ;
        RECT 613.950 95.550 634.050 96.450 ;
        RECT 613.950 94.950 616.050 95.550 ;
        RECT 622.950 94.950 625.050 95.550 ;
        RECT 631.950 94.950 634.050 95.550 ;
        RECT 635.700 93.600 636.900 100.950 ;
        RECT 650.400 93.600 651.300 100.950 ;
        RECT 655.950 99.150 657.750 100.950 ;
        RECT 665.550 100.050 666.450 103.950 ;
        RECT 671.100 103.050 672.900 104.850 ;
        RECT 677.100 103.050 678.900 104.850 ;
        RECT 680.100 103.050 681.000 106.800 ;
        RECT 692.100 103.050 693.900 104.850 ;
        RECT 695.100 103.050 696.300 107.400 ;
        RECT 698.100 103.050 699.900 104.850 ;
        RECT 713.400 103.050 714.300 110.400 ;
        RECT 734.100 107.400 735.900 117.000 ;
        RECT 740.700 108.000 742.500 116.400 ;
        RECT 755.100 110.400 756.900 116.400 ;
        RECT 755.700 108.300 756.900 110.400 ;
        RECT 758.100 111.300 759.900 116.400 ;
        RECT 761.100 112.200 762.900 117.000 ;
        RECT 764.100 111.300 765.900 116.400 ;
        RECT 758.100 109.950 765.900 111.300 ;
        RECT 776.100 111.300 777.900 116.400 ;
        RECT 779.100 112.200 780.900 117.000 ;
        RECT 782.100 111.300 783.900 116.400 ;
        RECT 776.100 109.950 783.900 111.300 ;
        RECT 785.100 110.400 786.900 116.400 ;
        RECT 797.700 113.400 799.500 117.000 ;
        RECT 800.700 111.600 802.500 116.400 ;
        RECT 797.400 110.400 802.500 111.600 ;
        RECT 805.200 110.400 807.000 117.000 ;
        RECT 785.100 108.300 786.300 110.400 ;
        RECT 740.700 106.800 744.000 108.000 ;
        RECT 755.700 107.400 759.300 108.300 ;
        RECT 715.950 103.050 717.750 104.850 ;
        RECT 722.100 103.050 723.900 104.850 ;
        RECT 734.100 103.050 735.900 104.850 ;
        RECT 740.100 103.050 741.900 104.850 ;
        RECT 743.100 103.050 744.000 106.800 ;
        RECT 755.100 103.050 756.900 104.850 ;
        RECT 758.100 103.050 759.300 107.400 ;
        RECT 782.700 107.400 786.300 108.300 ;
        RECT 771.000 105.450 775.050 106.050 ;
        RECT 761.100 103.050 762.900 104.850 ;
        RECT 770.550 103.950 775.050 105.450 ;
        RECT 670.950 100.950 673.050 103.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 742.950 100.950 745.050 103.050 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 760.950 100.950 763.050 103.050 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 661.950 98.550 666.450 100.050 ;
        RECT 674.100 99.150 675.900 100.950 ;
        RECT 661.950 97.950 666.000 98.550 ;
        RECT 652.950 96.450 655.050 97.050 ;
        RECT 670.950 96.450 673.050 97.050 ;
        RECT 652.950 95.550 673.050 96.450 ;
        RECT 652.950 94.950 655.050 95.550 ;
        RECT 670.950 94.950 673.050 95.550 ;
        RECT 611.100 92.100 613.500 93.600 ;
        RECT 609.000 89.100 610.800 90.900 ;
        RECT 551.100 81.000 552.900 87.600 ;
        RECT 554.100 81.600 555.900 87.600 ;
        RECT 557.100 81.000 558.900 87.600 ;
        RECT 569.100 81.000 570.900 87.600 ;
        RECT 572.100 81.600 573.900 87.600 ;
        RECT 575.100 81.000 576.900 87.600 ;
        RECT 587.100 81.000 588.900 87.600 ;
        RECT 590.100 81.600 591.900 87.600 ;
        RECT 593.100 81.000 594.900 87.600 ;
        RECT 608.700 81.000 610.500 87.600 ;
        RECT 611.700 81.600 613.500 92.100 ;
        RECT 616.800 81.000 618.600 93.600 ;
        RECT 629.400 81.000 631.200 93.600 ;
        RECT 634.500 92.100 636.900 93.600 ;
        RECT 634.500 81.600 636.300 92.100 ;
        RECT 637.200 89.100 639.000 90.900 ;
        RECT 637.500 81.000 639.300 87.600 ;
        RECT 650.100 81.600 651.900 93.600 ;
        RECT 653.100 92.700 660.900 93.600 ;
        RECT 653.100 81.600 654.900 92.700 ;
        RECT 656.100 81.000 657.900 91.800 ;
        RECT 659.100 81.600 660.900 92.700 ;
        RECT 680.100 88.800 681.000 100.950 ;
        RECT 695.100 93.600 696.300 100.950 ;
        RECT 701.100 99.150 702.900 100.950 ;
        RECT 713.400 93.600 714.300 100.950 ;
        RECT 718.950 99.150 720.750 100.950 ;
        RECT 737.100 99.150 738.900 100.950 ;
        RECT 695.100 92.100 697.500 93.600 ;
        RECT 693.000 89.100 694.800 90.900 ;
        RECT 674.400 87.900 681.000 88.800 ;
        RECT 674.400 87.600 675.900 87.900 ;
        RECT 671.100 81.000 672.900 87.600 ;
        RECT 674.100 81.600 675.900 87.600 ;
        RECT 680.100 87.600 681.000 87.900 ;
        RECT 677.100 81.000 678.900 87.000 ;
        RECT 680.100 81.600 681.900 87.600 ;
        RECT 692.700 81.000 694.500 87.600 ;
        RECT 695.700 81.600 697.500 92.100 ;
        RECT 700.800 81.000 702.600 93.600 ;
        RECT 713.100 81.600 714.900 93.600 ;
        RECT 716.100 92.700 723.900 93.600 ;
        RECT 716.100 81.600 717.900 92.700 ;
        RECT 719.100 81.000 720.900 91.800 ;
        RECT 722.100 81.600 723.900 92.700 ;
        RECT 743.100 88.800 744.000 100.950 ;
        RECT 758.100 93.600 759.300 100.950 ;
        RECT 764.100 99.150 765.900 100.950 ;
        RECT 770.550 100.050 771.450 103.950 ;
        RECT 779.100 103.050 780.900 104.850 ;
        RECT 782.700 103.050 783.900 107.400 ;
        RECT 785.100 103.050 786.900 104.850 ;
        RECT 797.400 103.050 798.300 110.400 ;
        RECT 818.100 107.400 819.900 117.000 ;
        RECT 824.700 108.000 826.500 116.400 ;
        RECT 841.500 108.000 843.300 116.400 ;
        RECT 824.700 106.800 828.000 108.000 ;
        RECT 813.000 105.450 817.050 106.050 ;
        RECT 799.950 103.050 801.750 104.850 ;
        RECT 806.100 103.050 807.900 104.850 ;
        RECT 812.550 103.950 817.050 105.450 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 770.550 98.550 775.050 100.050 ;
        RECT 776.100 99.150 777.900 100.950 ;
        RECT 771.000 97.950 775.050 98.550 ;
        RECT 782.700 93.600 783.900 100.950 ;
        RECT 797.400 93.600 798.300 100.950 ;
        RECT 802.950 99.150 804.750 100.950 ;
        RECT 812.550 99.450 813.450 103.950 ;
        RECT 818.100 103.050 819.900 104.850 ;
        RECT 824.100 103.050 825.900 104.850 ;
        RECT 827.100 103.050 828.000 106.800 ;
        RECT 840.000 106.800 843.300 108.000 ;
        RECT 848.100 107.400 849.900 117.000 ;
        RECT 860.100 113.400 861.900 116.400 ;
        RECT 863.100 113.400 864.900 117.000 ;
        RECT 829.950 105.450 834.000 106.050 ;
        RECT 829.950 103.950 834.450 105.450 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 809.550 98.550 813.450 99.450 ;
        RECT 821.100 99.150 822.900 100.950 ;
        RECT 799.950 96.450 802.050 97.050 ;
        RECT 809.550 96.450 810.450 98.550 ;
        RECT 799.950 95.550 810.450 96.450 ;
        RECT 799.950 94.950 802.050 95.550 ;
        RECT 758.100 92.100 760.500 93.600 ;
        RECT 756.000 89.100 757.800 90.900 ;
        RECT 737.400 87.900 744.000 88.800 ;
        RECT 737.400 87.600 738.900 87.900 ;
        RECT 734.100 81.000 735.900 87.600 ;
        RECT 737.100 81.600 738.900 87.600 ;
        RECT 743.100 87.600 744.000 87.900 ;
        RECT 740.100 81.000 741.900 87.000 ;
        RECT 743.100 81.600 744.900 87.600 ;
        RECT 755.700 81.000 757.500 87.600 ;
        RECT 758.700 81.600 760.500 92.100 ;
        RECT 763.800 81.000 765.600 93.600 ;
        RECT 776.400 81.000 778.200 93.600 ;
        RECT 781.500 92.100 783.900 93.600 ;
        RECT 781.500 81.600 783.300 92.100 ;
        RECT 784.200 89.100 786.000 90.900 ;
        RECT 784.500 81.000 786.300 87.600 ;
        RECT 797.100 81.600 798.900 93.600 ;
        RECT 800.100 92.700 807.900 93.600 ;
        RECT 800.100 81.600 801.900 92.700 ;
        RECT 803.100 81.000 804.900 91.800 ;
        RECT 806.100 81.600 807.900 92.700 ;
        RECT 827.100 88.800 828.000 100.950 ;
        RECT 833.550 100.050 834.450 103.950 ;
        RECT 840.000 103.050 840.900 106.800 ;
        RECT 842.100 103.050 843.900 104.850 ;
        RECT 848.100 103.050 849.900 104.850 ;
        RECT 860.700 103.050 861.900 113.400 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 859.950 100.950 862.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 829.950 98.550 834.450 100.050 ;
        RECT 829.950 97.950 834.000 98.550 ;
        RECT 821.400 87.900 828.000 88.800 ;
        RECT 821.400 87.600 822.900 87.900 ;
        RECT 818.100 81.000 819.900 87.600 ;
        RECT 821.100 81.600 822.900 87.600 ;
        RECT 827.100 87.600 828.000 87.900 ;
        RECT 840.000 88.800 840.900 100.950 ;
        RECT 845.100 99.150 846.900 100.950 ;
        RECT 840.000 87.900 846.600 88.800 ;
        RECT 840.000 87.600 840.900 87.900 ;
        RECT 824.100 81.000 825.900 87.000 ;
        RECT 827.100 81.600 828.900 87.600 ;
        RECT 839.100 81.600 840.900 87.600 ;
        RECT 845.100 87.600 846.600 87.900 ;
        RECT 860.700 87.600 861.900 100.950 ;
        RECT 863.100 99.150 864.900 100.950 ;
        RECT 842.100 81.000 843.900 87.000 ;
        RECT 845.100 81.600 846.900 87.600 ;
        RECT 848.100 81.000 849.900 87.600 ;
        RECT 860.100 81.600 861.900 87.600 ;
        RECT 863.100 81.000 864.900 87.600 ;
        RECT 14.100 71.400 15.900 77.400 ;
        RECT 17.100 72.000 18.900 78.000 ;
        RECT 15.000 71.100 15.900 71.400 ;
        RECT 20.100 71.400 21.900 77.400 ;
        RECT 23.100 71.400 24.900 78.000 ;
        RECT 35.100 71.400 36.900 77.400 ;
        RECT 38.100 72.000 39.900 78.000 ;
        RECT 20.100 71.100 21.600 71.400 ;
        RECT 15.000 70.200 21.600 71.100 ;
        RECT 36.000 71.100 36.900 71.400 ;
        RECT 41.100 71.400 42.900 77.400 ;
        RECT 44.100 71.400 45.900 78.000 ;
        RECT 59.100 71.400 60.900 77.400 ;
        RECT 62.100 72.000 63.900 78.000 ;
        RECT 41.100 71.100 42.600 71.400 ;
        RECT 36.000 70.200 42.600 71.100 ;
        RECT 60.000 71.100 60.900 71.400 ;
        RECT 65.100 71.400 66.900 77.400 ;
        RECT 68.100 71.400 69.900 78.000 ;
        RECT 80.700 71.400 82.500 78.000 ;
        RECT 65.100 71.100 66.600 71.400 ;
        RECT 60.000 70.200 66.600 71.100 ;
        RECT 15.000 58.050 15.900 70.200 ;
        RECT 30.000 60.450 34.050 61.050 ;
        RECT 20.100 58.050 21.900 59.850 ;
        RECT 29.550 58.950 34.050 60.450 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 15.000 52.200 15.900 55.950 ;
        RECT 17.100 54.150 18.900 55.950 ;
        RECT 23.100 54.150 24.900 55.950 ;
        RECT 29.550 55.050 30.450 58.950 ;
        RECT 36.000 58.050 36.900 70.200 ;
        RECT 37.950 63.450 40.050 64.050 ;
        RECT 52.950 63.450 55.050 64.050 ;
        RECT 37.950 62.550 55.050 63.450 ;
        RECT 37.950 61.950 40.050 62.550 ;
        RECT 52.950 61.950 55.050 62.550 ;
        RECT 41.100 58.050 42.900 59.850 ;
        RECT 60.000 58.050 60.900 70.200 ;
        RECT 81.000 68.100 82.800 69.900 ;
        RECT 83.700 66.900 85.500 77.400 ;
        RECT 83.100 65.400 85.500 66.900 ;
        RECT 88.800 65.400 90.600 78.000 ;
        RECT 101.700 71.400 103.500 78.000 ;
        RECT 102.000 68.100 103.800 69.900 ;
        RECT 104.700 66.900 106.500 77.400 ;
        RECT 104.100 65.400 106.500 66.900 ;
        RECT 109.800 65.400 111.600 78.000 ;
        RECT 122.100 71.400 123.900 77.400 ;
        RECT 125.100 72.000 126.900 78.000 ;
        RECT 123.000 71.100 123.900 71.400 ;
        RECT 128.100 71.400 129.900 77.400 ;
        RECT 131.100 71.400 132.900 78.000 ;
        RECT 128.100 71.100 129.600 71.400 ;
        RECT 123.000 70.200 129.600 71.100 ;
        RECT 65.100 58.050 66.900 59.850 ;
        RECT 83.100 58.050 84.300 65.400 ;
        RECT 89.100 58.050 90.900 59.850 ;
        RECT 104.100 58.050 105.300 65.400 ;
        RECT 110.100 58.050 111.900 59.850 ;
        RECT 123.000 58.050 123.900 70.200 ;
        RECT 143.100 65.400 144.900 77.400 ;
        RECT 146.100 66.300 147.900 77.400 ;
        RECT 149.100 67.200 150.900 78.000 ;
        RECT 152.100 66.300 153.900 77.400 ;
        RECT 164.700 71.400 166.500 78.000 ;
        RECT 165.000 68.100 166.800 69.900 ;
        RECT 167.700 66.900 169.500 77.400 ;
        RECT 146.100 65.400 153.900 66.300 ;
        RECT 167.100 65.400 169.500 66.900 ;
        RECT 172.800 65.400 174.600 78.000 ;
        RECT 185.700 71.400 187.500 78.000 ;
        RECT 186.000 68.100 187.800 69.900 ;
        RECT 188.700 66.900 190.500 77.400 ;
        RECT 188.100 65.400 190.500 66.900 ;
        RECT 193.800 65.400 195.600 78.000 ;
        RECT 206.100 71.400 207.900 78.000 ;
        RECT 209.100 71.400 210.900 77.400 ;
        RECT 212.100 72.000 213.900 78.000 ;
        RECT 209.400 71.100 210.900 71.400 ;
        RECT 215.100 71.400 216.900 77.400 ;
        RECT 215.100 71.100 216.000 71.400 ;
        RECT 209.400 70.200 216.000 71.100 ;
        RECT 124.950 63.450 127.050 64.050 ;
        RECT 133.950 63.450 136.050 64.050 ;
        RECT 124.950 62.550 136.050 63.450 ;
        RECT 124.950 61.950 127.050 62.550 ;
        RECT 133.950 61.950 136.050 62.550 ;
        RECT 128.100 58.050 129.900 59.850 ;
        RECT 143.400 58.050 144.300 65.400 ;
        RECT 148.950 58.050 150.750 59.850 ;
        RECT 167.100 58.050 168.300 65.400 ;
        RECT 175.950 63.450 178.050 64.050 ;
        RECT 181.950 63.450 184.050 64.050 ;
        RECT 175.950 62.550 184.050 63.450 ;
        RECT 175.950 61.950 178.050 62.550 ;
        RECT 181.950 61.950 184.050 62.550 ;
        RECT 173.100 58.050 174.900 59.850 ;
        RECT 188.100 58.050 189.300 65.400 ;
        RECT 194.100 58.050 195.900 59.850 ;
        RECT 209.100 58.050 210.900 59.850 ;
        RECT 215.100 58.050 216.000 70.200 ;
        RECT 227.100 66.300 228.900 77.400 ;
        RECT 230.100 67.200 231.900 78.000 ;
        RECT 233.100 66.300 234.900 77.400 ;
        RECT 227.100 65.400 234.900 66.300 ;
        RECT 236.100 65.400 237.900 77.400 ;
        RECT 248.400 65.400 250.200 78.000 ;
        RECT 253.500 66.900 255.300 77.400 ;
        RECT 256.500 71.400 258.300 78.000 ;
        RECT 269.100 71.400 270.900 78.000 ;
        RECT 272.100 71.400 273.900 77.400 ;
        RECT 256.200 68.100 258.000 69.900 ;
        RECT 253.500 65.400 255.900 66.900 ;
        RECT 229.950 63.450 232.050 64.050 ;
        RECT 224.550 62.550 232.050 63.450 ;
        RECT 224.550 60.450 225.450 62.550 ;
        RECT 229.950 61.950 232.050 62.550 ;
        RECT 221.550 59.550 225.450 60.450 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 43.950 55.950 46.050 58.050 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 29.550 53.550 34.050 55.050 ;
        RECT 30.000 52.950 34.050 53.550 ;
        RECT 36.000 52.200 36.900 55.950 ;
        RECT 38.100 54.150 39.900 55.950 ;
        RECT 44.100 54.150 45.900 55.950 ;
        RECT 60.000 52.200 60.900 55.950 ;
        RECT 62.100 54.150 63.900 55.950 ;
        RECT 68.100 54.150 69.900 55.950 ;
        RECT 80.100 54.150 81.900 55.950 ;
        RECT 15.000 51.000 18.300 52.200 ;
        RECT 16.500 42.600 18.300 51.000 ;
        RECT 23.100 42.000 24.900 51.600 ;
        RECT 36.000 51.000 39.300 52.200 ;
        RECT 37.500 42.600 39.300 51.000 ;
        RECT 44.100 42.000 45.900 51.600 ;
        RECT 60.000 51.000 63.300 52.200 ;
        RECT 83.100 51.600 84.300 55.950 ;
        RECT 86.100 54.150 87.900 55.950 ;
        RECT 101.100 54.150 102.900 55.950 ;
        RECT 104.100 51.600 105.300 55.950 ;
        RECT 107.100 54.150 108.900 55.950 ;
        RECT 61.500 42.600 63.300 51.000 ;
        RECT 68.100 42.000 69.900 51.600 ;
        RECT 80.700 50.700 84.300 51.600 ;
        RECT 101.700 50.700 105.300 51.600 ;
        RECT 123.000 52.200 123.900 55.950 ;
        RECT 125.100 54.150 126.900 55.950 ;
        RECT 131.100 54.150 132.900 55.950 ;
        RECT 123.000 51.000 126.300 52.200 ;
        RECT 80.700 48.600 81.900 50.700 ;
        RECT 80.100 42.600 81.900 48.600 ;
        RECT 83.100 47.700 90.900 49.050 ;
        RECT 101.700 48.600 102.900 50.700 ;
        RECT 83.100 42.600 84.900 47.700 ;
        RECT 86.100 42.000 87.900 46.800 ;
        RECT 89.100 42.600 90.900 47.700 ;
        RECT 101.100 42.600 102.900 48.600 ;
        RECT 104.100 47.700 111.900 49.050 ;
        RECT 104.100 42.600 105.900 47.700 ;
        RECT 107.100 42.000 108.900 46.800 ;
        RECT 110.100 42.600 111.900 47.700 ;
        RECT 124.500 42.600 126.300 51.000 ;
        RECT 131.100 42.000 132.900 51.600 ;
        RECT 143.400 48.600 144.300 55.950 ;
        RECT 145.950 54.150 147.750 55.950 ;
        RECT 152.100 54.150 153.900 55.950 ;
        RECT 164.100 54.150 165.900 55.950 ;
        RECT 167.100 51.600 168.300 55.950 ;
        RECT 170.100 54.150 171.900 55.950 ;
        RECT 185.100 54.150 186.900 55.950 ;
        RECT 188.100 51.600 189.300 55.950 ;
        RECT 191.100 54.150 192.900 55.950 ;
        RECT 206.100 54.150 207.900 55.950 ;
        RECT 212.100 54.150 213.900 55.950 ;
        RECT 215.100 52.200 216.000 55.950 ;
        RECT 221.550 55.050 222.450 59.550 ;
        RECT 230.250 58.050 232.050 59.850 ;
        RECT 236.700 58.050 237.600 65.400 ;
        RECT 250.950 63.450 253.050 64.050 ;
        RECT 245.550 62.550 253.050 63.450 ;
        RECT 245.550 60.450 246.450 62.550 ;
        RECT 250.950 61.950 253.050 62.550 ;
        RECT 242.550 59.550 246.450 60.450 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 217.950 53.550 222.450 55.050 ;
        RECT 227.100 54.150 228.900 55.950 ;
        RECT 233.250 54.150 235.050 55.950 ;
        RECT 217.950 52.950 222.000 53.550 ;
        RECT 164.700 50.700 168.300 51.600 ;
        RECT 185.700 50.700 189.300 51.600 ;
        RECT 164.700 48.600 165.900 50.700 ;
        RECT 143.400 47.400 148.500 48.600 ;
        RECT 143.700 42.000 145.500 45.600 ;
        RECT 146.700 42.600 148.500 47.400 ;
        RECT 151.200 42.000 153.000 48.600 ;
        RECT 164.100 42.600 165.900 48.600 ;
        RECT 167.100 47.700 174.900 49.050 ;
        RECT 185.700 48.600 186.900 50.700 ;
        RECT 167.100 42.600 168.900 47.700 ;
        RECT 170.100 42.000 171.900 46.800 ;
        RECT 173.100 42.600 174.900 47.700 ;
        RECT 185.100 42.600 186.900 48.600 ;
        RECT 188.100 47.700 195.900 49.050 ;
        RECT 188.100 42.600 189.900 47.700 ;
        RECT 191.100 42.000 192.900 46.800 ;
        RECT 194.100 42.600 195.900 47.700 ;
        RECT 206.100 42.000 207.900 51.600 ;
        RECT 212.700 51.000 216.000 52.200 ;
        RECT 212.700 42.600 214.500 51.000 ;
        RECT 236.700 48.600 237.600 55.950 ;
        RECT 242.550 55.050 243.450 59.550 ;
        RECT 248.100 58.050 249.900 59.850 ;
        RECT 254.700 58.050 255.900 65.400 ;
        RECT 269.100 58.050 270.900 59.850 ;
        RECT 272.100 58.050 273.300 71.400 ;
        RECT 284.100 66.300 285.900 77.400 ;
        RECT 287.100 67.200 288.900 78.000 ;
        RECT 290.100 66.300 291.900 77.400 ;
        RECT 284.100 65.400 291.900 66.300 ;
        RECT 293.100 65.400 294.900 77.400 ;
        RECT 308.100 71.400 309.900 77.400 ;
        RECT 311.100 72.000 312.900 78.000 ;
        RECT 309.000 71.100 309.900 71.400 ;
        RECT 314.100 71.400 315.900 77.400 ;
        RECT 317.100 71.400 318.900 78.000 ;
        RECT 314.100 71.100 315.600 71.400 ;
        RECT 309.000 70.200 315.600 71.100 ;
        RECT 274.950 60.450 279.000 61.050 ;
        RECT 274.950 58.950 279.450 60.450 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 238.950 53.550 243.450 55.050 ;
        RECT 251.100 54.150 252.900 55.950 ;
        RECT 238.950 52.950 243.000 53.550 ;
        RECT 254.700 51.600 255.900 55.950 ;
        RECT 257.100 54.150 258.900 55.950 ;
        RECT 254.700 50.700 258.300 51.600 ;
        RECT 228.000 42.000 229.800 48.600 ;
        RECT 232.500 47.400 237.600 48.600 ;
        RECT 248.100 47.700 255.900 49.050 ;
        RECT 232.500 42.600 234.300 47.400 ;
        RECT 235.500 42.000 237.300 45.600 ;
        RECT 248.100 42.600 249.900 47.700 ;
        RECT 251.100 42.000 252.900 46.800 ;
        RECT 254.100 42.600 255.900 47.700 ;
        RECT 257.100 48.600 258.300 50.700 ;
        RECT 257.100 42.600 258.900 48.600 ;
        RECT 272.100 45.600 273.300 55.950 ;
        RECT 278.550 55.050 279.450 58.950 ;
        RECT 287.250 58.050 289.050 59.850 ;
        RECT 293.700 58.050 294.600 65.400 ;
        RECT 309.000 58.050 309.900 70.200 ;
        RECT 329.100 66.300 330.900 77.400 ;
        RECT 332.100 67.200 333.900 78.000 ;
        RECT 335.100 66.300 336.900 77.400 ;
        RECT 329.100 65.400 336.900 66.300 ;
        RECT 338.100 65.400 339.900 77.400 ;
        RECT 350.700 71.400 352.500 78.000 ;
        RECT 351.000 68.100 352.800 69.900 ;
        RECT 353.700 66.900 355.500 77.400 ;
        RECT 353.100 65.400 355.500 66.900 ;
        RECT 358.800 65.400 360.600 78.000 ;
        RECT 371.400 65.400 373.200 78.000 ;
        RECT 376.500 66.900 378.300 77.400 ;
        RECT 379.500 71.400 381.300 78.000 ;
        RECT 392.100 71.400 393.900 77.400 ;
        RECT 395.100 72.000 396.900 78.000 ;
        RECT 393.000 71.100 393.900 71.400 ;
        RECT 398.100 71.400 399.900 77.400 ;
        RECT 401.100 71.400 402.900 78.000 ;
        RECT 413.100 71.400 414.900 77.400 ;
        RECT 416.100 72.000 417.900 78.000 ;
        RECT 398.100 71.100 399.600 71.400 ;
        RECT 393.000 70.200 399.600 71.100 ;
        RECT 414.000 71.100 414.900 71.400 ;
        RECT 419.100 71.400 420.900 77.400 ;
        RECT 422.100 71.400 423.900 78.000 ;
        RECT 419.100 71.100 420.600 71.400 ;
        RECT 414.000 70.200 420.600 71.100 ;
        RECT 379.200 68.100 381.000 69.900 ;
        RECT 376.500 65.400 378.900 66.900 ;
        RECT 316.950 63.450 319.050 64.050 ;
        RECT 334.950 63.450 337.050 64.050 ;
        RECT 316.950 62.550 337.050 63.450 ;
        RECT 316.950 61.950 319.050 62.550 ;
        RECT 334.950 61.950 337.050 62.550 ;
        RECT 314.100 58.050 315.900 59.850 ;
        RECT 332.250 58.050 334.050 59.850 ;
        RECT 338.700 58.050 339.600 65.400 ;
        RECT 345.000 60.450 349.050 61.050 ;
        RECT 344.550 58.950 349.050 60.450 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 274.950 53.550 279.450 55.050 ;
        RECT 284.100 54.150 285.900 55.950 ;
        RECT 290.250 54.150 292.050 55.950 ;
        RECT 274.950 52.950 279.000 53.550 ;
        RECT 293.700 48.600 294.600 55.950 ;
        RECT 309.000 52.200 309.900 55.950 ;
        RECT 311.100 54.150 312.900 55.950 ;
        RECT 317.100 54.150 318.900 55.950 ;
        RECT 329.100 54.150 330.900 55.950 ;
        RECT 335.250 54.150 337.050 55.950 ;
        RECT 309.000 51.000 312.300 52.200 ;
        RECT 269.100 42.000 270.900 45.600 ;
        RECT 272.100 42.600 273.900 45.600 ;
        RECT 285.000 42.000 286.800 48.600 ;
        RECT 289.500 47.400 294.600 48.600 ;
        RECT 289.500 42.600 291.300 47.400 ;
        RECT 292.500 42.000 294.300 45.600 ;
        RECT 310.500 42.600 312.300 51.000 ;
        RECT 317.100 42.000 318.900 51.600 ;
        RECT 338.700 48.600 339.600 55.950 ;
        RECT 344.550 55.050 345.450 58.950 ;
        RECT 353.100 58.050 354.300 65.400 ;
        RECT 359.100 58.050 360.900 59.850 ;
        RECT 371.100 58.050 372.900 59.850 ;
        RECT 377.700 58.050 378.900 65.400 ;
        RECT 393.000 58.050 393.900 70.200 ;
        RECT 398.100 58.050 399.900 59.850 ;
        RECT 414.000 58.050 414.900 70.200 ;
        RECT 434.100 65.400 435.900 77.400 ;
        RECT 437.100 66.300 438.900 77.400 ;
        RECT 440.100 67.200 441.900 78.000 ;
        RECT 443.100 66.300 444.900 77.400 ;
        RECT 437.100 65.400 444.900 66.300 ;
        RECT 455.100 65.400 456.900 77.400 ;
        RECT 458.100 66.300 459.900 77.400 ;
        RECT 461.100 67.200 462.900 78.000 ;
        RECT 464.100 66.300 465.900 77.400 ;
        RECT 479.100 71.400 480.900 77.400 ;
        RECT 482.100 72.000 483.900 78.000 ;
        RECT 458.100 65.400 465.900 66.300 ;
        RECT 480.000 71.100 480.900 71.400 ;
        RECT 485.100 71.400 486.900 77.400 ;
        RECT 488.100 71.400 489.900 78.000 ;
        RECT 500.100 71.400 501.900 78.000 ;
        RECT 503.100 71.400 504.900 77.400 ;
        RECT 485.100 71.100 486.600 71.400 ;
        RECT 480.000 70.200 486.600 71.100 ;
        RECT 419.100 58.050 420.900 59.850 ;
        RECT 434.400 58.050 435.300 65.400 ;
        RECT 445.950 60.450 450.000 61.050 ;
        RECT 439.950 58.050 441.750 59.850 ;
        RECT 445.950 58.950 450.450 60.450 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 355.950 55.950 358.050 58.050 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 400.950 55.950 403.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 344.550 53.550 349.050 55.050 ;
        RECT 350.100 54.150 351.900 55.950 ;
        RECT 345.000 52.950 349.050 53.550 ;
        RECT 353.100 51.600 354.300 55.950 ;
        RECT 356.100 54.150 357.900 55.950 ;
        RECT 374.100 54.150 375.900 55.950 ;
        RECT 350.700 50.700 354.300 51.600 ;
        RECT 377.700 51.600 378.900 55.950 ;
        RECT 380.100 54.150 381.900 55.950 ;
        RECT 393.000 52.200 393.900 55.950 ;
        RECT 395.100 54.150 396.900 55.950 ;
        RECT 401.100 54.150 402.900 55.950 ;
        RECT 414.000 52.200 414.900 55.950 ;
        RECT 416.100 54.150 417.900 55.950 ;
        RECT 422.100 54.150 423.900 55.950 ;
        RECT 377.700 50.700 381.300 51.600 ;
        RECT 393.000 51.000 396.300 52.200 ;
        RECT 350.700 48.600 351.900 50.700 ;
        RECT 330.000 42.000 331.800 48.600 ;
        RECT 334.500 47.400 339.600 48.600 ;
        RECT 334.500 42.600 336.300 47.400 ;
        RECT 337.500 42.000 339.300 45.600 ;
        RECT 350.100 42.600 351.900 48.600 ;
        RECT 353.100 47.700 360.900 49.050 ;
        RECT 353.100 42.600 354.900 47.700 ;
        RECT 356.100 42.000 357.900 46.800 ;
        RECT 359.100 42.600 360.900 47.700 ;
        RECT 371.100 47.700 378.900 49.050 ;
        RECT 371.100 42.600 372.900 47.700 ;
        RECT 374.100 42.000 375.900 46.800 ;
        RECT 377.100 42.600 378.900 47.700 ;
        RECT 380.100 48.600 381.300 50.700 ;
        RECT 380.100 42.600 381.900 48.600 ;
        RECT 394.500 42.600 396.300 51.000 ;
        RECT 401.100 42.000 402.900 51.600 ;
        RECT 414.000 51.000 417.300 52.200 ;
        RECT 415.500 42.600 417.300 51.000 ;
        RECT 422.100 42.000 423.900 51.600 ;
        RECT 434.400 48.600 435.300 55.950 ;
        RECT 436.950 54.150 438.750 55.950 ;
        RECT 443.100 54.150 444.900 55.950 ;
        RECT 449.550 55.050 450.450 58.950 ;
        RECT 455.400 58.050 456.300 65.400 ;
        RECT 460.950 63.450 463.050 64.050 ;
        RECT 460.950 62.550 468.450 63.450 ;
        RECT 460.950 61.950 463.050 62.550 ;
        RECT 467.550 60.450 468.450 62.550 ;
        RECT 460.950 58.050 462.750 59.850 ;
        RECT 467.550 59.550 471.450 60.450 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 445.950 53.550 450.450 55.050 ;
        RECT 445.950 52.950 450.000 53.550 ;
        RECT 455.400 48.600 456.300 55.950 ;
        RECT 457.950 54.150 459.750 55.950 ;
        RECT 464.100 54.150 465.900 55.950 ;
        RECT 463.950 51.450 466.050 52.050 ;
        RECT 470.550 51.450 471.450 59.550 ;
        RECT 480.000 58.050 480.900 70.200 ;
        RECT 485.100 58.050 486.900 59.850 ;
        RECT 500.100 58.050 501.900 59.850 ;
        RECT 503.100 58.050 504.300 71.400 ;
        RECT 515.100 66.300 516.900 77.400 ;
        RECT 518.100 67.200 519.900 78.000 ;
        RECT 521.100 66.300 522.900 77.400 ;
        RECT 515.100 65.400 522.900 66.300 ;
        RECT 524.100 65.400 525.900 77.400 ;
        RECT 536.100 71.400 537.900 78.000 ;
        RECT 539.100 71.400 540.900 77.400 ;
        RECT 542.100 71.400 543.900 78.000 ;
        RECT 554.100 71.400 555.900 77.400 ;
        RECT 557.100 72.000 558.900 78.000 ;
        RECT 518.250 58.050 520.050 59.850 ;
        RECT 524.700 58.050 525.600 65.400 ;
        RECT 539.700 58.050 540.900 71.400 ;
        RECT 555.000 71.100 555.900 71.400 ;
        RECT 560.100 71.400 561.900 77.400 ;
        RECT 563.100 71.400 564.900 78.000 ;
        RECT 575.100 71.400 576.900 78.000 ;
        RECT 578.100 71.400 579.900 77.400 ;
        RECT 560.100 71.100 561.600 71.400 ;
        RECT 555.000 70.200 561.600 71.100 ;
        RECT 555.000 58.050 555.900 70.200 ;
        RECT 560.100 58.050 561.900 59.850 ;
        RECT 575.100 58.050 576.900 59.850 ;
        RECT 578.100 58.050 579.300 71.400 ;
        RECT 593.400 65.400 595.200 78.000 ;
        RECT 598.500 66.900 600.300 77.400 ;
        RECT 601.500 71.400 603.300 78.000 ;
        RECT 601.200 68.100 603.000 69.900 ;
        RECT 598.500 65.400 600.900 66.900 ;
        RECT 614.100 65.400 615.900 77.400 ;
        RECT 617.100 66.300 618.900 77.400 ;
        RECT 620.100 67.200 621.900 78.000 ;
        RECT 623.100 66.300 624.900 77.400 ;
        RECT 635.100 71.400 636.900 77.400 ;
        RECT 638.100 72.000 639.900 78.000 ;
        RECT 617.100 65.400 624.900 66.300 ;
        RECT 636.000 71.100 636.900 71.400 ;
        RECT 641.100 71.400 642.900 77.400 ;
        RECT 644.100 71.400 645.900 78.000 ;
        RECT 659.100 71.400 660.900 78.000 ;
        RECT 662.100 71.400 663.900 77.400 ;
        RECT 665.100 72.000 666.900 78.000 ;
        RECT 641.100 71.100 642.600 71.400 ;
        RECT 636.000 70.200 642.600 71.100 ;
        RECT 662.400 71.100 663.900 71.400 ;
        RECT 668.100 71.400 669.900 77.400 ;
        RECT 680.100 71.400 681.900 77.400 ;
        RECT 683.100 72.000 684.900 78.000 ;
        RECT 668.100 71.100 669.000 71.400 ;
        RECT 662.400 70.200 669.000 71.100 ;
        RECT 593.100 58.050 594.900 59.850 ;
        RECT 599.700 58.050 600.900 65.400 ;
        RECT 614.400 58.050 615.300 65.400 ;
        RECT 619.950 58.050 621.750 59.850 ;
        RECT 636.000 58.050 636.900 70.200 ;
        RECT 641.100 58.050 642.900 59.850 ;
        RECT 662.100 58.050 663.900 59.850 ;
        RECT 668.100 58.050 669.000 70.200 ;
        RECT 681.000 71.100 681.900 71.400 ;
        RECT 686.100 71.400 687.900 77.400 ;
        RECT 689.100 71.400 690.900 78.000 ;
        RECT 686.100 71.100 687.600 71.400 ;
        RECT 681.000 70.200 687.600 71.100 ;
        RECT 681.000 58.050 681.900 70.200 ;
        RECT 701.100 66.300 702.900 77.400 ;
        RECT 704.100 67.200 705.900 78.000 ;
        RECT 707.100 66.300 708.900 77.400 ;
        RECT 701.100 65.400 708.900 66.300 ;
        RECT 710.100 65.400 711.900 77.400 ;
        RECT 722.100 71.400 723.900 78.000 ;
        RECT 725.100 71.400 726.900 77.400 ;
        RECT 728.100 71.400 729.900 78.000 ;
        RECT 740.100 71.400 741.900 78.000 ;
        RECT 743.100 71.400 744.900 77.400 ;
        RECT 758.100 71.400 759.900 78.000 ;
        RECT 761.100 71.400 762.900 77.400 ;
        RECT 764.100 72.000 765.900 78.000 ;
        RECT 682.950 63.450 685.050 64.050 ;
        RECT 700.950 63.450 703.050 64.050 ;
        RECT 682.950 62.550 703.050 63.450 ;
        RECT 682.950 61.950 685.050 62.550 ;
        RECT 700.950 61.950 703.050 62.550 ;
        RECT 686.100 58.050 687.900 59.850 ;
        RECT 704.250 58.050 706.050 59.850 ;
        RECT 710.700 58.050 711.600 65.400 ;
        RECT 725.700 58.050 726.900 71.400 ;
        RECT 740.100 58.050 741.900 59.850 ;
        RECT 743.100 58.050 744.300 71.400 ;
        RECT 761.400 71.100 762.900 71.400 ;
        RECT 767.100 71.400 768.900 77.400 ;
        RECT 767.100 71.100 768.000 71.400 ;
        RECT 761.400 70.200 768.000 71.100 ;
        RECT 761.100 58.050 762.900 59.850 ;
        RECT 767.100 58.050 768.000 70.200 ;
        RECT 779.400 65.400 781.200 78.000 ;
        RECT 784.500 66.900 786.300 77.400 ;
        RECT 787.500 71.400 789.300 78.000 ;
        RECT 787.200 68.100 789.000 69.900 ;
        RECT 784.500 65.400 786.900 66.900 ;
        RECT 800.100 65.400 801.900 77.400 ;
        RECT 803.100 66.300 804.900 77.400 ;
        RECT 806.100 67.200 807.900 78.000 ;
        RECT 809.100 66.300 810.900 77.400 ;
        RECT 821.700 71.400 823.500 78.000 ;
        RECT 822.000 68.100 823.800 69.900 ;
        RECT 824.700 66.900 826.500 77.400 ;
        RECT 803.100 65.400 810.900 66.300 ;
        RECT 824.100 65.400 826.500 66.900 ;
        RECT 829.800 65.400 831.600 78.000 ;
        RECT 842.100 65.400 843.900 77.400 ;
        RECT 845.100 66.300 846.900 77.400 ;
        RECT 848.100 67.200 849.900 78.000 ;
        RECT 851.100 66.300 852.900 77.400 ;
        RECT 863.100 71.400 864.900 77.400 ;
        RECT 866.100 71.400 867.900 78.000 ;
        RECT 845.100 65.400 852.900 66.300 ;
        RECT 769.950 60.450 772.050 64.050 ;
        RECT 769.950 60.000 774.450 60.450 ;
        RECT 770.550 59.550 774.450 60.000 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 481.950 55.950 484.050 58.050 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 517.950 55.950 520.050 58.050 ;
        RECT 520.950 55.950 523.050 58.050 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 556.950 55.950 559.050 58.050 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 667.950 55.950 670.050 58.050 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 700.950 55.950 703.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 721.950 55.950 724.050 58.050 ;
        RECT 724.950 55.950 727.050 58.050 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 739.950 55.950 742.050 58.050 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 463.950 50.550 471.450 51.450 ;
        RECT 480.000 52.200 480.900 55.950 ;
        RECT 482.100 54.150 483.900 55.950 ;
        RECT 488.100 54.150 489.900 55.950 ;
        RECT 480.000 51.000 483.300 52.200 ;
        RECT 463.950 49.950 466.050 50.550 ;
        RECT 469.950 48.900 474.000 49.050 ;
        RECT 434.400 47.400 439.500 48.600 ;
        RECT 434.700 42.000 436.500 45.600 ;
        RECT 437.700 42.600 439.500 47.400 ;
        RECT 442.200 42.000 444.000 48.600 ;
        RECT 455.400 47.400 460.500 48.600 ;
        RECT 455.700 42.000 457.500 45.600 ;
        RECT 458.700 42.600 460.500 47.400 ;
        RECT 463.200 42.000 465.000 48.600 ;
        RECT 469.950 46.950 475.050 48.900 ;
        RECT 472.950 46.800 475.050 46.950 ;
        RECT 481.500 42.600 483.300 51.000 ;
        RECT 488.100 42.000 489.900 51.600 ;
        RECT 503.100 45.600 504.300 55.950 ;
        RECT 515.100 54.150 516.900 55.950 ;
        RECT 521.250 54.150 523.050 55.950 ;
        RECT 508.950 51.450 511.050 52.050 ;
        RECT 517.950 51.450 520.050 51.750 ;
        RECT 508.950 50.550 520.050 51.450 ;
        RECT 508.950 49.950 511.050 50.550 ;
        RECT 517.950 49.650 520.050 50.550 ;
        RECT 524.700 48.600 525.600 55.950 ;
        RECT 536.100 54.150 537.900 55.950 ;
        RECT 539.700 50.700 540.900 55.950 ;
        RECT 541.950 54.150 543.750 55.950 ;
        RECT 555.000 52.200 555.900 55.950 ;
        RECT 557.100 54.150 558.900 55.950 ;
        RECT 563.100 54.150 564.900 55.950 ;
        RECT 555.000 51.000 558.300 52.200 ;
        RECT 500.100 42.000 501.900 45.600 ;
        RECT 503.100 42.600 504.900 45.600 ;
        RECT 516.000 42.000 517.800 48.600 ;
        RECT 520.500 47.400 525.600 48.600 ;
        RECT 536.700 49.800 540.900 50.700 ;
        RECT 520.500 42.600 522.300 47.400 ;
        RECT 523.500 42.000 525.300 45.600 ;
        RECT 536.700 42.600 538.500 49.800 ;
        RECT 541.800 42.000 543.600 48.600 ;
        RECT 556.500 42.600 558.300 51.000 ;
        RECT 563.100 42.000 564.900 51.600 ;
        RECT 578.100 45.600 579.300 55.950 ;
        RECT 596.100 54.150 597.900 55.950 ;
        RECT 599.700 51.600 600.900 55.950 ;
        RECT 602.100 54.150 603.900 55.950 ;
        RECT 599.700 50.700 603.300 51.600 ;
        RECT 593.100 47.700 600.900 49.050 ;
        RECT 575.100 42.000 576.900 45.600 ;
        RECT 578.100 42.600 579.900 45.600 ;
        RECT 593.100 42.600 594.900 47.700 ;
        RECT 596.100 42.000 597.900 46.800 ;
        RECT 599.100 42.600 600.900 47.700 ;
        RECT 602.100 48.600 603.300 50.700 ;
        RECT 614.400 48.600 615.300 55.950 ;
        RECT 616.950 54.150 618.750 55.950 ;
        RECT 623.100 54.150 624.900 55.950 ;
        RECT 636.000 52.200 636.900 55.950 ;
        RECT 638.100 54.150 639.900 55.950 ;
        RECT 644.100 54.150 645.900 55.950 ;
        RECT 659.100 54.150 660.900 55.950 ;
        RECT 665.100 54.150 666.900 55.950 ;
        RECT 668.100 52.200 669.000 55.950 ;
        RECT 636.000 51.000 639.300 52.200 ;
        RECT 602.100 42.600 603.900 48.600 ;
        RECT 614.400 47.400 619.500 48.600 ;
        RECT 614.700 42.000 616.500 45.600 ;
        RECT 617.700 42.600 619.500 47.400 ;
        RECT 622.200 42.000 624.000 48.600 ;
        RECT 637.500 42.600 639.300 51.000 ;
        RECT 644.100 42.000 645.900 51.600 ;
        RECT 659.100 42.000 660.900 51.600 ;
        RECT 665.700 51.000 669.000 52.200 ;
        RECT 681.000 52.200 681.900 55.950 ;
        RECT 683.100 54.150 684.900 55.950 ;
        RECT 689.100 54.150 690.900 55.950 ;
        RECT 701.100 54.150 702.900 55.950 ;
        RECT 707.250 54.150 709.050 55.950 ;
        RECT 681.000 51.000 684.300 52.200 ;
        RECT 665.700 42.600 667.500 51.000 ;
        RECT 682.500 42.600 684.300 51.000 ;
        RECT 689.100 42.000 690.900 51.600 ;
        RECT 710.700 48.600 711.600 55.950 ;
        RECT 722.100 54.150 723.900 55.950 ;
        RECT 725.700 50.700 726.900 55.950 ;
        RECT 727.950 54.150 729.750 55.950 ;
        RECT 702.000 42.000 703.800 48.600 ;
        RECT 706.500 47.400 711.600 48.600 ;
        RECT 722.700 49.800 726.900 50.700 ;
        RECT 706.500 42.600 708.300 47.400 ;
        RECT 709.500 42.000 711.300 45.600 ;
        RECT 722.700 42.600 724.500 49.800 ;
        RECT 727.800 42.000 729.600 48.600 ;
        RECT 743.100 45.600 744.300 55.950 ;
        RECT 758.100 54.150 759.900 55.950 ;
        RECT 764.100 54.150 765.900 55.950 ;
        RECT 767.100 52.200 768.000 55.950 ;
        RECT 773.550 55.050 774.450 59.550 ;
        RECT 779.100 58.050 780.900 59.850 ;
        RECT 785.700 58.050 786.900 65.400 ;
        RECT 800.400 58.050 801.300 65.400 ;
        RECT 814.950 61.950 817.050 64.050 ;
        RECT 805.950 58.050 807.750 59.850 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 769.950 53.550 774.450 55.050 ;
        RECT 782.100 54.150 783.900 55.950 ;
        RECT 769.950 52.950 774.000 53.550 ;
        RECT 740.100 42.000 741.900 45.600 ;
        RECT 743.100 42.600 744.900 45.600 ;
        RECT 758.100 42.000 759.900 51.600 ;
        RECT 764.700 51.000 768.000 52.200 ;
        RECT 785.700 51.600 786.900 55.950 ;
        RECT 788.100 54.150 789.900 55.950 ;
        RECT 764.700 42.600 766.500 51.000 ;
        RECT 785.700 50.700 789.300 51.600 ;
        RECT 779.100 47.700 786.900 49.050 ;
        RECT 779.100 42.600 780.900 47.700 ;
        RECT 782.100 42.000 783.900 46.800 ;
        RECT 785.100 42.600 786.900 47.700 ;
        RECT 788.100 48.600 789.300 50.700 ;
        RECT 800.400 48.600 801.300 55.950 ;
        RECT 802.950 54.150 804.750 55.950 ;
        RECT 809.100 54.150 810.900 55.950 ;
        RECT 815.550 54.450 816.450 61.950 ;
        RECT 824.100 58.050 825.300 65.400 ;
        RECT 830.100 58.050 831.900 59.850 ;
        RECT 842.400 58.050 843.300 65.400 ;
        RECT 847.950 58.050 849.750 59.850 ;
        RECT 863.700 58.050 864.900 71.400 ;
        RECT 866.100 58.050 867.900 59.850 ;
        RECT 820.950 55.950 823.050 58.050 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 844.950 55.950 847.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 812.550 53.550 816.450 54.450 ;
        RECT 821.100 54.150 822.900 55.950 ;
        RECT 805.950 51.450 808.050 52.050 ;
        RECT 812.550 51.450 813.450 53.550 ;
        RECT 824.100 51.600 825.300 55.950 ;
        RECT 827.100 54.150 828.900 55.950 ;
        RECT 805.950 50.550 813.450 51.450 ;
        RECT 821.700 50.700 825.300 51.600 ;
        RECT 805.950 49.950 808.050 50.550 ;
        RECT 821.700 48.600 822.900 50.700 ;
        RECT 788.100 42.600 789.900 48.600 ;
        RECT 800.400 47.400 805.500 48.600 ;
        RECT 800.700 42.000 802.500 45.600 ;
        RECT 803.700 42.600 805.500 47.400 ;
        RECT 808.200 42.000 810.000 48.600 ;
        RECT 821.100 42.600 822.900 48.600 ;
        RECT 824.100 47.700 831.900 49.050 ;
        RECT 824.100 42.600 825.900 47.700 ;
        RECT 827.100 42.000 828.900 46.800 ;
        RECT 830.100 42.600 831.900 47.700 ;
        RECT 842.400 48.600 843.300 55.950 ;
        RECT 844.950 54.150 846.750 55.950 ;
        RECT 851.100 54.150 852.900 55.950 ;
        RECT 842.400 47.400 847.500 48.600 ;
        RECT 842.700 42.000 844.500 45.600 ;
        RECT 845.700 42.600 847.500 47.400 ;
        RECT 850.200 42.000 852.000 48.600 ;
        RECT 863.700 45.600 864.900 55.950 ;
        RECT 863.100 42.600 864.900 45.600 ;
        RECT 866.100 42.000 867.900 45.600 ;
        RECT 14.100 35.400 15.900 39.000 ;
        RECT 17.100 35.400 18.900 38.400 ;
        RECT 29.100 35.400 30.900 39.000 ;
        RECT 32.100 35.400 33.900 38.400 ;
        RECT 17.100 25.050 18.300 35.400 ;
        RECT 32.100 25.050 33.300 35.400 ;
        RECT 45.000 32.400 46.800 39.000 ;
        RECT 49.500 33.600 51.300 38.400 ;
        RECT 52.500 35.400 54.300 39.000 ;
        RECT 49.500 32.400 54.600 33.600 ;
        RECT 44.100 25.050 45.900 26.850 ;
        RECT 50.250 25.050 52.050 26.850 ;
        RECT 53.700 25.050 54.600 32.400 ;
        RECT 67.500 30.000 69.300 38.400 ;
        RECT 66.000 28.800 69.300 30.000 ;
        RECT 74.100 29.400 75.900 39.000 ;
        RECT 87.000 32.400 88.800 39.000 ;
        RECT 91.500 33.600 93.300 38.400 ;
        RECT 94.500 35.400 96.300 39.000 ;
        RECT 91.500 32.400 96.600 33.600 ;
        RECT 107.100 32.400 108.900 38.400 ;
        RECT 66.000 25.050 66.900 28.800 ;
        RECT 68.100 25.050 69.900 26.850 ;
        RECT 74.100 25.050 75.900 26.850 ;
        RECT 86.100 25.050 87.900 26.850 ;
        RECT 92.250 25.050 94.050 26.850 ;
        RECT 95.700 25.050 96.600 32.400 ;
        RECT 107.700 30.300 108.900 32.400 ;
        RECT 110.100 33.300 111.900 38.400 ;
        RECT 113.100 34.200 114.900 39.000 ;
        RECT 116.100 33.300 117.900 38.400 ;
        RECT 128.700 35.400 130.500 39.000 ;
        RECT 131.700 33.600 133.500 38.400 ;
        RECT 110.100 31.950 117.900 33.300 ;
        RECT 128.400 32.400 133.500 33.600 ;
        RECT 136.200 32.400 138.000 39.000 ;
        RECT 107.700 29.400 111.300 30.300 ;
        RECT 107.100 25.050 108.900 26.850 ;
        RECT 110.100 25.050 111.300 29.400 ;
        RECT 113.100 25.050 114.900 26.850 ;
        RECT 128.400 25.050 129.300 32.400 ;
        RECT 151.500 30.000 153.300 38.400 ;
        RECT 150.000 28.800 153.300 30.000 ;
        RECT 158.100 29.400 159.900 39.000 ;
        RECT 170.100 35.400 171.900 39.000 ;
        RECT 173.100 35.400 174.900 38.400 ;
        RECT 130.950 25.050 132.750 26.850 ;
        RECT 137.100 25.050 138.900 26.850 ;
        RECT 150.000 25.050 150.900 28.800 ;
        RECT 165.000 27.450 169.050 28.050 ;
        RECT 152.100 25.050 153.900 26.850 ;
        RECT 158.100 25.050 159.900 26.850 ;
        RECT 164.550 25.950 169.050 27.450 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 28.950 22.950 31.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 43.950 22.950 46.050 25.050 ;
        RECT 46.950 22.950 49.050 25.050 ;
        RECT 49.950 22.950 52.050 25.050 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 115.950 22.950 118.050 25.050 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 14.100 21.150 15.900 22.950 ;
        RECT 17.100 9.600 18.300 22.950 ;
        RECT 29.100 21.150 30.900 22.950 ;
        RECT 32.100 9.600 33.300 22.950 ;
        RECT 47.250 21.150 49.050 22.950 ;
        RECT 53.700 15.600 54.600 22.950 ;
        RECT 44.100 14.700 51.900 15.600 ;
        RECT 14.100 3.000 15.900 9.600 ;
        RECT 17.100 3.600 18.900 9.600 ;
        RECT 29.100 3.000 30.900 9.600 ;
        RECT 32.100 3.600 33.900 9.600 ;
        RECT 44.100 3.600 45.900 14.700 ;
        RECT 47.100 3.000 48.900 13.800 ;
        RECT 50.100 3.600 51.900 14.700 ;
        RECT 53.100 3.600 54.900 15.600 ;
        RECT 66.000 10.800 66.900 22.950 ;
        RECT 71.100 21.150 72.900 22.950 ;
        RECT 89.250 21.150 91.050 22.950 ;
        RECT 67.950 18.450 70.050 19.050 ;
        RECT 91.950 18.450 94.050 19.050 ;
        RECT 67.950 17.550 94.050 18.450 ;
        RECT 67.950 16.950 70.050 17.550 ;
        RECT 91.950 16.950 94.050 17.550 ;
        RECT 95.700 15.600 96.600 22.950 ;
        RECT 86.100 14.700 93.900 15.600 ;
        RECT 66.000 9.900 72.600 10.800 ;
        RECT 66.000 9.600 66.900 9.900 ;
        RECT 65.100 3.600 66.900 9.600 ;
        RECT 71.100 9.600 72.600 9.900 ;
        RECT 68.100 3.000 69.900 9.000 ;
        RECT 71.100 3.600 72.900 9.600 ;
        RECT 74.100 3.000 75.900 9.600 ;
        RECT 86.100 3.600 87.900 14.700 ;
        RECT 89.100 3.000 90.900 13.800 ;
        RECT 92.100 3.600 93.900 14.700 ;
        RECT 95.100 3.600 96.900 15.600 ;
        RECT 100.950 15.450 103.050 16.050 ;
        RECT 106.950 15.450 109.050 16.050 ;
        RECT 100.950 14.550 109.050 15.450 ;
        RECT 100.950 13.950 103.050 14.550 ;
        RECT 106.950 13.950 109.050 14.550 ;
        RECT 110.100 15.600 111.300 22.950 ;
        RECT 116.100 21.150 117.900 22.950 ;
        RECT 128.400 15.600 129.300 22.950 ;
        RECT 133.950 21.150 135.750 22.950 ;
        RECT 110.100 14.100 112.500 15.600 ;
        RECT 108.000 11.100 109.800 12.900 ;
        RECT 107.700 3.000 109.500 9.600 ;
        RECT 110.700 3.600 112.500 14.100 ;
        RECT 115.800 3.000 117.600 15.600 ;
        RECT 128.100 3.600 129.900 15.600 ;
        RECT 131.100 14.700 138.900 15.600 ;
        RECT 131.100 3.600 132.900 14.700 ;
        RECT 134.100 3.000 135.900 13.800 ;
        RECT 137.100 3.600 138.900 14.700 ;
        RECT 150.000 10.800 150.900 22.950 ;
        RECT 155.100 21.150 156.900 22.950 ;
        RECT 164.550 21.450 165.450 25.950 ;
        RECT 173.100 25.050 174.300 35.400 ;
        RECT 187.500 30.000 189.300 38.400 ;
        RECT 186.000 28.800 189.300 30.000 ;
        RECT 194.100 29.400 195.900 39.000 ;
        RECT 206.100 35.400 207.900 39.000 ;
        RECT 209.100 35.400 210.900 38.400 ;
        RECT 212.100 35.400 213.900 39.000 ;
        RECT 196.950 33.450 199.050 34.050 ;
        RECT 205.950 33.450 208.050 34.050 ;
        RECT 196.950 32.550 208.050 33.450 ;
        RECT 196.950 31.950 199.050 32.550 ;
        RECT 205.950 31.950 208.050 32.550 ;
        RECT 186.000 25.050 186.900 28.800 ;
        RECT 188.100 25.050 189.900 26.850 ;
        RECT 194.100 25.050 195.900 26.850 ;
        RECT 209.400 25.050 210.300 35.400 ;
        RECT 224.100 32.400 225.900 38.400 ;
        RECT 227.400 33.300 229.200 39.000 ;
        RECT 231.900 33.000 233.700 38.400 ;
        RECT 236.100 33.300 237.900 39.000 ;
        RECT 224.100 31.500 228.600 32.400 ;
        RECT 226.500 29.100 228.600 31.500 ;
        RECT 231.900 30.900 232.800 33.000 ;
        RECT 239.100 32.400 240.900 38.400 ;
        RECT 239.400 31.500 240.900 32.400 ;
        RECT 254.100 33.300 255.900 38.400 ;
        RECT 257.100 34.200 258.900 39.000 ;
        RECT 260.100 33.300 261.900 38.400 ;
        RECT 254.100 31.950 261.900 33.300 ;
        RECT 263.100 32.400 264.900 38.400 ;
        RECT 275.400 32.400 277.200 39.000 ;
        RECT 229.800 28.800 232.800 30.900 ;
        RECT 236.400 30.000 240.900 31.500 ;
        RECT 263.100 30.300 264.300 32.400 ;
        RECT 280.500 31.200 282.300 38.400 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 224.100 22.950 226.200 25.050 ;
        RECT 228.900 24.900 231.000 27.000 ;
        RECT 229.200 23.100 231.000 24.900 ;
        RECT 161.550 20.550 165.450 21.450 ;
        RECT 170.100 21.150 171.900 22.950 ;
        RECT 151.950 18.450 154.050 19.050 ;
        RECT 161.550 18.450 162.450 20.550 ;
        RECT 151.950 17.550 162.450 18.450 ;
        RECT 151.950 16.950 154.050 17.550 ;
        RECT 150.000 9.900 156.600 10.800 ;
        RECT 150.000 9.600 150.900 9.900 ;
        RECT 149.100 3.600 150.900 9.600 ;
        RECT 155.100 9.600 156.600 9.900 ;
        RECT 173.100 9.600 174.300 22.950 ;
        RECT 186.000 10.800 186.900 22.950 ;
        RECT 191.100 21.150 192.900 22.950 ;
        RECT 206.250 21.150 208.050 22.950 ;
        RECT 209.400 15.600 210.300 22.950 ;
        RECT 212.100 21.150 213.900 22.950 ;
        RECT 224.400 21.150 226.200 22.950 ;
        RECT 231.900 22.050 232.800 28.800 ;
        RECT 233.700 27.900 235.500 29.700 ;
        RECT 236.400 29.400 238.500 30.000 ;
        RECT 260.700 29.400 264.300 30.300 ;
        RECT 278.100 30.300 282.300 31.200 ;
        RECT 234.000 27.000 236.100 27.900 ;
        RECT 234.000 25.800 240.600 27.000 ;
        RECT 238.800 25.200 240.600 25.800 ;
        RECT 234.000 22.800 236.100 24.900 ;
        RECT 238.800 22.950 240.900 25.200 ;
        RECT 257.100 25.050 258.900 26.850 ;
        RECT 260.700 25.050 261.900 29.400 ;
        RECT 263.100 25.050 264.900 26.850 ;
        RECT 275.250 25.050 277.050 26.850 ;
        RECT 278.100 25.050 279.300 30.300 ;
        RECT 293.100 29.400 294.900 39.000 ;
        RECT 299.700 30.000 301.500 38.400 ;
        RECT 316.500 30.000 318.300 38.400 ;
        RECT 299.700 28.800 303.000 30.000 ;
        RECT 281.100 25.050 282.900 26.850 ;
        RECT 293.100 25.050 294.900 26.850 ;
        RECT 299.100 25.050 300.900 26.850 ;
        RECT 302.100 25.050 303.000 28.800 ;
        RECT 315.000 28.800 318.300 30.000 ;
        RECT 323.100 29.400 324.900 39.000 ;
        RECT 335.100 32.400 336.900 38.400 ;
        RECT 335.700 30.300 336.900 32.400 ;
        RECT 338.100 33.300 339.900 38.400 ;
        RECT 341.100 34.200 342.900 39.000 ;
        RECT 344.100 33.300 345.900 38.400 ;
        RECT 346.950 36.450 349.050 37.050 ;
        RECT 352.950 36.450 355.050 37.050 ;
        RECT 346.950 35.550 355.050 36.450 ;
        RECT 346.950 34.950 349.050 35.550 ;
        RECT 352.950 34.950 355.050 35.550 ;
        RECT 356.700 35.400 358.500 39.000 ;
        RECT 359.700 33.600 361.500 38.400 ;
        RECT 338.100 31.950 345.900 33.300 ;
        RECT 356.400 32.400 361.500 33.600 ;
        RECT 364.200 32.400 366.000 39.000 ;
        RECT 335.700 29.400 339.300 30.300 ;
        RECT 315.000 25.050 315.900 28.800 ;
        RECT 330.000 27.450 334.050 28.050 ;
        RECT 317.100 25.050 318.900 26.850 ;
        RECT 323.100 25.050 324.900 26.850 ;
        RECT 329.550 25.950 334.050 27.450 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 313.950 22.950 316.050 25.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 229.800 20.700 232.800 22.050 ;
        RECT 234.300 21.000 236.100 22.800 ;
        RECT 254.100 21.150 255.900 22.950 ;
        RECT 229.800 19.950 231.900 20.700 ;
        RECT 227.100 15.600 229.200 16.500 ;
        RECT 186.000 9.900 192.600 10.800 ;
        RECT 186.000 9.600 186.900 9.900 ;
        RECT 152.100 3.000 153.900 9.000 ;
        RECT 155.100 3.600 156.900 9.600 ;
        RECT 158.100 3.000 159.900 9.600 ;
        RECT 170.100 3.000 171.900 9.600 ;
        RECT 173.100 3.600 174.900 9.600 ;
        RECT 185.100 3.600 186.900 9.600 ;
        RECT 191.100 9.600 192.600 9.900 ;
        RECT 188.100 3.000 189.900 9.000 ;
        RECT 191.100 3.600 192.900 9.600 ;
        RECT 194.100 3.000 195.900 9.600 ;
        RECT 206.100 3.000 207.900 15.600 ;
        RECT 209.400 14.400 213.000 15.600 ;
        RECT 211.200 3.600 213.000 14.400 ;
        RECT 224.100 14.400 229.200 15.600 ;
        RECT 230.100 15.600 231.300 19.950 ;
        RECT 232.800 17.700 234.600 19.500 ;
        RECT 232.800 16.800 238.200 17.700 ;
        RECT 236.100 15.900 238.200 16.800 ;
        RECT 230.100 14.700 233.400 15.600 ;
        RECT 236.100 14.700 240.900 15.900 ;
        RECT 260.700 15.600 261.900 22.950 ;
        RECT 224.100 3.600 225.900 14.400 ;
        RECT 227.100 3.000 229.200 13.500 ;
        RECT 231.600 3.600 233.400 14.700 ;
        RECT 236.100 3.000 237.900 13.500 ;
        RECT 239.100 3.600 240.900 14.700 ;
        RECT 254.400 3.000 256.200 15.600 ;
        RECT 259.500 14.100 261.900 15.600 ;
        RECT 259.500 3.600 261.300 14.100 ;
        RECT 262.200 11.100 264.000 12.900 ;
        RECT 278.100 9.600 279.300 22.950 ;
        RECT 296.100 21.150 297.900 22.950 ;
        RECT 302.100 10.800 303.000 22.950 ;
        RECT 296.400 9.900 303.000 10.800 ;
        RECT 296.400 9.600 297.900 9.900 ;
        RECT 262.500 3.000 264.300 9.600 ;
        RECT 275.100 3.000 276.900 9.600 ;
        RECT 278.100 3.600 279.900 9.600 ;
        RECT 281.100 3.000 282.900 9.600 ;
        RECT 293.100 3.000 294.900 9.600 ;
        RECT 296.100 3.600 297.900 9.600 ;
        RECT 302.100 9.600 303.000 9.900 ;
        RECT 315.000 10.800 315.900 22.950 ;
        RECT 320.100 21.150 321.900 22.950 ;
        RECT 329.550 21.450 330.450 25.950 ;
        RECT 335.100 25.050 336.900 26.850 ;
        RECT 338.100 25.050 339.300 29.400 ;
        RECT 341.100 25.050 342.900 26.850 ;
        RECT 356.400 25.050 357.300 32.400 ;
        RECT 379.500 30.000 381.300 38.400 ;
        RECT 378.000 28.800 381.300 30.000 ;
        RECT 386.100 29.400 387.900 39.000 ;
        RECT 399.000 32.400 400.800 39.000 ;
        RECT 403.500 33.600 405.300 38.400 ;
        RECT 406.500 35.400 408.300 39.000 ;
        RECT 419.100 35.400 420.900 38.400 ;
        RECT 422.100 35.400 423.900 39.000 ;
        RECT 403.500 32.400 408.600 33.600 ;
        RECT 358.950 25.050 360.750 26.850 ;
        RECT 365.100 25.050 366.900 26.850 ;
        RECT 378.000 25.050 378.900 28.800 ;
        RECT 380.100 25.050 381.900 26.850 ;
        RECT 386.100 25.050 387.900 26.850 ;
        RECT 398.100 25.050 399.900 26.850 ;
        RECT 404.250 25.050 406.050 26.850 ;
        RECT 407.700 25.050 408.600 32.400 ;
        RECT 409.950 27.450 414.000 28.050 ;
        RECT 409.950 27.000 414.450 27.450 ;
        RECT 409.950 25.950 415.050 27.000 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 376.950 22.950 379.050 25.050 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 382.950 22.950 385.050 25.050 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 326.550 20.550 330.450 21.450 ;
        RECT 316.950 18.450 319.050 19.050 ;
        RECT 326.550 18.450 327.450 20.550 ;
        RECT 316.950 17.550 327.450 18.450 ;
        RECT 316.950 16.950 319.050 17.550 ;
        RECT 338.100 15.600 339.300 22.950 ;
        RECT 344.100 21.150 345.900 22.950 ;
        RECT 356.400 15.600 357.300 22.950 ;
        RECT 361.950 21.150 363.750 22.950 ;
        RECT 338.100 14.100 340.500 15.600 ;
        RECT 336.000 11.100 337.800 12.900 ;
        RECT 315.000 9.900 321.600 10.800 ;
        RECT 315.000 9.600 315.900 9.900 ;
        RECT 299.100 3.000 300.900 9.000 ;
        RECT 302.100 3.600 303.900 9.600 ;
        RECT 314.100 3.600 315.900 9.600 ;
        RECT 320.100 9.600 321.600 9.900 ;
        RECT 317.100 3.000 318.900 9.000 ;
        RECT 320.100 3.600 321.900 9.600 ;
        RECT 323.100 3.000 324.900 9.600 ;
        RECT 335.700 3.000 337.500 9.600 ;
        RECT 338.700 3.600 340.500 14.100 ;
        RECT 343.800 3.000 345.600 15.600 ;
        RECT 356.100 3.600 357.900 15.600 ;
        RECT 359.100 14.700 366.900 15.600 ;
        RECT 359.100 3.600 360.900 14.700 ;
        RECT 362.100 3.000 363.900 13.800 ;
        RECT 365.100 3.600 366.900 14.700 ;
        RECT 378.000 10.800 378.900 22.950 ;
        RECT 383.100 21.150 384.900 22.950 ;
        RECT 401.250 21.150 403.050 22.950 ;
        RECT 379.950 18.450 382.050 19.050 ;
        RECT 391.950 18.450 394.050 19.050 ;
        RECT 379.950 17.550 394.050 18.450 ;
        RECT 379.950 16.950 382.050 17.550 ;
        RECT 391.950 16.950 394.050 17.550 ;
        RECT 379.950 15.450 382.050 15.900 ;
        RECT 391.950 15.450 394.050 15.900 ;
        RECT 407.700 15.600 408.600 22.950 ;
        RECT 412.950 22.800 415.050 25.950 ;
        RECT 419.700 25.050 420.900 35.400 ;
        RECT 434.100 33.300 435.900 38.400 ;
        RECT 437.100 34.200 438.900 39.000 ;
        RECT 440.100 33.300 441.900 38.400 ;
        RECT 434.100 31.950 441.900 33.300 ;
        RECT 443.100 32.400 444.900 38.400 ;
        RECT 443.100 30.300 444.300 32.400 ;
        RECT 440.700 29.400 444.300 30.300 ;
        RECT 455.100 29.400 456.900 39.000 ;
        RECT 461.700 30.000 463.500 38.400 ;
        RECT 476.700 31.200 478.500 38.400 ;
        RECT 481.800 32.400 483.600 39.000 ;
        RECT 495.600 34.200 497.400 38.400 ;
        RECT 494.700 32.400 497.400 34.200 ;
        RECT 498.600 32.400 500.400 39.000 ;
        RECT 476.700 30.300 480.900 31.200 ;
        RECT 437.100 25.050 438.900 26.850 ;
        RECT 440.700 25.050 441.900 29.400 ;
        RECT 461.700 28.800 465.000 30.000 ;
        RECT 443.100 25.050 444.900 26.850 ;
        RECT 455.100 25.050 456.900 26.850 ;
        RECT 461.100 25.050 462.900 26.850 ;
        RECT 464.100 25.050 465.000 28.800 ;
        RECT 476.100 25.050 477.900 26.850 ;
        RECT 479.700 25.050 480.900 30.300 ;
        RECT 481.950 25.050 483.750 26.850 ;
        RECT 494.700 25.050 495.600 32.400 ;
        RECT 496.500 30.600 498.300 31.500 ;
        RECT 503.100 30.600 504.900 38.400 ;
        RECT 515.400 32.400 517.200 39.000 ;
        RECT 520.500 31.200 522.300 38.400 ;
        RECT 496.500 29.700 504.900 30.600 ;
        RECT 518.100 30.300 522.300 31.200 ;
        RECT 418.950 22.950 421.050 25.050 ;
        RECT 421.950 22.950 424.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 475.950 22.950 478.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 494.100 22.950 496.200 25.050 ;
        RECT 497.400 22.950 499.500 25.050 ;
        RECT 379.950 14.550 394.050 15.450 ;
        RECT 379.950 13.800 382.050 14.550 ;
        RECT 391.950 13.800 394.050 14.550 ;
        RECT 398.100 14.700 405.900 15.600 ;
        RECT 378.000 9.900 384.600 10.800 ;
        RECT 378.000 9.600 378.900 9.900 ;
        RECT 377.100 3.600 378.900 9.600 ;
        RECT 383.100 9.600 384.600 9.900 ;
        RECT 380.100 3.000 381.900 9.000 ;
        RECT 383.100 3.600 384.900 9.600 ;
        RECT 386.100 3.000 387.900 9.600 ;
        RECT 398.100 3.600 399.900 14.700 ;
        RECT 401.100 3.000 402.900 13.800 ;
        RECT 404.100 3.600 405.900 14.700 ;
        RECT 407.100 3.600 408.900 15.600 ;
        RECT 419.700 9.600 420.900 22.950 ;
        RECT 422.100 21.150 423.900 22.950 ;
        RECT 434.100 21.150 435.900 22.950 ;
        RECT 440.700 15.600 441.900 22.950 ;
        RECT 458.100 21.150 459.900 22.950 ;
        RECT 419.100 3.600 420.900 9.600 ;
        RECT 422.100 3.000 423.900 9.600 ;
        RECT 434.400 3.000 436.200 15.600 ;
        RECT 439.500 14.100 441.900 15.600 ;
        RECT 439.500 3.600 441.300 14.100 ;
        RECT 442.200 11.100 444.000 12.900 ;
        RECT 464.100 10.800 465.000 22.950 ;
        RECT 458.400 9.900 465.000 10.800 ;
        RECT 458.400 9.600 459.900 9.900 ;
        RECT 442.500 3.000 444.300 9.600 ;
        RECT 455.100 3.000 456.900 9.600 ;
        RECT 458.100 3.600 459.900 9.600 ;
        RECT 464.100 9.600 465.000 9.900 ;
        RECT 479.700 9.600 480.900 22.950 ;
        RECT 494.700 15.600 495.600 22.950 ;
        RECT 498.000 21.150 499.800 22.950 ;
        RECT 461.100 3.000 462.900 9.000 ;
        RECT 464.100 3.600 465.900 9.600 ;
        RECT 476.100 3.000 477.900 9.600 ;
        RECT 479.100 3.600 480.900 9.600 ;
        RECT 482.100 3.000 483.900 9.600 ;
        RECT 494.100 3.600 495.900 15.600 ;
        RECT 497.100 3.000 498.900 15.000 ;
        RECT 501.000 9.600 501.900 29.700 ;
        RECT 502.950 25.050 504.750 26.850 ;
        RECT 515.250 25.050 517.050 26.850 ;
        RECT 518.100 25.050 519.300 30.300 ;
        RECT 535.500 30.000 537.300 38.400 ;
        RECT 534.000 28.800 537.300 30.000 ;
        RECT 542.100 29.400 543.900 39.000 ;
        RECT 557.100 32.400 558.900 38.400 ;
        RECT 557.700 30.300 558.900 32.400 ;
        RECT 560.100 33.300 561.900 38.400 ;
        RECT 563.100 34.200 564.900 39.000 ;
        RECT 566.100 33.300 567.900 38.400 ;
        RECT 578.700 35.400 580.500 39.000 ;
        RECT 581.700 33.600 583.500 38.400 ;
        RECT 560.100 31.950 567.900 33.300 ;
        RECT 578.400 32.400 583.500 33.600 ;
        RECT 586.200 32.400 588.000 39.000 ;
        RECT 599.700 35.400 601.500 39.000 ;
        RECT 602.700 33.600 604.500 38.400 ;
        RECT 599.400 32.400 604.500 33.600 ;
        RECT 607.200 32.400 609.000 39.000 ;
        RECT 557.700 29.400 561.300 30.300 ;
        RECT 521.100 25.050 522.900 26.850 ;
        RECT 534.000 25.050 534.900 28.800 ;
        RECT 536.100 25.050 537.900 26.850 ;
        RECT 542.100 25.050 543.900 26.850 ;
        RECT 557.100 25.050 558.900 26.850 ;
        RECT 560.100 25.050 561.300 29.400 ;
        RECT 573.000 27.450 577.050 28.050 ;
        RECT 563.100 25.050 564.900 26.850 ;
        RECT 572.550 25.950 577.050 27.450 ;
        RECT 502.800 22.950 504.900 25.050 ;
        RECT 514.950 22.950 517.050 25.050 ;
        RECT 517.950 22.950 520.050 25.050 ;
        RECT 520.950 22.950 523.050 25.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 518.100 9.600 519.300 22.950 ;
        RECT 520.950 18.450 523.050 19.050 ;
        RECT 526.950 18.450 529.050 19.050 ;
        RECT 520.950 17.550 529.050 18.450 ;
        RECT 520.950 16.950 523.050 17.550 ;
        RECT 526.950 16.950 529.050 17.550 ;
        RECT 534.000 10.800 534.900 22.950 ;
        RECT 539.100 21.150 540.900 22.950 ;
        RECT 560.100 15.600 561.300 22.950 ;
        RECT 566.100 21.150 567.900 22.950 ;
        RECT 572.550 21.450 573.450 25.950 ;
        RECT 578.400 25.050 579.300 32.400 ;
        RECT 580.950 25.050 582.750 26.850 ;
        RECT 587.100 25.050 588.900 26.850 ;
        RECT 599.400 25.050 600.300 32.400 ;
        RECT 622.500 30.000 624.300 38.400 ;
        RECT 621.000 28.800 624.300 30.000 ;
        RECT 629.100 29.400 630.900 39.000 ;
        RECT 643.500 30.000 645.300 38.400 ;
        RECT 642.000 28.800 645.300 30.000 ;
        RECT 650.100 29.400 651.900 39.000 ;
        RECT 662.100 32.400 663.900 38.400 ;
        RECT 662.700 30.300 663.900 32.400 ;
        RECT 665.100 33.300 666.900 38.400 ;
        RECT 668.100 34.200 669.900 39.000 ;
        RECT 671.100 33.300 672.900 38.400 ;
        RECT 665.100 31.950 672.900 33.300 ;
        RECT 683.100 32.400 684.900 38.400 ;
        RECT 683.700 30.300 684.900 32.400 ;
        RECT 686.100 33.300 687.900 38.400 ;
        RECT 689.100 34.200 690.900 39.000 ;
        RECT 692.100 33.300 693.900 38.400 ;
        RECT 704.700 35.400 706.500 39.000 ;
        RECT 707.700 33.600 709.500 38.400 ;
        RECT 686.100 31.950 693.900 33.300 ;
        RECT 704.400 32.400 709.500 33.600 ;
        RECT 712.200 32.400 714.000 39.000 ;
        RECT 662.700 29.400 666.300 30.300 ;
        RECT 683.700 29.400 687.300 30.300 ;
        RECT 615.000 27.450 619.050 28.050 ;
        RECT 601.950 25.050 603.750 26.850 ;
        RECT 608.100 25.050 609.900 26.850 ;
        RECT 614.550 25.950 619.050 27.450 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 572.550 21.000 576.450 21.450 ;
        RECT 572.550 20.550 577.050 21.000 ;
        RECT 574.950 16.950 577.050 20.550 ;
        RECT 578.400 15.600 579.300 22.950 ;
        RECT 583.950 21.150 585.750 22.950 ;
        RECT 599.400 15.600 600.300 22.950 ;
        RECT 604.950 21.150 606.750 22.950 ;
        RECT 614.550 22.050 615.450 25.950 ;
        RECT 621.000 25.050 621.900 28.800 ;
        RECT 623.100 25.050 624.900 26.850 ;
        RECT 629.100 25.050 630.900 26.850 ;
        RECT 642.000 25.050 642.900 28.800 ;
        RECT 644.100 25.050 645.900 26.850 ;
        RECT 650.100 25.050 651.900 26.850 ;
        RECT 662.100 25.050 663.900 26.850 ;
        RECT 665.100 25.050 666.300 29.400 ;
        RECT 668.100 25.050 669.900 26.850 ;
        RECT 683.100 25.050 684.900 26.850 ;
        RECT 686.100 25.050 687.300 29.400 ;
        RECT 699.000 27.450 703.050 28.050 ;
        RECT 689.100 25.050 690.900 26.850 ;
        RECT 698.550 25.950 703.050 27.450 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 640.950 22.950 643.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 646.950 22.950 649.050 25.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 667.950 22.950 670.050 25.050 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 688.950 22.950 691.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 610.950 20.550 615.450 22.050 ;
        RECT 610.950 19.950 615.000 20.550 ;
        RECT 560.100 14.100 562.500 15.600 ;
        RECT 558.000 11.100 559.800 12.900 ;
        RECT 534.000 9.900 540.600 10.800 ;
        RECT 534.000 9.600 534.900 9.900 ;
        RECT 500.100 3.600 501.900 9.600 ;
        RECT 503.100 3.000 504.900 9.600 ;
        RECT 515.100 3.000 516.900 9.600 ;
        RECT 518.100 3.600 519.900 9.600 ;
        RECT 521.100 3.000 522.900 9.600 ;
        RECT 533.100 3.600 534.900 9.600 ;
        RECT 539.100 9.600 540.600 9.900 ;
        RECT 536.100 3.000 537.900 9.000 ;
        RECT 539.100 3.600 540.900 9.600 ;
        RECT 542.100 3.000 543.900 9.600 ;
        RECT 557.700 3.000 559.500 9.600 ;
        RECT 560.700 3.600 562.500 14.100 ;
        RECT 565.800 3.000 567.600 15.600 ;
        RECT 578.100 3.600 579.900 15.600 ;
        RECT 581.100 14.700 588.900 15.600 ;
        RECT 581.100 3.600 582.900 14.700 ;
        RECT 584.100 3.000 585.900 13.800 ;
        RECT 587.100 3.600 588.900 14.700 ;
        RECT 599.100 3.600 600.900 15.600 ;
        RECT 602.100 14.700 609.900 15.600 ;
        RECT 602.100 3.600 603.900 14.700 ;
        RECT 605.100 3.000 606.900 13.800 ;
        RECT 608.100 3.600 609.900 14.700 ;
        RECT 621.000 10.800 621.900 22.950 ;
        RECT 626.100 21.150 627.900 22.950 ;
        RECT 622.950 18.450 625.050 19.050 ;
        RECT 634.950 18.450 637.050 19.050 ;
        RECT 622.950 17.550 637.050 18.450 ;
        RECT 622.950 16.950 625.050 17.550 ;
        RECT 634.950 16.950 637.050 17.550 ;
        RECT 642.000 10.800 642.900 22.950 ;
        RECT 647.100 21.150 648.900 22.950 ;
        RECT 665.100 15.600 666.300 22.950 ;
        RECT 671.100 21.150 672.900 22.950 ;
        RECT 686.100 15.600 687.300 22.950 ;
        RECT 692.100 21.150 693.900 22.950 ;
        RECT 698.550 21.450 699.450 25.950 ;
        RECT 704.400 25.050 705.300 32.400 ;
        RECT 725.100 30.600 726.900 38.400 ;
        RECT 729.600 32.400 731.400 39.000 ;
        RECT 732.600 34.200 734.400 38.400 ;
        RECT 732.600 32.400 735.300 34.200 ;
        RECT 731.700 30.600 733.500 31.500 ;
        RECT 725.100 29.700 733.500 30.600 ;
        RECT 706.950 25.050 708.750 26.850 ;
        RECT 713.100 25.050 714.900 26.850 ;
        RECT 725.250 25.050 727.050 26.850 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 725.100 22.950 727.200 25.050 ;
        RECT 695.550 20.550 699.450 21.450 ;
        RECT 688.950 18.450 691.050 19.050 ;
        RECT 695.550 18.450 696.450 20.550 ;
        RECT 688.950 17.550 696.450 18.450 ;
        RECT 688.950 16.950 691.050 17.550 ;
        RECT 704.400 15.600 705.300 22.950 ;
        RECT 709.950 21.150 711.750 22.950 ;
        RECT 665.100 14.100 667.500 15.600 ;
        RECT 663.000 11.100 664.800 12.900 ;
        RECT 621.000 9.900 627.600 10.800 ;
        RECT 621.000 9.600 621.900 9.900 ;
        RECT 620.100 3.600 621.900 9.600 ;
        RECT 626.100 9.600 627.600 9.900 ;
        RECT 642.000 9.900 648.600 10.800 ;
        RECT 642.000 9.600 642.900 9.900 ;
        RECT 623.100 3.000 624.900 9.000 ;
        RECT 626.100 3.600 627.900 9.600 ;
        RECT 629.100 3.000 630.900 9.600 ;
        RECT 641.100 3.600 642.900 9.600 ;
        RECT 647.100 9.600 648.600 9.900 ;
        RECT 644.100 3.000 645.900 9.000 ;
        RECT 647.100 3.600 648.900 9.600 ;
        RECT 650.100 3.000 651.900 9.600 ;
        RECT 662.700 3.000 664.500 9.600 ;
        RECT 665.700 3.600 667.500 14.100 ;
        RECT 670.800 3.000 672.600 15.600 ;
        RECT 686.100 14.100 688.500 15.600 ;
        RECT 684.000 11.100 685.800 12.900 ;
        RECT 683.700 3.000 685.500 9.600 ;
        RECT 686.700 3.600 688.500 14.100 ;
        RECT 691.800 3.000 693.600 15.600 ;
        RECT 704.100 3.600 705.900 15.600 ;
        RECT 707.100 14.700 714.900 15.600 ;
        RECT 707.100 3.600 708.900 14.700 ;
        RECT 710.100 3.000 711.900 13.800 ;
        RECT 713.100 3.600 714.900 14.700 ;
        RECT 728.100 9.600 729.000 29.700 ;
        RECT 734.400 25.050 735.300 32.400 ;
        RECT 748.500 30.000 750.300 38.400 ;
        RECT 747.000 28.800 750.300 30.000 ;
        RECT 755.100 29.400 756.900 39.000 ;
        RECT 768.000 32.400 769.800 39.000 ;
        RECT 772.500 33.600 774.300 38.400 ;
        RECT 775.500 35.400 777.300 39.000 ;
        RECT 788.100 35.400 789.900 38.400 ;
        RECT 791.100 35.400 792.900 39.000 ;
        RECT 803.100 35.400 804.900 39.000 ;
        RECT 806.100 35.400 807.900 38.400 ;
        RECT 809.100 35.400 810.900 39.000 ;
        RECT 772.500 32.400 777.600 33.600 ;
        RECT 757.950 30.450 760.050 31.050 ;
        RECT 769.950 30.450 772.050 31.050 ;
        RECT 757.950 29.550 772.050 30.450 ;
        RECT 757.950 28.950 760.050 29.550 ;
        RECT 769.950 28.950 772.050 29.550 ;
        RECT 747.000 25.050 747.900 28.800 ;
        RECT 749.100 25.050 750.900 26.850 ;
        RECT 755.100 25.050 756.900 26.850 ;
        RECT 767.100 25.050 768.900 26.850 ;
        RECT 773.250 25.050 775.050 26.850 ;
        RECT 776.700 25.050 777.600 32.400 ;
        RECT 788.700 25.050 789.900 35.400 ;
        RECT 796.950 33.450 799.050 34.050 ;
        RECT 802.950 33.450 805.050 34.050 ;
        RECT 796.950 32.550 805.050 33.450 ;
        RECT 796.950 31.950 799.050 32.550 ;
        RECT 802.950 31.950 805.050 32.550 ;
        RECT 806.700 25.050 807.600 35.400 ;
        RECT 823.500 30.000 825.300 38.400 ;
        RECT 822.000 28.800 825.300 30.000 ;
        RECT 830.100 29.400 831.900 39.000 ;
        RECT 844.500 30.000 846.300 38.400 ;
        RECT 843.000 28.800 846.300 30.000 ;
        RECT 851.100 29.400 852.900 39.000 ;
        RECT 863.100 35.400 864.900 38.400 ;
        RECT 866.100 35.400 867.900 39.000 ;
        RECT 822.000 25.050 822.900 28.800 ;
        RECT 824.100 25.050 825.900 26.850 ;
        RECT 830.100 25.050 831.900 26.850 ;
        RECT 843.000 25.050 843.900 28.800 ;
        RECT 845.100 25.050 846.900 26.850 ;
        RECT 851.100 25.050 852.900 26.850 ;
        RECT 863.700 25.050 864.900 35.400 ;
        RECT 730.500 22.950 732.600 25.050 ;
        RECT 733.800 22.950 735.900 25.050 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 787.950 22.950 790.050 25.050 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 808.950 22.950 811.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 829.950 22.950 832.050 25.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 850.950 22.950 853.050 25.050 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 730.200 21.150 732.000 22.950 ;
        RECT 734.400 15.600 735.300 22.950 ;
        RECT 725.100 3.000 726.900 9.600 ;
        RECT 728.100 3.600 729.900 9.600 ;
        RECT 731.100 3.000 732.900 15.000 ;
        RECT 734.100 3.600 735.900 15.600 ;
        RECT 747.000 10.800 747.900 22.950 ;
        RECT 752.100 21.150 753.900 22.950 ;
        RECT 770.250 21.150 772.050 22.950 ;
        RECT 748.950 18.450 751.050 18.750 ;
        RECT 766.950 18.450 769.050 19.050 ;
        RECT 748.950 17.550 769.050 18.450 ;
        RECT 748.950 16.650 751.050 17.550 ;
        RECT 766.950 16.950 769.050 17.550 ;
        RECT 776.700 15.600 777.600 22.950 ;
        RECT 767.100 14.700 774.900 15.600 ;
        RECT 747.000 9.900 753.600 10.800 ;
        RECT 747.000 9.600 747.900 9.900 ;
        RECT 746.100 3.600 747.900 9.600 ;
        RECT 752.100 9.600 753.600 9.900 ;
        RECT 749.100 3.000 750.900 9.000 ;
        RECT 752.100 3.600 753.900 9.600 ;
        RECT 755.100 3.000 756.900 9.600 ;
        RECT 767.100 3.600 768.900 14.700 ;
        RECT 770.100 3.000 771.900 13.800 ;
        RECT 773.100 3.600 774.900 14.700 ;
        RECT 776.100 3.600 777.900 15.600 ;
        RECT 788.700 9.600 789.900 22.950 ;
        RECT 791.100 21.150 792.900 22.950 ;
        RECT 803.100 21.150 804.900 22.950 ;
        RECT 806.700 15.600 807.600 22.950 ;
        RECT 808.950 21.150 810.750 22.950 ;
        RECT 804.000 14.400 807.600 15.600 ;
        RECT 788.100 3.600 789.900 9.600 ;
        RECT 791.100 3.000 792.900 9.600 ;
        RECT 804.000 3.600 805.800 14.400 ;
        RECT 809.100 3.000 810.900 15.600 ;
        RECT 822.000 10.800 822.900 22.950 ;
        RECT 827.100 21.150 828.900 22.950 ;
        RECT 823.950 18.450 826.050 19.050 ;
        RECT 835.950 18.450 838.050 19.050 ;
        RECT 823.950 17.550 838.050 18.450 ;
        RECT 823.950 16.950 826.050 17.550 ;
        RECT 835.950 16.950 838.050 17.550 ;
        RECT 843.000 10.800 843.900 22.950 ;
        RECT 848.100 21.150 849.900 22.950 ;
        RECT 822.000 9.900 828.600 10.800 ;
        RECT 822.000 9.600 822.900 9.900 ;
        RECT 821.100 3.600 822.900 9.600 ;
        RECT 827.100 9.600 828.600 9.900 ;
        RECT 843.000 9.900 849.600 10.800 ;
        RECT 843.000 9.600 843.900 9.900 ;
        RECT 824.100 3.000 825.900 9.000 ;
        RECT 827.100 3.600 828.900 9.600 ;
        RECT 830.100 3.000 831.900 9.600 ;
        RECT 842.100 3.600 843.900 9.600 ;
        RECT 848.100 9.600 849.600 9.900 ;
        RECT 863.700 9.600 864.900 22.950 ;
        RECT 866.100 21.150 867.900 22.950 ;
        RECT 845.100 3.000 846.900 9.000 ;
        RECT 848.100 3.600 849.900 9.600 ;
        RECT 851.100 3.000 852.900 9.600 ;
        RECT 863.100 3.600 864.900 9.600 ;
        RECT 866.100 3.000 867.900 9.600 ;
      LAYER metal2 ;
        RECT 454.950 817.950 457.050 820.050 ;
        RECT 484.950 817.950 487.050 820.050 ;
        RECT 8.850 813.300 10.950 815.400 ;
        RECT 26.550 813.300 28.650 815.400 ;
        RECT 61.350 813.300 63.450 815.400 ;
        RECT 79.050 813.300 81.150 815.400 ;
        RECT 173.850 813.300 175.950 815.400 ;
        RECT 191.550 813.300 193.650 815.400 ;
        RECT 4.950 802.950 7.050 805.050 ;
        RECT 5.400 800.400 6.600 802.650 ;
        RECT 5.400 787.050 6.450 800.400 ;
        RECT 9.150 794.700 10.350 813.300 ;
        RECT 14.100 802.950 16.200 805.050 ;
        RECT 14.400 801.450 15.600 802.650 ;
        RECT 14.400 800.400 18.450 801.450 ;
        RECT 9.150 793.500 13.350 794.700 ;
        RECT 11.250 792.600 13.350 793.500 ;
        RECT 4.950 784.950 7.050 787.050 ;
        RECT 17.400 778.050 18.450 800.400 ;
        RECT 26.550 800.400 27.750 813.300 ;
        RECT 31.950 806.100 34.050 808.200 ;
        RECT 49.950 806.100 52.050 808.200 ;
        RECT 55.950 806.100 58.050 808.200 ;
        RECT 32.400 805.350 33.600 806.100 ;
        RECT 50.400 805.350 51.600 806.100 ;
        RECT 56.400 805.350 57.600 806.100 ;
        RECT 31.950 802.950 34.050 805.050 ;
        RECT 40.950 802.950 43.050 805.050 ;
        RECT 46.950 802.950 49.050 805.050 ;
        RECT 49.950 802.950 52.050 805.050 ;
        RECT 55.950 802.950 58.050 805.050 ;
        RECT 26.550 798.300 28.650 800.400 ;
        RECT 26.550 791.700 27.750 798.300 ;
        RECT 26.550 789.600 28.650 791.700 ;
        RECT 10.950 775.950 13.050 778.050 ;
        RECT 16.950 775.950 19.050 778.050 ;
        RECT 7.950 761.100 10.050 763.200 ;
        RECT 11.400 763.050 12.450 775.950 ;
        RECT 41.400 772.050 42.450 802.950 ;
        RECT 47.400 801.000 48.600 802.650 ;
        RECT 46.950 796.950 49.050 801.000 ;
        RECT 52.950 798.450 55.050 802.050 ;
        RECT 62.250 800.400 63.450 813.300 ;
        RECT 73.800 802.950 75.900 805.050 ;
        RECT 74.400 801.900 75.600 802.650 ;
        RECT 50.400 798.000 55.050 798.450 ;
        RECT 61.350 798.300 63.450 800.400 ;
        RECT 73.950 799.800 76.050 801.900 ;
        RECT 50.400 797.400 54.450 798.000 ;
        RECT 40.950 769.950 43.050 772.050 ;
        RECT 8.400 730.050 9.450 761.100 ;
        RECT 10.950 760.950 13.050 763.050 ;
        RECT 16.950 761.100 19.050 763.200 ;
        RECT 22.950 761.100 25.050 763.200 ;
        RECT 28.950 761.100 31.050 763.200 ;
        RECT 34.950 761.100 37.050 763.200 ;
        RECT 41.400 762.600 42.450 769.950 ;
        RECT 17.400 760.350 18.600 761.100 ;
        RECT 23.400 760.350 24.600 761.100 ;
        RECT 13.950 757.950 16.050 760.050 ;
        RECT 16.950 757.950 19.050 760.050 ;
        RECT 19.950 757.950 22.050 760.050 ;
        RECT 22.950 757.950 25.050 760.050 ;
        RECT 10.950 751.950 13.050 757.050 ;
        RECT 14.400 755.400 15.600 757.650 ;
        RECT 20.400 756.900 21.600 757.650 ;
        RECT 14.400 742.050 15.450 755.400 ;
        RECT 19.950 754.800 22.050 756.900 ;
        RECT 29.400 751.050 30.450 761.100 ;
        RECT 35.400 760.350 36.600 761.100 ;
        RECT 41.400 760.350 42.600 762.600 ;
        RECT 46.950 760.950 49.050 763.050 ;
        RECT 34.950 757.950 37.050 760.050 ;
        RECT 37.950 757.950 40.050 760.050 ;
        RECT 40.950 757.950 43.050 760.050 ;
        RECT 31.950 754.950 34.050 757.050 ;
        RECT 38.400 755.400 39.600 757.650 ;
        RECT 28.950 748.950 31.050 751.050 ;
        RECT 32.400 742.050 33.450 754.950 ;
        RECT 38.400 751.050 39.450 755.400 ;
        RECT 37.950 748.950 40.050 751.050 ;
        RECT 13.950 739.950 16.050 742.050 ;
        RECT 31.950 739.950 34.050 742.050 ;
        RECT 47.400 736.050 48.450 760.950 ;
        RECT 50.400 757.050 51.450 797.400 ;
        RECT 62.250 791.700 63.450 798.300 ;
        RECT 79.650 794.700 80.850 813.300 ;
        RECT 91.950 806.100 94.050 808.200 ;
        RECT 97.950 807.000 100.050 811.050 ;
        RECT 112.950 808.950 115.050 811.050 ;
        RECT 82.950 802.950 85.050 805.050 ;
        RECT 76.650 793.500 80.850 794.700 ;
        RECT 83.400 800.400 84.600 802.650 ;
        RECT 92.400 802.050 93.450 806.100 ;
        RECT 98.400 805.350 99.600 807.000 ;
        RECT 103.950 806.100 106.050 808.200 ;
        RECT 104.400 805.350 105.600 806.100 ;
        RECT 97.950 802.950 100.050 805.050 ;
        RECT 100.950 802.950 103.050 805.050 ;
        RECT 103.950 802.950 106.050 805.050 ;
        RECT 106.950 802.950 109.050 805.050 ;
        RECT 76.650 792.600 78.750 793.500 ;
        RECT 61.350 789.600 63.450 791.700 ;
        RECT 83.400 787.050 84.450 800.400 ;
        RECT 91.950 799.950 94.050 802.050 ;
        RECT 101.400 800.400 102.600 802.650 ;
        RECT 107.400 801.900 108.600 802.650 ;
        RECT 101.400 799.050 102.450 800.400 ;
        RECT 106.950 799.800 109.050 801.900 ;
        RECT 100.950 796.950 103.050 799.050 ;
        RECT 101.400 793.050 102.450 796.950 ;
        RECT 113.400 793.050 114.450 808.950 ;
        RECT 121.950 806.100 124.050 808.200 ;
        RECT 122.400 805.350 123.600 806.100 ;
        RECT 118.950 802.950 121.050 805.050 ;
        RECT 121.950 802.950 124.050 805.050 ;
        RECT 124.950 802.950 127.050 805.050 ;
        RECT 143.100 802.950 145.200 805.050 ;
        RECT 161.100 802.950 163.200 805.050 ;
        RECT 169.950 802.950 172.050 805.050 ;
        RECT 119.400 800.400 120.600 802.650 ;
        RECT 125.400 800.400 126.600 802.650 ;
        RECT 143.400 801.000 144.600 802.650 ;
        RECT 170.400 801.000 171.600 802.650 ;
        RECT 119.400 793.050 120.450 800.400 ;
        RECT 100.950 790.950 103.050 793.050 ;
        RECT 106.950 790.950 109.050 793.050 ;
        RECT 112.950 790.950 115.050 793.050 ;
        RECT 118.950 790.950 121.050 793.050 ;
        RECT 82.950 784.950 85.050 787.050 ;
        RECT 88.950 784.950 91.050 787.050 ;
        RECT 103.950 784.950 106.050 787.050 ;
        RECT 58.950 761.100 61.050 763.200 ;
        RECT 67.950 761.100 70.050 763.200 ;
        RECT 76.950 761.100 79.050 763.200 ;
        RECT 82.950 762.000 85.050 766.050 ;
        RECT 89.400 762.600 90.450 784.950 ;
        RECT 95.250 769.500 97.350 770.400 ;
        RECT 93.150 768.300 97.350 769.500 ;
        RECT 59.400 760.350 60.600 761.100 ;
        RECT 55.950 757.950 58.050 760.050 ;
        RECT 58.950 757.950 61.050 760.050 ;
        RECT 61.950 757.950 64.050 760.050 ;
        RECT 49.950 754.950 52.050 757.050 ;
        RECT 56.400 756.900 57.600 757.650 ;
        RECT 55.950 754.800 58.050 756.900 ;
        RECT 62.400 755.400 63.600 757.650 ;
        RECT 68.400 756.450 69.450 761.100 ;
        RECT 77.400 760.350 78.600 761.100 ;
        RECT 83.400 760.350 84.600 762.000 ;
        RECT 89.400 760.350 90.600 762.600 ;
        RECT 73.950 757.950 76.050 760.050 ;
        RECT 76.950 757.950 79.050 760.050 ;
        RECT 79.950 757.950 82.050 760.050 ;
        RECT 82.950 757.950 85.050 760.050 ;
        RECT 88.950 757.950 91.050 760.050 ;
        RECT 68.400 755.400 72.450 756.450 ;
        RECT 62.400 748.050 63.450 755.400 ;
        RECT 61.950 745.950 64.050 748.050 ;
        RECT 34.950 733.950 37.050 736.050 ;
        RECT 40.950 733.950 43.050 736.050 ;
        RECT 46.950 733.950 49.050 736.050 ;
        RECT 7.950 727.950 10.050 730.050 ;
        RECT 13.950 728.100 16.050 730.200 ;
        RECT 14.400 727.350 15.600 728.100 ;
        RECT 22.950 727.950 25.050 730.050 ;
        RECT 28.950 728.100 31.050 730.200 ;
        RECT 35.400 729.600 36.450 733.950 ;
        RECT 10.950 724.950 13.050 727.050 ;
        RECT 13.950 724.950 16.050 727.050 ;
        RECT 16.950 724.950 19.050 727.050 ;
        RECT 7.950 721.950 10.050 724.050 ;
        RECT 11.400 722.400 12.600 724.650 ;
        RECT 17.400 723.000 18.600 724.650 ;
        RECT 8.400 658.050 9.450 721.950 ;
        RECT 11.400 685.050 12.450 722.400 ;
        RECT 16.950 718.950 19.050 723.000 ;
        RECT 23.400 718.050 24.450 727.950 ;
        RECT 29.400 727.350 30.600 728.100 ;
        RECT 35.400 727.350 36.600 729.600 ;
        RECT 28.950 724.950 31.050 727.050 ;
        RECT 31.950 724.950 34.050 727.050 ;
        RECT 34.950 724.950 37.050 727.050 ;
        RECT 32.400 722.400 33.600 724.650 ;
        RECT 41.400 723.900 42.450 733.950 ;
        RECT 46.950 728.100 49.050 730.200 ;
        RECT 52.950 728.100 55.050 730.200 ;
        RECT 47.400 727.350 48.600 728.100 ;
        RECT 53.400 727.350 54.600 728.100 ;
        RECT 61.950 727.950 64.050 730.050 ;
        RECT 71.400 729.600 72.450 755.400 ;
        RECT 74.400 755.400 75.600 757.650 ;
        RECT 80.400 756.900 81.600 757.650 ;
        RECT 74.400 742.050 75.450 755.400 ;
        RECT 79.950 754.800 82.050 756.900 ;
        RECT 93.150 749.700 94.350 768.300 ;
        RECT 97.950 761.100 100.050 763.200 ;
        RECT 98.400 760.350 99.600 761.100 ;
        RECT 98.100 757.950 100.200 760.050 ;
        RECT 104.400 751.050 105.450 784.950 ;
        RECT 92.850 747.600 94.950 749.700 ;
        RECT 103.950 748.950 106.050 751.050 ;
        RECT 97.950 745.950 100.050 748.050 ;
        RECT 73.950 739.950 76.050 742.050 ;
        RECT 46.950 724.950 49.050 727.050 ;
        RECT 49.950 724.950 52.050 727.050 ;
        RECT 52.950 724.950 55.050 727.050 ;
        RECT 55.950 724.950 58.050 727.050 ;
        RECT 50.400 723.900 51.600 724.650 ;
        RECT 32.400 721.050 33.450 722.400 ;
        RECT 40.950 721.800 43.050 723.900 ;
        RECT 49.950 721.800 52.050 723.900 ;
        RECT 56.400 722.400 57.600 724.650 ;
        RECT 62.400 723.900 63.450 727.950 ;
        RECT 71.400 727.350 72.600 729.600 ;
        RECT 85.950 729.000 88.050 733.050 ;
        RECT 86.400 727.350 87.600 729.000 ;
        RECT 91.950 728.100 94.050 730.200 ;
        RECT 92.400 727.350 93.600 728.100 ;
        RECT 67.950 724.950 70.050 727.050 ;
        RECT 70.950 724.950 73.050 727.050 ;
        RECT 73.950 724.950 76.050 727.050 ;
        RECT 85.950 724.950 88.050 727.050 ;
        RECT 88.950 724.950 91.050 727.050 ;
        RECT 91.950 724.950 94.050 727.050 ;
        RECT 68.400 723.900 69.600 724.650 ;
        RECT 28.950 719.400 33.450 721.050 ;
        RECT 28.950 718.950 33.000 719.400 ;
        RECT 22.950 715.950 25.050 718.050 ;
        RECT 56.400 691.050 57.450 722.400 ;
        RECT 61.950 721.800 64.050 723.900 ;
        RECT 67.950 721.800 70.050 723.900 ;
        RECT 74.400 722.400 75.600 724.650 ;
        RECT 89.400 723.900 90.600 724.650 ;
        RECT 74.400 718.050 75.450 722.400 ;
        RECT 88.950 721.800 91.050 723.900 ;
        RECT 73.950 715.950 76.050 718.050 ;
        RECT 98.400 709.050 99.450 745.950 ;
        RECT 107.400 745.050 108.450 790.950 ;
        RECT 110.550 771.300 112.650 773.400 ;
        RECT 110.550 764.700 111.750 771.300 ;
        RECT 110.550 762.600 112.650 764.700 ;
        RECT 121.950 763.950 124.050 766.050 ;
        RECT 110.550 749.700 111.750 762.600 ;
        RECT 115.950 757.950 118.050 760.050 ;
        RECT 116.400 756.900 117.600 757.650 ;
        RECT 115.950 754.800 118.050 756.900 ;
        RECT 122.400 754.050 123.450 763.950 ;
        RECT 121.950 751.950 124.050 754.050 ;
        RECT 110.550 747.600 112.650 749.700 ;
        RECT 118.950 748.950 121.050 751.050 ;
        RECT 106.950 742.950 109.050 745.050 ;
        RECT 112.950 742.950 115.050 745.050 ;
        RECT 106.950 736.950 109.050 739.050 ;
        RECT 107.400 729.600 108.450 736.950 ;
        RECT 113.400 733.050 114.450 742.950 ;
        RECT 107.400 727.350 108.600 729.600 ;
        RECT 112.950 729.000 115.050 733.050 ;
        RECT 113.400 727.350 114.600 729.000 ;
        RECT 103.950 724.950 106.050 727.050 ;
        RECT 106.950 724.950 109.050 727.050 ;
        RECT 109.950 724.950 112.050 727.050 ;
        RECT 112.950 724.950 115.050 727.050 ;
        RECT 104.400 722.400 105.600 724.650 ;
        RECT 110.400 723.900 111.600 724.650 ;
        RECT 104.400 718.050 105.450 722.400 ;
        RECT 109.950 721.800 112.050 723.900 ;
        RECT 103.950 715.950 106.050 718.050 ;
        RECT 119.400 715.050 120.450 748.950 ;
        RECT 125.400 733.050 126.450 800.400 ;
        RECT 142.950 796.950 145.050 801.000 ;
        RECT 169.950 796.950 172.050 801.000 ;
        RECT 143.400 787.050 144.450 796.950 ;
        RECT 170.400 790.050 171.450 796.950 ;
        RECT 174.150 794.700 175.350 813.300 ;
        RECT 179.100 802.950 181.200 805.050 ;
        RECT 179.400 801.900 180.600 802.650 ;
        RECT 178.950 799.800 181.050 801.900 ;
        RECT 191.550 800.400 192.750 813.300 ;
        RECT 205.950 811.950 208.050 814.050 ;
        RECT 196.950 806.100 199.050 808.200 ;
        RECT 197.400 805.350 198.600 806.100 ;
        RECT 196.950 802.950 199.050 805.050 ;
        RECT 206.400 802.050 207.450 811.950 ;
        RECT 217.950 808.950 220.050 814.050 ;
        RECT 277.950 811.950 280.050 814.050 ;
        RECT 313.950 811.950 316.050 814.050 ;
        RECT 344.850 813.300 346.950 815.400 ;
        RECT 362.550 813.300 364.650 815.400 ;
        RECT 394.950 814.950 397.050 817.050 ;
        RECT 409.950 814.950 412.050 817.050 ;
        RECT 385.950 813.450 388.050 814.050 ;
        RECT 391.950 813.450 394.050 814.050 ;
        RECT 223.950 810.450 226.050 811.050 ;
        RECT 223.950 809.400 234.450 810.450 ;
        RECT 223.950 808.950 226.050 809.400 ;
        RECT 211.950 806.100 214.050 808.200 ;
        RECT 220.950 806.100 223.050 808.200 ;
        RECT 226.950 806.100 229.050 808.200 ;
        RECT 233.400 807.600 234.450 809.400 ;
        RECT 212.400 805.350 213.600 806.100 ;
        RECT 211.950 802.950 214.050 805.050 ;
        RECT 214.950 802.950 217.050 805.050 ;
        RECT 191.550 798.300 193.650 800.400 ;
        RECT 205.950 799.950 208.050 802.050 ;
        RECT 215.400 801.900 216.600 802.650 ;
        RECT 214.950 799.800 217.050 801.900 ;
        RECT 174.150 793.500 178.350 794.700 ;
        RECT 176.250 792.600 178.350 793.500 ;
        RECT 191.550 791.700 192.750 798.300 ;
        RECT 221.400 793.050 222.450 806.100 ;
        RECT 227.400 805.350 228.600 806.100 ;
        RECT 233.400 805.350 234.600 807.600 ;
        RECT 241.950 805.950 244.050 808.050 ;
        RECT 250.950 806.100 253.050 808.200 ;
        RECT 268.950 806.100 271.050 808.200 ;
        RECT 226.950 802.950 229.050 805.050 ;
        RECT 229.950 802.950 232.050 805.050 ;
        RECT 232.950 802.950 235.050 805.050 ;
        RECT 235.950 802.950 238.050 805.050 ;
        RECT 230.400 801.900 231.600 802.650 ;
        RECT 236.400 801.900 237.600 802.650 ;
        RECT 242.400 801.900 243.450 805.950 ;
        RECT 251.400 805.350 252.600 806.100 ;
        RECT 269.400 805.350 270.600 806.100 ;
        RECT 247.950 802.950 250.050 805.050 ;
        RECT 250.950 802.950 253.050 805.050 ;
        RECT 253.950 802.950 256.050 805.050 ;
        RECT 259.950 802.950 262.050 805.050 ;
        RECT 265.950 802.950 268.050 805.050 ;
        RECT 268.950 802.950 271.050 805.050 ;
        RECT 271.950 802.950 274.050 805.050 ;
        RECT 229.950 799.800 232.050 801.900 ;
        RECT 235.950 799.800 238.050 801.900 ;
        RECT 241.950 799.800 244.050 801.900 ;
        RECT 248.400 800.400 249.600 802.650 ;
        RECT 254.400 800.400 255.600 802.650 ;
        RECT 169.950 787.950 172.050 790.050 ;
        RECT 191.550 789.600 193.650 791.700 ;
        RECT 220.950 790.950 223.050 793.050 ;
        RECT 221.400 787.050 222.450 790.950 ;
        RECT 248.400 787.050 249.450 800.400 ;
        RECT 254.400 793.050 255.450 800.400 ;
        RECT 260.400 796.050 261.450 802.950 ;
        RECT 266.400 800.400 267.600 802.650 ;
        RECT 272.400 801.900 273.600 802.650 ;
        RECT 278.400 801.900 279.450 811.950 ;
        RECT 289.950 806.100 292.050 808.200 ;
        RECT 290.400 805.350 291.600 806.100 ;
        RECT 301.950 805.950 304.050 808.050 ;
        RECT 314.400 807.600 315.450 811.950 ;
        RECT 287.100 802.950 289.200 805.050 ;
        RECT 290.400 802.950 292.500 805.050 ;
        RECT 295.800 802.950 297.900 805.050 ;
        RECT 266.400 796.050 267.450 800.400 ;
        RECT 271.950 799.800 274.050 801.900 ;
        RECT 277.950 799.800 280.050 801.900 ;
        RECT 287.400 800.400 288.600 802.650 ;
        RECT 296.400 801.900 297.600 802.650 ;
        RECT 274.950 796.950 277.050 799.050 ;
        RECT 259.950 793.950 262.050 796.050 ;
        RECT 265.950 793.950 268.050 796.050 ;
        RECT 275.400 793.050 276.450 796.950 ;
        RECT 253.950 790.950 256.050 793.050 ;
        RECT 267.000 792.900 270.000 793.050 ;
        RECT 265.950 790.950 271.050 792.900 ;
        RECT 274.950 790.950 277.050 793.050 ;
        RECT 265.950 790.800 268.050 790.950 ;
        RECT 268.950 790.800 271.050 790.950 ;
        RECT 142.950 784.950 145.050 787.050 ;
        RECT 193.950 784.950 196.050 787.050 ;
        RECT 220.950 784.950 223.050 787.050 ;
        RECT 247.950 784.950 250.050 787.050 ;
        RECT 268.950 784.950 271.050 787.050 ;
        RECT 154.950 781.950 157.050 784.050 ;
        RECT 145.950 769.950 148.050 772.050 ;
        RECT 130.950 761.100 133.050 763.200 ;
        RECT 146.400 763.050 147.450 769.950 ;
        RECT 148.950 766.950 151.050 769.050 ;
        RECT 137.400 762.450 138.600 762.600 ;
        RECT 137.400 761.400 144.450 762.450 ;
        RECT 131.400 760.350 132.600 761.100 ;
        RECT 137.400 760.350 138.600 761.400 ;
        RECT 130.950 757.950 133.050 760.050 ;
        RECT 133.950 757.950 136.050 760.050 ;
        RECT 136.950 757.950 139.050 760.050 ;
        RECT 134.400 756.000 135.600 757.650 ;
        RECT 133.950 751.950 136.050 756.000 ;
        RECT 139.950 754.950 142.050 757.050 ;
        RECT 140.400 748.050 141.450 754.950 ;
        RECT 127.950 745.950 130.050 748.050 ;
        RECT 139.950 745.950 142.050 748.050 ;
        RECT 124.950 730.950 127.050 733.050 ;
        RECT 128.400 729.600 129.450 745.950 ;
        RECT 143.400 742.050 144.450 761.400 ;
        RECT 145.950 760.950 148.050 763.050 ;
        RECT 149.400 762.600 150.450 766.950 ;
        RECT 155.400 762.600 156.450 781.950 ;
        RECT 194.400 781.050 195.450 784.950 ;
        RECT 193.950 778.950 196.050 781.050 ;
        RECT 181.950 775.950 184.050 778.050 ;
        RECT 169.950 769.950 172.050 772.050 ;
        RECT 170.400 763.200 171.450 769.950 ;
        RECT 175.950 766.950 178.050 769.050 ;
        RECT 149.400 760.350 150.600 762.600 ;
        RECT 155.400 760.350 156.600 762.600 ;
        RECT 160.950 761.100 163.050 763.200 ;
        RECT 169.950 761.100 172.050 763.200 ;
        RECT 176.400 762.600 177.450 766.950 ;
        RECT 182.400 762.600 183.450 775.950 ;
        RECT 187.950 769.950 190.050 772.050 ;
        RECT 188.400 762.600 189.450 769.950 ;
        RECT 194.400 762.600 195.450 778.950 ;
        RECT 200.250 769.500 202.350 770.400 ;
        RECT 211.950 769.950 214.050 772.050 ;
        RECT 215.550 771.300 217.650 773.400 ;
        RECT 198.150 768.300 202.350 769.500 ;
        RECT 161.400 760.350 162.600 761.100 ;
        RECT 148.950 757.950 151.050 760.050 ;
        RECT 151.950 757.950 154.050 760.050 ;
        RECT 154.950 757.950 157.050 760.050 ;
        RECT 157.950 757.950 160.050 760.050 ;
        RECT 160.950 757.950 163.050 760.050 ;
        RECT 152.400 756.900 153.600 757.650 ;
        RECT 151.950 754.800 154.050 756.900 ;
        RECT 158.400 756.000 159.600 757.650 ;
        RECT 148.950 751.950 151.050 754.050 ;
        RECT 157.950 751.950 160.050 756.000 ;
        RECT 170.400 754.050 171.450 761.100 ;
        RECT 176.400 760.350 177.600 762.600 ;
        RECT 182.400 760.350 183.600 762.600 ;
        RECT 188.400 760.350 189.600 762.600 ;
        RECT 194.400 760.350 195.600 762.600 ;
        RECT 175.950 757.950 178.050 760.050 ;
        RECT 178.950 757.950 181.050 760.050 ;
        RECT 181.950 757.950 184.050 760.050 ;
        RECT 184.950 757.950 187.050 760.050 ;
        RECT 187.950 757.950 190.050 760.050 ;
        RECT 193.950 757.950 196.050 760.050 ;
        RECT 179.400 755.400 180.600 757.650 ;
        RECT 185.400 755.400 186.600 757.650 ;
        RECT 169.950 751.950 172.050 754.050 ;
        RECT 145.950 742.950 148.050 745.050 ;
        RECT 142.950 739.950 145.050 742.050 ;
        RECT 146.400 738.450 147.450 742.950 ;
        RECT 143.400 737.400 147.450 738.450 ;
        RECT 139.350 735.300 141.450 737.400 ;
        RECT 128.400 727.350 129.600 729.600 ;
        RECT 133.950 729.000 136.050 733.050 ;
        RECT 134.400 727.350 135.600 729.000 ;
        RECT 124.950 724.950 127.050 727.050 ;
        RECT 127.950 724.950 130.050 727.050 ;
        RECT 133.950 724.950 136.050 727.050 ;
        RECT 125.400 723.900 126.600 724.650 ;
        RECT 124.950 721.800 127.050 723.900 ;
        RECT 140.250 722.400 141.450 735.300 ;
        RECT 139.350 720.300 141.450 722.400 ;
        RECT 118.950 712.950 121.050 715.050 ;
        RECT 140.250 713.700 141.450 720.300 ;
        RECT 97.950 706.950 100.050 709.050 ;
        RECT 103.950 697.950 106.050 700.050 ;
        RECT 16.950 688.950 19.050 691.050 ;
        RECT 55.950 688.950 58.050 691.050 ;
        RECT 64.950 688.950 67.050 691.050 ;
        RECT 10.950 682.950 13.050 685.050 ;
        RECT 17.400 684.600 18.450 688.950 ;
        RECT 17.400 682.350 18.600 684.600 ;
        RECT 22.950 682.950 25.050 685.050 ;
        RECT 31.950 683.100 34.050 685.200 ;
        RECT 40.950 683.100 43.050 685.200 ;
        RECT 46.950 683.100 49.050 685.200 ;
        RECT 52.950 683.100 55.050 685.200 ;
        RECT 58.950 683.100 61.050 685.200 ;
        RECT 65.400 684.600 66.450 688.950 ;
        RECT 13.950 679.950 16.050 682.050 ;
        RECT 16.950 679.950 19.050 682.050 ;
        RECT 14.400 678.900 15.600 679.650 ;
        RECT 23.400 678.900 24.450 682.950 ;
        RECT 32.400 682.350 33.600 683.100 ;
        RECT 28.950 679.950 31.050 682.050 ;
        RECT 31.950 679.950 34.050 682.050 ;
        RECT 34.950 679.950 37.050 682.050 ;
        RECT 13.950 676.800 16.050 678.900 ;
        RECT 22.950 676.800 25.050 678.900 ;
        RECT 29.400 677.400 30.600 679.650 ;
        RECT 35.400 678.900 36.600 679.650 ;
        RECT 41.400 679.050 42.450 683.100 ;
        RECT 47.400 682.350 48.600 683.100 ;
        RECT 53.400 682.350 54.600 683.100 ;
        RECT 46.950 679.950 49.050 682.050 ;
        RECT 49.950 679.950 52.050 682.050 ;
        RECT 52.950 679.950 55.050 682.050 ;
        RECT 29.400 673.050 30.450 677.400 ;
        RECT 34.950 676.800 37.050 678.900 ;
        RECT 40.950 676.950 43.050 679.050 ;
        RECT 50.400 678.900 51.600 679.650 ;
        RECT 28.950 670.950 31.050 673.050 ;
        RECT 41.400 667.050 42.450 676.950 ;
        RECT 49.950 676.800 52.050 678.900 ;
        RECT 59.400 673.050 60.450 683.100 ;
        RECT 65.400 682.350 66.600 684.600 ;
        RECT 70.950 683.100 73.050 685.200 ;
        RECT 76.950 683.100 79.050 685.200 ;
        RECT 85.950 683.100 88.050 685.200 ;
        RECT 91.950 683.100 94.050 685.200 ;
        RECT 97.950 683.100 100.050 685.200 ;
        RECT 104.400 684.600 105.450 697.950 ;
        RECT 109.950 694.950 112.050 697.050 ;
        RECT 119.400 696.450 120.450 712.950 ;
        RECT 139.350 711.600 141.450 713.700 ;
        RECT 133.950 706.950 136.050 709.050 ;
        RECT 116.400 695.400 120.450 696.450 ;
        RECT 110.400 685.200 111.450 694.950 ;
        RECT 71.400 682.350 72.600 683.100 ;
        RECT 64.950 679.950 67.050 682.050 ;
        RECT 67.950 679.950 70.050 682.050 ;
        RECT 70.950 679.950 73.050 682.050 ;
        RECT 68.400 678.900 69.600 679.650 ;
        RECT 77.400 679.050 78.450 683.100 ;
        RECT 86.400 682.350 87.600 683.100 ;
        RECT 92.400 682.350 93.600 683.100 ;
        RECT 82.950 679.950 85.050 682.050 ;
        RECT 85.950 679.950 88.050 682.050 ;
        RECT 88.950 679.950 91.050 682.050 ;
        RECT 91.950 679.950 94.050 682.050 ;
        RECT 67.950 676.800 70.050 678.900 ;
        RECT 76.950 676.950 79.050 679.050 ;
        RECT 83.400 677.400 84.600 679.650 ;
        RECT 89.400 678.000 90.600 679.650 ;
        RECT 58.950 670.950 61.050 673.050 ;
        RECT 40.950 664.950 43.050 667.050 ;
        RECT 55.950 664.950 58.050 667.050 ;
        RECT 7.950 655.950 10.050 658.050 ;
        RECT 46.950 655.950 49.050 658.050 ;
        RECT 13.950 650.100 16.050 652.200 ;
        RECT 33.000 651.600 37.050 652.050 ;
        RECT 14.400 649.350 15.600 650.100 ;
        RECT 32.400 649.950 37.050 651.600 ;
        RECT 37.950 649.950 40.050 652.050 ;
        RECT 47.400 651.600 48.450 655.950 ;
        RECT 32.400 649.350 33.600 649.950 ;
        RECT 10.950 646.950 13.050 649.050 ;
        RECT 13.950 646.950 16.050 649.050 ;
        RECT 16.950 646.950 19.050 649.050 ;
        RECT 28.950 646.950 31.050 649.050 ;
        RECT 31.950 646.950 34.050 649.050 ;
        RECT 11.400 645.900 12.600 646.650 ;
        RECT 10.950 643.800 13.050 645.900 ;
        RECT 17.400 644.400 18.600 646.650 ;
        RECT 29.400 645.900 30.600 646.650 ;
        RECT 38.400 645.900 39.450 649.950 ;
        RECT 47.400 649.350 48.600 651.600 ;
        RECT 43.950 646.950 46.050 649.050 ;
        RECT 46.950 646.950 49.050 649.050 ;
        RECT 49.950 646.950 52.050 649.050 ;
        RECT 17.400 619.050 18.450 644.400 ;
        RECT 28.950 643.800 31.050 645.900 ;
        RECT 37.950 643.800 40.050 645.900 ;
        RECT 40.950 643.950 43.050 646.050 ;
        RECT 44.400 645.900 45.600 646.650 ;
        RECT 16.950 616.950 19.050 619.050 ;
        RECT 41.400 607.200 42.450 643.950 ;
        RECT 43.950 643.800 46.050 645.900 ;
        RECT 50.400 644.400 51.600 646.650 ;
        RECT 50.400 642.450 51.450 644.400 ;
        RECT 52.950 643.950 55.050 646.050 ;
        RECT 47.400 641.400 51.450 642.450 ;
        RECT 14.400 606.450 15.600 606.600 ;
        RECT 11.400 605.400 15.600 606.450 ;
        RECT 11.400 597.450 12.450 605.400 ;
        RECT 14.400 604.350 15.600 605.400 ;
        RECT 22.950 605.100 25.050 607.200 ;
        RECT 23.400 604.350 24.600 605.100 ;
        RECT 28.950 604.950 31.050 607.050 ;
        RECT 34.950 605.100 37.050 607.200 ;
        RECT 40.950 605.100 43.050 607.200 ;
        RECT 14.100 601.950 16.200 604.050 ;
        RECT 19.500 601.950 21.600 604.050 ;
        RECT 22.800 601.950 24.900 604.050 ;
        RECT 20.400 599.400 21.600 601.650 ;
        RECT 29.400 600.900 30.450 604.950 ;
        RECT 35.400 604.350 36.600 605.100 ;
        RECT 41.400 604.350 42.600 605.100 ;
        RECT 34.950 601.950 37.050 604.050 ;
        RECT 37.950 601.950 40.050 604.050 ;
        RECT 40.950 601.950 43.050 604.050 ;
        RECT 11.400 596.400 15.450 597.450 ;
        RECT 14.400 573.600 15.450 596.400 ;
        RECT 20.400 595.050 21.450 599.400 ;
        RECT 28.950 598.800 31.050 600.900 ;
        RECT 38.400 599.400 39.600 601.650 ;
        RECT 38.400 598.050 39.450 599.400 ;
        RECT 43.950 598.950 46.050 601.050 ;
        RECT 37.950 595.950 40.050 598.050 ;
        RECT 19.950 592.950 22.050 595.050 ;
        RECT 34.950 583.950 37.050 586.050 ;
        RECT 14.400 571.350 15.600 573.600 ;
        RECT 22.950 572.100 25.050 574.200 ;
        RECT 28.950 572.100 31.050 574.200 ;
        RECT 35.400 573.600 36.450 583.950 ;
        RECT 38.400 580.050 39.450 595.950 ;
        RECT 44.400 586.050 45.450 598.950 ;
        RECT 47.400 598.050 48.450 641.400 ;
        RECT 53.400 627.450 54.450 643.950 ;
        RECT 50.400 626.400 54.450 627.450 ;
        RECT 50.400 607.050 51.450 626.400 ;
        RECT 56.400 625.050 57.450 664.950 ;
        RECT 59.400 661.050 60.450 670.950 ;
        RECT 83.400 664.050 84.450 677.400 ;
        RECT 88.950 673.950 91.050 678.000 ;
        RECT 98.400 670.050 99.450 683.100 ;
        RECT 104.400 682.350 105.600 684.600 ;
        RECT 109.950 683.100 112.050 685.200 ;
        RECT 116.400 684.600 117.450 695.400 ;
        RECT 122.250 691.500 124.350 692.400 ;
        RECT 120.150 690.300 124.350 691.500 ;
        RECT 110.400 682.350 111.600 683.100 ;
        RECT 116.400 682.350 117.600 684.600 ;
        RECT 103.950 679.950 106.050 682.050 ;
        RECT 106.950 679.950 109.050 682.050 ;
        RECT 109.950 679.950 112.050 682.050 ;
        RECT 115.950 679.950 118.050 682.050 ;
        RECT 107.400 677.400 108.600 679.650 ;
        RECT 97.950 667.950 100.050 670.050 ;
        RECT 82.950 661.950 85.050 664.050 ;
        RECT 58.950 658.950 61.050 661.050 ;
        RECT 73.950 658.950 76.050 661.050 ;
        RECT 61.950 650.100 64.050 652.200 ;
        RECT 68.400 651.450 69.600 651.600 ;
        RECT 70.950 651.450 73.050 655.050 ;
        RECT 68.400 651.000 73.050 651.450 ;
        RECT 68.400 650.400 72.450 651.000 ;
        RECT 62.400 649.350 63.600 650.100 ;
        RECT 68.400 649.350 69.600 650.400 ;
        RECT 61.950 646.950 64.050 649.050 ;
        RECT 64.950 646.950 67.050 649.050 ;
        RECT 67.950 646.950 70.050 649.050 ;
        RECT 65.400 645.900 66.600 646.650 ;
        RECT 64.950 643.800 67.050 645.900 ;
        RECT 55.950 622.950 58.050 625.050 ;
        RECT 61.950 622.950 64.050 625.050 ;
        RECT 55.950 616.950 58.050 619.050 ;
        RECT 56.400 607.050 57.450 616.950 ;
        RECT 49.950 604.950 52.050 607.050 ;
        RECT 56.400 604.950 61.050 607.050 ;
        RECT 56.400 604.350 57.600 604.950 ;
        RECT 52.950 601.950 55.050 604.050 ;
        RECT 55.950 601.950 58.050 604.050 ;
        RECT 53.400 600.900 54.600 601.650 ;
        RECT 52.950 598.800 55.050 600.900 ;
        RECT 46.950 595.950 49.050 598.050 ;
        RECT 46.950 592.800 49.050 594.900 ;
        RECT 43.950 583.950 46.050 586.050 ;
        RECT 37.950 577.950 40.050 580.050 ;
        RECT 43.950 577.950 46.050 580.050 ;
        RECT 10.950 568.950 13.050 571.050 ;
        RECT 13.950 568.950 16.050 571.050 ;
        RECT 16.950 568.950 19.050 571.050 ;
        RECT 11.400 566.400 12.600 568.650 ;
        RECT 17.400 567.900 18.600 568.650 ;
        RECT 23.400 568.050 24.450 572.100 ;
        RECT 29.400 571.350 30.600 572.100 ;
        RECT 35.400 571.350 36.600 573.600 ;
        RECT 28.950 568.950 31.050 571.050 ;
        RECT 31.950 568.950 34.050 571.050 ;
        RECT 34.950 568.950 37.050 571.050 ;
        RECT 37.950 568.950 40.050 571.050 ;
        RECT 11.400 556.050 12.450 566.400 ;
        RECT 16.950 565.800 19.050 567.900 ;
        RECT 22.950 565.950 25.050 568.050 ;
        RECT 32.400 566.400 33.600 568.650 ;
        RECT 38.400 567.900 39.600 568.650 ;
        RECT 44.400 567.900 45.450 577.950 ;
        RECT 47.400 577.050 48.450 592.800 ;
        RECT 52.950 583.950 55.050 586.050 ;
        RECT 46.950 574.950 49.050 577.050 ;
        RECT 10.950 555.450 13.050 556.050 ;
        RECT 8.400 554.400 13.050 555.450 ;
        RECT 1.950 541.950 4.050 544.050 ;
        RECT 2.400 418.050 3.450 541.950 ;
        RECT 8.400 529.050 9.450 554.400 ;
        RECT 10.950 553.950 13.050 554.400 ;
        RECT 17.400 529.050 18.450 565.800 ;
        RECT 28.950 559.950 31.050 562.050 ;
        RECT 25.350 537.300 27.450 539.400 ;
        RECT 26.250 530.700 27.450 537.300 ;
        RECT 7.950 526.950 10.050 529.050 ;
        RECT 14.400 528.450 15.600 528.600 ;
        RECT 16.950 528.450 19.050 529.050 ;
        RECT 25.350 528.600 27.450 530.700 ;
        RECT 14.400 527.400 19.050 528.450 ;
        RECT 14.400 526.350 15.600 527.400 ;
        RECT 16.950 526.950 19.050 527.400 ;
        RECT 10.950 523.950 13.050 526.050 ;
        RECT 13.950 523.950 16.050 526.050 ;
        RECT 19.950 523.950 22.050 526.050 ;
        RECT 7.950 520.950 10.050 523.050 ;
        RECT 11.400 521.400 12.600 523.650 ;
        RECT 20.400 522.000 21.600 523.650 ;
        RECT 8.400 496.050 9.450 520.950 ;
        RECT 11.400 520.050 12.450 521.400 ;
        RECT 10.950 517.950 13.050 520.050 ;
        RECT 19.950 517.950 22.050 522.000 ;
        RECT 11.400 499.050 12.450 517.950 ;
        RECT 26.250 515.700 27.450 528.600 ;
        RECT 25.350 513.600 27.450 515.700 ;
        RECT 25.950 508.950 28.050 511.050 ;
        RECT 13.950 502.950 16.050 505.050 ;
        RECT 10.950 496.950 13.050 499.050 ;
        RECT 7.950 493.950 10.050 496.050 ;
        RECT 14.400 495.600 15.450 502.950 ;
        RECT 14.400 493.350 15.600 495.600 ;
        RECT 22.950 493.950 25.050 496.050 ;
        RECT 10.950 490.950 13.050 493.050 ;
        RECT 13.950 490.950 16.050 493.050 ;
        RECT 16.950 490.950 19.050 493.050 ;
        RECT 7.950 487.950 10.050 490.050 ;
        RECT 11.400 489.000 12.600 490.650 ;
        RECT 4.950 451.950 7.050 454.050 ;
        RECT 5.400 421.050 6.450 451.950 ;
        RECT 8.400 430.050 9.450 487.950 ;
        RECT 10.950 484.950 13.050 489.000 ;
        RECT 17.400 488.400 18.600 490.650 ;
        RECT 23.400 489.900 24.450 493.950 ;
        RECT 17.400 454.050 18.450 488.400 ;
        RECT 22.950 487.800 25.050 489.900 ;
        RECT 19.950 478.950 22.050 481.050 ;
        RECT 16.950 451.950 19.050 454.050 ;
        RECT 20.400 451.050 21.450 478.950 ;
        RECT 26.400 462.450 27.450 508.950 ;
        RECT 29.400 505.050 30.450 559.950 ;
        RECT 32.400 556.050 33.450 566.400 ;
        RECT 37.950 565.800 40.050 567.900 ;
        RECT 43.950 565.800 46.050 567.900 ;
        RECT 47.400 562.050 48.450 574.950 ;
        RECT 53.400 573.600 54.450 583.950 ;
        RECT 58.950 580.950 61.050 583.050 ;
        RECT 59.400 574.050 60.450 580.950 ;
        RECT 53.400 571.350 54.600 573.600 ;
        RECT 58.950 571.950 61.050 574.050 ;
        RECT 52.950 568.950 55.050 571.050 ;
        RECT 55.950 568.950 58.050 571.050 ;
        RECT 56.400 566.400 57.600 568.650 ;
        RECT 56.400 562.050 57.450 566.400 ;
        RECT 58.950 565.950 61.050 568.050 ;
        RECT 46.950 559.950 49.050 562.050 ;
        RECT 55.950 559.950 58.050 562.050 ;
        RECT 31.950 553.950 34.050 556.050 ;
        RECT 59.400 550.050 60.450 565.950 ;
        RECT 58.950 547.950 61.050 550.050 ;
        RECT 40.650 535.500 42.750 536.400 ;
        RECT 40.650 534.300 44.850 535.500 ;
        RECT 31.950 526.950 34.050 529.050 ;
        RECT 37.950 527.100 40.050 529.200 ;
        RECT 28.950 502.950 31.050 505.050 ;
        RECT 32.400 498.450 33.450 526.950 ;
        RECT 38.400 526.350 39.600 527.100 ;
        RECT 37.800 523.950 39.900 526.050 ;
        RECT 37.950 517.950 40.050 520.050 ;
        RECT 29.400 498.000 33.450 498.450 ;
        RECT 28.950 497.400 33.450 498.000 ;
        RECT 28.950 493.950 31.050 497.400 ;
        RECT 31.950 494.100 34.050 496.200 ;
        RECT 38.400 495.600 39.450 517.950 ;
        RECT 43.650 515.700 44.850 534.300 ;
        RECT 46.950 528.000 49.050 532.050 ;
        RECT 52.950 529.950 55.050 532.050 ;
        RECT 62.400 531.450 63.450 622.950 ;
        RECT 70.950 610.950 73.050 613.050 ;
        RECT 71.400 606.600 72.450 610.950 ;
        RECT 74.400 610.050 75.450 658.950 ;
        RECT 82.950 655.950 85.050 658.050 ;
        RECT 91.950 655.950 94.050 658.050 ;
        RECT 83.400 651.600 84.450 655.950 ;
        RECT 83.400 649.350 84.600 651.600 ;
        RECT 88.950 650.100 91.050 652.200 ;
        RECT 92.400 652.050 93.450 655.950 ;
        RECT 94.950 652.950 97.050 655.050 ;
        RECT 89.400 649.350 90.600 650.100 ;
        RECT 91.950 649.950 94.050 652.050 ;
        RECT 79.950 646.950 82.050 649.050 ;
        RECT 82.950 646.950 85.050 649.050 ;
        RECT 85.950 646.950 88.050 649.050 ;
        RECT 88.950 646.950 91.050 649.050 ;
        RECT 80.400 645.900 81.600 646.650 ;
        RECT 79.950 643.800 82.050 645.900 ;
        RECT 86.400 644.400 87.600 646.650 ;
        RECT 86.400 631.050 87.450 644.400 ;
        RECT 85.950 628.950 88.050 631.050 ;
        RECT 73.950 607.950 76.050 610.050 ;
        RECT 82.950 607.950 85.050 610.050 ;
        RECT 71.400 604.350 72.600 606.600 ;
        RECT 67.950 601.950 70.050 604.050 ;
        RECT 70.950 601.950 73.050 604.050 ;
        RECT 73.950 601.950 76.050 604.050 ;
        RECT 64.950 598.950 67.050 601.050 ;
        RECT 68.400 600.000 69.600 601.650 ;
        RECT 65.400 574.050 66.450 598.950 ;
        RECT 67.950 595.950 70.050 600.000 ;
        RECT 74.400 599.400 75.600 601.650 ;
        RECT 74.400 589.050 75.450 599.400 ;
        RECT 73.950 586.950 76.050 589.050 ;
        RECT 73.950 580.950 76.050 583.050 ;
        RECT 79.950 580.950 82.050 583.050 ;
        RECT 64.950 571.950 67.050 574.050 ;
        RECT 67.950 573.000 70.050 577.050 ;
        RECT 74.400 573.600 75.450 580.950 ;
        RECT 80.400 574.050 81.450 580.950 ;
        RECT 68.400 571.350 69.600 573.000 ;
        RECT 74.400 571.350 75.600 573.600 ;
        RECT 79.950 571.950 82.050 574.050 ;
        RECT 67.950 568.950 70.050 571.050 ;
        RECT 70.950 568.950 73.050 571.050 ;
        RECT 73.950 568.950 76.050 571.050 ;
        RECT 76.950 568.950 79.050 571.050 ;
        RECT 64.950 565.950 67.050 568.050 ;
        RECT 71.400 567.900 72.600 568.650 ;
        RECT 77.400 568.050 78.600 568.650 ;
        RECT 65.400 535.050 66.450 565.950 ;
        RECT 70.950 565.800 73.050 567.900 ;
        RECT 77.400 566.400 82.050 568.050 ;
        RECT 78.000 565.950 82.050 566.400 ;
        RECT 79.950 553.950 82.050 556.050 ;
        RECT 80.400 544.050 81.450 553.950 ;
        RECT 79.950 541.950 82.050 544.050 ;
        RECT 76.350 537.300 78.450 539.400 ;
        RECT 64.950 532.950 67.050 535.050 ;
        RECT 62.400 530.400 66.450 531.450 ;
        RECT 77.250 530.700 78.450 537.300 ;
        RECT 79.950 532.950 82.050 535.050 ;
        RECT 47.400 526.350 48.600 528.000 ;
        RECT 46.950 523.950 49.050 526.050 ;
        RECT 43.050 513.600 45.150 515.700 ;
        RECT 53.400 511.050 54.450 529.950 ;
        RECT 65.400 529.200 66.450 530.400 ;
        RECT 64.950 527.100 67.050 529.200 ;
        RECT 76.350 528.600 78.450 530.700 ;
        RECT 65.400 526.350 66.600 527.100 ;
        RECT 61.950 523.950 64.050 526.050 ;
        RECT 64.950 523.950 67.050 526.050 ;
        RECT 70.950 523.950 73.050 526.050 ;
        RECT 62.400 522.900 63.600 523.650 ;
        RECT 71.400 523.050 72.600 523.650 ;
        RECT 69.000 522.900 72.600 523.050 ;
        RECT 61.950 520.800 64.050 522.900 ;
        RECT 67.950 521.400 72.600 522.900 ;
        RECT 67.950 520.950 72.000 521.400 ;
        RECT 67.950 520.800 70.050 520.950 ;
        RECT 77.250 515.700 78.450 528.600 ;
        RECT 76.350 513.600 78.450 515.700 ;
        RECT 52.950 508.950 55.050 511.050 ;
        RECT 80.400 510.450 81.450 532.950 ;
        RECT 77.400 509.400 81.450 510.450 ;
        RECT 70.950 505.950 73.050 508.050 ;
        RECT 71.400 496.200 72.450 505.950 ;
        RECT 32.400 493.350 33.600 494.100 ;
        RECT 38.400 493.350 39.600 495.600 ;
        RECT 46.950 493.950 49.050 496.050 ;
        RECT 55.950 494.100 58.050 496.200 ;
        RECT 64.950 494.100 67.050 496.200 ;
        RECT 70.950 494.100 73.050 496.200 ;
        RECT 77.400 495.600 78.450 509.400 ;
        RECT 31.950 490.950 34.050 493.050 ;
        RECT 34.950 490.950 37.050 493.050 ;
        RECT 37.950 490.950 40.050 493.050 ;
        RECT 40.950 490.950 43.050 493.050 ;
        RECT 35.400 489.900 36.600 490.650 ;
        RECT 34.950 487.800 37.050 489.900 ;
        RECT 41.400 489.000 42.600 490.650 ;
        RECT 40.950 484.950 43.050 489.000 ;
        RECT 47.400 487.050 48.450 493.950 ;
        RECT 56.400 493.350 57.600 494.100 ;
        RECT 52.950 490.950 55.050 493.050 ;
        RECT 55.950 490.950 58.050 493.050 ;
        RECT 58.950 490.950 61.050 493.050 ;
        RECT 53.400 489.900 54.600 490.650 ;
        RECT 52.950 487.800 55.050 489.900 ;
        RECT 59.400 488.400 60.600 490.650 ;
        RECT 46.950 484.950 49.050 487.050 ;
        RECT 53.400 481.050 54.450 487.800 ;
        RECT 52.950 478.950 55.050 481.050 ;
        RECT 59.400 475.050 60.450 488.400 ;
        RECT 58.950 472.950 61.050 475.050 ;
        RECT 65.400 469.050 66.450 494.100 ;
        RECT 71.400 493.350 72.600 494.100 ;
        RECT 77.400 493.350 78.600 495.600 ;
        RECT 83.400 495.450 84.450 607.950 ;
        RECT 85.950 605.100 88.050 607.200 ;
        RECT 95.400 606.600 96.450 652.950 ;
        RECT 103.950 651.000 106.050 655.050 ;
        RECT 107.400 652.050 108.450 677.400 ;
        RECT 112.950 676.950 115.050 679.050 ;
        RECT 113.400 663.450 114.450 676.950 ;
        RECT 120.150 671.700 121.350 690.300 ;
        RECT 124.950 683.100 127.050 685.200 ;
        RECT 125.400 682.350 126.600 683.100 ;
        RECT 125.100 679.950 127.200 682.050 ;
        RECT 119.850 669.600 121.950 671.700 ;
        RECT 134.400 666.450 135.450 706.950 ;
        RECT 143.400 697.050 144.450 737.400 ;
        RECT 149.400 735.450 150.450 751.950 ;
        RECT 179.400 745.050 180.450 755.400 ;
        RECT 181.950 751.950 184.050 754.050 ;
        RECT 178.950 742.950 181.050 745.050 ;
        RECT 146.400 734.400 150.450 735.450 ;
        RECT 157.050 735.300 159.150 737.400 ;
        RECT 169.950 736.950 172.050 739.050 ;
        RECT 146.400 723.450 147.450 734.400 ;
        RECT 151.800 724.950 153.900 727.050 ;
        RECT 146.400 722.400 150.450 723.450 ;
        RECT 152.400 723.000 153.600 724.650 ;
        RECT 137.550 693.300 139.650 695.400 ;
        RECT 142.950 694.950 145.050 697.050 ;
        RECT 137.550 686.700 138.750 693.300 ;
        RECT 149.400 691.050 150.450 722.400 ;
        RECT 151.950 718.950 154.050 723.000 ;
        RECT 157.650 716.700 158.850 735.300 ;
        RECT 166.950 730.950 169.050 736.050 ;
        RECT 166.950 727.800 169.050 729.900 ;
        RECT 160.950 724.950 163.050 727.050 ;
        RECT 154.650 715.500 158.850 716.700 ;
        RECT 161.400 722.400 162.600 724.650 ;
        RECT 154.650 714.600 156.750 715.500 ;
        RECT 161.400 715.050 162.450 722.400 ;
        RECT 167.400 718.050 168.450 727.800 ;
        RECT 166.950 715.950 169.050 718.050 ;
        RECT 160.950 712.950 163.050 715.050 ;
        RECT 151.950 697.950 154.050 700.050 ;
        RECT 148.950 688.950 151.050 691.050 ;
        RECT 137.550 684.600 139.650 686.700 ;
        RECT 137.550 671.700 138.750 684.600 ;
        RECT 142.950 679.950 145.050 682.050 ;
        RECT 143.400 678.900 144.600 679.650 ;
        RECT 149.400 678.900 150.450 688.950 ;
        RECT 152.400 685.200 153.450 697.950 ;
        RECT 163.950 688.950 166.050 691.050 ;
        RECT 151.950 683.100 154.050 685.200 ;
        RECT 157.950 683.100 160.050 685.200 ;
        RECT 164.400 684.600 165.450 688.950 ;
        RECT 142.950 676.800 145.050 678.900 ;
        RECT 148.950 676.800 151.050 678.900 ;
        RECT 137.550 669.600 139.650 671.700 ;
        RECT 134.400 665.400 138.450 666.450 ;
        RECT 110.400 662.400 114.450 663.450 ;
        RECT 104.400 649.350 105.600 651.000 ;
        RECT 106.950 649.950 109.050 652.050 ;
        RECT 110.400 651.600 111.450 662.400 ;
        RECT 115.350 657.300 117.450 659.400 ;
        RECT 133.050 657.300 135.150 659.400 ;
        RECT 110.400 649.350 111.600 651.600 ;
        RECT 100.950 646.950 103.050 649.050 ;
        RECT 103.950 646.950 106.050 649.050 ;
        RECT 109.950 646.950 112.050 649.050 ;
        RECT 97.950 643.950 100.050 646.050 ;
        RECT 101.400 644.400 102.600 646.650 ;
        RECT 116.250 644.400 117.450 657.300 ;
        RECT 127.800 646.950 129.900 649.050 ;
        RECT 128.400 645.450 129.600 646.650 ;
        RECT 98.400 640.050 99.450 643.950 ;
        RECT 97.950 637.950 100.050 640.050 ;
        RECT 97.950 628.950 100.050 631.050 ;
        RECT 86.400 604.350 87.600 605.100 ;
        RECT 95.400 604.350 96.600 606.600 ;
        RECT 86.100 601.950 88.200 604.050 ;
        RECT 91.500 601.950 93.600 604.050 ;
        RECT 94.800 601.950 96.900 604.050 ;
        RECT 92.400 599.400 93.600 601.650 ;
        RECT 85.950 586.950 88.050 589.050 ;
        RECT 86.400 574.050 87.450 586.950 ;
        RECT 92.400 583.050 93.450 599.400 ;
        RECT 98.400 597.450 99.450 628.950 ;
        RECT 101.400 615.450 102.450 644.400 ;
        RECT 115.350 642.300 117.450 644.400 ;
        RECT 116.250 635.700 117.450 642.300 ;
        RECT 125.400 644.400 129.600 645.450 ;
        RECT 125.400 640.050 126.450 644.400 ;
        RECT 124.950 637.950 127.050 640.050 ;
        RECT 133.650 638.700 134.850 657.300 ;
        RECT 137.400 655.050 138.450 665.400 ;
        RECT 142.950 661.950 145.050 664.050 ;
        RECT 143.400 655.050 144.450 661.950 ;
        RECT 152.400 655.050 153.450 683.100 ;
        RECT 158.400 682.350 159.600 683.100 ;
        RECT 164.400 682.350 165.600 684.600 ;
        RECT 157.950 679.950 160.050 682.050 ;
        RECT 160.950 679.950 163.050 682.050 ;
        RECT 163.950 679.950 166.050 682.050 ;
        RECT 161.400 677.400 162.600 679.650 ;
        RECT 161.400 670.050 162.450 677.400 ;
        RECT 170.400 676.050 171.450 736.950 ;
        RECT 172.950 733.950 175.050 736.050 ;
        RECT 173.400 730.050 174.450 733.950 ;
        RECT 172.950 727.950 175.050 730.050 ;
        RECT 175.950 729.000 178.050 733.050 ;
        RECT 182.400 730.200 183.450 751.950 ;
        RECT 185.400 748.050 186.450 755.400 ;
        RECT 198.150 749.700 199.350 768.300 ;
        RECT 208.950 766.950 211.050 769.050 ;
        RECT 202.950 761.100 205.050 763.200 ;
        RECT 203.400 760.350 204.600 761.100 ;
        RECT 203.100 757.950 205.200 760.050 ;
        RECT 184.950 745.950 187.050 748.050 ;
        RECT 197.850 747.600 199.950 749.700 ;
        RECT 193.950 733.950 196.050 736.050 ;
        RECT 199.950 733.950 202.050 736.050 ;
        RECT 176.400 727.350 177.600 729.000 ;
        RECT 181.950 728.100 184.050 730.200 ;
        RECT 187.950 728.100 190.050 730.200 ;
        RECT 194.400 729.600 195.450 733.950 ;
        RECT 200.400 729.600 201.450 733.950 ;
        RECT 182.400 727.350 183.600 728.100 ;
        RECT 175.950 724.950 178.050 727.050 ;
        RECT 178.950 724.950 181.050 727.050 ;
        RECT 181.950 724.950 184.050 727.050 ;
        RECT 179.400 723.900 180.600 724.650 ;
        RECT 178.950 721.800 181.050 723.900 ;
        RECT 188.400 709.050 189.450 728.100 ;
        RECT 194.400 727.350 195.600 729.600 ;
        RECT 200.400 727.350 201.600 729.600 ;
        RECT 193.950 724.950 196.050 727.050 ;
        RECT 196.950 724.950 199.050 727.050 ;
        RECT 199.950 724.950 202.050 727.050 ;
        RECT 202.950 724.950 205.050 727.050 ;
        RECT 197.400 723.900 198.600 724.650 ;
        RECT 196.950 721.800 199.050 723.900 ;
        RECT 203.400 722.400 204.600 724.650 ;
        RECT 199.950 718.950 202.050 721.050 ;
        RECT 187.950 706.950 190.050 709.050 ;
        RECT 184.950 684.000 187.050 688.050 ;
        RECT 190.950 685.950 193.050 688.050 ;
        RECT 185.400 682.350 186.600 684.000 ;
        RECT 179.100 679.950 181.200 682.050 ;
        RECT 185.100 679.950 187.200 682.050 ;
        RECT 179.400 677.400 180.600 679.650 ;
        RECT 169.950 673.950 172.050 676.050 ;
        RECT 179.400 670.050 180.450 677.400 ;
        RECT 160.950 667.950 163.050 670.050 ;
        RECT 172.950 667.950 175.050 670.050 ;
        RECT 178.950 667.950 181.050 670.050 ;
        RECT 169.350 657.300 171.450 659.400 ;
        RECT 136.950 652.950 139.050 655.050 ;
        RECT 142.950 652.950 145.050 655.050 ;
        RECT 145.950 652.950 148.050 655.050 ;
        RECT 151.950 652.950 154.050 655.050 ;
        RECT 136.950 646.950 139.050 649.050 ;
        RECT 130.650 637.500 134.850 638.700 ;
        RECT 137.400 644.400 138.600 646.650 ;
        RECT 130.650 636.600 132.750 637.500 ;
        RECT 115.350 633.600 117.450 635.700 ;
        RECT 137.400 619.050 138.450 644.400 ;
        RECT 143.400 640.050 144.450 652.950 ;
        RECT 146.400 645.900 147.450 652.950 ;
        RECT 154.950 650.100 157.050 652.200 ;
        RECT 163.950 651.000 166.050 655.050 ;
        RECT 155.400 649.350 156.600 650.100 ;
        RECT 164.400 649.350 165.600 651.000 ;
        RECT 151.950 646.950 154.050 649.050 ;
        RECT 154.950 646.950 157.050 649.050 ;
        RECT 157.950 646.950 160.050 649.050 ;
        RECT 163.950 646.950 166.050 649.050 ;
        RECT 152.400 645.900 153.600 646.650 ;
        RECT 145.950 643.800 148.050 645.900 ;
        RECT 151.950 643.800 154.050 645.900 ;
        RECT 158.400 644.400 159.600 646.650 ;
        RECT 170.250 644.400 171.450 657.300 ;
        RECT 158.400 640.050 159.450 644.400 ;
        RECT 169.350 642.300 171.450 644.400 ;
        RECT 142.950 637.950 145.050 640.050 ;
        RECT 148.950 637.950 151.050 640.050 ;
        RECT 157.950 637.950 160.050 640.050 ;
        RECT 136.950 616.950 139.050 619.050 ;
        RECT 101.400 614.400 105.450 615.450 ;
        RECT 145.350 615.300 147.450 617.400 ;
        RECT 100.950 610.950 103.050 613.050 ;
        RECT 95.400 596.400 99.450 597.450 ;
        RECT 91.950 580.950 94.050 583.050 ;
        RECT 95.400 579.450 96.450 596.400 ;
        RECT 97.950 586.950 100.050 589.050 ;
        RECT 92.400 578.400 96.450 579.450 ;
        RECT 85.950 571.950 88.050 574.050 ;
        RECT 92.400 573.600 93.450 578.400 ;
        RECT 98.400 573.600 99.450 586.950 ;
        RECT 101.400 574.050 102.450 610.950 ;
        RECT 104.400 589.050 105.450 614.400 ;
        RECT 146.250 608.700 147.450 615.300 ;
        RECT 106.950 605.100 109.050 607.200 ;
        RECT 115.950 605.100 118.050 607.200 ;
        RECT 121.950 605.100 124.050 607.200 ;
        RECT 127.950 605.100 130.050 607.200 ;
        RECT 133.950 605.100 136.050 607.200 ;
        RECT 145.350 606.600 147.450 608.700 ;
        RECT 107.400 604.350 108.600 605.100 ;
        RECT 116.400 604.350 117.600 605.100 ;
        RECT 107.100 601.950 109.200 604.050 ;
        RECT 112.500 601.950 114.600 604.050 ;
        RECT 115.800 601.950 117.900 604.050 ;
        RECT 113.400 600.000 114.600 601.650 ;
        RECT 112.950 595.950 115.050 600.000 ;
        RECT 122.400 598.050 123.450 605.100 ;
        RECT 128.400 604.350 129.600 605.100 ;
        RECT 134.400 604.350 135.600 605.100 ;
        RECT 127.950 601.950 130.050 604.050 ;
        RECT 130.950 601.950 133.050 604.050 ;
        RECT 133.950 601.950 136.050 604.050 ;
        RECT 139.950 601.950 142.050 604.050 ;
        RECT 131.400 599.400 132.600 601.650 ;
        RECT 140.400 600.000 141.600 601.650 ;
        RECT 121.950 595.950 124.050 598.050 ;
        RECT 103.950 586.950 106.050 589.050 ;
        RECT 109.950 586.950 112.050 589.050 ;
        RECT 103.950 580.950 106.050 583.050 ;
        RECT 92.400 571.350 93.600 573.600 ;
        RECT 98.400 571.350 99.600 573.600 ;
        RECT 100.950 571.950 103.050 574.050 ;
        RECT 88.950 568.950 91.050 571.050 ;
        RECT 91.950 568.950 94.050 571.050 ;
        RECT 94.950 568.950 97.050 571.050 ;
        RECT 97.950 568.950 100.050 571.050 ;
        RECT 89.400 567.900 90.600 568.650 ;
        RECT 88.950 565.800 91.050 567.900 ;
        RECT 95.400 566.400 96.600 568.650 ;
        RECT 95.400 565.050 96.450 566.400 ;
        RECT 104.400 565.050 105.450 580.950 ;
        RECT 106.950 577.950 109.050 580.050 ;
        RECT 107.400 574.050 108.450 577.950 ;
        RECT 106.950 571.950 109.050 574.050 ;
        RECT 110.400 573.600 111.450 586.950 ;
        RECT 115.950 577.950 118.050 580.050 ;
        RECT 116.400 573.600 117.450 577.950 ;
        RECT 122.400 574.050 123.450 595.950 ;
        RECT 131.400 583.050 132.450 599.400 ;
        RECT 139.950 595.950 142.050 600.000 ;
        RECT 146.250 593.700 147.450 606.600 ;
        RECT 145.350 591.600 147.450 593.700 ;
        RECT 130.950 580.950 133.050 583.050 ;
        RECT 149.400 580.050 150.450 637.950 ;
        RECT 170.250 635.700 171.450 642.300 ;
        RECT 169.350 633.600 171.450 635.700 ;
        RECT 166.950 616.950 169.050 619.050 ;
        RECT 160.650 613.500 162.750 614.400 ;
        RECT 160.650 612.300 164.850 613.500 ;
        RECT 157.950 605.100 160.050 607.200 ;
        RECT 158.400 604.350 159.600 605.100 ;
        RECT 151.950 601.950 154.050 604.050 ;
        RECT 157.800 601.950 159.900 604.050 ;
        RECT 152.400 595.050 153.450 601.950 ;
        RECT 154.950 598.950 157.050 601.050 ;
        RECT 151.950 592.950 154.050 595.050 ;
        RECT 124.950 577.950 127.050 580.050 ;
        RECT 148.950 577.950 151.050 580.050 ;
        RECT 110.400 571.350 111.600 573.600 ;
        RECT 116.400 571.350 117.600 573.600 ;
        RECT 121.950 571.950 124.050 574.050 ;
        RECT 109.950 568.950 112.050 571.050 ;
        RECT 112.950 568.950 115.050 571.050 ;
        RECT 115.950 568.950 118.050 571.050 ;
        RECT 118.950 568.950 121.050 571.050 ;
        RECT 106.950 565.950 109.050 568.050 ;
        RECT 113.400 567.000 114.600 568.650 ;
        RECT 119.400 567.000 120.600 568.650 ;
        RECT 125.400 567.900 126.450 577.950 ;
        RECT 155.400 576.450 156.450 598.950 ;
        RECT 163.650 593.700 164.850 612.300 ;
        RECT 167.400 606.600 168.450 616.950 ;
        RECT 167.400 604.350 168.600 606.600 ;
        RECT 166.950 601.950 169.050 604.050 ;
        RECT 163.050 591.600 165.150 593.700 ;
        RECT 157.950 577.950 160.050 580.050 ;
        RECT 167.850 579.300 169.950 581.400 ;
        RECT 152.400 575.400 156.450 576.450 ;
        RECT 133.950 572.100 136.050 574.200 ;
        RECT 134.400 571.350 135.600 572.100 ;
        RECT 142.950 571.950 145.050 574.050 ;
        RECT 152.400 573.600 153.450 575.400 ;
        RECT 158.400 573.600 159.450 577.950 ;
        RECT 130.950 568.950 133.050 571.050 ;
        RECT 133.950 568.950 136.050 571.050 ;
        RECT 136.950 568.950 139.050 571.050 ;
        RECT 94.950 559.950 97.050 565.050 ;
        RECT 103.950 562.950 106.050 565.050 ;
        RECT 85.950 538.950 88.050 541.050 ;
        RECT 103.950 538.950 106.050 541.050 ;
        RECT 86.400 531.450 87.450 538.950 ;
        RECT 91.650 535.500 93.750 536.400 ;
        RECT 91.650 534.300 95.850 535.500 ;
        RECT 86.400 530.400 90.450 531.450 ;
        RECT 89.400 528.600 90.450 530.400 ;
        RECT 89.400 526.350 90.600 528.600 ;
        RECT 88.800 523.950 90.900 526.050 ;
        RECT 94.650 515.700 95.850 534.300 ;
        RECT 97.950 528.000 100.050 532.050 ;
        RECT 98.400 526.350 99.600 528.000 ;
        RECT 97.950 523.950 100.050 526.050 ;
        RECT 104.400 522.900 105.450 538.950 ;
        RECT 107.400 538.050 108.450 565.950 ;
        RECT 112.950 562.950 115.050 567.000 ;
        RECT 118.950 562.950 121.050 567.000 ;
        RECT 124.950 565.800 127.050 567.900 ;
        RECT 127.950 565.950 130.050 568.050 ;
        RECT 131.400 567.900 132.600 568.650 ;
        RECT 128.400 562.050 129.450 565.950 ;
        RECT 130.950 565.800 133.050 567.900 ;
        RECT 137.400 566.400 138.600 568.650 ;
        RECT 143.400 567.900 144.450 571.950 ;
        RECT 152.400 571.350 153.600 573.600 ;
        RECT 158.400 571.350 159.600 573.600 ;
        RECT 148.950 568.950 151.050 571.050 ;
        RECT 151.950 568.950 154.050 571.050 ;
        RECT 154.950 568.950 157.050 571.050 ;
        RECT 157.950 568.950 160.050 571.050 ;
        RECT 163.950 568.950 166.050 571.050 ;
        RECT 149.400 567.900 150.600 568.650 ;
        RECT 133.950 562.950 136.050 565.050 ;
        RECT 127.950 559.950 130.050 562.050 ;
        RECT 106.950 535.950 109.050 538.050 ;
        RECT 115.950 527.100 118.050 529.200 ;
        RECT 121.950 527.100 124.050 529.200 ;
        RECT 127.950 527.100 130.050 529.200 ;
        RECT 134.400 528.600 135.450 562.950 ;
        RECT 137.400 562.050 138.450 566.400 ;
        RECT 142.950 565.800 145.050 567.900 ;
        RECT 148.950 565.800 151.050 567.900 ;
        RECT 155.400 566.400 156.600 568.650 ;
        RECT 164.400 566.400 165.600 568.650 ;
        RECT 136.950 559.950 139.050 562.050 ;
        RECT 155.400 556.050 156.450 566.400 ;
        RECT 154.950 553.950 157.050 556.050 ;
        RECT 154.950 547.950 157.050 550.050 ;
        RECT 151.950 538.950 154.050 541.050 ;
        RECT 148.950 535.950 151.050 538.050 ;
        RECT 139.950 532.950 142.050 535.050 ;
        RECT 140.400 528.600 141.450 532.950 ;
        RECT 116.400 526.350 117.600 527.100 ;
        RECT 122.400 526.350 123.600 527.100 ;
        RECT 112.950 523.950 115.050 526.050 ;
        RECT 115.950 523.950 118.050 526.050 ;
        RECT 118.950 523.950 121.050 526.050 ;
        RECT 121.950 523.950 124.050 526.050 ;
        RECT 103.950 520.800 106.050 522.900 ;
        RECT 113.400 521.400 114.600 523.650 ;
        RECT 119.400 522.900 120.600 523.650 ;
        RECT 113.400 517.050 114.450 521.400 ;
        RECT 118.950 520.800 121.050 522.900 ;
        RECT 94.050 513.600 96.150 515.700 ;
        RECT 112.950 514.950 115.050 517.050 ;
        RECT 118.950 514.950 121.050 517.050 ;
        RECT 106.950 505.950 109.050 508.050 ;
        RECT 88.950 502.950 91.050 505.050 ;
        RECT 89.400 496.050 90.450 502.950 ;
        RECT 83.400 494.400 87.450 495.450 ;
        RECT 70.950 490.950 73.050 493.050 ;
        RECT 73.950 490.950 76.050 493.050 ;
        RECT 76.950 490.950 79.050 493.050 ;
        RECT 79.950 490.950 82.050 493.050 ;
        RECT 74.400 489.900 75.600 490.650 ;
        RECT 80.400 489.900 81.600 490.650 ;
        RECT 73.950 487.800 76.050 489.900 ;
        RECT 79.950 487.800 82.050 489.900 ;
        RECT 55.950 466.950 58.050 469.050 ;
        RECT 64.950 466.950 67.050 469.050 ;
        RECT 23.400 461.400 27.450 462.450 ;
        RECT 23.400 454.050 24.450 461.400 ;
        RECT 44.550 459.300 46.650 461.400 ;
        RECT 29.250 457.500 31.350 458.400 ;
        RECT 27.150 456.300 31.350 457.500 ;
        RECT 22.950 451.950 25.050 454.050 ;
        RECT 19.950 448.950 22.050 451.050 ;
        RECT 23.400 450.600 24.450 451.950 ;
        RECT 23.400 448.350 24.600 450.600 ;
        RECT 11.100 445.950 13.200 448.050 ;
        RECT 16.500 445.950 18.600 448.050 ;
        RECT 22.950 445.950 25.050 448.050 ;
        RECT 17.400 444.900 18.600 445.650 ;
        RECT 16.950 442.800 19.050 444.900 ;
        RECT 27.150 437.700 28.350 456.300 ;
        RECT 40.950 451.950 43.050 454.050 ;
        RECT 44.550 452.700 45.750 459.300 ;
        RECT 31.950 449.100 34.050 451.200 ;
        RECT 32.400 448.350 33.600 449.100 ;
        RECT 32.100 445.950 34.200 448.050 ;
        RECT 26.850 435.600 28.950 437.700 ;
        RECT 31.950 430.950 34.050 433.050 ;
        RECT 7.950 427.950 10.050 430.050 ;
        RECT 19.950 427.950 22.050 430.050 ;
        RECT 8.850 423.300 10.950 425.400 ;
        RECT 4.950 418.950 7.050 421.050 ;
        RECT 1.950 415.950 4.050 418.050 ;
        RECT 4.950 412.950 7.050 415.050 ;
        RECT 1.950 409.950 4.050 412.050 ;
        RECT 5.400 410.400 6.600 412.650 ;
        RECT 2.400 286.050 3.450 409.950 ;
        RECT 5.400 403.050 6.450 410.400 ;
        RECT 9.150 404.700 10.350 423.300 ;
        RECT 14.100 412.950 16.200 415.050 ;
        RECT 9.150 403.500 13.350 404.700 ;
        RECT 4.950 400.950 7.050 403.050 ;
        RECT 11.250 402.600 13.350 403.500 ;
        RECT 20.400 376.050 21.450 427.950 ;
        RECT 26.550 423.300 28.650 425.400 ;
        RECT 22.950 418.950 25.050 421.050 ;
        RECT 23.400 388.050 24.450 418.950 ;
        RECT 26.550 410.400 27.750 423.300 ;
        RECT 32.400 417.600 33.450 430.950 ;
        RECT 32.400 415.350 33.600 417.600 ;
        RECT 31.950 412.950 34.050 415.050 ;
        RECT 26.550 408.300 28.650 410.400 ;
        RECT 26.550 401.700 27.750 408.300 ;
        RECT 41.400 403.050 42.450 451.950 ;
        RECT 44.550 450.600 46.650 452.700 ;
        RECT 44.550 437.700 45.750 450.600 ;
        RECT 49.950 445.950 52.050 448.050 ;
        RECT 50.400 444.900 51.600 445.650 ;
        RECT 49.950 442.800 52.050 444.900 ;
        RECT 44.550 435.600 46.650 437.700 ;
        RECT 50.400 420.450 51.450 442.800 ;
        RECT 56.400 435.450 57.450 466.950 ;
        RECT 86.400 460.050 87.450 494.400 ;
        RECT 88.950 493.950 91.050 496.050 ;
        RECT 94.950 495.000 97.050 499.050 ;
        RECT 95.400 493.350 96.600 495.000 ;
        RECT 100.950 494.100 103.050 499.050 ;
        RECT 107.400 495.600 108.450 505.950 ;
        RECT 91.950 490.950 94.050 493.050 ;
        RECT 94.950 490.950 97.050 493.050 ;
        RECT 92.400 489.900 93.600 490.650 ;
        RECT 91.950 487.800 94.050 489.900 ;
        RECT 73.950 457.950 76.050 460.050 ;
        RECT 85.950 457.950 88.050 460.050 ;
        RECT 58.950 448.950 61.050 451.050 ;
        RECT 67.950 449.100 70.050 451.200 ;
        RECT 59.400 439.050 60.450 448.950 ;
        RECT 68.400 448.350 69.600 449.100 ;
        RECT 64.950 445.950 67.050 448.050 ;
        RECT 67.950 445.950 70.050 448.050 ;
        RECT 65.400 444.900 66.600 445.650 ;
        RECT 64.950 442.800 67.050 444.900 ;
        RECT 58.950 436.950 61.050 439.050 ;
        RECT 56.400 434.400 60.450 435.450 ;
        RECT 47.400 419.400 51.450 420.450 ;
        RECT 47.400 417.600 48.450 419.400 ;
        RECT 47.400 415.350 48.600 417.600 ;
        RECT 52.950 416.100 55.050 418.200 ;
        RECT 53.400 415.350 54.600 416.100 ;
        RECT 46.950 412.950 49.050 415.050 ;
        RECT 49.950 412.950 52.050 415.050 ;
        RECT 52.950 412.950 55.050 415.050 ;
        RECT 50.400 411.900 51.600 412.650 ;
        RECT 59.400 412.050 60.450 434.400 ;
        RECT 74.400 421.050 75.450 457.950 ;
        RECT 101.400 457.050 102.450 494.100 ;
        RECT 107.400 493.350 108.600 495.600 ;
        RECT 112.950 494.100 115.050 496.200 ;
        RECT 113.400 493.350 114.600 494.100 ;
        RECT 106.950 490.950 109.050 493.050 ;
        RECT 109.950 490.950 112.050 493.050 ;
        RECT 112.950 490.950 115.050 493.050 ;
        RECT 110.400 489.000 111.600 490.650 ;
        RECT 109.950 484.950 112.050 489.000 ;
        RECT 119.400 481.050 120.450 514.950 ;
        RECT 128.400 508.050 129.450 527.100 ;
        RECT 134.400 526.350 135.600 528.600 ;
        RECT 140.400 526.350 141.600 528.600 ;
        RECT 133.950 523.950 136.050 526.050 ;
        RECT 136.950 523.950 139.050 526.050 ;
        RECT 139.950 523.950 142.050 526.050 ;
        RECT 142.950 523.950 145.050 526.050 ;
        RECT 137.400 521.400 138.600 523.650 ;
        RECT 143.400 522.900 144.600 523.650 ;
        RECT 137.400 517.050 138.450 521.400 ;
        RECT 142.950 520.800 145.050 522.900 ;
        RECT 136.950 514.950 139.050 517.050 ;
        RECT 130.950 508.950 133.050 511.050 ;
        RECT 127.950 505.950 130.050 508.050 ;
        RECT 131.400 501.450 132.450 508.950 ;
        RECT 142.950 502.950 145.050 505.050 ;
        RECT 127.800 498.300 129.900 500.400 ;
        RECT 131.400 499.200 132.600 501.450 ;
        RECT 125.400 495.450 126.600 495.600 ;
        RECT 122.400 494.400 126.600 495.450 ;
        RECT 122.400 487.050 123.450 494.400 ;
        RECT 125.400 493.350 126.600 494.400 ;
        RECT 125.100 490.950 127.200 493.050 ;
        RECT 128.100 492.900 129.000 498.300 ;
        RECT 131.100 496.800 133.200 498.900 ;
        RECT 135.000 495.900 137.100 497.700 ;
        RECT 129.900 494.700 138.600 495.900 ;
        RECT 129.900 493.800 132.000 494.700 ;
        RECT 128.100 491.700 135.000 492.900 ;
        RECT 121.950 484.950 124.050 487.050 ;
        RECT 128.100 484.500 129.300 491.700 ;
        RECT 131.100 487.950 133.200 490.050 ;
        RECT 134.100 489.300 135.000 491.700 ;
        RECT 131.400 485.400 132.600 487.650 ;
        RECT 134.100 487.200 136.200 489.300 ;
        RECT 137.700 485.700 138.600 494.700 ;
        RECT 139.800 490.950 141.900 493.050 ;
        RECT 140.400 489.450 141.600 490.650 ;
        RECT 143.400 489.450 144.450 502.950 ;
        RECT 145.950 499.950 148.050 502.050 ;
        RECT 146.400 490.050 147.450 499.950 ;
        RECT 149.400 496.050 150.450 535.950 ;
        RECT 152.400 529.050 153.450 538.950 ;
        RECT 151.950 526.950 154.050 529.050 ;
        RECT 155.400 528.600 156.450 547.950 ;
        RECT 160.950 535.950 163.050 538.050 ;
        RECT 161.400 528.600 162.450 535.950 ;
        RECT 164.400 532.050 165.450 566.400 ;
        RECT 168.150 560.700 169.350 579.300 ;
        RECT 173.400 577.050 174.450 667.950 ;
        RECT 191.400 667.050 192.450 685.950 ;
        RECT 200.400 684.600 201.450 718.950 ;
        RECT 203.400 709.050 204.450 722.400 ;
        RECT 209.400 715.050 210.450 766.950 ;
        RECT 212.400 756.900 213.450 769.950 ;
        RECT 215.550 764.700 216.750 771.300 ;
        RECT 262.950 769.950 265.050 772.050 ;
        RECT 229.950 766.950 232.050 769.050 ;
        RECT 241.950 766.950 244.050 769.050 ;
        RECT 215.550 762.600 217.650 764.700 ;
        RECT 211.950 754.800 214.050 756.900 ;
        RECT 211.950 748.950 214.050 751.050 ;
        RECT 215.550 749.700 216.750 762.600 ;
        RECT 226.950 761.100 229.050 763.200 ;
        RECT 220.950 757.950 223.050 760.050 ;
        RECT 221.400 756.900 222.600 757.650 ;
        RECT 227.400 757.050 228.450 761.100 ;
        RECT 220.950 754.800 223.050 756.900 ;
        RECT 226.950 754.950 229.050 757.050 ;
        RECT 230.400 756.450 231.450 766.950 ;
        RECT 235.950 761.100 238.050 763.200 ;
        RECT 242.400 762.600 243.450 766.950 ;
        RECT 247.950 763.200 250.050 766.050 ;
        RECT 236.400 760.350 237.600 761.100 ;
        RECT 242.400 760.350 243.600 762.600 ;
        RECT 247.800 762.000 250.050 763.200 ;
        RECT 247.800 761.100 249.900 762.000 ;
        RECT 250.950 761.100 253.050 763.200 ;
        RECT 256.950 761.100 259.050 763.200 ;
        RECT 263.400 762.600 264.450 769.950 ;
        RECT 235.950 757.950 238.050 760.050 ;
        RECT 238.950 757.950 241.050 760.050 ;
        RECT 241.950 757.950 244.050 760.050 ;
        RECT 244.950 757.950 247.050 760.050 ;
        RECT 239.400 756.900 240.600 757.650 ;
        RECT 245.400 756.900 246.600 757.650 ;
        RECT 230.400 755.400 234.450 756.450 ;
        RECT 212.400 742.050 213.450 748.950 ;
        RECT 215.550 747.600 217.650 749.700 ;
        RECT 214.950 742.950 217.050 745.050 ;
        RECT 211.950 739.950 214.050 742.050 ;
        RECT 212.400 730.050 213.450 739.950 ;
        RECT 215.400 730.200 216.450 742.950 ;
        RECT 223.950 733.950 226.050 736.050 ;
        RECT 211.950 727.950 214.050 730.050 ;
        RECT 214.950 728.100 217.050 730.200 ;
        RECT 215.400 727.350 216.600 728.100 ;
        RECT 214.950 724.950 217.050 727.050 ;
        RECT 217.950 724.950 220.050 727.050 ;
        RECT 218.400 723.000 219.600 724.650 ;
        RECT 217.950 718.950 220.050 723.000 ;
        RECT 220.950 721.950 223.050 724.050 ;
        RECT 208.950 712.950 211.050 715.050 ;
        RECT 202.950 706.950 205.050 709.050 ;
        RECT 208.950 706.950 211.050 709.050 ;
        RECT 200.400 682.350 201.600 684.600 ;
        RECT 200.100 679.950 202.200 682.050 ;
        RECT 205.500 679.950 207.600 682.050 ;
        RECT 206.400 677.400 207.600 679.650 ;
        RECT 199.950 673.950 202.050 676.050 ;
        RECT 190.950 664.950 193.050 667.050 ;
        RECT 175.950 655.950 178.050 658.050 ;
        RECT 187.050 657.300 189.150 659.400 ;
        RECT 176.400 646.050 177.450 655.950 ;
        RECT 181.800 646.950 183.900 649.050 ;
        RECT 175.950 643.950 178.050 646.050 ;
        RECT 182.400 645.900 183.600 646.650 ;
        RECT 181.950 643.800 184.050 645.900 ;
        RECT 187.650 638.700 188.850 657.300 ;
        RECT 196.950 649.950 199.050 652.050 ;
        RECT 190.950 646.950 193.050 649.050 ;
        RECT 184.650 637.500 188.850 638.700 ;
        RECT 191.400 644.400 192.600 646.650 ;
        RECT 184.650 636.600 186.750 637.500 ;
        RECT 191.400 619.050 192.450 644.400 ;
        RECT 193.950 643.950 196.050 646.050 ;
        RECT 194.400 640.050 195.450 643.950 ;
        RECT 197.400 643.050 198.450 649.950 ;
        RECT 196.950 640.950 199.050 643.050 ;
        RECT 193.950 637.950 196.050 640.050 ;
        RECT 190.950 616.950 193.050 619.050 ;
        RECT 196.350 615.300 198.450 617.400 ;
        RECT 184.950 610.950 187.050 613.050 ;
        RECT 185.400 606.600 186.450 610.950 ;
        RECT 197.250 608.700 198.450 615.300 ;
        RECT 196.350 606.600 198.450 608.700 ;
        RECT 200.400 609.450 201.450 673.950 ;
        RECT 206.400 667.050 207.450 677.400 ;
        RECT 205.950 664.950 208.050 667.050 ;
        RECT 209.400 661.050 210.450 706.950 ;
        RECT 221.400 703.050 222.450 721.950 ;
        RECT 220.950 700.950 223.050 703.050 ;
        RECT 211.950 685.950 214.050 688.050 ;
        RECT 212.400 678.900 213.450 685.950 ;
        RECT 217.950 683.100 220.050 685.200 ;
        RECT 224.400 685.050 225.450 733.950 ;
        RECT 233.400 729.600 234.450 755.400 ;
        RECT 238.950 754.800 241.050 756.900 ;
        RECT 244.950 754.800 247.050 756.900 ;
        RECT 247.950 751.950 250.050 754.050 ;
        RECT 248.400 745.050 249.450 751.950 ;
        RECT 251.400 751.050 252.450 761.100 ;
        RECT 257.400 760.350 258.600 761.100 ;
        RECT 263.400 760.350 264.600 762.600 ;
        RECT 256.950 757.950 259.050 760.050 ;
        RECT 259.950 757.950 262.050 760.050 ;
        RECT 262.950 757.950 265.050 760.050 ;
        RECT 253.950 751.950 256.050 757.050 ;
        RECT 260.400 756.900 261.600 757.650 ;
        RECT 259.950 754.800 262.050 756.900 ;
        RECT 250.950 748.950 253.050 751.050 ;
        RECT 247.950 742.950 250.050 745.050 ;
        RECT 251.400 742.050 252.450 748.950 ;
        RECT 250.950 739.950 253.050 742.050 ;
        RECT 238.950 733.950 241.050 736.050 ;
        RECT 250.950 733.950 253.050 736.050 ;
        RECT 239.400 729.600 240.450 733.950 ;
        RECT 251.400 729.600 252.450 733.950 ;
        RECT 233.400 727.350 234.600 729.600 ;
        RECT 239.400 727.350 240.600 729.600 ;
        RECT 251.400 727.350 252.600 729.600 ;
        RECT 256.950 728.100 259.050 730.200 ;
        RECT 257.400 727.350 258.600 728.100 ;
        RECT 265.950 727.950 268.050 730.050 ;
        RECT 229.950 724.950 232.050 727.050 ;
        RECT 232.950 724.950 235.050 727.050 ;
        RECT 235.950 724.950 238.050 727.050 ;
        RECT 238.950 724.950 241.050 727.050 ;
        RECT 250.950 724.950 253.050 727.050 ;
        RECT 253.950 724.950 256.050 727.050 ;
        RECT 256.950 724.950 259.050 727.050 ;
        RECT 259.950 724.950 262.050 727.050 ;
        RECT 230.400 723.450 231.600 724.650 ;
        RECT 227.400 722.400 231.600 723.450 ;
        RECT 236.400 723.000 237.600 724.650 ;
        RECT 254.400 723.000 255.600 724.650 ;
        RECT 260.400 723.900 261.600 724.650 ;
        RECT 259.950 723.450 262.050 723.900 ;
        RECT 227.400 709.050 228.450 722.400 ;
        RECT 235.950 718.950 238.050 723.000 ;
        RECT 253.950 718.950 256.050 723.000 ;
        RECT 259.950 722.400 264.450 723.450 ;
        RECT 259.950 721.800 262.050 722.400 ;
        RECT 244.950 712.950 247.050 715.050 ;
        RECT 253.950 712.950 256.050 715.050 ;
        RECT 226.950 706.950 229.050 709.050 ;
        RECT 218.400 682.350 219.600 683.100 ;
        RECT 223.950 682.950 226.050 685.050 ;
        RECT 217.950 679.950 220.050 682.050 ;
        RECT 220.950 679.950 223.050 682.050 ;
        RECT 221.400 678.900 222.600 679.650 ;
        RECT 211.950 676.800 214.050 678.900 ;
        RECT 220.950 676.800 223.050 678.900 ;
        RECT 227.400 670.050 228.450 706.950 ;
        RECT 235.950 683.100 238.050 685.200 ;
        RECT 236.400 682.350 237.600 683.100 ;
        RECT 241.950 682.950 244.050 688.050 ;
        RECT 232.950 679.950 235.050 682.050 ;
        RECT 235.950 679.950 238.050 682.050 ;
        RECT 238.950 679.950 241.050 682.050 ;
        RECT 229.950 676.950 232.050 679.050 ;
        RECT 233.400 678.900 234.600 679.650 ;
        RECT 239.400 679.050 240.600 679.650 ;
        RECT 230.400 673.050 231.450 676.950 ;
        RECT 232.950 676.800 235.050 678.900 ;
        RECT 239.400 677.400 244.050 679.050 ;
        RECT 240.000 676.950 244.050 677.400 ;
        RECT 229.950 670.950 232.050 673.050 ;
        RECT 220.950 667.950 223.050 670.050 ;
        RECT 226.950 667.950 229.050 670.050 ;
        RECT 208.950 658.950 211.050 661.050 ;
        RECT 208.950 655.800 211.050 657.900 ;
        RECT 209.400 651.600 210.450 655.800 ;
        RECT 209.400 649.350 210.600 651.600 ;
        RECT 214.950 650.100 217.050 652.200 ;
        RECT 215.400 649.350 216.600 650.100 ;
        RECT 205.950 646.950 208.050 649.050 ;
        RECT 208.950 646.950 211.050 649.050 ;
        RECT 211.950 646.950 214.050 649.050 ;
        RECT 214.950 646.950 217.050 649.050 ;
        RECT 206.400 645.000 207.600 646.650 ;
        RECT 205.950 640.950 208.050 645.000 ;
        RECT 212.400 644.400 213.600 646.650 ;
        RECT 212.400 634.050 213.450 644.400 ;
        RECT 221.400 640.050 222.450 667.950 ;
        RECT 232.950 664.950 235.050 667.050 ;
        RECT 233.400 651.600 234.450 664.950 ;
        RECT 238.950 658.950 241.050 661.050 ;
        RECT 233.400 651.450 234.600 651.600 ;
        RECT 233.400 650.400 237.450 651.450 ;
        RECT 233.400 649.350 234.600 650.400 ;
        RECT 227.100 646.950 229.200 649.050 ;
        RECT 232.500 646.950 234.600 649.050 ;
        RECT 227.400 645.900 228.600 646.650 ;
        RECT 226.950 643.800 229.050 645.900 ;
        RECT 220.950 637.950 223.050 640.050 ;
        RECT 226.950 637.950 229.050 640.050 ;
        RECT 205.950 631.950 208.050 634.050 ;
        RECT 211.950 631.950 214.050 634.050 ;
        RECT 206.400 610.050 207.450 631.950 ;
        RECT 217.950 616.950 220.050 619.050 ;
        RECT 211.650 613.500 213.750 614.400 ;
        RECT 211.650 612.300 215.850 613.500 ;
        RECT 200.400 608.400 204.450 609.450 ;
        RECT 185.400 604.350 186.600 606.600 ;
        RECT 181.950 601.950 184.050 604.050 ;
        RECT 184.950 601.950 187.050 604.050 ;
        RECT 190.950 601.950 193.050 604.050 ;
        RECT 182.400 599.400 183.600 601.650 ;
        RECT 191.400 599.400 192.600 601.650 ;
        RECT 182.400 595.050 183.450 599.400 ;
        RECT 191.400 595.050 192.450 599.400 ;
        RECT 181.950 592.950 184.050 595.050 ;
        RECT 190.950 592.950 193.050 595.050 ;
        RECT 197.250 593.700 198.450 606.600 ;
        RECT 199.950 604.950 202.050 607.050 ;
        RECT 196.350 591.600 198.450 593.700 ;
        RECT 200.400 589.050 201.450 604.950 ;
        RECT 181.950 586.950 184.050 589.050 ;
        RECT 199.950 586.950 202.050 589.050 ;
        RECT 172.950 574.950 175.050 577.050 ;
        RECT 178.950 571.950 181.050 574.050 ;
        RECT 173.100 568.950 175.200 571.050 ;
        RECT 173.400 567.900 174.600 568.650 ;
        RECT 179.400 567.900 180.450 571.950 ;
        RECT 172.950 565.800 175.050 567.900 ;
        RECT 178.950 565.800 181.050 567.900 ;
        RECT 168.150 559.500 172.350 560.700 ;
        RECT 170.250 558.600 172.350 559.500 ;
        RECT 182.400 553.050 183.450 586.950 ;
        RECT 185.550 579.300 187.650 581.400 ;
        RECT 193.950 580.950 196.050 583.050 ;
        RECT 185.550 566.400 186.750 579.300 ;
        RECT 190.950 577.950 193.050 580.050 ;
        RECT 191.400 573.600 192.450 577.950 ;
        RECT 194.400 574.050 195.450 580.950 ;
        RECT 191.400 571.350 192.600 573.600 ;
        RECT 193.950 571.950 196.050 574.050 ;
        RECT 196.950 571.950 199.050 574.050 ;
        RECT 199.950 572.100 202.050 574.200 ;
        RECT 203.400 574.050 204.450 608.400 ;
        RECT 205.950 607.950 208.050 610.050 ;
        RECT 208.950 605.100 211.050 607.200 ;
        RECT 209.400 604.350 210.600 605.100 ;
        RECT 208.800 601.950 210.900 604.050 ;
        RECT 214.650 593.700 215.850 612.300 ;
        RECT 218.400 606.600 219.450 616.950 ;
        RECT 218.400 604.350 219.600 606.600 ;
        RECT 217.950 601.950 220.050 604.050 ;
        RECT 227.400 601.050 228.450 637.950 ;
        RECT 236.400 637.050 237.450 650.400 ;
        RECT 239.400 643.050 240.450 658.950 ;
        RECT 238.950 640.950 241.050 643.050 ;
        RECT 235.950 634.950 238.050 637.050 ;
        RECT 245.400 631.050 246.450 712.950 ;
        RECT 254.400 684.600 255.450 712.950 ;
        RECT 256.950 700.950 259.050 703.050 ;
        RECT 257.400 685.050 258.450 700.950 ;
        RECT 259.950 685.950 262.050 688.050 ;
        RECT 254.400 682.350 255.600 684.600 ;
        RECT 256.950 682.950 259.050 685.050 ;
        RECT 260.400 682.050 261.450 685.950 ;
        RECT 263.400 685.050 264.450 722.400 ;
        RECT 266.400 721.050 267.450 727.950 ;
        RECT 265.950 718.950 268.050 721.050 ;
        RECT 269.400 709.050 270.450 784.950 ;
        RECT 277.950 761.100 280.050 763.200 ;
        RECT 287.400 763.050 288.450 800.400 ;
        RECT 295.950 799.800 298.050 801.900 ;
        RECT 302.400 774.450 303.450 805.950 ;
        RECT 314.400 805.350 315.600 807.600 ;
        RECT 322.950 805.950 325.050 808.050 ;
        RECT 328.950 806.100 331.050 808.200 ;
        RECT 308.100 802.950 310.200 805.050 ;
        RECT 313.500 802.950 315.600 805.050 ;
        RECT 316.800 802.950 318.900 805.050 ;
        RECT 308.400 801.900 309.600 802.650 ;
        RECT 307.950 799.800 310.050 801.900 ;
        RECT 317.400 800.400 318.600 802.650 ;
        RECT 317.400 796.050 318.450 800.400 ;
        RECT 316.950 793.950 319.050 796.050 ;
        RECT 307.950 778.950 310.050 781.050 ;
        RECT 302.400 773.400 306.450 774.450 ;
        RECT 298.950 769.950 301.050 772.050 ;
        RECT 299.400 766.050 300.450 769.950 ;
        RECT 301.950 766.950 304.050 769.050 ;
        RECT 298.950 763.950 301.050 766.050 ;
        RECT 278.400 760.350 279.600 761.100 ;
        RECT 286.950 760.950 289.050 763.050 ;
        RECT 295.950 761.100 298.050 763.200 ;
        RECT 296.400 760.350 297.600 761.100 ;
        RECT 274.950 757.950 277.050 760.050 ;
        RECT 277.950 757.950 280.050 760.050 ;
        RECT 280.950 757.950 283.050 760.050 ;
        RECT 286.950 757.800 289.050 759.900 ;
        RECT 292.950 757.950 295.050 760.050 ;
        RECT 295.950 757.950 298.050 760.050 ;
        RECT 275.400 756.000 276.600 757.650 ;
        RECT 281.400 757.050 282.600 757.650 ;
        RECT 274.950 751.950 277.050 756.000 ;
        RECT 281.400 755.400 286.050 757.050 ;
        RECT 282.000 754.950 286.050 755.400 ;
        RECT 287.400 733.050 288.450 757.800 ;
        RECT 293.400 757.050 294.600 757.650 ;
        RECT 289.950 755.400 294.600 757.050 ;
        RECT 289.950 754.950 294.000 755.400 ;
        RECT 289.950 736.950 292.050 739.050 ;
        RECT 274.950 729.000 277.050 733.050 ;
        RECT 286.950 730.950 289.050 733.050 ;
        RECT 281.400 729.450 282.600 729.600 ;
        RECT 275.400 727.350 276.600 729.000 ;
        RECT 281.400 728.400 288.450 729.450 ;
        RECT 281.400 727.350 282.600 728.400 ;
        RECT 274.950 724.950 277.050 727.050 ;
        RECT 277.950 724.950 280.050 727.050 ;
        RECT 280.950 724.950 283.050 727.050 ;
        RECT 278.400 722.400 279.600 724.650 ;
        RECT 268.950 706.950 271.050 709.050 ;
        RECT 262.950 682.950 265.050 685.050 ;
        RECT 268.950 683.100 271.050 688.050 ;
        RECT 274.950 684.000 277.050 688.050 ;
        RECT 278.400 684.450 279.450 722.400 ;
        RECT 287.400 715.050 288.450 728.400 ;
        RECT 290.400 727.050 291.450 736.950 ;
        RECT 302.400 735.450 303.450 766.950 ;
        RECT 305.400 739.050 306.450 773.400 ;
        RECT 308.400 739.050 309.450 778.950 ;
        RECT 311.100 757.950 313.200 760.050 ;
        RECT 316.500 757.950 318.600 760.050 ;
        RECT 317.400 756.900 318.600 757.650 ;
        RECT 316.950 754.800 319.050 756.900 ;
        RECT 304.800 736.950 306.900 739.050 ;
        RECT 307.950 736.950 310.050 739.050 ;
        RECT 313.950 736.950 316.050 739.050 ;
        RECT 302.400 733.200 303.600 735.450 ;
        RECT 297.900 729.900 300.000 731.700 ;
        RECT 301.800 730.800 303.900 732.900 ;
        RECT 305.100 732.300 307.200 734.400 ;
        RECT 296.400 728.700 305.100 729.900 ;
        RECT 289.950 724.950 292.050 727.050 ;
        RECT 293.100 724.950 295.200 727.050 ;
        RECT 293.400 723.450 294.600 724.650 ;
        RECT 290.400 723.000 294.600 723.450 ;
        RECT 289.950 722.400 294.600 723.000 ;
        RECT 289.950 718.950 292.050 722.400 ;
        RECT 296.400 719.700 297.300 728.700 ;
        RECT 303.000 727.800 305.100 728.700 ;
        RECT 306.000 726.900 306.900 732.300 ;
        RECT 308.400 729.450 309.600 729.600 ;
        RECT 308.400 728.400 312.450 729.450 ;
        RECT 308.400 727.350 309.600 728.400 ;
        RECT 300.000 725.700 306.900 726.900 ;
        RECT 300.000 723.300 300.900 725.700 ;
        RECT 298.800 721.200 300.900 723.300 ;
        RECT 301.800 721.950 303.900 724.050 ;
        RECT 295.500 717.600 297.600 719.700 ;
        RECT 302.400 719.400 303.600 721.650 ;
        RECT 305.700 718.500 306.900 725.700 ;
        RECT 307.800 724.950 309.900 727.050 ;
        RECT 305.100 716.400 307.200 718.500 ;
        RECT 311.400 715.050 312.450 728.400 ;
        RECT 286.950 712.950 289.050 715.050 ;
        RECT 310.950 712.950 313.050 715.050 ;
        RECT 307.950 703.950 310.050 706.050 ;
        RECT 301.950 688.950 304.050 691.050 ;
        RECT 298.950 685.950 301.050 688.050 ;
        RECT 269.400 682.350 270.600 683.100 ;
        RECT 275.400 682.350 276.600 684.000 ;
        RECT 278.400 683.400 282.450 684.450 ;
        RECT 250.950 679.950 253.050 682.050 ;
        RECT 253.950 679.950 256.050 682.050 ;
        RECT 259.950 679.950 262.050 682.050 ;
        RECT 265.950 679.950 268.050 682.050 ;
        RECT 268.950 679.950 271.050 682.050 ;
        RECT 271.950 679.950 274.050 682.050 ;
        RECT 274.950 679.950 277.050 682.050 ;
        RECT 251.400 679.050 252.600 679.650 ;
        RECT 247.950 677.400 252.600 679.050 ;
        RECT 266.400 678.900 267.600 679.650 ;
        RECT 247.950 676.950 252.000 677.400 ;
        RECT 259.950 676.800 262.050 678.900 ;
        RECT 265.950 676.800 268.050 678.900 ;
        RECT 272.400 677.400 273.600 679.650 ;
        RECT 253.950 670.950 256.050 673.050 ;
        RECT 248.100 646.950 250.200 649.050 ;
        RECT 248.400 644.400 249.600 646.650 ;
        RECT 244.950 628.950 247.050 631.050 ;
        RECT 248.400 619.050 249.450 644.400 ;
        RECT 254.400 625.050 255.450 670.950 ;
        RECT 260.400 634.050 261.450 676.800 ;
        RECT 266.100 646.950 268.200 649.050 ;
        RECT 272.400 643.050 273.450 677.400 ;
        RECT 281.400 654.450 282.450 683.400 ;
        RECT 289.950 683.100 292.050 685.200 ;
        RECT 290.400 682.350 291.600 683.100 ;
        RECT 286.950 679.950 289.050 682.050 ;
        RECT 289.950 679.950 292.050 682.050 ;
        RECT 292.950 679.950 295.050 682.050 ;
        RECT 287.400 677.400 288.600 679.650 ;
        RECT 293.400 678.900 294.600 679.650 ;
        RECT 299.400 679.050 300.450 685.950 ;
        RECT 287.400 655.050 288.450 677.400 ;
        RECT 292.950 676.800 295.050 678.900 ;
        RECT 298.950 676.950 301.050 679.050 ;
        RECT 289.950 670.950 292.050 673.050 ;
        RECT 281.400 653.400 285.450 654.450 ;
        RECT 284.400 651.600 285.450 653.400 ;
        RECT 286.950 652.950 289.050 655.050 ;
        RECT 290.400 651.600 291.450 670.950 ;
        RECT 302.400 655.050 303.450 688.950 ;
        RECT 308.400 685.200 309.450 703.950 ;
        RECT 314.400 697.050 315.450 736.950 ;
        RECT 323.400 729.600 324.450 805.950 ;
        RECT 329.400 805.350 330.600 806.100 ;
        RECT 329.400 802.950 331.500 805.050 ;
        RECT 334.800 802.950 336.900 805.050 ;
        RECT 340.950 802.950 343.050 805.050 ;
        RECT 341.400 800.400 342.600 802.650 ;
        RECT 328.950 781.950 331.050 784.050 ;
        RECT 329.400 762.600 330.450 781.950 ;
        RECT 341.400 781.050 342.450 800.400 ;
        RECT 345.150 794.700 346.350 813.300 ;
        RECT 350.100 802.950 352.200 805.050 ;
        RECT 350.400 801.900 351.600 802.650 ;
        RECT 349.950 799.800 352.050 801.900 ;
        RECT 362.550 800.400 363.750 813.300 ;
        RECT 385.950 812.400 394.050 813.450 ;
        RECT 385.950 811.950 388.050 812.400 ;
        RECT 391.950 811.950 394.050 812.400 ;
        RECT 395.400 811.050 396.450 814.950 ;
        RECT 367.950 806.100 370.050 808.200 ;
        RECT 382.950 806.100 385.050 808.200 ;
        RECT 388.950 807.000 391.050 811.050 ;
        RECT 394.950 808.950 397.050 811.050 ;
        RECT 406.950 808.950 409.050 814.050 ;
        RECT 368.400 805.350 369.600 806.100 ;
        RECT 383.400 805.350 384.600 806.100 ;
        RECT 389.400 805.350 390.600 807.000 ;
        RECT 367.950 802.950 370.050 805.050 ;
        RECT 382.950 802.950 385.050 805.050 ;
        RECT 385.950 802.950 388.050 805.050 ;
        RECT 388.950 802.950 391.050 805.050 ;
        RECT 386.400 801.900 387.600 802.650 ;
        RECT 362.550 798.300 364.650 800.400 ;
        RECT 385.950 799.800 388.050 801.900 ;
        RECT 345.150 793.500 349.350 794.700 ;
        RECT 347.250 792.600 349.350 793.500 ;
        RECT 362.550 791.700 363.750 798.300 ;
        RECT 395.400 796.050 396.450 808.950 ;
        RECT 403.950 806.100 406.050 808.200 ;
        RECT 410.400 807.600 411.450 814.950 ;
        RECT 418.950 808.950 421.050 811.050 ;
        RECT 421.950 808.950 424.050 814.050 ;
        RECT 440.850 813.300 442.950 815.400 ;
        RECT 404.400 805.350 405.600 806.100 ;
        RECT 410.400 805.350 411.600 807.600 ;
        RECT 403.950 802.950 406.050 805.050 ;
        RECT 406.950 802.950 409.050 805.050 ;
        RECT 409.950 802.950 412.050 805.050 ;
        RECT 412.950 802.950 415.050 805.050 ;
        RECT 407.400 801.900 408.600 802.650 ;
        RECT 413.400 801.900 414.600 802.650 ;
        RECT 406.950 799.800 409.050 801.900 ;
        RECT 412.950 799.800 415.050 801.900 ;
        RECT 373.950 793.950 376.050 796.050 ;
        RECT 394.950 793.950 397.050 796.050 ;
        RECT 400.950 793.950 403.050 796.050 ;
        RECT 362.550 789.600 364.650 791.700 ;
        RECT 340.950 778.950 343.050 781.050 ;
        RECT 364.950 769.950 367.050 772.050 ;
        RECT 352.950 768.450 355.050 769.050 ;
        RECT 358.950 768.450 361.050 769.050 ;
        RECT 352.950 767.400 361.050 768.450 ;
        RECT 352.950 766.950 355.050 767.400 ;
        RECT 358.950 766.950 361.050 767.400 ;
        RECT 329.400 760.350 330.600 762.600 ;
        RECT 334.950 761.100 337.050 763.200 ;
        RECT 343.950 761.100 346.050 763.200 ;
        RECT 349.950 761.100 352.050 763.200 ;
        RECT 355.950 762.000 358.050 766.050 ;
        RECT 335.400 760.350 336.600 761.100 ;
        RECT 328.950 757.950 331.050 760.050 ;
        RECT 331.950 757.950 334.050 760.050 ;
        RECT 334.950 757.950 337.050 760.050 ;
        RECT 337.950 757.950 340.050 760.050 ;
        RECT 332.400 756.900 333.600 757.650 ;
        RECT 331.950 754.800 334.050 756.900 ;
        RECT 338.400 755.400 339.600 757.650 ;
        RECT 338.400 751.050 339.450 755.400 ;
        RECT 337.950 748.950 340.050 751.050 ;
        RECT 328.950 736.950 331.050 739.050 ;
        RECT 334.950 736.950 337.050 739.050 ;
        RECT 329.400 729.600 330.450 736.950 ;
        RECT 323.400 727.350 324.600 729.600 ;
        RECT 329.400 727.350 330.600 729.600 ;
        RECT 319.950 724.950 322.050 727.050 ;
        RECT 322.950 724.950 325.050 727.050 ;
        RECT 325.950 724.950 328.050 727.050 ;
        RECT 328.950 724.950 331.050 727.050 ;
        RECT 320.400 722.400 321.600 724.650 ;
        RECT 326.400 722.400 327.600 724.650 ;
        RECT 335.400 723.900 336.450 736.950 ;
        RECT 344.400 730.200 345.450 761.100 ;
        RECT 350.400 760.350 351.600 761.100 ;
        RECT 356.400 760.350 357.600 762.000 ;
        RECT 349.950 757.950 352.050 760.050 ;
        RECT 352.950 757.950 355.050 760.050 ;
        RECT 355.950 757.950 358.050 760.050 ;
        RECT 358.950 757.950 361.050 760.050 ;
        RECT 353.400 756.900 354.600 757.650 ;
        RECT 359.400 756.900 360.600 757.650 ;
        RECT 352.950 754.800 355.050 756.900 ;
        RECT 358.950 754.800 361.050 756.900 ;
        RECT 359.400 753.450 360.450 754.800 ;
        RECT 356.400 752.400 360.450 753.450 ;
        RECT 349.950 733.950 352.050 736.050 ;
        RECT 343.950 728.100 346.050 730.200 ;
        RECT 344.400 727.350 345.600 728.100 ;
        RECT 340.950 724.950 343.050 727.050 ;
        RECT 343.950 724.950 346.050 727.050 ;
        RECT 341.400 723.900 342.600 724.650 ;
        RECT 320.400 715.050 321.450 722.400 ;
        RECT 326.400 718.050 327.450 722.400 ;
        RECT 334.950 721.800 337.050 723.900 ;
        RECT 340.950 721.800 343.050 723.900 ;
        RECT 350.400 718.050 351.450 733.950 ;
        RECT 356.400 730.200 357.450 752.400 ;
        RECT 365.400 751.050 366.450 769.950 ;
        RECT 374.400 763.200 375.450 793.950 ;
        RECT 388.950 775.950 391.050 778.050 ;
        RECT 373.950 761.100 376.050 763.200 ;
        RECT 374.400 760.350 375.600 761.100 ;
        RECT 382.950 760.950 385.050 763.050 ;
        RECT 389.400 762.600 390.450 775.950 ;
        RECT 401.400 763.200 402.450 793.950 ;
        RECT 403.950 778.950 406.050 781.050 ;
        RECT 370.950 757.950 373.050 760.050 ;
        RECT 373.950 757.950 376.050 760.050 ;
        RECT 376.950 757.950 379.050 760.050 ;
        RECT 371.400 755.400 372.600 757.650 ;
        RECT 377.400 756.900 378.600 757.650 ;
        RECT 371.400 751.050 372.450 755.400 ;
        RECT 376.950 754.800 379.050 756.900 ;
        RECT 364.950 748.950 367.050 751.050 ;
        RECT 370.950 748.950 373.050 751.050 ;
        RECT 371.400 739.050 372.450 748.950 ;
        RECT 377.400 745.050 378.450 754.800 ;
        RECT 376.950 742.950 379.050 745.050 ;
        RECT 370.950 736.950 373.050 739.050 ;
        RECT 361.950 733.950 364.050 736.050 ;
        RECT 355.950 728.100 358.050 730.200 ;
        RECT 362.400 729.600 363.450 733.950 ;
        RECT 383.400 733.050 384.450 760.950 ;
        RECT 389.400 760.350 390.600 762.600 ;
        RECT 394.950 761.100 397.050 763.200 ;
        RECT 400.950 761.100 403.050 763.200 ;
        RECT 395.400 760.350 396.600 761.100 ;
        RECT 388.950 757.950 391.050 760.050 ;
        RECT 391.950 757.950 394.050 760.050 ;
        RECT 394.950 757.950 397.050 760.050 ;
        RECT 397.950 757.950 400.050 760.050 ;
        RECT 392.400 756.900 393.600 757.650 ;
        RECT 391.950 754.800 394.050 756.900 ;
        RECT 398.400 755.400 399.600 757.650 ;
        RECT 404.400 756.900 405.450 778.950 ;
        RECT 412.950 769.950 415.050 772.050 ;
        RECT 413.400 762.600 414.450 769.950 ;
        RECT 419.400 763.050 420.450 808.950 ;
        RECT 425.400 807.450 426.600 807.600 ;
        RECT 422.400 806.400 426.600 807.450 ;
        RECT 422.400 781.050 423.450 806.400 ;
        RECT 425.400 805.350 426.600 806.400 ;
        RECT 425.400 802.950 427.500 805.050 ;
        RECT 430.800 802.950 432.900 805.050 ;
        RECT 436.950 802.950 439.050 805.050 ;
        RECT 437.400 800.400 438.600 802.650 ;
        RECT 437.400 781.050 438.450 800.400 ;
        RECT 441.150 794.700 442.350 813.300 ;
        RECT 446.100 802.950 448.200 805.050 ;
        RECT 446.400 801.450 447.600 802.650 ;
        RECT 446.400 800.400 450.450 801.450 ;
        RECT 441.150 793.500 445.350 794.700 ;
        RECT 443.250 792.600 445.350 793.500 ;
        RECT 449.400 790.050 450.450 800.400 ;
        RECT 455.400 796.050 456.450 817.950 ;
        RECT 458.550 813.300 460.650 815.400 ;
        RECT 458.550 800.400 459.750 813.300 ;
        RECT 469.950 811.950 475.050 814.050 ;
        RECT 475.950 813.450 478.050 814.050 ;
        RECT 481.950 813.450 484.050 814.050 ;
        RECT 475.950 812.400 484.050 813.450 ;
        RECT 475.950 811.950 478.050 812.400 ;
        RECT 481.950 811.950 484.050 812.400 ;
        RECT 463.950 806.100 466.050 808.200 ;
        RECT 469.950 806.100 472.050 808.200 ;
        RECT 478.950 806.100 481.050 811.050 ;
        RECT 485.400 807.600 486.450 817.950 ;
        RECT 565.950 811.950 568.050 814.050 ;
        RECT 574.950 811.950 577.050 814.050 ;
        RECT 589.350 813.300 591.450 815.400 ;
        RECT 464.400 805.350 465.600 806.100 ;
        RECT 463.950 802.950 466.050 805.050 ;
        RECT 458.550 798.300 460.650 800.400 ;
        RECT 466.950 798.450 469.050 799.050 ;
        RECT 470.400 798.450 471.450 806.100 ;
        RECT 479.400 805.350 480.600 806.100 ;
        RECT 485.400 805.350 486.600 807.600 ;
        RECT 496.950 805.950 499.050 811.050 ;
        RECT 566.400 808.200 567.450 811.950 ;
        RECT 502.950 806.100 505.050 808.200 ;
        RECT 503.400 805.350 504.600 806.100 ;
        RECT 511.950 805.950 514.050 808.050 ;
        RECT 559.950 805.950 562.050 808.050 ;
        RECT 565.950 806.100 568.050 808.200 ;
        RECT 575.400 807.600 576.450 811.950 ;
        RECT 472.950 802.950 475.050 805.050 ;
        RECT 478.950 802.950 481.050 805.050 ;
        RECT 481.950 802.950 484.050 805.050 ;
        RECT 484.950 802.950 487.050 805.050 ;
        RECT 487.950 802.950 490.050 805.050 ;
        RECT 499.950 802.950 502.050 805.050 ;
        RECT 502.950 802.950 505.050 805.050 ;
        RECT 505.950 802.950 508.050 805.050 ;
        RECT 454.950 793.950 457.050 796.050 ;
        RECT 458.550 791.700 459.750 798.300 ;
        RECT 466.950 797.400 471.450 798.450 ;
        RECT 466.950 796.950 469.050 797.400 ;
        RECT 442.950 787.950 445.050 790.050 ;
        RECT 448.950 787.950 451.050 790.050 ;
        RECT 458.550 789.600 460.650 791.700 ;
        RECT 421.950 778.950 424.050 781.050 ;
        RECT 436.950 778.950 439.050 781.050 ;
        RECT 421.950 772.950 424.050 775.050 ;
        RECT 413.400 760.350 414.600 762.600 ;
        RECT 418.950 760.950 421.050 763.050 ;
        RECT 409.950 757.950 412.050 760.050 ;
        RECT 412.950 757.950 415.050 760.050 ;
        RECT 415.950 757.950 418.050 760.050 ;
        RECT 398.400 751.050 399.450 755.400 ;
        RECT 403.950 754.800 406.050 756.900 ;
        RECT 410.400 755.400 411.600 757.650 ;
        RECT 416.400 756.900 417.600 757.650 ;
        RECT 422.400 756.900 423.450 772.950 ;
        RECT 428.100 757.950 430.200 760.050 ;
        RECT 433.500 757.950 435.600 760.050 ;
        RECT 410.400 751.050 411.450 755.400 ;
        RECT 415.950 754.800 418.050 756.900 ;
        RECT 421.950 754.800 424.050 756.900 ;
        RECT 434.400 755.400 435.600 757.650 ;
        RECT 430.950 751.950 433.050 754.050 ;
        RECT 397.950 748.950 400.050 751.050 ;
        RECT 409.950 748.950 412.050 751.050 ;
        RECT 418.950 748.950 421.050 751.050 ;
        RECT 394.950 742.950 397.050 745.050 ;
        RECT 412.950 742.950 415.050 745.050 ;
        RECT 382.950 730.950 385.050 733.050 ;
        RECT 388.950 730.950 391.050 733.050 ;
        RECT 356.400 727.350 357.600 728.100 ;
        RECT 362.400 727.350 363.600 729.600 ;
        RECT 370.950 728.100 373.050 730.200 ;
        RECT 379.950 728.100 382.050 730.200 ;
        RECT 355.950 724.950 358.050 727.050 ;
        RECT 358.950 724.950 361.050 727.050 ;
        RECT 361.950 724.950 364.050 727.050 ;
        RECT 364.950 724.950 367.050 727.050 ;
        RECT 359.400 722.400 360.600 724.650 ;
        RECT 365.400 723.900 366.600 724.650 ;
        RECT 359.400 720.450 360.450 722.400 ;
        RECT 364.950 721.800 367.050 723.900 ;
        RECT 359.400 719.400 363.450 720.450 ;
        RECT 325.950 715.950 328.050 718.050 ;
        RECT 349.950 715.950 352.050 718.050 ;
        RECT 319.950 712.950 322.050 715.050 ;
        RECT 337.950 712.950 340.050 715.050 ;
        RECT 313.950 694.950 316.050 697.050 ;
        RECT 319.950 694.950 322.050 697.050 ;
        RECT 313.950 688.950 316.050 691.050 ;
        RECT 307.950 683.100 310.050 685.200 ;
        RECT 314.400 684.600 315.450 688.950 ;
        RECT 320.400 684.600 321.450 694.950 ;
        RECT 326.250 691.500 328.350 692.400 ;
        RECT 324.150 690.300 328.350 691.500 ;
        RECT 308.400 682.350 309.600 683.100 ;
        RECT 314.400 682.350 315.600 684.600 ;
        RECT 320.400 682.350 321.600 684.600 ;
        RECT 307.950 679.950 310.050 682.050 ;
        RECT 310.950 679.950 313.050 682.050 ;
        RECT 313.950 679.950 316.050 682.050 ;
        RECT 319.950 679.950 322.050 682.050 ;
        RECT 311.400 678.900 312.600 679.650 ;
        RECT 310.950 676.800 313.050 678.900 ;
        RECT 324.150 671.700 325.350 690.300 ;
        RECT 328.950 683.100 331.050 685.200 ;
        RECT 334.950 683.100 337.050 685.200 ;
        RECT 329.400 682.350 330.600 683.100 ;
        RECT 329.100 679.950 331.200 682.050 ;
        RECT 335.400 673.050 336.450 683.100 ;
        RECT 323.850 669.600 325.950 671.700 ;
        RECT 334.950 670.950 337.050 673.050 ;
        RECT 316.350 657.300 318.450 659.400 ;
        RECT 284.400 649.350 285.600 651.600 ;
        RECT 290.400 649.350 291.600 651.600 ;
        RECT 301.950 651.000 304.050 655.050 ;
        RECT 310.950 651.000 313.050 655.050 ;
        RECT 302.400 649.350 303.600 651.000 ;
        RECT 311.400 649.350 312.600 651.000 ;
        RECT 280.950 646.950 283.050 649.050 ;
        RECT 283.950 646.950 286.050 649.050 ;
        RECT 286.950 646.950 289.050 649.050 ;
        RECT 289.950 646.950 292.050 649.050 ;
        RECT 301.950 646.950 304.050 649.050 ;
        RECT 304.950 646.950 307.050 649.050 ;
        RECT 310.950 646.950 313.050 649.050 ;
        RECT 281.400 644.400 282.600 646.650 ;
        RECT 287.400 645.000 288.600 646.650 ;
        RECT 271.950 640.950 274.050 643.050 ;
        RECT 281.400 634.050 282.450 644.400 ;
        RECT 283.950 640.950 286.050 643.050 ;
        RECT 286.950 640.950 289.050 645.000 ;
        RECT 305.400 644.400 306.600 646.650 ;
        RECT 317.250 644.400 318.450 657.300 ;
        RECT 319.950 655.950 322.050 658.050 ;
        RECT 334.050 657.300 336.150 659.400 ;
        RECT 338.400 658.050 339.450 712.950 ;
        RECT 341.550 693.300 343.650 695.400 ;
        RECT 341.550 686.700 342.750 693.300 ;
        RECT 355.950 688.950 358.050 691.050 ;
        RECT 341.550 684.600 343.650 686.700 ;
        RECT 352.950 685.950 355.050 688.050 ;
        RECT 341.550 671.700 342.750 684.600 ;
        RECT 346.950 679.950 349.050 682.050 ;
        RECT 347.400 678.900 348.600 679.650 ;
        RECT 353.400 678.900 354.450 685.950 ;
        RECT 346.950 676.800 349.050 678.900 ;
        RECT 352.950 676.800 355.050 678.900 ;
        RECT 356.400 676.050 357.450 688.950 ;
        RECT 362.400 688.050 363.450 719.400 ;
        RECT 367.950 709.950 370.050 712.050 ;
        RECT 361.950 685.950 364.050 688.050 ;
        RECT 362.400 684.600 363.450 685.950 ;
        RECT 368.400 684.600 369.450 709.950 ;
        RECT 371.400 709.050 372.450 728.100 ;
        RECT 380.400 727.350 381.600 728.100 ;
        RECT 376.950 724.950 379.050 727.050 ;
        RECT 379.950 724.950 382.050 727.050 ;
        RECT 382.950 724.950 385.050 727.050 ;
        RECT 377.400 722.400 378.600 724.650 ;
        RECT 383.400 722.400 384.600 724.650 ;
        RECT 377.400 709.050 378.450 722.400 ;
        RECT 383.400 718.050 384.450 722.400 ;
        RECT 382.950 715.950 385.050 718.050 ;
        RECT 370.950 706.950 373.050 709.050 ;
        RECT 376.950 706.950 379.050 709.050 ;
        RECT 389.400 700.050 390.450 730.950 ;
        RECT 395.400 729.600 396.450 742.950 ;
        RECT 403.950 733.950 406.050 736.050 ;
        RECT 395.400 727.350 396.600 729.600 ;
        RECT 394.950 724.950 397.050 727.050 ;
        RECT 397.950 724.950 400.050 727.050 ;
        RECT 398.400 722.400 399.600 724.650 ;
        RECT 394.950 718.950 397.050 721.050 ;
        RECT 373.950 697.950 376.050 700.050 ;
        RECT 388.950 697.950 391.050 700.050 ;
        RECT 362.400 682.350 363.600 684.600 ;
        RECT 368.400 682.350 369.600 684.600 ;
        RECT 361.950 679.950 364.050 682.050 ;
        RECT 364.950 679.950 367.050 682.050 ;
        RECT 367.950 679.950 370.050 682.050 ;
        RECT 365.400 678.900 366.600 679.650 ;
        RECT 364.950 676.800 367.050 678.900 ;
        RECT 355.950 673.950 358.050 676.050 ;
        RECT 352.950 672.900 357.000 673.050 ;
        RECT 341.550 669.600 343.650 671.700 ;
        RECT 352.950 670.950 358.050 672.900 ;
        RECT 358.950 670.950 364.050 673.050 ;
        RECT 355.950 670.800 358.050 670.950 ;
        RECT 364.950 664.950 367.050 667.050 ;
        RECT 349.950 658.950 352.050 661.050 ;
        RECT 259.950 631.950 262.050 634.050 ;
        RECT 265.950 631.950 268.050 634.050 ;
        RECT 280.950 631.950 283.050 634.050 ;
        RECT 253.950 622.950 256.050 625.050 ;
        RECT 247.950 616.950 250.050 619.050 ;
        RECT 235.950 610.950 238.050 613.050 ;
        RECT 236.400 606.600 237.450 610.950 ;
        RECT 236.400 604.350 237.600 606.600 ;
        RECT 241.950 605.100 244.050 607.200 ;
        RECT 248.400 606.600 249.450 616.950 ;
        RECT 254.250 613.500 256.350 614.400 ;
        RECT 252.150 612.300 256.350 613.500 ;
        RECT 242.400 604.350 243.600 605.100 ;
        RECT 248.400 604.350 249.600 606.600 ;
        RECT 232.950 601.950 235.050 604.050 ;
        RECT 235.950 601.950 238.050 604.050 ;
        RECT 238.950 601.950 241.050 604.050 ;
        RECT 241.950 601.950 244.050 604.050 ;
        RECT 247.950 601.950 250.050 604.050 ;
        RECT 226.950 598.950 229.050 601.050 ;
        RECT 233.400 600.900 234.600 601.650 ;
        RECT 239.400 600.900 240.600 601.650 ;
        RECT 232.950 598.800 235.050 600.900 ;
        RECT 238.950 598.800 241.050 600.900 ;
        RECT 214.050 591.600 216.150 593.700 ;
        RECT 211.950 580.950 214.050 583.050 ;
        RECT 190.950 568.950 193.050 571.050 ;
        RECT 185.550 564.300 187.650 566.400 ;
        RECT 185.550 557.700 186.750 564.300 ;
        RECT 185.550 555.600 187.650 557.700 ;
        RECT 181.950 550.950 184.050 553.050 ;
        RECT 187.950 550.950 190.050 553.050 ;
        RECT 181.950 538.950 184.050 541.050 ;
        RECT 169.950 535.950 172.050 538.050 ;
        RECT 163.950 529.950 166.050 532.050 ;
        RECT 155.400 526.350 156.600 528.600 ;
        RECT 161.400 526.350 162.600 528.600 ;
        RECT 154.950 523.950 157.050 526.050 ;
        RECT 157.950 523.950 160.050 526.050 ;
        RECT 160.950 523.950 163.050 526.050 ;
        RECT 163.950 523.950 166.050 526.050 ;
        RECT 158.400 521.400 159.600 523.650 ;
        RECT 164.400 522.900 165.600 523.650 ;
        RECT 158.400 517.050 159.450 521.400 ;
        RECT 163.950 520.800 166.050 522.900 ;
        RECT 170.400 522.450 171.450 535.950 ;
        RECT 175.950 527.100 178.050 529.200 ;
        RECT 182.400 528.600 183.450 538.950 ;
        RECT 176.400 526.350 177.600 527.100 ;
        RECT 182.400 526.350 183.600 528.600 ;
        RECT 175.950 523.950 178.050 526.050 ;
        RECT 178.950 523.950 181.050 526.050 ;
        RECT 181.950 523.950 184.050 526.050 ;
        RECT 167.400 521.400 171.450 522.450 ;
        RECT 179.400 522.000 180.600 523.650 ;
        RECT 157.950 514.950 160.050 517.050 ;
        RECT 158.400 502.050 159.450 514.950 ;
        RECT 157.950 499.950 160.050 502.050 ;
        RECT 148.950 495.450 151.050 496.050 ;
        RECT 152.400 495.450 153.600 495.600 ;
        RECT 148.950 494.400 153.600 495.450 ;
        RECT 148.950 493.950 151.050 494.400 ;
        RECT 152.400 493.350 153.600 494.400 ;
        RECT 157.950 494.100 160.050 496.200 ;
        RECT 163.950 494.100 166.050 496.200 ;
        RECT 158.400 493.350 159.600 494.100 ;
        RECT 151.950 490.950 154.050 493.050 ;
        RECT 154.950 490.950 157.050 493.050 ;
        RECT 157.950 490.950 160.050 493.050 ;
        RECT 140.400 488.400 144.450 489.450 ;
        RECT 145.950 487.950 148.050 490.050 ;
        RECT 155.400 489.900 156.600 490.650 ;
        RECT 154.950 487.800 157.050 489.900 ;
        RECT 127.800 482.400 129.900 484.500 ;
        RECT 137.400 483.600 139.500 485.700 ;
        RECT 142.950 484.950 145.050 487.050 ;
        RECT 118.950 478.950 121.050 481.050 ;
        RECT 127.950 478.950 130.050 481.050 ;
        RECT 118.950 463.950 121.050 466.050 ;
        RECT 85.950 454.800 88.050 456.900 ;
        RECT 100.950 454.950 103.050 457.050 ;
        RECT 86.400 450.600 87.450 454.800 ;
        RECT 86.400 448.350 87.600 450.600 ;
        RECT 94.950 449.100 97.050 451.200 ;
        RECT 103.950 449.100 106.050 451.200 ;
        RECT 109.950 449.100 112.050 451.200 ;
        RECT 115.950 449.100 118.050 451.200 ;
        RECT 82.950 445.950 85.050 448.050 ;
        RECT 85.950 445.950 88.050 448.050 ;
        RECT 88.950 445.950 91.050 448.050 ;
        RECT 83.400 443.400 84.600 445.650 ;
        RECT 89.400 444.900 90.600 445.650 ;
        RECT 95.400 445.050 96.450 449.100 ;
        RECT 104.400 448.350 105.600 449.100 ;
        RECT 110.400 448.350 111.600 449.100 ;
        RECT 100.950 445.950 103.050 448.050 ;
        RECT 103.950 445.950 106.050 448.050 ;
        RECT 106.950 445.950 109.050 448.050 ;
        RECT 109.950 445.950 112.050 448.050 ;
        RECT 79.350 423.300 81.450 425.400 ;
        RECT 73.950 418.950 76.050 421.050 ;
        RECT 64.950 416.100 67.050 418.200 ;
        RECT 70.950 417.600 75.000 418.050 ;
        RECT 65.400 415.350 66.600 416.100 ;
        RECT 70.950 415.950 75.600 417.600 ;
        RECT 74.400 415.350 75.600 415.950 ;
        RECT 64.950 412.950 67.050 415.050 ;
        RECT 67.950 412.950 70.050 415.050 ;
        RECT 73.950 412.950 76.050 415.050 ;
        RECT 49.950 409.800 52.050 411.900 ;
        RECT 58.950 409.950 61.050 412.050 ;
        RECT 68.400 411.900 69.600 412.650 ;
        RECT 67.950 409.800 70.050 411.900 ;
        RECT 80.250 410.400 81.450 423.300 ;
        RECT 83.400 423.450 84.450 443.400 ;
        RECT 88.950 442.800 91.050 444.900 ;
        RECT 94.950 442.950 97.050 445.050 ;
        RECT 101.400 444.900 102.600 445.650 ;
        RECT 100.950 442.800 103.050 444.900 ;
        RECT 107.400 443.400 108.600 445.650 ;
        RECT 107.400 439.050 108.450 443.400 ;
        RECT 116.400 439.050 117.450 449.100 ;
        RECT 119.400 444.450 120.450 463.950 ;
        RECT 128.400 451.200 129.450 478.950 ;
        RECT 136.950 451.950 139.050 454.050 ;
        RECT 127.950 450.450 130.050 451.200 ;
        RECT 127.950 449.400 132.450 450.450 ;
        RECT 127.950 449.100 130.050 449.400 ;
        RECT 128.400 448.350 129.600 449.100 ;
        RECT 122.400 445.950 124.500 448.050 ;
        RECT 127.800 445.950 129.900 448.050 ;
        RECT 122.400 444.450 123.600 445.650 ;
        RECT 131.400 445.050 132.450 449.400 ;
        RECT 119.400 443.400 123.600 444.450 ;
        RECT 106.950 436.950 109.050 439.050 ;
        RECT 115.950 436.950 118.050 439.050 ;
        RECT 83.400 422.400 87.450 423.450 ;
        RECT 97.050 423.300 99.150 425.400 ;
        RECT 82.950 418.950 85.050 421.050 ;
        RECT 26.550 399.600 28.650 401.700 ;
        RECT 40.950 400.950 43.050 403.050 ;
        RECT 22.950 385.950 25.050 388.050 ;
        RECT 28.950 385.950 31.050 388.050 ;
        RECT 25.350 381.300 27.450 383.400 ;
        RECT 10.950 371.100 13.050 376.050 ;
        RECT 19.950 373.950 22.050 376.050 ;
        RECT 26.250 374.700 27.450 381.300 ;
        RECT 25.350 372.600 27.450 374.700 ;
        RECT 11.400 370.350 12.600 371.100 ;
        RECT 10.950 367.950 13.050 370.050 ;
        RECT 13.950 367.950 16.050 370.050 ;
        RECT 19.950 367.950 22.050 370.050 ;
        RECT 14.400 366.900 15.600 367.650 ;
        RECT 20.400 366.900 21.600 367.650 ;
        RECT 13.950 364.800 16.050 366.900 ;
        RECT 19.950 364.800 22.050 366.900 ;
        RECT 10.950 361.950 13.050 364.050 ;
        RECT 11.400 339.600 12.450 361.950 ;
        RECT 26.250 359.700 27.450 372.600 ;
        RECT 29.400 366.900 30.450 385.950 ;
        RECT 41.400 385.050 42.450 400.950 ;
        RECT 40.950 382.950 43.050 385.050 ;
        RECT 46.950 382.950 49.050 385.050 ;
        RECT 55.950 382.950 58.050 385.050 ;
        RECT 40.650 379.500 42.750 380.400 ;
        RECT 40.650 378.300 44.850 379.500 ;
        RECT 31.950 370.950 34.050 373.050 ;
        RECT 37.950 371.100 40.050 373.200 ;
        RECT 28.950 364.800 31.050 366.900 ;
        RECT 25.350 357.600 27.450 359.700 ;
        RECT 32.400 346.050 33.450 370.950 ;
        RECT 38.400 370.350 39.600 371.100 ;
        RECT 37.800 367.950 39.900 370.050 ;
        RECT 43.650 359.700 44.850 378.300 ;
        RECT 47.400 372.600 48.450 382.950 ;
        RECT 56.400 372.600 57.450 382.950 ;
        RECT 62.250 379.500 64.350 380.400 ;
        RECT 60.150 378.300 64.350 379.500 ;
        RECT 47.400 370.350 48.600 372.600 ;
        RECT 56.400 370.350 57.600 372.600 ;
        RECT 46.950 367.950 49.050 370.050 ;
        RECT 55.950 367.950 58.050 370.050 ;
        RECT 60.150 359.700 61.350 378.300 ;
        RECT 68.400 376.050 69.450 409.800 ;
        RECT 79.350 408.300 81.450 410.400 ;
        RECT 80.250 401.700 81.450 408.300 ;
        RECT 79.350 399.600 81.450 401.700 ;
        RECT 77.550 381.300 79.650 383.400 ;
        RECT 67.950 373.950 70.050 376.050 ;
        RECT 73.950 373.950 76.050 376.050 ;
        RECT 77.550 374.700 78.750 381.300 ;
        RECT 83.400 376.050 84.450 418.950 ;
        RECT 86.400 411.900 87.450 422.400 ;
        RECT 91.800 412.950 93.900 415.050 ;
        RECT 85.950 409.800 88.050 411.900 ;
        RECT 92.400 410.400 93.600 412.650 ;
        RECT 92.400 408.450 93.450 410.400 ;
        RECT 89.400 407.400 93.450 408.450 ;
        RECT 64.950 371.100 67.050 373.200 ;
        RECT 65.400 370.350 66.600 371.100 ;
        RECT 65.100 367.950 67.200 370.050 ;
        RECT 43.050 357.600 45.150 359.700 ;
        RECT 59.850 357.600 61.950 359.700 ;
        RECT 16.950 343.950 19.050 346.050 ;
        RECT 31.950 343.950 34.050 346.050 ;
        RECT 17.400 339.600 18.450 343.950 ;
        RECT 11.400 337.350 12.600 339.600 ;
        RECT 17.400 337.350 18.600 339.600 ;
        RECT 22.950 338.100 25.050 340.200 ;
        RECT 28.800 338.100 30.900 340.200 ;
        RECT 23.400 337.350 24.600 338.100 ;
        RECT 10.950 334.950 13.050 337.050 ;
        RECT 13.950 334.950 16.050 337.050 ;
        RECT 16.950 334.950 19.050 337.050 ;
        RECT 19.950 334.950 22.050 337.050 ;
        RECT 22.950 334.950 25.050 337.050 ;
        RECT 14.400 332.400 15.600 334.650 ;
        RECT 20.400 333.900 21.600 334.650 ;
        RECT 14.400 316.050 15.450 332.400 ;
        RECT 19.950 331.800 22.050 333.900 ;
        RECT 13.950 313.950 16.050 316.050 ;
        RECT 4.950 293.100 7.050 295.200 ;
        RECT 10.950 293.100 13.050 295.200 ;
        RECT 16.950 294.000 19.050 298.050 ;
        RECT 22.950 295.950 28.050 298.050 ;
        RECT 29.400 294.450 30.450 338.100 ;
        RECT 31.950 337.950 34.050 340.050 ;
        RECT 40.950 338.100 43.050 340.200 ;
        RECT 58.950 338.100 61.050 340.200 ;
        RECT 32.400 333.900 33.450 337.950 ;
        RECT 41.400 337.350 42.600 338.100 ;
        RECT 59.400 337.350 60.600 338.100 ;
        RECT 67.950 337.950 70.050 340.050 ;
        RECT 74.400 339.600 75.450 373.950 ;
        RECT 77.550 372.600 79.650 374.700 ;
        RECT 82.950 373.950 85.050 376.050 ;
        RECT 77.550 359.700 78.750 372.600 ;
        RECT 82.950 367.950 85.050 370.050 ;
        RECT 83.400 366.900 84.600 367.650 ;
        RECT 82.950 364.800 85.050 366.900 ;
        RECT 77.550 357.600 79.650 359.700 ;
        RECT 89.400 343.050 90.450 407.400 ;
        RECT 97.650 404.700 98.850 423.300 ;
        RECT 122.400 417.600 123.450 443.400 ;
        RECT 130.950 442.950 133.050 445.050 ;
        RECT 137.400 442.050 138.450 451.950 ;
        RECT 143.400 450.600 144.450 484.950 ;
        RECT 164.400 481.050 165.450 494.100 ;
        RECT 148.950 478.950 151.050 481.050 ;
        RECT 163.950 478.950 166.050 481.050 ;
        RECT 149.400 454.050 150.450 478.950 ;
        RECT 154.950 475.950 157.050 478.050 ;
        RECT 143.400 448.350 144.600 450.600 ;
        RECT 148.950 450.000 151.050 454.050 ;
        RECT 149.400 448.350 150.600 450.000 ;
        RECT 142.950 445.950 145.050 448.050 ;
        RECT 145.950 445.950 148.050 448.050 ;
        RECT 148.950 445.950 151.050 448.050 ;
        RECT 146.400 444.900 147.600 445.650 ;
        RECT 145.950 442.800 148.050 444.900 ;
        RECT 155.400 444.450 156.450 475.950 ;
        RECT 160.950 460.950 163.050 463.050 ;
        RECT 161.400 451.200 162.450 460.950 ;
        RECT 167.400 460.050 168.450 521.400 ;
        RECT 178.950 517.950 181.050 522.000 ;
        RECT 181.950 514.950 184.050 517.050 ;
        RECT 182.400 508.050 183.450 514.950 ;
        RECT 181.950 505.950 184.050 508.050 ;
        RECT 184.950 502.950 187.050 505.050 ;
        RECT 169.950 499.950 172.050 502.050 ;
        RECT 170.400 489.450 171.450 499.950 ;
        RECT 175.950 494.100 178.050 496.200 ;
        RECT 176.400 493.350 177.600 494.100 ;
        RECT 185.400 493.050 186.450 502.950 ;
        RECT 173.100 490.950 175.200 493.050 ;
        RECT 176.400 490.950 178.500 493.050 ;
        RECT 181.800 490.950 183.900 493.050 ;
        RECT 184.950 490.950 187.050 493.050 ;
        RECT 173.400 489.450 174.600 490.650 ;
        RECT 170.400 488.400 174.600 489.450 ;
        RECT 182.400 488.400 183.600 490.650 ;
        RECT 172.950 484.950 175.050 487.050 ;
        RECT 166.950 457.950 169.050 460.050 ;
        RECT 160.950 449.100 163.050 451.200 ;
        RECT 166.950 449.100 169.050 451.200 ;
        RECT 161.400 448.350 162.600 449.100 ;
        RECT 167.400 448.350 168.600 449.100 ;
        RECT 160.950 445.950 163.050 448.050 ;
        RECT 163.950 445.950 166.050 448.050 ;
        RECT 166.950 445.950 169.050 448.050 ;
        RECT 152.400 443.400 156.450 444.450 ;
        RECT 164.400 444.000 165.600 445.650 ;
        RECT 136.950 439.950 139.050 442.050 ;
        RECT 142.950 439.950 145.050 442.050 ;
        RECT 133.950 433.950 136.050 436.050 ;
        RECT 134.400 421.050 135.450 433.950 ;
        RECT 143.400 423.450 144.450 439.950 ;
        RECT 143.400 421.200 144.600 423.450 ;
        RECT 133.950 418.950 136.050 421.050 ;
        RECT 138.900 417.900 141.000 419.700 ;
        RECT 142.800 418.800 144.900 420.900 ;
        RECT 146.100 420.300 148.200 422.400 ;
        RECT 122.400 415.350 123.600 417.600 ;
        RECT 137.400 416.700 146.100 417.900 ;
        RECT 100.950 412.950 103.050 415.050 ;
        RECT 116.100 412.950 118.200 415.050 ;
        RECT 121.500 412.950 123.600 415.050 ;
        RECT 134.100 412.950 136.200 415.050 ;
        RECT 94.650 403.500 98.850 404.700 ;
        RECT 101.400 410.400 102.600 412.650 ;
        RECT 116.400 410.400 117.600 412.650 ;
        RECT 134.400 411.900 135.600 412.650 ;
        RECT 94.650 402.600 96.750 403.500 ;
        RECT 101.400 403.050 102.450 410.400 ;
        RECT 100.950 400.950 103.050 403.050 ;
        RECT 116.400 382.050 117.450 410.400 ;
        RECT 133.950 409.800 136.050 411.900 ;
        RECT 137.400 407.700 138.300 416.700 ;
        RECT 144.000 415.800 146.100 416.700 ;
        RECT 147.000 414.900 147.900 420.300 ;
        RECT 148.950 416.100 151.050 418.200 ;
        RECT 149.400 415.350 150.600 416.100 ;
        RECT 141.000 413.700 147.900 414.900 ;
        RECT 141.000 411.300 141.900 413.700 ;
        RECT 139.800 409.200 141.900 411.300 ;
        RECT 142.800 409.950 144.900 412.050 ;
        RECT 136.500 405.600 138.600 407.700 ;
        RECT 143.400 407.400 144.600 409.650 ;
        RECT 146.700 406.500 147.900 413.700 ;
        RECT 148.800 412.950 150.900 415.050 ;
        RECT 146.100 404.400 148.200 406.500 ;
        RECT 127.950 400.950 130.050 403.050 ;
        RECT 115.950 379.950 118.050 382.050 ;
        RECT 91.950 370.950 94.050 373.050 ;
        RECT 100.950 372.000 103.050 376.050 ;
        RECT 106.950 373.950 109.050 376.050 ;
        RECT 92.400 358.050 93.450 370.950 ;
        RECT 101.400 370.350 102.600 372.000 ;
        RECT 97.950 367.950 100.050 370.050 ;
        RECT 100.950 367.950 103.050 370.050 ;
        RECT 98.400 366.900 99.600 367.650 ;
        RECT 107.400 366.900 108.450 373.950 ;
        RECT 116.400 372.600 117.450 379.950 ;
        RECT 116.400 370.350 117.600 372.600 ;
        RECT 121.950 371.100 124.050 373.200 ;
        RECT 128.400 372.600 129.450 400.950 ;
        RECT 152.400 400.050 153.450 443.400 ;
        RECT 163.950 439.950 166.050 444.000 ;
        RECT 173.400 442.050 174.450 484.950 ;
        RECT 182.400 484.050 183.450 488.400 ;
        RECT 181.950 481.950 184.050 484.050 ;
        RECT 182.400 478.050 183.450 481.950 ;
        RECT 188.400 481.050 189.450 550.950 ;
        RECT 197.400 538.050 198.450 571.950 ;
        RECT 200.400 568.050 201.450 572.100 ;
        RECT 202.950 571.950 205.050 574.050 ;
        RECT 205.950 572.100 208.050 574.200 ;
        RECT 212.400 573.600 213.450 580.950 ;
        RECT 233.400 577.050 234.450 598.800 ;
        RECT 252.150 593.700 253.350 612.300 ;
        RECT 256.950 605.100 259.050 607.200 ;
        RECT 262.950 605.100 265.050 607.200 ;
        RECT 257.400 604.350 258.600 605.100 ;
        RECT 257.100 601.950 259.200 604.050 ;
        RECT 251.850 591.600 253.950 593.700 ;
        RECT 263.400 589.050 264.450 605.100 ;
        RECT 262.950 586.950 265.050 589.050 ;
        RECT 238.950 583.950 241.050 586.050 ;
        RECT 239.400 580.050 240.450 583.950 ;
        RECT 266.400 583.050 267.450 631.950 ;
        RECT 269.550 615.300 271.650 617.400 ;
        RECT 269.550 608.700 270.750 615.300 ;
        RECT 269.550 606.600 271.650 608.700 ;
        RECT 284.400 607.200 285.450 640.950 ;
        RECT 295.950 637.950 298.050 640.050 ;
        RECT 269.550 593.700 270.750 606.600 ;
        RECT 283.950 605.100 286.050 607.200 ;
        RECT 289.950 605.100 292.050 607.200 ;
        RECT 296.400 606.600 297.450 637.950 ;
        RECT 305.400 634.050 306.450 644.400 ;
        RECT 316.350 642.300 318.450 644.400 ;
        RECT 317.250 635.700 318.450 642.300 ;
        RECT 304.950 631.950 307.050 634.050 ;
        RECT 316.350 633.600 318.450 635.700 ;
        RECT 301.950 628.950 304.050 631.050 ;
        RECT 302.400 607.200 303.450 628.950 ;
        RECT 313.350 615.300 315.450 617.400 ;
        RECT 314.250 608.700 315.450 615.300 ;
        RECT 274.950 601.950 277.050 604.050 ;
        RECT 275.400 599.400 276.600 601.650 ;
        RECT 269.550 591.600 271.650 593.700 ;
        RECT 271.950 586.950 274.050 589.050 ;
        RECT 241.950 580.950 244.050 583.050 ;
        RECT 265.950 580.950 268.050 583.050 ;
        RECT 238.950 577.950 241.050 580.050 ;
        RECT 206.400 571.350 207.600 572.100 ;
        RECT 212.400 571.350 213.600 573.600 ;
        RECT 217.950 571.950 220.050 577.050 ;
        RECT 232.950 574.950 235.050 577.050 ;
        RECT 229.950 572.100 232.050 574.200 ;
        RECT 230.400 571.350 231.600 572.100 ;
        RECT 205.950 568.950 208.050 571.050 ;
        RECT 208.950 568.950 211.050 571.050 ;
        RECT 211.950 568.950 214.050 571.050 ;
        RECT 214.950 568.950 217.050 571.050 ;
        RECT 226.950 568.950 229.050 571.050 ;
        RECT 229.950 568.950 232.050 571.050 ;
        RECT 232.950 568.950 235.050 571.050 ;
        RECT 199.950 565.950 202.050 568.050 ;
        RECT 209.400 566.400 210.600 568.650 ;
        RECT 215.400 568.050 216.600 568.650 ;
        RECT 215.400 566.400 220.050 568.050 ;
        RECT 227.400 567.900 228.600 568.650 ;
        RECT 233.400 567.900 234.600 568.650 ;
        RECT 239.400 568.050 240.450 577.950 ;
        RECT 196.950 535.950 199.050 538.050 ;
        RECT 190.950 529.950 193.050 532.050 ;
        RECT 191.400 505.050 192.450 529.950 ;
        RECT 196.950 528.000 199.050 532.050 ;
        RECT 197.400 526.350 198.600 528.000 ;
        RECT 197.100 523.950 199.200 526.050 ;
        RECT 209.400 511.050 210.450 566.400 ;
        RECT 216.000 565.950 220.050 566.400 ;
        RECT 226.950 565.800 229.050 567.900 ;
        RECT 232.950 565.800 235.050 567.900 ;
        RECT 238.950 565.950 241.050 568.050 ;
        RECT 227.400 556.050 228.450 565.800 ;
        RECT 235.950 556.950 238.050 559.050 ;
        RECT 226.950 553.950 229.050 556.050 ;
        RECT 229.950 553.950 232.050 556.050 ;
        RECT 223.950 544.950 226.050 547.050 ;
        RECT 215.100 523.950 217.200 526.050 ;
        RECT 208.950 508.950 211.050 511.050 ;
        RECT 190.950 502.950 193.050 505.050 ;
        RECT 193.950 499.950 196.050 502.050 ;
        RECT 212.850 501.300 214.950 503.400 ;
        RECT 194.400 495.600 195.450 499.950 ;
        RECT 194.400 493.350 195.600 495.600 ;
        RECT 199.950 494.100 202.050 496.200 ;
        RECT 200.400 493.350 201.600 494.100 ;
        RECT 193.950 490.950 196.050 493.050 ;
        RECT 196.950 490.950 199.050 493.050 ;
        RECT 199.950 490.950 202.050 493.050 ;
        RECT 202.950 490.950 205.050 493.050 ;
        RECT 208.950 490.950 211.050 493.050 ;
        RECT 197.400 489.900 198.600 490.650 ;
        RECT 196.950 487.800 199.050 489.900 ;
        RECT 203.400 488.400 204.600 490.650 ;
        RECT 209.400 489.900 210.600 490.650 ;
        RECT 203.400 481.050 204.450 488.400 ;
        RECT 208.950 487.800 211.050 489.900 ;
        RECT 213.150 482.700 214.350 501.300 ;
        RECT 218.100 490.950 220.200 493.050 ;
        RECT 218.400 489.900 219.600 490.650 ;
        RECT 217.950 487.800 220.050 489.900 ;
        RECT 213.150 481.500 217.350 482.700 ;
        RECT 187.950 478.950 190.050 481.050 ;
        RECT 193.950 478.950 196.050 481.050 ;
        RECT 202.950 478.950 205.050 481.050 ;
        RECT 215.250 480.600 217.350 481.500 ;
        RECT 181.950 475.950 184.050 478.050 ;
        RECT 190.950 457.950 193.050 460.050 ;
        RECT 178.950 449.100 181.050 451.200 ;
        RECT 184.950 449.100 187.050 451.200 ;
        RECT 191.400 451.050 192.450 457.950 ;
        RECT 179.400 448.350 180.600 449.100 ;
        RECT 185.400 448.350 186.600 449.100 ;
        RECT 190.950 448.950 193.050 451.050 ;
        RECT 178.950 445.950 181.050 448.050 ;
        RECT 181.950 445.950 184.050 448.050 ;
        RECT 184.950 445.950 187.050 448.050 ;
        RECT 187.950 445.950 190.050 448.050 ;
        RECT 175.950 442.950 178.050 445.050 ;
        RECT 182.400 443.400 183.600 445.650 ;
        RECT 188.400 444.900 189.600 445.650 ;
        RECT 172.950 439.950 175.050 442.050 ;
        RECT 169.950 433.950 172.050 436.050 ;
        RECT 154.950 415.950 157.050 418.050 ;
        RECT 163.950 417.000 166.050 421.050 ;
        RECT 170.400 418.050 171.450 433.950 ;
        RECT 176.400 418.050 177.450 442.950 ;
        RECT 182.400 430.050 183.450 443.400 ;
        RECT 187.950 442.800 190.050 444.900 ;
        RECT 190.950 442.950 193.050 445.050 ;
        RECT 181.950 427.950 184.050 430.050 ;
        RECT 191.400 427.050 192.450 442.950 ;
        RECT 184.950 424.950 187.050 427.050 ;
        RECT 190.950 424.950 193.050 427.050 ;
        RECT 155.400 411.900 156.450 415.950 ;
        RECT 164.400 415.350 165.600 417.000 ;
        RECT 169.950 415.950 172.050 418.050 ;
        RECT 175.950 415.950 178.050 418.050 ;
        RECT 178.950 417.000 181.050 421.050 ;
        RECT 185.400 417.600 186.450 424.950 ;
        RECT 179.400 415.350 180.600 417.000 ;
        RECT 185.400 415.350 186.600 417.600 ;
        RECT 160.950 412.950 163.050 415.050 ;
        RECT 163.950 412.950 166.050 415.050 ;
        RECT 166.950 412.950 169.050 415.050 ;
        RECT 178.950 412.950 181.050 415.050 ;
        RECT 181.950 412.950 184.050 415.050 ;
        RECT 184.950 412.950 187.050 415.050 ;
        RECT 187.950 412.950 190.050 415.050 ;
        RECT 161.400 411.900 162.600 412.650 ;
        RECT 167.400 411.900 168.600 412.650 ;
        RECT 154.950 409.800 157.050 411.900 ;
        RECT 160.950 409.800 163.050 411.900 ;
        RECT 166.950 409.800 169.050 411.900 ;
        RECT 175.950 409.950 178.050 412.050 ;
        RECT 182.400 411.900 183.600 412.650 ;
        RECT 151.950 397.950 154.050 400.050 ;
        RECT 149.550 381.300 151.650 383.400 ;
        RECT 134.250 379.500 136.350 380.400 ;
        RECT 132.150 378.300 136.350 379.500 ;
        RECT 122.400 370.350 123.600 371.100 ;
        RECT 128.400 370.350 129.600 372.600 ;
        RECT 112.950 367.950 115.050 370.050 ;
        RECT 115.950 367.950 118.050 370.050 ;
        RECT 118.950 367.950 121.050 370.050 ;
        RECT 121.950 367.950 124.050 370.050 ;
        RECT 127.950 367.950 130.050 370.050 ;
        RECT 113.400 366.900 114.600 367.650 ;
        RECT 97.950 364.800 100.050 366.900 ;
        RECT 106.950 364.800 109.050 366.900 ;
        RECT 112.950 364.800 115.050 366.900 ;
        RECT 119.400 365.400 120.600 367.650 ;
        RECT 119.400 358.050 120.450 365.400 ;
        RECT 132.150 359.700 133.350 378.300 ;
        RECT 149.550 374.700 150.750 381.300 ;
        RECT 136.950 371.100 139.050 373.200 ;
        RECT 142.950 371.100 145.050 373.200 ;
        RECT 149.550 372.600 151.650 374.700 ;
        RECT 137.400 370.350 138.600 371.100 ;
        RECT 137.100 367.950 139.200 370.050 ;
        RECT 143.400 361.050 144.450 371.100 ;
        RECT 145.950 364.950 148.050 367.050 ;
        RECT 91.950 355.950 94.050 358.050 ;
        RECT 118.950 355.950 121.050 358.050 ;
        RECT 131.850 357.600 133.950 359.700 ;
        RECT 142.950 358.950 145.050 361.050 ;
        RECT 146.400 358.050 147.450 364.950 ;
        RECT 149.550 359.700 150.750 372.600 ;
        RECT 154.950 367.950 157.050 370.050 ;
        RECT 155.400 366.900 156.600 367.650 ;
        RECT 161.400 366.900 162.450 409.800 ;
        RECT 163.950 379.950 166.050 382.050 ;
        RECT 154.950 364.800 157.050 366.900 ;
        RECT 160.950 364.800 163.050 366.900 ;
        RECT 145.950 355.950 148.050 358.050 ;
        RECT 149.550 357.600 151.650 359.700 ;
        RECT 160.950 349.950 163.050 352.050 ;
        RECT 91.950 343.950 94.050 346.050 ;
        RECT 151.950 343.950 154.050 346.050 ;
        RECT 37.950 334.950 40.050 337.050 ;
        RECT 40.950 334.950 43.050 337.050 ;
        RECT 43.950 334.950 46.050 337.050 ;
        RECT 55.950 334.950 58.050 337.050 ;
        RECT 58.950 334.950 61.050 337.050 ;
        RECT 61.950 334.950 64.050 337.050 ;
        RECT 31.950 331.800 34.050 333.900 ;
        RECT 38.400 332.400 39.600 334.650 ;
        RECT 44.400 333.450 45.600 334.650 ;
        RECT 44.400 332.400 48.450 333.450 ;
        RECT 38.400 316.050 39.450 332.400 ;
        RECT 37.950 313.950 40.050 316.050 ;
        RECT 1.950 283.950 4.050 286.050 ;
        RECT 1.950 253.800 4.050 255.900 ;
        RECT 2.400 211.050 3.450 253.800 ;
        RECT 5.400 247.050 6.450 293.100 ;
        RECT 11.400 292.350 12.600 293.100 ;
        RECT 17.400 292.350 18.600 294.000 ;
        RECT 26.400 293.400 30.450 294.450 ;
        RECT 10.950 289.950 13.050 292.050 ;
        RECT 13.950 289.950 16.050 292.050 ;
        RECT 16.950 289.950 19.050 292.050 ;
        RECT 19.950 289.950 22.050 292.050 ;
        RECT 14.400 287.400 15.600 289.650 ;
        RECT 20.400 288.450 21.600 289.650 ;
        RECT 26.400 288.450 27.450 293.400 ;
        RECT 31.950 293.100 34.050 295.200 ;
        RECT 37.950 293.100 40.050 298.050 ;
        RECT 32.400 292.350 33.600 293.100 ;
        RECT 38.400 292.350 39.600 293.100 ;
        RECT 31.950 289.950 34.050 292.050 ;
        RECT 34.950 289.950 37.050 292.050 ;
        RECT 37.950 289.950 40.050 292.050 ;
        RECT 40.950 289.950 43.050 292.050 ;
        RECT 20.400 287.400 27.450 288.450 ;
        RECT 35.400 287.400 36.600 289.650 ;
        RECT 41.400 288.000 42.600 289.650 ;
        RECT 14.400 280.050 15.450 287.400 ;
        RECT 19.950 283.950 22.050 286.050 ;
        RECT 28.950 283.950 31.050 286.050 ;
        RECT 35.400 285.450 36.450 287.400 ;
        RECT 32.400 284.400 36.450 285.450 ;
        RECT 13.950 277.950 16.050 280.050 ;
        RECT 20.400 267.450 21.450 283.950 ;
        RECT 13.500 263.400 15.600 265.500 ;
        RECT 20.400 265.200 21.600 267.450 ;
        RECT 7.950 260.100 10.050 262.200 ;
        RECT 4.950 244.950 7.050 247.050 ;
        RECT 8.400 243.450 9.450 260.100 ;
        RECT 11.100 256.950 13.200 259.050 ;
        RECT 11.400 255.900 12.600 256.650 ;
        RECT 10.950 253.800 13.050 255.900 ;
        RECT 14.100 250.800 15.000 263.400 ;
        RECT 20.100 262.800 22.200 264.900 ;
        RECT 23.400 263.100 25.500 265.200 ;
        RECT 15.900 261.000 18.000 261.900 ;
        RECT 15.900 259.800 23.100 261.000 ;
        RECT 21.000 258.900 23.100 259.800 ;
        RECT 15.900 258.000 18.000 258.900 ;
        RECT 24.000 258.000 24.900 263.100 ;
        RECT 25.950 260.100 28.050 262.200 ;
        RECT 26.400 259.350 27.600 260.100 ;
        RECT 15.900 257.100 24.900 258.000 ;
        RECT 15.900 256.800 18.000 257.100 ;
        RECT 20.100 253.950 22.200 256.050 ;
        RECT 20.400 251.400 21.600 253.650 ;
        RECT 13.800 248.700 15.900 250.800 ;
        RECT 24.000 250.500 24.900 257.100 ;
        RECT 25.800 256.950 27.900 259.050 ;
        RECT 22.800 248.400 24.900 250.500 ;
        RECT 10.950 244.950 13.050 247.050 ;
        RECT 22.950 244.950 25.050 247.050 ;
        RECT 5.400 242.400 9.450 243.450 ;
        RECT 1.950 208.950 4.050 211.050 ;
        RECT 5.400 205.050 6.450 242.400 ;
        RECT 11.400 226.050 12.450 244.950 ;
        RECT 10.950 223.950 13.050 226.050 ;
        RECT 11.400 216.600 12.450 223.950 ;
        RECT 11.400 214.350 12.600 216.600 ;
        RECT 16.950 215.100 19.050 220.050 ;
        RECT 17.400 214.350 18.600 215.100 ;
        RECT 10.950 211.950 13.050 214.050 ;
        RECT 13.950 211.950 16.050 214.050 ;
        RECT 16.950 211.950 19.050 214.050 ;
        RECT 14.400 210.900 15.600 211.650 ;
        RECT 13.950 208.800 16.050 210.900 ;
        RECT 4.950 202.950 7.050 205.050 ;
        RECT 13.950 202.950 16.050 205.050 ;
        RECT 1.950 193.950 4.050 196.050 ;
        RECT 2.400 133.050 3.450 193.950 ;
        RECT 4.950 184.950 7.050 187.050 ;
        RECT 5.400 177.900 6.450 184.950 ;
        RECT 14.400 183.600 15.450 202.950 ;
        RECT 23.400 202.050 24.450 244.950 ;
        RECT 29.400 220.050 30.450 283.950 ;
        RECT 32.400 280.050 33.450 284.400 ;
        RECT 40.950 283.950 43.050 288.000 ;
        RECT 47.400 286.050 48.450 332.400 ;
        RECT 56.400 332.400 57.600 334.650 ;
        RECT 62.400 332.400 63.600 334.650 ;
        RECT 56.400 316.050 57.450 332.400 ;
        RECT 62.400 325.050 63.450 332.400 ;
        RECT 68.400 328.050 69.450 337.950 ;
        RECT 74.400 337.350 75.600 339.600 ;
        RECT 79.950 339.000 82.050 343.050 ;
        RECT 88.950 340.950 91.050 343.050 ;
        RECT 80.400 337.350 81.600 339.000 ;
        RECT 85.950 338.100 88.050 340.200 ;
        RECT 86.400 337.350 87.600 338.100 ;
        RECT 73.950 334.950 76.050 337.050 ;
        RECT 76.950 334.950 79.050 337.050 ;
        RECT 79.950 334.950 82.050 337.050 ;
        RECT 82.950 334.950 85.050 337.050 ;
        RECT 85.950 334.950 88.050 337.050 ;
        RECT 77.400 332.400 78.600 334.650 ;
        RECT 83.400 332.400 84.600 334.650 ;
        RECT 67.950 325.950 70.050 328.050 ;
        RECT 61.950 322.950 64.050 325.050 ;
        RECT 55.950 313.950 58.050 316.050 ;
        RECT 55.950 293.100 58.050 295.200 ;
        RECT 62.400 295.050 63.450 322.950 ;
        RECT 77.400 322.050 78.450 332.400 ;
        RECT 83.400 328.050 84.450 332.400 ;
        RECT 82.950 325.950 85.050 328.050 ;
        RECT 92.400 322.050 93.450 343.950 ;
        RECT 97.950 338.100 100.050 340.200 ;
        RECT 103.950 338.100 106.050 340.200 ;
        RECT 98.400 337.350 99.600 338.100 ;
        RECT 104.400 337.350 105.600 338.100 ;
        RECT 112.950 337.950 115.050 340.050 ;
        RECT 118.950 338.100 121.050 340.200 ;
        RECT 124.950 338.100 127.050 340.200 ;
        RECT 133.950 338.100 136.050 340.200 ;
        RECT 142.950 339.000 145.050 343.050 ;
        RECT 97.950 334.950 100.050 337.050 ;
        RECT 100.950 334.950 103.050 337.050 ;
        RECT 103.950 334.950 106.050 337.050 ;
        RECT 106.950 334.950 109.050 337.050 ;
        RECT 101.400 333.000 102.600 334.650 ;
        RECT 100.950 328.950 103.050 333.000 ;
        RECT 107.400 332.400 108.600 334.650 ;
        RECT 103.950 325.950 106.050 328.050 ;
        RECT 76.950 319.950 79.050 322.050 ;
        RECT 91.950 319.950 94.050 322.050 ;
        RECT 77.400 316.050 78.450 319.950 ;
        RECT 76.950 313.950 79.050 316.050 ;
        RECT 79.950 304.950 82.050 307.050 ;
        RECT 56.400 292.350 57.600 293.100 ;
        RECT 61.800 292.950 63.900 295.050 ;
        RECT 64.950 292.950 67.050 295.050 ;
        RECT 70.950 293.100 73.050 295.200 ;
        RECT 55.950 289.950 58.050 292.050 ;
        RECT 58.950 289.950 61.050 292.050 ;
        RECT 59.400 288.900 60.600 289.650 ;
        RECT 58.950 286.800 61.050 288.900 ;
        RECT 46.950 283.950 49.050 286.050 ;
        RECT 31.950 277.950 34.050 280.050 ;
        RECT 43.950 277.950 46.050 280.050 ;
        RECT 32.400 247.050 33.450 277.950 ;
        RECT 37.950 260.100 40.050 262.200 ;
        RECT 44.400 261.600 45.450 277.950 ;
        RECT 55.950 274.950 58.050 277.050 ;
        RECT 52.950 262.950 55.050 265.050 ;
        RECT 38.400 259.350 39.600 260.100 ;
        RECT 44.400 259.350 45.600 261.600 ;
        RECT 37.950 256.950 40.050 259.050 ;
        RECT 40.950 256.950 43.050 259.050 ;
        RECT 43.950 256.950 46.050 259.050 ;
        RECT 46.950 256.950 49.050 259.050 ;
        RECT 41.400 255.000 42.600 256.650 ;
        RECT 47.400 255.450 48.600 256.650 ;
        RECT 53.400 255.450 54.450 262.950 ;
        RECT 37.950 250.950 40.050 253.050 ;
        RECT 40.950 250.950 43.050 255.000 ;
        RECT 47.400 254.400 54.450 255.450 ;
        RECT 31.950 244.950 34.050 247.050 ;
        RECT 28.950 217.950 31.050 220.050 ;
        RECT 31.950 215.100 34.050 217.200 ;
        RECT 38.400 216.600 39.450 250.950 ;
        RECT 43.950 223.950 46.050 226.050 ;
        RECT 32.400 214.350 33.600 215.100 ;
        RECT 38.400 214.350 39.600 216.600 ;
        RECT 28.950 211.950 31.050 214.050 ;
        RECT 31.950 211.950 34.050 214.050 ;
        RECT 34.950 211.950 37.050 214.050 ;
        RECT 37.950 211.950 40.050 214.050 ;
        RECT 25.950 208.950 28.050 211.050 ;
        RECT 29.400 209.400 30.600 211.650 ;
        RECT 35.400 209.400 36.600 211.650 ;
        RECT 44.400 210.450 45.450 223.950 ;
        RECT 49.950 215.100 52.050 217.200 ;
        RECT 56.400 216.450 57.450 274.950 ;
        RECT 61.950 271.950 64.050 274.050 ;
        RECT 62.400 261.600 63.450 271.950 ;
        RECT 65.400 271.050 66.450 292.950 ;
        RECT 71.400 292.350 72.600 293.100 ;
        RECT 70.950 289.950 73.050 292.050 ;
        RECT 73.950 289.950 76.050 292.050 ;
        RECT 74.400 288.900 75.600 289.650 ;
        RECT 80.400 288.900 81.450 304.950 ;
        RECT 85.950 293.100 88.050 295.200 ;
        RECT 91.950 293.100 94.050 295.200 ;
        RECT 100.950 293.100 103.050 295.200 ;
        RECT 104.400 295.050 105.450 325.950 ;
        RECT 107.400 304.050 108.450 332.400 ;
        RECT 113.400 325.050 114.450 337.950 ;
        RECT 119.400 337.350 120.600 338.100 ;
        RECT 125.400 337.350 126.600 338.100 ;
        RECT 118.950 334.950 121.050 337.050 ;
        RECT 121.950 334.950 124.050 337.050 ;
        RECT 124.950 334.950 127.050 337.050 ;
        RECT 127.950 334.950 130.050 337.050 ;
        RECT 122.400 333.900 123.600 334.650 ;
        RECT 128.400 333.900 129.600 334.650 ;
        RECT 121.950 331.800 124.050 333.900 ;
        RECT 122.400 328.050 123.450 331.800 ;
        RECT 127.950 328.950 130.050 333.900 ;
        RECT 121.950 325.950 124.050 328.050 ;
        RECT 112.950 322.950 115.050 325.050 ;
        RECT 134.400 322.050 135.450 338.100 ;
        RECT 143.400 337.350 144.600 339.000 ;
        RECT 139.950 334.950 142.050 337.050 ;
        RECT 142.950 334.950 145.050 337.050 ;
        RECT 140.400 333.900 141.600 334.650 ;
        RECT 152.400 333.900 153.450 343.950 ;
        RECT 161.400 339.600 162.450 349.950 ;
        RECT 164.400 346.050 165.450 379.950 ;
        RECT 172.950 371.100 175.050 373.200 ;
        RECT 176.400 372.450 177.450 409.950 ;
        RECT 181.950 409.800 184.050 411.900 ;
        RECT 188.400 411.000 189.600 412.650 ;
        RECT 187.950 406.950 190.050 411.000 ;
        RECT 194.400 406.050 195.450 478.950 ;
        RECT 199.950 466.950 202.050 469.050 ;
        RECT 200.400 451.200 201.450 466.950 ;
        RECT 224.400 466.050 225.450 544.950 ;
        RECT 230.400 528.600 231.450 553.950 ;
        RECT 236.400 532.050 237.450 556.950 ;
        RECT 238.950 535.950 241.050 538.050 ;
        RECT 235.950 529.950 238.050 532.050 ;
        RECT 236.400 528.600 237.450 529.950 ;
        RECT 239.400 529.200 240.450 535.950 ;
        RECT 230.400 526.350 231.600 528.600 ;
        RECT 236.400 526.350 237.600 528.600 ;
        RECT 238.950 527.100 241.050 529.200 ;
        RECT 229.950 523.950 232.050 526.050 ;
        RECT 232.950 523.950 235.050 526.050 ;
        RECT 235.950 523.950 238.050 526.050 ;
        RECT 233.400 521.400 234.600 523.650 ;
        RECT 233.400 511.050 234.450 521.400 ;
        RECT 238.950 520.950 241.050 523.050 ;
        RECT 226.950 508.950 229.050 511.050 ;
        RECT 232.950 508.950 235.050 511.050 ;
        RECT 227.400 481.050 228.450 508.950 ;
        RECT 230.550 501.300 232.650 503.400 ;
        RECT 230.550 488.400 231.750 501.300 ;
        RECT 236.400 495.450 237.600 495.600 ;
        RECT 239.400 495.450 240.450 520.950 ;
        RECT 242.400 520.050 243.450 580.950 ;
        RECT 244.950 574.950 247.050 577.050 ;
        RECT 245.400 567.450 246.450 574.950 ;
        RECT 272.400 573.600 273.450 586.950 ;
        RECT 275.400 580.050 276.450 599.400 ;
        RECT 277.950 598.950 280.050 601.050 ;
        RECT 274.950 577.950 277.050 580.050 ;
        RECT 278.400 574.050 279.450 598.950 ;
        RECT 284.400 589.050 285.450 605.100 ;
        RECT 290.400 604.350 291.600 605.100 ;
        RECT 296.400 604.350 297.600 606.600 ;
        RECT 301.950 605.100 304.050 607.200 ;
        RECT 313.350 606.600 315.450 608.700 ;
        RECT 302.400 604.350 303.600 605.100 ;
        RECT 289.950 601.950 292.050 604.050 ;
        RECT 292.950 601.950 295.050 604.050 ;
        RECT 295.950 601.950 298.050 604.050 ;
        RECT 298.950 601.950 301.050 604.050 ;
        RECT 301.950 601.950 304.050 604.050 ;
        RECT 307.950 601.950 310.050 604.050 ;
        RECT 293.400 599.400 294.600 601.650 ;
        RECT 299.400 599.400 300.600 601.650 ;
        RECT 283.950 586.950 286.050 589.050 ;
        RECT 293.400 586.050 294.450 599.400 ;
        RECT 299.400 595.050 300.450 599.400 ;
        RECT 304.950 598.950 307.050 601.050 ;
        RECT 308.400 599.400 309.600 601.650 ;
        RECT 298.950 592.950 301.050 595.050 ;
        RECT 292.950 583.950 295.050 586.050 ;
        RECT 295.950 577.950 298.050 580.050 ;
        RECT 296.400 574.200 297.450 577.950 ;
        RECT 254.400 573.450 255.600 573.600 ;
        RECT 266.400 573.450 267.600 573.600 ;
        RECT 254.400 572.400 258.450 573.450 ;
        RECT 254.400 571.350 255.600 572.400 ;
        RECT 248.100 568.950 250.200 571.050 ;
        RECT 253.500 568.950 255.600 571.050 ;
        RECT 248.400 567.450 249.600 568.650 ;
        RECT 245.400 566.400 249.600 567.450 ;
        RECT 257.400 547.050 258.450 572.400 ;
        RECT 260.400 572.400 267.600 573.450 ;
        RECT 260.400 556.050 261.450 572.400 ;
        RECT 266.400 571.350 267.600 572.400 ;
        RECT 272.400 571.350 273.600 573.600 ;
        RECT 277.950 571.950 280.050 574.050 ;
        RECT 280.950 572.100 283.050 574.200 ;
        RECT 289.950 572.100 292.050 574.200 ;
        RECT 295.950 572.100 298.050 574.200 ;
        RECT 265.950 568.950 268.050 571.050 ;
        RECT 268.950 568.950 271.050 571.050 ;
        RECT 271.950 568.950 274.050 571.050 ;
        RECT 274.950 568.950 277.050 571.050 ;
        RECT 269.400 566.400 270.600 568.650 ;
        RECT 275.400 566.400 276.600 568.650 ;
        RECT 259.950 553.950 262.050 556.050 ;
        RECT 256.950 544.950 259.050 547.050 ;
        RECT 244.950 538.950 247.050 541.050 ;
        RECT 241.950 517.950 244.050 520.050 ;
        RECT 245.400 502.050 246.450 538.950 ;
        RECT 257.400 538.050 258.450 544.950 ;
        RECT 260.400 544.050 261.450 553.950 ;
        RECT 259.950 541.950 262.050 544.050 ;
        RECT 265.950 541.950 268.050 544.050 ;
        RECT 256.950 535.950 259.050 538.050 ;
        RECT 250.800 532.200 252.900 534.300 ;
        RECT 259.800 532.500 261.900 534.600 ;
        RECT 247.950 527.100 250.050 529.200 ;
        RECT 248.400 526.350 249.600 527.100 ;
        RECT 248.100 523.950 250.200 526.050 ;
        RECT 251.100 519.600 252.000 532.200 ;
        RECT 257.400 529.350 258.600 531.600 ;
        RECT 257.100 526.950 259.200 529.050 ;
        RECT 252.900 525.900 255.000 526.200 ;
        RECT 261.000 525.900 261.900 532.500 ;
        RECT 252.900 525.000 261.900 525.900 ;
        RECT 252.900 524.100 255.000 525.000 ;
        RECT 258.000 523.200 260.100 524.100 ;
        RECT 252.900 522.000 260.100 523.200 ;
        RECT 252.900 521.100 255.000 522.000 ;
        RECT 250.500 517.500 252.600 519.600 ;
        RECT 257.100 518.100 259.200 520.200 ;
        RECT 261.000 519.900 261.900 525.000 ;
        RECT 262.800 523.950 264.900 526.050 ;
        RECT 263.400 522.900 264.600 523.650 ;
        RECT 262.950 520.800 265.050 522.900 ;
        RECT 260.400 517.800 262.500 519.900 ;
        RECT 257.400 515.550 258.600 517.800 ;
        RECT 257.400 508.050 258.450 515.550 ;
        RECT 266.400 511.050 267.450 541.950 ;
        RECT 265.950 508.950 268.050 511.050 ;
        RECT 269.400 508.050 270.450 566.400 ;
        RECT 275.400 556.050 276.450 566.400 ;
        RECT 281.400 559.050 282.450 572.100 ;
        RECT 290.400 571.350 291.600 572.100 ;
        RECT 296.400 571.350 297.600 572.100 ;
        RECT 286.950 568.950 289.050 571.050 ;
        RECT 289.950 568.950 292.050 571.050 ;
        RECT 292.950 568.950 295.050 571.050 ;
        RECT 295.950 568.950 298.050 571.050 ;
        RECT 298.950 568.950 301.050 571.050 ;
        RECT 283.950 565.950 286.050 568.050 ;
        RECT 287.400 567.000 288.600 568.650 ;
        RECT 293.400 567.900 294.600 568.650 ;
        RECT 280.950 556.950 283.050 559.050 ;
        RECT 274.950 553.950 277.050 556.050 ;
        RECT 284.400 553.050 285.450 565.950 ;
        RECT 286.950 562.950 289.050 567.000 ;
        RECT 292.950 565.800 295.050 567.900 ;
        RECT 299.400 566.400 300.600 568.650 ;
        RECT 299.400 562.050 300.450 566.400 ;
        RECT 301.950 562.950 304.050 568.050 ;
        RECT 305.400 564.450 306.450 598.950 ;
        RECT 308.400 595.050 309.450 599.400 ;
        RECT 307.950 592.950 310.050 595.050 ;
        RECT 314.250 593.700 315.450 606.600 ;
        RECT 313.350 591.600 315.450 593.700 ;
        RECT 320.400 586.050 321.450 655.950 ;
        RECT 328.800 646.950 330.900 649.050 ;
        RECT 329.400 645.900 330.600 646.650 ;
        RECT 328.950 643.800 331.050 645.900 ;
        RECT 334.650 638.700 335.850 657.300 ;
        RECT 337.950 655.950 340.050 658.050 ;
        RECT 346.950 650.100 349.050 652.200 ;
        RECT 337.950 646.950 340.050 649.050 ;
        RECT 331.650 637.500 335.850 638.700 ;
        RECT 338.400 644.400 339.600 646.650 ;
        RECT 347.400 646.050 348.450 650.100 ;
        RECT 331.650 636.600 333.750 637.500 ;
        RECT 338.400 633.450 339.450 644.400 ;
        RECT 346.800 643.950 348.900 646.050 ;
        RECT 350.400 645.900 351.450 658.950 ;
        RECT 365.400 652.200 366.450 664.950 ;
        RECT 358.950 650.100 361.050 652.200 ;
        RECT 364.950 650.100 367.050 652.200 ;
        RECT 374.400 651.450 375.450 697.950 ;
        RECT 379.950 683.100 382.050 685.200 ;
        RECT 385.950 684.000 388.050 688.050 ;
        RECT 380.400 682.350 381.600 683.100 ;
        RECT 386.400 682.350 387.600 684.000 ;
        RECT 379.950 679.950 382.050 682.050 ;
        RECT 382.950 679.950 385.050 682.050 ;
        RECT 385.950 679.950 388.050 682.050 ;
        RECT 388.950 679.950 391.050 682.050 ;
        RECT 383.400 677.400 384.600 679.650 ;
        RECT 389.400 677.400 390.600 679.650 ;
        RECT 383.400 673.050 384.450 677.400 ;
        RECT 389.400 673.050 390.450 677.400 ;
        RECT 382.950 670.950 385.050 673.050 ;
        RECT 388.950 670.950 391.050 673.050 ;
        RECT 395.400 670.050 396.450 718.950 ;
        RECT 398.400 715.050 399.450 722.400 ;
        RECT 397.950 712.950 400.050 715.050 ;
        RECT 397.950 700.950 400.050 703.050 ;
        RECT 398.400 691.050 399.450 700.950 ;
        RECT 404.400 697.050 405.450 733.950 ;
        RECT 413.400 729.600 414.450 742.950 ;
        RECT 413.400 727.350 414.600 729.600 ;
        RECT 409.950 724.950 412.050 727.050 ;
        RECT 412.950 724.950 415.050 727.050 ;
        RECT 410.400 723.900 411.600 724.650 ;
        RECT 409.950 721.800 412.050 723.900 ;
        RECT 410.400 718.050 411.450 721.800 ;
        RECT 409.950 715.950 412.050 718.050 ;
        RECT 419.400 715.050 420.450 748.950 ;
        RECT 424.950 728.100 427.050 730.200 ;
        RECT 431.400 729.600 432.450 751.950 ;
        RECT 434.400 736.050 435.450 755.400 ;
        RECT 433.950 733.950 436.050 736.050 ;
        RECT 437.400 733.200 438.450 778.950 ;
        RECT 439.950 769.950 442.050 772.050 ;
        RECT 440.400 754.050 441.450 769.950 ;
        RECT 443.400 763.050 444.450 787.950 ;
        RECT 445.950 771.450 448.050 772.050 ;
        RECT 451.950 771.450 454.050 772.050 ;
        RECT 445.950 770.400 454.050 771.450 ;
        RECT 445.950 769.950 448.050 770.400 ;
        RECT 451.950 769.950 454.050 770.400 ;
        RECT 448.950 766.950 451.050 769.050 ;
        RECT 460.950 766.950 463.050 769.050 ;
        RECT 442.950 760.950 445.050 763.050 ;
        RECT 449.400 762.600 450.450 766.950 ;
        RECT 449.400 760.350 450.600 762.600 ;
        RECT 454.950 761.100 457.050 763.200 ;
        RECT 455.400 760.350 456.600 761.100 ;
        RECT 445.950 757.950 448.050 760.050 ;
        RECT 448.950 757.950 451.050 760.050 ;
        RECT 451.950 757.950 454.050 760.050 ;
        RECT 454.950 757.950 457.050 760.050 ;
        RECT 446.400 755.400 447.600 757.650 ;
        RECT 452.400 756.900 453.600 757.650 ;
        RECT 439.950 751.950 442.050 754.050 ;
        RECT 446.400 742.050 447.450 755.400 ;
        RECT 451.950 754.800 454.050 756.900 ;
        RECT 461.400 745.050 462.450 766.950 ;
        RECT 467.400 762.600 468.450 796.950 ;
        RECT 473.400 787.050 474.450 802.950 ;
        RECT 482.400 801.000 483.600 802.650 ;
        RECT 488.400 801.000 489.600 802.650 ;
        RECT 500.400 801.900 501.600 802.650 ;
        RECT 506.400 801.900 507.600 802.650 ;
        RECT 512.400 801.900 513.450 805.950 ;
        RECT 520.950 802.950 523.050 805.050 ;
        RECT 523.950 802.950 526.050 805.050 ;
        RECT 538.800 802.950 540.900 805.050 ;
        RECT 556.800 802.950 558.900 805.050 ;
        RECT 481.950 796.950 484.050 801.000 ;
        RECT 487.950 796.950 490.050 801.000 ;
        RECT 499.950 799.800 502.050 801.900 ;
        RECT 505.950 799.800 508.050 801.900 ;
        RECT 511.950 799.800 514.050 801.900 ;
        RECT 524.400 800.400 525.600 802.650 ;
        RECT 557.400 801.000 558.600 802.650 ;
        RECT 472.950 784.950 475.050 787.050 ;
        RECT 524.400 784.050 525.450 800.400 ;
        RECT 556.950 796.950 559.050 801.000 ;
        RECT 523.950 781.950 526.050 784.050 ;
        RECT 532.950 781.950 535.050 784.050 ;
        RECT 514.950 778.950 517.050 781.050 ;
        RECT 487.950 775.950 490.050 778.050 ;
        RECT 484.350 771.300 486.450 773.400 ;
        RECT 475.950 766.950 478.050 769.050 ;
        RECT 467.400 760.350 468.600 762.600 ;
        RECT 472.800 761.100 474.900 763.200 ;
        RECT 476.400 763.050 477.450 766.950 ;
        RECT 485.250 764.700 486.450 771.300 ;
        RECT 473.400 760.350 474.600 761.100 ;
        RECT 475.950 760.950 478.050 763.050 ;
        RECT 484.350 762.600 486.450 764.700 ;
        RECT 466.950 757.950 469.050 760.050 ;
        RECT 469.950 757.950 472.050 760.050 ;
        RECT 472.950 757.950 475.050 760.050 ;
        RECT 478.950 757.950 481.050 760.050 ;
        RECT 470.400 756.900 471.600 757.650 ;
        RECT 469.950 754.800 472.050 756.900 ;
        RECT 475.800 754.950 477.900 757.050 ;
        RECT 479.400 756.900 480.600 757.650 ;
        RECT 460.950 742.950 463.050 745.050 ;
        RECT 445.950 739.950 448.050 742.050 ;
        RECT 442.950 733.950 445.050 736.050 ;
        RECT 460.950 733.950 466.050 736.050 ;
        RECT 466.950 733.950 469.050 736.050 ;
        RECT 469.950 733.950 472.050 739.050 ;
        RECT 436.950 731.100 439.050 733.200 ;
        RECT 425.400 727.350 426.600 728.100 ;
        RECT 431.400 727.350 432.600 729.600 ;
        RECT 436.950 727.950 439.050 730.050 ;
        RECT 437.400 727.350 438.600 727.950 ;
        RECT 424.950 724.950 427.050 727.050 ;
        RECT 427.950 724.950 430.050 727.050 ;
        RECT 430.950 724.950 433.050 727.050 ;
        RECT 433.950 724.950 436.050 727.050 ;
        RECT 436.950 724.950 439.050 727.050 ;
        RECT 428.400 723.000 429.600 724.650 ;
        RECT 434.400 723.900 435.600 724.650 ;
        RECT 427.950 718.950 430.050 723.000 ;
        RECT 433.950 721.800 436.050 723.900 ;
        RECT 439.950 721.950 442.050 724.050 ;
        RECT 443.400 723.900 444.450 733.950 ;
        RECT 451.950 728.100 454.050 730.200 ;
        RECT 457.950 728.100 460.050 730.200 ;
        RECT 467.400 730.050 468.450 733.950 ;
        RECT 452.400 727.350 453.600 728.100 ;
        RECT 458.400 727.350 459.600 728.100 ;
        RECT 463.950 727.950 466.050 730.050 ;
        RECT 466.950 727.950 469.050 730.050 ;
        RECT 469.950 728.100 472.050 730.200 ;
        RECT 476.400 730.050 477.450 754.950 ;
        RECT 478.950 754.800 481.050 756.900 ;
        RECT 485.250 749.700 486.450 762.600 ;
        RECT 478.950 745.950 481.050 748.050 ;
        RECT 484.350 747.600 486.450 749.700 ;
        RECT 488.400 748.050 489.450 775.950 ;
        RECT 493.950 769.950 496.050 772.050 ;
        RECT 494.400 762.450 495.450 769.950 ;
        RECT 499.650 769.500 501.750 770.400 ;
        RECT 499.650 768.300 503.850 769.500 ;
        RECT 497.400 762.450 498.600 762.600 ;
        RECT 494.400 761.400 498.600 762.450 ;
        RECT 497.400 760.350 498.600 761.400 ;
        RECT 496.800 757.950 498.900 760.050 ;
        RECT 493.950 748.950 496.050 751.050 ;
        RECT 502.650 749.700 503.850 768.300 ;
        RECT 515.400 763.200 516.450 778.950 ;
        RECT 526.950 775.950 529.050 778.050 ;
        RECT 521.250 769.500 523.350 770.400 ;
        RECT 519.150 768.300 523.350 769.500 ;
        RECT 505.950 761.100 508.050 763.200 ;
        RECT 514.950 761.100 517.050 763.200 ;
        RECT 506.400 760.350 507.600 761.100 ;
        RECT 515.400 760.350 516.600 761.100 ;
        RECT 505.950 757.950 508.050 760.050 ;
        RECT 514.950 757.950 517.050 760.050 ;
        RECT 508.950 754.950 511.050 757.050 ;
        RECT 487.950 745.950 490.050 748.050 ;
        RECT 448.950 724.950 451.050 727.050 ;
        RECT 451.950 724.950 454.050 727.050 ;
        RECT 454.950 724.950 457.050 727.050 ;
        RECT 457.950 724.950 460.050 727.050 ;
        RECT 418.950 712.950 421.050 715.050 ;
        RECT 415.950 706.950 418.050 709.050 ;
        RECT 403.950 694.950 406.050 697.050 ;
        RECT 404.400 692.400 411.450 693.450 ;
        RECT 397.950 688.950 400.050 691.050 ;
        RECT 400.950 688.050 403.050 688.200 ;
        RECT 404.400 688.050 405.450 692.400 ;
        RECT 406.950 688.950 409.050 691.050 ;
        RECT 400.950 686.700 405.450 688.050 ;
        RECT 400.950 686.100 405.000 686.700 ;
        RECT 402.000 685.950 405.000 686.100 ;
        RECT 400.950 682.950 403.050 685.050 ;
        RECT 407.400 684.600 408.450 688.950 ;
        RECT 410.400 688.050 411.450 692.400 ;
        RECT 409.950 685.950 412.050 688.050 ;
        RECT 401.400 682.350 402.600 682.950 ;
        RECT 407.400 682.350 408.600 684.600 ;
        RECT 400.950 679.950 403.050 682.050 ;
        RECT 403.950 679.950 406.050 682.050 ;
        RECT 406.950 679.950 409.050 682.050 ;
        RECT 409.950 679.950 412.050 682.050 ;
        RECT 397.950 676.950 400.050 679.050 ;
        RECT 404.400 677.400 405.600 679.650 ;
        RECT 410.400 678.900 411.600 679.650 ;
        RECT 388.950 667.800 391.050 669.900 ;
        RECT 394.950 667.950 397.050 670.050 ;
        RECT 379.950 658.950 382.050 661.050 ;
        RECT 371.400 650.400 375.450 651.450 ;
        RECT 380.400 651.600 381.450 658.950 ;
        RECT 359.400 649.350 360.600 650.100 ;
        RECT 365.400 649.350 366.600 650.100 ;
        RECT 355.950 646.950 358.050 649.050 ;
        RECT 358.950 646.950 361.050 649.050 ;
        RECT 361.950 646.950 364.050 649.050 ;
        RECT 364.950 646.950 367.050 649.050 ;
        RECT 356.400 645.900 357.600 646.650 ;
        RECT 349.950 643.800 352.050 645.900 ;
        RECT 355.950 643.800 358.050 645.900 ;
        RECT 362.400 644.400 363.600 646.650 ;
        RECT 362.400 642.450 363.450 644.400 ;
        RECT 359.400 641.400 363.450 642.450 ;
        RECT 359.400 634.050 360.450 641.400 ;
        RECT 361.950 634.950 364.050 637.050 ;
        RECT 335.400 632.400 339.450 633.450 ;
        RECT 335.400 628.050 336.450 632.400 ;
        RECT 358.950 631.950 361.050 634.050 ;
        RECT 334.950 625.950 337.050 628.050 ;
        RECT 335.400 619.050 336.450 625.950 ;
        RECT 334.950 616.950 337.050 619.050 ;
        RECT 328.650 613.500 330.750 614.400 ;
        RECT 328.650 612.300 332.850 613.500 ;
        RECT 325.950 605.100 328.050 607.200 ;
        RECT 326.400 604.350 327.600 605.100 ;
        RECT 325.800 601.950 327.900 604.050 ;
        RECT 331.650 593.700 332.850 612.300 ;
        RECT 335.400 606.600 336.450 616.950 ;
        RECT 340.950 613.950 343.050 616.050 ;
        RECT 335.400 604.350 336.600 606.600 ;
        RECT 334.950 601.950 337.050 604.050 ;
        RECT 341.400 600.900 342.450 613.950 ;
        RECT 352.950 605.100 355.050 607.200 ;
        RECT 353.400 604.350 354.600 605.100 ;
        RECT 349.950 601.950 352.050 604.050 ;
        RECT 352.950 601.950 355.050 604.050 ;
        RECT 355.950 601.950 358.050 604.050 ;
        RECT 340.950 598.800 343.050 600.900 ;
        RECT 350.400 599.400 351.600 601.650 ;
        RECT 356.400 599.400 357.600 601.650 ;
        RECT 334.950 595.950 337.050 598.050 ;
        RECT 331.050 591.600 333.150 593.700 ;
        RECT 307.950 583.950 310.050 586.050 ;
        RECT 319.950 583.950 322.050 586.050 ;
        RECT 308.400 574.050 309.450 583.950 ;
        RECT 307.950 571.950 310.050 574.050 ;
        RECT 313.950 572.100 316.050 574.200 ;
        RECT 322.950 572.100 325.050 574.200 ;
        RECT 328.950 572.100 331.050 574.200 ;
        RECT 335.400 573.600 336.450 595.950 ;
        RECT 346.950 592.950 349.050 595.050 ;
        RECT 314.400 571.350 315.600 572.100 ;
        RECT 310.950 568.950 313.050 571.050 ;
        RECT 313.950 568.950 316.050 571.050 ;
        RECT 316.950 568.950 319.050 571.050 ;
        RECT 311.400 567.900 312.600 568.650 ;
        RECT 310.950 565.800 313.050 567.900 ;
        RECT 317.400 566.400 318.600 568.650 ;
        RECT 307.950 564.450 310.050 565.050 ;
        RECT 305.400 563.400 310.050 564.450 ;
        RECT 307.950 562.950 310.050 563.400 ;
        RECT 289.950 559.950 292.050 562.050 ;
        RECT 298.950 559.950 301.050 562.050 ;
        RECT 283.950 550.950 286.050 553.050 ;
        RECT 274.950 527.100 277.050 529.200 ;
        RECT 280.950 527.100 283.050 529.200 ;
        RECT 275.400 526.350 276.600 527.100 ;
        RECT 281.400 526.350 282.600 527.100 ;
        RECT 274.950 523.950 277.050 526.050 ;
        RECT 277.950 523.950 280.050 526.050 ;
        RECT 280.950 523.950 283.050 526.050 ;
        RECT 283.950 523.950 286.050 526.050 ;
        RECT 278.400 522.900 279.600 523.650 ;
        RECT 277.950 517.950 280.050 522.900 ;
        RECT 284.400 521.400 285.600 523.650 ;
        RECT 271.950 508.950 274.050 511.050 ;
        RECT 256.950 505.950 259.050 508.050 ;
        RECT 268.950 505.950 271.050 508.050 ;
        RECT 244.950 499.950 247.050 502.050 ;
        RECT 259.950 499.950 262.050 502.050 ;
        RECT 253.500 497.400 255.600 499.500 ;
        RECT 260.400 499.200 261.600 499.950 ;
        RECT 236.400 494.400 240.450 495.450 ;
        RECT 236.400 493.350 237.600 494.400 ;
        RECT 235.950 490.950 238.050 493.050 ;
        RECT 251.100 490.950 253.200 493.050 ;
        RECT 251.400 489.900 252.600 490.650 ;
        RECT 230.550 486.300 232.650 488.400 ;
        RECT 241.950 487.800 244.050 489.900 ;
        RECT 250.950 487.800 253.050 489.900 ;
        RECT 226.950 478.950 229.050 481.050 ;
        RECT 230.550 479.700 231.750 486.300 ;
        RECT 230.550 477.600 232.650 479.700 ;
        RECT 235.950 475.950 238.050 478.050 ;
        RECT 223.950 463.950 226.050 466.050 ;
        RECT 214.350 459.300 216.450 461.400 ;
        RECT 215.250 452.700 216.450 459.300 ;
        RECT 229.650 457.500 231.750 458.400 ;
        RECT 229.650 456.300 233.850 457.500 ;
        RECT 199.950 449.100 202.050 451.200 ;
        RECT 214.350 450.600 216.450 452.700 ;
        RECT 200.400 448.350 201.600 449.100 ;
        RECT 199.950 445.950 202.050 448.050 ;
        RECT 202.950 445.950 205.050 448.050 ;
        RECT 208.950 445.950 211.050 448.050 ;
        RECT 203.400 443.400 204.600 445.650 ;
        RECT 209.400 443.400 210.600 445.650 ;
        RECT 203.400 436.050 204.450 443.400 ;
        RECT 209.400 436.050 210.450 443.400 ;
        RECT 215.250 437.700 216.450 450.600 ;
        RECT 220.950 448.950 223.050 451.050 ;
        RECT 226.950 449.100 229.050 451.200 ;
        RECT 221.400 439.050 222.450 448.950 ;
        RECT 227.400 448.350 228.600 449.100 ;
        RECT 226.800 445.950 228.900 448.050 ;
        RECT 223.950 439.950 226.050 442.050 ;
        RECT 202.950 433.950 205.050 436.050 ;
        RECT 208.950 433.950 211.050 436.050 ;
        RECT 214.350 435.600 216.450 437.700 ;
        RECT 220.950 436.950 223.050 439.050 ;
        RECT 224.400 436.050 225.450 439.950 ;
        RECT 232.650 437.700 233.850 456.300 ;
        RECT 236.400 450.600 237.450 475.950 ;
        RECT 236.400 448.350 237.600 450.600 ;
        RECT 235.950 445.950 238.050 448.050 ;
        RECT 223.950 433.950 226.050 436.050 ;
        RECT 232.050 435.600 234.150 437.700 ;
        RECT 242.400 430.050 243.450 487.800 ;
        RECT 254.100 484.800 255.000 497.400 ;
        RECT 260.100 496.800 262.200 498.900 ;
        RECT 263.400 497.100 265.500 499.200 ;
        RECT 255.900 495.000 258.000 495.900 ;
        RECT 255.900 493.800 263.100 495.000 ;
        RECT 261.000 492.900 263.100 493.800 ;
        RECT 255.900 492.000 258.000 492.900 ;
        RECT 264.000 492.000 264.900 497.100 ;
        RECT 266.400 495.450 267.600 495.600 ;
        RECT 266.400 494.400 270.450 495.450 ;
        RECT 266.400 493.350 267.600 494.400 ;
        RECT 255.900 491.100 264.900 492.000 ;
        RECT 255.900 490.800 258.000 491.100 ;
        RECT 260.100 487.950 262.200 490.050 ;
        RECT 260.400 485.400 261.600 487.650 ;
        RECT 253.800 482.700 255.900 484.800 ;
        RECT 264.000 484.500 264.900 491.100 ;
        RECT 265.800 490.950 267.900 493.050 ;
        RECT 262.800 482.400 264.900 484.500 ;
        RECT 269.400 484.050 270.450 494.400 ;
        RECT 268.950 481.950 271.050 484.050 ;
        RECT 253.950 466.950 256.050 469.050 ;
        RECT 244.950 460.950 247.050 463.050 ;
        RECT 245.400 444.900 246.450 460.950 ;
        RECT 254.400 450.600 255.450 466.950 ;
        RECT 272.400 460.050 273.450 508.950 ;
        RECT 277.950 505.950 280.050 508.050 ;
        RECT 274.950 493.950 277.050 496.050 ;
        RECT 271.950 457.950 274.050 460.050 ;
        RECT 272.400 450.600 273.450 457.950 ;
        RECT 275.400 457.050 276.450 493.950 ;
        RECT 274.950 454.950 277.050 457.050 ;
        RECT 278.400 451.200 279.450 505.950 ;
        RECT 284.400 505.050 285.450 521.400 ;
        RECT 286.950 520.800 289.050 522.900 ;
        RECT 283.950 502.950 286.050 505.050 ;
        RECT 287.400 501.450 288.450 520.800 ;
        RECT 290.400 514.050 291.450 559.950 ;
        RECT 299.400 547.050 300.450 559.950 ;
        RECT 298.950 544.950 301.050 547.050 ;
        RECT 298.950 527.100 301.050 529.200 ;
        RECT 299.400 526.350 300.600 527.100 ;
        RECT 295.950 523.950 298.050 526.050 ;
        RECT 298.950 523.950 301.050 526.050 ;
        RECT 301.950 523.950 304.050 526.050 ;
        RECT 296.400 521.400 297.600 523.650 ;
        RECT 302.400 522.900 303.600 523.650 ;
        RECT 308.400 523.050 309.450 562.950 ;
        RECT 317.400 562.050 318.450 566.400 ;
        RECT 319.950 565.950 322.050 568.050 ;
        RECT 316.950 559.950 319.050 562.050 ;
        RECT 320.400 556.050 321.450 565.950 ;
        RECT 323.400 562.050 324.450 572.100 ;
        RECT 329.400 571.350 330.600 572.100 ;
        RECT 335.400 571.350 336.600 573.600 ;
        RECT 340.950 571.950 343.050 577.050 ;
        RECT 347.400 574.050 348.450 592.950 ;
        RECT 350.400 589.050 351.450 599.400 ;
        RECT 349.950 586.950 352.050 589.050 ;
        RECT 356.400 583.050 357.450 599.400 ;
        RECT 355.950 580.950 358.050 583.050 ;
        RECT 349.950 576.450 354.000 577.050 ;
        RECT 349.950 574.950 354.450 576.450 ;
        RECT 346.950 571.950 349.050 574.050 ;
        RECT 353.400 573.600 354.450 574.950 ;
        RECT 362.400 574.200 363.450 634.950 ;
        RECT 371.400 616.050 372.450 650.400 ;
        RECT 380.400 649.350 381.600 651.600 ;
        RECT 376.950 646.950 379.050 649.050 ;
        RECT 379.950 646.950 382.050 649.050 ;
        RECT 382.950 646.950 385.050 649.050 ;
        RECT 377.400 645.900 378.600 646.650 ;
        RECT 376.950 643.800 379.050 645.900 ;
        RECT 383.400 644.400 384.600 646.650 ;
        RECT 383.400 642.450 384.450 644.400 ;
        RECT 380.400 641.400 384.450 642.450 ;
        RECT 370.950 613.950 373.050 616.050 ;
        RECT 372.000 609.450 376.050 610.050 ;
        RECT 371.400 607.950 376.050 609.450 ;
        RECT 371.400 606.600 372.450 607.950 ;
        RECT 371.400 604.350 372.600 606.600 ;
        RECT 367.950 601.950 370.050 604.050 ;
        RECT 370.950 601.950 373.050 604.050 ;
        RECT 373.950 601.950 376.050 604.050 ;
        RECT 368.400 600.900 369.600 601.650 ;
        RECT 367.950 595.950 370.050 600.900 ;
        RECT 374.400 599.400 375.600 601.650 ;
        RECT 364.950 586.950 367.050 589.050 ;
        RECT 353.400 571.350 354.600 573.600 ;
        RECT 361.950 572.100 364.050 574.200 ;
        RECT 328.950 568.950 331.050 571.050 ;
        RECT 331.950 568.950 334.050 571.050 ;
        RECT 334.950 568.950 337.050 571.050 ;
        RECT 337.950 568.950 340.050 571.050 ;
        RECT 349.950 568.950 352.050 571.050 ;
        RECT 352.950 568.950 355.050 571.050 ;
        RECT 355.950 568.950 358.050 571.050 ;
        RECT 332.400 566.400 333.600 568.650 ;
        RECT 338.400 567.900 339.600 568.650 ;
        RECT 350.400 567.900 351.600 568.650 ;
        RECT 322.950 559.950 325.050 562.050 ;
        RECT 319.950 553.950 322.050 556.050 ;
        RECT 310.950 550.950 313.050 553.050 ;
        RECT 289.950 511.950 292.050 514.050 ;
        RECT 296.400 508.050 297.450 521.400 ;
        RECT 301.950 520.800 304.050 522.900 ;
        RECT 307.950 520.950 310.050 523.050 ;
        RECT 307.950 511.950 310.050 514.050 ;
        RECT 295.950 505.950 298.050 508.050 ;
        RECT 308.400 507.450 309.450 511.950 ;
        RECT 311.400 511.050 312.450 550.950 ;
        RECT 332.400 541.050 333.450 566.400 ;
        RECT 337.950 565.800 340.050 567.900 ;
        RECT 349.950 565.800 352.050 567.900 ;
        RECT 356.400 566.400 357.600 568.650 ;
        RECT 356.400 562.050 357.450 566.400 ;
        RECT 358.950 562.950 361.050 565.050 ;
        RECT 355.950 559.950 358.050 562.050 ;
        RECT 359.400 544.050 360.450 562.950 ;
        RECT 361.950 550.950 364.050 553.050 ;
        RECT 358.950 541.950 361.050 544.050 ;
        RECT 331.950 538.950 334.050 541.050 ;
        RECT 362.400 538.050 363.450 550.950 ;
        RECT 365.400 547.050 366.450 586.950 ;
        RECT 374.400 577.050 375.450 599.400 ;
        RECT 380.400 577.050 381.450 641.400 ;
        RECT 385.950 622.950 388.050 625.050 ;
        RECT 386.400 606.600 387.450 622.950 ;
        RECT 389.400 610.050 390.450 667.800 ;
        RECT 398.400 667.050 399.450 676.950 ;
        RECT 404.400 673.050 405.450 677.400 ;
        RECT 409.950 676.800 412.050 678.900 ;
        RECT 416.400 678.450 417.450 706.950 ;
        RECT 413.400 677.400 417.450 678.450 ;
        RECT 403.950 670.950 406.050 673.050 ;
        RECT 397.950 664.950 400.050 667.050 ;
        RECT 397.950 658.950 400.050 661.050 ;
        RECT 398.400 651.600 399.450 658.950 ;
        RECT 398.400 649.350 399.600 651.600 ;
        RECT 403.950 650.100 406.050 652.200 ;
        RECT 409.950 650.100 412.050 652.200 ;
        RECT 404.400 649.350 405.600 650.100 ;
        RECT 394.950 646.950 397.050 649.050 ;
        RECT 397.950 646.950 400.050 649.050 ;
        RECT 400.950 646.950 403.050 649.050 ;
        RECT 403.950 646.950 406.050 649.050 ;
        RECT 395.400 644.400 396.600 646.650 ;
        RECT 401.400 644.400 402.600 646.650 ;
        RECT 395.400 640.050 396.450 644.400 ;
        RECT 401.400 642.450 402.450 644.400 ;
        RECT 406.950 643.950 409.050 646.050 ;
        RECT 401.400 641.400 405.450 642.450 ;
        RECT 394.950 637.950 397.050 640.050 ;
        RECT 404.400 631.050 405.450 641.400 ;
        RECT 407.400 634.050 408.450 643.950 ;
        RECT 410.400 643.050 411.450 650.100 ;
        RECT 409.950 640.950 412.050 643.050 ;
        RECT 406.950 631.950 409.050 634.050 ;
        RECT 403.950 628.950 406.050 631.050 ;
        RECT 400.950 625.950 403.050 628.050 ;
        RECT 388.950 607.950 391.050 610.050 ;
        RECT 386.400 604.350 387.600 606.600 ;
        RECT 391.950 606.000 394.050 610.050 ;
        RECT 401.400 607.200 402.450 625.950 ;
        RECT 413.400 622.050 414.450 677.400 ;
        RECT 419.400 652.200 420.450 712.950 ;
        RECT 424.950 703.950 427.050 706.050 ;
        RECT 421.950 694.950 424.050 697.050 ;
        RECT 422.400 661.050 423.450 694.950 ;
        RECT 425.400 694.050 426.450 703.950 ;
        RECT 433.950 700.950 436.050 703.050 ;
        RECT 424.950 691.950 427.050 694.050 ;
        RECT 434.400 691.050 435.450 700.950 ;
        RECT 433.950 688.950 436.050 691.050 ;
        RECT 424.950 684.000 427.050 688.050 ;
        RECT 434.400 684.600 435.450 688.950 ;
        RECT 425.400 682.350 426.600 684.000 ;
        RECT 434.400 682.350 435.600 684.600 ;
        RECT 425.100 679.950 427.200 682.050 ;
        RECT 428.400 679.950 430.500 682.050 ;
        RECT 433.800 679.950 435.900 682.050 ;
        RECT 428.400 678.900 429.600 679.650 ;
        RECT 427.950 676.800 430.050 678.900 ;
        RECT 424.950 667.950 427.050 670.050 ;
        RECT 421.950 658.950 424.050 661.050 ;
        RECT 418.950 650.100 421.050 652.200 ;
        RECT 425.400 651.600 426.450 667.950 ;
        RECT 434.850 657.300 436.950 659.400 ;
        RECT 419.400 649.350 420.600 650.100 ;
        RECT 425.400 649.350 426.600 651.600 ;
        RECT 418.950 646.950 421.050 649.050 ;
        RECT 421.950 646.950 424.050 649.050 ;
        RECT 424.950 646.950 427.050 649.050 ;
        RECT 430.950 646.950 433.050 649.050 ;
        RECT 422.400 644.400 423.600 646.650 ;
        RECT 431.400 645.000 432.600 646.650 ;
        RECT 418.950 640.950 421.050 643.050 ;
        RECT 412.950 619.950 415.050 622.050 ;
        RECT 407.250 613.500 409.350 614.400 ;
        RECT 405.150 612.300 409.350 613.500 ;
        RECT 392.400 604.350 393.600 606.000 ;
        RECT 400.950 605.100 403.050 607.200 ;
        RECT 401.400 604.350 402.600 605.100 ;
        RECT 385.950 601.950 388.050 604.050 ;
        RECT 388.950 601.950 391.050 604.050 ;
        RECT 391.950 601.950 394.050 604.050 ;
        RECT 394.950 601.950 397.050 604.050 ;
        RECT 400.950 601.950 403.050 604.050 ;
        RECT 389.400 600.000 390.600 601.650 ;
        RECT 388.950 595.950 391.050 600.000 ;
        RECT 395.400 599.400 396.600 601.650 ;
        RECT 385.350 579.300 387.450 581.400 ;
        RECT 373.950 574.950 376.050 577.050 ;
        RECT 367.950 572.100 370.050 574.200 ;
        RECT 379.950 573.000 382.050 577.050 ;
        RECT 368.400 571.350 369.600 572.100 ;
        RECT 380.400 571.350 381.600 573.000 ;
        RECT 368.400 568.950 370.500 571.050 ;
        RECT 373.800 568.950 375.900 571.050 ;
        RECT 379.950 568.950 382.050 571.050 ;
        RECT 374.400 567.000 375.600 568.650 ;
        RECT 373.950 562.950 376.050 567.000 ;
        RECT 386.250 566.400 387.450 579.300 ;
        RECT 395.400 573.450 396.450 599.400 ;
        RECT 405.150 593.700 406.350 612.300 ;
        RECT 412.950 610.950 415.050 613.050 ;
        RECT 410.400 606.450 411.600 606.600 ;
        RECT 413.400 606.450 414.450 610.950 ;
        RECT 410.400 605.400 414.450 606.450 ;
        RECT 410.400 604.350 411.600 605.400 ;
        RECT 415.950 604.950 418.050 607.050 ;
        RECT 410.100 601.950 412.200 604.050 ;
        RECT 404.850 591.600 406.950 593.700 ;
        RECT 403.050 579.300 405.150 581.400 ;
        RECT 392.400 572.400 396.450 573.450 ;
        RECT 392.400 567.900 393.450 572.400 ;
        RECT 397.800 568.950 399.900 571.050 ;
        RECT 398.400 567.900 399.600 568.650 ;
        RECT 385.350 564.300 387.450 566.400 ;
        RECT 391.950 565.800 394.050 567.900 ;
        RECT 397.950 565.800 400.050 567.900 ;
        RECT 386.250 557.700 387.450 564.300 ;
        RECT 403.650 560.700 404.850 579.300 ;
        RECT 416.400 577.050 417.450 604.950 ;
        RECT 419.400 601.050 420.450 640.950 ;
        RECT 422.400 634.050 423.450 644.400 ;
        RECT 430.950 640.950 433.050 645.000 ;
        RECT 435.150 638.700 436.350 657.300 ;
        RECT 440.400 655.050 441.450 721.950 ;
        RECT 442.950 721.800 445.050 723.900 ;
        RECT 449.400 722.400 450.600 724.650 ;
        RECT 455.400 723.900 456.600 724.650 ;
        RECT 449.400 721.050 450.450 722.400 ;
        RECT 454.950 721.800 457.050 723.900 ;
        RECT 448.950 718.950 451.050 721.050 ;
        RECT 445.950 709.950 448.050 712.050 ;
        RECT 442.950 697.950 445.050 700.050 ;
        RECT 443.400 661.050 444.450 697.950 ;
        RECT 446.400 684.600 447.450 709.950 ;
        RECT 449.400 688.050 450.450 718.950 ;
        RECT 455.400 718.050 456.450 721.800 ;
        RECT 454.950 715.950 457.050 718.050 ;
        RECT 464.400 706.050 465.450 727.950 ;
        RECT 470.400 727.350 471.600 728.100 ;
        RECT 475.950 727.950 478.050 730.050 ;
        RECT 469.950 724.950 472.050 727.050 ;
        RECT 472.950 724.950 475.050 727.050 ;
        RECT 466.950 718.950 469.050 724.050 ;
        RECT 473.400 723.000 474.600 724.650 ;
        RECT 472.950 718.950 475.050 723.000 ;
        RECT 475.950 721.950 478.050 724.050 ;
        RECT 476.400 712.050 477.450 721.950 ;
        RECT 475.950 709.950 478.050 712.050 ;
        RECT 463.950 703.950 466.050 706.050 ;
        RECT 448.950 685.950 451.050 688.050 ;
        RECT 454.950 685.950 457.050 688.050 ;
        RECT 446.400 682.350 447.600 684.600 ;
        RECT 446.100 679.950 448.200 682.050 ;
        RECT 451.500 679.950 453.600 682.050 ;
        RECT 452.400 677.400 453.600 679.650 ;
        RECT 452.400 675.450 453.450 677.400 ;
        RECT 449.400 674.400 453.450 675.450 ;
        RECT 442.950 658.950 445.050 661.050 ;
        RECT 439.950 652.950 442.050 655.050 ;
        RECT 445.950 652.950 448.050 655.050 ;
        RECT 440.100 646.950 442.200 649.050 ;
        RECT 440.400 645.450 441.600 646.650 ;
        RECT 440.400 644.400 444.450 645.450 ;
        RECT 435.150 637.500 439.350 638.700 ;
        RECT 437.250 636.600 439.350 637.500 ;
        RECT 421.950 631.950 424.050 634.050 ;
        RECT 436.950 628.950 439.050 631.050 ;
        RECT 422.550 615.300 424.650 617.400 ;
        RECT 422.550 608.700 423.750 615.300 ;
        RECT 433.950 610.950 436.050 613.050 ;
        RECT 422.550 606.600 424.650 608.700 ;
        RECT 418.950 598.950 421.050 601.050 ;
        RECT 422.550 593.700 423.750 606.600 ;
        RECT 427.950 601.950 430.050 604.050 ;
        RECT 428.400 600.900 429.600 601.650 ;
        RECT 427.950 598.800 430.050 600.900 ;
        RECT 422.550 591.600 424.650 593.700 ;
        RECT 419.850 579.300 421.950 581.400 ;
        RECT 415.950 574.950 418.050 577.050 ;
        RECT 406.950 568.950 409.050 571.050 ;
        RECT 415.950 568.950 418.050 571.050 ;
        RECT 407.400 567.900 408.600 568.650 ;
        RECT 416.400 567.900 417.600 568.650 ;
        RECT 406.950 565.800 409.050 567.900 ;
        RECT 415.950 565.800 418.050 567.900 ;
        RECT 400.650 559.500 404.850 560.700 ;
        RECT 420.150 560.700 421.350 579.300 ;
        RECT 428.400 573.450 429.450 598.800 ;
        RECT 434.400 583.050 435.450 610.950 ;
        RECT 437.400 601.050 438.450 628.950 ;
        RECT 443.400 616.050 444.450 644.400 ;
        RECT 446.400 643.050 447.450 652.950 ;
        RECT 445.950 640.950 448.050 643.050 ;
        RECT 449.400 637.050 450.450 674.400 ;
        RECT 455.400 667.050 456.450 685.950 ;
        RECT 464.400 685.200 465.450 703.950 ;
        RECT 479.400 688.050 480.450 745.950 ;
        RECT 481.950 736.950 484.050 739.050 ;
        RECT 482.400 724.050 483.450 736.950 ;
        RECT 487.950 733.950 490.050 736.050 ;
        RECT 488.400 730.200 489.450 733.950 ;
        RECT 494.400 733.050 495.450 748.950 ;
        RECT 502.050 747.600 504.150 749.700 ;
        RECT 493.950 730.950 496.050 733.050 ;
        RECT 499.950 730.950 502.050 733.050 ;
        RECT 487.950 728.100 490.050 730.200 ;
        RECT 494.400 729.600 495.450 730.950 ;
        RECT 488.400 727.350 489.600 728.100 ;
        RECT 494.400 727.350 495.600 729.600 ;
        RECT 487.950 724.950 490.050 727.050 ;
        RECT 490.950 724.950 493.050 727.050 ;
        RECT 493.950 724.950 496.050 727.050 ;
        RECT 481.950 721.950 484.050 724.050 ;
        RECT 491.400 723.900 492.600 724.650 ;
        RECT 490.950 721.800 493.050 723.900 ;
        RECT 500.400 723.450 501.450 730.950 ;
        RECT 509.400 729.600 510.450 754.950 ;
        RECT 519.150 749.700 520.350 768.300 ;
        RECT 527.400 765.450 528.450 775.950 ;
        RECT 524.400 764.400 528.450 765.450 ;
        RECT 524.400 762.600 525.450 764.400 ;
        RECT 524.400 760.350 525.600 762.600 ;
        RECT 524.100 757.950 526.200 760.050 ;
        RECT 518.850 747.600 520.950 749.700 ;
        RECT 529.950 733.950 532.050 736.050 ;
        RECT 509.400 727.350 510.600 729.600 ;
        RECT 514.950 728.100 517.050 730.200 ;
        RECT 530.400 729.600 531.450 733.950 ;
        RECT 533.400 733.050 534.450 781.950 ;
        RECT 557.400 781.050 558.450 796.950 ;
        RECT 560.400 796.050 561.450 805.950 ;
        RECT 566.400 802.050 567.450 806.100 ;
        RECT 575.400 805.350 576.600 807.600 ;
        RECT 583.950 806.100 586.050 808.200 ;
        RECT 584.400 805.350 585.600 806.100 ;
        RECT 571.950 802.950 574.050 805.050 ;
        RECT 574.950 802.950 577.050 805.050 ;
        RECT 577.950 802.950 580.050 805.050 ;
        RECT 583.950 802.950 586.050 805.050 ;
        RECT 565.950 799.950 568.050 802.050 ;
        RECT 572.400 801.900 573.600 802.650 ;
        RECT 571.950 799.800 574.050 801.900 ;
        RECT 578.400 800.400 579.600 802.650 ;
        RECT 590.250 800.400 591.450 813.300 ;
        RECT 595.950 811.950 598.050 814.050 ;
        RECT 607.050 813.300 609.150 815.400 ;
        RECT 640.350 813.300 642.450 815.400 ;
        RECT 658.050 813.300 660.150 815.400 ;
        RECT 592.950 802.950 595.050 805.050 ;
        RECT 559.950 793.950 562.050 796.050 ;
        RECT 571.950 790.950 574.050 793.050 ;
        RECT 556.950 778.950 559.050 781.050 ;
        RECT 565.950 778.950 568.050 781.050 ;
        RECT 536.550 771.300 538.650 773.400 ;
        RECT 536.550 764.700 537.750 771.300 ;
        RECT 536.550 762.600 538.650 764.700 ;
        RECT 536.550 749.700 537.750 762.600 ;
        RECT 550.950 761.100 553.050 763.200 ;
        RECT 556.950 761.100 559.050 763.200 ;
        RECT 541.950 757.950 544.050 760.050 ;
        RECT 542.400 755.400 543.600 757.650 ;
        RECT 551.400 756.450 552.450 761.100 ;
        RECT 557.400 760.350 558.600 761.100 ;
        RECT 556.950 757.950 559.050 760.050 ;
        RECT 559.950 757.950 562.050 760.050 ;
        RECT 551.400 755.400 555.450 756.450 ;
        RECT 542.400 751.050 543.450 755.400 ;
        RECT 536.550 747.600 538.650 749.700 ;
        RECT 541.950 748.950 544.050 751.050 ;
        RECT 542.400 745.050 543.450 748.950 ;
        RECT 541.950 742.950 544.050 745.050 ;
        RECT 532.950 730.950 535.050 733.050 ;
        RECT 538.800 730.950 540.900 733.050 ;
        RECT 515.400 727.350 516.600 728.100 ;
        RECT 530.400 727.350 531.600 729.600 ;
        RECT 505.950 724.950 508.050 727.050 ;
        RECT 508.950 724.950 511.050 727.050 ;
        RECT 511.950 724.950 514.050 727.050 ;
        RECT 514.950 724.950 517.050 727.050 ;
        RECT 520.950 724.950 523.050 727.050 ;
        RECT 526.950 724.950 529.050 727.050 ;
        RECT 529.950 724.950 532.050 727.050 ;
        RECT 532.950 724.950 535.050 727.050 ;
        RECT 506.400 723.450 507.600 724.650 ;
        RECT 512.400 723.900 513.600 724.650 ;
        RECT 500.400 722.400 507.600 723.450 ;
        RECT 511.950 721.800 514.050 723.900 ;
        RECT 508.950 709.950 511.050 712.050 ;
        RECT 496.950 700.950 499.050 703.050 ;
        RECT 490.950 694.950 493.050 697.050 ;
        RECT 478.950 685.950 481.050 688.050 ;
        RECT 463.950 683.100 466.050 685.200 ;
        RECT 469.950 683.100 472.050 685.200 ;
        RECT 477.000 684.900 480.000 685.050 ;
        RECT 477.000 684.600 481.050 684.900 ;
        RECT 470.400 682.350 471.600 683.100 ;
        RECT 476.400 682.950 481.050 684.600 ;
        RECT 476.400 682.350 477.600 682.950 ;
        RECT 478.950 682.800 481.050 682.950 ;
        RECT 491.400 684.600 492.450 694.950 ;
        RECT 491.400 682.350 492.600 684.600 ;
        RECT 466.950 679.950 469.050 682.050 ;
        RECT 469.950 679.950 472.050 682.050 ;
        RECT 472.950 679.950 475.050 682.050 ;
        RECT 475.950 679.950 478.050 682.050 ;
        RECT 487.950 679.950 490.050 682.050 ;
        RECT 490.950 679.950 493.050 682.050 ;
        RECT 457.950 676.800 460.050 678.900 ;
        RECT 467.400 677.400 468.600 679.650 ;
        RECT 473.400 678.900 474.600 679.650 ;
        RECT 454.950 664.950 457.050 667.050 ;
        RECT 458.400 664.050 459.450 676.800 ;
        RECT 467.400 667.050 468.450 677.400 ;
        RECT 472.950 676.800 475.050 678.900 ;
        RECT 478.950 675.450 481.050 679.050 ;
        RECT 476.400 675.000 481.050 675.450 ;
        RECT 476.400 674.400 480.450 675.000 ;
        RECT 466.950 664.950 469.050 667.050 ;
        RECT 457.950 661.950 460.050 664.050 ;
        RECT 452.550 657.300 454.650 659.400 ;
        RECT 452.550 644.400 453.750 657.300 ;
        RECT 458.400 651.450 459.600 651.600 ;
        RECT 458.400 650.400 465.450 651.450 ;
        RECT 458.400 649.350 459.600 650.400 ;
        RECT 457.950 646.950 460.050 649.050 ;
        RECT 452.550 642.300 454.650 644.400 ;
        RECT 448.950 634.950 451.050 637.050 ;
        RECT 452.550 635.700 453.750 642.300 ;
        RECT 449.400 631.050 450.450 634.950 ;
        RECT 452.550 633.600 454.650 635.700 ;
        RECT 448.950 628.950 451.050 631.050 ;
        RECT 464.400 628.050 465.450 650.400 ;
        RECT 467.400 643.050 468.450 664.950 ;
        RECT 476.400 651.600 477.450 674.400 ;
        RECT 497.400 673.050 498.450 700.950 ;
        RECT 509.400 685.200 510.450 709.950 ;
        RECT 521.400 706.050 522.450 724.950 ;
        RECT 527.400 723.000 528.600 724.650 ;
        RECT 533.400 724.050 534.600 724.650 ;
        RECT 526.950 718.950 529.050 723.000 ;
        RECT 533.400 722.400 538.050 724.050 ;
        RECT 534.000 721.950 538.050 722.400 ;
        RECT 520.950 703.950 523.050 706.050 ;
        RECT 539.400 700.050 540.450 730.950 ;
        RECT 541.950 727.950 544.050 733.050 ;
        RECT 554.400 730.200 555.450 755.400 ;
        RECT 560.400 755.400 561.600 757.650 ;
        RECT 560.400 745.050 561.450 755.400 ;
        RECT 559.950 742.950 562.050 745.050 ;
        RECT 559.950 733.950 562.050 736.050 ;
        RECT 547.950 728.100 550.050 730.200 ;
        RECT 553.950 728.100 556.050 730.200 ;
        RECT 548.400 727.350 549.600 728.100 ;
        RECT 554.400 727.350 555.600 728.100 ;
        RECT 544.950 724.950 547.050 727.050 ;
        RECT 547.950 724.950 550.050 727.050 ;
        RECT 550.950 724.950 553.050 727.050 ;
        RECT 553.950 724.950 556.050 727.050 ;
        RECT 545.400 723.900 546.600 724.650 ;
        RECT 544.950 721.800 547.050 723.900 ;
        RECT 551.400 722.400 552.600 724.650 ;
        RECT 551.400 718.050 552.450 722.400 ;
        RECT 550.950 715.950 553.050 718.050 ;
        RECT 553.950 700.950 556.050 703.050 ;
        RECT 538.950 697.950 541.050 700.050 ;
        RECT 550.950 697.950 553.050 700.050 ;
        RECT 517.950 694.950 520.050 697.050 ;
        RECT 529.950 694.950 532.050 697.050 ;
        RECT 514.950 688.950 517.050 691.050 ;
        RECT 502.950 683.100 505.050 685.200 ;
        RECT 508.950 683.100 511.050 685.200 ;
        RECT 503.400 682.350 504.600 683.100 ;
        RECT 509.400 682.350 510.600 683.100 ;
        RECT 502.950 679.950 505.050 682.050 ;
        RECT 505.950 679.950 508.050 682.050 ;
        RECT 508.950 679.950 511.050 682.050 ;
        RECT 499.950 676.950 502.050 679.050 ;
        RECT 506.400 678.900 507.600 679.650 ;
        RECT 496.950 670.950 499.050 673.050 ;
        RECT 500.400 670.050 501.450 676.950 ;
        RECT 505.950 676.800 508.050 678.900 ;
        RECT 511.950 673.950 514.050 679.050 ;
        RECT 499.950 667.950 502.050 670.050 ;
        RECT 515.400 664.050 516.450 688.950 ;
        RECT 514.950 661.950 517.050 664.050 ;
        RECT 484.950 658.950 487.050 661.050 ;
        RECT 493.950 658.950 496.050 661.050 ;
        RECT 476.400 649.350 477.600 651.600 ;
        RECT 472.950 646.950 475.050 649.050 ;
        RECT 475.950 646.950 478.050 649.050 ;
        RECT 478.950 646.950 481.050 649.050 ;
        RECT 473.400 645.000 474.600 646.650 ;
        RECT 466.950 640.950 469.050 643.050 ;
        RECT 472.950 640.950 475.050 645.000 ;
        RECT 479.400 644.400 480.600 646.650 ;
        RECT 479.400 628.050 480.450 644.400 ;
        RECT 463.950 625.950 466.050 628.050 ;
        RECT 478.950 625.950 481.050 628.050 ;
        RECT 475.950 619.950 478.050 622.050 ;
        RECT 442.950 613.950 445.050 616.050 ;
        RECT 442.950 605.100 445.050 610.050 ;
        RECT 448.950 605.100 451.050 607.200 ;
        RECT 457.950 605.100 460.050 607.200 ;
        RECT 460.950 606.600 465.000 607.050 ;
        RECT 443.400 604.350 444.600 605.100 ;
        RECT 449.400 604.350 450.600 605.100 ;
        RECT 442.950 601.950 445.050 604.050 ;
        RECT 445.950 601.950 448.050 604.050 ;
        RECT 448.950 601.950 451.050 604.050 ;
        RECT 451.950 601.950 454.050 604.050 ;
        RECT 436.950 598.950 439.050 601.050 ;
        RECT 446.400 600.900 447.600 601.650 ;
        RECT 452.400 600.900 453.600 601.650 ;
        RECT 445.950 598.800 448.050 600.900 ;
        RECT 451.950 598.800 454.050 600.900 ;
        RECT 458.400 586.050 459.450 605.100 ;
        RECT 460.950 604.950 465.600 606.600 ;
        RECT 469.950 606.000 472.050 610.050 ;
        RECT 476.400 607.050 477.450 619.950 ;
        RECT 478.950 613.950 481.050 616.050 ;
        RECT 464.400 604.350 465.600 604.950 ;
        RECT 470.400 604.350 471.600 606.000 ;
        RECT 475.950 604.950 478.050 607.050 ;
        RECT 463.950 601.950 466.050 604.050 ;
        RECT 466.950 601.950 469.050 604.050 ;
        RECT 469.950 601.950 472.050 604.050 ;
        RECT 472.950 601.950 475.050 604.050 ;
        RECT 460.950 598.950 463.050 601.050 ;
        RECT 467.400 600.900 468.600 601.650 ;
        RECT 457.950 583.950 460.050 586.050 ;
        RECT 433.950 580.950 436.050 583.050 ;
        RECT 428.400 572.400 432.450 573.450 ;
        RECT 425.100 568.950 427.200 571.050 ;
        RECT 425.400 567.900 426.600 568.650 ;
        RECT 431.400 567.900 432.450 572.400 ;
        RECT 424.950 565.800 427.050 567.900 ;
        RECT 430.950 565.800 433.050 567.900 ;
        RECT 420.150 559.500 424.350 560.700 ;
        RECT 400.650 558.600 402.750 559.500 ;
        RECT 422.250 558.600 424.350 559.500 ;
        RECT 385.350 555.600 387.450 557.700 ;
        RECT 364.950 544.950 367.050 547.050 ;
        RECT 434.400 538.050 435.450 580.950 ;
        RECT 437.550 579.300 439.650 581.400 ;
        RECT 451.950 580.950 454.050 583.050 ;
        RECT 437.550 566.400 438.750 579.300 ;
        RECT 442.950 572.100 445.050 574.200 ;
        RECT 452.400 573.600 453.450 580.950 ;
        RECT 457.350 579.300 459.450 581.400 ;
        RECT 443.400 571.350 444.600 572.100 ;
        RECT 452.400 571.350 453.600 573.600 ;
        RECT 442.950 568.950 445.050 571.050 ;
        RECT 451.950 568.950 454.050 571.050 ;
        RECT 458.250 566.400 459.450 579.300 ;
        RECT 461.400 574.200 462.450 598.950 ;
        RECT 466.950 598.800 469.050 600.900 ;
        RECT 473.400 599.400 474.600 601.650 ;
        RECT 479.400 601.050 480.450 613.950 ;
        RECT 485.400 610.050 486.450 658.950 ;
        RECT 494.400 651.600 495.450 658.950 ;
        RECT 509.850 657.300 511.950 659.400 ;
        RECT 494.400 649.350 495.600 651.600 ;
        RECT 499.950 650.100 502.050 652.200 ;
        RECT 500.400 649.350 501.600 650.100 ;
        RECT 490.950 646.950 493.050 649.050 ;
        RECT 493.950 646.950 496.050 649.050 ;
        RECT 496.950 646.950 499.050 649.050 ;
        RECT 499.950 646.950 502.050 649.050 ;
        RECT 505.950 646.950 508.050 649.050 ;
        RECT 491.400 644.400 492.600 646.650 ;
        RECT 497.400 644.400 498.600 646.650 ;
        RECT 506.400 645.000 507.600 646.650 ;
        RECT 491.400 637.050 492.450 644.400 ;
        RECT 497.400 642.450 498.450 644.400 ;
        RECT 494.400 641.400 498.450 642.450 ;
        RECT 490.950 634.950 493.050 637.050 ;
        RECT 494.400 622.050 495.450 641.400 ;
        RECT 505.950 640.950 508.050 645.000 ;
        RECT 510.150 638.700 511.350 657.300 ;
        RECT 518.400 651.450 519.450 694.950 ;
        RECT 520.950 684.600 525.000 685.050 ;
        RECT 530.400 684.600 531.450 694.950 ;
        RECT 538.950 691.950 541.050 694.050 ;
        RECT 544.350 693.300 546.450 695.400 ;
        RECT 539.400 688.050 540.450 691.950 ;
        RECT 538.950 685.950 541.050 688.050 ;
        RECT 545.250 686.700 546.450 693.300 ;
        RECT 547.950 688.950 550.050 691.050 ;
        RECT 544.350 684.600 546.450 686.700 ;
        RECT 520.950 682.950 525.600 684.600 ;
        RECT 524.400 682.350 525.600 682.950 ;
        RECT 530.400 682.350 531.600 684.600 ;
        RECT 523.950 679.950 526.050 682.050 ;
        RECT 526.950 679.950 529.050 682.050 ;
        RECT 529.950 679.950 532.050 682.050 ;
        RECT 532.950 679.950 535.050 682.050 ;
        RECT 538.950 679.950 541.050 682.050 ;
        RECT 527.400 677.400 528.600 679.650 ;
        RECT 533.400 678.900 534.600 679.650 ;
        RECT 527.400 673.050 528.450 677.400 ;
        RECT 532.950 676.800 535.050 678.900 ;
        RECT 539.400 677.400 540.600 679.650 ;
        RECT 526.950 670.950 529.050 673.050 ;
        RECT 539.400 670.050 540.450 677.400 ;
        RECT 545.250 671.700 546.450 684.600 ;
        RECT 548.400 679.050 549.450 688.950 ;
        RECT 547.950 676.950 550.050 679.050 ;
        RECT 538.950 667.950 541.050 670.050 ;
        RECT 544.350 669.600 546.450 671.700 ;
        RECT 547.950 661.950 550.050 664.050 ;
        RECT 527.550 657.300 529.650 659.400 ;
        RECT 518.400 650.400 522.450 651.450 ;
        RECT 515.100 646.950 517.200 649.050 ;
        RECT 515.400 645.900 516.600 646.650 ;
        RECT 514.950 643.800 517.050 645.900 ;
        RECT 510.150 637.500 514.350 638.700 ;
        RECT 499.950 634.950 502.050 637.050 ;
        RECT 512.250 636.600 514.350 637.500 ;
        RECT 496.950 628.950 499.050 631.050 ;
        RECT 493.950 619.950 496.050 622.050 ;
        RECT 487.950 613.950 490.050 616.050 ;
        RECT 484.950 607.950 487.050 610.050 ;
        RECT 488.400 606.600 489.450 613.950 ;
        RECT 488.400 604.350 489.600 606.600 ;
        RECT 493.950 606.000 496.050 610.050 ;
        RECT 497.400 607.050 498.450 628.950 ;
        RECT 494.400 604.350 495.600 606.000 ;
        RECT 496.950 604.950 499.050 607.050 ;
        RECT 484.950 601.950 487.050 604.050 ;
        RECT 487.950 601.950 490.050 604.050 ;
        RECT 490.950 601.950 493.050 604.050 ;
        RECT 493.950 601.950 496.050 604.050 ;
        RECT 473.400 595.050 474.450 599.400 ;
        RECT 478.950 598.950 481.050 601.050 ;
        RECT 485.400 599.400 486.600 601.650 ;
        RECT 491.400 600.900 492.600 601.650 ;
        RECT 472.950 592.950 475.050 595.050 ;
        RECT 485.400 592.050 486.450 599.400 ;
        RECT 490.950 598.800 493.050 600.900 ;
        RECT 493.950 595.950 496.050 598.050 ;
        RECT 484.950 589.950 487.050 592.050 ;
        RECT 463.950 580.950 466.050 583.050 ;
        RECT 460.950 572.100 463.050 574.200 ;
        RECT 461.400 567.900 462.450 572.100 ;
        RECT 437.550 564.300 439.650 566.400 ;
        RECT 457.350 564.300 459.450 566.400 ;
        RECT 460.950 565.800 463.050 567.900 ;
        RECT 437.550 557.700 438.750 564.300 ;
        RECT 458.250 557.700 459.450 564.300 ;
        RECT 437.550 555.600 439.650 557.700 ;
        RECT 457.350 555.600 459.450 557.700 ;
        RECT 464.400 553.050 465.450 580.950 ;
        RECT 475.050 579.300 477.150 581.400 ;
        RECT 469.800 568.950 471.900 571.050 ;
        RECT 470.400 567.900 471.600 568.650 ;
        RECT 469.950 565.800 472.050 567.900 ;
        RECT 475.650 560.700 476.850 579.300 ;
        RECT 494.400 573.600 495.450 595.950 ;
        RECT 500.400 592.050 501.450 634.950 ;
        RECT 505.950 625.950 508.050 628.050 ;
        RECT 502.950 604.950 505.050 610.050 ;
        RECT 506.400 606.600 507.450 625.950 ;
        RECT 511.950 613.950 514.050 616.050 ;
        RECT 512.400 610.050 513.450 613.950 ;
        RECT 521.400 613.050 522.450 650.400 ;
        RECT 527.550 644.400 528.750 657.300 ;
        RECT 538.950 652.950 541.050 655.050 ;
        RECT 532.950 650.100 535.050 652.200 ;
        RECT 533.400 649.350 534.600 650.100 ;
        RECT 532.950 646.950 535.050 649.050 ;
        RECT 527.550 642.300 529.650 644.400 ;
        RECT 527.550 635.700 528.750 642.300 ;
        RECT 539.400 637.050 540.450 652.950 ;
        RECT 548.400 651.600 549.450 661.950 ;
        RECT 551.400 655.050 552.450 697.950 ;
        RECT 554.400 684.450 555.450 700.950 ;
        RECT 560.400 697.050 561.450 733.950 ;
        RECT 566.400 733.050 567.450 778.950 ;
        RECT 572.400 763.050 573.450 790.950 ;
        RECT 578.400 781.050 579.450 800.400 ;
        RECT 589.350 798.300 591.450 800.400 ;
        RECT 590.250 791.700 591.450 798.300 ;
        RECT 593.400 796.050 594.450 802.950 ;
        RECT 592.950 793.950 595.050 796.050 ;
        RECT 589.350 789.600 591.450 791.700 ;
        RECT 577.950 778.950 580.050 781.050 ;
        RECT 596.400 769.050 597.450 811.950 ;
        RECT 601.800 802.950 603.900 805.050 ;
        RECT 602.400 801.450 603.600 802.650 ;
        RECT 599.400 800.400 603.600 801.450 ;
        RECT 599.400 793.050 600.450 800.400 ;
        RECT 607.650 794.700 608.850 813.300 ;
        RECT 628.950 806.100 631.050 808.200 ;
        RECT 634.950 806.100 637.050 808.200 ;
        RECT 629.400 805.350 630.600 806.100 ;
        RECT 635.400 805.350 636.600 806.100 ;
        RECT 610.950 802.950 613.050 805.050 ;
        RECT 625.950 802.950 628.050 805.050 ;
        RECT 628.950 802.950 631.050 805.050 ;
        RECT 634.950 802.950 637.050 805.050 ;
        RECT 611.400 801.000 612.600 802.650 ;
        RECT 626.400 801.900 627.600 802.650 ;
        RECT 610.950 796.950 613.050 801.000 ;
        RECT 625.950 799.800 628.050 801.900 ;
        RECT 641.250 800.400 642.450 813.300 ;
        RECT 646.950 808.950 649.050 811.050 ;
        RECT 647.400 801.900 648.450 808.950 ;
        RECT 652.800 802.950 654.900 805.050 ;
        RECT 653.400 801.900 654.600 802.650 ;
        RECT 640.350 798.300 642.450 800.400 ;
        RECT 646.950 799.800 649.050 801.900 ;
        RECT 652.950 799.800 655.050 801.900 ;
        RECT 604.650 793.500 608.850 794.700 ;
        RECT 598.950 790.950 601.050 793.050 ;
        RECT 604.650 792.600 606.750 793.500 ;
        RECT 641.250 791.700 642.450 798.300 ;
        RECT 658.650 794.700 659.850 813.300 ;
        RECT 817.950 811.950 820.050 814.050 ;
        RECT 853.950 811.950 856.050 814.050 ;
        RECT 670.950 808.950 673.050 811.050 ;
        RECT 661.950 802.950 664.050 805.050 ;
        RECT 667.950 802.950 670.050 805.050 ;
        RECT 662.400 801.000 663.600 802.650 ;
        RECT 661.950 796.950 664.050 801.000 ;
        RECT 668.400 796.050 669.450 802.950 ;
        RECT 671.400 802.050 672.450 808.950 ;
        RECT 700.950 806.100 703.050 808.200 ;
        RECT 709.950 806.100 712.050 808.200 ;
        RECT 715.950 806.100 718.050 808.200 ;
        RECT 730.950 806.100 733.050 808.200 ;
        RECT 736.950 806.100 739.050 808.200 ;
        RECT 745.950 806.100 748.050 808.200 ;
        RECT 757.950 806.100 760.050 808.200 ;
        RECT 769.950 806.100 772.050 808.200 ;
        RECT 775.950 806.100 778.050 808.200 ;
        RECT 781.950 806.100 784.050 808.200 ;
        RECT 818.400 807.600 819.450 811.950 ;
        RECT 800.400 807.450 801.600 807.600 ;
        RECT 800.400 806.400 807.450 807.450 ;
        RECT 676.950 802.950 679.050 805.050 ;
        RECT 679.950 802.950 682.050 805.050 ;
        RECT 691.950 802.950 694.050 805.050 ;
        RECT 694.950 802.950 697.050 805.050 ;
        RECT 670.950 799.950 673.050 802.050 ;
        RECT 677.400 800.400 678.600 802.650 ;
        RECT 692.400 800.400 693.600 802.650 ;
        RECT 655.650 793.500 659.850 794.700 ;
        RECT 667.950 793.950 670.050 796.050 ;
        RECT 655.650 792.600 657.750 793.500 ;
        RECT 640.350 789.600 642.450 791.700 ;
        RECT 640.950 784.950 643.050 787.050 ;
        RECT 601.950 772.950 604.050 775.050 ;
        RECT 574.950 766.950 577.050 769.050 ;
        RECT 595.950 766.950 598.050 769.050 ;
        RECT 571.950 760.950 574.050 763.050 ;
        RECT 575.400 762.600 576.450 766.950 ;
        RECT 602.400 763.200 603.450 772.950 ;
        RECT 613.350 771.300 615.450 773.400 ;
        RECT 614.250 764.700 615.450 771.300 ;
        RECT 616.950 769.950 619.050 772.050 ;
        RECT 575.400 760.350 576.600 762.600 ;
        RECT 580.950 761.100 583.050 763.200 ;
        RECT 589.950 761.100 592.050 763.200 ;
        RECT 595.950 761.100 598.050 763.200 ;
        RECT 601.950 761.100 604.050 763.200 ;
        RECT 613.350 762.600 615.450 764.700 ;
        RECT 581.400 760.350 582.600 761.100 ;
        RECT 574.950 757.950 577.050 760.050 ;
        RECT 577.950 757.950 580.050 760.050 ;
        RECT 580.950 757.950 583.050 760.050 ;
        RECT 583.950 757.950 586.050 760.050 ;
        RECT 568.950 754.950 571.050 757.050 ;
        RECT 578.400 756.900 579.600 757.650 ;
        RECT 565.950 730.950 568.050 733.050 ;
        RECT 569.400 730.200 570.450 754.950 ;
        RECT 577.950 754.800 580.050 756.900 ;
        RECT 584.400 756.450 585.600 757.650 ;
        RECT 586.950 756.450 589.050 757.050 ;
        RECT 584.400 755.400 589.050 756.450 ;
        RECT 586.950 754.950 589.050 755.400 ;
        RECT 580.350 735.300 582.450 737.400 ;
        RECT 568.950 728.100 571.050 730.200 ;
        RECT 574.950 728.100 577.050 730.200 ;
        RECT 569.400 727.350 570.600 728.100 ;
        RECT 575.400 727.350 576.600 728.100 ;
        RECT 565.950 724.950 568.050 727.050 ;
        RECT 568.950 724.950 571.050 727.050 ;
        RECT 574.950 724.950 577.050 727.050 ;
        RECT 566.400 724.050 567.600 724.650 ;
        RECT 562.950 722.400 567.600 724.050 ;
        RECT 581.250 722.400 582.450 735.300 ;
        RECT 583.950 730.950 586.050 733.050 ;
        RECT 584.400 727.050 585.450 730.950 ;
        RECT 583.950 724.950 586.050 727.050 ;
        RECT 562.950 721.950 567.450 722.400 ;
        RECT 566.400 706.050 567.450 721.950 ;
        RECT 571.950 718.950 574.050 721.050 ;
        RECT 580.350 720.300 582.450 722.400 ;
        RECT 565.950 703.950 568.050 706.050 ;
        RECT 568.950 697.950 571.050 700.050 ;
        RECT 559.950 694.950 562.050 697.050 ;
        RECT 559.650 691.500 561.750 692.400 ;
        RECT 559.650 690.300 563.850 691.500 ;
        RECT 557.400 684.450 558.600 684.600 ;
        RECT 554.400 683.400 558.600 684.450 ;
        RECT 557.400 682.350 558.600 683.400 ;
        RECT 556.800 679.950 558.900 682.050 ;
        RECT 562.650 671.700 563.850 690.300 ;
        RECT 565.950 688.950 568.050 691.050 ;
        RECT 566.400 684.600 567.450 688.950 ;
        RECT 569.400 685.050 570.450 697.950 ;
        RECT 566.400 682.350 567.600 684.600 ;
        RECT 568.950 682.950 571.050 685.050 ;
        RECT 565.950 679.950 568.050 682.050 ;
        RECT 562.050 669.600 564.150 671.700 ;
        RECT 559.950 664.950 562.050 667.050 ;
        RECT 550.950 652.950 553.050 655.050 ;
        RECT 560.400 652.200 561.450 664.950 ;
        RECT 548.400 649.350 549.600 651.600 ;
        RECT 553.950 650.100 556.050 652.200 ;
        RECT 559.950 650.100 562.050 652.200 ;
        RECT 565.950 650.100 568.050 652.200 ;
        RECT 572.400 651.600 573.450 718.950 ;
        RECT 581.250 713.700 582.450 720.300 ;
        RECT 580.350 711.600 582.450 713.700 ;
        RECT 574.950 703.950 577.050 706.050 ;
        RECT 575.400 655.050 576.450 703.950 ;
        RECT 584.400 696.450 585.450 724.950 ;
        RECT 587.400 712.050 588.450 754.950 ;
        RECT 590.400 751.050 591.450 761.100 ;
        RECT 596.400 760.350 597.600 761.100 ;
        RECT 602.400 760.350 603.600 761.100 ;
        RECT 595.950 757.950 598.050 760.050 ;
        RECT 598.950 757.950 601.050 760.050 ;
        RECT 601.950 757.950 604.050 760.050 ;
        RECT 607.950 757.950 610.050 760.050 ;
        RECT 599.400 756.000 600.600 757.650 ;
        RECT 608.400 756.900 609.600 757.650 ;
        RECT 598.950 751.950 601.050 756.000 ;
        RECT 607.950 754.800 610.050 756.900 ;
        RECT 604.950 753.450 607.050 754.050 ;
        RECT 610.950 753.450 613.050 754.050 ;
        RECT 604.950 752.400 613.050 753.450 ;
        RECT 604.950 751.950 607.050 752.400 ;
        RECT 610.950 751.950 613.050 752.400 ;
        RECT 589.950 748.950 592.050 751.050 ;
        RECT 607.950 748.950 610.050 751.050 ;
        RECT 614.250 749.700 615.450 762.600 ;
        RECT 598.050 735.300 600.150 737.400 ;
        RECT 592.800 724.950 594.900 727.050 ;
        RECT 593.400 723.000 594.600 724.650 ;
        RECT 592.950 718.950 595.050 723.000 ;
        RECT 598.650 716.700 599.850 735.300 ;
        RECT 601.950 724.950 604.050 727.050 ;
        RECT 602.400 723.900 603.600 724.650 ;
        RECT 601.950 721.800 604.050 723.900 ;
        RECT 595.650 715.500 599.850 716.700 ;
        RECT 595.650 714.600 597.750 715.500 ;
        RECT 586.950 709.950 589.050 712.050 ;
        RECT 581.400 695.400 585.450 696.450 ;
        RECT 581.400 688.050 582.450 695.400 ;
        RECT 592.950 691.950 595.050 694.050 ;
        RECT 580.950 685.950 583.050 688.050 ;
        RECT 583.950 683.100 586.050 685.200 ;
        RECT 584.400 682.350 585.600 683.100 ;
        RECT 589.950 682.950 592.050 688.050 ;
        RECT 580.950 679.950 583.050 682.050 ;
        RECT 583.950 679.950 586.050 682.050 ;
        RECT 586.950 679.950 589.050 682.050 ;
        RECT 581.400 677.400 582.600 679.650 ;
        RECT 587.400 678.900 588.600 679.650 ;
        RECT 593.400 678.900 594.450 691.950 ;
        RECT 601.950 684.000 604.050 688.050 ;
        RECT 608.400 685.050 609.450 748.950 ;
        RECT 613.350 747.600 615.450 749.700 ;
        RECT 617.400 729.450 618.450 769.950 ;
        RECT 628.650 769.500 630.750 770.400 ;
        RECT 628.650 768.300 632.850 769.500 ;
        RECT 619.950 761.100 622.050 763.200 ;
        RECT 625.950 761.100 628.050 763.200 ;
        RECT 620.400 751.050 621.450 761.100 ;
        RECT 626.400 760.350 627.600 761.100 ;
        RECT 625.800 757.950 627.900 760.050 ;
        RECT 619.950 748.950 622.050 751.050 ;
        RECT 631.650 749.700 632.850 768.300 ;
        RECT 634.950 762.000 637.050 766.050 ;
        RECT 635.400 760.350 636.600 762.000 ;
        RECT 634.950 757.950 637.050 760.050 ;
        RECT 631.050 747.600 633.150 749.700 ;
        RECT 614.400 728.400 618.450 729.450 ;
        RECT 602.400 682.350 603.600 684.000 ;
        RECT 607.950 682.950 610.050 685.050 ;
        RECT 598.950 679.950 601.050 682.050 ;
        RECT 601.950 679.950 604.050 682.050 ;
        RECT 604.950 679.950 607.050 682.050 ;
        RECT 599.400 679.050 600.600 679.650 ;
        RECT 581.400 673.050 582.450 677.400 ;
        RECT 586.950 676.800 589.050 678.900 ;
        RECT 592.950 676.800 595.050 678.900 ;
        RECT 595.950 677.400 600.600 679.050 ;
        RECT 605.400 677.400 606.600 679.650 ;
        RECT 595.950 676.950 600.000 677.400 ;
        RECT 580.950 672.450 583.050 673.050 ;
        RECT 580.950 671.400 585.450 672.450 ;
        RECT 580.950 670.950 583.050 671.400 ;
        RECT 580.950 658.950 583.050 661.050 ;
        RECT 574.950 652.950 577.050 655.050 ;
        RECT 554.400 649.350 555.600 650.100 ;
        RECT 541.950 646.950 544.050 649.050 ;
        RECT 547.950 646.950 550.050 649.050 ;
        RECT 550.950 646.950 553.050 649.050 ;
        RECT 553.950 646.950 556.050 649.050 ;
        RECT 527.550 633.600 529.650 635.700 ;
        RECT 538.950 634.950 541.050 637.050 ;
        RECT 538.950 628.950 541.050 631.050 ;
        RECT 535.950 622.950 538.050 625.050 ;
        RECT 520.950 610.950 523.050 613.050 ;
        RECT 532.950 610.950 535.050 613.050 ;
        RECT 506.400 604.350 507.600 606.600 ;
        RECT 511.950 606.000 514.050 610.050 ;
        RECT 517.950 607.950 520.050 610.050 ;
        RECT 512.400 604.350 513.600 606.000 ;
        RECT 505.950 601.950 508.050 604.050 ;
        RECT 508.950 601.950 511.050 604.050 ;
        RECT 511.950 601.950 514.050 604.050 ;
        RECT 509.400 600.900 510.600 601.650 ;
        RECT 518.400 600.900 519.450 607.950 ;
        RECT 520.950 607.800 523.050 609.900 ;
        RECT 508.950 598.800 511.050 600.900 ;
        RECT 517.950 598.800 520.050 600.900 ;
        RECT 521.400 595.050 522.450 607.800 ;
        RECT 529.950 606.000 532.050 610.050 ;
        RECT 530.400 604.350 531.600 606.000 ;
        RECT 524.400 601.950 526.500 604.050 ;
        RECT 529.800 601.950 531.900 604.050 ;
        RECT 524.400 599.400 525.600 601.650 ;
        RECT 520.950 592.950 523.050 595.050 ;
        RECT 499.950 591.450 502.050 592.050 ;
        RECT 499.950 590.400 504.450 591.450 ;
        RECT 499.950 589.950 502.050 590.400 ;
        RECT 494.400 571.350 495.600 573.600 ;
        RECT 478.950 568.950 481.050 571.050 ;
        RECT 494.400 568.950 496.500 571.050 ;
        RECT 499.800 568.950 501.900 571.050 ;
        RECT 472.650 559.500 476.850 560.700 ;
        RECT 479.400 566.400 480.600 568.650 ;
        RECT 500.400 567.900 501.600 568.650 ;
        RECT 472.650 558.600 474.750 559.500 ;
        RECT 463.950 550.950 466.050 553.050 ;
        RECT 457.950 547.950 460.050 550.050 ;
        RECT 361.950 535.950 364.050 538.050 ;
        RECT 319.950 527.100 322.050 529.200 ;
        RECT 325.950 527.100 328.050 529.200 ;
        RECT 334.950 527.100 337.050 529.200 ;
        RECT 340.950 527.100 343.050 529.200 ;
        RECT 346.950 527.100 349.050 529.200 ;
        RECT 358.950 527.100 361.050 529.200 ;
        RECT 320.400 526.350 321.600 527.100 ;
        RECT 316.950 523.950 319.050 526.050 ;
        RECT 319.950 523.950 322.050 526.050 ;
        RECT 313.950 520.950 316.050 523.050 ;
        RECT 317.400 521.400 318.600 523.650 ;
        RECT 326.400 523.050 327.450 527.100 ;
        RECT 335.400 526.350 336.600 527.100 ;
        RECT 341.400 526.350 342.600 527.100 ;
        RECT 331.950 523.950 334.050 526.050 ;
        RECT 334.950 523.950 337.050 526.050 ;
        RECT 337.950 523.950 340.050 526.050 ;
        RECT 340.950 523.950 343.050 526.050 ;
        RECT 310.950 508.950 313.050 511.050 ;
        RECT 308.400 506.400 312.450 507.450 ;
        RECT 301.950 502.950 304.050 505.050 ;
        RECT 283.800 498.300 285.900 500.400 ;
        RECT 287.400 499.200 288.600 501.450 ;
        RECT 280.950 494.100 283.050 496.200 ;
        RECT 281.400 493.350 282.600 494.100 ;
        RECT 281.100 490.950 283.200 493.050 ;
        RECT 284.100 492.900 285.000 498.300 ;
        RECT 287.100 496.800 289.200 498.900 ;
        RECT 291.000 495.900 293.100 497.700 ;
        RECT 302.400 496.200 303.450 502.950 ;
        RECT 307.350 501.300 309.450 503.400 ;
        RECT 285.900 494.700 294.600 495.900 ;
        RECT 285.900 493.800 288.000 494.700 ;
        RECT 284.100 491.700 291.000 492.900 ;
        RECT 284.100 484.500 285.300 491.700 ;
        RECT 287.100 487.950 289.200 490.050 ;
        RECT 290.100 489.300 291.000 491.700 ;
        RECT 287.400 485.400 288.600 487.650 ;
        RECT 290.100 487.200 292.200 489.300 ;
        RECT 293.700 485.700 294.600 494.700 ;
        RECT 301.950 494.100 304.050 496.200 ;
        RECT 302.400 493.350 303.600 494.100 ;
        RECT 295.800 490.950 297.900 493.050 ;
        RECT 301.950 490.950 304.050 493.050 ;
        RECT 296.400 489.900 297.600 490.650 ;
        RECT 295.950 487.800 298.050 489.900 ;
        RECT 308.250 488.400 309.450 501.300 ;
        RECT 307.350 486.300 309.450 488.400 ;
        RECT 283.800 482.400 285.900 484.500 ;
        RECT 293.400 483.600 295.500 485.700 ;
        RECT 308.250 479.700 309.450 486.300 ;
        RECT 307.350 477.600 309.450 479.700 ;
        RECT 311.400 472.050 312.450 506.400 ;
        RECT 304.950 469.950 307.050 472.050 ;
        RECT 310.950 469.950 313.050 472.050 ;
        RECT 301.950 457.950 304.050 460.050 ;
        RECT 283.950 454.950 286.050 457.050 ;
        RECT 254.400 448.350 255.600 450.600 ;
        RECT 260.400 450.450 261.600 450.600 ;
        RECT 260.400 449.400 267.450 450.450 ;
        RECT 260.400 448.350 261.600 449.400 ;
        RECT 250.950 445.950 253.050 448.050 ;
        RECT 253.950 445.950 256.050 448.050 ;
        RECT 256.950 445.950 259.050 448.050 ;
        RECT 259.950 445.950 262.050 448.050 ;
        RECT 251.400 444.900 252.600 445.650 ;
        RECT 244.950 442.800 247.050 444.900 ;
        RECT 250.950 442.800 253.050 444.900 ;
        RECT 257.400 443.400 258.600 445.650 ;
        RECT 253.950 439.950 256.050 442.050 ;
        RECT 254.400 436.050 255.450 439.950 ;
        RECT 257.400 439.050 258.450 443.400 ;
        RECT 256.950 436.950 259.050 439.050 ;
        RECT 266.400 436.050 267.450 449.400 ;
        RECT 272.400 448.350 273.600 450.600 ;
        RECT 277.950 449.100 280.050 451.200 ;
        RECT 278.400 448.350 279.600 449.100 ;
        RECT 271.950 445.950 274.050 448.050 ;
        RECT 274.950 445.950 277.050 448.050 ;
        RECT 277.950 445.950 280.050 448.050 ;
        RECT 275.400 443.400 276.600 445.650 ;
        RECT 284.400 444.900 285.450 454.950 ;
        RECT 292.950 449.100 295.050 451.200 ;
        RECT 293.400 448.350 294.600 449.100 ;
        RECT 289.950 445.950 292.050 448.050 ;
        RECT 292.950 445.950 295.050 448.050 ;
        RECT 290.400 444.900 291.600 445.650 ;
        RECT 253.950 433.950 256.050 436.050 ;
        RECT 265.950 433.950 268.050 436.050 ;
        RECT 241.950 427.950 244.050 430.050 ;
        RECT 271.350 423.300 273.450 425.400 ;
        RECT 211.950 418.950 214.050 421.050 ;
        RECT 199.950 416.100 202.050 418.200 ;
        RECT 208.950 416.100 211.050 418.200 ;
        RECT 200.400 415.350 201.600 416.100 ;
        RECT 199.950 412.950 202.050 415.050 ;
        RECT 202.950 412.950 205.050 415.050 ;
        RECT 203.400 412.050 204.600 412.650 ;
        RECT 203.400 410.400 208.050 412.050 ;
        RECT 204.000 409.950 208.050 410.400 ;
        RECT 209.400 409.050 210.450 416.100 ;
        RECT 212.400 411.900 213.450 418.950 ;
        RECT 214.950 417.600 219.000 418.050 ;
        RECT 214.950 415.950 219.600 417.600 ;
        RECT 223.950 417.000 226.050 421.050 ;
        RECT 218.400 415.350 219.600 415.950 ;
        RECT 224.400 415.350 225.600 417.000 ;
        RECT 229.950 415.950 232.050 418.050 ;
        RECT 238.950 416.100 241.050 418.200 ;
        RECT 217.950 412.950 220.050 415.050 ;
        RECT 220.950 412.950 223.050 415.050 ;
        RECT 223.950 412.950 226.050 415.050 ;
        RECT 211.950 409.800 214.050 411.900 ;
        RECT 221.400 410.400 222.600 412.650 ;
        RECT 208.950 406.950 211.050 409.050 ;
        RECT 193.950 403.950 196.050 406.050 ;
        RECT 202.950 403.950 205.050 406.050 ;
        RECT 187.950 379.950 190.050 382.050 ;
        RECT 178.950 372.450 181.050 373.200 ;
        RECT 176.400 371.400 181.050 372.450 ;
        RECT 178.950 371.100 181.050 371.400 ;
        RECT 188.400 372.600 189.450 379.950 ;
        RECT 173.400 370.350 174.600 371.100 ;
        RECT 169.950 367.950 172.050 370.050 ;
        RECT 172.950 367.950 175.050 370.050 ;
        RECT 170.400 366.900 171.600 367.650 ;
        RECT 179.400 367.050 180.450 371.100 ;
        RECT 188.400 370.350 189.600 372.600 ;
        RECT 193.950 371.100 196.050 373.200 ;
        RECT 194.400 370.350 195.600 371.100 ;
        RECT 184.950 367.950 187.050 370.050 ;
        RECT 187.950 367.950 190.050 370.050 ;
        RECT 190.950 367.950 193.050 370.050 ;
        RECT 193.950 367.950 196.050 370.050 ;
        RECT 196.950 367.950 199.050 370.050 ;
        RECT 169.950 364.800 172.050 366.900 ;
        RECT 178.950 364.950 181.050 367.050 ;
        RECT 185.400 366.900 186.600 367.650 ;
        RECT 184.950 364.800 187.050 366.900 ;
        RECT 191.400 365.400 192.600 367.650 ;
        RECT 197.400 366.900 198.600 367.650 ;
        RECT 191.400 361.050 192.450 365.400 ;
        RECT 196.950 364.800 199.050 366.900 ;
        RECT 203.400 361.050 204.450 403.950 ;
        RECT 221.400 400.050 222.450 410.400 ;
        RECT 230.400 409.050 231.450 415.950 ;
        RECT 239.400 415.350 240.600 416.100 ;
        RECT 244.950 415.950 247.050 421.050 ;
        RECT 247.950 415.950 250.050 418.050 ;
        RECT 253.950 416.100 256.050 418.200 ;
        RECT 259.950 416.100 262.050 418.200 ;
        RECT 265.950 416.100 268.050 418.200 ;
        RECT 235.950 412.950 238.050 415.050 ;
        RECT 238.950 412.950 241.050 415.050 ;
        RECT 241.950 412.950 244.050 415.050 ;
        RECT 236.400 410.400 237.600 412.650 ;
        RECT 242.400 411.900 243.600 412.650 ;
        RECT 248.400 411.900 249.450 415.950 ;
        RECT 254.400 415.350 255.600 416.100 ;
        RECT 260.400 415.350 261.600 416.100 ;
        RECT 266.400 415.350 267.600 416.100 ;
        RECT 253.950 412.950 256.050 415.050 ;
        RECT 256.950 412.950 259.050 415.050 ;
        RECT 259.950 412.950 262.050 415.050 ;
        RECT 265.950 412.950 268.050 415.050 ;
        RECT 229.950 406.950 232.050 409.050 ;
        RECT 236.400 403.050 237.450 410.400 ;
        RECT 241.950 409.800 244.050 411.900 ;
        RECT 247.800 409.800 249.900 411.900 ;
        RECT 248.400 406.050 249.450 409.800 ;
        RECT 250.950 406.950 253.050 412.050 ;
        RECT 257.400 411.900 258.600 412.650 ;
        RECT 256.950 409.800 259.050 411.900 ;
        RECT 272.250 410.400 273.450 423.300 ;
        RECT 271.350 408.300 273.450 410.400 ;
        RECT 247.950 403.950 250.050 406.050 ;
        RECT 235.950 400.950 238.050 403.050 ;
        RECT 272.250 401.700 273.450 408.300 ;
        RECT 220.950 397.950 223.050 400.050 ;
        RECT 271.350 399.600 273.450 401.700 ;
        RECT 268.950 388.950 271.050 391.050 ;
        RECT 259.950 382.950 262.050 385.050 ;
        RECT 208.950 379.950 211.050 382.050 ;
        RECT 209.400 372.600 210.450 379.950 ;
        RECT 229.800 376.200 231.900 378.300 ;
        RECT 238.800 376.500 240.900 378.600 ;
        RECT 209.400 370.350 210.600 372.600 ;
        RECT 214.950 371.100 217.050 373.200 ;
        RECT 223.800 371.100 225.900 373.200 ;
        RECT 226.950 371.100 229.050 373.200 ;
        RECT 215.400 370.350 216.600 371.100 ;
        RECT 208.950 367.950 211.050 370.050 ;
        RECT 211.950 367.950 214.050 370.050 ;
        RECT 214.950 367.950 217.050 370.050 ;
        RECT 220.950 367.950 223.050 370.050 ;
        RECT 212.400 366.900 213.600 367.650 ;
        RECT 211.950 364.800 214.050 366.900 ;
        RECT 221.400 364.050 222.450 367.950 ;
        RECT 214.950 361.950 217.050 364.050 ;
        RECT 220.950 361.950 223.050 364.050 ;
        RECT 190.950 358.950 193.050 361.050 ;
        RECT 202.950 358.950 205.050 361.050 ;
        RECT 187.950 357.450 190.050 358.050 ;
        RECT 193.950 357.450 196.050 358.050 ;
        RECT 187.950 356.400 196.050 357.450 ;
        RECT 187.950 355.950 190.050 356.400 ;
        RECT 193.950 355.950 196.050 356.400 ;
        RECT 163.950 343.950 166.050 346.050 ;
        RECT 178.950 343.050 181.050 343.200 ;
        RECT 181.950 343.050 184.050 343.200 ;
        RECT 178.950 341.100 184.050 343.050 ;
        RECT 196.950 342.450 201.000 343.050 ;
        RECT 180.000 340.950 183.000 341.100 ;
        RECT 196.950 340.950 201.450 342.450 ;
        RECT 161.400 337.350 162.600 339.600 ;
        RECT 166.950 338.100 169.050 340.200 ;
        RECT 167.400 337.350 168.600 338.100 ;
        RECT 178.950 337.950 181.050 340.050 ;
        RECT 184.950 338.100 187.050 340.200 ;
        RECT 193.950 338.100 196.050 340.200 ;
        RECT 200.400 339.600 201.450 340.950 ;
        RECT 179.400 337.350 180.600 337.950 ;
        RECT 185.400 337.350 186.600 338.100 ;
        RECT 157.950 334.950 160.050 337.050 ;
        RECT 160.950 334.950 163.050 337.050 ;
        RECT 163.950 334.950 166.050 337.050 ;
        RECT 166.950 334.950 169.050 337.050 ;
        RECT 178.950 334.950 181.050 337.050 ;
        RECT 181.950 334.950 184.050 337.050 ;
        RECT 184.950 334.950 187.050 337.050 ;
        RECT 187.950 334.950 190.050 337.050 ;
        RECT 158.400 333.900 159.600 334.650 ;
        RECT 139.950 331.800 142.050 333.900 ;
        RECT 151.950 331.800 154.050 333.900 ;
        RECT 157.950 331.800 160.050 333.900 ;
        RECT 164.400 332.400 165.600 334.650 ;
        RECT 182.400 333.000 183.600 334.650 ;
        RECT 188.400 333.900 189.600 334.650 ;
        RECT 140.400 328.050 141.450 331.800 ;
        RECT 164.400 328.050 165.450 332.400 ;
        RECT 181.950 328.950 184.050 333.000 ;
        RECT 187.950 331.800 190.050 333.900 ;
        RECT 139.950 325.950 142.050 328.050 ;
        RECT 163.950 325.950 166.050 328.050 ;
        RECT 121.950 319.950 124.050 322.050 ;
        RECT 133.950 319.950 136.050 322.050 ;
        RECT 122.400 304.050 123.450 319.950 ;
        RECT 127.950 313.950 130.050 316.050 ;
        RECT 128.400 307.050 129.450 313.950 ;
        RECT 133.950 307.950 136.050 310.050 ;
        RECT 160.950 307.950 163.050 310.050 ;
        RECT 181.950 307.950 184.050 310.050 ;
        RECT 127.950 304.950 130.050 307.050 ;
        RECT 106.950 301.950 109.050 304.050 ;
        RECT 121.950 301.950 124.050 304.050 ;
        RECT 86.400 292.350 87.600 293.100 ;
        RECT 92.400 292.350 93.600 293.100 ;
        RECT 85.950 289.950 88.050 292.050 ;
        RECT 88.950 289.950 91.050 292.050 ;
        RECT 91.950 289.950 94.050 292.050 ;
        RECT 94.950 289.950 97.050 292.050 ;
        RECT 73.950 286.800 76.050 288.900 ;
        RECT 79.950 286.800 82.050 288.900 ;
        RECT 89.400 287.400 90.600 289.650 ;
        RECT 95.400 289.050 96.600 289.650 ;
        RECT 95.400 287.400 100.050 289.050 ;
        RECT 74.400 277.050 75.450 286.800 ;
        RECT 73.950 274.950 76.050 277.050 ;
        RECT 89.400 274.050 90.450 287.400 ;
        RECT 96.000 286.950 100.050 287.400 ;
        RECT 101.400 280.050 102.450 293.100 ;
        RECT 103.950 292.950 106.050 295.050 ;
        RECT 106.950 293.100 109.050 295.200 ;
        RECT 112.950 293.100 115.050 295.200 ;
        RECT 107.400 292.350 108.600 293.100 ;
        RECT 113.400 292.350 114.600 293.100 ;
        RECT 106.950 289.950 109.050 292.050 ;
        RECT 109.950 289.950 112.050 292.050 ;
        RECT 112.950 289.950 115.050 292.050 ;
        RECT 115.950 289.950 118.050 292.050 ;
        RECT 103.950 286.950 106.050 289.050 ;
        RECT 110.400 287.400 111.600 289.650 ;
        RECT 116.400 288.000 117.600 289.650 ;
        RECT 122.400 289.050 123.450 301.950 ;
        RECT 128.400 294.600 129.450 304.950 ;
        RECT 134.400 294.600 135.450 307.950 ;
        RECT 142.950 301.950 145.050 304.050 ;
        RECT 128.400 292.350 129.600 294.600 ;
        RECT 134.400 292.350 135.600 294.600 ;
        RECT 127.950 289.950 130.050 292.050 ;
        RECT 130.950 289.950 133.050 292.050 ;
        RECT 133.950 289.950 136.050 292.050 ;
        RECT 136.950 289.950 139.050 292.050 ;
        RECT 100.950 277.950 103.050 280.050 ;
        RECT 104.400 274.050 105.450 286.950 ;
        RECT 70.950 271.950 73.050 274.050 ;
        RECT 88.800 271.950 90.900 274.050 ;
        RECT 91.950 271.950 94.050 274.050 ;
        RECT 103.950 271.950 106.050 274.050 ;
        RECT 64.950 268.950 67.050 271.050 ;
        RECT 65.400 265.050 66.450 268.950 ;
        RECT 64.950 262.950 67.050 265.050 ;
        RECT 62.400 259.350 63.600 261.600 ;
        RECT 61.950 256.950 64.050 259.050 ;
        RECT 64.950 256.950 67.050 259.050 ;
        RECT 65.400 254.400 66.600 256.650 ;
        RECT 65.400 253.050 66.450 254.400 ;
        RECT 61.950 251.400 66.450 253.050 ;
        RECT 61.950 250.950 66.000 251.400 ;
        RECT 71.400 223.050 72.450 271.950 ;
        RECT 89.400 268.050 90.450 271.950 ;
        RECT 88.950 265.950 91.050 268.050 ;
        RECT 92.400 262.200 93.450 271.950 ;
        RECT 97.950 265.950 100.050 268.050 ;
        RECT 76.950 260.100 79.050 262.200 ;
        RECT 82.950 260.100 85.050 262.200 ;
        RECT 91.950 260.100 94.050 262.200 ;
        RECT 98.400 261.600 99.450 265.950 ;
        RECT 104.400 261.600 105.450 271.950 ;
        RECT 110.400 262.050 111.450 287.400 ;
        RECT 115.950 283.950 118.050 288.000 ;
        RECT 121.950 286.950 124.050 289.050 ;
        RECT 131.400 288.000 132.600 289.650 ;
        RECT 137.400 288.900 138.600 289.650 ;
        RECT 130.950 283.950 133.050 288.000 ;
        RECT 136.950 286.800 139.050 288.900 ;
        RECT 143.400 286.050 144.450 301.950 ;
        RECT 151.950 294.000 154.050 298.050 ;
        RECT 152.400 292.350 153.600 294.000 ;
        RECT 157.950 293.100 160.050 295.200 ;
        RECT 161.400 295.050 162.450 307.950 ;
        RECT 158.400 292.350 159.600 293.100 ;
        RECT 160.950 292.950 163.050 295.050 ;
        RECT 163.950 293.100 166.050 295.200 ;
        RECT 172.950 293.100 175.050 298.050 ;
        RECT 148.950 289.950 151.050 292.050 ;
        RECT 151.950 289.950 154.050 292.050 ;
        RECT 154.950 289.950 157.050 292.050 ;
        RECT 157.950 289.950 160.050 292.050 ;
        RECT 149.400 288.900 150.600 289.650 ;
        RECT 148.950 286.800 151.050 288.900 ;
        RECT 155.400 288.000 156.600 289.650 ;
        RECT 142.950 283.950 145.050 286.050 ;
        RECT 142.950 277.950 145.050 280.050 ;
        RECT 127.950 268.950 130.050 271.050 ;
        RECT 77.400 259.350 78.600 260.100 ;
        RECT 83.400 259.350 84.600 260.100 ;
        RECT 76.950 256.950 79.050 259.050 ;
        RECT 79.950 256.950 82.050 259.050 ;
        RECT 82.950 256.950 85.050 259.050 ;
        RECT 85.950 256.950 88.050 259.050 ;
        RECT 73.950 253.950 76.050 256.050 ;
        RECT 80.400 254.400 81.600 256.650 ;
        RECT 86.400 255.900 87.600 256.650 ;
        RECT 64.950 220.950 67.050 223.050 ;
        RECT 70.950 220.950 73.050 223.050 ;
        RECT 65.400 216.600 66.450 220.950 ;
        RECT 74.400 219.450 75.450 253.950 ;
        RECT 80.400 250.050 81.450 254.400 ;
        RECT 85.950 253.800 88.050 255.900 ;
        RECT 79.950 247.950 82.050 250.050 ;
        RECT 92.400 244.050 93.450 260.100 ;
        RECT 98.400 259.350 99.600 261.600 ;
        RECT 104.400 259.350 105.600 261.600 ;
        RECT 109.800 259.950 111.900 262.050 ;
        RECT 112.950 259.950 115.050 262.050 ;
        RECT 121.950 260.100 124.050 262.200 ;
        RECT 128.400 262.050 129.450 268.950 ;
        RECT 133.950 265.950 136.050 268.050 ;
        RECT 97.950 256.950 100.050 259.050 ;
        RECT 100.950 256.950 103.050 259.050 ;
        RECT 103.950 256.950 106.050 259.050 ;
        RECT 106.950 256.950 109.050 259.050 ;
        RECT 101.400 255.900 102.600 256.650 ;
        RECT 100.950 253.800 103.050 255.900 ;
        RECT 107.400 255.000 108.600 256.650 ;
        RECT 79.950 241.950 82.050 244.050 ;
        RECT 91.950 241.950 94.050 244.050 ;
        RECT 71.400 218.400 75.450 219.450 ;
        RECT 71.400 216.600 72.450 218.400 ;
        RECT 56.400 215.400 60.450 216.450 ;
        RECT 50.400 214.350 51.600 215.100 ;
        RECT 49.950 211.950 52.050 214.050 ;
        RECT 52.950 211.950 55.050 214.050 ;
        RECT 41.400 209.400 45.450 210.450 ;
        RECT 53.400 209.400 54.600 211.650 ;
        RECT 59.400 210.900 60.450 215.400 ;
        RECT 65.400 214.350 66.600 216.600 ;
        RECT 71.400 214.350 72.600 216.600 ;
        RECT 64.950 211.950 67.050 214.050 ;
        RECT 67.950 211.950 70.050 214.050 ;
        RECT 70.950 211.950 73.050 214.050 ;
        RECT 73.950 211.950 76.050 214.050 ;
        RECT 22.950 199.950 25.050 202.050 ;
        RECT 19.950 184.950 25.050 187.050 ;
        RECT 26.400 184.050 27.450 208.950 ;
        RECT 29.400 196.050 30.450 209.400 ;
        RECT 35.400 202.050 36.450 209.400 ;
        RECT 34.950 199.950 37.050 202.050 ;
        RECT 28.950 193.950 31.050 196.050 ;
        RECT 14.400 181.350 15.600 183.600 ;
        RECT 25.950 181.950 28.050 184.050 ;
        RECT 34.950 183.000 37.050 187.050 ;
        RECT 41.400 184.200 42.450 209.400 ;
        RECT 53.400 207.450 54.450 209.400 ;
        RECT 58.950 208.800 61.050 210.900 ;
        RECT 68.400 209.400 69.600 211.650 ;
        RECT 74.400 210.900 75.600 211.650 ;
        RECT 80.400 211.050 81.450 241.950 ;
        RECT 88.950 226.950 91.050 229.050 ;
        RECT 89.400 216.600 90.450 226.950 ;
        RECT 89.400 214.350 90.600 216.600 ;
        RECT 94.950 215.100 97.050 217.200 ;
        RECT 95.400 214.350 96.600 215.100 ;
        RECT 85.950 211.950 88.050 214.050 ;
        RECT 88.950 211.950 91.050 214.050 ;
        RECT 91.950 211.950 94.050 214.050 ;
        RECT 94.950 211.950 97.050 214.050 ;
        RECT 50.400 206.400 54.450 207.450 ;
        RECT 35.400 181.350 36.600 183.000 ;
        RECT 40.950 182.100 43.050 184.200 ;
        RECT 41.400 181.350 42.600 182.100 ;
        RECT 10.950 178.950 13.050 181.050 ;
        RECT 13.950 178.950 16.050 181.050 ;
        RECT 16.950 178.950 19.050 181.050 ;
        RECT 31.950 178.950 34.050 181.050 ;
        RECT 34.950 178.950 37.050 181.050 ;
        RECT 37.950 178.950 40.050 181.050 ;
        RECT 40.950 178.950 43.050 181.050 ;
        RECT 43.950 178.950 46.050 181.050 ;
        RECT 11.400 177.900 12.600 178.650 ;
        RECT 17.400 177.900 18.600 178.650 ;
        RECT 32.400 177.900 33.600 178.650 ;
        RECT 4.950 175.800 7.050 177.900 ;
        RECT 10.950 175.800 13.050 177.900 ;
        RECT 16.950 175.800 19.050 177.900 ;
        RECT 25.950 175.800 28.050 177.900 ;
        RECT 31.950 175.800 34.050 177.900 ;
        RECT 38.400 176.400 39.600 178.650 ;
        RECT 44.400 177.900 45.600 178.650 ;
        RECT 1.950 130.950 4.050 133.050 ;
        RECT 5.400 55.050 6.450 175.800 ;
        RECT 13.950 137.100 16.050 142.050 ;
        RECT 20.400 138.450 21.600 138.600 ;
        RECT 22.950 138.450 25.050 142.050 ;
        RECT 20.400 138.000 25.050 138.450 ;
        RECT 20.400 137.400 24.450 138.000 ;
        RECT 14.400 136.350 15.600 137.100 ;
        RECT 20.400 136.350 21.600 137.400 ;
        RECT 26.400 136.050 27.450 175.800 ;
        RECT 38.400 169.050 39.450 176.400 ;
        RECT 43.950 175.800 46.050 177.900 ;
        RECT 50.400 175.050 51.450 206.400 ;
        RECT 68.400 184.200 69.450 209.400 ;
        RECT 73.950 208.800 76.050 210.900 ;
        RECT 79.950 208.950 82.050 211.050 ;
        RECT 86.400 210.900 87.600 211.650 ;
        RECT 85.950 208.800 88.050 210.900 ;
        RECT 92.400 209.400 93.600 211.650 ;
        RECT 92.400 193.050 93.450 209.400 ;
        RECT 97.950 208.950 100.050 211.050 ;
        RECT 98.400 199.050 99.450 208.950 ;
        RECT 97.950 196.950 100.050 199.050 ;
        RECT 101.400 196.050 102.450 253.800 ;
        RECT 106.950 250.950 109.050 255.000 ;
        RECT 113.400 238.050 114.450 259.950 ;
        RECT 122.400 259.350 123.600 260.100 ;
        RECT 127.950 259.950 130.050 262.050 ;
        RECT 118.950 256.950 121.050 259.050 ;
        RECT 121.950 256.950 124.050 259.050 ;
        RECT 124.950 256.950 127.050 259.050 ;
        RECT 119.400 254.400 120.600 256.650 ;
        RECT 125.400 255.900 126.600 256.650 ;
        RECT 134.400 255.900 135.450 265.950 ;
        RECT 143.400 261.600 144.450 277.950 ;
        RECT 149.400 268.050 150.450 286.800 ;
        RECT 154.950 283.950 157.050 288.000 ;
        RECT 164.400 277.050 165.450 293.100 ;
        RECT 173.400 292.350 174.600 293.100 ;
        RECT 169.950 289.950 172.050 292.050 ;
        RECT 172.950 289.950 175.050 292.050 ;
        RECT 175.950 289.950 178.050 292.050 ;
        RECT 166.950 286.950 169.050 289.050 ;
        RECT 170.400 287.400 171.600 289.650 ;
        RECT 176.400 288.450 177.600 289.650 ;
        RECT 182.400 288.450 183.450 307.950 ;
        RECT 188.400 301.050 189.450 331.800 ;
        RECT 194.400 328.050 195.450 338.100 ;
        RECT 200.400 337.350 201.600 339.600 ;
        RECT 205.950 338.100 208.050 340.200 ;
        RECT 206.400 337.350 207.600 338.100 ;
        RECT 199.950 334.950 202.050 337.050 ;
        RECT 202.950 334.950 205.050 337.050 ;
        RECT 205.950 334.950 208.050 337.050 ;
        RECT 208.950 334.950 211.050 337.050 ;
        RECT 203.400 333.900 204.600 334.650 ;
        RECT 209.400 333.900 210.600 334.650 ;
        RECT 202.950 331.800 205.050 333.900 ;
        RECT 208.950 328.950 211.050 333.900 ;
        RECT 193.950 325.950 196.050 328.050 ;
        RECT 199.950 325.950 202.050 328.050 ;
        RECT 187.950 298.950 190.050 301.050 ;
        RECT 190.950 293.100 193.050 295.200 ;
        RECT 196.950 293.100 199.050 295.200 ;
        RECT 200.400 295.050 201.450 325.950 ;
        RECT 215.400 298.050 216.450 361.950 ;
        RECT 224.400 355.050 225.450 371.100 ;
        RECT 227.400 370.350 228.600 371.100 ;
        RECT 227.100 367.950 229.200 370.050 ;
        RECT 230.100 363.600 231.000 376.200 ;
        RECT 236.400 373.350 237.600 375.600 ;
        RECT 236.100 370.950 238.200 373.050 ;
        RECT 231.900 369.900 234.000 370.200 ;
        RECT 240.000 369.900 240.900 376.500 ;
        RECT 260.400 376.050 261.450 382.950 ;
        RECT 259.950 373.950 262.050 376.050 ;
        RECT 254.400 372.450 255.600 372.600 ;
        RECT 251.400 371.400 255.600 372.450 ;
        RECT 231.900 369.000 240.900 369.900 ;
        RECT 231.900 368.100 234.000 369.000 ;
        RECT 237.000 367.200 239.100 368.100 ;
        RECT 231.900 366.000 239.100 367.200 ;
        RECT 231.900 365.100 234.000 366.000 ;
        RECT 229.500 361.500 231.600 363.600 ;
        RECT 232.950 361.950 235.050 364.050 ;
        RECT 236.100 362.100 238.200 364.200 ;
        RECT 240.000 363.900 240.900 369.000 ;
        RECT 241.800 367.950 243.900 370.050 ;
        RECT 242.400 366.450 243.600 367.650 ;
        RECT 242.400 365.400 246.450 366.450 ;
        RECT 223.950 352.950 226.050 355.050 ;
        RECT 220.950 343.950 223.050 346.050 ;
        RECT 221.400 339.600 222.450 343.950 ;
        RECT 221.400 337.350 222.600 339.600 ;
        RECT 226.950 338.100 229.050 340.200 ;
        RECT 233.400 340.050 234.450 361.950 ;
        RECT 239.400 361.800 241.500 363.900 ;
        RECT 236.400 361.050 237.600 361.800 ;
        RECT 235.950 358.950 238.050 361.050 ;
        RECT 245.400 346.050 246.450 365.400 ;
        RECT 251.400 352.050 252.450 371.400 ;
        RECT 254.400 370.350 255.600 371.400 ;
        RECT 262.950 371.100 265.050 373.200 ;
        RECT 269.400 372.600 270.450 388.950 ;
        RECT 275.400 385.050 276.450 443.400 ;
        RECT 283.950 442.800 286.050 444.900 ;
        RECT 289.950 442.800 292.050 444.900 ;
        RECT 295.950 442.950 298.050 445.050 ;
        RECT 284.400 421.050 285.450 442.800 ;
        RECT 296.400 436.050 297.450 442.950 ;
        RECT 302.400 436.050 303.450 457.950 ;
        RECT 305.400 450.600 306.450 469.950 ;
        RECT 305.400 448.350 306.600 450.600 ;
        RECT 305.100 445.950 307.200 448.050 ;
        RECT 310.500 445.950 312.600 448.050 ;
        RECT 311.400 443.400 312.600 445.650 ;
        RECT 295.950 433.950 298.050 436.050 ;
        RECT 301.950 433.950 304.050 436.050 ;
        RECT 307.950 433.950 310.050 436.050 ;
        RECT 289.050 423.300 291.150 425.400 ;
        RECT 304.950 424.950 307.050 427.050 ;
        RECT 283.950 418.950 286.050 421.050 ;
        RECT 277.950 416.100 280.050 418.200 ;
        RECT 278.400 403.050 279.450 416.100 ;
        RECT 283.800 412.950 285.900 415.050 ;
        RECT 284.400 411.900 285.600 412.650 ;
        RECT 283.950 409.800 286.050 411.900 ;
        RECT 289.650 404.700 290.850 423.300 ;
        RECT 301.950 418.950 304.050 421.050 ;
        RECT 292.950 412.950 295.050 415.050 ;
        RECT 286.650 403.500 290.850 404.700 ;
        RECT 293.400 410.400 294.600 412.650 ;
        RECT 277.950 400.950 280.050 403.050 ;
        RECT 286.650 402.600 288.750 403.500 ;
        RECT 293.400 400.050 294.450 410.400 ;
        RECT 292.950 397.950 295.050 400.050 ;
        RECT 293.400 391.050 294.450 397.950 ;
        RECT 292.950 388.950 295.050 391.050 ;
        RECT 283.950 385.950 286.050 388.050 ;
        RECT 274.950 382.950 277.050 385.050 ;
        RECT 275.250 379.500 277.350 380.400 ;
        RECT 273.150 378.300 277.350 379.500 ;
        RECT 263.400 370.350 264.600 371.100 ;
        RECT 269.400 370.350 270.600 372.600 ;
        RECT 254.100 367.950 256.200 370.050 ;
        RECT 259.500 367.950 261.600 370.050 ;
        RECT 262.800 367.950 264.900 370.050 ;
        RECT 268.950 367.950 271.050 370.050 ;
        RECT 260.400 366.900 261.600 367.650 ;
        RECT 259.950 364.800 262.050 366.900 ;
        RECT 273.150 359.700 274.350 378.300 ;
        RECT 277.950 371.100 280.050 373.200 ;
        RECT 278.400 370.350 279.600 371.100 ;
        RECT 278.100 367.950 280.200 370.050 ;
        RECT 272.850 357.600 274.950 359.700 ;
        RECT 284.400 355.050 285.450 385.950 ;
        RECT 290.550 381.300 292.650 383.400 ;
        RECT 290.550 374.700 291.750 381.300 ;
        RECT 290.550 372.600 292.650 374.700 ;
        RECT 286.950 361.950 289.050 364.050 ;
        RECT 274.950 352.950 277.050 355.050 ;
        RECT 283.950 352.950 286.050 355.050 ;
        RECT 250.950 349.950 253.050 352.050 ;
        RECT 235.950 343.950 238.050 346.050 ;
        RECT 244.950 343.950 247.050 346.050 ;
        RECT 262.950 343.950 265.050 346.050 ;
        RECT 271.950 343.950 274.050 346.050 ;
        RECT 227.400 337.350 228.600 338.100 ;
        RECT 232.950 337.950 235.050 340.050 ;
        RECT 220.950 334.950 223.050 337.050 ;
        RECT 223.950 334.950 226.050 337.050 ;
        RECT 226.950 334.950 229.050 337.050 ;
        RECT 224.400 333.900 225.600 334.650 ;
        RECT 223.950 331.800 226.050 333.900 ;
        RECT 229.950 325.950 232.050 328.050 ;
        RECT 217.950 301.950 220.050 304.050 ;
        RECT 214.950 295.950 217.050 298.050 ;
        RECT 218.400 295.200 219.450 301.950 ;
        RECT 191.400 292.350 192.600 293.100 ;
        RECT 197.400 292.350 198.600 293.100 ;
        RECT 199.950 292.950 202.050 295.050 ;
        RECT 211.950 293.100 214.050 295.200 ;
        RECT 217.950 293.100 220.050 295.200 ;
        RECT 223.950 293.100 226.050 295.200 ;
        RECT 230.400 294.600 231.450 325.950 ;
        RECT 236.400 310.050 237.450 343.950 ;
        RECT 244.950 338.100 247.050 340.200 ;
        RECT 263.400 339.600 264.450 343.950 ;
        RECT 245.400 337.350 246.600 338.100 ;
        RECT 263.400 337.350 264.600 339.600 ;
        RECT 241.950 334.950 244.050 337.050 ;
        RECT 244.950 334.950 247.050 337.050 ;
        RECT 247.950 334.950 250.050 337.050 ;
        RECT 259.950 334.950 262.050 337.050 ;
        RECT 262.950 334.950 265.050 337.050 ;
        RECT 265.950 334.950 268.050 337.050 ;
        RECT 242.400 332.400 243.600 334.650 ;
        RECT 248.400 333.450 249.600 334.650 ;
        RECT 248.400 332.400 252.450 333.450 ;
        RECT 242.400 328.050 243.450 332.400 ;
        RECT 241.950 325.950 244.050 328.050 ;
        RECT 247.950 316.950 250.050 319.050 ;
        RECT 235.950 307.950 238.050 310.050 ;
        RECT 244.950 301.950 247.050 304.050 ;
        RECT 245.400 295.050 246.450 301.950 ;
        RECT 248.400 295.200 249.450 316.950 ;
        RECT 251.400 298.050 252.450 332.400 ;
        RECT 260.400 332.400 261.600 334.650 ;
        RECT 266.400 333.900 267.600 334.650 ;
        RECT 272.400 333.900 273.450 343.950 ;
        RECT 260.400 325.050 261.450 332.400 ;
        RECT 265.950 331.800 268.050 333.900 ;
        RECT 271.950 331.800 274.050 333.900 ;
        RECT 259.950 322.950 262.050 325.050 ;
        RECT 253.950 301.950 256.050 304.050 ;
        RECT 250.950 295.950 253.050 298.050 ;
        RECT 212.400 292.350 213.600 293.100 ;
        RECT 218.400 292.350 219.600 293.100 ;
        RECT 187.950 289.950 190.050 292.050 ;
        RECT 190.950 289.950 193.050 292.050 ;
        RECT 193.950 289.950 196.050 292.050 ;
        RECT 196.950 289.950 199.050 292.050 ;
        RECT 202.950 289.950 205.050 292.050 ;
        RECT 208.950 289.950 211.050 292.050 ;
        RECT 211.950 289.950 214.050 292.050 ;
        RECT 214.950 289.950 217.050 292.050 ;
        RECT 217.950 289.950 220.050 292.050 ;
        RECT 176.400 287.400 183.450 288.450 ;
        RECT 188.400 287.400 189.600 289.650 ;
        RECT 194.400 288.900 195.600 289.650 ;
        RECT 163.950 274.950 166.050 277.050 ;
        RECT 148.950 265.950 151.050 268.050 ;
        RECT 143.400 259.350 144.600 261.600 ;
        RECT 148.950 260.100 151.050 262.200 ;
        RECT 154.950 260.100 157.050 262.200 ;
        RECT 160.950 260.100 163.050 262.200 ;
        RECT 167.400 261.600 168.450 286.950 ;
        RECT 170.400 283.050 171.450 287.400 ;
        RECT 169.950 280.950 172.050 283.050 ;
        RECT 175.950 280.950 178.050 283.050 ;
        RECT 181.950 280.950 184.050 283.050 ;
        RECT 149.400 259.350 150.600 260.100 ;
        RECT 139.950 256.950 142.050 259.050 ;
        RECT 142.950 256.950 145.050 259.050 ;
        RECT 145.950 256.950 148.050 259.050 ;
        RECT 148.950 256.950 151.050 259.050 ;
        RECT 140.400 255.900 141.600 256.650 ;
        RECT 112.950 235.950 115.050 238.050 ;
        RECT 119.400 235.050 120.450 254.400 ;
        RECT 124.950 253.800 127.050 255.900 ;
        RECT 133.950 253.800 136.050 255.900 ;
        RECT 139.950 253.800 142.050 255.900 ;
        RECT 146.400 254.400 147.600 256.650 ;
        RECT 124.950 244.950 127.050 247.050 ;
        RECT 118.950 232.950 121.050 235.050 ;
        RECT 112.950 220.950 115.050 223.050 ;
        RECT 121.950 220.950 124.050 223.050 ;
        RECT 106.950 215.100 109.050 217.200 ;
        RECT 113.400 216.600 114.450 220.950 ;
        RECT 107.400 214.350 108.600 215.100 ;
        RECT 113.400 214.350 114.600 216.600 ;
        RECT 106.950 211.950 109.050 214.050 ;
        RECT 109.950 211.950 112.050 214.050 ;
        RECT 112.950 211.950 115.050 214.050 ;
        RECT 115.950 211.950 118.050 214.050 ;
        RECT 103.950 208.950 106.050 211.050 ;
        RECT 110.400 209.400 111.600 211.650 ;
        RECT 116.400 209.400 117.600 211.650 ;
        RECT 104.400 205.050 105.450 208.950 ;
        RECT 103.950 202.950 106.050 205.050 ;
        RECT 100.950 193.950 103.050 196.050 ;
        RECT 91.950 190.950 94.050 193.050 ;
        RECT 79.950 187.950 82.050 190.050 ;
        RECT 80.400 184.200 81.450 187.950 ;
        RECT 88.950 184.950 91.050 187.050 ;
        RECT 55.950 182.100 58.050 184.200 ;
        RECT 61.950 182.100 64.050 184.200 ;
        RECT 67.950 182.100 70.050 184.200 ;
        RECT 73.950 182.100 76.050 184.200 ;
        RECT 79.950 182.100 82.050 184.200 ;
        RECT 56.400 181.350 57.600 182.100 ;
        RECT 62.400 181.350 63.600 182.100 ;
        RECT 55.950 178.950 58.050 181.050 ;
        RECT 58.950 178.950 61.050 181.050 ;
        RECT 61.950 178.950 64.050 181.050 ;
        RECT 64.950 178.950 67.050 181.050 ;
        RECT 59.400 176.400 60.600 178.650 ;
        RECT 65.400 177.000 66.600 178.650 ;
        RECT 49.950 172.950 52.050 175.050 ;
        RECT 37.950 166.950 40.050 169.050 ;
        RECT 31.950 138.000 34.050 142.050 ;
        RECT 32.400 136.350 33.600 138.000 ;
        RECT 37.950 137.100 40.050 142.050 ;
        RECT 46.950 137.100 49.050 139.200 ;
        RECT 50.400 139.050 51.450 172.950 ;
        RECT 59.400 172.050 60.450 176.400 ;
        RECT 64.950 172.950 67.050 177.000 ;
        RECT 58.950 169.950 61.050 172.050 ;
        RECT 64.950 169.800 67.050 171.900 ;
        RECT 61.950 151.950 64.050 154.050 ;
        RECT 62.400 139.200 63.450 151.950 ;
        RECT 38.400 136.350 39.600 137.100 ;
        RECT 10.950 133.950 13.050 136.050 ;
        RECT 13.950 133.950 16.050 136.050 ;
        RECT 16.950 133.950 19.050 136.050 ;
        RECT 19.950 133.950 22.050 136.050 ;
        RECT 25.950 133.950 28.050 136.050 ;
        RECT 31.950 133.950 34.050 136.050 ;
        RECT 34.950 133.950 37.050 136.050 ;
        RECT 37.950 133.950 40.050 136.050 ;
        RECT 40.950 133.950 43.050 136.050 ;
        RECT 11.400 132.900 12.600 133.650 ;
        RECT 10.950 130.800 13.050 132.900 ;
        RECT 17.400 132.000 18.600 133.650 ;
        RECT 16.950 127.950 19.050 132.000 ;
        RECT 28.950 130.950 31.050 133.050 ;
        RECT 35.400 131.400 36.600 133.650 ;
        RECT 41.400 133.050 42.600 133.650 ;
        RECT 41.400 131.400 46.050 133.050 ;
        RECT 19.950 127.950 22.050 130.050 ;
        RECT 25.950 127.950 28.050 130.050 ;
        RECT 16.950 115.950 19.050 118.050 ;
        RECT 17.400 112.050 18.450 115.950 ;
        RECT 10.950 109.950 13.050 112.050 ;
        RECT 16.950 109.950 19.050 112.050 ;
        RECT 11.400 105.600 12.450 109.950 ;
        RECT 20.400 109.050 21.450 127.950 ;
        RECT 22.950 121.950 25.050 124.050 ;
        RECT 19.950 106.950 22.050 109.050 ;
        RECT 11.400 103.350 12.600 105.600 ;
        RECT 10.950 100.950 13.050 103.050 ;
        RECT 13.950 100.950 16.050 103.050 ;
        RECT 14.400 99.900 15.600 100.650 ;
        RECT 20.400 100.050 21.450 106.950 ;
        RECT 23.400 106.050 24.450 121.950 ;
        RECT 26.400 121.050 27.450 127.950 ;
        RECT 25.950 118.950 28.050 121.050 ;
        RECT 29.400 118.050 30.450 130.950 ;
        RECT 31.950 127.950 34.050 130.050 ;
        RECT 28.950 115.950 31.050 118.050 ;
        RECT 32.400 112.050 33.450 127.950 ;
        RECT 35.400 121.050 36.450 131.400 ;
        RECT 42.000 130.950 46.050 131.400 ;
        RECT 34.950 118.950 37.050 121.050 ;
        RECT 40.950 118.950 43.050 121.050 ;
        RECT 47.400 120.450 48.450 137.100 ;
        RECT 49.950 136.950 52.050 139.050 ;
        RECT 55.950 137.100 58.050 139.200 ;
        RECT 61.800 137.100 63.900 139.200 ;
        RECT 65.400 139.050 66.450 169.800 ;
        RECT 74.400 169.050 75.450 182.100 ;
        RECT 80.400 181.350 81.600 182.100 ;
        RECT 79.950 178.950 82.050 181.050 ;
        RECT 82.950 178.950 85.050 181.050 ;
        RECT 83.400 177.900 84.600 178.650 ;
        RECT 82.950 175.800 85.050 177.900 ;
        RECT 67.950 166.950 70.050 169.050 ;
        RECT 73.950 166.950 76.050 169.050 ;
        RECT 56.400 136.350 57.600 137.100 ;
        RECT 62.400 136.350 63.600 137.100 ;
        RECT 64.950 136.950 67.050 139.050 ;
        RECT 52.950 133.950 55.050 136.050 ;
        RECT 55.950 133.950 58.050 136.050 ;
        RECT 58.950 133.950 61.050 136.050 ;
        RECT 61.950 133.950 64.050 136.050 ;
        RECT 49.950 130.950 52.050 133.050 ;
        RECT 53.400 131.400 54.600 133.650 ;
        RECT 59.400 132.900 60.600 133.650 ;
        RECT 50.400 124.050 51.450 130.950 ;
        RECT 49.950 121.950 52.050 124.050 ;
        RECT 47.400 119.400 51.450 120.450 ;
        RECT 31.950 109.950 34.050 112.050 ;
        RECT 22.950 103.950 25.050 106.050 ;
        RECT 28.950 105.000 31.050 109.050 ;
        RECT 29.400 103.350 30.600 105.000 ;
        RECT 34.950 104.100 37.050 106.200 ;
        RECT 35.400 103.350 36.600 104.100 ;
        RECT 25.950 100.950 28.050 103.050 ;
        RECT 28.950 100.950 31.050 103.050 ;
        RECT 31.950 100.950 34.050 103.050 ;
        RECT 34.950 100.950 37.050 103.050 ;
        RECT 13.950 97.800 16.050 99.900 ;
        RECT 19.950 97.950 22.050 100.050 ;
        RECT 22.950 97.950 25.050 100.050 ;
        RECT 26.400 99.900 27.600 100.650 ;
        RECT 32.400 99.900 33.600 100.650 ;
        RECT 23.400 78.450 24.450 97.950 ;
        RECT 25.950 97.800 28.050 99.900 ;
        RECT 31.950 97.800 34.050 99.900 ;
        RECT 37.950 97.950 40.050 100.050 ;
        RECT 41.400 99.450 42.450 118.950 ;
        RECT 47.400 109.050 48.450 119.400 ;
        RECT 50.400 111.450 51.450 119.400 ;
        RECT 53.400 115.050 54.450 131.400 ;
        RECT 58.950 130.800 61.050 132.900 ;
        RECT 68.400 130.050 69.450 166.950 ;
        RECT 89.400 145.050 90.450 184.950 ;
        RECT 92.400 184.050 93.450 190.950 ;
        RECT 91.950 181.950 94.050 184.050 ;
        RECT 97.950 183.000 100.050 187.050 ;
        RECT 104.400 183.600 105.450 202.950 ;
        RECT 110.400 196.050 111.450 209.400 ;
        RECT 109.950 193.950 112.050 196.050 ;
        RECT 116.400 190.050 117.450 209.400 ;
        RECT 122.400 198.450 123.450 220.950 ;
        RECT 125.400 217.050 126.450 244.950 ;
        RECT 146.400 244.050 147.450 254.400 ;
        RECT 155.400 247.050 156.450 260.100 ;
        RECT 161.400 259.350 162.600 260.100 ;
        RECT 167.400 259.350 168.600 261.600 ;
        RECT 160.950 256.950 163.050 259.050 ;
        RECT 163.950 256.950 166.050 259.050 ;
        RECT 166.950 256.950 169.050 259.050 ;
        RECT 169.950 256.950 172.050 259.050 ;
        RECT 164.400 254.400 165.600 256.650 ;
        RECT 170.400 255.900 171.600 256.650 ;
        RECT 154.950 244.950 157.050 247.050 ;
        RECT 164.400 244.050 165.450 254.400 ;
        RECT 169.950 250.950 172.050 255.900 ;
        RECT 176.400 255.450 177.450 280.950 ;
        RECT 182.400 277.050 183.450 280.950 ;
        RECT 181.950 274.950 184.050 277.050 ;
        RECT 188.400 271.050 189.450 287.400 ;
        RECT 193.950 286.800 196.050 288.900 ;
        RECT 196.950 283.950 199.050 286.050 ;
        RECT 190.950 274.950 193.050 277.050 ;
        RECT 187.950 268.950 190.050 271.050 ;
        RECT 184.950 260.100 187.050 262.200 ;
        RECT 191.400 261.600 192.450 274.950 ;
        RECT 193.950 268.950 196.050 271.050 ;
        RECT 194.400 262.050 195.450 268.950 ;
        RECT 197.400 265.050 198.450 283.950 ;
        RECT 203.400 277.050 204.450 289.950 ;
        RECT 209.400 289.050 210.600 289.650 ;
        RECT 205.950 287.400 210.600 289.050 ;
        RECT 215.400 287.400 216.600 289.650 ;
        RECT 205.950 286.950 210.000 287.400 ;
        RECT 215.400 283.050 216.450 287.400 ;
        RECT 220.950 286.950 223.050 289.050 ;
        RECT 214.950 280.950 217.050 283.050 ;
        RECT 211.950 277.950 214.050 280.050 ;
        RECT 202.950 274.950 205.050 277.050 ;
        RECT 196.950 262.950 199.050 265.050 ;
        RECT 185.400 259.350 186.600 260.100 ;
        RECT 191.400 259.350 192.600 261.600 ;
        RECT 193.950 259.950 196.050 262.050 ;
        RECT 181.950 256.950 184.050 259.050 ;
        RECT 184.950 256.950 187.050 259.050 ;
        RECT 187.950 256.950 190.050 259.050 ;
        RECT 190.950 256.950 193.050 259.050 ;
        RECT 176.400 254.400 180.450 255.450 ;
        RECT 145.950 241.950 148.050 244.050 ;
        RECT 163.950 241.950 166.050 244.050 ;
        RECT 142.950 235.950 145.050 238.050 ;
        RECT 166.950 235.950 169.050 238.050 ;
        RECT 136.950 223.950 139.050 226.050 ;
        RECT 124.950 214.950 127.050 217.050 ;
        RECT 130.950 215.100 133.050 217.200 ;
        RECT 137.400 216.600 138.450 223.950 ;
        RECT 131.400 214.350 132.600 215.100 ;
        RECT 137.400 214.350 138.600 216.600 ;
        RECT 127.950 211.950 130.050 214.050 ;
        RECT 130.950 211.950 133.050 214.050 ;
        RECT 133.950 211.950 136.050 214.050 ;
        RECT 136.950 211.950 139.050 214.050 ;
        RECT 128.400 211.050 129.600 211.650 ;
        RECT 124.950 209.400 129.600 211.050 ;
        RECT 134.400 209.400 135.600 211.650 ;
        RECT 124.950 208.950 129.000 209.400 ;
        RECT 127.950 205.950 130.050 208.050 ;
        RECT 128.400 199.050 129.450 205.950 ;
        RECT 122.400 197.400 126.450 198.450 ;
        RECT 121.950 190.950 124.050 193.050 ;
        RECT 115.950 187.950 118.050 190.050 ;
        RECT 98.400 181.350 99.600 183.000 ;
        RECT 104.400 181.350 105.600 183.600 ;
        RECT 109.950 181.950 112.050 184.050 ;
        RECT 115.950 182.100 118.050 184.200 ;
        RECT 122.400 183.600 123.450 190.950 ;
        RECT 125.400 187.050 126.450 197.400 ;
        RECT 127.950 196.950 130.050 199.050 ;
        RECT 124.950 184.950 127.050 187.050 ;
        RECT 128.400 184.050 129.450 196.950 ;
        RECT 134.400 193.050 135.450 209.400 ;
        RECT 139.950 202.950 142.050 205.050 ;
        RECT 140.400 199.050 141.450 202.950 ;
        RECT 139.950 196.950 142.050 199.050 ;
        RECT 133.950 190.950 136.050 193.050 ;
        RECT 130.950 184.950 133.050 187.050 ;
        RECT 94.950 178.950 97.050 181.050 ;
        RECT 97.950 178.950 100.050 181.050 ;
        RECT 100.950 178.950 103.050 181.050 ;
        RECT 103.950 178.950 106.050 181.050 ;
        RECT 95.400 176.400 96.600 178.650 ;
        RECT 101.400 176.400 102.600 178.650 ;
        RECT 95.400 166.050 96.450 176.400 ;
        RECT 101.400 169.050 102.450 176.400 ;
        RECT 100.950 166.950 103.050 169.050 ;
        RECT 94.950 163.950 97.050 166.050 ;
        RECT 110.400 151.050 111.450 181.950 ;
        RECT 116.400 181.350 117.600 182.100 ;
        RECT 122.400 181.350 123.600 183.600 ;
        RECT 127.950 181.950 130.050 184.050 ;
        RECT 115.950 178.950 118.050 181.050 ;
        RECT 118.950 178.950 121.050 181.050 ;
        RECT 121.950 178.950 124.050 181.050 ;
        RECT 124.950 178.950 127.050 181.050 ;
        RECT 119.400 177.000 120.600 178.650 ;
        RECT 125.400 177.900 126.600 178.650 ;
        RECT 118.950 172.950 121.050 177.000 ;
        RECT 124.950 175.800 127.050 177.900 ;
        RECT 131.400 175.050 132.450 184.950 ;
        RECT 140.400 183.600 141.450 196.950 ;
        RECT 140.400 181.350 141.600 183.600 ;
        RECT 143.400 183.450 144.450 235.950 ;
        RECT 160.950 223.950 163.050 226.050 ;
        RECT 151.950 220.950 154.050 223.050 ;
        RECT 152.400 216.600 153.450 220.950 ;
        RECT 152.400 214.350 153.600 216.600 ;
        RECT 148.950 211.950 151.050 214.050 ;
        RECT 151.950 211.950 154.050 214.050 ;
        RECT 154.950 211.950 157.050 214.050 ;
        RECT 149.400 210.000 150.600 211.650 ;
        RECT 148.950 205.950 151.050 210.000 ;
        RECT 155.400 209.400 156.600 211.650 ;
        RECT 155.400 196.050 156.450 209.400 ;
        RECT 161.400 205.050 162.450 223.950 ;
        RECT 167.400 216.600 168.450 235.950 ;
        RECT 172.950 220.950 175.050 223.050 ;
        RECT 173.400 216.600 174.450 220.950 ;
        RECT 167.400 214.350 168.600 216.600 ;
        RECT 173.400 214.350 174.600 216.600 ;
        RECT 166.950 211.950 169.050 214.050 ;
        RECT 169.950 211.950 172.050 214.050 ;
        RECT 172.950 211.950 175.050 214.050 ;
        RECT 170.400 210.000 171.600 211.650 ;
        RECT 163.950 205.950 166.050 208.050 ;
        RECT 169.950 205.950 172.050 210.000 ;
        RECT 179.400 208.050 180.450 254.400 ;
        RECT 182.400 254.400 183.600 256.650 ;
        RECT 188.400 255.900 189.600 256.650 ;
        RECT 182.400 250.050 183.450 254.400 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 197.400 250.050 198.450 262.950 ;
        RECT 203.400 261.600 204.450 274.950 ;
        RECT 203.400 259.350 204.600 261.600 ;
        RECT 202.950 256.950 205.050 259.050 ;
        RECT 205.950 256.950 208.050 259.050 ;
        RECT 206.400 256.050 207.600 256.650 ;
        RECT 206.400 254.400 211.050 256.050 ;
        RECT 207.000 253.950 211.050 254.400 ;
        RECT 181.950 247.950 184.050 250.050 ;
        RECT 196.950 247.950 199.050 250.050 ;
        RECT 212.400 247.050 213.450 277.950 ;
        RECT 215.400 262.050 216.450 280.950 ;
        RECT 221.400 280.050 222.450 286.950 ;
        RECT 220.950 277.950 223.050 280.050 ;
        RECT 224.400 274.050 225.450 293.100 ;
        RECT 230.400 292.350 231.600 294.600 ;
        RECT 244.950 292.950 247.050 295.050 ;
        RECT 247.950 293.100 250.050 295.200 ;
        RECT 254.400 294.600 255.450 301.950 ;
        RECT 260.400 298.050 261.450 322.950 ;
        RECT 266.400 319.050 267.450 331.800 ;
        RECT 275.400 331.050 276.450 352.950 ;
        RECT 280.950 343.950 283.050 346.050 ;
        RECT 287.400 345.450 288.450 361.950 ;
        RECT 290.550 359.700 291.750 372.600 ;
        RECT 295.950 367.950 298.050 370.050 ;
        RECT 296.400 366.900 297.600 367.650 ;
        RECT 302.400 366.900 303.450 418.950 ;
        RECT 305.400 418.050 306.450 424.950 ;
        RECT 308.400 421.050 309.450 433.950 ;
        RECT 311.400 430.050 312.450 443.400 ;
        RECT 314.400 436.050 315.450 520.950 ;
        RECT 317.400 505.050 318.450 521.400 ;
        RECT 325.950 520.950 328.050 523.050 ;
        RECT 332.400 521.400 333.600 523.650 ;
        RECT 338.400 521.400 339.600 523.650 ;
        RECT 332.400 519.450 333.450 521.400 ;
        RECT 332.400 518.400 336.450 519.450 ;
        RECT 316.950 502.950 319.050 505.050 ;
        RECT 325.050 501.300 327.150 503.400 ;
        RECT 319.800 490.950 321.900 493.050 ;
        RECT 320.400 489.900 321.600 490.650 ;
        RECT 319.950 487.800 322.050 489.900 ;
        RECT 325.650 482.700 326.850 501.300 ;
        RECT 328.950 490.950 331.050 493.050 ;
        RECT 329.400 489.000 330.600 490.650 ;
        RECT 328.950 484.950 331.050 489.000 ;
        RECT 322.650 481.500 326.850 482.700 ;
        RECT 322.650 480.600 324.750 481.500 ;
        RECT 329.400 478.050 330.450 484.950 ;
        RECT 328.950 475.950 331.050 478.050 ;
        RECT 335.400 463.050 336.450 518.400 ;
        RECT 338.400 493.050 339.450 521.400 ;
        RECT 347.400 514.050 348.450 527.100 ;
        RECT 359.400 526.350 360.600 527.100 ;
        RECT 353.400 523.950 355.500 526.050 ;
        RECT 358.800 523.950 360.900 526.050 ;
        RECT 353.400 522.900 354.600 523.650 ;
        RECT 362.400 522.900 363.450 535.950 ;
        RECT 425.250 535.500 427.350 536.400 ;
        RECT 433.950 535.950 436.050 538.050 ;
        RECT 440.550 537.300 442.650 539.400 ;
        RECT 423.150 534.300 427.350 535.500 ;
        RECT 364.950 526.950 367.050 529.050 ;
        RECT 370.950 527.100 373.050 532.050 ;
        RECT 376.950 527.100 379.050 529.200 ;
        RECT 382.950 527.100 385.050 529.200 ;
        RECT 388.950 528.000 391.050 532.050 ;
        RECT 352.950 520.800 355.050 522.900 ;
        RECT 361.950 520.800 364.050 522.900 ;
        RECT 346.950 511.950 349.050 514.050 ;
        RECT 365.400 507.450 366.450 526.950 ;
        RECT 371.400 526.350 372.600 527.100 ;
        RECT 377.400 526.350 378.600 527.100 ;
        RECT 370.950 523.950 373.050 526.050 ;
        RECT 373.950 523.950 376.050 526.050 ;
        RECT 376.950 523.950 379.050 526.050 ;
        RECT 374.400 521.400 375.600 523.650 ;
        RECT 374.400 511.050 375.450 521.400 ;
        RECT 373.950 508.950 376.050 511.050 ;
        RECT 365.400 506.400 369.450 507.450 ;
        RECT 337.950 490.950 340.050 493.050 ;
        RECT 346.800 490.950 348.900 493.050 ;
        RECT 364.800 490.950 366.900 493.050 ;
        RECT 365.400 489.000 366.600 490.650 ;
        RECT 364.950 484.950 367.050 489.000 ;
        RECT 346.950 466.950 349.050 469.050 ;
        RECT 334.950 460.950 337.050 463.050 ;
        RECT 328.950 454.950 331.050 457.050 ;
        RECT 334.950 454.950 337.050 457.050 ;
        RECT 322.950 450.000 325.050 454.050 ;
        RECT 329.400 450.600 330.450 454.950 ;
        RECT 323.400 448.350 324.600 450.000 ;
        RECT 329.400 448.350 330.600 450.600 ;
        RECT 322.950 445.950 325.050 448.050 ;
        RECT 325.950 445.950 328.050 448.050 ;
        RECT 328.950 445.950 331.050 448.050 ;
        RECT 326.400 444.900 327.600 445.650 ;
        RECT 335.400 444.900 336.450 454.950 ;
        RECT 340.950 450.000 343.050 454.050 ;
        RECT 347.400 450.600 348.450 466.950 ;
        RECT 358.350 459.300 360.450 461.400 ;
        RECT 359.250 452.700 360.450 459.300 ;
        RECT 358.350 450.600 360.450 452.700 ;
        RECT 361.950 451.950 364.050 454.050 ;
        RECT 341.400 448.350 342.600 450.000 ;
        RECT 347.400 448.350 348.600 450.600 ;
        RECT 340.950 445.950 343.050 448.050 ;
        RECT 343.950 445.950 346.050 448.050 ;
        RECT 346.950 445.950 349.050 448.050 ;
        RECT 352.950 445.950 355.050 448.050 ;
        RECT 325.950 442.800 328.050 444.900 ;
        RECT 334.950 442.800 337.050 444.900 ;
        RECT 344.400 443.400 345.600 445.650 ;
        RECT 353.400 444.900 354.600 445.650 ;
        RECT 344.400 439.050 345.450 443.400 ;
        RECT 352.950 442.800 355.050 444.900 ;
        RECT 343.950 436.950 346.050 439.050 ;
        RECT 359.250 437.700 360.450 450.600 ;
        RECT 313.950 433.950 316.050 436.050 ;
        RECT 358.350 435.600 360.450 437.700 ;
        RECT 362.400 430.050 363.450 451.950 ;
        RECT 310.950 427.950 313.050 430.050 ;
        RECT 355.950 427.950 358.050 430.050 ;
        RECT 361.950 427.950 364.050 430.050 ;
        RECT 313.950 424.950 316.050 427.050 ;
        RECT 307.950 418.950 310.050 421.050 ;
        RECT 304.950 415.950 307.050 418.050 ;
        RECT 308.400 417.600 309.450 418.950 ;
        RECT 314.400 417.600 315.450 424.950 ;
        RECT 356.400 424.050 357.450 427.950 ;
        RECT 355.950 421.950 358.050 424.050 ;
        RECT 361.350 423.300 363.450 425.400 ;
        RECT 322.950 418.950 325.050 421.050 ;
        RECT 308.400 415.350 309.600 417.600 ;
        RECT 314.400 415.350 315.600 417.600 ;
        RECT 307.950 412.950 310.050 415.050 ;
        RECT 310.950 412.950 313.050 415.050 ;
        RECT 313.950 412.950 316.050 415.050 ;
        RECT 316.950 412.950 319.050 415.050 ;
        RECT 311.400 411.900 312.600 412.650 ;
        RECT 317.400 412.050 318.600 412.650 ;
        RECT 304.950 409.800 307.050 411.900 ;
        RECT 310.950 409.800 313.050 411.900 ;
        RECT 317.400 410.400 322.050 412.050 ;
        RECT 323.400 411.900 324.450 418.950 ;
        RECT 325.950 415.950 328.050 421.050 ;
        RECT 331.950 416.100 334.050 418.200 ;
        RECT 340.950 416.100 343.050 418.200 ;
        RECT 346.950 416.100 349.050 418.200 ;
        RECT 355.950 416.100 358.050 418.200 ;
        RECT 332.400 415.350 333.600 416.100 ;
        RECT 328.950 412.950 331.050 415.050 ;
        RECT 331.950 412.950 334.050 415.050 ;
        RECT 334.950 412.950 337.050 415.050 ;
        RECT 318.000 409.950 322.050 410.400 ;
        RECT 322.950 409.800 325.050 411.900 ;
        RECT 329.400 410.400 330.600 412.650 ;
        RECT 335.400 411.900 336.600 412.650 ;
        RECT 295.950 364.800 298.050 366.900 ;
        RECT 301.950 364.800 304.050 366.900 ;
        RECT 305.400 366.450 306.450 409.800 ;
        RECT 329.400 403.050 330.450 410.400 ;
        RECT 334.950 409.800 337.050 411.900 ;
        RECT 341.400 406.050 342.450 416.100 ;
        RECT 347.400 415.350 348.600 416.100 ;
        RECT 356.400 415.350 357.600 416.100 ;
        RECT 346.950 412.950 349.050 415.050 ;
        RECT 349.950 412.950 352.050 415.050 ;
        RECT 355.950 412.950 358.050 415.050 ;
        RECT 350.400 410.400 351.600 412.650 ;
        RECT 362.250 410.400 363.450 423.300 ;
        RECT 350.400 406.050 351.450 410.400 ;
        RECT 361.350 408.300 363.450 410.400 ;
        RECT 365.400 409.050 366.450 484.950 ;
        RECT 368.400 454.050 369.450 506.400 ;
        RECT 379.350 501.300 381.450 503.400 ;
        RECT 373.950 495.000 376.050 499.050 ;
        RECT 374.400 493.350 375.600 495.000 ;
        RECT 373.950 490.950 376.050 493.050 ;
        RECT 380.250 488.400 381.450 501.300 ;
        RECT 383.400 499.050 384.450 527.100 ;
        RECT 389.400 526.350 390.600 528.000 ;
        RECT 394.950 527.100 397.050 529.200 ;
        RECT 400.950 527.100 403.050 529.200 ;
        RECT 406.950 528.000 409.050 532.050 ;
        RECT 395.400 526.350 396.600 527.100 ;
        RECT 388.950 523.950 391.050 526.050 ;
        RECT 391.950 523.950 394.050 526.050 ;
        RECT 394.950 523.950 397.050 526.050 ;
        RECT 392.400 521.400 393.600 523.650 ;
        RECT 385.950 517.950 388.050 520.050 ;
        RECT 382.950 496.950 385.050 499.050 ;
        RECT 379.350 486.300 381.450 488.400 ;
        RECT 386.400 487.050 387.450 517.950 ;
        RECT 392.400 514.050 393.450 521.400 ;
        RECT 391.950 511.950 394.050 514.050 ;
        RECT 401.400 508.050 402.450 527.100 ;
        RECT 407.400 526.350 408.600 528.000 ;
        RECT 412.950 527.100 415.050 529.200 ;
        RECT 418.950 527.100 421.050 529.200 ;
        RECT 413.400 526.350 414.600 527.100 ;
        RECT 419.400 526.350 420.600 527.100 ;
        RECT 406.950 523.950 409.050 526.050 ;
        RECT 409.950 523.950 412.050 526.050 ;
        RECT 412.950 523.950 415.050 526.050 ;
        RECT 418.950 523.950 421.050 526.050 ;
        RECT 410.400 521.400 411.600 523.650 ;
        RECT 410.400 517.050 411.450 521.400 ;
        RECT 415.950 520.950 418.050 523.050 ;
        RECT 409.950 514.950 412.050 517.050 ;
        RECT 416.400 514.050 417.450 520.950 ;
        RECT 423.150 515.700 424.350 534.300 ;
        RECT 440.550 530.700 441.750 537.300 ;
        RECT 454.950 535.950 457.050 538.050 ;
        RECT 427.950 527.100 430.050 529.200 ;
        RECT 433.950 527.100 436.050 529.200 ;
        RECT 440.550 528.600 442.650 530.700 ;
        RECT 455.400 529.200 456.450 535.950 ;
        RECT 428.400 526.350 429.600 527.100 ;
        RECT 428.100 523.950 430.200 526.050 ;
        RECT 434.400 520.050 435.450 527.100 ;
        RECT 433.950 517.950 436.050 520.050 ;
        RECT 415.950 511.950 418.050 514.050 ;
        RECT 422.850 513.600 424.950 515.700 ;
        RECT 400.950 505.950 403.050 508.050 ;
        RECT 397.050 501.300 399.150 503.400 ;
        RECT 391.800 490.950 393.900 493.050 ;
        RECT 392.400 489.900 393.600 490.650 ;
        RECT 391.950 487.800 394.050 489.900 ;
        RECT 385.950 486.450 388.050 487.050 ;
        RECT 380.250 479.700 381.450 486.300 ;
        RECT 379.350 477.600 381.450 479.700 ;
        RECT 383.400 485.400 388.050 486.450 ;
        RECT 373.650 457.500 375.750 458.400 ;
        RECT 373.650 456.300 377.850 457.500 ;
        RECT 367.950 451.950 370.050 454.050 ;
        RECT 370.950 449.100 373.050 451.200 ;
        RECT 371.400 448.350 372.600 449.100 ;
        RECT 370.800 445.950 372.900 448.050 ;
        RECT 376.650 437.700 377.850 456.300 ;
        RECT 380.400 450.450 381.600 450.600 ;
        RECT 383.400 450.450 384.450 485.400 ;
        RECT 385.950 484.950 388.050 485.400 ;
        RECT 397.650 482.700 398.850 501.300 ;
        RECT 406.950 499.950 409.050 502.050 ;
        RECT 407.400 493.050 408.450 499.950 ;
        RECT 409.950 496.950 412.050 499.050 ;
        RECT 400.950 490.950 403.050 493.050 ;
        RECT 406.950 490.950 409.050 493.050 ;
        RECT 401.400 489.000 402.600 490.650 ;
        RECT 410.400 490.050 411.450 496.950 ;
        RECT 418.950 494.100 421.050 496.200 ;
        RECT 424.950 494.100 427.050 496.200 ;
        RECT 430.950 495.450 433.050 496.200 ;
        RECT 434.400 495.450 435.450 517.950 ;
        RECT 440.550 515.700 441.750 528.600 ;
        RECT 454.950 527.100 457.050 529.200 ;
        RECT 445.950 523.950 448.050 526.050 ;
        RECT 446.400 522.900 447.600 523.650 ;
        RECT 455.400 523.050 456.450 527.100 ;
        RECT 445.950 520.800 448.050 522.900 ;
        RECT 454.950 520.950 457.050 523.050 ;
        RECT 440.550 513.600 442.650 515.700 ;
        RECT 458.400 511.050 459.450 547.950 ;
        RECT 479.400 547.050 480.450 566.400 ;
        RECT 499.950 565.800 502.050 567.900 ;
        RECT 472.950 544.950 475.050 547.050 ;
        RECT 478.950 544.950 481.050 547.050 ;
        RECT 463.950 527.100 466.050 529.200 ;
        RECT 464.400 526.350 465.600 527.100 ;
        RECT 463.950 523.950 466.050 526.050 ;
        RECT 466.950 523.950 469.050 526.050 ;
        RECT 467.400 521.400 468.600 523.650 ;
        RECT 467.400 519.450 468.450 521.400 ;
        RECT 464.400 518.400 468.450 519.450 ;
        RECT 445.950 508.950 448.050 511.050 ;
        RECT 457.950 508.950 460.050 511.050 ;
        RECT 439.950 499.950 442.050 502.050 ;
        RECT 430.950 494.400 435.450 495.450 ;
        RECT 440.400 495.600 441.450 499.950 ;
        RECT 446.400 495.600 447.450 508.950 ;
        RECT 457.350 501.300 459.450 503.400 ;
        RECT 430.950 494.100 433.050 494.400 ;
        RECT 419.400 493.350 420.600 494.100 ;
        RECT 425.400 493.350 426.600 494.100 ;
        RECT 415.950 490.950 418.050 493.050 ;
        RECT 418.950 490.950 421.050 493.050 ;
        RECT 421.950 490.950 424.050 493.050 ;
        RECT 424.950 490.950 427.050 493.050 ;
        RECT 400.950 484.950 403.050 489.000 ;
        RECT 409.950 487.950 412.050 490.050 ;
        RECT 416.400 489.900 417.600 490.650 ;
        RECT 415.950 487.800 418.050 489.900 ;
        RECT 422.400 488.400 423.600 490.650 ;
        RECT 394.650 481.500 398.850 482.700 ;
        RECT 394.650 480.600 396.750 481.500 ;
        RECT 422.400 463.050 423.450 488.400 ;
        RECT 400.950 460.950 403.050 463.050 ;
        RECT 421.950 460.950 424.050 463.050 ;
        RECT 394.950 454.950 397.050 457.050 ;
        RECT 380.400 449.400 384.450 450.450 ;
        RECT 395.400 450.600 396.450 454.950 ;
        RECT 401.400 450.600 402.450 460.950 ;
        RECT 380.400 448.350 381.600 449.400 ;
        RECT 395.400 448.350 396.600 450.600 ;
        RECT 401.400 448.350 402.600 450.600 ;
        RECT 409.950 449.100 412.050 451.200 ;
        RECT 415.950 449.100 418.050 451.200 ;
        RECT 421.950 449.100 424.050 451.200 ;
        RECT 379.950 445.950 382.050 448.050 ;
        RECT 394.950 445.950 397.050 448.050 ;
        RECT 397.950 445.950 400.050 448.050 ;
        RECT 400.950 445.950 403.050 448.050 ;
        RECT 403.950 445.950 406.050 448.050 ;
        RECT 398.400 444.900 399.600 445.650 ;
        RECT 397.950 442.800 400.050 444.900 ;
        RECT 404.400 443.400 405.600 445.650 ;
        RECT 410.400 445.050 411.450 449.100 ;
        RECT 416.400 448.350 417.600 449.100 ;
        RECT 422.400 448.350 423.600 449.100 ;
        RECT 415.950 445.950 418.050 448.050 ;
        RECT 418.950 445.950 421.050 448.050 ;
        RECT 421.950 445.950 424.050 448.050 ;
        RECT 424.950 445.950 427.050 448.050 ;
        RECT 404.400 439.050 405.450 443.400 ;
        RECT 409.950 442.950 412.050 445.050 ;
        RECT 419.400 444.900 420.600 445.650 ;
        RECT 425.400 444.900 426.600 445.650 ;
        RECT 418.950 442.800 421.050 444.900 ;
        RECT 424.950 442.800 427.050 444.900 ;
        RECT 431.400 439.050 432.450 494.100 ;
        RECT 440.400 493.350 441.600 495.600 ;
        RECT 446.400 493.350 447.600 495.600 ;
        RECT 451.950 494.100 454.050 496.200 ;
        RECT 452.400 493.350 453.600 494.100 ;
        RECT 436.950 490.950 439.050 493.050 ;
        RECT 439.950 490.950 442.050 493.050 ;
        RECT 442.950 490.950 445.050 493.050 ;
        RECT 445.950 490.950 448.050 493.050 ;
        RECT 451.950 490.950 454.050 493.050 ;
        RECT 437.400 489.900 438.600 490.650 ;
        RECT 436.950 487.800 439.050 489.900 ;
        RECT 443.400 488.400 444.600 490.650 ;
        RECT 458.250 488.400 459.450 501.300 ;
        RECT 460.950 494.100 463.050 496.200 ;
        RECT 443.400 486.450 444.450 488.400 ;
        RECT 440.400 485.400 444.450 486.450 ;
        RECT 457.350 486.300 459.450 488.400 ;
        RECT 433.950 454.950 436.050 457.050 ;
        RECT 434.400 444.900 435.450 454.950 ;
        RECT 440.400 451.200 441.450 485.400 ;
        RECT 458.250 479.700 459.450 486.300 ;
        RECT 461.400 484.050 462.450 494.100 ;
        RECT 460.950 481.950 463.050 484.050 ;
        RECT 457.350 477.600 459.450 479.700 ;
        RECT 461.400 475.050 462.450 481.950 ;
        RECT 460.950 472.950 463.050 475.050 ;
        RECT 460.950 462.450 463.050 463.050 ;
        RECT 464.400 462.450 465.450 518.400 ;
        RECT 473.400 511.050 474.450 544.950 ;
        RECT 503.400 541.050 504.450 590.400 ;
        RECT 524.400 589.050 525.450 599.400 ;
        RECT 505.950 586.950 508.050 589.050 ;
        RECT 523.950 586.950 526.050 589.050 ;
        RECT 506.400 583.050 507.450 586.950 ;
        RECT 520.950 583.950 523.050 586.050 ;
        RECT 505.950 580.950 508.050 583.050 ;
        RECT 505.950 571.950 508.050 574.050 ;
        RECT 514.950 572.100 517.050 574.200 ;
        RECT 521.400 573.450 522.450 583.950 ;
        RECT 529.350 579.300 531.450 581.400 ;
        RECT 523.950 573.450 526.050 574.200 ;
        RECT 521.400 572.400 526.050 573.450 ;
        RECT 523.950 572.100 526.050 572.400 ;
        RECT 506.400 556.050 507.450 571.950 ;
        RECT 515.400 571.350 516.600 572.100 ;
        RECT 524.400 571.350 525.600 572.100 ;
        RECT 511.950 568.950 514.050 571.050 ;
        RECT 514.950 568.950 517.050 571.050 ;
        RECT 517.950 568.950 520.050 571.050 ;
        RECT 523.950 568.950 526.050 571.050 ;
        RECT 512.400 567.900 513.600 568.650 ;
        RECT 518.400 567.900 519.600 568.650 ;
        RECT 511.950 565.800 514.050 567.900 ;
        RECT 517.950 565.800 520.050 567.900 ;
        RECT 530.250 566.400 531.450 579.300 ;
        RECT 512.400 562.050 513.450 565.800 ;
        RECT 529.350 564.300 531.450 566.400 ;
        RECT 511.950 559.950 514.050 562.050 ;
        RECT 517.950 556.950 520.050 559.050 ;
        RECT 530.250 557.700 531.450 564.300 ;
        RECT 505.950 553.950 508.050 556.050 ;
        RECT 518.400 547.050 519.450 556.950 ;
        RECT 529.350 555.600 531.450 557.700 ;
        RECT 517.950 544.950 520.050 547.050 ;
        RECT 496.350 537.300 498.450 539.400 ;
        RECT 502.950 538.950 505.050 541.050 ;
        RECT 481.950 532.950 484.050 535.050 ;
        RECT 482.400 528.600 483.450 532.950 ;
        RECT 497.250 530.700 498.450 537.300 ;
        RECT 496.350 528.600 498.450 530.700 ;
        RECT 482.400 526.350 483.600 528.600 ;
        RECT 478.950 523.950 481.050 526.050 ;
        RECT 481.950 523.950 484.050 526.050 ;
        RECT 484.950 523.950 487.050 526.050 ;
        RECT 490.950 523.950 493.050 526.050 ;
        RECT 479.400 522.000 480.600 523.650 ;
        RECT 485.400 522.900 486.600 523.650 ;
        RECT 491.400 522.900 492.600 523.650 ;
        RECT 478.950 517.950 481.050 522.000 ;
        RECT 484.950 520.800 487.050 522.900 ;
        RECT 490.950 520.800 493.050 522.900 ;
        RECT 485.400 514.050 486.450 520.800 ;
        RECT 497.250 515.700 498.450 528.600 ;
        RECT 484.950 511.950 487.050 514.050 ;
        RECT 496.350 513.600 498.450 515.700 ;
        RECT 472.950 508.950 475.050 511.050 ;
        RECT 484.950 508.800 487.050 510.900 ;
        RECT 475.050 501.300 477.150 503.400 ;
        RECT 469.800 490.950 471.900 493.050 ;
        RECT 470.400 489.900 471.600 490.650 ;
        RECT 469.950 487.800 472.050 489.900 ;
        RECT 475.650 482.700 476.850 501.300 ;
        RECT 478.950 490.950 481.050 493.050 ;
        RECT 479.400 489.450 480.600 490.650 ;
        RECT 485.400 489.450 486.450 508.800 ;
        RECT 493.950 502.950 496.050 505.050 ;
        RECT 494.400 495.600 495.450 502.950 ;
        RECT 503.400 499.050 504.450 538.950 ;
        RECT 511.650 535.500 513.750 536.400 ;
        RECT 511.650 534.300 515.850 535.500 ;
        RECT 508.950 527.100 511.050 529.200 ;
        RECT 509.400 526.350 510.600 527.100 ;
        RECT 508.800 523.950 510.900 526.050 ;
        RECT 514.650 515.700 515.850 534.300 ;
        RECT 518.400 528.600 519.450 544.950 ;
        RECT 533.400 532.050 534.450 610.950 ;
        RECT 536.400 550.050 537.450 622.950 ;
        RECT 539.400 600.450 540.450 628.950 ;
        RECT 542.400 628.050 543.450 646.950 ;
        RECT 551.400 644.400 552.600 646.650 ;
        RECT 547.950 628.950 550.050 631.050 ;
        RECT 541.950 625.950 544.050 628.050 ;
        RECT 548.400 606.600 549.450 628.950 ;
        RECT 551.400 622.050 552.450 644.400 ;
        RECT 550.950 619.950 553.050 622.050 ;
        RECT 556.950 610.950 559.050 613.050 ;
        RECT 548.400 604.350 549.600 606.600 ;
        RECT 557.400 606.450 558.450 610.950 ;
        RECT 560.400 610.050 561.450 650.100 ;
        RECT 566.400 649.350 567.600 650.100 ;
        RECT 572.400 649.350 573.600 651.600 ;
        RECT 565.950 646.950 568.050 649.050 ;
        RECT 568.950 646.950 571.050 649.050 ;
        RECT 571.950 646.950 574.050 649.050 ;
        RECT 574.950 646.950 577.050 649.050 ;
        RECT 569.400 645.900 570.600 646.650 ;
        RECT 568.950 643.800 571.050 645.900 ;
        RECT 575.400 644.400 576.600 646.650 ;
        RECT 581.400 645.900 582.450 658.950 ;
        RECT 584.400 652.050 585.450 671.400 ;
        RECT 586.950 670.950 589.050 673.050 ;
        RECT 598.950 670.950 604.050 673.050 ;
        RECT 587.400 661.050 588.450 670.950 ;
        RECT 589.950 664.950 592.050 667.050 ;
        RECT 601.950 664.950 604.050 667.050 ;
        RECT 586.950 658.950 589.050 661.050 ;
        RECT 590.400 654.450 591.450 664.950 ;
        RECT 592.950 658.950 595.050 661.050 ;
        RECT 587.400 653.400 591.450 654.450 ;
        RECT 583.950 649.950 586.050 652.050 ;
        RECT 587.400 651.600 588.450 653.400 ;
        RECT 593.400 651.600 594.450 658.950 ;
        RECT 587.400 649.350 588.600 651.600 ;
        RECT 593.400 649.350 594.600 651.600 ;
        RECT 586.950 646.950 589.050 649.050 ;
        RECT 589.950 646.950 592.050 649.050 ;
        RECT 592.950 646.950 595.050 649.050 ;
        RECT 595.950 646.950 598.050 649.050 ;
        RECT 559.950 607.950 562.050 610.050 ;
        RECT 560.400 606.450 561.600 606.600 ;
        RECT 557.400 605.400 561.600 606.450 ;
        RECT 565.950 606.000 568.050 610.050 ;
        RECT 560.400 604.350 561.600 605.400 ;
        RECT 566.400 604.350 567.600 606.000 ;
        RECT 542.400 601.950 544.500 604.050 ;
        RECT 547.800 601.950 549.900 604.050 ;
        RECT 559.950 601.950 562.050 604.050 ;
        RECT 562.950 601.950 565.050 604.050 ;
        RECT 565.950 601.950 568.050 604.050 ;
        RECT 568.950 601.950 571.050 604.050 ;
        RECT 542.400 600.450 543.600 601.650 ;
        RECT 563.400 600.900 564.600 601.650 ;
        RECT 569.400 600.900 570.600 601.650 ;
        RECT 539.400 599.400 543.600 600.450 ;
        RECT 562.950 595.950 565.050 600.900 ;
        RECT 568.950 598.800 571.050 600.900 ;
        RECT 559.950 586.950 562.050 589.050 ;
        RECT 547.050 579.300 549.150 581.400 ;
        RECT 541.800 568.950 543.900 571.050 ;
        RECT 542.400 567.900 543.600 568.650 ;
        RECT 541.950 565.800 544.050 567.900 ;
        RECT 547.650 560.700 548.850 579.300 ;
        RECT 556.950 571.950 559.050 574.050 ;
        RECT 550.950 568.950 553.050 571.050 ;
        RECT 544.650 559.500 548.850 560.700 ;
        RECT 551.400 566.400 552.600 568.650 ;
        RECT 557.400 567.900 558.450 571.950 ;
        RECT 544.650 558.600 546.750 559.500 ;
        RECT 551.400 559.050 552.450 566.400 ;
        RECT 556.950 565.800 559.050 567.900 ;
        RECT 550.950 556.950 553.050 559.050 ;
        RECT 535.950 547.950 538.050 550.050 ;
        RECT 560.400 538.050 561.450 586.950 ;
        RECT 575.400 583.050 576.450 644.400 ;
        RECT 580.950 643.800 583.050 645.900 ;
        RECT 590.400 644.400 591.600 646.650 ;
        RECT 596.400 645.900 597.600 646.650 ;
        RECT 590.400 642.450 591.450 644.400 ;
        RECT 595.950 643.800 598.050 645.900 ;
        RECT 598.950 643.950 601.050 646.050 ;
        RECT 592.950 642.450 595.050 643.050 ;
        RECT 590.400 641.400 595.050 642.450 ;
        RECT 592.950 640.950 595.050 641.400 ;
        RECT 589.950 637.950 592.050 640.050 ;
        RECT 586.950 628.950 589.050 631.050 ;
        RECT 577.950 619.950 580.050 622.050 ;
        RECT 578.400 607.050 579.450 619.950 ;
        RECT 587.400 610.050 588.450 628.950 ;
        RECT 577.950 604.950 580.050 607.050 ;
        RECT 583.950 606.000 586.050 610.050 ;
        RECT 586.950 607.950 589.050 610.050 ;
        RECT 590.400 607.050 591.450 637.950 ;
        RECT 584.400 604.350 585.600 606.000 ;
        RECT 589.950 604.950 592.050 607.050 ;
        RECT 580.950 601.950 583.050 604.050 ;
        RECT 583.950 601.950 586.050 604.050 ;
        RECT 586.950 601.950 589.050 604.050 ;
        RECT 581.400 600.000 582.600 601.650 ;
        RECT 587.400 600.900 588.600 601.650 ;
        RECT 580.950 595.950 583.050 600.000 ;
        RECT 586.950 598.800 589.050 600.900 ;
        RECT 589.950 598.950 592.050 601.050 ;
        RECT 586.950 592.950 589.050 595.050 ;
        RECT 583.950 589.950 586.050 592.050 ;
        RECT 574.950 580.950 577.050 583.050 ;
        RECT 568.950 572.100 571.050 574.200 ;
        RECT 574.950 572.100 577.050 574.200 ;
        RECT 580.950 572.100 583.050 574.200 ;
        RECT 584.400 574.050 585.450 589.950 ;
        RECT 587.400 583.050 588.450 592.950 ;
        RECT 590.400 592.050 591.450 598.950 ;
        RECT 593.400 595.050 594.450 640.950 ;
        RECT 599.400 640.050 600.450 643.950 ;
        RECT 595.950 637.950 598.050 640.050 ;
        RECT 598.950 637.950 601.050 640.050 ;
        RECT 596.400 622.050 597.450 637.950 ;
        RECT 598.950 625.950 601.050 628.050 ;
        RECT 595.950 619.950 598.050 622.050 ;
        RECT 599.400 616.050 600.450 625.950 ;
        RECT 602.400 625.050 603.450 664.950 ;
        RECT 605.400 664.050 606.450 677.400 ;
        RECT 607.950 676.950 610.050 679.050 ;
        RECT 604.950 661.950 607.050 664.050 ;
        RECT 608.400 660.450 609.450 676.950 ;
        RECT 610.950 670.950 613.050 673.050 ;
        RECT 605.400 659.400 609.450 660.450 ;
        RECT 605.400 652.050 606.450 659.400 ;
        RECT 604.950 649.950 607.050 652.050 ;
        RECT 611.400 651.600 612.450 670.950 ;
        RECT 614.400 667.050 615.450 728.400 ;
        RECT 622.950 727.950 625.050 730.050 ;
        RECT 619.800 724.950 621.900 727.050 ;
        RECT 623.400 718.050 624.450 727.950 ;
        RECT 637.800 724.950 639.900 727.050 ;
        RECT 638.400 723.900 639.600 724.650 ;
        RECT 637.950 721.800 640.050 723.900 ;
        RECT 622.950 715.950 625.050 718.050 ;
        RECT 619.500 687.300 621.600 689.400 ;
        RECT 629.100 688.500 631.200 690.600 ;
        RECT 616.950 683.100 619.050 685.200 ;
        RECT 617.400 682.350 618.600 683.100 ;
        RECT 617.100 679.950 619.200 682.050 ;
        RECT 620.400 678.300 621.300 687.300 ;
        RECT 622.800 683.700 624.900 685.800 ;
        RECT 626.400 685.350 627.600 687.600 ;
        RECT 624.000 681.300 624.900 683.700 ;
        RECT 625.800 682.950 627.900 685.050 ;
        RECT 629.700 681.300 630.900 688.500 ;
        RECT 641.400 685.050 642.450 784.950 ;
        RECT 677.400 772.050 678.450 800.400 ;
        RECT 692.400 787.050 693.450 800.400 ;
        RECT 691.950 784.950 694.050 787.050 ;
        RECT 701.400 781.050 702.450 806.100 ;
        RECT 710.400 805.350 711.600 806.100 ;
        RECT 716.400 805.350 717.600 806.100 ;
        RECT 731.400 805.350 732.600 806.100 ;
        RECT 737.400 805.350 738.600 806.100 ;
        RECT 706.950 802.950 709.050 805.050 ;
        RECT 709.950 802.950 712.050 805.050 ;
        RECT 712.950 802.950 715.050 805.050 ;
        RECT 715.950 802.950 718.050 805.050 ;
        RECT 718.950 802.950 721.050 805.050 ;
        RECT 730.950 802.950 733.050 805.050 ;
        RECT 733.950 802.950 736.050 805.050 ;
        RECT 736.950 802.950 739.050 805.050 ;
        RECT 739.950 802.950 742.050 805.050 ;
        RECT 707.400 800.400 708.600 802.650 ;
        RECT 713.400 801.900 714.600 802.650 ;
        RECT 707.400 796.050 708.450 800.400 ;
        RECT 712.950 799.800 715.050 801.900 ;
        RECT 719.400 800.400 720.600 802.650 ;
        RECT 734.400 800.400 735.600 802.650 ;
        RECT 740.400 801.900 741.600 802.650 ;
        RECT 706.950 793.950 709.050 796.050 ;
        RECT 719.400 793.050 720.450 800.400 ;
        RECT 718.950 790.950 721.050 793.050 ;
        RECT 727.950 784.950 730.050 787.050 ;
        RECT 700.950 778.950 703.050 781.050 ;
        RECT 676.950 769.950 679.050 772.050 ;
        RECT 691.950 769.950 694.050 772.050 ;
        RECT 682.950 766.950 685.050 769.050 ;
        RECT 643.950 763.950 646.050 766.050 ;
        RECT 644.400 724.050 645.450 763.950 ;
        RECT 649.950 761.100 652.050 763.200 ;
        RECT 655.950 761.100 658.050 763.200 ;
        RECT 650.400 760.350 651.600 761.100 ;
        RECT 656.400 760.350 657.600 761.100 ;
        RECT 664.950 760.950 667.050 763.050 ;
        RECT 673.950 761.100 676.050 763.200 ;
        RECT 649.950 757.950 652.050 760.050 ;
        RECT 652.950 757.950 655.050 760.050 ;
        RECT 655.950 757.950 658.050 760.050 ;
        RECT 658.950 757.950 661.050 760.050 ;
        RECT 653.400 755.400 654.600 757.650 ;
        RECT 659.400 756.450 660.600 757.650 ;
        RECT 665.400 756.450 666.450 760.950 ;
        RECT 674.400 760.350 675.600 761.100 ;
        RECT 670.950 757.950 673.050 760.050 ;
        RECT 673.950 757.950 676.050 760.050 ;
        RECT 676.950 757.950 679.050 760.050 ;
        RECT 659.400 755.400 666.450 756.450 ;
        RECT 671.400 755.400 672.600 757.650 ;
        RECT 677.400 756.450 678.600 757.650 ;
        RECT 683.400 756.450 684.450 766.950 ;
        RECT 692.400 762.600 693.450 769.950 ;
        RECT 692.400 760.350 693.600 762.600 ;
        RECT 697.950 761.100 700.050 763.200 ;
        RECT 688.950 757.950 691.050 760.050 ;
        RECT 691.950 757.950 694.050 760.050 ;
        RECT 677.400 755.400 684.450 756.450 ;
        RECT 653.400 751.050 654.450 755.400 ;
        RECT 652.950 748.950 655.050 751.050 ;
        RECT 671.400 739.050 672.450 755.400 ;
        RECT 685.950 754.950 688.050 757.050 ;
        RECT 689.400 755.400 690.600 757.650 ;
        RECT 676.950 742.950 679.050 745.050 ;
        RECT 670.950 736.950 673.050 739.050 ;
        RECT 667.950 730.950 670.050 733.050 ;
        RECT 652.950 728.100 655.050 730.200 ;
        RECT 658.950 728.100 661.050 730.200 ;
        RECT 653.400 727.350 654.600 728.100 ;
        RECT 659.400 727.350 660.600 728.100 ;
        RECT 652.950 724.950 655.050 727.050 ;
        RECT 655.950 724.950 658.050 727.050 ;
        RECT 658.950 724.950 661.050 727.050 ;
        RECT 661.950 724.950 664.050 727.050 ;
        RECT 643.950 721.950 646.050 724.050 ;
        RECT 656.400 723.000 657.600 724.650 ;
        RECT 644.400 712.050 645.450 721.950 ;
        RECT 655.950 718.950 658.050 723.000 ;
        RECT 662.400 722.400 663.600 724.650 ;
        RECT 662.400 715.050 663.450 722.400 ;
        RECT 661.950 712.950 664.050 715.050 ;
        RECT 643.950 709.950 646.050 712.050 ;
        RECT 643.950 691.950 646.050 694.050 ;
        RECT 634.950 682.950 637.050 685.050 ;
        RECT 640.950 682.950 643.050 685.050 ;
        RECT 644.400 684.600 645.450 691.950 ;
        RECT 662.400 691.050 663.450 712.950 ;
        RECT 668.400 709.050 669.450 730.950 ;
        RECT 677.400 729.600 678.450 742.950 ;
        RECT 682.950 736.950 685.050 739.050 ;
        RECT 677.400 727.350 678.600 729.600 ;
        RECT 673.950 724.950 676.050 727.050 ;
        RECT 676.950 724.950 679.050 727.050 ;
        RECT 674.400 723.000 675.600 724.650 ;
        RECT 673.950 718.950 676.050 723.000 ;
        RECT 683.400 715.050 684.450 736.950 ;
        RECT 686.400 733.050 687.450 754.950 ;
        RECT 689.400 739.050 690.450 755.400 ;
        RECT 698.400 742.050 699.450 761.100 ;
        RECT 701.400 757.050 702.450 778.950 ;
        RECT 721.950 772.950 724.050 775.050 ;
        RECT 712.950 769.950 715.050 772.050 ;
        RECT 713.400 766.050 714.450 769.950 ;
        RECT 722.400 769.050 723.450 772.950 ;
        RECT 724.950 769.950 727.050 772.050 ;
        RECT 721.950 766.950 724.050 769.050 ;
        RECT 725.400 766.050 726.450 769.950 ;
        RECT 712.950 763.950 715.050 766.050 ;
        RECT 724.950 763.950 727.050 766.050 ;
        RECT 706.950 761.100 709.050 763.200 ;
        RECT 713.400 762.600 714.450 763.950 ;
        RECT 728.400 763.200 729.450 784.950 ;
        RECT 734.400 781.050 735.450 800.400 ;
        RECT 739.950 799.800 742.050 801.900 ;
        RECT 746.400 801.450 747.450 806.100 ;
        RECT 758.400 805.350 759.600 806.100 ;
        RECT 755.100 802.950 757.200 805.050 ;
        RECT 758.400 802.950 760.500 805.050 ;
        RECT 763.800 802.950 765.900 805.050 ;
        RECT 755.400 801.900 756.600 802.650 ;
        RECT 743.400 800.400 747.450 801.450 ;
        RECT 733.950 778.950 736.050 781.050 ;
        RECT 736.950 772.950 739.050 775.050 ;
        RECT 707.400 760.350 708.600 761.100 ;
        RECT 713.400 760.350 714.600 762.600 ;
        RECT 721.950 760.950 724.050 763.050 ;
        RECT 727.950 761.100 730.050 763.200 ;
        RECT 706.950 757.950 709.050 760.050 ;
        RECT 709.950 757.950 712.050 760.050 ;
        RECT 712.950 757.950 715.050 760.050 ;
        RECT 715.950 757.950 718.050 760.050 ;
        RECT 700.950 754.950 703.050 757.050 ;
        RECT 710.400 755.400 711.600 757.650 ;
        RECT 716.400 756.900 717.600 757.650 ;
        RECT 722.400 756.900 723.450 760.950 ;
        RECT 728.400 760.350 729.600 761.100 ;
        RECT 727.950 757.950 730.050 760.050 ;
        RECT 730.950 757.950 733.050 760.050 ;
        RECT 731.400 756.900 732.600 757.650 ;
        RECT 737.400 756.900 738.450 772.950 ;
        RECT 743.400 763.200 744.450 800.400 ;
        RECT 754.950 799.800 757.050 801.900 ;
        RECT 764.400 800.400 765.600 802.650 ;
        RECT 764.400 793.050 765.450 800.400 ;
        RECT 763.950 790.950 766.050 793.050 ;
        RECT 770.400 787.050 771.450 806.100 ;
        RECT 776.400 805.350 777.600 806.100 ;
        RECT 782.400 805.350 783.600 806.100 ;
        RECT 800.400 805.350 801.600 806.400 ;
        RECT 775.950 802.950 778.050 805.050 ;
        RECT 778.950 802.950 781.050 805.050 ;
        RECT 781.950 802.950 784.050 805.050 ;
        RECT 784.950 802.950 787.050 805.050 ;
        RECT 796.950 802.950 799.050 805.050 ;
        RECT 799.950 802.950 802.050 805.050 ;
        RECT 779.400 800.400 780.600 802.650 ;
        RECT 785.400 801.900 786.600 802.650 ;
        RECT 797.400 801.900 798.600 802.650 ;
        RECT 806.400 802.050 807.450 806.400 ;
        RECT 818.400 805.350 819.600 807.600 ;
        RECT 826.950 806.100 829.050 808.200 ;
        RECT 832.950 806.100 835.050 808.200 ;
        RECT 838.950 806.100 841.050 808.200 ;
        RECT 844.950 806.100 847.050 808.200 ;
        RECT 854.400 807.600 855.450 811.950 ;
        RECT 812.100 802.950 814.200 805.050 ;
        RECT 817.500 802.950 819.600 805.050 ;
        RECT 820.800 802.950 822.900 805.050 ;
        RECT 769.950 784.950 772.050 787.050 ;
        RECT 772.950 775.950 775.050 778.050 ;
        RECT 751.950 763.950 754.050 766.050 ;
        RECT 742.950 761.100 745.050 763.200 ;
        RECT 743.400 760.350 744.600 761.100 ;
        RECT 742.950 757.950 745.050 760.050 ;
        RECT 745.950 757.950 748.050 760.050 ;
        RECT 710.400 751.050 711.450 755.400 ;
        RECT 715.950 754.800 718.050 756.900 ;
        RECT 721.950 754.800 724.050 756.900 ;
        RECT 730.950 754.800 733.050 756.900 ;
        RECT 736.800 754.800 738.900 756.900 ;
        RECT 739.950 754.950 742.050 757.050 ;
        RECT 746.400 756.900 747.600 757.650 ;
        RECT 752.400 756.900 753.450 763.950 ;
        RECT 760.950 761.100 763.050 763.200 ;
        RECT 766.950 761.100 769.050 766.050 ;
        RECT 761.400 760.350 762.600 761.100 ;
        RECT 767.400 760.350 768.600 761.100 ;
        RECT 757.950 757.950 760.050 760.050 ;
        RECT 760.950 757.950 763.050 760.050 ;
        RECT 763.950 757.950 766.050 760.050 ;
        RECT 766.950 757.950 769.050 760.050 ;
        RECT 709.950 748.950 712.050 751.050 ;
        RECT 697.950 739.950 700.050 742.050 ;
        RECT 688.950 736.950 691.050 739.050 ;
        RECT 691.950 733.950 694.050 736.050 ;
        RECT 685.950 730.950 688.050 733.050 ;
        RECT 692.400 729.600 693.450 733.950 ;
        RECT 698.400 729.600 699.450 739.950 ;
        RECT 703.950 733.950 706.050 736.050 ;
        RECT 715.950 733.950 718.050 736.050 ;
        RECT 692.400 727.350 693.600 729.600 ;
        RECT 698.400 727.350 699.600 729.600 ;
        RECT 688.950 724.950 691.050 727.050 ;
        RECT 691.950 724.950 694.050 727.050 ;
        RECT 694.950 724.950 697.050 727.050 ;
        RECT 697.950 724.950 700.050 727.050 ;
        RECT 689.400 723.450 690.600 724.650 ;
        RECT 686.400 722.400 690.600 723.450 ;
        RECT 695.400 723.000 696.600 724.650 ;
        RECT 704.400 724.050 705.450 733.950 ;
        RECT 709.950 729.000 712.050 733.050 ;
        RECT 716.400 729.600 717.450 733.950 ;
        RECT 722.400 733.050 723.450 754.800 ;
        RECT 736.950 748.950 739.050 751.050 ;
        RECT 737.400 742.050 738.450 748.950 ;
        RECT 736.950 739.950 739.050 742.050 ;
        RECT 725.850 735.300 727.950 737.400 ;
        RECT 721.950 730.950 724.050 733.050 ;
        RECT 710.400 727.350 711.600 729.000 ;
        RECT 716.400 727.350 717.600 729.600 ;
        RECT 709.950 724.950 712.050 727.050 ;
        RECT 712.950 724.950 715.050 727.050 ;
        RECT 715.950 724.950 718.050 727.050 ;
        RECT 721.950 724.950 724.050 727.050 ;
        RECT 682.950 712.950 685.050 715.050 ;
        RECT 667.950 706.950 670.050 709.050 ;
        RECT 673.950 706.950 676.050 709.050 ;
        RECT 670.950 697.950 673.050 700.050 ;
        RECT 667.950 691.950 670.050 694.050 ;
        RECT 661.950 688.950 664.050 691.050 ;
        RECT 664.950 688.950 667.050 691.050 ;
        RECT 665.400 685.200 666.450 688.950 ;
        RECT 624.000 680.100 630.900 681.300 ;
        RECT 627.000 678.300 629.100 679.200 ;
        RECT 620.400 677.100 629.100 678.300 ;
        RECT 621.900 675.300 624.000 677.100 ;
        RECT 625.800 674.100 627.900 676.200 ;
        RECT 630.000 674.700 630.900 680.100 ;
        RECT 631.800 679.950 633.900 682.050 ;
        RECT 632.400 678.900 633.600 679.650 ;
        RECT 631.950 676.800 634.050 678.900 ;
        RECT 626.400 671.550 627.600 673.800 ;
        RECT 629.100 672.600 631.200 674.700 ;
        RECT 613.950 664.950 616.050 667.050 ;
        RECT 626.400 663.450 627.450 671.550 ;
        RECT 626.400 662.400 630.450 663.450 ;
        RECT 616.950 658.950 619.050 661.050 ;
        RECT 617.400 655.050 618.450 658.950 ;
        RECT 625.350 657.300 627.450 659.400 ;
        RECT 616.950 652.950 619.050 655.050 ;
        RECT 611.400 649.350 612.600 651.600 ;
        RECT 619.950 650.100 622.050 652.200 ;
        RECT 620.400 649.350 621.600 650.100 ;
        RECT 607.950 646.950 610.050 649.050 ;
        RECT 610.950 646.950 613.050 649.050 ;
        RECT 613.950 646.950 616.050 649.050 ;
        RECT 619.950 646.950 622.050 649.050 ;
        RECT 608.400 645.000 609.600 646.650 ;
        RECT 614.400 645.900 615.600 646.650 ;
        RECT 607.950 640.950 610.050 645.000 ;
        RECT 613.950 643.800 616.050 645.900 ;
        RECT 626.250 644.400 627.450 657.300 ;
        RECT 614.400 640.050 615.450 643.800 ;
        RECT 625.350 642.300 627.450 644.400 ;
        RECT 607.950 637.800 610.050 639.900 ;
        RECT 613.950 637.950 616.050 640.050 ;
        RECT 604.950 634.950 607.050 637.050 ;
        RECT 601.950 622.950 604.050 625.050 ;
        RECT 598.950 613.950 601.050 616.050 ;
        RECT 595.950 610.950 598.050 613.050 ;
        RECT 596.400 607.050 597.450 610.950 ;
        RECT 595.950 604.950 598.050 607.050 ;
        RECT 598.950 606.000 601.050 610.050 ;
        RECT 605.400 607.200 606.450 634.950 ;
        RECT 608.400 619.050 609.450 637.800 ;
        RECT 626.250 635.700 627.450 642.300 ;
        RECT 625.350 633.600 627.450 635.700 ;
        RECT 607.950 616.950 610.050 619.050 ;
        RECT 622.950 616.950 625.050 619.050 ;
        RECT 617.250 613.500 619.350 614.400 ;
        RECT 615.150 612.300 619.350 613.500 ;
        RECT 599.400 604.350 600.600 606.000 ;
        RECT 604.950 605.100 607.050 607.200 ;
        RECT 610.950 605.100 613.050 607.200 ;
        RECT 605.400 604.350 606.600 605.100 ;
        RECT 611.400 604.350 612.600 605.100 ;
        RECT 598.950 601.950 601.050 604.050 ;
        RECT 601.950 601.950 604.050 604.050 ;
        RECT 604.950 601.950 607.050 604.050 ;
        RECT 610.950 601.950 613.050 604.050 ;
        RECT 602.400 599.400 603.600 601.650 ;
        RECT 592.950 592.950 595.050 595.050 ;
        RECT 589.950 589.950 592.050 592.050 ;
        RECT 593.400 589.050 594.450 592.950 ;
        RECT 595.950 589.950 598.050 595.050 ;
        RECT 592.950 586.950 595.050 589.050 ;
        RECT 602.400 588.450 603.450 599.400 ;
        RECT 607.950 598.950 610.050 601.050 ;
        RECT 599.400 587.400 603.450 588.450 ;
        RECT 586.950 580.950 589.050 583.050 ;
        RECT 569.400 571.350 570.600 572.100 ;
        RECT 575.400 571.350 576.600 572.100 ;
        RECT 565.950 568.950 568.050 571.050 ;
        RECT 568.950 568.950 571.050 571.050 ;
        RECT 571.950 568.950 574.050 571.050 ;
        RECT 574.950 568.950 577.050 571.050 ;
        RECT 566.400 566.400 567.600 568.650 ;
        RECT 572.400 566.400 573.600 568.650 ;
        RECT 566.400 556.050 567.450 566.400 ;
        RECT 572.400 564.450 573.450 566.400 ;
        RECT 572.400 563.400 576.450 564.450 ;
        RECT 571.950 556.950 574.050 559.050 ;
        RECT 565.950 553.950 568.050 556.050 ;
        RECT 572.400 553.050 573.450 556.950 ;
        RECT 575.400 556.050 576.450 563.400 ;
        RECT 581.400 562.050 582.450 572.100 ;
        RECT 583.950 571.950 586.050 574.050 ;
        RECT 586.950 572.100 589.050 574.200 ;
        RECT 592.950 573.000 595.050 577.050 ;
        RECT 599.400 574.050 600.450 587.400 ;
        RECT 608.400 586.050 609.450 598.950 ;
        RECT 615.150 593.700 616.350 612.300 ;
        RECT 620.400 606.450 621.600 606.600 ;
        RECT 623.400 606.450 624.450 616.950 ;
        RECT 629.400 606.450 630.450 662.400 ;
        RECT 635.400 651.450 636.450 682.950 ;
        RECT 644.400 682.350 645.600 684.600 ;
        RECT 652.950 683.100 655.050 685.200 ;
        RECT 658.950 683.100 661.050 685.200 ;
        RECT 664.950 683.100 667.050 685.200 ;
        RECT 668.400 685.050 669.450 691.950 ;
        RECT 643.950 679.950 646.050 682.050 ;
        RECT 646.950 679.950 649.050 682.050 ;
        RECT 647.400 677.400 648.600 679.650 ;
        RECT 647.400 673.050 648.450 677.400 ;
        RECT 653.400 673.050 654.450 683.100 ;
        RECT 659.400 682.350 660.600 683.100 ;
        RECT 665.400 682.350 666.600 683.100 ;
        RECT 667.950 682.950 670.050 685.050 ;
        RECT 658.950 679.950 661.050 682.050 ;
        RECT 661.950 679.950 664.050 682.050 ;
        RECT 664.950 679.950 667.050 682.050 ;
        RECT 662.400 678.900 663.600 679.650 ;
        RECT 661.950 676.800 664.050 678.900 ;
        RECT 664.950 673.950 667.050 676.050 ;
        RECT 646.950 670.950 649.050 673.050 ;
        RECT 652.950 670.950 655.050 673.050 ;
        RECT 655.950 667.950 658.050 670.050 ;
        RECT 643.050 657.300 645.150 659.400 ;
        RECT 632.400 650.400 636.450 651.450 ;
        RECT 632.400 622.050 633.450 650.400 ;
        RECT 637.800 646.950 639.900 649.050 ;
        RECT 638.400 645.900 639.600 646.650 ;
        RECT 637.950 643.800 640.050 645.900 ;
        RECT 643.650 638.700 644.850 657.300 ;
        RECT 646.950 646.950 649.050 649.050 ;
        RECT 647.400 645.000 648.600 646.650 ;
        RECT 646.950 640.950 649.050 645.000 ;
        RECT 640.650 637.500 644.850 638.700 ;
        RECT 640.650 636.600 642.750 637.500 ;
        RECT 656.400 637.050 657.450 667.950 ;
        RECT 665.400 651.600 666.450 673.950 ;
        RECT 671.400 670.050 672.450 697.950 ;
        RECT 674.400 670.050 675.450 706.950 ;
        RECT 676.950 694.950 679.050 697.050 ;
        RECT 677.400 691.050 678.450 694.950 ;
        RECT 686.400 694.050 687.450 722.400 ;
        RECT 694.950 718.950 697.050 723.000 ;
        RECT 700.800 721.950 702.900 724.050 ;
        RECT 703.950 721.950 706.050 724.050 ;
        RECT 713.400 722.400 714.600 724.650 ;
        RECT 722.400 722.400 723.600 724.650 ;
        RECT 701.400 718.050 702.450 721.950 ;
        RECT 713.400 718.050 714.450 722.400 ;
        RECT 700.950 715.950 703.050 718.050 ;
        RECT 712.950 715.950 715.050 718.050 ;
        RECT 722.400 712.050 723.450 722.400 ;
        RECT 726.150 716.700 727.350 735.300 ;
        RECT 731.100 724.950 733.200 727.050 ;
        RECT 731.400 723.900 732.600 724.650 ;
        RECT 730.950 721.800 733.050 723.900 ;
        RECT 726.150 715.500 730.350 716.700 ;
        RECT 728.250 714.600 730.350 715.500 ;
        RECT 694.950 709.950 697.050 712.050 ;
        RECT 721.950 709.950 724.050 712.050 ;
        RECT 685.950 691.950 688.050 694.050 ;
        RECT 676.950 688.950 679.050 691.050 ;
        RECT 688.950 688.950 691.050 691.050 ;
        RECT 682.950 684.000 685.050 688.050 ;
        RECT 689.400 684.600 690.450 688.950 ;
        RECT 683.400 682.350 684.600 684.000 ;
        RECT 689.400 682.350 690.600 684.600 ;
        RECT 679.950 679.950 682.050 682.050 ;
        RECT 682.950 679.950 685.050 682.050 ;
        RECT 685.950 679.950 688.050 682.050 ;
        RECT 688.950 679.950 691.050 682.050 ;
        RECT 676.950 676.950 679.050 679.050 ;
        RECT 680.400 678.900 681.600 679.650 ;
        RECT 686.400 678.900 687.600 679.650 ;
        RECT 670.800 667.950 672.900 670.050 ;
        RECT 673.950 667.950 676.050 670.050 ;
        RECT 677.400 666.450 678.450 676.950 ;
        RECT 679.950 676.800 682.050 678.900 ;
        RECT 685.950 676.800 688.050 678.900 ;
        RECT 691.950 676.950 694.050 679.050 ;
        RECT 685.950 672.450 688.050 673.050 ;
        RECT 692.400 672.450 693.450 676.950 ;
        RECT 685.950 671.400 693.450 672.450 ;
        RECT 685.950 670.950 688.050 671.400 ;
        RECT 688.950 667.950 691.050 670.050 ;
        RECT 674.400 665.400 678.450 666.450 ;
        RECT 674.400 661.050 675.450 665.400 ;
        RECT 673.950 658.950 676.050 661.050 ;
        RECT 677.850 657.300 679.950 659.400 ;
        RECT 665.400 649.350 666.600 651.600 ;
        RECT 661.950 646.950 664.050 649.050 ;
        RECT 664.950 646.950 667.050 649.050 ;
        RECT 667.950 646.950 670.050 649.050 ;
        RECT 673.950 646.950 676.050 649.050 ;
        RECT 662.400 644.400 663.600 646.650 ;
        RECT 668.400 644.400 669.600 646.650 ;
        RECT 674.400 645.900 675.600 646.650 ;
        RECT 662.400 640.050 663.450 644.400 ;
        RECT 661.950 637.950 664.050 640.050 ;
        RECT 655.950 634.950 658.050 637.050 ;
        RECT 668.400 634.050 669.450 644.400 ;
        RECT 673.950 640.950 676.050 645.900 ;
        RECT 678.150 638.700 679.350 657.300 ;
        RECT 683.100 646.950 685.200 649.050 ;
        RECT 683.400 645.450 684.600 646.650 ;
        RECT 683.400 644.400 687.450 645.450 ;
        RECT 678.150 637.500 682.350 638.700 ;
        RECT 680.250 636.600 682.350 637.500 ;
        RECT 667.950 631.950 670.050 634.050 ;
        RECT 631.950 619.950 634.050 622.050 ;
        RECT 646.950 619.950 649.050 622.050 ;
        RECT 620.400 605.400 624.450 606.450 ;
        RECT 626.400 605.400 630.450 606.450 ;
        RECT 632.550 615.300 634.650 617.400 ;
        RECT 632.550 608.700 633.750 615.300 ;
        RECT 643.950 610.950 646.050 613.050 ;
        RECT 632.550 606.600 634.650 608.700 ;
        RECT 620.400 604.350 621.600 605.400 ;
        RECT 620.100 601.950 622.200 604.050 ;
        RECT 614.850 591.600 616.950 593.700 ;
        RECT 626.400 592.050 627.450 605.400 ;
        RECT 628.950 601.950 631.050 604.050 ;
        RECT 619.950 589.950 622.050 592.050 ;
        RECT 625.950 589.950 628.050 592.050 ;
        RECT 601.950 583.950 604.050 586.050 ;
        RECT 607.950 583.950 610.050 586.050 ;
        RECT 587.400 571.350 588.600 572.100 ;
        RECT 593.400 571.350 594.600 573.000 ;
        RECT 598.950 571.950 601.050 574.050 ;
        RECT 602.400 573.600 603.450 583.950 ;
        RECT 607.350 579.300 609.450 581.400 ;
        RECT 602.400 571.350 603.600 573.600 ;
        RECT 586.950 568.950 589.050 571.050 ;
        RECT 589.950 568.950 592.050 571.050 ;
        RECT 592.950 568.950 595.050 571.050 ;
        RECT 595.950 568.950 598.050 571.050 ;
        RECT 601.950 568.950 604.050 571.050 ;
        RECT 583.950 565.950 586.050 568.050 ;
        RECT 590.400 566.400 591.600 568.650 ;
        RECT 596.400 567.900 597.600 568.650 ;
        RECT 580.950 559.950 583.050 562.050 ;
        RECT 574.950 553.950 577.050 556.050 ;
        RECT 571.950 550.950 574.050 553.050 ;
        RECT 559.950 535.950 562.050 538.050 ;
        RECT 535.950 532.950 538.050 535.050 ;
        RECT 547.950 532.950 550.050 535.050 ;
        RECT 556.950 532.950 559.050 535.050 ;
        RECT 565.950 532.950 568.050 535.050 ;
        RECT 523.950 529.950 526.050 532.050 ;
        RECT 532.950 529.950 535.050 532.050 ;
        RECT 518.400 526.350 519.600 528.600 ;
        RECT 517.950 523.950 520.050 526.050 ;
        RECT 514.050 513.600 516.150 515.700 ;
        RECT 524.400 502.050 525.450 529.950 ;
        RECT 536.400 528.600 537.450 532.950 ;
        RECT 536.400 526.350 537.600 528.600 ;
        RECT 541.950 527.100 544.050 529.200 ;
        RECT 542.400 526.350 543.600 527.100 ;
        RECT 532.950 523.950 535.050 526.050 ;
        RECT 535.950 523.950 538.050 526.050 ;
        RECT 538.950 523.950 541.050 526.050 ;
        RECT 541.950 523.950 544.050 526.050 ;
        RECT 533.400 522.900 534.600 523.650 ;
        RECT 532.950 520.800 535.050 522.900 ;
        RECT 539.400 521.400 540.600 523.650 ;
        RECT 532.950 511.950 535.050 514.050 ;
        RECT 523.950 499.950 526.050 502.050 ;
        RECT 502.950 496.950 505.050 499.050 ;
        RECT 508.950 496.950 511.050 499.050 ;
        RECT 494.400 493.350 495.600 495.600 ;
        RECT 499.950 494.100 502.050 496.200 ;
        RECT 500.400 493.350 501.600 494.100 ;
        RECT 493.950 490.950 496.050 493.050 ;
        RECT 496.950 490.950 499.050 493.050 ;
        RECT 499.950 490.950 502.050 493.050 ;
        RECT 502.950 490.950 505.050 493.050 ;
        RECT 479.400 488.400 486.450 489.450 ;
        RECT 497.400 489.000 498.600 490.650 ;
        RECT 503.400 489.900 504.600 490.650 ;
        RECT 484.950 484.950 487.050 487.050 ;
        RECT 496.950 484.950 499.050 489.000 ;
        RECT 502.950 487.800 505.050 489.900 ;
        RECT 472.650 481.500 476.850 482.700 ;
        RECT 472.650 480.600 474.750 481.500 ;
        RECT 460.950 461.400 465.450 462.450 ;
        RECT 460.950 460.950 463.050 461.400 ;
        RECT 439.950 449.100 442.050 451.200 ;
        RECT 440.400 448.350 441.600 449.100 ;
        RECT 448.950 448.950 451.050 451.050 ;
        RECT 454.950 449.100 457.050 451.200 ;
        RECT 461.400 450.600 462.450 460.950 ;
        RECT 485.400 454.050 486.450 484.950 ;
        RECT 493.950 478.950 496.050 481.050 ;
        RECT 439.950 445.950 442.050 448.050 ;
        RECT 442.950 445.950 445.050 448.050 ;
        RECT 433.950 442.800 436.050 444.900 ;
        RECT 443.400 443.400 444.600 445.650 ;
        RECT 376.050 435.600 378.150 437.700 ;
        RECT 403.950 436.950 406.050 439.050 ;
        RECT 412.950 436.950 415.050 439.050 ;
        RECT 430.950 436.950 433.050 439.050 ;
        RECT 370.950 427.950 373.050 430.050 ;
        RECT 371.400 418.200 372.450 427.950 ;
        RECT 379.050 423.300 381.150 425.400 ;
        RECT 370.950 416.100 373.050 418.200 ;
        RECT 373.800 412.950 375.900 415.050 ;
        RECT 374.400 411.900 375.600 412.650 ;
        RECT 373.950 409.800 376.050 411.900 ;
        RECT 340.950 403.950 343.050 406.050 ;
        RECT 349.950 403.950 352.050 406.050 ;
        RECT 328.950 400.950 331.050 403.050 ;
        RECT 362.250 401.700 363.450 408.300 ;
        RECT 364.950 406.950 367.050 409.050 ;
        RECT 367.950 406.950 370.050 409.050 ;
        RECT 361.350 399.600 363.450 401.700 ;
        RECT 368.400 400.050 369.450 406.950 ;
        RECT 379.650 404.700 380.850 423.300 ;
        RECT 388.950 418.950 391.050 421.050 ;
        RECT 394.950 420.450 397.050 421.050 ;
        RECT 394.950 419.400 405.450 420.450 ;
        RECT 394.950 418.950 397.050 419.400 ;
        RECT 389.400 415.050 390.450 418.950 ;
        RECT 391.950 415.950 394.050 418.050 ;
        RECT 397.950 416.100 400.050 418.200 ;
        RECT 404.400 417.600 405.450 419.400 ;
        RECT 382.950 412.950 385.050 415.050 ;
        RECT 388.950 412.950 391.050 415.050 ;
        RECT 383.400 411.000 384.600 412.650 ;
        RECT 382.950 406.950 385.050 411.000 ;
        RECT 392.400 409.050 393.450 415.950 ;
        RECT 398.400 415.350 399.600 416.100 ;
        RECT 404.400 415.350 405.600 417.600 ;
        RECT 397.950 412.950 400.050 415.050 ;
        RECT 400.950 412.950 403.050 415.050 ;
        RECT 403.950 412.950 406.050 415.050 ;
        RECT 406.950 412.950 409.050 415.050 ;
        RECT 401.400 410.400 402.600 412.650 ;
        RECT 407.400 411.900 408.600 412.650 ;
        RECT 391.950 406.950 394.050 409.050 ;
        RECT 376.650 403.500 380.850 404.700 ;
        RECT 376.650 402.600 378.750 403.500 ;
        RECT 367.950 397.950 370.050 400.050 ;
        RECT 349.950 391.950 352.050 394.050 ;
        RECT 346.350 381.300 348.450 383.400 ;
        RECT 313.950 376.950 316.050 379.050 ;
        RECT 314.400 372.600 315.450 376.950 ;
        RECT 347.250 374.700 348.450 381.300 ;
        RECT 314.400 370.350 315.600 372.600 ;
        RECT 319.950 371.100 322.050 373.200 ;
        RECT 325.950 371.100 328.050 373.200 ;
        RECT 334.950 371.100 337.050 373.200 ;
        RECT 346.350 372.600 348.450 374.700 ;
        RECT 320.400 370.350 321.600 371.100 ;
        RECT 310.950 367.950 313.050 370.050 ;
        RECT 313.950 367.950 316.050 370.050 ;
        RECT 316.950 367.950 319.050 370.050 ;
        RECT 319.950 367.950 322.050 370.050 ;
        RECT 305.400 365.400 309.450 366.450 ;
        RECT 290.550 357.600 292.650 359.700 ;
        RECT 287.400 344.400 291.450 345.450 ;
        RECT 281.400 339.600 282.450 343.950 ;
        RECT 281.400 337.350 282.600 339.600 ;
        RECT 280.950 334.950 283.050 337.050 ;
        RECT 283.950 334.950 286.050 337.050 ;
        RECT 284.400 332.400 285.600 334.650 ;
        RECT 274.950 328.950 277.050 331.050 ;
        RECT 265.950 316.950 268.050 319.050 ;
        RECT 274.950 313.950 277.050 316.050 ;
        RECT 262.950 307.950 265.050 310.050 ;
        RECT 259.950 295.950 262.050 298.050 ;
        RECT 263.400 295.050 264.450 307.950 ;
        RECT 275.400 307.050 276.450 313.950 ;
        RECT 274.950 304.950 277.050 307.050 ;
        RECT 284.400 304.050 285.450 332.400 ;
        RECT 286.950 328.950 289.050 331.050 ;
        RECT 283.950 301.950 286.050 304.050 ;
        RECT 261.000 294.600 265.050 295.050 ;
        RECT 248.400 292.350 249.600 293.100 ;
        RECT 254.400 292.350 255.600 294.600 ;
        RECT 260.400 292.950 265.050 294.600 ;
        RECT 274.950 293.100 277.050 295.200 ;
        RECT 280.950 293.100 283.050 298.050 ;
        RECT 284.400 295.050 285.450 301.950 ;
        RECT 287.400 298.050 288.450 328.950 ;
        RECT 290.400 325.050 291.450 344.400 ;
        RECT 298.950 338.100 301.050 340.200 ;
        RECT 299.400 337.350 300.600 338.100 ;
        RECT 295.950 334.950 298.050 337.050 ;
        RECT 298.950 334.950 301.050 337.050 ;
        RECT 301.950 334.950 304.050 337.050 ;
        RECT 296.400 332.400 297.600 334.650 ;
        RECT 302.400 333.450 303.600 334.650 ;
        RECT 302.400 332.400 306.450 333.450 ;
        RECT 296.400 325.050 297.450 332.400 ;
        RECT 298.950 328.950 301.050 331.050 ;
        RECT 301.950 328.950 304.050 331.050 ;
        RECT 289.950 322.950 292.050 325.050 ;
        RECT 295.950 322.950 298.050 325.050 ;
        RECT 296.400 301.050 297.450 322.950 ;
        RECT 295.950 298.950 298.050 301.050 ;
        RECT 286.950 295.950 289.050 298.050 ;
        RECT 260.400 292.350 261.600 292.950 ;
        RECT 275.400 292.350 276.600 293.100 ;
        RECT 229.950 289.950 232.050 292.050 ;
        RECT 232.950 289.950 235.050 292.050 ;
        RECT 235.950 289.950 238.050 292.050 ;
        RECT 247.950 289.950 250.050 292.050 ;
        RECT 250.950 289.950 253.050 292.050 ;
        RECT 253.950 289.950 256.050 292.050 ;
        RECT 256.950 289.950 259.050 292.050 ;
        RECT 259.950 289.950 262.050 292.050 ;
        RECT 271.950 289.950 274.050 292.050 ;
        RECT 274.950 289.950 277.050 292.050 ;
        RECT 233.400 287.400 234.600 289.650 ;
        RECT 233.400 277.050 234.450 287.400 ;
        RECT 238.950 286.950 241.050 289.050 ;
        RECT 244.950 286.950 247.050 289.050 ;
        RECT 251.400 288.900 252.600 289.650 ;
        RECT 257.400 288.900 258.600 289.650 ;
        RECT 272.400 288.900 273.600 289.650 ;
        RECT 239.400 277.050 240.450 286.950 ;
        RECT 232.950 274.950 235.050 277.050 ;
        RECT 238.950 274.950 241.050 277.050 ;
        RECT 223.950 271.950 226.050 274.050 ;
        RECT 245.400 271.050 246.450 286.950 ;
        RECT 250.950 286.800 253.050 288.900 ;
        RECT 256.950 286.800 259.050 288.900 ;
        RECT 262.950 286.800 265.050 288.900 ;
        RECT 271.950 286.800 274.050 288.900 ;
        RECT 251.400 283.050 252.450 286.800 ;
        RECT 263.400 283.050 264.450 286.800 ;
        RECT 281.400 286.050 282.450 293.100 ;
        RECT 283.950 292.950 286.050 295.050 ;
        RECT 289.950 294.000 292.050 298.050 ;
        RECT 296.400 294.450 297.600 294.600 ;
        RECT 299.400 294.450 300.450 328.950 ;
        RECT 290.400 292.350 291.600 294.000 ;
        RECT 296.400 293.400 300.450 294.450 ;
        RECT 296.400 292.350 297.600 293.400 ;
        RECT 286.950 289.950 289.050 292.050 ;
        RECT 289.950 289.950 292.050 292.050 ;
        RECT 292.950 289.950 295.050 292.050 ;
        RECT 295.950 289.950 298.050 292.050 ;
        RECT 287.400 289.050 288.600 289.650 ;
        RECT 283.950 287.400 288.600 289.050 ;
        RECT 293.400 287.400 294.600 289.650 ;
        RECT 283.950 286.950 288.000 287.400 ;
        RECT 271.950 283.650 274.050 285.750 ;
        RECT 274.950 283.950 277.050 286.050 ;
        RECT 280.950 283.950 283.050 286.050 ;
        RECT 250.950 280.950 253.050 283.050 ;
        RECT 262.950 280.950 265.050 283.050 ;
        RECT 247.950 274.950 250.050 277.050 ;
        RECT 244.950 268.950 247.050 271.050 ;
        RECT 214.950 259.950 217.050 262.050 ;
        RECT 220.950 261.000 223.050 265.050 ;
        RECT 221.400 259.350 222.600 261.000 ;
        RECT 238.950 260.100 241.050 262.200 ;
        RECT 239.400 259.350 240.600 260.100 ;
        RECT 217.950 256.950 220.050 259.050 ;
        RECT 220.950 256.950 223.050 259.050 ;
        RECT 223.950 256.950 226.050 259.050 ;
        RECT 236.100 256.950 238.200 259.050 ;
        RECT 239.400 256.950 241.500 259.050 ;
        RECT 244.800 256.950 246.900 259.050 ;
        RECT 218.400 254.400 219.600 256.650 ;
        RECT 224.400 255.900 225.600 256.650 ;
        RECT 236.400 255.900 237.600 256.650 ;
        RECT 199.950 244.950 202.050 247.050 ;
        RECT 211.950 244.950 214.050 247.050 ;
        RECT 190.950 226.950 193.050 229.050 ;
        RECT 184.950 215.100 187.050 217.200 ;
        RECT 191.400 216.600 192.450 226.950 ;
        RECT 196.950 220.950 199.050 223.050 ;
        RECT 185.400 214.350 186.600 215.100 ;
        RECT 191.400 214.350 192.600 216.600 ;
        RECT 184.950 211.950 187.050 214.050 ;
        RECT 187.950 211.950 190.050 214.050 ;
        RECT 190.950 211.950 193.050 214.050 ;
        RECT 181.950 208.950 184.050 211.050 ;
        RECT 188.400 209.400 189.600 211.650 ;
        RECT 178.950 205.950 181.050 208.050 ;
        RECT 160.950 202.950 163.050 205.050 ;
        RECT 154.950 193.950 157.050 196.050 ;
        RECT 143.400 182.400 147.450 183.450 ;
        RECT 154.950 183.000 157.050 187.050 ;
        RECT 160.950 184.950 163.050 187.050 ;
        RECT 136.950 178.950 139.050 181.050 ;
        RECT 139.950 178.950 142.050 181.050 ;
        RECT 137.400 177.900 138.600 178.650 ;
        RECT 136.950 175.800 139.050 177.900 ;
        RECT 130.950 172.950 133.050 175.050 ;
        RECT 94.950 148.950 97.050 151.050 ;
        RECT 109.950 148.950 112.050 151.050 ;
        RECT 76.950 142.950 79.050 145.050 ;
        RECT 82.950 142.950 85.050 145.050 ;
        RECT 88.950 142.950 91.050 145.050 ;
        RECT 77.400 138.600 78.450 142.950 ;
        RECT 83.400 139.200 84.450 142.950 ;
        RECT 95.400 142.050 96.450 148.950 ;
        RECT 146.400 148.050 147.450 182.400 ;
        RECT 155.400 181.350 156.600 183.000 ;
        RECT 151.950 178.950 154.050 181.050 ;
        RECT 154.950 178.950 157.050 181.050 ;
        RECT 152.400 176.400 153.600 178.650 ;
        RECT 145.950 145.950 148.050 148.050 ;
        RECT 103.950 142.950 106.050 145.050 ;
        RECT 130.950 142.950 133.050 145.050 ;
        RECT 88.950 139.800 91.050 141.900 ;
        RECT 94.950 139.950 97.050 142.050 ;
        RECT 77.400 136.350 78.600 138.600 ;
        RECT 82.950 137.100 85.050 139.200 ;
        RECT 83.400 136.350 84.600 137.100 ;
        RECT 73.950 133.950 76.050 136.050 ;
        RECT 76.950 133.950 79.050 136.050 ;
        RECT 79.950 133.950 82.050 136.050 ;
        RECT 82.950 133.950 85.050 136.050 ;
        RECT 74.400 131.400 75.600 133.650 ;
        RECT 80.400 132.900 81.600 133.650 ;
        RECT 55.950 127.950 58.050 130.050 ;
        RECT 61.950 127.950 64.050 130.050 ;
        RECT 67.950 127.950 70.050 130.050 ;
        RECT 52.950 112.950 55.050 115.050 ;
        RECT 50.400 111.000 54.450 111.450 ;
        RECT 50.400 110.400 55.050 111.000 ;
        RECT 46.950 106.950 49.050 109.050 ;
        RECT 52.950 106.950 55.050 110.400 ;
        RECT 49.950 104.100 52.050 106.200 ;
        RECT 56.400 105.600 57.450 127.950 ;
        RECT 58.950 112.950 61.050 115.050 ;
        RECT 59.400 106.050 60.450 112.950 ;
        RECT 50.400 103.350 51.600 104.100 ;
        RECT 56.400 103.350 57.600 105.600 ;
        RECT 58.950 103.950 61.050 106.050 ;
        RECT 46.950 100.950 49.050 103.050 ;
        RECT 49.950 100.950 52.050 103.050 ;
        RECT 52.950 100.950 55.050 103.050 ;
        RECT 55.950 100.950 58.050 103.050 ;
        RECT 47.400 99.450 48.600 100.650 ;
        RECT 41.400 98.400 48.600 99.450 ;
        RECT 53.400 99.000 54.600 100.650 ;
        RECT 23.400 77.400 27.450 78.450 ;
        RECT 22.950 70.950 25.050 73.050 ;
        RECT 16.950 59.100 19.050 61.200 ;
        RECT 23.400 60.600 24.450 70.950 ;
        RECT 26.400 61.050 27.450 77.400 ;
        RECT 38.400 76.050 39.450 97.950 ;
        RECT 52.950 94.950 55.050 99.000 ;
        RECT 62.400 85.050 63.450 127.950 ;
        RECT 74.400 121.050 75.450 131.400 ;
        RECT 79.950 130.800 82.050 132.900 ;
        RECT 89.400 130.050 90.450 139.800 ;
        RECT 104.400 139.200 105.450 142.950 ;
        RECT 97.950 137.100 100.050 139.200 ;
        RECT 103.950 137.100 106.050 139.200 ;
        RECT 109.950 137.100 112.050 139.200 ;
        RECT 118.950 137.100 121.050 139.200 ;
        RECT 124.950 137.100 127.050 139.200 ;
        RECT 98.400 136.350 99.600 137.100 ;
        RECT 104.400 136.350 105.600 137.100 ;
        RECT 94.950 133.950 97.050 136.050 ;
        RECT 97.950 133.950 100.050 136.050 ;
        RECT 100.950 133.950 103.050 136.050 ;
        RECT 103.950 133.950 106.050 136.050 ;
        RECT 95.400 131.400 96.600 133.650 ;
        RECT 101.400 132.900 102.600 133.650 ;
        RECT 82.950 127.950 85.050 130.050 ;
        RECT 88.950 127.950 91.050 130.050 ;
        RECT 73.950 118.950 76.050 121.050 ;
        RECT 67.950 105.000 70.050 109.050 ;
        RECT 73.950 105.000 76.050 109.050 ;
        RECT 68.400 103.350 69.600 105.000 ;
        RECT 74.400 103.350 75.600 105.000 ;
        RECT 67.950 100.950 70.050 103.050 ;
        RECT 70.950 100.950 73.050 103.050 ;
        RECT 73.950 100.950 76.050 103.050 ;
        RECT 76.950 100.950 79.050 103.050 ;
        RECT 71.400 99.000 72.600 100.650 ;
        RECT 70.950 94.950 73.050 99.000 ;
        RECT 77.400 98.400 78.600 100.650 ;
        RECT 77.400 94.050 78.450 98.400 ;
        RECT 79.950 97.950 82.050 100.050 ;
        RECT 76.950 91.950 79.050 94.050 ;
        RECT 61.950 82.950 64.050 85.050 ;
        RECT 37.950 73.950 40.050 76.050 ;
        RECT 61.950 73.950 64.050 76.050 ;
        RECT 76.950 73.950 79.050 76.050 ;
        RECT 28.950 70.950 31.050 73.050 ;
        RECT 17.400 58.350 18.600 59.100 ;
        RECT 23.400 58.350 24.600 60.600 ;
        RECT 25.950 58.950 28.050 61.050 ;
        RECT 13.950 55.950 16.050 58.050 ;
        RECT 16.950 55.950 19.050 58.050 ;
        RECT 19.950 55.950 22.050 58.050 ;
        RECT 22.950 55.950 25.050 58.050 ;
        RECT 4.950 52.950 7.050 55.050 ;
        RECT 14.400 54.900 15.600 55.650 ;
        RECT 13.950 52.800 16.050 54.900 ;
        RECT 20.400 53.400 21.600 55.650 ;
        RECT 16.950 49.950 19.050 52.050 ;
        RECT 17.400 46.050 18.450 49.950 ;
        RECT 16.950 43.950 19.050 46.050 ;
        RECT 20.400 40.050 21.450 53.400 ;
        RECT 13.950 37.950 16.050 40.050 ;
        RECT 19.950 37.950 22.050 40.050 ;
        RECT 14.400 27.600 15.450 37.950 ;
        RECT 29.400 27.600 30.450 70.950 ;
        RECT 31.950 64.950 34.050 67.050 ;
        RECT 49.950 64.950 52.050 67.050 ;
        RECT 32.400 61.050 33.450 64.950 ;
        RECT 31.950 58.950 34.050 61.050 ;
        RECT 37.950 60.000 40.050 64.050 ;
        RECT 38.400 58.350 39.600 60.000 ;
        RECT 43.950 59.100 46.050 61.200 ;
        RECT 44.400 58.350 45.600 59.100 ;
        RECT 34.950 55.950 37.050 58.050 ;
        RECT 37.950 55.950 40.050 58.050 ;
        RECT 40.950 55.950 43.050 58.050 ;
        RECT 43.950 55.950 46.050 58.050 ;
        RECT 31.950 52.950 34.050 55.050 ;
        RECT 35.400 54.900 36.600 55.650 ;
        RECT 32.400 49.050 33.450 52.950 ;
        RECT 34.950 52.800 37.050 54.900 ;
        RECT 41.400 53.400 42.600 55.650 ;
        RECT 50.400 55.050 51.450 64.950 ;
        RECT 52.950 61.950 55.050 64.050 ;
        RECT 37.950 49.950 40.050 52.050 ;
        RECT 31.950 46.950 34.050 49.050 ;
        RECT 14.400 25.350 15.600 27.600 ;
        RECT 29.400 25.350 30.600 27.600 ;
        RECT 13.950 22.950 16.050 25.050 ;
        RECT 16.950 22.950 19.050 25.050 ;
        RECT 28.950 22.950 31.050 25.050 ;
        RECT 31.950 22.950 34.050 25.050 ;
        RECT 17.400 20.400 18.600 22.650 ;
        RECT 32.400 21.900 33.600 22.650 ;
        RECT 38.400 22.050 39.450 49.950 ;
        RECT 41.400 49.050 42.450 53.400 ;
        RECT 49.950 52.950 52.050 55.050 ;
        RECT 46.950 49.950 49.050 52.050 ;
        RECT 40.950 46.950 43.050 49.050 ;
        RECT 47.400 46.050 48.450 49.950 ;
        RECT 53.400 49.050 54.450 61.950 ;
        RECT 62.400 60.600 63.450 73.950 ;
        RECT 62.400 58.350 63.600 60.600 ;
        RECT 67.950 59.100 70.050 61.200 ;
        RECT 73.950 59.100 76.050 61.200 ;
        RECT 77.400 60.450 78.450 73.950 ;
        RECT 80.400 64.050 81.450 97.950 ;
        RECT 83.400 97.050 84.450 127.950 ;
        RECT 88.950 121.950 91.050 124.050 ;
        RECT 89.400 105.600 90.450 121.950 ;
        RECT 95.400 115.050 96.450 131.400 ;
        RECT 100.950 130.800 103.050 132.900 ;
        RECT 101.400 127.050 102.450 130.800 ;
        RECT 100.950 124.950 103.050 127.050 ;
        RECT 103.950 121.950 106.050 124.050 ;
        RECT 94.950 112.950 97.050 115.050 ;
        RECT 104.400 109.050 105.450 121.950 ;
        RECT 110.400 121.050 111.450 137.100 ;
        RECT 119.400 136.350 120.600 137.100 ;
        RECT 125.400 136.350 126.600 137.100 ;
        RECT 115.950 133.950 118.050 136.050 ;
        RECT 118.950 133.950 121.050 136.050 ;
        RECT 121.950 133.950 124.050 136.050 ;
        RECT 124.950 133.950 127.050 136.050 ;
        RECT 112.950 130.950 115.050 133.050 ;
        RECT 116.400 131.400 117.600 133.650 ;
        RECT 122.400 131.400 123.600 133.650 ;
        RECT 109.950 118.950 112.050 121.050 ;
        RECT 113.400 112.050 114.450 130.950 ;
        RECT 116.400 129.450 117.450 131.400 ;
        RECT 116.400 128.400 120.450 129.450 ;
        RECT 112.950 109.950 115.050 112.050 ;
        RECT 89.400 103.350 90.600 105.600 ;
        RECT 94.950 104.100 97.050 106.200 ;
        RECT 100.950 104.100 103.050 109.050 ;
        RECT 103.950 106.950 106.050 109.050 ;
        RECT 95.400 103.350 96.600 104.100 ;
        RECT 88.950 100.950 91.050 103.050 ;
        RECT 91.950 100.950 94.050 103.050 ;
        RECT 94.950 100.950 97.050 103.050 ;
        RECT 97.950 100.950 100.050 103.050 ;
        RECT 92.400 99.000 93.600 100.650 ;
        RECT 98.400 99.900 99.600 100.650 ;
        RECT 82.950 94.950 85.050 97.050 ;
        RECT 91.950 94.950 94.050 99.000 ;
        RECT 97.950 97.800 100.050 99.900 ;
        RECT 100.950 97.950 103.050 100.050 ;
        RECT 104.400 99.900 105.450 106.950 ;
        RECT 106.950 103.950 109.050 109.050 ;
        RECT 119.400 106.200 120.450 128.400 ;
        RECT 122.400 121.050 123.450 131.400 ;
        RECT 127.950 121.950 130.050 124.050 ;
        RECT 121.950 118.950 124.050 121.050 ;
        RECT 124.950 112.950 127.050 115.050 ;
        RECT 121.950 109.950 124.050 112.050 ;
        RECT 112.950 104.100 115.050 106.200 ;
        RECT 118.950 104.100 121.050 106.200 ;
        RECT 122.400 106.050 123.450 109.950 ;
        RECT 113.400 103.350 114.600 104.100 ;
        RECT 119.400 103.350 120.600 104.100 ;
        RECT 121.950 103.950 124.050 106.050 ;
        RECT 109.950 100.950 112.050 103.050 ;
        RECT 112.950 100.950 115.050 103.050 ;
        RECT 115.950 100.950 118.050 103.050 ;
        RECT 118.950 100.950 121.050 103.050 ;
        RECT 101.400 94.050 102.450 97.950 ;
        RECT 103.950 97.800 106.050 99.900 ;
        RECT 110.400 99.000 111.600 100.650 ;
        RECT 109.950 94.950 112.050 99.000 ;
        RECT 116.400 98.400 117.600 100.650 ;
        RECT 100.950 91.950 103.050 94.050 ;
        RECT 116.400 91.050 117.450 98.400 ;
        RECT 121.950 97.950 124.050 100.050 ;
        RECT 122.400 91.050 123.450 97.950 ;
        RECT 125.400 97.050 126.450 112.950 ;
        RECT 128.400 112.050 129.450 121.950 ;
        RECT 131.400 115.050 132.450 142.950 ;
        RECT 145.950 142.800 148.050 144.900 ;
        RECT 139.950 137.100 142.050 139.200 ;
        RECT 146.400 138.600 147.450 142.800 ;
        RECT 140.400 136.350 141.600 137.100 ;
        RECT 146.400 136.350 147.600 138.600 ;
        RECT 136.950 133.950 139.050 136.050 ;
        RECT 139.950 133.950 142.050 136.050 ;
        RECT 142.950 133.950 145.050 136.050 ;
        RECT 145.950 133.950 148.050 136.050 ;
        RECT 133.950 130.950 136.050 133.050 ;
        RECT 137.400 131.400 138.600 133.650 ;
        RECT 143.400 132.900 144.600 133.650 ;
        RECT 152.400 132.900 153.450 176.400 ;
        RECT 161.400 172.050 162.450 184.950 ;
        RECT 160.950 169.950 163.050 172.050 ;
        RECT 154.950 145.950 157.050 148.050 ;
        RECT 134.400 121.050 135.450 130.950 ;
        RECT 137.400 127.050 138.450 131.400 ;
        RECT 142.950 130.800 145.050 132.900 ;
        RECT 151.950 130.800 154.050 132.900 ;
        RECT 136.950 124.950 139.050 127.050 ;
        RECT 133.950 118.950 136.050 121.050 ;
        RECT 130.950 112.950 133.050 115.050 ;
        RECT 127.950 109.950 130.050 112.050 ;
        RECT 134.400 105.600 135.450 118.950 ;
        RECT 145.950 115.950 148.050 118.050 ;
        RECT 146.400 105.600 147.450 115.950 ;
        RECT 134.400 103.350 135.600 105.600 ;
        RECT 146.400 103.350 147.600 105.600 ;
        RECT 151.950 105.000 154.050 109.050 ;
        RECT 155.400 106.050 156.450 145.950 ;
        RECT 164.400 142.200 165.450 205.950 ;
        RECT 179.400 196.050 180.450 205.950 ;
        RECT 178.950 193.950 181.050 196.050 ;
        RECT 182.400 193.050 183.450 208.950 ;
        RECT 188.400 205.050 189.450 209.400 ;
        RECT 187.950 202.950 190.050 205.050 ;
        RECT 181.950 190.950 184.050 193.050 ;
        RECT 178.950 184.950 181.050 187.050 ;
        RECT 172.950 182.100 175.050 184.200 ;
        RECT 173.400 181.350 174.600 182.100 ;
        RECT 167.100 178.950 169.200 181.050 ;
        RECT 172.500 178.950 174.600 181.050 ;
        RECT 175.800 178.950 177.900 181.050 ;
        RECT 167.400 177.900 168.600 178.650 ;
        RECT 166.950 175.800 169.050 177.900 ;
        RECT 176.400 176.400 177.600 178.650 ;
        RECT 176.400 148.050 177.450 176.400 ;
        RECT 179.400 166.050 180.450 184.950 ;
        RECT 178.950 163.950 181.050 166.050 ;
        RECT 182.400 148.050 183.450 190.950 ;
        RECT 188.400 187.050 189.450 202.950 ;
        RECT 197.400 202.050 198.450 220.950 ;
        RECT 200.400 208.050 201.450 244.950 ;
        RECT 205.950 229.950 208.050 232.050 ;
        RECT 206.400 217.050 207.450 229.950 ;
        RECT 218.400 226.050 219.450 254.400 ;
        RECT 223.950 253.800 226.050 255.900 ;
        RECT 235.950 253.800 238.050 255.900 ;
        RECT 245.400 255.450 246.600 256.650 ;
        RECT 248.400 255.450 249.450 274.950 ;
        RECT 253.950 262.950 256.050 265.050 ;
        RECT 250.950 260.100 253.050 262.200 ;
        RECT 245.400 254.400 249.450 255.450 ;
        RECT 229.950 250.950 232.050 253.050 ;
        RECT 230.400 232.050 231.450 250.950 ;
        RECT 235.950 241.950 238.050 244.050 ;
        RECT 229.950 229.950 232.050 232.050 ;
        RECT 217.950 223.950 220.050 226.050 ;
        RECT 211.950 220.950 214.050 223.050 ;
        RECT 232.950 220.950 235.050 223.050 ;
        RECT 202.950 216.600 207.450 217.050 ;
        RECT 212.400 216.600 213.450 220.950 ;
        RECT 233.400 216.600 234.450 220.950 ;
        RECT 236.400 217.050 237.450 241.950 ;
        RECT 238.950 235.950 241.050 238.050 ;
        RECT 202.950 214.950 207.600 216.600 ;
        RECT 206.400 214.350 207.600 214.950 ;
        RECT 212.400 214.350 213.600 216.600 ;
        RECT 233.400 214.350 234.600 216.600 ;
        RECT 235.950 214.950 238.050 217.050 ;
        RECT 205.950 211.950 208.050 214.050 ;
        RECT 208.950 211.950 211.050 214.050 ;
        RECT 211.950 211.950 214.050 214.050 ;
        RECT 226.950 211.950 229.050 214.050 ;
        RECT 229.950 211.950 232.050 214.050 ;
        RECT 232.950 211.950 235.050 214.050 ;
        RECT 202.950 208.950 205.050 211.050 ;
        RECT 209.400 210.900 210.600 211.650 ;
        RECT 230.400 210.900 231.600 211.650 ;
        RECT 199.950 205.950 202.050 208.050 ;
        RECT 190.950 199.950 193.050 202.050 ;
        RECT 196.950 199.950 199.050 202.050 ;
        RECT 187.950 184.950 190.050 187.050 ;
        RECT 191.400 184.200 192.450 199.950 ;
        RECT 190.950 182.100 193.050 184.200 ;
        RECT 196.950 183.000 199.050 187.050 ;
        RECT 203.400 184.050 204.450 208.950 ;
        RECT 208.950 208.800 211.050 210.900 ;
        RECT 229.950 208.800 232.050 210.900 ;
        RECT 205.950 205.950 208.050 208.050 ;
        RECT 191.400 181.350 192.600 182.100 ;
        RECT 197.400 181.350 198.600 183.000 ;
        RECT 202.950 181.950 205.050 184.050 ;
        RECT 187.950 178.950 190.050 181.050 ;
        RECT 190.950 178.950 193.050 181.050 ;
        RECT 193.950 178.950 196.050 181.050 ;
        RECT 196.950 178.950 199.050 181.050 ;
        RECT 199.950 178.950 202.050 181.050 ;
        RECT 188.400 177.900 189.600 178.650 ;
        RECT 187.950 175.800 190.050 177.900 ;
        RECT 194.400 176.400 195.600 178.650 ;
        RECT 200.400 177.900 201.600 178.650 ;
        RECT 199.950 177.450 202.050 177.900 ;
        RECT 199.950 176.400 204.450 177.450 ;
        RECT 188.400 148.050 189.450 175.800 ;
        RECT 194.400 169.050 195.450 176.400 ;
        RECT 199.950 175.800 202.050 176.400 ;
        RECT 196.950 169.950 199.050 172.050 ;
        RECT 193.950 166.950 196.050 169.050 ;
        RECT 190.950 148.950 193.050 151.050 ;
        RECT 175.950 145.950 178.050 148.050 ;
        RECT 181.950 145.950 184.050 148.050 ;
        RECT 187.950 145.950 190.050 148.050 ;
        RECT 163.950 140.100 166.050 142.200 ;
        RECT 175.950 139.950 178.050 142.050 ;
        RECT 163.950 136.950 166.050 139.050 ;
        RECT 169.950 137.100 172.050 139.200 ;
        RECT 164.400 136.350 165.600 136.950 ;
        RECT 170.400 136.350 171.600 137.100 ;
        RECT 160.950 133.950 163.050 136.050 ;
        RECT 163.950 133.950 166.050 136.050 ;
        RECT 166.950 133.950 169.050 136.050 ;
        RECT 169.950 133.950 172.050 136.050 ;
        RECT 161.400 131.400 162.600 133.650 ;
        RECT 167.400 132.000 168.600 133.650 ;
        RECT 161.400 115.050 162.450 131.400 ;
        RECT 166.950 127.950 169.050 132.000 ;
        RECT 176.400 123.450 177.450 139.950 ;
        RECT 182.400 138.600 183.450 145.950 ;
        RECT 182.400 136.350 183.600 138.600 ;
        RECT 188.400 138.450 189.600 138.600 ;
        RECT 191.400 138.450 192.450 148.950 ;
        RECT 188.400 137.400 192.450 138.450 ;
        RECT 188.400 136.350 189.600 137.400 ;
        RECT 181.950 133.950 184.050 136.050 ;
        RECT 184.950 133.950 187.050 136.050 ;
        RECT 187.950 133.950 190.050 136.050 ;
        RECT 193.950 133.950 196.050 136.050 ;
        RECT 185.400 132.000 186.600 133.650 ;
        RECT 184.950 127.950 187.050 132.000 ;
        RECT 173.400 122.400 177.450 123.450 ;
        RECT 173.400 115.050 174.450 122.400 ;
        RECT 194.400 118.050 195.450 133.950 ;
        RECT 175.950 115.950 178.050 118.050 ;
        RECT 193.950 115.950 196.050 118.050 ;
        RECT 160.800 112.950 162.900 115.050 ;
        RECT 163.950 112.950 166.050 115.050 ;
        RECT 172.950 112.950 175.050 115.050 ;
        RECT 157.950 109.950 160.050 112.050 ;
        RECT 152.400 103.350 153.600 105.000 ;
        RECT 154.950 103.950 157.050 106.050 ;
        RECT 130.950 100.950 133.050 103.050 ;
        RECT 133.950 100.950 136.050 103.050 ;
        RECT 139.950 100.950 142.050 103.050 ;
        RECT 145.950 100.950 148.050 103.050 ;
        RECT 148.950 100.950 151.050 103.050 ;
        RECT 151.950 100.950 154.050 103.050 ;
        RECT 131.400 99.000 132.600 100.650 ;
        RECT 124.950 94.950 127.050 97.050 ;
        RECT 130.950 94.950 133.050 99.000 ;
        RECT 140.400 94.050 141.450 100.950 ;
        RECT 142.950 97.950 145.050 100.050 ;
        RECT 149.400 98.400 150.600 100.650 ;
        RECT 139.950 91.950 142.050 94.050 ;
        RECT 115.950 88.950 118.050 91.050 ;
        RECT 121.950 88.950 124.050 91.050 ;
        RECT 115.950 70.950 118.050 73.050 ;
        RECT 127.950 70.950 130.050 73.050 ;
        RECT 116.400 67.050 117.450 70.950 ;
        RECT 115.950 64.950 118.050 67.050 ;
        RECT 79.950 61.950 82.050 64.050 ;
        RECT 94.950 61.950 97.050 64.050 ;
        RECT 80.400 60.450 81.600 60.600 ;
        RECT 77.400 59.400 81.600 60.450 ;
        RECT 68.400 58.350 69.600 59.100 ;
        RECT 58.950 55.950 61.050 58.050 ;
        RECT 61.950 55.950 64.050 58.050 ;
        RECT 64.950 55.950 67.050 58.050 ;
        RECT 67.950 55.950 70.050 58.050 ;
        RECT 59.400 54.900 60.600 55.650 ;
        RECT 58.950 52.800 61.050 54.900 ;
        RECT 65.400 53.400 66.600 55.650 ;
        RECT 52.950 46.950 55.050 49.050 ;
        RECT 61.950 46.950 64.050 49.050 ;
        RECT 46.950 43.950 49.050 46.050 ;
        RECT 47.400 27.600 48.450 43.950 ;
        RECT 62.400 42.450 63.450 46.950 ;
        RECT 65.400 46.050 66.450 53.400 ;
        RECT 64.950 43.950 67.050 46.050 ;
        RECT 70.950 43.950 73.050 46.050 ;
        RECT 67.950 42.450 70.050 43.050 ;
        RECT 62.400 41.400 70.050 42.450 ;
        RECT 67.950 40.950 70.050 41.400 ;
        RECT 64.950 37.950 67.050 40.050 ;
        RECT 65.400 34.050 66.450 37.950 ;
        RECT 64.950 31.950 67.050 34.050 ;
        RECT 47.400 25.350 48.600 27.600 ;
        RECT 52.950 26.100 55.050 28.200 ;
        RECT 65.400 27.600 66.450 31.950 ;
        RECT 71.400 27.600 72.450 43.950 ;
        RECT 74.400 31.050 75.450 59.100 ;
        RECT 80.400 58.350 81.600 59.400 ;
        RECT 85.950 59.100 88.050 61.200 ;
        RECT 86.400 58.350 87.600 59.100 ;
        RECT 79.950 55.950 82.050 58.050 ;
        RECT 82.950 55.950 85.050 58.050 ;
        RECT 85.950 55.950 88.050 58.050 ;
        RECT 88.950 55.950 91.050 58.050 ;
        RECT 83.400 54.000 84.600 55.650 ;
        RECT 89.400 54.000 90.600 55.650 ;
        RECT 82.950 49.950 85.050 54.000 ;
        RECT 88.950 49.950 91.050 54.000 ;
        RECT 91.950 48.450 94.050 49.050 ;
        RECT 86.400 47.400 94.050 48.450 ;
        RECT 86.400 43.050 87.450 47.400 ;
        RECT 91.950 46.950 94.050 47.400 ;
        RECT 88.950 43.950 91.050 46.050 ;
        RECT 85.950 40.950 88.050 43.050 ;
        RECT 73.950 28.950 76.050 31.050 ;
        RECT 53.400 25.350 54.600 26.100 ;
        RECT 65.400 25.350 66.600 27.600 ;
        RECT 71.400 25.350 72.600 27.600 ;
        RECT 79.950 25.950 82.050 28.050 ;
        RECT 89.400 27.600 90.450 43.950 ;
        RECT 95.400 31.050 96.450 61.950 ;
        RECT 100.950 60.000 103.050 64.050 ;
        RECT 101.400 58.350 102.600 60.000 ;
        RECT 106.950 59.100 109.050 61.200 ;
        RECT 107.400 58.350 108.600 59.100 ;
        RECT 100.950 55.950 103.050 58.050 ;
        RECT 103.950 55.950 106.050 58.050 ;
        RECT 106.950 55.950 109.050 58.050 ;
        RECT 109.950 55.950 112.050 58.050 ;
        RECT 104.400 53.400 105.600 55.650 ;
        RECT 110.400 53.400 111.600 55.650 ;
        RECT 104.400 49.050 105.450 53.400 ;
        RECT 110.400 49.050 111.450 53.400 ;
        RECT 112.950 52.950 115.050 55.050 ;
        RECT 103.950 46.950 106.050 49.050 ;
        RECT 109.950 46.950 112.050 49.050 ;
        RECT 113.400 37.050 114.450 52.950 ;
        RECT 112.950 34.950 115.050 37.050 ;
        RECT 103.950 31.950 106.050 34.050 ;
        RECT 109.950 31.950 112.050 34.050 ;
        RECT 94.950 28.950 97.050 31.050 ;
        RECT 104.400 28.050 105.450 31.950 ;
        RECT 43.950 22.950 46.050 25.050 ;
        RECT 46.950 22.950 49.050 25.050 ;
        RECT 49.950 22.950 52.050 25.050 ;
        RECT 52.950 22.950 55.050 25.050 ;
        RECT 64.950 22.950 67.050 25.050 ;
        RECT 67.950 22.950 70.050 25.050 ;
        RECT 70.950 22.950 73.050 25.050 ;
        RECT 73.950 22.950 76.050 25.050 ;
        RECT 17.400 16.050 18.450 20.400 ;
        RECT 31.950 19.800 34.050 21.900 ;
        RECT 37.950 19.950 40.050 22.050 ;
        RECT 44.400 21.900 45.600 22.650 ;
        RECT 43.950 19.800 46.050 21.900 ;
        RECT 50.400 20.400 51.600 22.650 ;
        RECT 68.400 21.000 69.600 22.650 ;
        RECT 50.400 16.050 51.450 20.400 ;
        RECT 67.950 16.950 70.050 21.000 ;
        RECT 74.400 20.400 75.600 22.650 ;
        RECT 74.400 16.050 75.450 20.400 ;
        RECT 16.950 13.950 19.050 16.050 ;
        RECT 49.950 13.950 52.050 16.050 ;
        RECT 73.950 13.950 76.050 16.050 ;
        RECT 80.400 7.050 81.450 25.950 ;
        RECT 89.400 25.350 90.600 27.600 ;
        RECT 95.400 27.450 96.600 27.600 ;
        RECT 95.400 26.400 102.450 27.450 ;
        RECT 95.400 25.350 96.600 26.400 ;
        RECT 85.950 22.950 88.050 25.050 ;
        RECT 88.950 22.950 91.050 25.050 ;
        RECT 91.950 22.950 94.050 25.050 ;
        RECT 94.950 22.950 97.050 25.050 ;
        RECT 86.400 21.900 87.600 22.650 ;
        RECT 92.400 21.900 93.600 22.650 ;
        RECT 85.950 19.800 88.050 21.900 ;
        RECT 86.400 16.050 87.450 19.800 ;
        RECT 91.950 16.950 94.050 21.900 ;
        RECT 101.400 16.050 102.450 26.400 ;
        RECT 103.950 25.950 106.050 28.050 ;
        RECT 110.400 27.600 111.450 31.950 ;
        RECT 116.400 27.600 117.450 64.950 ;
        RECT 128.400 64.050 129.450 70.950 ;
        RECT 143.400 67.050 144.450 97.950 ;
        RECT 149.400 91.050 150.450 98.400 ;
        RECT 158.400 97.050 159.450 109.950 ;
        RECT 164.400 105.600 165.450 112.950 ;
        RECT 169.950 109.950 172.050 112.050 ;
        RECT 170.400 105.600 171.450 109.950 ;
        RECT 176.400 105.600 177.450 115.950 ;
        RECT 197.400 112.050 198.450 169.950 ;
        RECT 203.400 138.600 204.450 176.400 ;
        RECT 206.400 175.050 207.450 205.950 ;
        RECT 214.950 199.950 217.050 202.050 ;
        RECT 208.950 181.950 211.050 187.050 ;
        RECT 215.400 183.600 216.450 199.950 ;
        RECT 230.400 199.050 231.450 208.800 ;
        RECT 229.950 196.950 232.050 199.050 ;
        RECT 239.400 196.050 240.450 235.950 ;
        RECT 245.400 223.050 246.450 254.400 ;
        RECT 251.400 244.050 252.450 260.100 ;
        RECT 250.950 241.950 253.050 244.050 ;
        RECT 247.950 238.950 250.050 241.050 ;
        RECT 248.400 235.050 249.450 238.950 ;
        RECT 254.400 238.050 255.450 262.950 ;
        RECT 263.400 262.200 264.450 280.950 ;
        RECT 262.950 260.100 265.050 262.200 ;
        RECT 268.950 260.100 271.050 262.200 ;
        RECT 263.400 259.350 264.600 260.100 ;
        RECT 257.100 256.950 259.200 259.050 ;
        RECT 262.500 256.950 264.600 259.050 ;
        RECT 265.800 256.950 267.900 259.050 ;
        RECT 257.400 255.000 258.600 256.650 ;
        RECT 256.950 250.950 259.050 255.000 ;
        RECT 266.400 254.400 267.600 256.650 ;
        RECT 253.950 235.950 256.050 238.050 ;
        RECT 247.950 232.950 250.050 235.050 ;
        RECT 266.400 226.050 267.450 254.400 ;
        RECT 265.950 223.950 268.050 226.050 ;
        RECT 269.400 223.050 270.450 260.100 ;
        RECT 272.400 253.050 273.450 283.650 ;
        RECT 271.950 250.950 274.050 253.050 ;
        RECT 275.400 234.450 276.450 283.950 ;
        RECT 284.400 280.050 285.450 286.950 ;
        RECT 286.950 283.950 289.050 286.050 ;
        RECT 283.950 277.950 286.050 280.050 ;
        RECT 278.400 256.950 280.500 259.050 ;
        RECT 283.800 256.950 285.900 259.050 ;
        RECT 284.400 254.400 285.600 256.650 ;
        RECT 280.950 247.950 283.050 250.050 ;
        RECT 277.950 234.450 280.050 235.050 ;
        RECT 275.400 233.400 280.050 234.450 ;
        RECT 277.950 232.950 280.050 233.400 ;
        RECT 244.950 220.950 247.050 223.050 ;
        RECT 268.950 220.950 271.050 223.050 ;
        RECT 278.400 217.200 279.450 232.950 ;
        RECT 247.950 215.100 250.050 217.200 ;
        RECT 253.950 215.100 256.050 217.200 ;
        RECT 259.950 215.100 262.050 217.200 ;
        RECT 265.950 215.100 268.050 217.200 ;
        RECT 271.950 215.100 274.050 217.200 ;
        RECT 277.950 215.100 280.050 217.200 ;
        RECT 248.400 214.350 249.600 215.100 ;
        RECT 254.400 214.350 255.600 215.100 ;
        RECT 244.950 211.950 247.050 214.050 ;
        RECT 247.950 211.950 250.050 214.050 ;
        RECT 250.950 211.950 253.050 214.050 ;
        RECT 253.950 211.950 256.050 214.050 ;
        RECT 245.400 211.050 246.600 211.650 ;
        RECT 241.950 209.400 246.600 211.050 ;
        RECT 251.400 209.400 252.600 211.650 ;
        RECT 241.950 208.950 246.000 209.400 ;
        RECT 251.400 199.050 252.450 209.400 ;
        RECT 250.950 196.950 253.050 199.050 ;
        RECT 232.950 193.950 235.050 196.050 ;
        RECT 238.950 193.950 241.050 196.050 ;
        RECT 215.400 181.350 216.600 183.600 ;
        RECT 220.950 182.100 223.050 186.900 ;
        RECT 229.950 184.950 232.050 187.050 ;
        RECT 221.400 181.350 222.600 182.100 ;
        RECT 211.950 178.950 214.050 181.050 ;
        RECT 214.950 178.950 217.050 181.050 ;
        RECT 217.950 178.950 220.050 181.050 ;
        RECT 220.950 178.950 223.050 181.050 ;
        RECT 223.950 178.950 226.050 181.050 ;
        RECT 212.400 176.400 213.600 178.650 ;
        RECT 218.400 176.400 219.600 178.650 ;
        RECT 224.400 177.000 225.600 178.650 ;
        RECT 205.950 172.950 208.050 175.050 ;
        RECT 212.400 166.050 213.450 176.400 ;
        RECT 214.950 172.950 217.050 175.050 ;
        RECT 211.950 163.950 214.050 166.050 ;
        RECT 203.400 136.350 204.600 138.600 ;
        RECT 202.950 133.950 205.050 136.050 ;
        RECT 205.950 133.950 208.050 136.050 ;
        RECT 208.950 133.950 211.050 136.050 ;
        RECT 206.400 131.400 207.600 133.650 ;
        RECT 202.950 127.950 205.050 130.050 ;
        RECT 199.950 121.950 202.050 124.050 ;
        RECT 184.950 109.950 187.050 112.050 ;
        RECT 196.950 109.950 199.050 112.050 ;
        RECT 164.400 103.350 165.600 105.600 ;
        RECT 170.400 103.350 171.600 105.600 ;
        RECT 176.400 103.350 177.600 105.600 ;
        RECT 181.950 103.950 184.050 106.050 ;
        RECT 163.950 100.950 166.050 103.050 ;
        RECT 166.950 100.950 169.050 103.050 ;
        RECT 169.950 100.950 172.050 103.050 ;
        RECT 172.950 100.950 175.050 103.050 ;
        RECT 175.950 100.950 178.050 103.050 ;
        RECT 167.400 99.900 168.600 100.650 ;
        RECT 173.400 99.900 174.600 100.650 ;
        RECT 166.950 97.800 169.050 99.900 ;
        RECT 172.950 97.800 175.050 99.900 ;
        RECT 157.950 94.950 160.050 97.050 ;
        RECT 163.950 94.950 166.050 97.050 ;
        RECT 148.950 88.950 151.050 91.050 ;
        RECT 157.950 82.950 160.050 85.050 ;
        RECT 151.950 73.950 154.050 76.050 ;
        RECT 145.950 67.950 148.050 70.050 ;
        RECT 142.950 64.950 145.050 67.050 ;
        RECT 124.950 60.000 127.050 64.050 ;
        RECT 127.950 61.950 130.050 64.050 ;
        RECT 125.400 58.350 126.600 60.000 ;
        RECT 130.800 59.100 132.900 61.200 ;
        RECT 131.400 58.350 132.600 59.100 ;
        RECT 133.950 58.950 136.050 64.050 ;
        RECT 146.400 60.600 147.450 67.950 ;
        RECT 152.400 61.200 153.450 73.950 ;
        RECT 146.400 58.350 147.600 60.600 ;
        RECT 151.950 59.100 154.050 61.200 ;
        RECT 152.400 58.350 153.600 59.100 ;
        RECT 121.950 55.950 124.050 58.050 ;
        RECT 124.950 55.950 127.050 58.050 ;
        RECT 127.950 55.950 130.050 58.050 ;
        RECT 130.950 55.950 133.050 58.050 ;
        RECT 142.950 55.950 145.050 58.050 ;
        RECT 145.950 55.950 148.050 58.050 ;
        RECT 148.950 55.950 151.050 58.050 ;
        RECT 151.950 55.950 154.050 58.050 ;
        RECT 122.400 53.400 123.600 55.650 ;
        RECT 128.400 54.900 129.600 55.650 ;
        RECT 122.400 46.050 123.450 53.400 ;
        RECT 127.950 52.800 130.050 54.900 ;
        RECT 143.400 53.400 144.600 55.650 ;
        RECT 149.400 54.900 150.600 55.650 ;
        RECT 143.400 49.050 144.450 53.400 ;
        RECT 148.950 52.800 151.050 54.900 ;
        RECT 142.950 46.950 145.050 49.050 ;
        RECT 149.400 46.050 150.450 52.800 ;
        RECT 121.950 43.950 124.050 46.050 ;
        RECT 148.950 43.950 151.050 46.050 ;
        RECT 158.400 43.050 159.450 82.950 ;
        RECT 164.400 64.050 165.450 94.950 ;
        RECT 167.400 82.050 168.450 97.800 ;
        RECT 173.400 94.050 174.450 97.800 ;
        RECT 172.950 91.950 175.050 94.050 ;
        RECT 178.950 88.950 181.050 91.050 ;
        RECT 166.950 79.950 169.050 82.050 ;
        RECT 179.400 70.050 180.450 88.950 ;
        RECT 178.950 67.950 181.050 70.050 ;
        RECT 169.950 64.950 172.050 67.050 ;
        RECT 163.950 60.000 166.050 64.050 ;
        RECT 170.400 60.600 171.450 64.950 ;
        RECT 182.400 64.050 183.450 103.950 ;
        RECT 185.400 99.900 186.450 109.950 ;
        RECT 200.400 109.050 201.450 121.950 ;
        RECT 199.950 106.950 202.050 109.050 ;
        RECT 203.400 106.200 204.450 127.950 ;
        RECT 206.400 118.050 207.450 131.400 ;
        RECT 215.400 127.050 216.450 172.950 ;
        RECT 218.400 172.050 219.450 176.400 ;
        RECT 223.950 174.450 226.050 177.000 ;
        RECT 221.400 173.400 226.050 174.450 ;
        RECT 217.950 169.950 220.050 172.050 ;
        RECT 221.400 148.050 222.450 173.400 ;
        RECT 223.950 172.950 226.050 173.400 ;
        RECT 223.950 169.800 226.050 171.900 ;
        RECT 224.400 166.050 225.450 169.800 ;
        RECT 223.950 163.950 226.050 166.050 ;
        RECT 230.400 160.050 231.450 184.950 ;
        RECT 233.400 184.050 234.450 193.950 ;
        RECT 260.400 193.050 261.450 215.100 ;
        RECT 266.400 214.350 267.600 215.100 ;
        RECT 272.400 214.350 273.600 215.100 ;
        RECT 265.950 211.950 268.050 214.050 ;
        RECT 268.950 211.950 271.050 214.050 ;
        RECT 271.950 211.950 274.050 214.050 ;
        RECT 274.950 211.950 277.050 214.050 ;
        RECT 269.400 210.900 270.600 211.650 ;
        RECT 275.400 210.900 276.600 211.650 ;
        RECT 268.950 208.800 271.050 210.900 ;
        RECT 274.950 208.800 277.050 210.900 ;
        RECT 271.950 202.950 274.050 205.050 ;
        RECT 259.950 190.950 262.050 193.050 ;
        RECT 232.950 181.950 235.050 184.050 ;
        RECT 238.950 182.100 241.050 184.200 ;
        RECT 247.950 182.100 250.050 184.200 ;
        RECT 239.400 181.350 240.600 182.100 ;
        RECT 235.950 178.950 238.050 181.050 ;
        RECT 238.950 178.950 241.050 181.050 ;
        RECT 241.950 178.950 244.050 181.050 ;
        RECT 236.400 177.900 237.600 178.650 ;
        RECT 235.950 172.950 238.050 177.900 ;
        RECT 244.950 169.950 247.050 172.050 ;
        RECT 235.950 166.950 238.050 169.050 ;
        RECT 229.950 159.450 232.050 160.050 ;
        RECT 229.950 158.400 234.450 159.450 ;
        RECT 229.950 157.950 232.050 158.400 ;
        RECT 223.950 154.950 226.050 157.050 ;
        RECT 220.950 145.950 223.050 148.050 ;
        RECT 224.400 138.600 225.450 154.950 ;
        RECT 224.400 136.350 225.600 138.600 ;
        RECT 229.950 138.000 232.050 142.050 ;
        RECT 233.400 139.050 234.450 158.400 ;
        RECT 230.400 136.350 231.600 138.000 ;
        RECT 232.950 136.950 235.050 139.050 ;
        RECT 220.950 133.950 223.050 136.050 ;
        RECT 223.950 133.950 226.050 136.050 ;
        RECT 226.950 133.950 229.050 136.050 ;
        RECT 229.950 133.950 232.050 136.050 ;
        RECT 221.400 132.000 222.600 133.650 ;
        RECT 227.400 132.900 228.600 133.650 ;
        RECT 220.950 127.950 223.050 132.000 ;
        RECT 226.950 130.800 229.050 132.900 ;
        RECT 236.400 127.050 237.450 166.950 ;
        RECT 241.950 141.450 244.050 141.900 ;
        RECT 245.400 141.450 246.450 169.950 ;
        RECT 248.400 169.050 249.450 182.100 ;
        RECT 257.100 178.950 259.200 181.050 ;
        RECT 262.500 178.950 264.600 181.050 ;
        RECT 253.950 175.800 256.050 177.900 ;
        RECT 257.400 176.400 258.600 178.650 ;
        RECT 247.950 166.950 250.050 169.050 ;
        RECT 250.950 145.950 253.050 148.050 ;
        RECT 241.950 140.400 246.450 141.450 ;
        RECT 241.950 139.800 244.050 140.400 ;
        RECT 238.950 136.950 241.050 139.050 ;
        RECT 242.400 138.600 243.450 139.800 ;
        RECT 251.400 138.600 252.450 145.950 ;
        RECT 239.400 132.900 240.450 136.950 ;
        RECT 242.400 136.350 243.600 138.600 ;
        RECT 251.400 136.350 252.600 138.600 ;
        RECT 242.100 133.950 244.200 136.050 ;
        RECT 247.500 133.950 249.600 136.050 ;
        RECT 250.800 133.950 252.900 136.050 ;
        RECT 248.400 132.900 249.600 133.650 ;
        RECT 238.950 130.800 241.050 132.900 ;
        RECT 247.950 130.800 250.050 132.900 ;
        RECT 214.950 124.950 217.050 127.050 ;
        RECT 229.950 124.950 232.050 127.050 ;
        RECT 235.950 124.950 238.050 127.050 ;
        RECT 205.950 115.950 208.050 118.050 ;
        RECT 211.950 112.950 214.050 115.050 ;
        RECT 220.950 112.950 223.050 115.050 ;
        RECT 208.950 109.950 211.050 112.050 ;
        RECT 190.950 104.100 193.050 106.200 ;
        RECT 196.950 104.100 199.050 106.200 ;
        RECT 202.800 104.100 204.900 106.200 ;
        RECT 205.950 104.100 208.050 106.200 ;
        RECT 191.400 103.350 192.600 104.100 ;
        RECT 197.400 103.350 198.600 104.100 ;
        RECT 190.950 100.950 193.050 103.050 ;
        RECT 193.950 100.950 196.050 103.050 ;
        RECT 196.950 100.950 199.050 103.050 ;
        RECT 199.950 100.950 202.050 103.050 ;
        RECT 194.400 99.900 195.600 100.650 ;
        RECT 184.950 97.800 187.050 99.900 ;
        RECT 193.950 97.800 196.050 99.900 ;
        RECT 200.400 98.400 201.600 100.650 ;
        RECT 206.400 99.450 207.450 104.100 ;
        RECT 203.400 98.400 207.450 99.450 ;
        RECT 209.400 99.450 210.450 109.950 ;
        RECT 212.400 106.050 213.450 112.950 ;
        RECT 211.950 103.950 214.050 106.050 ;
        RECT 214.950 104.100 217.050 106.200 ;
        RECT 221.400 105.600 222.450 112.950 ;
        RECT 215.400 103.350 216.600 104.100 ;
        RECT 221.400 103.350 222.600 105.600 ;
        RECT 214.950 100.950 217.050 103.050 ;
        RECT 217.950 100.950 220.050 103.050 ;
        RECT 220.950 100.950 223.050 103.050 ;
        RECT 223.950 100.950 226.050 103.050 ;
        RECT 218.400 99.900 219.600 100.650 ;
        RECT 224.400 99.900 225.600 100.650 ;
        RECT 209.400 98.400 213.450 99.450 ;
        RECT 200.400 97.050 201.450 98.400 ;
        RECT 199.950 94.950 202.050 97.050 ;
        RECT 190.950 85.950 193.050 88.050 ;
        RECT 191.400 67.050 192.450 85.950 ;
        RECT 200.400 79.050 201.450 94.950 ;
        RECT 199.950 76.950 202.050 79.050 ;
        RECT 190.950 64.950 193.050 67.050 ;
        RECT 164.400 58.350 165.600 60.000 ;
        RECT 170.400 58.350 171.600 60.600 ;
        RECT 175.950 58.950 178.050 64.050 ;
        RECT 181.950 61.950 184.050 64.050 ;
        RECT 191.400 60.600 192.450 64.950 ;
        RECT 199.950 61.950 202.050 64.050 ;
        RECT 185.400 60.450 186.600 60.600 ;
        RECT 179.400 59.400 186.600 60.450 ;
        RECT 163.950 55.950 166.050 58.050 ;
        RECT 166.950 55.950 169.050 58.050 ;
        RECT 169.950 55.950 172.050 58.050 ;
        RECT 172.950 55.950 175.050 58.050 ;
        RECT 167.400 53.400 168.600 55.650 ;
        RECT 173.400 54.900 174.600 55.650 ;
        RECT 157.950 40.950 160.050 43.050 ;
        RECT 133.950 37.950 136.050 40.050 ;
        RECT 154.950 37.950 157.050 40.050 ;
        RECT 127.950 34.950 130.050 37.050 ;
        RECT 121.950 28.950 124.050 31.050 ;
        RECT 110.400 25.350 111.600 27.600 ;
        RECT 116.400 25.350 117.600 27.600 ;
        RECT 106.950 22.950 109.050 25.050 ;
        RECT 109.950 22.950 112.050 25.050 ;
        RECT 112.950 22.950 115.050 25.050 ;
        RECT 115.950 22.950 118.050 25.050 ;
        RECT 107.400 21.900 108.600 22.650 ;
        RECT 106.950 19.800 109.050 21.900 ;
        RECT 113.400 20.400 114.600 22.650 ;
        RECT 113.400 18.450 114.450 20.400 ;
        RECT 110.400 17.400 114.450 18.450 ;
        RECT 110.400 16.050 111.450 17.400 ;
        RECT 122.400 16.050 123.450 28.950 ;
        RECT 128.400 27.600 129.450 34.950 ;
        RECT 134.400 27.600 135.450 37.950 ;
        RECT 155.400 34.050 156.450 37.950 ;
        RECT 154.950 31.950 157.050 34.050 ;
        RECT 128.400 25.350 129.600 27.600 ;
        RECT 134.400 25.350 135.600 27.600 ;
        RECT 148.950 27.000 151.050 31.050 ;
        RECT 155.400 27.600 156.450 31.950 ;
        RECT 167.400 28.050 168.450 53.400 ;
        RECT 172.950 52.800 175.050 54.900 ;
        RECT 175.950 46.950 178.050 49.050 ;
        RECT 172.950 37.950 175.050 40.050 ;
        RECT 173.400 30.450 174.450 37.950 ;
        RECT 170.400 29.400 174.450 30.450 ;
        RECT 149.400 25.350 150.600 27.000 ;
        RECT 155.400 25.350 156.600 27.600 ;
        RECT 163.950 25.950 166.050 28.050 ;
        RECT 166.950 25.950 169.050 28.050 ;
        RECT 170.400 27.600 171.450 29.400 ;
        RECT 176.400 28.050 177.450 46.950 ;
        RECT 127.950 22.950 130.050 25.050 ;
        RECT 130.950 22.950 133.050 25.050 ;
        RECT 133.950 22.950 136.050 25.050 ;
        RECT 136.950 22.950 139.050 25.050 ;
        RECT 148.950 22.950 151.050 25.050 ;
        RECT 151.950 22.950 154.050 25.050 ;
        RECT 154.950 22.950 157.050 25.050 ;
        RECT 157.950 22.950 160.050 25.050 ;
        RECT 131.400 21.900 132.600 22.650 ;
        RECT 130.950 19.800 133.050 21.900 ;
        RECT 137.400 21.000 138.600 22.650 ;
        RECT 152.400 21.000 153.600 22.650 ;
        RECT 158.400 21.900 159.600 22.650 ;
        RECT 164.400 21.900 165.450 25.950 ;
        RECT 170.400 25.350 171.600 27.600 ;
        RECT 175.950 25.950 178.050 28.050 ;
        RECT 169.950 22.950 172.050 25.050 ;
        RECT 172.950 22.950 175.050 25.050 ;
        RECT 173.400 21.900 174.600 22.650 ;
        RECT 179.400 22.050 180.450 59.400 ;
        RECT 185.400 58.350 186.600 59.400 ;
        RECT 191.400 58.350 192.600 60.600 ;
        RECT 184.950 55.950 187.050 58.050 ;
        RECT 187.950 55.950 190.050 58.050 ;
        RECT 190.950 55.950 193.050 58.050 ;
        RECT 193.950 55.950 196.050 58.050 ;
        RECT 188.400 54.000 189.600 55.650 ;
        RECT 194.400 54.900 195.600 55.650 ;
        RECT 187.950 49.950 190.050 54.000 ;
        RECT 193.950 52.800 196.050 54.900 ;
        RECT 196.950 40.950 199.050 43.050 ;
        RECT 197.400 34.050 198.450 40.950 ;
        RECT 200.400 40.050 201.450 61.950 ;
        RECT 203.400 61.050 204.450 98.400 ;
        RECT 202.950 58.950 205.050 61.050 ;
        RECT 205.950 60.000 208.050 64.050 ;
        RECT 212.400 61.200 213.450 98.400 ;
        RECT 217.950 97.800 220.050 99.900 ;
        RECT 223.950 97.800 226.050 99.900 ;
        RECT 223.950 91.950 226.050 94.050 ;
        RECT 224.400 85.050 225.450 91.950 ;
        RECT 223.800 82.950 225.900 85.050 ;
        RECT 230.400 64.050 231.450 124.950 ;
        RECT 236.400 121.050 237.450 124.950 ;
        RECT 254.400 121.050 255.450 175.800 ;
        RECT 257.400 160.050 258.450 176.400 ;
        RECT 256.950 157.950 259.050 160.050 ;
        RECT 256.950 142.950 259.050 145.050 ;
        RECT 235.950 118.950 238.050 121.050 ;
        RECT 253.950 118.950 256.050 121.050 ;
        RECT 257.400 115.050 258.450 142.950 ;
        RECT 259.950 138.600 264.000 139.050 ;
        RECT 259.950 136.950 264.600 138.600 ;
        RECT 263.400 136.350 264.600 136.950 ;
        RECT 262.950 133.950 265.050 136.050 ;
        RECT 265.950 133.950 268.050 136.050 ;
        RECT 266.400 131.400 267.600 133.650 ;
        RECT 266.400 127.050 267.450 131.400 ;
        RECT 265.950 124.950 268.050 127.050 ;
        RECT 266.400 115.050 267.450 124.950 ;
        RECT 268.950 115.950 271.050 118.050 ;
        RECT 250.950 112.950 253.050 115.050 ;
        RECT 256.950 112.950 259.050 115.050 ;
        RECT 265.950 112.950 268.050 115.050 ;
        RECT 235.950 109.950 238.050 112.050 ;
        RECT 241.950 109.950 244.050 112.050 ;
        RECT 236.400 105.600 237.450 109.950 ;
        RECT 242.400 105.600 243.450 109.950 ;
        RECT 236.400 103.350 237.600 105.600 ;
        RECT 242.400 103.350 243.600 105.600 ;
        RECT 235.950 100.950 238.050 103.050 ;
        RECT 238.950 100.950 241.050 103.050 ;
        RECT 241.950 100.950 244.050 103.050 ;
        RECT 244.950 100.950 247.050 103.050 ;
        RECT 239.400 99.900 240.600 100.650 ;
        RECT 245.400 99.900 246.600 100.650 ;
        RECT 238.950 97.800 241.050 99.900 ;
        RECT 244.950 97.800 247.050 99.900 ;
        RECT 247.950 97.950 250.050 100.050 ;
        RECT 248.400 88.050 249.450 97.950 ;
        RECT 251.400 91.050 252.450 112.950 ;
        RECT 262.950 109.950 265.050 112.050 ;
        RECT 253.950 105.600 258.000 106.050 ;
        RECT 263.400 105.600 264.450 109.950 ;
        RECT 266.400 109.050 267.450 112.950 ;
        RECT 265.950 106.950 268.050 109.050 ;
        RECT 269.400 106.050 270.450 115.950 ;
        RECT 253.950 103.950 258.600 105.600 ;
        RECT 257.400 103.350 258.600 103.950 ;
        RECT 263.400 103.350 264.600 105.600 ;
        RECT 268.950 103.950 271.050 106.050 ;
        RECT 256.950 100.950 259.050 103.050 ;
        RECT 259.950 100.950 262.050 103.050 ;
        RECT 262.950 100.950 265.050 103.050 ;
        RECT 265.950 100.950 268.050 103.050 ;
        RECT 260.400 99.900 261.600 100.650 ;
        RECT 266.400 99.900 267.600 100.650 ;
        RECT 259.950 97.800 262.050 99.900 ;
        RECT 265.950 97.800 268.050 99.900 ;
        RECT 268.950 97.950 271.050 100.050 ;
        RECT 260.400 96.450 261.450 97.800 ;
        RECT 257.400 95.400 261.450 96.450 ;
        RECT 250.950 88.950 253.050 91.050 ;
        RECT 247.950 85.950 250.050 88.050 ;
        RECT 251.400 76.050 252.450 88.950 ;
        RECT 257.400 88.050 258.450 95.400 ;
        RECT 262.950 94.950 265.050 97.050 ;
        RECT 259.950 91.950 262.050 94.050 ;
        RECT 256.950 85.950 259.050 88.050 ;
        RECT 260.400 82.050 261.450 91.950 ;
        RECT 259.950 79.950 262.050 82.050 ;
        RECT 238.950 73.950 241.050 76.050 ;
        RECT 250.950 73.950 253.050 76.050 ;
        RECT 239.400 67.050 240.450 73.950 ;
        RECT 241.950 70.950 244.050 73.050 ;
        RECT 238.950 64.950 241.050 67.050 ;
        RECT 229.950 61.950 232.050 64.050 ;
        RECT 206.400 58.350 207.600 60.000 ;
        RECT 211.950 59.100 214.050 61.200 ;
        RECT 212.400 58.350 213.600 59.100 ;
        RECT 220.950 58.950 223.050 61.050 ;
        RECT 226.950 59.100 229.050 61.200 ;
        RECT 232.950 60.000 235.050 64.050 ;
        RECT 205.950 55.950 208.050 58.050 ;
        RECT 208.950 55.950 211.050 58.050 ;
        RECT 211.950 55.950 214.050 58.050 ;
        RECT 214.950 55.950 217.050 58.050 ;
        RECT 209.400 54.900 210.600 55.650 ;
        RECT 215.400 54.900 216.600 55.650 ;
        RECT 208.950 52.800 211.050 54.900 ;
        RECT 214.950 52.800 217.050 54.900 ;
        RECT 217.950 52.950 220.050 55.050 ;
        RECT 209.400 40.050 210.450 52.800 ;
        RECT 211.950 46.950 214.050 49.050 ;
        RECT 212.400 43.050 213.450 46.950 ;
        RECT 215.400 46.050 216.450 52.800 ;
        RECT 214.950 43.950 217.050 46.050 ;
        RECT 211.950 40.950 214.050 43.050 ;
        RECT 218.400 42.450 219.450 52.950 ;
        RECT 215.400 41.400 219.450 42.450 ;
        RECT 199.800 37.950 201.900 40.050 ;
        RECT 202.950 37.950 205.050 40.050 ;
        RECT 208.950 37.950 211.050 40.050 ;
        RECT 184.950 31.950 187.050 34.050 ;
        RECT 196.950 31.950 199.050 34.050 ;
        RECT 199.950 31.950 202.050 34.050 ;
        RECT 185.400 27.600 186.450 31.950 ;
        RECT 185.400 25.350 186.600 27.600 ;
        RECT 190.950 27.000 193.050 31.050 ;
        RECT 191.400 25.350 192.600 27.000 ;
        RECT 184.950 22.950 187.050 25.050 ;
        RECT 187.950 22.950 190.050 25.050 ;
        RECT 190.950 22.950 193.050 25.050 ;
        RECT 193.950 22.950 196.050 25.050 ;
        RECT 136.950 16.950 139.050 21.000 ;
        RECT 151.950 16.950 154.050 21.000 ;
        RECT 157.950 19.800 160.050 21.900 ;
        RECT 163.950 19.800 166.050 21.900 ;
        RECT 172.950 19.800 175.050 21.900 ;
        RECT 178.950 19.950 181.050 22.050 ;
        RECT 188.400 21.900 189.600 22.650 ;
        RECT 194.400 21.900 195.600 22.650 ;
        RECT 200.400 22.050 201.450 31.950 ;
        RECT 203.400 28.050 204.450 37.950 ;
        RECT 215.400 34.050 216.450 41.400 ;
        RECT 217.950 34.950 220.050 37.050 ;
        RECT 205.950 31.950 208.050 34.050 ;
        RECT 214.950 31.950 217.050 34.050 ;
        RECT 202.950 25.950 205.050 28.050 ;
        RECT 206.400 27.600 207.450 31.950 ;
        RECT 206.400 25.350 207.600 27.600 ;
        RECT 211.950 26.100 214.050 28.200 ;
        RECT 218.400 27.450 219.450 34.950 ;
        RECT 221.400 31.050 222.450 58.950 ;
        RECT 227.400 58.350 228.600 59.100 ;
        RECT 233.400 58.350 234.600 60.000 ;
        RECT 226.950 55.950 229.050 58.050 ;
        RECT 229.950 55.950 232.050 58.050 ;
        RECT 232.950 55.950 235.050 58.050 ;
        RECT 235.950 55.950 238.050 58.050 ;
        RECT 230.400 53.400 231.600 55.650 ;
        RECT 236.400 55.050 237.600 55.650 ;
        RECT 236.400 53.400 241.050 55.050 ;
        RECT 223.950 46.950 226.050 49.050 ;
        RECT 224.400 43.050 225.450 46.950 ;
        RECT 223.950 40.950 226.050 43.050 ;
        RECT 230.400 40.050 231.450 53.400 ;
        RECT 237.000 52.950 241.050 53.400 ;
        RECT 242.400 49.050 243.450 70.950 ;
        RECT 250.950 60.000 253.050 64.050 ;
        RECT 251.400 58.350 252.600 60.000 ;
        RECT 256.950 59.100 259.050 61.200 ;
        RECT 257.400 58.350 258.600 59.100 ;
        RECT 247.950 55.950 250.050 58.050 ;
        RECT 250.950 55.950 253.050 58.050 ;
        RECT 253.950 55.950 256.050 58.050 ;
        RECT 256.950 55.950 259.050 58.050 ;
        RECT 248.400 53.400 249.600 55.650 ;
        RECT 254.400 53.400 255.600 55.650 ;
        RECT 263.400 54.450 264.450 94.950 ;
        RECT 269.400 88.050 270.450 97.950 ;
        RECT 272.400 93.450 273.450 202.950 ;
        RECT 275.400 175.050 276.450 208.800 ;
        RECT 281.400 205.050 282.450 247.950 ;
        RECT 284.400 244.050 285.450 254.400 ;
        RECT 287.400 250.050 288.450 283.950 ;
        RECT 293.400 274.050 294.450 287.400 ;
        RECT 292.950 271.950 295.050 274.050 ;
        RECT 289.950 260.100 292.050 262.200 ;
        RECT 298.950 260.100 301.050 262.200 ;
        RECT 302.400 262.050 303.450 328.950 ;
        RECT 305.400 310.050 306.450 332.400 ;
        RECT 304.950 307.950 307.050 310.050 ;
        RECT 304.950 304.800 307.050 306.900 ;
        RECT 305.400 289.050 306.450 304.800 ;
        RECT 304.950 286.950 307.050 289.050 ;
        RECT 286.950 247.950 289.050 250.050 ;
        RECT 283.950 241.950 286.050 244.050 ;
        RECT 280.950 202.950 283.050 205.050 ;
        RECT 284.400 202.050 285.450 241.950 ;
        RECT 286.950 220.950 289.050 223.050 ;
        RECT 287.400 216.600 288.450 220.950 ;
        RECT 290.400 220.050 291.450 260.100 ;
        RECT 299.400 259.350 300.600 260.100 ;
        RECT 301.950 259.950 304.050 262.050 ;
        RECT 295.950 256.950 298.050 259.050 ;
        RECT 298.950 256.950 301.050 259.050 ;
        RECT 296.400 254.400 297.600 256.650 ;
        RECT 296.400 253.050 297.450 254.400 ;
        RECT 301.950 253.950 304.050 256.050 ;
        RECT 295.950 250.950 298.050 253.050 ;
        RECT 296.400 238.050 297.450 250.950 ;
        RECT 298.950 247.950 301.050 250.050 ;
        RECT 295.950 235.950 298.050 238.050 ;
        RECT 295.950 220.950 298.050 223.050 ;
        RECT 289.950 217.950 292.050 220.050 ;
        RECT 287.400 214.350 288.600 216.600 ;
        RECT 287.100 211.950 289.200 214.050 ;
        RECT 292.500 211.950 294.600 214.050 ;
        RECT 286.950 205.950 289.050 208.050 ;
        RECT 283.950 199.950 286.050 202.050 ;
        RECT 287.400 189.450 288.450 205.950 ;
        RECT 287.400 187.200 288.600 189.450 ;
        RECT 282.900 183.900 285.000 185.700 ;
        RECT 286.800 184.800 288.900 186.900 ;
        RECT 290.100 186.300 292.200 188.400 ;
        RECT 281.400 182.700 290.100 183.900 ;
        RECT 278.100 178.950 280.200 181.050 ;
        RECT 278.400 177.900 279.600 178.650 ;
        RECT 277.950 175.800 280.050 177.900 ;
        RECT 274.950 172.950 277.050 175.050 ;
        RECT 281.400 173.700 282.300 182.700 ;
        RECT 288.000 181.800 290.100 182.700 ;
        RECT 291.000 180.900 291.900 186.300 ;
        RECT 293.400 183.450 294.600 183.600 ;
        RECT 296.400 183.450 297.450 220.950 ;
        RECT 299.400 208.050 300.450 247.950 ;
        RECT 302.400 244.050 303.450 253.950 ;
        RECT 308.400 250.050 309.450 365.400 ;
        RECT 311.400 365.400 312.600 367.650 ;
        RECT 317.400 366.000 318.600 367.650 ;
        RECT 326.400 367.050 327.450 371.100 ;
        RECT 335.400 370.350 336.600 371.100 ;
        RECT 331.950 367.950 334.050 370.050 ;
        RECT 334.950 367.950 337.050 370.050 ;
        RECT 340.950 367.950 343.050 370.050 ;
        RECT 325.950 366.450 328.050 367.050 ;
        RECT 332.400 366.900 333.600 367.650 ;
        RECT 341.400 366.900 342.600 367.650 ;
        RECT 311.400 358.050 312.450 365.400 ;
        RECT 316.950 361.950 319.050 366.000 ;
        RECT 325.950 365.400 330.450 366.450 ;
        RECT 325.950 364.950 328.050 365.400 ;
        RECT 310.950 355.950 313.050 358.050 ;
        RECT 325.950 355.950 328.050 358.050 ;
        RECT 313.950 352.950 316.050 355.050 ;
        RECT 310.950 346.950 313.050 349.050 ;
        RECT 311.400 340.050 312.450 346.950 ;
        RECT 314.400 343.050 315.450 352.950 ;
        RECT 313.950 340.950 316.050 343.050 ;
        RECT 310.950 337.950 313.050 340.050 ;
        RECT 316.950 338.100 319.050 340.200 ;
        RECT 317.400 337.350 318.600 338.100 ;
        RECT 313.950 334.950 316.050 337.050 ;
        RECT 316.950 334.950 319.050 337.050 ;
        RECT 319.950 334.950 322.050 337.050 ;
        RECT 314.400 333.900 315.600 334.650 ;
        RECT 313.950 331.800 316.050 333.900 ;
        RECT 320.400 333.000 321.600 334.650 ;
        RECT 314.400 328.050 315.450 331.800 ;
        RECT 319.950 328.950 322.050 333.000 ;
        RECT 326.400 331.050 327.450 355.950 ;
        RECT 329.400 333.900 330.450 365.400 ;
        RECT 331.950 364.800 334.050 366.900 ;
        RECT 340.950 364.800 343.050 366.900 ;
        RECT 334.950 361.950 337.050 364.050 ;
        RECT 335.400 339.600 336.450 361.950 ;
        RECT 347.250 359.700 348.450 372.600 ;
        RECT 346.350 357.600 348.450 359.700 ;
        RECT 350.400 358.050 351.450 391.950 ;
        RECT 361.650 379.500 363.750 380.400 ;
        RECT 361.650 378.300 365.850 379.500 ;
        RECT 352.950 371.100 355.050 373.200 ;
        RECT 358.950 371.100 361.050 373.200 ;
        RECT 353.400 367.050 354.450 371.100 ;
        RECT 359.400 370.350 360.600 371.100 ;
        RECT 358.800 367.950 360.900 370.050 ;
        RECT 352.950 364.950 355.050 367.050 ;
        RECT 364.650 359.700 365.850 378.300 ;
        RECT 368.400 372.600 369.450 397.950 ;
        RECT 392.400 379.050 393.450 406.950 ;
        RECT 401.400 406.050 402.450 410.400 ;
        RECT 406.950 409.800 409.050 411.900 ;
        RECT 400.950 403.950 403.050 406.050 ;
        RECT 413.400 379.050 414.450 436.950 ;
        RECT 443.400 433.050 444.450 443.400 ;
        RECT 442.950 430.950 445.050 433.050 ;
        RECT 443.400 421.050 444.450 430.950 ;
        RECT 445.950 421.950 448.050 424.050 ;
        RECT 436.950 418.950 439.050 421.050 ;
        RECT 442.950 418.950 445.050 421.050 ;
        RECT 415.950 415.950 418.050 418.050 ;
        RECT 424.950 416.100 427.050 418.200 ;
        RECT 416.400 411.900 417.450 415.950 ;
        RECT 425.400 415.350 426.600 416.100 ;
        RECT 433.950 415.950 436.050 418.050 ;
        RECT 421.950 412.950 424.050 415.050 ;
        RECT 424.950 412.950 427.050 415.050 ;
        RECT 427.950 412.950 430.050 415.050 ;
        RECT 415.950 409.800 418.050 411.900 ;
        RECT 422.400 411.000 423.600 412.650 ;
        RECT 428.400 411.900 429.600 412.650 ;
        RECT 434.400 411.900 435.450 415.950 ;
        RECT 421.950 406.950 424.050 411.000 ;
        RECT 427.950 409.800 430.050 411.900 ;
        RECT 433.950 409.800 436.050 411.900 ;
        RECT 437.400 382.050 438.450 418.950 ;
        RECT 446.400 417.600 447.450 421.950 ;
        RECT 449.400 418.050 450.450 448.950 ;
        RECT 455.400 448.350 456.600 449.100 ;
        RECT 461.400 448.350 462.600 450.600 ;
        RECT 472.950 449.100 475.050 451.200 ;
        RECT 478.950 449.100 481.050 451.200 ;
        RECT 484.950 450.000 487.050 454.050 ;
        RECT 454.950 445.950 457.050 448.050 ;
        RECT 457.950 445.950 460.050 448.050 ;
        RECT 460.950 445.950 463.050 448.050 ;
        RECT 463.950 445.950 466.050 448.050 ;
        RECT 458.400 444.900 459.600 445.650 ;
        RECT 457.950 442.800 460.050 444.900 ;
        RECT 464.400 443.400 465.600 445.650 ;
        RECT 473.400 445.050 474.450 449.100 ;
        RECT 479.400 448.350 480.600 449.100 ;
        RECT 485.400 448.350 486.600 450.000 ;
        RECT 478.950 445.950 481.050 448.050 ;
        RECT 481.950 445.950 484.050 448.050 ;
        RECT 484.950 445.950 487.050 448.050 ;
        RECT 487.950 445.950 490.050 448.050 ;
        RECT 464.400 439.050 465.450 443.400 ;
        RECT 472.950 442.950 475.050 445.050 ;
        RECT 482.400 443.400 483.600 445.650 ;
        RECT 488.400 443.400 489.600 445.650 ;
        RECT 463.950 436.950 466.050 439.050 ;
        RECT 457.350 423.300 459.450 425.400 ;
        RECT 446.400 415.350 447.600 417.600 ;
        RECT 448.950 417.450 451.050 418.050 ;
        RECT 452.400 417.450 453.600 417.600 ;
        RECT 448.950 416.400 453.600 417.450 ;
        RECT 448.950 415.950 451.050 416.400 ;
        RECT 452.400 415.350 453.600 416.400 ;
        RECT 440.100 412.950 442.200 415.050 ;
        RECT 445.500 412.950 447.600 415.050 ;
        RECT 451.950 412.950 454.050 415.050 ;
        RECT 440.400 410.400 441.600 412.650 ;
        RECT 458.250 410.400 459.450 423.300 ;
        RECT 440.400 394.050 441.450 410.400 ;
        RECT 457.350 408.300 459.450 410.400 ;
        RECT 458.250 401.700 459.450 408.300 ;
        RECT 464.400 406.050 465.450 436.950 ;
        RECT 475.050 423.300 477.150 425.400 ;
        RECT 469.800 412.950 471.900 415.050 ;
        RECT 470.400 411.900 471.600 412.650 ;
        RECT 469.950 409.800 472.050 411.900 ;
        RECT 463.950 403.950 466.050 406.050 ;
        RECT 475.650 404.700 476.850 423.300 ;
        RECT 482.400 418.050 483.450 443.400 ;
        RECT 488.400 439.050 489.450 443.400 ;
        RECT 487.950 436.950 490.050 439.050 ;
        RECT 494.400 420.450 495.450 478.950 ;
        RECT 496.950 466.950 499.050 469.050 ;
        RECT 497.400 442.050 498.450 466.950 ;
        RECT 509.400 457.050 510.450 496.950 ;
        RECT 517.950 494.100 520.050 496.200 ;
        RECT 523.950 494.100 526.050 496.200 ;
        RECT 518.400 493.350 519.600 494.100 ;
        RECT 524.400 493.350 525.600 494.100 ;
        RECT 514.950 490.950 517.050 493.050 ;
        RECT 517.950 490.950 520.050 493.050 ;
        RECT 520.950 490.950 523.050 493.050 ;
        RECT 523.950 490.950 526.050 493.050 ;
        RECT 515.400 488.400 516.600 490.650 ;
        RECT 521.400 488.400 522.600 490.650 ;
        RECT 515.400 484.050 516.450 488.400 ;
        RECT 514.950 481.950 517.050 484.050 ;
        RECT 514.950 475.950 517.050 478.050 ;
        RECT 508.950 454.950 511.050 457.050 ;
        RECT 507.000 453.900 510.000 454.050 ;
        RECT 507.000 453.450 511.050 453.900 ;
        RECT 506.400 451.950 511.050 453.450 ;
        RECT 506.400 450.600 507.450 451.950 ;
        RECT 508.950 451.800 511.050 451.950 ;
        RECT 506.400 448.350 507.600 450.600 ;
        RECT 502.950 445.950 505.050 448.050 ;
        RECT 505.950 445.950 508.050 448.050 ;
        RECT 508.950 445.950 511.050 448.050 ;
        RECT 503.400 443.400 504.600 445.650 ;
        RECT 509.400 444.900 510.600 445.650 ;
        RECT 503.400 442.050 504.450 443.400 ;
        RECT 508.950 442.800 511.050 444.900 ;
        RECT 496.950 439.950 499.050 442.050 ;
        RECT 502.950 439.950 505.050 442.050 ;
        RECT 499.950 421.950 502.050 424.050 ;
        RECT 491.400 419.400 495.450 420.450 ;
        RECT 481.950 415.950 484.050 418.050 ;
        RECT 478.950 412.950 481.050 415.050 ;
        RECT 479.400 411.900 480.600 412.650 ;
        RECT 491.400 411.900 492.450 419.400 ;
        RECT 500.400 417.600 501.450 421.950 ;
        RECT 500.400 415.350 501.600 417.600 ;
        RECT 503.400 417.450 504.450 439.950 ;
        RECT 511.350 423.300 513.450 425.400 ;
        RECT 506.400 417.450 507.600 417.600 ;
        RECT 503.400 416.400 507.600 417.450 ;
        RECT 506.400 415.350 507.600 416.400 ;
        RECT 494.100 412.950 496.200 415.050 ;
        RECT 499.500 412.950 501.600 415.050 ;
        RECT 505.950 412.950 508.050 415.050 ;
        RECT 478.950 409.800 481.050 411.900 ;
        RECT 490.950 409.800 493.050 411.900 ;
        RECT 494.400 410.400 495.600 412.650 ;
        RECT 512.250 410.400 513.450 423.300 ;
        RECT 472.650 403.500 476.850 404.700 ;
        RECT 472.650 402.600 474.750 403.500 ;
        RECT 457.350 399.600 459.450 401.700 ;
        RECT 479.400 397.050 480.450 409.800 ;
        RECT 454.950 394.950 457.050 397.050 ;
        RECT 478.950 394.950 481.050 397.050 ;
        RECT 439.950 391.950 442.050 394.050 ;
        RECT 391.950 376.950 394.050 379.050 ;
        RECT 397.950 376.950 400.050 379.050 ;
        RECT 403.950 376.950 406.050 379.050 ;
        RECT 412.950 376.950 415.050 379.050 ;
        RECT 427.950 376.950 430.050 379.050 ;
        RECT 436.950 376.950 439.050 382.050 ;
        RECT 445.950 379.950 448.050 382.050 ;
        RECT 368.400 370.350 369.600 372.600 ;
        RECT 376.950 371.100 379.050 373.200 ;
        RECT 382.950 371.100 385.050 373.200 ;
        RECT 388.950 371.100 391.050 373.200 ;
        RECT 367.950 367.950 370.050 370.050 ;
        RECT 377.400 361.050 378.450 371.100 ;
        RECT 383.400 370.350 384.600 371.100 ;
        RECT 389.400 370.350 390.600 371.100 ;
        RECT 382.950 367.950 385.050 370.050 ;
        RECT 385.950 367.950 388.050 370.050 ;
        RECT 388.950 367.950 391.050 370.050 ;
        RECT 391.950 367.950 394.050 370.050 ;
        RECT 386.400 366.900 387.600 367.650 ;
        RECT 392.400 366.900 393.600 367.650 ;
        RECT 398.400 366.900 399.450 376.950 ;
        RECT 404.400 372.600 405.450 376.950 ;
        RECT 428.400 372.600 429.450 376.950 ;
        RECT 446.400 376.050 447.450 379.950 ;
        RECT 445.950 373.950 448.050 376.050 ;
        RECT 404.400 370.350 405.600 372.600 ;
        RECT 428.400 370.350 429.600 372.600 ;
        RECT 439.950 371.100 442.050 373.200 ;
        RECT 446.400 372.600 447.450 373.950 ;
        RECT 455.400 372.600 456.450 394.950 ;
        RECT 472.950 388.950 475.050 391.050 ;
        RECT 461.250 379.500 463.350 380.400 ;
        RECT 459.150 378.300 463.350 379.500 ;
        RECT 440.400 370.350 441.600 371.100 ;
        RECT 446.400 370.350 447.600 372.600 ;
        RECT 455.400 370.350 456.600 372.600 ;
        RECT 403.950 367.950 406.050 370.050 ;
        RECT 406.950 367.950 409.050 370.050 ;
        RECT 409.950 367.950 412.050 370.050 ;
        RECT 421.950 367.950 424.050 370.050 ;
        RECT 424.950 367.950 427.050 370.050 ;
        RECT 427.950 367.950 430.050 370.050 ;
        RECT 439.950 367.950 442.050 370.050 ;
        RECT 442.950 367.950 445.050 370.050 ;
        RECT 445.950 367.950 448.050 370.050 ;
        RECT 448.950 367.950 451.050 370.050 ;
        RECT 454.950 367.950 457.050 370.050 ;
        RECT 385.950 364.800 388.050 366.900 ;
        RECT 391.950 364.800 394.050 366.900 ;
        RECT 397.950 364.800 400.050 366.900 ;
        RECT 407.400 365.400 408.600 367.650 ;
        RECT 425.400 366.900 426.600 367.650 ;
        RECT 407.400 361.050 408.450 365.400 ;
        RECT 424.950 364.800 427.050 366.900 ;
        RECT 433.950 364.950 436.050 367.050 ;
        RECT 443.400 366.000 444.600 367.650 ;
        RECT 349.950 355.950 352.050 358.050 ;
        RECT 355.950 355.950 358.050 358.050 ;
        RECT 364.050 357.600 366.150 359.700 ;
        RECT 376.950 358.950 379.050 361.050 ;
        RECT 406.950 358.950 409.050 361.050 ;
        RECT 349.950 349.950 352.050 352.050 ;
        RECT 340.950 346.950 343.050 349.050 ;
        RECT 341.400 339.600 342.450 346.950 ;
        RECT 335.400 337.350 336.600 339.600 ;
        RECT 341.400 337.350 342.600 339.600 ;
        RECT 350.400 337.050 351.450 349.950 ;
        RECT 356.400 339.600 357.450 355.950 ;
        RECT 388.950 352.950 391.050 355.050 ;
        RECT 361.950 343.950 364.050 346.050 ;
        RECT 362.400 339.600 363.450 343.950 ;
        RECT 389.400 340.200 390.450 352.950 ;
        RECT 430.950 349.950 433.050 352.050 ;
        RECT 394.350 345.300 396.450 347.400 ;
        RECT 356.400 337.350 357.600 339.600 ;
        RECT 362.400 337.350 363.600 339.600 ;
        RECT 370.950 337.950 373.050 340.050 ;
        RECT 379.950 338.100 382.050 340.200 ;
        RECT 388.950 338.100 391.050 340.200 ;
        RECT 334.950 334.950 337.050 337.050 ;
        RECT 337.950 334.950 340.050 337.050 ;
        RECT 340.950 334.950 343.050 337.050 ;
        RECT 343.950 334.950 346.050 337.050 ;
        RECT 349.950 334.950 352.050 337.050 ;
        RECT 355.950 334.950 358.050 337.050 ;
        RECT 358.950 334.950 361.050 337.050 ;
        RECT 361.950 334.950 364.050 337.050 ;
        RECT 364.950 334.950 367.050 337.050 ;
        RECT 328.950 331.800 331.050 333.900 ;
        RECT 338.400 332.400 339.600 334.650 ;
        RECT 344.400 332.400 345.600 334.650 ;
        RECT 325.950 328.950 328.050 331.050 ;
        RECT 313.950 325.950 316.050 328.050 ;
        RECT 326.400 322.050 327.450 328.950 ;
        RECT 325.950 319.950 328.050 322.050 ;
        RECT 316.950 316.950 319.050 319.050 ;
        RECT 310.950 298.950 313.050 301.050 ;
        RECT 311.400 294.600 312.450 298.950 ;
        RECT 317.400 297.450 318.450 316.950 ;
        RECT 319.950 310.950 322.050 313.050 ;
        RECT 320.400 307.050 321.450 310.950 ;
        RECT 329.400 307.050 330.450 331.800 ;
        RECT 338.400 325.050 339.450 332.400 ;
        RECT 337.950 324.450 340.050 325.050 ;
        RECT 337.950 323.400 342.450 324.450 ;
        RECT 337.950 322.950 340.050 323.400 ;
        RECT 319.950 304.950 322.050 307.050 ;
        RECT 328.950 304.950 331.050 307.050 ;
        RECT 334.950 304.950 337.050 307.050 ;
        RECT 317.400 296.400 321.450 297.450 ;
        RECT 311.400 292.350 312.600 294.600 ;
        RECT 311.100 289.950 313.200 292.050 ;
        RECT 316.500 289.950 318.600 292.050 ;
        RECT 320.400 268.050 321.450 296.400 ;
        RECT 335.400 294.600 336.450 304.950 ;
        RECT 335.400 292.350 336.600 294.600 ;
        RECT 328.950 289.950 331.050 292.050 ;
        RECT 331.950 289.950 334.050 292.050 ;
        RECT 334.950 289.950 337.050 292.050 ;
        RECT 332.400 288.900 333.600 289.650 ;
        RECT 331.950 286.800 334.050 288.900 ;
        RECT 319.950 265.950 322.050 268.050 ;
        RECT 325.950 265.950 328.050 268.050 ;
        RECT 311.100 256.950 313.200 259.050 ;
        RECT 316.500 256.950 318.600 259.050 ;
        RECT 319.800 256.950 321.900 259.050 ;
        RECT 311.400 254.400 312.600 256.650 ;
        RECT 320.400 255.900 321.600 256.650 ;
        RECT 326.400 256.050 327.450 265.950 ;
        RECT 332.400 261.450 333.450 286.800 ;
        RECT 334.950 277.950 337.050 280.050 ;
        RECT 329.400 260.400 333.450 261.450 ;
        RECT 335.400 261.600 336.450 277.950 ;
        RECT 341.400 270.450 342.450 323.400 ;
        RECT 344.400 295.050 345.450 332.400 ;
        RECT 346.950 331.950 349.050 334.050 ;
        RECT 352.950 331.950 355.050 334.050 ;
        RECT 359.400 332.400 360.600 334.650 ;
        RECT 365.400 333.900 366.600 334.650 ;
        RECT 371.400 333.900 372.450 337.950 ;
        RECT 380.400 337.350 381.600 338.100 ;
        RECT 389.400 337.350 390.600 338.100 ;
        RECT 376.950 334.950 379.050 337.050 ;
        RECT 379.950 334.950 382.050 337.050 ;
        RECT 382.950 334.950 385.050 337.050 ;
        RECT 388.950 334.950 391.050 337.050 ;
        RECT 343.950 292.950 346.050 295.050 ;
        RECT 347.400 294.600 348.450 331.950 ;
        RECT 353.400 294.600 354.450 331.950 ;
        RECT 359.400 313.050 360.450 332.400 ;
        RECT 364.950 331.800 367.050 333.900 ;
        RECT 370.950 331.800 373.050 333.900 ;
        RECT 377.400 332.400 378.600 334.650 ;
        RECT 395.250 332.400 396.450 345.300 ;
        RECT 400.950 343.950 403.050 346.050 ;
        RECT 412.050 345.300 414.150 347.400 ;
        RECT 397.950 337.950 400.050 340.050 ;
        RECT 377.400 322.050 378.450 332.400 ;
        RECT 394.350 330.300 396.450 332.400 ;
        RECT 388.950 325.950 391.050 328.050 ;
        RECT 361.950 319.950 364.050 322.050 ;
        RECT 376.950 319.950 379.050 322.050 ;
        RECT 358.950 310.950 361.050 313.050 ;
        RECT 347.400 292.350 348.600 294.600 ;
        RECT 353.400 292.350 354.600 294.600 ;
        RECT 346.950 289.950 349.050 292.050 ;
        RECT 349.950 289.950 352.050 292.050 ;
        RECT 352.950 289.950 355.050 292.050 ;
        RECT 355.950 289.950 358.050 292.050 ;
        RECT 350.400 287.400 351.600 289.650 ;
        RECT 356.400 288.900 357.600 289.650 ;
        RECT 362.400 288.900 363.450 319.950 ;
        RECT 382.950 316.950 385.050 319.050 ;
        RECT 383.400 313.050 384.450 316.950 ;
        RECT 382.950 310.950 385.050 313.050 ;
        RECT 367.950 304.950 370.050 307.050 ;
        RECT 368.400 294.600 369.450 304.950 ;
        RECT 389.400 294.600 390.450 325.950 ;
        RECT 395.250 323.700 396.450 330.300 ;
        RECT 394.350 321.600 396.450 323.700 ;
        RECT 398.400 298.050 399.450 337.950 ;
        RECT 401.400 333.900 402.450 343.950 ;
        RECT 406.800 334.950 408.900 337.050 ;
        RECT 407.400 333.900 408.600 334.650 ;
        RECT 400.950 331.800 403.050 333.900 ;
        RECT 406.950 331.800 409.050 333.900 ;
        RECT 412.650 326.700 413.850 345.300 ;
        RECT 421.950 340.950 424.050 343.050 ;
        RECT 415.950 334.950 418.050 337.050 ;
        RECT 409.650 325.500 413.850 326.700 ;
        RECT 416.400 332.400 417.600 334.650 ;
        RECT 400.950 322.950 403.050 325.050 ;
        RECT 409.650 324.600 411.750 325.500 ;
        RECT 397.950 295.950 400.050 298.050 ;
        RECT 368.400 292.350 369.600 294.600 ;
        RECT 389.400 292.350 390.600 294.600 ;
        RECT 394.950 293.100 397.050 295.200 ;
        RECT 395.400 292.350 396.600 293.100 ;
        RECT 367.950 289.950 370.050 292.050 ;
        RECT 370.950 289.950 373.050 292.050 ;
        RECT 373.950 289.950 376.050 292.050 ;
        RECT 385.950 289.950 388.050 292.050 ;
        RECT 388.950 289.950 391.050 292.050 ;
        RECT 391.950 289.950 394.050 292.050 ;
        RECT 394.950 289.950 397.050 292.050 ;
        RECT 346.950 283.950 349.050 286.050 ;
        RECT 338.400 269.400 342.450 270.450 ;
        RECT 338.400 265.050 339.450 269.400 ;
        RECT 340.950 265.950 343.050 268.050 ;
        RECT 337.950 262.950 340.050 265.050 ;
        RECT 341.400 261.600 342.450 265.950 ;
        RECT 347.400 262.050 348.450 283.950 ;
        RECT 350.400 280.050 351.450 287.400 ;
        RECT 355.950 286.800 358.050 288.900 ;
        RECT 361.950 286.800 364.050 288.900 ;
        RECT 371.400 287.400 372.600 289.650 ;
        RECT 386.400 288.900 387.600 289.650 ;
        RECT 349.950 277.950 352.050 280.050 ;
        RECT 364.950 277.950 367.050 280.050 ;
        RECT 352.950 268.950 355.050 271.050 ;
        RECT 353.400 262.050 354.450 268.950 ;
        RECT 307.950 247.950 310.050 250.050 ;
        RECT 301.950 241.950 304.050 244.050 ;
        RECT 311.400 238.050 312.450 254.400 ;
        RECT 319.950 253.800 322.050 255.900 ;
        RECT 325.950 253.950 328.050 256.050 ;
        RECT 325.950 241.950 328.050 244.050 ;
        RECT 310.950 235.950 313.050 238.050 ;
        RECT 316.950 232.950 319.050 235.050 ;
        RECT 304.950 223.800 307.050 225.900 ;
        RECT 305.400 216.600 306.450 223.800 ;
        RECT 305.400 214.350 306.600 216.600 ;
        RECT 310.950 215.100 313.050 217.200 ;
        RECT 317.400 217.050 318.450 232.950 ;
        RECT 319.950 217.950 322.050 220.050 ;
        RECT 311.400 214.350 312.600 215.100 ;
        RECT 316.950 214.950 319.050 217.050 ;
        RECT 304.950 211.950 307.050 214.050 ;
        RECT 307.950 211.950 310.050 214.050 ;
        RECT 310.950 211.950 313.050 214.050 ;
        RECT 313.950 211.950 316.050 214.050 ;
        RECT 301.950 208.950 304.050 211.050 ;
        RECT 308.400 209.400 309.600 211.650 ;
        RECT 314.400 210.450 315.600 211.650 ;
        RECT 314.400 209.400 318.450 210.450 ;
        RECT 298.950 205.950 301.050 208.050 ;
        RECT 293.400 182.400 297.450 183.450 ;
        RECT 293.400 181.350 294.600 182.400 ;
        RECT 285.000 179.700 291.900 180.900 ;
        RECT 285.000 177.300 285.900 179.700 ;
        RECT 283.800 175.200 285.900 177.300 ;
        RECT 286.800 175.950 288.900 178.050 ;
        RECT 280.500 171.600 282.600 173.700 ;
        RECT 287.400 173.400 288.600 175.650 ;
        RECT 290.700 172.500 291.900 179.700 ;
        RECT 292.800 178.950 294.900 181.050 ;
        RECT 290.100 170.400 292.200 172.500 ;
        RECT 283.950 166.950 286.050 169.050 ;
        RECT 277.950 145.950 280.050 148.050 ;
        RECT 278.400 138.600 279.450 145.950 ;
        RECT 284.400 138.600 285.450 166.950 ;
        RECT 302.400 163.050 303.450 208.950 ;
        RECT 308.400 199.050 309.450 209.400 ;
        RECT 307.950 196.950 310.050 199.050 ;
        RECT 313.950 196.950 316.050 199.050 ;
        RECT 314.400 187.050 315.450 196.950 ;
        RECT 317.400 196.050 318.450 209.400 ;
        RECT 320.400 202.050 321.450 217.950 ;
        RECT 326.400 216.600 327.450 241.950 ;
        RECT 329.400 220.050 330.450 260.400 ;
        RECT 335.400 259.350 336.600 261.600 ;
        RECT 341.400 259.350 342.600 261.600 ;
        RECT 346.950 259.950 349.050 262.050 ;
        RECT 352.950 259.950 355.050 262.050 ;
        RECT 358.950 260.100 361.050 262.200 ;
        RECT 365.400 262.050 366.450 277.950 ;
        RECT 371.400 274.050 372.450 287.400 ;
        RECT 385.950 286.800 388.050 288.900 ;
        RECT 392.400 287.400 393.600 289.650 ;
        RECT 392.400 283.050 393.450 287.400 ;
        RECT 385.950 280.950 388.050 283.050 ;
        RECT 391.950 280.950 394.050 283.050 ;
        RECT 370.950 271.950 373.050 274.050 ;
        RECT 376.950 271.950 379.050 274.050 ;
        RECT 377.400 262.200 378.450 271.950 ;
        RECT 359.400 259.350 360.600 260.100 ;
        RECT 364.950 259.950 367.050 262.050 ;
        RECT 367.950 259.950 370.050 262.050 ;
        RECT 376.950 260.100 379.050 262.200 ;
        RECT 386.400 262.050 387.450 280.950 ;
        RECT 391.950 265.950 394.050 268.050 ;
        RECT 334.950 256.950 337.050 259.050 ;
        RECT 337.950 256.950 340.050 259.050 ;
        RECT 340.950 256.950 343.050 259.050 ;
        RECT 343.950 256.950 346.050 259.050 ;
        RECT 355.950 256.950 358.050 259.050 ;
        RECT 358.950 256.950 361.050 259.050 ;
        RECT 361.950 256.950 364.050 259.050 ;
        RECT 338.400 255.900 339.600 256.650 ;
        RECT 344.400 255.900 345.600 256.650 ;
        RECT 337.950 253.800 340.050 255.900 ;
        RECT 343.950 253.800 346.050 255.900 ;
        RECT 356.400 255.450 357.600 256.650 ;
        RECT 362.400 255.900 363.600 256.650 ;
        RECT 353.400 254.400 357.600 255.450 ;
        RECT 343.950 250.650 346.050 252.750 ;
        RECT 328.950 217.950 331.050 220.050 ;
        RECT 326.400 214.350 327.600 216.600 ;
        RECT 331.950 215.100 334.050 217.200 ;
        RECT 344.400 217.050 345.450 250.650 ;
        RECT 353.400 247.050 354.450 254.400 ;
        RECT 361.950 253.800 364.050 255.900 ;
        RECT 364.950 253.950 367.050 256.050 ;
        RECT 355.950 250.950 358.050 253.050 ;
        RECT 352.950 244.950 355.050 247.050 ;
        RECT 353.400 241.050 354.450 244.950 ;
        RECT 352.950 238.950 355.050 241.050 ;
        RECT 332.400 214.350 333.600 215.100 ;
        RECT 343.950 214.950 346.050 217.050 ;
        RECT 353.400 216.450 354.600 216.600 ;
        RECT 356.400 216.450 357.450 250.950 ;
        RECT 358.950 220.950 361.050 223.050 ;
        RECT 353.400 215.400 357.450 216.450 ;
        RECT 353.400 214.350 354.600 215.400 ;
        RECT 325.950 211.950 328.050 214.050 ;
        RECT 328.950 211.950 331.050 214.050 ;
        RECT 331.950 211.950 334.050 214.050 ;
        RECT 334.950 211.950 337.050 214.050 ;
        RECT 346.950 211.950 349.050 214.050 ;
        RECT 349.950 211.950 352.050 214.050 ;
        RECT 352.950 211.950 355.050 214.050 ;
        RECT 322.950 208.950 325.050 211.050 ;
        RECT 329.400 209.400 330.600 211.650 ;
        RECT 335.400 209.400 336.600 211.650 ;
        RECT 350.400 210.900 351.600 211.650 ;
        RECT 319.950 199.950 322.050 202.050 ;
        RECT 316.950 193.950 319.050 196.050 ;
        RECT 316.950 187.950 319.050 190.050 ;
        RECT 307.950 183.000 310.050 187.050 ;
        RECT 313.950 184.950 316.050 187.050 ;
        RECT 308.400 181.350 309.600 183.000 ;
        RECT 305.100 178.950 307.200 181.050 ;
        RECT 308.400 178.950 310.500 181.050 ;
        RECT 313.800 178.950 315.900 181.050 ;
        RECT 305.400 176.400 306.600 178.650 ;
        RECT 314.400 177.000 315.600 178.650 ;
        RECT 301.950 160.950 304.050 163.050 ;
        RECT 289.950 145.950 292.050 148.050 ;
        RECT 278.400 136.350 279.600 138.600 ;
        RECT 284.400 136.350 285.600 138.600 ;
        RECT 277.950 133.950 280.050 136.050 ;
        RECT 280.950 133.950 283.050 136.050 ;
        RECT 283.950 133.950 286.050 136.050 ;
        RECT 281.400 131.400 282.600 133.650 ;
        RECT 290.400 132.900 291.450 145.950 ;
        RECT 305.400 145.050 306.450 176.400 ;
        RECT 313.950 172.950 316.050 177.000 ;
        RECT 310.950 162.450 315.000 163.050 ;
        RECT 310.950 160.950 315.450 162.450 ;
        RECT 310.950 154.950 313.050 157.050 ;
        RECT 304.950 142.950 307.050 145.050 ;
        RECT 295.950 137.100 298.050 139.200 ;
        RECT 301.950 137.100 304.050 139.200 ;
        RECT 296.400 136.350 297.600 137.100 ;
        RECT 302.400 136.350 303.600 137.100 ;
        RECT 295.950 133.950 298.050 136.050 ;
        RECT 298.950 133.950 301.050 136.050 ;
        RECT 301.950 133.950 304.050 136.050 ;
        RECT 304.950 133.950 307.050 136.050 ;
        RECT 299.400 132.900 300.600 133.650 ;
        RECT 277.950 127.950 280.050 130.050 ;
        RECT 274.950 118.950 277.050 121.050 ;
        RECT 275.400 97.050 276.450 118.950 ;
        RECT 278.400 106.050 279.450 127.950 ;
        RECT 281.400 118.050 282.450 131.400 ;
        RECT 289.950 130.800 292.050 132.900 ;
        RECT 298.950 130.800 301.050 132.900 ;
        RECT 305.400 131.400 306.600 133.650 ;
        RECT 311.400 132.450 312.450 154.950 ;
        RECT 314.400 145.050 315.450 160.950 ;
        RECT 317.400 154.050 318.450 187.950 ;
        RECT 319.950 182.100 322.050 184.200 ;
        RECT 323.400 184.050 324.450 208.950 ;
        RECT 329.400 190.050 330.450 209.400 ;
        RECT 335.400 202.050 336.450 209.400 ;
        RECT 349.950 208.800 352.050 210.900 ;
        RECT 334.950 199.950 337.050 202.050 ;
        RECT 334.950 196.800 337.050 198.900 ;
        RECT 328.950 187.950 331.050 190.050 ;
        RECT 320.400 177.450 321.450 182.100 ;
        RECT 322.950 181.950 325.050 184.050 ;
        RECT 328.950 182.100 331.050 184.200 ;
        RECT 335.400 184.050 336.450 196.800 ;
        RECT 350.400 190.050 351.450 208.800 ;
        RECT 359.400 196.050 360.450 220.950 ;
        RECT 365.400 217.050 366.450 253.950 ;
        RECT 368.400 219.450 369.450 259.950 ;
        RECT 377.400 259.350 378.600 260.100 ;
        RECT 382.950 259.950 385.050 262.050 ;
        RECT 385.950 259.950 388.050 262.050 ;
        RECT 392.400 261.600 393.450 265.950 ;
        RECT 401.400 265.050 402.450 322.950 ;
        RECT 409.950 319.950 412.050 322.050 ;
        RECT 410.400 301.050 411.450 319.950 ;
        RECT 416.400 316.050 417.450 332.400 ;
        RECT 422.400 328.050 423.450 340.950 ;
        RECT 431.400 339.600 432.450 349.950 ;
        RECT 434.400 343.050 435.450 364.950 ;
        RECT 442.950 361.950 445.050 366.000 ;
        RECT 449.400 365.400 450.600 367.650 ;
        RECT 449.400 352.050 450.450 365.400 ;
        RECT 459.150 359.700 460.350 378.300 ;
        RECT 463.950 371.100 466.050 373.200 ;
        RECT 464.400 370.350 465.600 371.100 ;
        RECT 469.950 370.950 472.050 373.050 ;
        RECT 464.100 367.950 466.200 370.050 ;
        RECT 470.400 364.050 471.450 370.950 ;
        RECT 469.950 361.950 472.050 364.050 ;
        RECT 458.850 357.600 460.950 359.700 ;
        RECT 448.950 349.950 451.050 352.050 ;
        RECT 469.950 349.950 472.050 352.050 ;
        RECT 445.350 345.300 447.450 347.400 ;
        RECT 433.950 340.950 436.050 343.050 ;
        RECT 431.400 337.350 432.600 339.600 ;
        RECT 439.950 338.100 442.050 340.200 ;
        RECT 440.400 337.350 441.600 338.100 ;
        RECT 430.950 334.950 433.050 337.050 ;
        RECT 433.950 334.950 436.050 337.050 ;
        RECT 439.950 334.950 442.050 337.050 ;
        RECT 434.400 332.400 435.600 334.650 ;
        RECT 421.950 325.950 424.050 328.050 ;
        RECT 415.950 313.950 418.050 316.050 ;
        RECT 415.950 301.950 418.050 304.050 ;
        RECT 409.950 298.950 412.050 301.050 ;
        RECT 410.400 294.600 411.450 298.950 ;
        RECT 416.400 295.200 417.450 301.950 ;
        RECT 410.400 292.350 411.600 294.600 ;
        RECT 415.950 293.100 418.050 295.200 ;
        RECT 416.400 292.350 417.600 293.100 ;
        RECT 409.950 289.950 412.050 292.050 ;
        RECT 412.950 289.950 415.050 292.050 ;
        RECT 415.950 289.950 418.050 292.050 ;
        RECT 413.400 288.900 414.600 289.650 ;
        RECT 412.950 286.800 415.050 288.900 ;
        RECT 418.950 277.950 421.050 280.050 ;
        RECT 400.950 262.950 403.050 265.050 ;
        RECT 373.950 256.950 376.050 259.050 ;
        RECT 376.950 256.950 379.050 259.050 ;
        RECT 374.400 254.400 375.600 256.650 ;
        RECT 374.400 220.050 375.450 254.400 ;
        RECT 383.400 235.050 384.450 259.950 ;
        RECT 392.400 259.350 393.600 261.600 ;
        RECT 397.950 260.100 400.050 262.200 ;
        RECT 398.400 259.350 399.600 260.100 ;
        RECT 403.950 259.950 406.050 262.050 ;
        RECT 412.950 260.100 415.050 262.200 ;
        RECT 419.400 262.050 420.450 277.950 ;
        RECT 422.400 271.050 423.450 325.950 ;
        RECT 434.400 325.050 435.450 332.400 ;
        RECT 436.950 331.950 439.050 334.050 ;
        RECT 446.250 332.400 447.450 345.300 ;
        RECT 449.400 334.050 450.450 349.950 ;
        RECT 463.050 345.300 465.150 347.400 ;
        RECT 451.950 337.950 454.050 340.050 ;
        RECT 433.950 322.950 436.050 325.050 ;
        RECT 437.400 313.050 438.450 331.950 ;
        RECT 445.350 330.300 447.450 332.400 ;
        RECT 448.950 331.950 451.050 334.050 ;
        RECT 446.250 323.700 447.450 330.300 ;
        RECT 452.400 325.050 453.450 337.950 ;
        RECT 457.800 334.950 459.900 337.050 ;
        RECT 458.400 333.450 459.600 334.650 ;
        RECT 455.400 332.400 459.600 333.450 ;
        RECT 455.400 325.050 456.450 332.400 ;
        RECT 463.650 326.700 464.850 345.300 ;
        RECT 470.400 340.050 471.450 349.950 ;
        RECT 473.400 346.050 474.450 388.950 ;
        RECT 476.550 381.300 478.650 383.400 ;
        RECT 476.550 374.700 477.750 381.300 ;
        RECT 476.550 372.600 478.650 374.700 ;
        RECT 476.550 359.700 477.750 372.600 ;
        RECT 481.950 367.950 484.050 370.050 ;
        RECT 482.400 365.400 483.600 367.650 ;
        RECT 491.400 367.050 492.450 409.800 ;
        RECT 494.400 406.050 495.450 410.400 ;
        RECT 511.350 408.300 513.450 410.400 ;
        RECT 493.950 403.950 496.050 406.050 ;
        RECT 512.250 401.700 513.450 408.300 ;
        RECT 515.400 406.050 516.450 475.950 ;
        RECT 521.400 469.050 522.450 488.400 ;
        RECT 533.400 478.050 534.450 511.950 ;
        RECT 539.400 505.050 540.450 521.400 ;
        RECT 548.400 514.050 549.450 532.950 ;
        RECT 557.400 528.600 558.450 532.950 ;
        RECT 557.400 526.350 558.600 528.600 ;
        RECT 553.950 523.950 556.050 526.050 ;
        RECT 556.950 523.950 559.050 526.050 ;
        RECT 559.950 523.950 562.050 526.050 ;
        RECT 554.400 521.400 555.600 523.650 ;
        RECT 560.400 522.900 561.600 523.650 ;
        RECT 547.950 511.950 550.050 514.050 ;
        RECT 538.950 502.950 541.050 505.050 ;
        RECT 535.950 499.950 538.050 502.050 ;
        RECT 532.950 475.950 535.050 478.050 ;
        RECT 520.950 466.950 523.050 469.050 ;
        RECT 521.400 463.050 522.450 466.950 ;
        RECT 520.950 460.950 523.050 463.050 ;
        RECT 520.950 449.100 523.050 451.200 ;
        RECT 526.950 450.000 529.050 454.050 ;
        RECT 521.400 448.350 522.600 449.100 ;
        RECT 527.400 448.350 528.600 450.000 ;
        RECT 520.950 445.950 523.050 448.050 ;
        RECT 523.950 445.950 526.050 448.050 ;
        RECT 526.950 445.950 529.050 448.050 ;
        RECT 529.950 445.950 532.050 448.050 ;
        RECT 524.400 444.000 525.600 445.650 ;
        RECT 523.950 439.950 526.050 444.000 ;
        RECT 530.400 443.400 531.600 445.650 ;
        RECT 530.400 430.050 531.450 443.400 ;
        RECT 536.400 442.050 537.450 499.950 ;
        RECT 544.950 494.100 547.050 496.200 ;
        RECT 539.100 490.950 541.200 493.050 ;
        RECT 539.400 488.400 540.600 490.650 ;
        RECT 539.400 481.050 540.450 488.400 ;
        RECT 538.950 478.950 541.050 481.050 ;
        RECT 538.950 472.950 541.050 475.050 ;
        RECT 535.950 439.950 538.050 442.050 ;
        RECT 517.950 427.950 520.050 430.050 ;
        RECT 529.950 427.950 532.050 430.050 ;
        RECT 518.400 411.900 519.450 427.950 ;
        RECT 529.050 423.300 531.150 425.400 ;
        RECT 523.800 412.950 525.900 415.050 ;
        RECT 524.400 411.900 525.600 412.650 ;
        RECT 517.950 409.800 520.050 411.900 ;
        RECT 523.950 409.800 526.050 411.900 ;
        RECT 514.950 403.950 517.050 406.050 ;
        RECT 520.950 403.950 523.050 406.050 ;
        RECT 529.650 404.700 530.850 423.300 ;
        RECT 532.950 412.950 535.050 415.050 ;
        RECT 533.400 411.900 534.600 412.650 ;
        RECT 532.950 409.800 535.050 411.900 ;
        RECT 539.400 408.450 540.450 472.950 ;
        RECT 541.950 454.950 544.050 457.050 ;
        RECT 536.400 407.400 540.450 408.450 ;
        RECT 511.350 399.600 513.450 401.700 ;
        RECT 521.400 391.050 522.450 403.950 ;
        RECT 526.650 403.500 530.850 404.700 ;
        RECT 532.950 403.950 535.050 406.050 ;
        RECT 526.650 402.600 528.750 403.500 ;
        RECT 529.950 397.950 532.050 400.050 ;
        RECT 520.950 388.950 523.050 391.050 ;
        RECT 521.400 376.050 522.450 388.950 ;
        RECT 526.950 376.950 529.050 379.050 ;
        RECT 502.950 372.000 505.050 376.050 ;
        RECT 503.400 370.350 504.600 372.000 ;
        RECT 508.950 371.100 511.050 373.200 ;
        RECT 514.950 371.100 517.050 373.200 ;
        RECT 520.950 372.000 523.050 376.050 ;
        RECT 527.400 373.050 528.450 376.950 ;
        RECT 496.950 367.950 499.050 370.050 ;
        RECT 499.950 367.950 502.050 370.050 ;
        RECT 502.950 367.950 505.050 370.050 ;
        RECT 476.550 357.600 478.650 359.700 ;
        RECT 482.400 352.050 483.450 365.400 ;
        RECT 484.950 364.950 487.050 367.050 ;
        RECT 490.950 364.950 493.050 367.050 ;
        RECT 500.400 366.000 501.600 367.650 ;
        RECT 481.950 349.950 484.050 352.050 ;
        RECT 472.950 343.950 475.050 346.050 ;
        RECT 481.350 345.300 483.450 347.400 ;
        RECT 469.950 337.950 472.050 340.050 ;
        RECT 475.950 338.100 478.050 340.200 ;
        RECT 476.400 337.350 477.600 338.100 ;
        RECT 466.950 334.950 469.050 337.050 ;
        RECT 475.950 334.950 478.050 337.050 ;
        RECT 467.400 333.000 468.600 334.650 ;
        RECT 466.950 328.950 469.050 333.000 ;
        RECT 469.950 331.950 472.050 334.050 ;
        RECT 482.250 332.400 483.450 345.300 ;
        RECT 460.650 325.500 464.850 326.700 ;
        RECT 445.350 321.600 447.450 323.700 ;
        RECT 451.800 322.950 453.900 325.050 ;
        RECT 454.950 322.950 457.050 325.050 ;
        RECT 460.650 324.600 462.750 325.500 ;
        RECT 467.400 316.050 468.450 328.950 ;
        RECT 466.950 313.950 469.050 316.050 ;
        RECT 470.400 313.050 471.450 331.950 ;
        RECT 481.350 330.300 483.450 332.400 ;
        RECT 485.400 331.050 486.450 364.950 ;
        RECT 499.950 361.950 502.050 366.000 ;
        RECT 509.400 364.050 510.450 371.100 ;
        RECT 515.400 370.350 516.600 371.100 ;
        RECT 521.400 370.350 522.600 372.000 ;
        RECT 526.950 370.950 529.050 373.050 ;
        RECT 514.950 367.950 517.050 370.050 ;
        RECT 517.950 367.950 520.050 370.050 ;
        RECT 520.950 367.950 523.050 370.050 ;
        RECT 523.950 367.950 526.050 370.050 ;
        RECT 518.400 365.400 519.600 367.650 ;
        RECT 524.400 366.900 525.600 367.650 ;
        RECT 508.950 361.950 511.050 364.050 ;
        RECT 518.400 361.050 519.450 365.400 ;
        RECT 523.950 364.800 526.050 366.900 ;
        RECT 526.950 363.450 529.050 367.050 ;
        RECT 524.400 363.000 529.050 363.450 ;
        RECT 524.400 362.400 528.450 363.000 ;
        RECT 505.950 358.950 508.050 361.050 ;
        RECT 517.950 358.950 520.050 361.050 ;
        RECT 487.950 349.950 490.050 352.050 ;
        RECT 482.250 323.700 483.450 330.300 ;
        RECT 484.950 328.950 487.050 331.050 ;
        RECT 481.350 321.600 483.450 323.700 ;
        RECT 472.950 313.950 475.050 316.050 ;
        RECT 436.950 310.950 439.050 313.050 ;
        RECT 469.950 310.950 472.050 313.050 ;
        RECT 433.950 306.450 436.050 307.050 ;
        RECT 437.400 306.450 438.450 310.950 ;
        RECT 457.950 307.950 460.050 310.050 ;
        RECT 433.950 305.400 438.450 306.450 ;
        RECT 433.950 304.950 436.050 305.400 ;
        RECT 434.400 294.600 435.450 304.950 ;
        RECT 445.950 303.450 448.050 304.050 ;
        RECT 443.400 302.400 448.050 303.450 ;
        RECT 434.400 292.350 435.600 294.600 ;
        RECT 430.950 289.950 433.050 292.050 ;
        RECT 433.950 289.950 436.050 292.050 ;
        RECT 431.400 288.900 432.600 289.650 ;
        RECT 430.950 286.800 433.050 288.900 ;
        RECT 443.400 277.050 444.450 302.400 ;
        RECT 445.950 300.450 448.050 302.400 ;
        RECT 445.950 300.000 450.450 300.450 ;
        RECT 446.400 299.400 450.450 300.000 ;
        RECT 449.400 294.600 450.450 299.400 ;
        RECT 458.400 295.050 459.450 307.950 ;
        RECT 473.400 307.050 474.450 313.950 ;
        RECT 472.800 304.950 474.900 307.050 ;
        RECT 475.950 304.950 478.050 307.050 ;
        RECT 485.400 306.450 486.450 328.950 ;
        RECT 488.400 307.050 489.450 349.950 ;
        RECT 499.050 345.300 501.150 347.400 ;
        RECT 493.800 334.950 495.900 337.050 ;
        RECT 490.800 331.950 492.900 334.050 ;
        RECT 494.400 333.900 495.600 334.650 ;
        RECT 491.400 321.450 492.450 331.950 ;
        RECT 493.950 331.800 496.050 333.900 ;
        RECT 499.650 326.700 500.850 345.300 ;
        RECT 506.400 340.050 507.450 358.950 ;
        RECT 511.950 355.950 514.050 358.050 ;
        RECT 508.950 343.950 511.050 346.050 ;
        RECT 505.950 337.950 508.050 340.050 ;
        RECT 502.950 334.950 505.050 337.050 ;
        RECT 503.400 332.400 504.600 334.650 ;
        RECT 503.400 328.050 504.450 332.400 ;
        RECT 509.400 331.050 510.450 343.950 ;
        RECT 512.400 333.450 513.450 355.950 ;
        RECT 517.950 338.100 520.050 340.200 ;
        RECT 524.400 339.600 525.450 362.400 ;
        RECT 526.950 358.950 529.050 361.050 ;
        RECT 527.400 349.050 528.450 358.950 ;
        RECT 526.950 346.950 529.050 349.050 ;
        RECT 530.400 340.050 531.450 397.950 ;
        RECT 533.400 358.050 534.450 403.950 ;
        RECT 536.400 373.050 537.450 407.400 ;
        RECT 542.400 406.050 543.450 454.950 ;
        RECT 545.400 451.200 546.450 494.100 ;
        RECT 554.400 469.050 555.450 521.400 ;
        RECT 559.950 520.800 562.050 522.900 ;
        RECT 556.950 511.950 559.050 514.050 ;
        RECT 557.400 502.050 558.450 511.950 ;
        RECT 556.950 499.950 559.050 502.050 ;
        RECT 560.400 496.050 561.450 520.800 ;
        RECT 562.950 508.950 565.050 511.050 ;
        RECT 559.950 493.950 562.050 496.050 ;
        RECT 563.400 495.450 564.450 508.950 ;
        RECT 566.400 505.050 567.450 532.950 ;
        RECT 574.950 528.000 577.050 532.050 ;
        RECT 575.400 526.350 576.600 528.000 ;
        RECT 571.950 523.950 574.050 526.050 ;
        RECT 574.950 523.950 577.050 526.050 ;
        RECT 577.950 523.950 580.050 526.050 ;
        RECT 572.400 521.400 573.600 523.650 ;
        RECT 578.400 522.900 579.600 523.650 ;
        RECT 572.400 511.050 573.450 521.400 ;
        RECT 577.950 520.800 580.050 522.900 ;
        RECT 577.950 514.950 580.050 517.050 ;
        RECT 571.950 508.950 574.050 511.050 ;
        RECT 565.950 502.950 568.050 505.050 ;
        RECT 571.350 501.300 573.450 503.400 ;
        RECT 566.400 495.450 567.600 495.600 ;
        RECT 563.400 494.400 567.600 495.450 ;
        RECT 566.400 493.350 567.600 494.400 ;
        RECT 557.100 490.950 559.200 493.050 ;
        RECT 565.950 490.950 568.050 493.050 ;
        RECT 572.250 488.400 573.450 501.300 ;
        RECT 578.400 489.900 579.450 514.950 ;
        RECT 584.400 511.050 585.450 565.950 ;
        RECT 590.400 547.050 591.450 566.400 ;
        RECT 595.950 565.800 598.050 567.900 ;
        RECT 608.250 566.400 609.450 579.300 ;
        RECT 610.950 577.950 613.050 580.050 ;
        RECT 607.350 564.300 609.450 566.400 ;
        RECT 608.250 557.700 609.450 564.300 ;
        RECT 607.350 555.600 609.450 557.700 ;
        RECT 589.950 544.950 592.050 547.050 ;
        RECT 607.950 544.950 610.050 547.050 ;
        RECT 604.950 538.950 607.050 541.050 ;
        RECT 592.950 528.000 595.050 532.050 ;
        RECT 593.400 526.350 594.600 528.000 ;
        RECT 598.950 527.100 601.050 529.200 ;
        RECT 599.400 526.350 600.600 527.100 ;
        RECT 589.950 523.950 592.050 526.050 ;
        RECT 592.950 523.950 595.050 526.050 ;
        RECT 595.950 523.950 598.050 526.050 ;
        RECT 598.950 523.950 601.050 526.050 ;
        RECT 590.400 521.400 591.600 523.650 ;
        RECT 596.400 522.000 597.600 523.650 ;
        RECT 590.400 517.050 591.450 521.400 ;
        RECT 595.950 517.950 598.050 522.000 ;
        RECT 601.950 520.950 604.050 523.050 ;
        RECT 589.950 514.950 592.050 517.050 ;
        RECT 583.950 508.950 586.050 511.050 ;
        RECT 589.050 501.300 591.150 503.400 ;
        RECT 583.800 490.950 585.900 493.050 ;
        RECT 584.400 489.900 585.600 490.650 ;
        RECT 571.350 486.300 573.450 488.400 ;
        RECT 577.950 487.800 580.050 489.900 ;
        RECT 583.950 487.800 586.050 489.900 ;
        RECT 572.250 479.700 573.450 486.300 ;
        RECT 580.950 481.950 583.050 484.050 ;
        RECT 589.650 482.700 590.850 501.300 ;
        RECT 602.400 496.050 603.450 520.950 ;
        RECT 605.400 520.050 606.450 538.950 ;
        RECT 608.400 529.050 609.450 544.950 ;
        RECT 611.400 535.050 612.450 577.950 ;
        RECT 620.400 577.050 621.450 589.950 ;
        RECT 625.050 579.300 627.150 581.400 ;
        RECT 613.950 574.950 616.050 577.050 ;
        RECT 619.950 574.950 622.050 577.050 ;
        RECT 614.400 567.900 615.450 574.950 ;
        RECT 619.800 568.950 621.900 571.050 ;
        RECT 620.400 567.900 621.600 568.650 ;
        RECT 613.950 565.800 616.050 567.900 ;
        RECT 619.950 565.800 622.050 567.900 ;
        RECT 625.650 560.700 626.850 579.300 ;
        RECT 629.400 577.050 630.450 601.950 ;
        RECT 632.550 593.700 633.750 606.600 ;
        RECT 637.950 601.950 640.050 604.050 ;
        RECT 638.400 600.900 639.600 601.650 ;
        RECT 644.400 600.900 645.450 610.950 ;
        RECT 637.950 598.800 640.050 600.900 ;
        RECT 643.950 598.800 646.050 600.900 ;
        RECT 632.550 591.600 634.650 593.700 ;
        RECT 637.950 589.950 640.050 592.050 ;
        RECT 634.950 586.950 637.050 589.050 ;
        RECT 628.950 574.950 631.050 577.050 ;
        RECT 628.950 568.950 631.050 571.050 ;
        RECT 629.400 567.900 630.600 568.650 ;
        RECT 628.950 565.800 631.050 567.900 ;
        RECT 622.650 559.500 626.850 560.700 ;
        RECT 613.950 556.950 616.050 559.050 ;
        RECT 622.650 558.600 624.750 559.500 ;
        RECT 610.950 532.950 613.050 535.050 ;
        RECT 607.950 526.950 610.050 529.050 ;
        RECT 614.400 528.600 615.450 556.950 ;
        RECT 629.400 553.050 630.450 565.800 ;
        RECT 635.400 559.050 636.450 586.950 ;
        RECT 634.950 556.950 637.050 559.050 ;
        RECT 628.800 550.950 630.900 553.050 ;
        RECT 625.950 544.950 628.050 547.050 ;
        RECT 622.950 538.950 625.050 541.050 ;
        RECT 614.400 526.350 615.600 528.600 ;
        RECT 619.950 527.100 622.050 529.200 ;
        RECT 623.400 528.450 624.450 538.950 ;
        RECT 626.400 538.050 627.450 544.950 ;
        RECT 629.400 541.050 630.450 550.950 ;
        RECT 635.400 541.050 636.450 556.950 ;
        RECT 638.400 556.050 639.450 589.950 ;
        RECT 647.400 577.050 648.450 619.950 ;
        RECT 673.950 616.950 676.050 619.050 ;
        RECT 670.950 613.950 673.050 616.050 ;
        RECT 652.950 610.950 655.050 613.050 ;
        RECT 653.400 606.600 654.450 610.950 ;
        RECT 664.950 607.950 667.050 610.050 ;
        RECT 653.400 604.350 654.600 606.600 ;
        RECT 658.950 605.100 661.050 607.200 ;
        RECT 659.400 604.350 660.600 605.100 ;
        RECT 652.950 601.950 655.050 604.050 ;
        RECT 655.950 601.950 658.050 604.050 ;
        RECT 658.950 601.950 661.050 604.050 ;
        RECT 656.400 600.900 657.600 601.650 ;
        RECT 665.400 601.050 666.450 607.950 ;
        RECT 671.400 606.600 672.450 613.950 ;
        RECT 674.400 610.050 675.450 616.950 ;
        RECT 686.400 616.050 687.450 644.400 ;
        RECT 689.400 628.050 690.450 667.950 ;
        RECT 695.400 663.450 696.450 709.950 ;
        RECT 737.400 706.050 738.450 739.950 ;
        RECT 740.400 736.050 741.450 754.950 ;
        RECT 745.950 754.800 748.050 756.900 ;
        RECT 751.950 754.800 754.050 756.900 ;
        RECT 758.400 755.400 759.600 757.650 ;
        RECT 764.400 756.900 765.600 757.650 ;
        RECT 773.400 756.900 774.450 775.950 ;
        RECT 779.400 772.050 780.450 800.400 ;
        RECT 784.950 799.800 787.050 801.900 ;
        RECT 796.950 799.800 799.050 801.900 ;
        RECT 805.950 799.950 808.050 802.050 ;
        RECT 812.400 801.000 813.600 802.650 ;
        RECT 797.400 799.050 798.450 799.800 ;
        RECT 797.400 797.400 802.050 799.050 ;
        RECT 798.000 796.950 802.050 797.400 ;
        RECT 806.400 778.050 807.450 799.950 ;
        RECT 811.950 796.950 814.050 801.000 ;
        RECT 821.400 800.400 822.600 802.650 ;
        RECT 805.950 775.950 808.050 778.050 ;
        RECT 821.400 775.050 822.450 800.400 ;
        RECT 820.950 772.950 823.050 775.050 ;
        RECT 778.950 769.950 781.050 772.050 ;
        RECT 827.400 769.050 828.450 806.100 ;
        RECT 833.400 805.350 834.600 806.100 ;
        RECT 839.400 805.350 840.600 806.100 ;
        RECT 832.950 802.950 835.050 805.050 ;
        RECT 835.950 802.950 838.050 805.050 ;
        RECT 838.950 802.950 841.050 805.050 ;
        RECT 836.400 801.900 837.600 802.650 ;
        RECT 845.400 801.900 846.450 806.100 ;
        RECT 854.400 805.350 855.600 807.600 ;
        RECT 850.950 802.950 853.050 805.050 ;
        RECT 853.950 802.950 856.050 805.050 ;
        RECT 856.950 802.950 859.050 805.050 ;
        RECT 851.400 801.900 852.600 802.650 ;
        RECT 835.950 799.800 838.050 801.900 ;
        RECT 844.950 799.800 847.050 801.900 ;
        RECT 850.950 799.800 853.050 801.900 ;
        RECT 857.400 800.400 858.600 802.650 ;
        RECT 836.250 769.500 838.350 770.400 ;
        RECT 817.950 766.950 820.050 769.050 ;
        RECT 826.950 766.950 829.050 769.050 ;
        RECT 834.150 768.300 838.350 769.500 ;
        RECT 781.950 761.100 784.050 763.200 ;
        RECT 782.400 760.350 783.600 761.100 ;
        RECT 790.950 760.950 793.050 763.050 ;
        RECT 799.950 761.100 802.050 763.200 ;
        RECT 808.950 761.100 811.050 763.200 ;
        RECT 818.400 762.600 819.450 766.950 ;
        RECT 778.950 757.950 781.050 760.050 ;
        RECT 781.950 757.950 784.050 760.050 ;
        RECT 784.950 757.950 787.050 760.050 ;
        RECT 758.400 745.050 759.450 755.400 ;
        RECT 763.950 754.800 766.050 756.900 ;
        RECT 772.800 754.800 774.900 756.900 ;
        RECT 775.950 756.450 778.050 757.050 ;
        RECT 779.400 756.450 780.600 757.650 ;
        RECT 785.400 756.900 786.600 757.650 ;
        RECT 791.400 756.900 792.450 760.950 ;
        RECT 800.400 760.350 801.600 761.100 ;
        RECT 796.950 757.950 799.050 760.050 ;
        RECT 799.950 757.950 802.050 760.050 ;
        RECT 802.950 757.950 805.050 760.050 ;
        RECT 775.950 755.400 780.600 756.450 ;
        RECT 775.950 754.950 778.050 755.400 ;
        RECT 757.950 742.950 760.050 745.050 ;
        RECT 739.950 733.950 742.050 736.050 ;
        RECT 743.550 735.300 745.650 737.400 ;
        RECT 748.950 736.950 751.050 739.050 ;
        RECT 739.950 727.950 742.050 730.050 ;
        RECT 740.400 721.050 741.450 727.950 ;
        RECT 743.550 722.400 744.750 735.300 ;
        RECT 749.400 729.600 750.450 736.950 ;
        RECT 757.950 733.950 760.050 736.050 ;
        RECT 769.950 733.950 772.050 736.050 ;
        RECT 749.400 727.350 750.600 729.600 ;
        RECT 748.950 724.950 751.050 727.050 ;
        RECT 739.950 718.950 742.050 721.050 ;
        RECT 743.550 720.300 745.650 722.400 ;
        RECT 743.550 713.700 744.750 720.300 ;
        RECT 758.400 718.050 759.450 733.950 ;
        RECT 763.950 728.100 766.050 730.200 ;
        RECT 770.400 729.600 771.450 733.950 ;
        RECT 764.400 727.350 765.600 728.100 ;
        RECT 770.400 727.350 771.600 729.600 ;
        RECT 763.950 724.950 766.050 727.050 ;
        RECT 766.950 724.950 769.050 727.050 ;
        RECT 769.950 724.950 772.050 727.050 ;
        RECT 767.400 723.900 768.600 724.650 ;
        RECT 776.400 724.050 777.450 754.950 ;
        RECT 784.950 754.800 787.050 756.900 ;
        RECT 790.950 754.800 793.050 756.900 ;
        RECT 797.400 755.400 798.600 757.650 ;
        RECT 803.400 755.400 804.600 757.650 ;
        RECT 784.950 745.950 787.050 748.050 ;
        RECT 790.950 745.950 793.050 748.050 ;
        RECT 785.400 729.600 786.450 745.950 ;
        RECT 785.400 727.350 786.600 729.600 ;
        RECT 781.950 724.950 784.050 727.050 ;
        RECT 784.950 724.950 787.050 727.050 ;
        RECT 766.950 721.800 769.050 723.900 ;
        RECT 775.950 721.950 778.050 724.050 ;
        RECT 782.400 722.400 783.600 724.650 ;
        RECT 782.400 718.050 783.450 722.400 ;
        RECT 751.950 715.950 754.050 718.050 ;
        RECT 757.950 715.950 760.050 718.050 ;
        RECT 781.950 715.950 784.050 718.050 ;
        RECT 743.550 711.600 745.650 713.700 ;
        RECT 730.950 703.950 733.050 706.050 ;
        RECT 736.950 703.950 739.050 706.050 ;
        RECT 727.950 694.950 730.050 697.050 ;
        RECT 703.950 683.100 706.050 685.200 ;
        RECT 704.400 682.350 705.600 683.100 ;
        RECT 712.950 682.950 715.050 685.050 ;
        RECT 721.950 683.100 724.050 685.200 ;
        RECT 728.400 685.050 729.450 694.950 ;
        RECT 700.950 679.950 703.050 682.050 ;
        RECT 703.950 679.950 706.050 682.050 ;
        RECT 706.950 679.950 709.050 682.050 ;
        RECT 701.400 678.000 702.600 679.650 ;
        RECT 707.400 678.900 708.600 679.650 ;
        RECT 713.400 678.900 714.450 682.950 ;
        RECT 722.400 682.350 723.600 683.100 ;
        RECT 727.950 682.950 730.050 685.050 ;
        RECT 718.950 679.950 721.050 682.050 ;
        RECT 721.950 679.950 724.050 682.050 ;
        RECT 724.950 679.950 727.050 682.050 ;
        RECT 700.950 673.950 703.050 678.000 ;
        RECT 706.950 676.800 709.050 678.900 ;
        RECT 712.950 676.800 715.050 678.900 ;
        RECT 719.400 677.400 720.600 679.650 ;
        RECT 725.400 677.400 726.600 679.650 ;
        RECT 701.400 664.050 702.450 673.950 ;
        RECT 692.400 662.400 696.450 663.450 ;
        RECT 692.400 645.900 693.450 662.400 ;
        RECT 700.950 661.950 703.050 664.050 ;
        RECT 695.550 657.300 697.650 659.400 ;
        RECT 691.950 643.800 694.050 645.900 ;
        RECT 695.550 644.400 696.750 657.300 ;
        RECT 700.950 655.950 703.050 658.050 ;
        RECT 701.400 651.600 702.450 655.950 ;
        RECT 719.400 652.200 720.450 677.400 ;
        RECT 725.400 664.050 726.450 677.400 ;
        RECT 731.400 670.050 732.450 703.950 ;
        RECT 733.950 688.950 736.050 691.050 ;
        RECT 739.950 688.950 742.050 691.050 ;
        RECT 734.400 685.050 735.450 688.950 ;
        RECT 733.950 682.950 736.050 685.050 ;
        RECT 740.400 684.600 741.450 688.950 ;
        RECT 740.400 682.350 741.600 684.600 ;
        RECT 745.950 683.100 748.050 685.200 ;
        RECT 746.400 682.350 747.600 683.100 ;
        RECT 736.950 679.950 739.050 682.050 ;
        RECT 739.950 679.950 742.050 682.050 ;
        RECT 742.950 679.950 745.050 682.050 ;
        RECT 745.950 679.950 748.050 682.050 ;
        RECT 737.400 679.050 738.600 679.650 ;
        RECT 733.950 677.400 738.600 679.050 ;
        RECT 743.400 677.400 744.600 679.650 ;
        RECT 733.950 676.950 738.000 677.400 ;
        RECT 743.400 676.050 744.450 677.400 ;
        RECT 748.950 676.950 751.050 679.050 ;
        RECT 742.950 673.950 745.050 676.050 ;
        RECT 730.950 667.950 733.050 670.050 ;
        RECT 724.950 661.950 727.050 664.050 ;
        RECT 725.400 658.050 726.450 661.950 ;
        RECT 724.950 655.950 727.050 658.050 ;
        RECT 743.400 655.050 744.450 673.950 ;
        RECT 745.950 667.950 748.050 670.050 ;
        RECT 742.950 652.950 745.050 655.050 ;
        RECT 701.400 649.350 702.600 651.600 ;
        RECT 718.950 650.100 721.050 652.200 ;
        RECT 719.400 649.350 720.600 650.100 ;
        RECT 724.950 649.950 727.050 652.050 ;
        RECT 730.950 650.100 733.050 652.200 ;
        RECT 737.400 651.450 738.600 651.600 ;
        RECT 737.400 650.400 744.450 651.450 ;
        RECT 700.950 646.950 703.050 649.050 ;
        RECT 715.950 646.950 718.050 649.050 ;
        RECT 718.950 646.950 721.050 649.050 ;
        RECT 716.400 645.900 717.600 646.650 ;
        RECT 695.550 642.300 697.650 644.400 ;
        RECT 715.950 643.800 718.050 645.900 ;
        RECT 695.550 635.700 696.750 642.300 ;
        RECT 703.950 640.950 706.050 643.050 ;
        RECT 695.550 633.600 697.650 635.700 ;
        RECT 688.950 625.950 691.050 628.050 ;
        RECT 694.950 622.950 697.050 625.050 ;
        RECT 685.950 613.950 688.050 616.050 ;
        RECT 676.950 610.950 679.050 613.050 ;
        RECT 673.950 607.950 676.050 610.050 ;
        RECT 677.400 607.200 678.450 610.950 ;
        RECT 671.400 604.350 672.600 606.600 ;
        RECT 676.950 605.100 679.050 607.200 ;
        RECT 682.950 605.100 685.050 607.200 ;
        RECT 688.950 605.100 691.050 607.200 ;
        RECT 695.400 606.600 696.450 622.950 ;
        RECT 704.400 622.050 705.450 640.950 ;
        RECT 716.400 625.050 717.450 643.800 ;
        RECT 715.950 622.950 718.050 625.050 ;
        RECT 703.950 619.950 706.050 622.050 ;
        RECT 725.400 621.450 726.450 649.950 ;
        RECT 731.400 649.350 732.600 650.100 ;
        RECT 737.400 649.350 738.600 650.400 ;
        RECT 730.950 646.950 733.050 649.050 ;
        RECT 733.950 646.950 736.050 649.050 ;
        RECT 736.950 646.950 739.050 649.050 ;
        RECT 734.400 645.900 735.600 646.650 ;
        RECT 743.400 646.050 744.450 650.400 ;
        RECT 733.950 643.800 736.050 645.900 ;
        RECT 742.950 645.450 745.050 646.050 ;
        RECT 740.400 644.400 745.050 645.450 ;
        RECT 736.950 640.950 739.050 643.050 ;
        RECT 722.400 620.400 726.450 621.450 ;
        RECT 704.400 606.600 705.450 619.950 ;
        RECT 710.250 613.500 712.350 614.400 ;
        RECT 718.950 613.950 721.050 616.050 ;
        RECT 708.150 612.300 712.350 613.500 ;
        RECT 677.400 604.350 678.600 605.100 ;
        RECT 670.950 601.950 673.050 604.050 ;
        RECT 673.950 601.950 676.050 604.050 ;
        RECT 676.950 601.950 679.050 604.050 ;
        RECT 655.950 598.800 658.050 600.900 ;
        RECT 664.950 598.950 667.050 601.050 ;
        RECT 674.400 599.400 675.600 601.650 ;
        RECT 674.400 595.050 675.450 599.400 ;
        RECT 683.400 595.050 684.450 605.100 ;
        RECT 689.400 604.350 690.600 605.100 ;
        RECT 695.400 604.350 696.600 606.600 ;
        RECT 704.400 604.350 705.600 606.600 ;
        RECT 688.950 601.950 691.050 604.050 ;
        RECT 691.950 601.950 694.050 604.050 ;
        RECT 694.950 601.950 697.050 604.050 ;
        RECT 697.950 601.950 700.050 604.050 ;
        RECT 703.950 601.950 706.050 604.050 ;
        RECT 692.400 600.900 693.600 601.650 ;
        RECT 691.950 598.800 694.050 600.900 ;
        RECT 698.400 600.000 699.600 601.650 ;
        RECT 688.950 595.950 691.050 598.050 ;
        RECT 697.950 595.950 700.050 600.000 ;
        RECT 673.950 592.950 676.050 595.050 ;
        RECT 682.950 592.950 685.050 595.050 ;
        RECT 640.950 574.950 643.050 577.050 ;
        RECT 646.950 574.950 649.050 577.050 ;
        RECT 641.400 568.050 642.450 574.950 ;
        RECT 649.950 571.950 652.050 574.050 ;
        RECT 680.400 573.450 681.600 573.600 ;
        RECT 677.400 572.400 681.600 573.450 ;
        RECT 646.800 568.950 648.900 571.050 ;
        RECT 640.950 565.950 643.050 568.050 ;
        RECT 650.400 565.050 651.450 571.950 ;
        RECT 664.800 568.950 666.900 571.050 ;
        RECT 665.400 567.900 666.600 568.650 ;
        RECT 664.950 567.450 667.050 567.900 ;
        RECT 662.400 566.400 667.050 567.450 ;
        RECT 643.950 562.950 646.050 565.050 ;
        RECT 649.950 562.950 652.050 565.050 ;
        RECT 637.950 553.950 640.050 556.050 ;
        RECT 628.950 538.950 631.050 541.050 ;
        RECT 634.950 538.950 637.050 541.050 ;
        RECT 625.950 535.950 628.050 538.050 ;
        RECT 632.250 535.500 634.350 536.400 ;
        RECT 630.150 534.300 634.350 535.500 ;
        RECT 626.400 528.450 627.600 528.600 ;
        RECT 623.400 527.400 627.600 528.450 ;
        RECT 620.400 526.350 621.600 527.100 ;
        RECT 626.400 526.350 627.600 527.400 ;
        RECT 610.950 523.950 613.050 526.050 ;
        RECT 613.950 523.950 616.050 526.050 ;
        RECT 616.950 523.950 619.050 526.050 ;
        RECT 619.950 523.950 622.050 526.050 ;
        RECT 625.950 523.950 628.050 526.050 ;
        RECT 611.400 521.400 612.600 523.650 ;
        RECT 617.400 522.900 618.600 523.650 ;
        RECT 604.950 517.950 607.050 520.050 ;
        RECT 611.400 514.050 612.450 521.400 ;
        RECT 616.950 520.800 619.050 522.900 ;
        RECT 613.950 517.950 616.050 520.050 ;
        RECT 610.950 511.950 613.050 514.050 ;
        RECT 614.400 501.450 615.450 517.950 ;
        RECT 630.150 515.700 631.350 534.300 ;
        RECT 634.950 528.000 637.050 532.050 ;
        RECT 640.950 529.950 643.050 532.050 ;
        RECT 635.400 526.350 636.600 528.000 ;
        RECT 635.100 523.950 637.200 526.050 ;
        RECT 641.400 523.050 642.450 529.950 ;
        RECT 640.950 520.950 643.050 523.050 ;
        RECT 644.400 517.050 645.450 562.950 ;
        RECT 647.550 537.300 649.650 539.400 ;
        RECT 647.550 530.700 648.750 537.300 ;
        RECT 647.550 528.600 649.650 530.700 ;
        RECT 629.850 513.600 631.950 515.700 ;
        RECT 643.950 514.950 646.050 517.050 ;
        RECT 647.550 515.700 648.750 528.600 ;
        RECT 658.950 527.100 661.050 529.200 ;
        RECT 652.950 523.950 655.050 526.050 ;
        RECT 653.400 522.900 654.600 523.650 ;
        RECT 659.400 523.050 660.450 527.100 ;
        RECT 652.950 520.800 655.050 522.900 ;
        RECT 658.950 520.950 661.050 523.050 ;
        RECT 647.550 513.600 649.650 515.700 ;
        RECT 643.950 508.950 646.050 511.050 ;
        RECT 610.800 498.300 612.900 500.400 ;
        RECT 614.400 499.200 615.600 501.450 ;
        RECT 628.950 499.950 631.050 502.050 ;
        RECT 644.400 501.450 645.450 508.950 ;
        RECT 662.400 502.050 663.450 566.400 ;
        RECT 664.950 565.800 667.050 566.400 ;
        RECT 673.950 565.950 676.050 568.050 ;
        RECT 674.400 559.050 675.450 565.950 ;
        RECT 673.950 556.950 676.050 559.050 ;
        RECT 677.400 547.050 678.450 572.400 ;
        RECT 680.400 571.350 681.600 572.400 ;
        RECT 680.400 568.950 682.500 571.050 ;
        RECT 685.800 568.950 687.900 571.050 ;
        RECT 686.400 566.400 687.600 568.650 ;
        RECT 686.400 562.050 687.450 566.400 ;
        RECT 685.950 559.950 688.050 562.050 ;
        RECT 676.950 544.950 679.050 547.050 ;
        RECT 689.400 535.050 690.450 595.950 ;
        RECT 708.150 593.700 709.350 612.300 ;
        RECT 712.950 605.100 715.050 607.200 ;
        RECT 713.400 604.350 714.600 605.100 ;
        RECT 713.100 601.950 715.200 604.050 ;
        RECT 719.400 595.050 720.450 613.950 ;
        RECT 722.400 600.900 723.450 620.400 ;
        RECT 725.550 615.300 727.650 617.400 ;
        RECT 725.550 608.700 726.750 615.300 ;
        RECT 725.550 606.600 727.650 608.700 ;
        RECT 721.950 598.800 724.050 600.900 ;
        RECT 707.850 591.600 709.950 593.700 ;
        RECT 718.950 592.950 721.050 595.050 ;
        RECT 725.550 593.700 726.750 606.600 ;
        RECT 730.950 601.950 733.050 604.050 ;
        RECT 731.400 600.900 732.600 601.650 ;
        RECT 730.950 598.800 733.050 600.900 ;
        RECT 725.550 591.600 727.650 593.700 ;
        RECT 737.400 589.050 738.450 640.950 ;
        RECT 740.400 600.900 741.450 644.400 ;
        RECT 742.950 643.950 745.050 644.400 ;
        RECT 746.400 634.050 747.450 667.950 ;
        RECT 749.400 652.050 750.450 676.950 ;
        RECT 752.400 673.050 753.450 715.950 ;
        RECT 772.950 709.950 775.050 712.050 ;
        RECT 769.950 700.950 772.050 703.050 ;
        RECT 754.950 688.950 757.050 691.050 ;
        RECT 755.400 678.900 756.450 688.950 ;
        RECT 763.950 683.100 766.050 685.200 ;
        RECT 770.400 685.050 771.450 700.950 ;
        RECT 764.400 682.350 765.600 683.100 ;
        RECT 769.950 682.950 772.050 685.050 ;
        RECT 773.400 684.600 774.450 709.950 ;
        RECT 779.250 691.500 781.350 692.400 ;
        RECT 777.150 690.300 781.350 691.500 ;
        RECT 773.400 682.350 774.600 684.600 ;
        RECT 760.950 679.950 763.050 682.050 ;
        RECT 763.950 679.950 766.050 682.050 ;
        RECT 766.950 679.950 769.050 682.050 ;
        RECT 772.950 679.950 775.050 682.050 ;
        RECT 754.950 676.800 757.050 678.900 ;
        RECT 761.400 677.400 762.600 679.650 ;
        RECT 767.400 678.900 768.600 679.650 ;
        RECT 761.400 675.450 762.450 677.400 ;
        RECT 766.950 676.800 769.050 678.900 ;
        RECT 761.400 674.400 765.450 675.450 ;
        RECT 751.950 670.950 754.050 673.050 ;
        RECT 760.950 670.950 763.050 673.050 ;
        RECT 754.950 661.950 757.050 664.050 ;
        RECT 748.950 649.950 751.050 652.050 ;
        RECT 755.400 651.600 756.450 661.950 ;
        RECT 755.400 649.350 756.600 651.600 ;
        RECT 751.950 646.950 754.050 649.050 ;
        RECT 754.950 646.950 757.050 649.050 ;
        RECT 752.400 645.900 753.600 646.650 ;
        RECT 751.950 643.800 754.050 645.900 ;
        RECT 745.950 631.950 748.050 634.050 ;
        RECT 748.950 610.950 751.050 613.050 ;
        RECT 749.400 606.600 750.450 610.950 ;
        RECT 761.400 610.050 762.450 670.950 ;
        RECT 764.400 664.050 765.450 674.400 ;
        RECT 777.150 671.700 778.350 690.300 ;
        RECT 781.950 683.100 784.050 685.200 ;
        RECT 787.950 683.100 790.050 685.200 ;
        RECT 782.400 682.350 783.600 683.100 ;
        RECT 782.100 679.950 784.200 682.050 ;
        RECT 776.850 669.600 778.950 671.700 ;
        RECT 781.950 670.950 784.050 673.050 ;
        RECT 778.950 664.950 781.050 667.050 ;
        RECT 763.950 661.950 766.050 664.050 ;
        RECT 769.950 650.100 772.050 652.200 ;
        RECT 770.400 649.350 771.600 650.100 ;
        RECT 775.950 649.950 778.050 655.050 ;
        RECT 766.950 646.950 769.050 649.050 ;
        RECT 769.950 646.950 772.050 649.050 ;
        RECT 772.950 646.950 775.050 649.050 ;
        RECT 767.400 644.400 768.600 646.650 ;
        RECT 773.400 645.900 774.600 646.650 ;
        RECT 767.400 628.050 768.450 644.400 ;
        RECT 772.950 643.800 775.050 645.900 ;
        RECT 779.400 643.050 780.450 664.950 ;
        RECT 782.400 652.050 783.450 670.950 ;
        RECT 788.400 667.050 789.450 683.100 ;
        RECT 791.400 678.900 792.450 745.950 ;
        RECT 797.400 739.050 798.450 755.400 ;
        RECT 803.400 748.050 804.450 755.400 ;
        RECT 802.950 745.950 805.050 748.050 ;
        RECT 809.400 745.050 810.450 761.100 ;
        RECT 818.400 760.350 819.600 762.600 ;
        RECT 823.950 761.100 826.050 763.200 ;
        RECT 829.950 761.100 832.050 763.200 ;
        RECT 824.400 760.350 825.600 761.100 ;
        RECT 830.400 760.350 831.600 761.100 ;
        RECT 814.950 757.950 817.050 760.050 ;
        RECT 817.950 757.950 820.050 760.050 ;
        RECT 820.950 757.950 823.050 760.050 ;
        RECT 823.950 757.950 826.050 760.050 ;
        RECT 829.950 757.950 832.050 760.050 ;
        RECT 815.400 755.400 816.600 757.650 ;
        RECT 821.400 755.400 822.600 757.650 ;
        RECT 815.400 751.050 816.450 755.400 ;
        RECT 821.400 751.050 822.450 755.400 ;
        RECT 823.950 751.950 826.050 754.050 ;
        RECT 814.950 748.950 817.050 751.050 ;
        RECT 820.950 748.950 823.050 751.050 ;
        RECT 808.950 742.950 811.050 745.050 ;
        RECT 820.950 742.950 823.050 745.050 ;
        RECT 796.950 736.950 799.050 739.050 ;
        RECT 797.400 729.600 798.450 736.950 ;
        RECT 809.850 735.300 811.950 737.400 ;
        RECT 797.400 727.350 798.600 729.600 ;
        RECT 796.950 724.950 799.050 727.050 ;
        RECT 799.950 724.950 802.050 727.050 ;
        RECT 805.950 724.950 808.050 727.050 ;
        RECT 800.400 723.900 801.600 724.650 ;
        RECT 806.400 723.900 807.600 724.650 ;
        RECT 799.950 721.800 802.050 723.900 ;
        RECT 805.950 721.800 808.050 723.900 ;
        RECT 806.400 712.050 807.450 721.800 ;
        RECT 810.150 716.700 811.350 735.300 ;
        RECT 815.100 724.950 817.200 727.050 ;
        RECT 815.400 723.450 816.600 724.650 ;
        RECT 815.400 722.400 819.450 723.450 ;
        RECT 810.150 715.500 814.350 716.700 ;
        RECT 812.250 714.600 814.350 715.500 ;
        RECT 805.950 709.950 808.050 712.050 ;
        RECT 818.400 709.050 819.450 722.400 ;
        RECT 808.950 706.950 811.050 709.050 ;
        RECT 817.950 706.950 820.050 709.050 ;
        RECT 794.550 693.300 796.650 695.400 ;
        RECT 794.550 686.700 795.750 693.300 ;
        RECT 794.550 684.600 796.650 686.700 ;
        RECT 790.950 676.800 793.050 678.900 ;
        RECT 794.550 671.700 795.750 684.600 ;
        RECT 799.950 679.950 802.050 682.050 ;
        RECT 805.950 679.950 808.050 682.050 ;
        RECT 800.400 678.900 801.600 679.650 ;
        RECT 799.950 676.800 802.050 678.900 ;
        RECT 794.550 669.600 796.650 671.700 ;
        RECT 787.950 664.950 790.050 667.050 ;
        RECT 806.400 664.050 807.450 679.950 ;
        RECT 805.950 661.950 808.050 664.050 ;
        RECT 781.950 649.950 784.050 652.050 ;
        RECT 787.950 650.100 790.050 652.200 ;
        RECT 788.400 649.350 789.600 650.100 ;
        RECT 796.950 649.950 799.050 652.050 ;
        RECT 802.950 650.100 805.050 652.200 ;
        RECT 809.400 651.600 810.450 706.950 ;
        RECT 821.400 706.050 822.450 742.950 ;
        RECT 824.400 724.050 825.450 751.950 ;
        RECT 834.150 749.700 835.350 768.300 ;
        RECT 838.950 761.100 841.050 763.200 ;
        RECT 839.400 760.350 840.600 761.100 ;
        RECT 839.100 757.950 841.200 760.050 ;
        RECT 845.400 756.450 846.450 799.800 ;
        RECT 851.550 771.300 853.650 773.400 ;
        RECT 851.550 764.700 852.750 771.300 ;
        RECT 857.400 769.050 858.450 800.400 ;
        RECT 856.950 766.950 859.050 769.050 ;
        RECT 862.950 766.950 865.050 769.050 ;
        RECT 847.950 760.950 850.050 763.050 ;
        RECT 851.550 762.600 853.650 764.700 ;
        RECT 842.400 755.400 846.450 756.450 ;
        RECT 833.850 747.600 835.950 749.700 ;
        RECT 827.550 735.300 829.650 737.400 ;
        RECT 823.950 721.950 826.050 724.050 ;
        RECT 827.550 722.400 828.750 735.300 ;
        RECT 832.950 733.950 835.050 736.050 ;
        RECT 833.400 729.600 834.450 733.950 ;
        RECT 833.400 727.350 834.600 729.600 ;
        RECT 832.950 724.950 835.050 727.050 ;
        RECT 842.400 724.050 843.450 755.400 ;
        RECT 848.400 751.050 849.450 760.950 ;
        RECT 847.950 748.950 850.050 751.050 ;
        RECT 851.550 749.700 852.750 762.600 ;
        RECT 856.950 757.950 859.050 760.050 ;
        RECT 857.400 755.400 858.600 757.650 ;
        RECT 851.550 747.600 853.650 749.700 ;
        RECT 857.400 739.050 858.450 755.400 ;
        RECT 856.950 736.950 859.050 739.050 ;
        RECT 853.950 735.900 858.000 736.050 ;
        RECT 853.950 733.950 859.050 735.900 ;
        RECT 863.400 735.450 864.450 766.950 ;
        RECT 874.950 736.950 877.050 739.050 ;
        RECT 856.950 733.800 859.050 733.950 ;
        RECT 860.400 734.400 864.450 735.450 ;
        RECT 850.950 728.100 853.050 730.200 ;
        RECT 851.400 727.350 852.600 728.100 ;
        RECT 856.950 727.950 859.050 732.900 ;
        RECT 847.950 724.950 850.050 727.050 ;
        RECT 850.950 724.950 853.050 727.050 ;
        RECT 853.950 724.950 856.050 727.050 ;
        RECT 827.550 720.300 829.650 722.400 ;
        RECT 841.950 721.950 844.050 724.050 ;
        RECT 848.400 723.450 849.600 724.650 ;
        RECT 845.400 722.400 849.600 723.450 ;
        RECT 854.400 722.400 855.600 724.650 ;
        RECT 827.550 713.700 828.750 720.300 ;
        RECT 827.550 711.600 829.650 713.700 ;
        RECT 820.950 703.950 823.050 706.050 ;
        RECT 826.950 703.950 829.050 706.050 ;
        RECT 817.950 683.100 820.050 685.200 ;
        RECT 818.400 682.350 819.600 683.100 ;
        RECT 814.950 679.950 817.050 682.050 ;
        RECT 817.950 679.950 820.050 682.050 ;
        RECT 820.950 679.950 823.050 682.050 ;
        RECT 815.400 678.900 816.600 679.650 ;
        RECT 814.950 676.800 817.050 678.900 ;
        RECT 821.400 677.400 822.600 679.650 ;
        RECT 815.400 673.050 816.450 676.800 ;
        RECT 814.950 670.950 817.050 673.050 ;
        RECT 815.400 664.050 816.450 670.950 ;
        RECT 821.400 670.050 822.450 677.400 ;
        RECT 820.950 667.950 823.050 670.050 ;
        RECT 827.400 667.050 828.450 703.950 ;
        RECT 835.950 688.950 838.050 691.050 ;
        RECT 841.950 688.950 844.050 691.050 ;
        RECT 836.400 684.600 837.450 688.950 ;
        RECT 836.400 682.350 837.600 684.600 ;
        RECT 832.950 679.950 835.050 682.050 ;
        RECT 835.950 679.950 838.050 682.050 ;
        RECT 833.400 677.400 834.600 679.650 ;
        RECT 833.400 673.050 834.450 677.400 ;
        RECT 838.950 676.950 841.050 679.050 ;
        RECT 832.950 670.950 835.050 673.050 ;
        RECT 835.950 667.950 838.050 670.050 ;
        RECT 826.950 664.950 829.050 667.050 ;
        RECT 832.950 664.950 835.050 667.050 ;
        RECT 814.950 661.950 817.050 664.050 ;
        RECT 814.950 655.950 817.050 658.050 ;
        RECT 824.850 657.300 826.950 659.400 ;
        RECT 815.400 651.600 816.450 655.950 ;
        RECT 784.950 646.950 787.050 649.050 ;
        RECT 787.950 646.950 790.050 649.050 ;
        RECT 790.950 646.950 793.050 649.050 ;
        RECT 785.400 646.050 786.600 646.650 ;
        RECT 781.950 644.400 786.600 646.050 ;
        RECT 791.400 644.400 792.600 646.650 ;
        RECT 781.950 643.950 786.000 644.400 ;
        RECT 772.950 640.650 775.050 642.750 ;
        RECT 778.950 640.950 781.050 643.050 ;
        RECT 766.950 625.950 769.050 628.050 ;
        RECT 760.950 607.950 763.050 610.050 ;
        RECT 749.400 604.350 750.600 606.600 ;
        RECT 754.950 605.100 757.050 607.200 ;
        RECT 755.400 604.350 756.600 605.100 ;
        RECT 760.950 604.800 763.050 606.900 ;
        RECT 766.950 606.000 769.050 610.050 ;
        RECT 773.400 606.600 774.450 640.650 ;
        RECT 775.950 625.950 778.050 628.050 ;
        RECT 776.400 610.050 777.450 625.950 ;
        RECT 787.950 616.950 790.050 619.050 ;
        RECT 775.950 607.950 778.050 610.050 ;
        RECT 745.950 601.950 748.050 604.050 ;
        RECT 748.950 601.950 751.050 604.050 ;
        RECT 751.950 601.950 754.050 604.050 ;
        RECT 754.950 601.950 757.050 604.050 ;
        RECT 746.400 600.900 747.600 601.650 ;
        RECT 739.950 598.800 742.050 600.900 ;
        RECT 745.950 598.800 748.050 600.900 ;
        RECT 752.400 599.400 753.600 601.650 ;
        RECT 752.400 595.050 753.450 599.400 ;
        RECT 751.950 592.950 754.050 595.050 ;
        RECT 727.950 586.950 730.050 589.050 ;
        RECT 736.950 586.950 739.050 589.050 ;
        RECT 691.950 568.950 694.050 574.050 ;
        RECT 697.950 573.000 700.050 577.050 ;
        RECT 698.400 571.350 699.600 573.000 ;
        RECT 703.950 572.100 706.050 574.200 ;
        RECT 704.400 571.350 705.600 572.100 ;
        RECT 712.950 571.950 715.050 574.050 ;
        RECT 721.950 572.100 724.050 574.200 ;
        RECT 728.400 574.050 729.450 586.950 ;
        RECT 761.400 586.050 762.450 604.800 ;
        RECT 767.400 604.350 768.600 606.000 ;
        RECT 773.400 604.350 774.600 606.600 ;
        RECT 778.950 606.000 781.050 610.050 ;
        RECT 784.950 607.950 787.050 610.050 ;
        RECT 779.400 604.350 780.600 606.000 ;
        RECT 766.950 601.950 769.050 604.050 ;
        RECT 769.950 601.950 772.050 604.050 ;
        RECT 772.950 601.950 775.050 604.050 ;
        RECT 775.950 601.950 778.050 604.050 ;
        RECT 778.950 601.950 781.050 604.050 ;
        RECT 770.400 600.900 771.600 601.650 ;
        RECT 769.950 598.800 772.050 600.900 ;
        RECT 776.400 599.400 777.600 601.650 ;
        RECT 766.950 595.950 769.050 598.050 ;
        RECT 748.950 583.950 751.050 586.050 ;
        RECT 760.950 583.950 763.050 586.050 ;
        RECT 734.850 579.300 736.950 581.400 ;
        RECT 697.950 568.950 700.050 571.050 ;
        RECT 700.950 568.950 703.050 571.050 ;
        RECT 703.950 568.950 706.050 571.050 ;
        RECT 706.950 568.950 709.050 571.050 ;
        RECT 691.950 565.800 694.050 567.900 ;
        RECT 694.950 565.950 697.050 568.050 ;
        RECT 701.400 567.900 702.600 568.650 ;
        RECT 707.400 567.900 708.600 568.650 ;
        RECT 713.400 567.900 714.450 571.950 ;
        RECT 722.400 571.350 723.600 572.100 ;
        RECT 727.950 571.950 730.050 574.050 ;
        RECT 718.950 568.950 721.050 571.050 ;
        RECT 721.950 568.950 724.050 571.050 ;
        RECT 724.950 568.950 727.050 571.050 ;
        RECT 730.950 568.950 733.050 571.050 ;
        RECT 692.400 541.050 693.450 565.800 ;
        RECT 695.400 556.050 696.450 565.950 ;
        RECT 700.950 562.950 703.050 567.900 ;
        RECT 706.950 565.800 709.050 567.900 ;
        RECT 712.950 565.800 715.050 567.900 ;
        RECT 719.400 567.000 720.600 568.650 ;
        RECT 725.400 567.000 726.600 568.650 ;
        RECT 718.950 562.950 721.050 567.000 ;
        RECT 724.950 562.950 727.050 567.000 ;
        RECT 727.950 565.950 730.050 568.050 ;
        RECT 731.400 566.400 732.600 568.650 ;
        RECT 694.950 553.950 697.050 556.050 ;
        RECT 728.400 550.050 729.450 565.950 ;
        RECT 731.400 559.050 732.450 566.400 ;
        RECT 735.150 560.700 736.350 579.300 ;
        RECT 745.950 572.100 748.050 574.200 ;
        RECT 740.100 568.950 742.200 571.050 ;
        RECT 740.400 567.450 741.600 568.650 ;
        RECT 740.400 566.400 744.450 567.450 ;
        RECT 735.150 559.500 739.350 560.700 ;
        RECT 730.950 556.950 733.050 559.050 ;
        RECT 737.250 558.600 739.350 559.500 ;
        RECT 743.400 556.050 744.450 566.400 ;
        RECT 746.400 565.050 747.450 572.100 ;
        RECT 745.950 562.950 748.050 565.050 ;
        RECT 742.950 553.950 745.050 556.050 ;
        RECT 749.400 552.450 750.450 583.950 ;
        RECT 752.550 579.300 754.650 581.400 ;
        RECT 752.550 566.400 753.750 579.300 ;
        RECT 757.950 572.100 760.050 574.200 ;
        RECT 758.400 571.350 759.600 572.100 ;
        RECT 757.950 568.950 760.050 571.050 ;
        RECT 752.550 564.300 754.650 566.400 ;
        RECT 763.950 565.800 766.050 567.900 ;
        RECT 752.550 557.700 753.750 564.300 ;
        RECT 760.950 562.950 763.050 565.050 ;
        RECT 752.550 555.600 754.650 557.700 ;
        RECT 761.400 556.050 762.450 562.950 ;
        RECT 760.950 553.950 763.050 556.050 ;
        RECT 749.400 551.400 753.450 552.450 ;
        RECT 727.950 547.950 730.050 550.050 ;
        RECT 748.950 547.950 751.050 550.050 ;
        RECT 700.950 544.950 703.050 547.050 ;
        RECT 691.950 538.950 694.050 541.050 ;
        RECT 673.950 532.950 676.050 535.050 ;
        RECT 688.950 532.950 691.050 535.050 ;
        RECT 667.950 527.100 670.050 529.200 ;
        RECT 674.400 528.600 675.450 532.950 ;
        RECT 668.400 526.350 669.600 527.100 ;
        RECT 674.400 526.350 675.600 528.600 ;
        RECT 685.950 527.100 688.050 529.200 ;
        RECT 692.400 528.600 693.450 538.950 ;
        RECT 686.400 526.350 687.600 527.100 ;
        RECT 692.400 526.350 693.600 528.600 ;
        RECT 667.950 523.950 670.050 526.050 ;
        RECT 670.950 523.950 673.050 526.050 ;
        RECT 673.950 523.950 676.050 526.050 ;
        RECT 685.950 523.950 688.050 526.050 ;
        RECT 688.950 523.950 691.050 526.050 ;
        RECT 691.950 523.950 694.050 526.050 ;
        RECT 671.400 521.400 672.600 523.650 ;
        RECT 689.400 522.900 690.600 523.650 ;
        RECT 671.400 517.050 672.450 521.400 ;
        RECT 688.950 520.800 691.050 522.900 ;
        RECT 701.400 522.450 702.450 544.950 ;
        RECT 709.950 538.950 712.050 541.050 ;
        RECT 710.400 535.050 711.450 538.950 ;
        RECT 712.950 535.950 715.050 538.050 ;
        RECT 709.950 532.950 712.050 535.050 ;
        RECT 710.400 528.600 711.450 532.950 ;
        RECT 710.400 526.350 711.600 528.600 ;
        RECT 704.400 523.950 706.500 526.050 ;
        RECT 709.800 523.950 711.900 526.050 ;
        RECT 704.400 522.450 705.600 523.650 ;
        RECT 701.400 521.400 705.600 522.450 ;
        RECT 670.950 514.950 673.050 517.050 ;
        RECT 706.950 511.950 709.050 514.050 ;
        RECT 691.950 508.950 694.050 511.050 ;
        RECT 601.950 493.950 604.050 496.050 ;
        RECT 608.400 495.450 609.600 495.600 ;
        RECT 605.400 494.400 609.600 495.450 ;
        RECT 592.950 490.950 595.050 493.050 ;
        RECT 593.400 489.900 594.600 490.650 ;
        RECT 592.950 487.800 595.050 489.900 ;
        RECT 571.350 477.600 573.450 479.700 ;
        RECT 553.950 466.950 556.050 469.050 ;
        RECT 565.950 454.950 568.050 457.050 ;
        RECT 544.950 449.100 547.050 451.200 ;
        RECT 566.400 450.600 567.450 454.950 ;
        RECT 545.400 448.350 546.600 449.100 ;
        RECT 566.400 448.350 567.600 450.600 ;
        RECT 571.950 449.100 574.050 451.200 ;
        RECT 572.400 448.350 573.600 449.100 ;
        RECT 545.100 445.950 547.200 448.050 ;
        RECT 550.500 445.950 552.600 448.050 ;
        RECT 565.950 445.950 568.050 448.050 ;
        RECT 568.950 445.950 571.050 448.050 ;
        RECT 571.950 445.950 574.050 448.050 ;
        RECT 574.950 445.950 577.050 448.050 ;
        RECT 551.400 443.400 552.600 445.650 ;
        RECT 569.400 443.400 570.600 445.650 ;
        RECT 575.400 444.900 576.600 445.650 ;
        RECT 581.400 445.050 582.450 481.950 ;
        RECT 586.650 481.500 590.850 482.700 ;
        RECT 586.650 480.600 588.750 481.500 ;
        RECT 605.400 463.050 606.450 494.400 ;
        RECT 608.400 493.350 609.600 494.400 ;
        RECT 608.100 490.950 610.200 493.050 ;
        RECT 611.100 492.900 612.000 498.300 ;
        RECT 614.100 496.800 616.200 498.900 ;
        RECT 618.000 495.900 620.100 497.700 ;
        RECT 612.900 494.700 621.600 495.900 ;
        RECT 612.900 493.800 615.000 494.700 ;
        RECT 611.100 491.700 618.000 492.900 ;
        RECT 611.100 484.500 612.300 491.700 ;
        RECT 614.100 487.950 616.200 490.050 ;
        RECT 617.100 489.300 618.000 491.700 ;
        RECT 614.400 485.400 615.600 487.650 ;
        RECT 617.100 487.200 619.200 489.300 ;
        RECT 620.700 485.700 621.600 494.700 ;
        RECT 622.800 490.950 624.900 493.050 ;
        RECT 623.400 489.450 624.600 490.650 ;
        RECT 629.400 489.900 630.450 499.950 ;
        RECT 644.400 499.200 645.600 501.450 ;
        RECT 639.900 495.900 642.000 497.700 ;
        RECT 643.800 496.800 645.900 498.900 ;
        RECT 647.100 498.300 649.200 500.400 ;
        RECT 661.950 499.950 664.050 502.050 ;
        RECT 638.400 494.700 647.100 495.900 ;
        RECT 635.100 490.950 637.200 493.050 ;
        RECT 623.400 488.400 627.450 489.450 ;
        RECT 610.800 482.400 612.900 484.500 ;
        RECT 620.400 483.600 622.500 485.700 ;
        RECT 626.400 469.050 627.450 488.400 ;
        RECT 628.950 487.800 631.050 489.900 ;
        RECT 635.400 489.450 636.600 490.650 ;
        RECT 632.400 488.400 636.600 489.450 ;
        RECT 632.400 475.050 633.450 488.400 ;
        RECT 638.400 485.700 639.300 494.700 ;
        RECT 645.000 493.800 647.100 494.700 ;
        RECT 648.000 492.900 648.900 498.300 ;
        RECT 692.400 496.200 693.450 508.950 ;
        RECT 700.950 499.950 703.050 502.050 ;
        RECT 701.400 496.200 702.450 499.950 ;
        RECT 649.950 494.100 652.050 496.200 ;
        RECT 655.950 494.100 658.050 496.200 ;
        RECT 664.950 494.100 667.050 496.200 ;
        RECT 670.950 494.100 673.050 496.200 ;
        RECT 650.400 493.350 651.600 494.100 ;
        RECT 642.000 491.700 648.900 492.900 ;
        RECT 642.000 489.300 642.900 491.700 ;
        RECT 640.800 487.200 642.900 489.300 ;
        RECT 643.800 487.950 645.900 490.050 ;
        RECT 637.500 483.600 639.600 485.700 ;
        RECT 644.400 485.400 645.600 487.650 ;
        RECT 647.700 484.500 648.900 491.700 ;
        RECT 649.800 490.950 651.900 493.050 ;
        RECT 647.100 482.400 649.200 484.500 ;
        RECT 631.950 472.950 634.050 475.050 ;
        RECT 616.950 466.950 619.050 469.050 ;
        RECT 625.950 466.950 628.050 469.050 ;
        RECT 589.950 460.950 592.050 463.050 ;
        RECT 604.950 460.950 607.050 463.050 ;
        RECT 590.400 450.600 591.450 460.950 ;
        RECT 601.950 454.950 604.050 457.050 ;
        RECT 602.400 451.200 603.450 454.950 ;
        RECT 590.400 448.350 591.600 450.600 ;
        RECT 595.950 449.100 598.050 451.200 ;
        RECT 601.950 449.100 604.050 451.200 ;
        RECT 610.950 449.100 613.050 451.200 ;
        RECT 596.400 448.350 597.600 449.100 ;
        RECT 586.950 445.950 589.050 448.050 ;
        RECT 589.950 445.950 592.050 448.050 ;
        RECT 592.950 445.950 595.050 448.050 ;
        RECT 595.950 445.950 598.050 448.050 ;
        RECT 551.400 424.050 552.450 443.400 ;
        RECT 550.950 421.950 553.050 424.050 ;
        RECT 553.950 421.950 556.050 424.050 ;
        RECT 565.350 423.300 567.450 425.400 ;
        RECT 554.400 417.600 555.450 421.950 ;
        RECT 554.400 415.350 555.600 417.600 ;
        RECT 559.950 416.100 562.050 418.200 ;
        RECT 560.400 415.350 561.600 416.100 ;
        RECT 548.100 412.950 550.200 415.050 ;
        RECT 553.500 412.950 555.600 415.050 ;
        RECT 559.950 412.950 562.050 415.050 ;
        RECT 548.400 410.400 549.600 412.650 ;
        RECT 566.250 410.400 567.450 423.300 ;
        RECT 541.950 403.950 544.050 406.050 ;
        RECT 548.400 382.050 549.450 410.400 ;
        RECT 565.350 408.300 567.450 410.400 ;
        RECT 550.950 403.950 553.050 406.050 ;
        RECT 538.950 379.950 541.050 382.050 ;
        RECT 547.950 379.950 550.050 382.050 ;
        RECT 535.950 370.950 538.050 373.050 ;
        RECT 539.400 372.600 540.450 379.950 ;
        RECT 539.400 370.350 540.600 372.600 ;
        RECT 548.400 372.450 549.450 379.950 ;
        RECT 551.400 379.050 552.450 403.950 ;
        RECT 566.250 401.700 567.450 408.300 ;
        RECT 565.350 399.600 567.450 401.700 ;
        RECT 569.400 400.050 570.450 443.400 ;
        RECT 574.950 442.800 577.050 444.900 ;
        RECT 580.950 442.950 583.050 445.050 ;
        RECT 587.400 443.400 588.600 445.650 ;
        RECT 593.400 443.400 594.600 445.650 ;
        RECT 587.400 439.050 588.450 443.400 ;
        RECT 586.950 436.950 589.050 439.050 ;
        RECT 593.400 433.050 594.450 443.400 ;
        RECT 602.400 439.050 603.450 449.100 ;
        RECT 611.400 448.350 612.600 449.100 ;
        RECT 607.950 445.950 610.050 448.050 ;
        RECT 610.950 445.950 613.050 448.050 ;
        RECT 608.400 443.400 609.600 445.650 ;
        RECT 617.400 445.050 618.450 466.950 ;
        RECT 625.950 449.100 628.050 451.200 ;
        RECT 632.400 450.600 633.450 472.950 ;
        RECT 649.950 454.950 652.050 457.050 ;
        RECT 626.400 448.350 627.600 449.100 ;
        RECT 632.400 448.350 633.600 450.600 ;
        RECT 637.950 449.100 640.050 451.200 ;
        RECT 643.950 449.100 646.050 451.200 ;
        RECT 650.400 450.600 651.450 454.950 ;
        RECT 622.950 445.950 625.050 448.050 ;
        RECT 625.950 445.950 628.050 448.050 ;
        RECT 628.950 445.950 631.050 448.050 ;
        RECT 631.950 445.950 634.050 448.050 ;
        RECT 608.400 439.050 609.450 443.400 ;
        RECT 616.950 442.950 619.050 445.050 ;
        RECT 623.400 444.900 624.600 445.650 ;
        RECT 622.950 442.800 625.050 444.900 ;
        RECT 629.400 443.400 630.600 445.650 ;
        RECT 595.950 436.950 598.050 439.050 ;
        RECT 601.950 436.950 604.050 439.050 ;
        RECT 607.950 436.950 610.050 439.050 ;
        RECT 592.950 430.950 595.050 433.050 ;
        RECT 571.950 421.950 574.050 424.050 ;
        RECT 583.050 423.300 585.150 425.400 ;
        RECT 572.400 412.050 573.450 421.950 ;
        RECT 577.800 412.950 579.900 415.050 ;
        RECT 571.950 409.950 574.050 412.050 ;
        RECT 578.400 411.900 579.600 412.650 ;
        RECT 577.950 409.800 580.050 411.900 ;
        RECT 583.650 404.700 584.850 423.300 ;
        RECT 592.950 416.100 595.050 418.200 ;
        RECT 586.950 412.950 589.050 415.050 ;
        RECT 587.400 411.900 588.600 412.650 ;
        RECT 586.950 409.800 589.050 411.900 ;
        RECT 580.650 403.500 584.850 404.700 ;
        RECT 580.650 402.600 582.750 403.500 ;
        RECT 568.950 397.950 571.050 400.050 ;
        RECT 583.950 391.950 586.050 394.050 ;
        RECT 562.950 388.950 565.050 391.050 ;
        RECT 550.950 376.950 553.050 379.050 ;
        RECT 563.400 376.050 564.450 388.950 ;
        RECT 584.400 376.050 585.450 391.950 ;
        RECT 587.400 382.050 588.450 409.800 ;
        RECT 589.950 406.950 592.050 409.050 ;
        RECT 586.950 379.950 589.050 382.050 ;
        RECT 562.950 373.950 565.050 376.050 ;
        RECT 563.400 372.600 564.450 373.950 ;
        RECT 548.400 371.400 552.450 372.450 ;
        RECT 538.950 367.950 541.050 370.050 ;
        RECT 541.950 367.950 544.050 370.050 ;
        RECT 544.950 367.950 547.050 370.050 ;
        RECT 542.400 365.400 543.600 367.650 ;
        RECT 532.950 355.950 535.050 358.050 ;
        RECT 542.400 346.050 543.450 365.400 ;
        RECT 551.400 346.050 552.450 371.400 ;
        RECT 563.400 370.350 564.600 372.600 ;
        RECT 571.950 371.100 574.050 373.200 ;
        RECT 577.950 371.100 580.050 373.200 ;
        RECT 583.950 372.000 586.050 376.050 ;
        RECT 590.400 373.050 591.450 406.950 ;
        RECT 593.400 400.050 594.450 416.100 ;
        RECT 596.400 409.050 597.450 436.950 ;
        RECT 629.400 433.050 630.450 443.400 ;
        RECT 638.400 433.050 639.450 449.100 ;
        RECT 644.400 448.350 645.600 449.100 ;
        RECT 650.400 448.350 651.600 450.600 ;
        RECT 643.950 445.950 646.050 448.050 ;
        RECT 646.950 445.950 649.050 448.050 ;
        RECT 649.950 445.950 652.050 448.050 ;
        RECT 647.400 444.900 648.600 445.650 ;
        RECT 656.400 445.050 657.450 494.100 ;
        RECT 665.400 493.350 666.600 494.100 ;
        RECT 671.400 493.350 672.600 494.100 ;
        RECT 676.950 493.950 679.050 496.050 ;
        RECT 685.950 494.100 688.050 496.200 ;
        RECT 691.950 494.100 694.050 496.200 ;
        RECT 700.950 494.100 703.050 496.200 ;
        RECT 661.950 490.950 664.050 493.050 ;
        RECT 664.950 490.950 667.050 493.050 ;
        RECT 667.950 490.950 670.050 493.050 ;
        RECT 670.950 490.950 673.050 493.050 ;
        RECT 662.400 488.400 663.600 490.650 ;
        RECT 668.400 489.900 669.600 490.650 ;
        RECT 662.400 475.050 663.450 488.400 ;
        RECT 667.950 487.800 670.050 489.900 ;
        RECT 664.950 484.950 667.050 487.050 ;
        RECT 661.950 472.950 664.050 475.050 ;
        RECT 665.400 450.600 666.450 484.950 ;
        RECT 677.400 481.050 678.450 493.950 ;
        RECT 686.400 493.350 687.600 494.100 ;
        RECT 682.950 490.950 685.050 493.050 ;
        RECT 685.950 490.950 688.050 493.050 ;
        RECT 683.400 489.900 684.600 490.650 ;
        RECT 682.950 487.800 685.050 489.900 ;
        RECT 676.950 478.950 679.050 481.050 ;
        RECT 692.400 471.450 693.450 494.100 ;
        RECT 701.400 493.350 702.600 494.100 ;
        RECT 697.950 490.950 700.050 493.050 ;
        RECT 700.950 490.950 703.050 493.050 ;
        RECT 698.400 489.000 699.600 490.650 ;
        RECT 707.400 490.050 708.450 511.950 ;
        RECT 713.400 508.050 714.450 535.950 ;
        RECT 736.950 532.950 739.050 535.050 ;
        RECT 715.950 527.100 718.050 529.200 ;
        RECT 724.950 527.100 727.050 529.200 ;
        RECT 730.950 527.100 733.050 529.200 ;
        RECT 716.400 517.050 717.450 527.100 ;
        RECT 725.400 526.350 726.600 527.100 ;
        RECT 731.400 526.350 732.600 527.100 ;
        RECT 721.950 523.950 724.050 526.050 ;
        RECT 724.950 523.950 727.050 526.050 ;
        RECT 727.950 523.950 730.050 526.050 ;
        RECT 730.950 523.950 733.050 526.050 ;
        RECT 722.400 521.400 723.600 523.650 ;
        RECT 728.400 522.900 729.600 523.650 ;
        RECT 737.400 523.050 738.450 532.950 ;
        RECT 742.950 527.100 745.050 529.200 ;
        RECT 749.400 529.050 750.450 547.950 ;
        RECT 743.400 526.350 744.600 527.100 ;
        RECT 748.950 526.950 751.050 529.050 ;
        RECT 742.950 523.950 745.050 526.050 ;
        RECT 745.950 523.950 748.050 526.050 ;
        RECT 715.950 514.950 718.050 517.050 ;
        RECT 722.400 514.050 723.450 521.400 ;
        RECT 727.950 520.800 730.050 522.900 ;
        RECT 736.950 520.950 739.050 523.050 ;
        RECT 746.400 521.400 747.600 523.650 ;
        RECT 746.400 517.050 747.450 521.400 ;
        RECT 748.950 520.950 751.050 523.050 ;
        RECT 727.950 514.950 730.050 517.050 ;
        RECT 745.950 514.950 748.050 517.050 ;
        RECT 721.950 511.950 724.050 514.050 ;
        RECT 712.950 505.950 715.050 508.050 ;
        RECT 721.950 505.950 724.050 508.050 ;
        RECT 715.950 495.000 718.050 499.050 ;
        RECT 722.400 495.600 723.450 505.950 ;
        RECT 716.400 493.350 717.600 495.000 ;
        RECT 722.400 493.350 723.600 495.600 ;
        RECT 712.950 490.950 715.050 493.050 ;
        RECT 715.950 490.950 718.050 493.050 ;
        RECT 718.950 490.950 721.050 493.050 ;
        RECT 721.950 490.950 724.050 493.050 ;
        RECT 697.950 484.950 700.050 489.000 ;
        RECT 703.950 484.950 706.050 490.050 ;
        RECT 706.950 487.950 709.050 490.050 ;
        RECT 713.400 488.400 714.600 490.650 ;
        RECT 719.400 489.900 720.600 490.650 ;
        RECT 713.400 484.050 714.450 488.400 ;
        RECT 718.950 487.800 721.050 489.900 ;
        RECT 724.950 484.950 727.050 489.900 ;
        RECT 728.400 484.050 729.450 514.950 ;
        RECT 733.950 508.950 736.050 511.050 ;
        RECT 730.950 493.950 733.050 499.050 ;
        RECT 734.400 495.600 735.450 508.950 ;
        RECT 749.400 507.450 750.450 520.950 ;
        RECT 752.400 520.050 753.450 551.400 ;
        RECT 760.950 544.950 763.050 547.050 ;
        RECT 761.400 535.050 762.450 544.950 ;
        RECT 760.950 532.950 763.050 535.050 ;
        RECT 761.400 528.600 762.450 532.950 ;
        RECT 764.400 532.050 765.450 565.800 ;
        RECT 767.400 562.050 768.450 595.950 ;
        RECT 776.400 580.050 777.450 599.400 ;
        RECT 785.400 589.050 786.450 607.950 ;
        RECT 788.400 606.450 789.450 616.950 ;
        RECT 791.400 616.050 792.450 644.400 ;
        RECT 797.400 640.050 798.450 649.950 ;
        RECT 803.400 649.350 804.600 650.100 ;
        RECT 809.400 649.350 810.600 651.600 ;
        RECT 815.400 649.350 816.600 651.600 ;
        RECT 802.950 646.950 805.050 649.050 ;
        RECT 805.950 646.950 808.050 649.050 ;
        RECT 808.950 646.950 811.050 649.050 ;
        RECT 811.950 646.950 814.050 649.050 ;
        RECT 814.950 646.950 817.050 649.050 ;
        RECT 820.950 646.950 823.050 649.050 ;
        RECT 806.400 644.400 807.600 646.650 ;
        RECT 812.400 645.000 813.600 646.650 ;
        RECT 802.950 640.950 805.050 643.050 ;
        RECT 796.950 637.950 799.050 640.050 ;
        RECT 803.400 634.050 804.450 640.950 ;
        RECT 802.950 631.950 805.050 634.050 ;
        RECT 790.950 613.950 793.050 616.050 ;
        RECT 791.400 606.450 792.600 606.600 ;
        RECT 788.400 605.400 792.600 606.450 ;
        RECT 791.400 604.350 792.600 605.400 ;
        RECT 796.950 605.100 799.050 607.200 ;
        RECT 803.400 607.050 804.450 631.950 ;
        RECT 797.400 604.350 798.600 605.100 ;
        RECT 802.950 604.950 805.050 607.050 ;
        RECT 790.950 601.950 793.050 604.050 ;
        RECT 793.950 601.950 796.050 604.050 ;
        RECT 796.950 601.950 799.050 604.050 ;
        RECT 799.950 601.950 802.050 604.050 ;
        RECT 794.400 600.900 795.600 601.650 ;
        RECT 800.400 601.050 801.600 601.650 ;
        RECT 793.950 598.800 796.050 600.900 ;
        RECT 800.400 600.000 805.050 601.050 ;
        RECT 799.950 598.950 805.050 600.000 ;
        RECT 806.400 600.450 807.450 644.400 ;
        RECT 811.950 640.950 814.050 645.000 ;
        RECT 817.950 643.950 820.050 646.050 ;
        RECT 821.400 644.400 822.600 646.650 ;
        RECT 808.950 639.450 811.050 640.050 ;
        RECT 814.950 639.450 817.050 640.050 ;
        RECT 808.950 638.400 817.050 639.450 ;
        RECT 808.950 637.950 811.050 638.400 ;
        RECT 814.950 637.950 817.050 638.400 ;
        RECT 808.950 607.050 811.050 607.200 ;
        RECT 818.400 607.050 819.450 643.950 ;
        RECT 821.400 622.050 822.450 644.400 ;
        RECT 825.150 638.700 826.350 657.300 ;
        RECT 833.400 652.050 834.450 664.950 ;
        RECT 832.950 649.950 835.050 652.050 ;
        RECT 830.100 646.950 832.200 649.050 ;
        RECT 830.400 645.000 831.600 646.650 ;
        RECT 836.400 645.450 837.450 667.950 ;
        RECT 829.950 640.950 832.050 645.000 ;
        RECT 833.400 644.400 837.450 645.450 ;
        RECT 825.150 637.500 829.350 638.700 ;
        RECT 827.250 636.600 829.350 637.500 ;
        RECT 820.950 619.950 823.050 622.050 ;
        RECT 808.950 606.600 813.000 607.050 ;
        RECT 808.950 605.100 813.600 606.600 ;
        RECT 810.000 604.950 813.600 605.100 ;
        RECT 817.950 604.950 820.050 607.050 ;
        RECT 821.400 606.600 822.450 619.950 ;
        RECT 827.250 613.500 829.350 614.400 ;
        RECT 825.150 612.300 829.350 613.500 ;
        RECT 812.400 604.350 813.600 604.950 ;
        RECT 821.400 604.350 822.600 606.600 ;
        RECT 811.950 601.950 814.050 604.050 ;
        RECT 814.950 601.950 817.050 604.050 ;
        RECT 820.950 601.950 823.050 604.050 ;
        RECT 815.400 600.900 816.600 601.650 ;
        RECT 806.400 599.400 810.450 600.450 ;
        RECT 799.950 595.950 802.050 598.950 ;
        RECT 805.950 595.950 808.050 598.050 ;
        RECT 784.950 586.950 787.050 589.050 ;
        RECT 802.950 586.950 805.050 589.050 ;
        RECT 787.950 580.950 790.050 583.050 ;
        RECT 775.950 577.950 778.050 580.050 ;
        RECT 784.950 577.950 787.050 580.050 ;
        RECT 769.950 572.100 772.050 574.200 ;
        RECT 778.950 572.100 781.050 574.200 ;
        RECT 766.950 559.950 769.050 562.050 ;
        RECT 767.400 550.050 768.450 559.950 ;
        RECT 766.950 547.950 769.050 550.050 ;
        RECT 766.950 540.450 769.050 541.050 ;
        RECT 770.400 540.450 771.450 572.100 ;
        RECT 779.400 571.350 780.600 572.100 ;
        RECT 773.100 568.950 775.200 571.050 ;
        RECT 778.500 568.950 780.600 571.050 ;
        RECT 781.800 568.950 783.900 571.050 ;
        RECT 773.400 567.900 774.600 568.650 ;
        RECT 772.950 565.800 775.050 567.900 ;
        RECT 782.400 567.450 783.600 568.650 ;
        RECT 785.400 567.450 786.450 577.950 ;
        RECT 782.400 566.400 786.450 567.450 ;
        RECT 788.400 567.450 789.450 580.950 ;
        RECT 796.950 572.100 799.050 574.200 ;
        RECT 803.400 573.600 804.450 586.950 ;
        RECT 806.400 574.050 807.450 595.950 ;
        RECT 797.400 571.350 798.600 572.100 ;
        RECT 803.400 571.350 804.600 573.600 ;
        RECT 805.950 571.950 808.050 574.050 ;
        RECT 793.950 568.950 796.050 571.050 ;
        RECT 796.950 568.950 799.050 571.050 ;
        RECT 799.950 568.950 802.050 571.050 ;
        RECT 802.950 568.950 805.050 571.050 ;
        RECT 794.400 567.450 795.600 568.650 ;
        RECT 788.400 566.400 795.600 567.450 ;
        RECT 800.400 566.400 801.600 568.650 ;
        RECT 772.950 559.950 775.050 562.050 ;
        RECT 766.950 539.400 771.450 540.450 ;
        RECT 766.950 538.950 769.050 539.400 ;
        RECT 763.950 529.950 766.050 532.050 ;
        RECT 767.400 528.600 768.450 538.950 ;
        RECT 761.400 526.350 762.600 528.600 ;
        RECT 767.400 526.350 768.600 528.600 ;
        RECT 757.950 523.950 760.050 526.050 ;
        RECT 760.950 523.950 763.050 526.050 ;
        RECT 763.950 523.950 766.050 526.050 ;
        RECT 766.950 523.950 769.050 526.050 ;
        RECT 758.400 522.000 759.600 523.650 ;
        RECT 764.400 522.900 765.600 523.650 ;
        RECT 751.950 517.950 754.050 520.050 ;
        RECT 757.950 517.950 760.050 522.000 ;
        RECT 763.950 520.800 766.050 522.900 ;
        RECT 769.950 519.450 772.050 523.050 ;
        RECT 767.400 519.000 772.050 519.450 ;
        RECT 767.400 518.400 771.450 519.000 ;
        RECT 749.400 506.400 753.450 507.450 ;
        RECT 734.400 493.350 735.600 495.600 ;
        RECT 739.950 495.000 742.050 499.050 ;
        RECT 740.400 493.350 741.600 495.000 ;
        RECT 748.950 494.100 751.050 496.200 ;
        RECT 733.950 490.950 736.050 493.050 ;
        RECT 736.950 490.950 739.050 493.050 ;
        RECT 739.950 490.950 742.050 493.050 ;
        RECT 742.950 490.950 745.050 493.050 ;
        RECT 737.400 489.900 738.600 490.650 ;
        RECT 736.950 487.800 739.050 489.900 ;
        RECT 743.400 489.000 744.600 490.650 ;
        RECT 742.950 484.950 745.050 489.000 ;
        RECT 712.950 481.950 715.050 484.050 ;
        RECT 727.950 481.950 730.050 484.050 ;
        RECT 692.400 470.400 696.450 471.450 ;
        RECT 679.950 460.950 682.050 463.050 ;
        RECT 680.400 450.600 681.450 460.950 ;
        RECT 691.950 454.950 694.050 457.050 ;
        RECT 665.400 448.350 666.600 450.600 ;
        RECT 680.400 448.350 681.600 450.600 ;
        RECT 689.400 450.450 690.600 450.600 ;
        RECT 692.400 450.450 693.450 454.950 ;
        RECT 689.400 449.400 693.450 450.450 ;
        RECT 689.400 448.350 690.600 449.400 ;
        RECT 661.950 445.950 664.050 448.050 ;
        RECT 664.950 445.950 667.050 448.050 ;
        RECT 667.950 445.950 670.050 448.050 ;
        RECT 680.100 445.950 682.200 448.050 ;
        RECT 683.400 445.950 685.500 448.050 ;
        RECT 688.800 445.950 690.900 448.050 ;
        RECT 691.950 445.950 694.050 448.050 ;
        RECT 646.950 442.800 649.050 444.900 ;
        RECT 655.950 442.950 658.050 445.050 ;
        RECT 662.400 444.900 663.600 445.650 ;
        RECT 668.400 444.900 669.600 445.650 ;
        RECT 683.400 444.900 684.600 445.650 ;
        RECT 661.950 442.800 664.050 444.900 ;
        RECT 667.950 442.800 670.050 444.900 ;
        RECT 682.950 442.800 685.050 444.900 ;
        RECT 628.950 430.950 631.050 433.050 ;
        RECT 637.950 430.950 640.050 433.050 ;
        RECT 655.950 424.950 658.050 427.050 ;
        RECT 598.950 423.450 601.050 424.050 ;
        RECT 598.950 422.400 606.450 423.450 ;
        RECT 598.950 421.950 601.050 422.400 ;
        RECT 601.950 417.000 604.050 421.050 ;
        RECT 605.400 420.450 606.450 422.400 ;
        RECT 656.400 421.050 657.450 424.950 ;
        RECT 605.400 419.400 609.450 420.450 ;
        RECT 608.400 417.600 609.450 419.400 ;
        RECT 634.950 418.950 637.050 421.050 ;
        RECT 649.950 418.950 652.050 421.050 ;
        RECT 602.400 415.350 603.600 417.000 ;
        RECT 608.400 415.350 609.600 417.600 ;
        RECT 616.950 415.950 619.050 418.050 ;
        RECT 625.950 416.100 628.050 418.200 ;
        RECT 601.950 412.950 604.050 415.050 ;
        RECT 604.950 412.950 607.050 415.050 ;
        RECT 607.950 412.950 610.050 415.050 ;
        RECT 610.950 412.950 613.050 415.050 ;
        RECT 605.400 411.900 606.600 412.650 ;
        RECT 604.950 409.800 607.050 411.900 ;
        RECT 611.400 411.000 612.600 412.650 ;
        RECT 595.950 406.950 598.050 409.050 ;
        RECT 592.950 397.950 595.050 400.050 ;
        RECT 605.400 394.050 606.450 409.800 ;
        RECT 607.950 406.950 610.050 409.050 ;
        RECT 610.950 406.950 613.050 411.000 ;
        RECT 617.400 409.050 618.450 415.950 ;
        RECT 626.400 415.350 627.600 416.100 ;
        RECT 622.950 412.950 625.050 415.050 ;
        RECT 625.950 412.950 628.050 415.050 ;
        RECT 628.950 412.950 631.050 415.050 ;
        RECT 623.400 411.900 624.600 412.650 ;
        RECT 622.950 409.800 625.050 411.900 ;
        RECT 616.950 406.950 619.050 409.050 ;
        RECT 608.400 400.050 609.450 406.950 ;
        RECT 613.950 403.950 616.050 406.050 ;
        RECT 607.800 397.950 609.900 400.050 ;
        RECT 610.950 397.950 613.050 400.050 ;
        RECT 604.950 391.950 607.050 394.050 ;
        RECT 592.950 379.950 595.050 382.050 ;
        RECT 556.950 367.950 559.050 370.050 ;
        RECT 559.950 367.950 562.050 370.050 ;
        RECT 562.950 367.950 565.050 370.050 ;
        RECT 560.400 366.900 561.600 367.650 ;
        RECT 572.400 367.050 573.450 371.100 ;
        RECT 578.400 370.350 579.600 371.100 ;
        RECT 584.400 370.350 585.600 372.000 ;
        RECT 589.950 370.950 592.050 373.050 ;
        RECT 593.400 372.600 594.450 379.950 ;
        RECT 599.250 379.500 601.350 380.400 ;
        RECT 597.150 378.300 601.350 379.500 ;
        RECT 593.400 370.350 594.600 372.600 ;
        RECT 577.950 367.950 580.050 370.050 ;
        RECT 580.950 367.950 583.050 370.050 ;
        RECT 583.950 367.950 586.050 370.050 ;
        RECT 586.950 367.950 589.050 370.050 ;
        RECT 592.950 367.950 595.050 370.050 ;
        RECT 559.950 364.800 562.050 366.900 ;
        RECT 571.800 364.950 573.900 367.050 ;
        RECT 574.950 363.450 577.050 367.050 ;
        RECT 581.400 366.000 582.600 367.650 ;
        RECT 587.400 366.450 588.600 367.650 ;
        RECT 589.950 366.450 592.050 367.050 ;
        RECT 572.400 363.000 577.050 363.450 ;
        RECT 572.400 362.400 576.450 363.000 ;
        RECT 562.950 349.950 565.050 352.050 ;
        RECT 541.950 343.950 544.050 346.050 ;
        RECT 550.950 343.950 553.050 346.050 ;
        RECT 532.950 340.950 535.050 343.050 ;
        RECT 538.950 342.450 543.000 343.050 ;
        RECT 538.950 340.950 543.450 342.450 ;
        RECT 518.400 337.350 519.600 338.100 ;
        RECT 524.400 337.350 525.600 339.600 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 517.950 334.950 520.050 337.050 ;
        RECT 520.950 334.950 523.050 337.050 ;
        RECT 523.950 334.950 526.050 337.050 ;
        RECT 526.950 334.950 529.050 337.050 ;
        RECT 512.400 332.400 516.450 333.450 ;
        RECT 521.400 333.000 522.600 334.650 ;
        RECT 527.400 333.900 528.600 334.650 ;
        RECT 508.950 328.950 511.050 331.050 ;
        RECT 511.950 328.950 514.050 331.050 ;
        RECT 496.650 325.500 500.850 326.700 ;
        RECT 502.950 325.950 505.050 328.050 ;
        RECT 496.650 324.600 498.750 325.500 ;
        RECT 491.400 320.400 495.450 321.450 ;
        RECT 482.400 305.400 486.450 306.450 ;
        RECT 460.950 298.950 463.050 301.050 ;
        RECT 449.400 292.350 450.600 294.600 ;
        RECT 457.950 292.950 460.050 295.050 ;
        RECT 448.950 289.950 451.050 292.050 ;
        RECT 451.950 289.950 454.050 292.050 ;
        RECT 454.950 289.950 457.050 292.050 ;
        RECT 445.950 286.950 448.050 289.050 ;
        RECT 452.400 287.400 453.600 289.650 ;
        RECT 461.400 288.900 462.450 298.950 ;
        RECT 469.950 293.100 472.050 295.200 ;
        RECT 476.400 294.600 477.450 304.950 ;
        RECT 482.400 294.600 483.450 305.400 ;
        RECT 487.950 304.950 490.050 307.050 ;
        RECT 488.250 301.500 490.350 302.400 ;
        RECT 486.150 300.300 490.350 301.500 ;
        RECT 470.400 292.350 471.600 293.100 ;
        RECT 476.400 292.350 477.600 294.600 ;
        RECT 482.400 292.350 483.600 294.600 ;
        RECT 466.950 289.950 469.050 292.050 ;
        RECT 469.950 289.950 472.050 292.050 ;
        RECT 472.950 289.950 475.050 292.050 ;
        RECT 475.950 289.950 478.050 292.050 ;
        RECT 481.950 289.950 484.050 292.050 ;
        RECT 467.400 288.900 468.600 289.650 ;
        RECT 427.950 274.950 430.050 277.050 ;
        RECT 442.950 274.950 445.050 277.050 ;
        RECT 421.950 268.950 424.050 271.050 ;
        RECT 428.400 265.050 429.450 274.950 ;
        RECT 442.950 268.950 445.050 271.050 ;
        RECT 427.950 262.950 430.050 265.050 ;
        RECT 388.950 256.950 391.050 259.050 ;
        RECT 391.950 256.950 394.050 259.050 ;
        RECT 394.950 256.950 397.050 259.050 ;
        RECT 397.950 256.950 400.050 259.050 ;
        RECT 385.950 253.950 388.050 256.050 ;
        RECT 389.400 255.900 390.600 256.650 ;
        RECT 382.950 232.950 385.050 235.050 ;
        RECT 368.400 218.400 372.450 219.450 ;
        RECT 364.950 214.950 367.050 217.050 ;
        RECT 371.400 216.600 372.450 218.400 ;
        RECT 373.950 217.950 376.050 220.050 ;
        RECT 371.400 214.350 372.600 216.600 ;
        RECT 376.950 215.100 379.050 217.200 ;
        RECT 382.950 215.100 385.050 217.200 ;
        RECT 386.400 217.050 387.450 253.950 ;
        RECT 388.950 253.800 391.050 255.900 ;
        RECT 395.400 254.400 396.600 256.650 ;
        RECT 395.400 250.050 396.450 254.400 ;
        RECT 397.950 250.950 400.050 253.050 ;
        RECT 394.950 247.950 397.050 250.050 ;
        RECT 398.400 220.050 399.450 250.950 ;
        RECT 404.400 250.050 405.450 259.950 ;
        RECT 413.400 259.350 414.600 260.100 ;
        RECT 419.400 259.950 424.050 262.050 ;
        RECT 419.400 259.350 420.600 259.950 ;
        RECT 409.950 256.950 412.050 259.050 ;
        RECT 412.950 256.950 415.050 259.050 ;
        RECT 415.950 256.950 418.050 259.050 ;
        RECT 418.950 256.950 421.050 259.050 ;
        RECT 431.100 256.950 433.200 259.050 ;
        RECT 436.500 256.950 438.600 259.050 ;
        RECT 439.800 256.950 441.900 259.050 ;
        RECT 410.400 254.400 411.600 256.650 ;
        RECT 416.400 254.400 417.600 256.650 ;
        RECT 410.400 250.050 411.450 254.400 ;
        RECT 403.950 247.950 406.050 250.050 ;
        RECT 409.950 247.950 412.050 250.050 ;
        RECT 412.950 244.950 415.050 247.050 ;
        RECT 406.950 235.950 409.050 238.050 ;
        RECT 407.400 229.050 408.450 235.950 ;
        RECT 406.950 226.950 409.050 229.050 ;
        RECT 400.950 223.950 403.050 226.050 ;
        RECT 377.400 214.350 378.600 215.100 ;
        RECT 367.950 211.950 370.050 214.050 ;
        RECT 370.950 211.950 373.050 214.050 ;
        RECT 373.950 211.950 376.050 214.050 ;
        RECT 376.950 211.950 379.050 214.050 ;
        RECT 364.950 208.950 367.050 211.050 ;
        RECT 368.400 209.400 369.600 211.650 ;
        RECT 374.400 210.900 375.600 211.650 ;
        RECT 352.950 193.950 355.050 196.050 ;
        RECT 358.950 193.950 361.050 196.050 ;
        RECT 343.950 187.950 346.050 190.050 ;
        RECT 349.950 187.950 352.050 190.050 ;
        RECT 329.400 181.350 330.600 182.100 ;
        RECT 334.950 181.950 337.050 184.050 ;
        RECT 340.950 182.100 343.050 187.050 ;
        RECT 344.400 183.600 345.450 187.950 ;
        RECT 353.400 187.050 354.450 193.950 ;
        RECT 361.950 190.950 364.050 193.050 ;
        RECT 352.950 184.950 355.050 187.050 ;
        RECT 344.400 181.350 345.600 183.600 ;
        RECT 349.950 182.100 352.050 184.200 ;
        RECT 350.400 181.350 351.600 182.100 ;
        RECT 325.950 178.950 328.050 181.050 ;
        RECT 328.950 178.950 331.050 181.050 ;
        RECT 331.950 178.950 334.050 181.050 ;
        RECT 343.950 178.950 346.050 181.050 ;
        RECT 346.950 178.950 349.050 181.050 ;
        RECT 349.950 178.950 352.050 181.050 ;
        RECT 352.950 178.950 355.050 181.050 ;
        RECT 320.400 176.400 324.450 177.450 ;
        RECT 326.400 177.000 327.600 178.650 ;
        RECT 332.400 177.900 333.600 178.650 ;
        RECT 319.950 166.950 322.050 169.050 ;
        RECT 320.400 154.050 321.450 166.950 ;
        RECT 316.800 151.950 318.900 154.050 ;
        RECT 319.950 151.950 322.050 154.050 ;
        RECT 313.950 142.950 316.050 145.050 ;
        RECT 323.400 142.050 324.450 176.400 ;
        RECT 325.950 172.950 328.050 177.000 ;
        RECT 331.950 175.800 334.050 177.900 ;
        RECT 334.950 175.950 337.050 178.050 ;
        RECT 347.400 177.900 348.600 178.650 ;
        RECT 332.400 172.050 333.450 175.800 ;
        RECT 325.950 169.800 328.050 171.900 ;
        RECT 331.950 169.950 334.050 172.050 ;
        RECT 326.400 151.050 327.450 169.800 ;
        RECT 335.400 169.050 336.450 175.950 ;
        RECT 346.950 175.800 349.050 177.900 ;
        RECT 353.400 177.000 354.600 178.650 ;
        RECT 352.950 169.950 355.050 177.000 ;
        RECT 362.400 175.050 363.450 190.950 ;
        RECT 365.400 183.600 366.450 208.950 ;
        RECT 368.400 193.050 369.450 209.400 ;
        RECT 373.950 208.800 376.050 210.900 ;
        RECT 379.950 208.950 382.050 211.050 ;
        RECT 380.400 202.050 381.450 208.950 ;
        RECT 383.400 205.050 384.450 215.100 ;
        RECT 385.950 214.950 388.050 217.050 ;
        RECT 388.950 215.100 391.050 217.200 ;
        RECT 394.950 216.000 397.050 220.050 ;
        RECT 397.950 217.950 400.050 220.050 ;
        RECT 401.400 217.050 402.450 223.950 ;
        RECT 409.950 219.450 412.050 220.050 ;
        RECT 413.400 219.450 414.450 244.950 ;
        RECT 416.400 220.050 417.450 254.400 ;
        RECT 421.950 253.950 424.050 256.050 ;
        RECT 431.400 255.000 432.600 256.650 ;
        RECT 418.950 250.950 421.050 253.050 ;
        RECT 419.400 226.050 420.450 250.950 ;
        RECT 422.400 244.050 423.450 253.950 ;
        RECT 430.950 250.950 433.050 255.000 ;
        RECT 440.400 254.400 441.600 256.650 ;
        RECT 431.400 247.050 432.450 250.950 ;
        RECT 440.400 250.050 441.450 254.400 ;
        RECT 439.950 247.950 442.050 250.050 ;
        RECT 430.950 244.950 433.050 247.050 ;
        RECT 421.950 241.950 424.050 244.050 ;
        RECT 443.400 235.050 444.450 268.950 ;
        RECT 446.400 241.050 447.450 286.950 ;
        RECT 452.400 264.450 453.450 287.400 ;
        RECT 460.950 286.800 463.050 288.900 ;
        RECT 466.950 286.800 469.050 288.900 ;
        RECT 473.400 288.000 474.600 289.650 ;
        RECT 472.950 283.950 475.050 288.000 ;
        RECT 478.950 286.950 481.050 289.050 ;
        RECT 472.950 280.800 475.050 282.900 ;
        RECT 457.950 277.950 460.050 280.050 ;
        RECT 458.400 274.050 459.450 277.950 ;
        RECT 457.950 271.950 460.050 274.050 ;
        RECT 452.400 263.400 456.450 264.450 ;
        RECT 455.400 262.200 456.450 263.400 ;
        RECT 454.950 260.100 457.050 262.200 ;
        RECT 460.950 260.100 463.050 262.200 ;
        RECT 466.950 260.100 469.050 262.200 ;
        RECT 473.400 261.600 474.450 280.800 ;
        RECT 479.400 274.050 480.450 286.950 ;
        RECT 486.150 281.700 487.350 300.300 ;
        RECT 490.800 293.100 492.900 295.200 ;
        RECT 494.400 295.050 495.450 320.400 ;
        RECT 512.400 319.050 513.450 328.950 ;
        RECT 499.950 316.950 502.050 319.050 ;
        RECT 511.950 316.950 514.050 319.050 ;
        RECT 496.950 313.950 499.050 316.050 ;
        RECT 491.400 292.350 492.600 293.100 ;
        RECT 493.950 292.950 496.050 295.050 ;
        RECT 491.100 289.950 493.200 292.050 ;
        RECT 493.950 286.950 496.050 289.050 ;
        RECT 485.850 279.600 487.950 281.700 ;
        RECT 490.950 280.950 493.050 283.050 ;
        RECT 481.950 274.950 484.050 277.050 ;
        RECT 478.950 271.950 481.050 274.050 ;
        RECT 479.400 262.200 480.450 271.950 ;
        RECT 455.400 259.350 456.600 260.100 ;
        RECT 451.950 256.950 454.050 259.050 ;
        RECT 454.950 256.950 457.050 259.050 ;
        RECT 452.400 254.400 453.600 256.650 ;
        RECT 448.950 250.950 451.050 253.050 ;
        RECT 445.950 238.950 448.050 241.050 ;
        RECT 421.950 232.950 424.050 235.050 ;
        RECT 442.950 232.950 445.050 235.050 ;
        RECT 418.950 223.950 421.050 226.050 ;
        RECT 409.950 218.400 414.450 219.450 ;
        RECT 409.950 217.950 412.050 218.400 ;
        RECT 415.950 217.950 418.050 220.050 ;
        RECT 389.400 214.350 390.600 215.100 ;
        RECT 395.400 214.350 396.600 216.000 ;
        RECT 400.950 214.950 403.050 217.050 ;
        RECT 410.400 216.600 411.450 217.950 ;
        RECT 410.400 214.350 411.600 216.600 ;
        RECT 388.950 211.950 391.050 214.050 ;
        RECT 391.950 211.950 394.050 214.050 ;
        RECT 394.950 211.950 397.050 214.050 ;
        RECT 397.950 211.950 400.050 214.050 ;
        RECT 409.950 211.950 412.050 214.050 ;
        RECT 412.950 211.950 415.050 214.050 ;
        RECT 415.950 211.950 418.050 214.050 ;
        RECT 385.950 207.450 388.050 211.050 ;
        RECT 392.400 209.400 393.600 211.650 ;
        RECT 398.400 210.900 399.600 211.650 ;
        RECT 385.950 207.000 390.450 207.450 ;
        RECT 386.400 206.400 390.450 207.000 ;
        RECT 382.950 202.950 385.050 205.050 ;
        RECT 379.950 199.950 382.050 202.050 ;
        RECT 373.950 193.950 376.050 196.050 ;
        RECT 367.950 190.950 370.050 193.050 ;
        RECT 365.400 181.350 366.600 183.600 ;
        RECT 365.400 178.950 367.500 181.050 ;
        RECT 370.800 178.950 372.900 181.050 ;
        RECT 361.950 172.950 364.050 175.050 ;
        RECT 328.950 166.950 331.050 169.050 ;
        RECT 334.950 166.950 337.050 169.050 ;
        RECT 325.950 148.950 328.050 151.050 ;
        RECT 322.950 139.950 325.050 142.050 ;
        RECT 319.950 137.100 322.050 139.200 ;
        RECT 320.400 136.350 321.600 137.100 ;
        RECT 316.950 133.950 319.050 136.050 ;
        RECT 319.950 133.950 322.050 136.050 ;
        RECT 322.950 133.950 325.050 136.050 ;
        RECT 317.400 132.450 318.600 133.650 ;
        RECT 311.400 131.400 318.600 132.450 ;
        RECT 323.400 131.400 324.600 133.650 ;
        RECT 280.950 115.950 283.050 118.050 ;
        RECT 280.950 112.800 283.050 114.900 ;
        RECT 277.950 103.950 280.050 106.050 ;
        RECT 281.400 105.600 282.450 112.800 ;
        RECT 290.400 112.050 291.450 130.800 ;
        RECT 305.400 121.050 306.450 131.400 ;
        RECT 304.950 118.950 307.050 121.050 ;
        RECT 292.950 115.950 295.050 118.050 ;
        RECT 289.950 109.950 292.050 112.050 ;
        RECT 281.400 103.350 282.600 105.600 ;
        RECT 286.950 104.100 289.050 106.200 ;
        RECT 293.400 106.050 294.450 115.950 ;
        RECT 295.950 112.950 298.050 115.050 ;
        RECT 287.400 103.350 288.600 104.100 ;
        RECT 292.950 103.950 295.050 106.050 ;
        RECT 280.950 100.950 283.050 103.050 ;
        RECT 283.950 100.950 286.050 103.050 ;
        RECT 286.950 100.950 289.050 103.050 ;
        RECT 289.950 100.950 292.050 103.050 ;
        RECT 277.950 97.950 280.050 100.050 ;
        RECT 284.400 98.400 285.600 100.650 ;
        RECT 290.400 99.900 291.600 100.650 ;
        RECT 274.950 94.950 277.050 97.050 ;
        RECT 272.400 92.400 276.450 93.450 ;
        RECT 271.950 88.950 274.050 91.050 ;
        RECT 268.950 85.950 271.050 88.050 ;
        RECT 272.400 70.050 273.450 88.950 ;
        RECT 271.950 67.950 274.050 70.050 ;
        RECT 271.950 59.100 274.050 61.200 ;
        RECT 275.400 61.050 276.450 92.400 ;
        RECT 278.400 88.050 279.450 97.950 ;
        RECT 284.400 94.050 285.450 98.400 ;
        RECT 289.950 97.800 292.050 99.900 ;
        RECT 292.950 97.950 295.050 100.050 ;
        RECT 296.400 99.900 297.450 112.950 ;
        RECT 298.950 105.600 303.000 106.050 ;
        RECT 298.950 103.950 303.600 105.600 ;
        RECT 307.950 105.000 310.050 109.050 ;
        RECT 314.400 106.050 315.450 131.400 ;
        RECT 316.950 127.950 319.050 130.050 ;
        RECT 302.400 103.350 303.600 103.950 ;
        RECT 308.400 103.350 309.600 105.000 ;
        RECT 313.950 103.950 316.050 106.050 ;
        RECT 301.950 100.950 304.050 103.050 ;
        RECT 304.950 100.950 307.050 103.050 ;
        RECT 307.950 100.950 310.050 103.050 ;
        RECT 310.950 100.950 313.050 103.050 ;
        RECT 305.400 99.900 306.600 100.650 ;
        RECT 283.950 91.950 286.050 94.050 ;
        RECT 277.950 85.950 280.050 88.050 ;
        RECT 293.400 79.050 294.450 97.950 ;
        RECT 295.950 97.800 298.050 99.900 ;
        RECT 304.950 97.800 307.050 99.900 ;
        RECT 311.400 99.000 312.600 100.650 ;
        RECT 310.950 94.950 313.050 99.000 ;
        RECT 292.950 76.950 295.050 79.050 ;
        RECT 283.950 73.950 286.050 76.050 ;
        RECT 277.950 64.950 280.050 67.050 ;
        RECT 272.400 58.350 273.600 59.100 ;
        RECT 274.950 58.950 277.050 61.050 ;
        RECT 268.950 55.950 271.050 58.050 ;
        RECT 271.950 55.950 274.050 58.050 ;
        RECT 269.400 54.900 270.600 55.650 ;
        RECT 260.400 53.400 264.450 54.450 ;
        RECT 248.400 49.050 249.450 53.400 ;
        RECT 254.400 49.050 255.450 53.400 ;
        RECT 241.950 46.950 244.050 49.050 ;
        RECT 247.950 46.950 250.050 49.050 ;
        RECT 253.950 46.950 256.050 49.050 ;
        RECT 229.950 37.950 232.050 40.050 ;
        RECT 244.950 34.950 247.050 37.050 ;
        RECT 229.950 31.950 232.050 34.050 ;
        RECT 230.400 31.200 231.600 31.950 ;
        RECT 220.950 28.950 223.050 31.050 ;
        RECT 226.500 29.100 228.600 31.200 ;
        RECT 224.400 27.450 225.600 27.600 ;
        RECT 218.400 26.400 225.600 27.450 ;
        RECT 212.400 25.350 213.600 26.100 ;
        RECT 205.950 22.950 208.050 25.050 ;
        RECT 208.950 22.950 211.050 25.050 ;
        RECT 211.950 22.950 214.050 25.050 ;
        RECT 187.950 19.800 190.050 21.900 ;
        RECT 193.950 19.800 196.050 21.900 ;
        RECT 199.950 19.950 202.050 22.050 ;
        RECT 209.400 21.900 210.600 22.650 ;
        RECT 208.950 19.800 211.050 21.900 ;
        RECT 214.950 16.950 217.050 19.050 ;
        RECT 85.950 13.950 88.050 16.050 ;
        RECT 100.950 13.950 103.050 16.050 ;
        RECT 106.950 14.400 111.450 16.050 ;
        RECT 106.950 13.950 111.000 14.400 ;
        RECT 121.950 13.950 124.050 16.050 ;
        RECT 215.400 7.050 216.450 16.950 ;
        RECT 221.400 7.050 222.450 26.400 ;
        RECT 224.400 25.350 225.600 26.400 ;
        RECT 224.100 22.950 226.200 25.050 ;
        RECT 227.100 24.000 228.000 29.100 ;
        RECT 229.800 28.800 231.900 30.900 ;
        RECT 236.400 29.400 238.500 31.500 ;
        RECT 234.000 27.000 236.100 27.900 ;
        RECT 228.900 25.800 236.100 27.000 ;
        RECT 228.900 24.900 231.000 25.800 ;
        RECT 234.000 24.000 236.100 24.900 ;
        RECT 227.100 23.100 236.100 24.000 ;
        RECT 227.100 16.500 228.000 23.100 ;
        RECT 234.000 22.800 236.100 23.100 ;
        RECT 229.800 19.950 231.900 22.050 ;
        RECT 230.400 17.400 231.600 19.650 ;
        RECT 237.000 16.800 237.900 29.400 ;
        RECT 241.950 28.950 244.050 31.050 ;
        RECT 238.800 22.950 240.900 25.050 ;
        RECT 239.400 21.450 240.600 22.650 ;
        RECT 242.400 21.900 243.450 28.950 ;
        RECT 241.950 21.450 244.050 21.900 ;
        RECT 239.400 20.400 244.050 21.450 ;
        RECT 241.950 19.800 244.050 20.400 ;
        RECT 227.100 14.400 229.200 16.500 ;
        RECT 236.100 14.700 238.200 16.800 ;
        RECT 245.400 13.050 246.450 34.950 ;
        RECT 247.950 26.100 250.050 28.200 ;
        RECT 253.950 26.100 256.050 28.200 ;
        RECT 260.400 27.600 261.450 53.400 ;
        RECT 268.950 52.800 271.050 54.900 ;
        RECT 274.950 52.950 277.050 55.050 ;
        RECT 278.400 54.900 279.450 64.950 ;
        RECT 284.400 60.600 285.450 73.950 ;
        RECT 317.400 73.050 318.450 127.950 ;
        RECT 319.950 118.950 322.050 121.050 ;
        RECT 320.400 106.050 321.450 118.950 ;
        RECT 323.400 115.050 324.450 131.400 ;
        RECT 325.950 130.950 328.050 133.050 ;
        RECT 322.950 112.950 325.050 115.050 ;
        RECT 326.400 109.050 327.450 130.950 ;
        RECT 329.400 124.050 330.450 166.950 ;
        RECT 352.950 166.800 355.050 168.900 ;
        RECT 345.000 165.450 349.050 166.050 ;
        RECT 344.400 163.950 349.050 165.450 ;
        RECT 334.950 154.950 337.050 157.050 ;
        RECT 335.400 139.200 336.450 154.950 ;
        RECT 334.950 137.100 337.050 139.200 ;
        RECT 344.400 139.050 345.450 163.950 ;
        RECT 349.950 160.950 352.050 163.050 ;
        RECT 350.400 154.050 351.450 160.950 ;
        RECT 353.400 157.050 354.450 166.800 ;
        RECT 374.400 157.050 375.450 193.950 ;
        RECT 389.400 183.600 390.450 206.400 ;
        RECT 392.400 202.050 393.450 209.400 ;
        RECT 397.950 208.800 400.050 210.900 ;
        RECT 413.400 209.400 414.600 211.650 ;
        RECT 391.950 199.950 394.050 202.050 ;
        RECT 391.950 187.950 394.050 190.050 ;
        RECT 389.400 181.350 390.600 183.600 ;
        RECT 383.100 178.950 385.200 181.050 ;
        RECT 388.500 178.950 390.600 181.050 ;
        RECT 388.950 166.950 391.050 169.050 ;
        RECT 376.950 157.950 379.050 160.050 ;
        RECT 352.950 154.950 355.050 157.050 ;
        RECT 365.400 156.000 372.450 156.450 ;
        RECT 365.400 155.400 373.050 156.000 ;
        RECT 349.800 151.950 351.900 154.050 ;
        RECT 352.950 151.800 355.050 153.900 ;
        RECT 349.950 148.800 352.050 150.900 ;
        RECT 350.400 139.050 351.450 148.800 ;
        RECT 342.000 138.600 346.050 139.050 ;
        RECT 335.400 136.350 336.600 137.100 ;
        RECT 341.400 136.950 346.050 138.600 ;
        RECT 349.950 136.950 352.050 139.050 ;
        RECT 353.400 138.600 354.450 151.800 ;
        RECT 358.950 142.950 361.050 148.050 ;
        RECT 361.950 145.950 364.050 148.050 ;
        RECT 341.400 136.350 342.600 136.950 ;
        RECT 353.400 136.350 354.600 138.600 ;
        RECT 358.950 137.100 361.050 139.200 ;
        RECT 362.400 139.050 363.450 145.950 ;
        RECT 359.400 136.350 360.600 137.100 ;
        RECT 361.950 136.950 364.050 139.050 ;
        RECT 365.400 136.050 366.450 155.400 ;
        RECT 367.800 151.950 369.900 154.050 ;
        RECT 370.950 151.950 373.050 155.400 ;
        RECT 373.950 154.950 376.050 157.050 ;
        RECT 368.400 148.050 369.450 151.950 ;
        RECT 367.950 145.950 370.050 148.050 ;
        RECT 377.400 145.050 378.450 157.950 ;
        RECT 370.950 142.950 376.050 145.050 ;
        RECT 376.950 142.950 379.050 145.050 ;
        RECT 370.950 137.100 373.050 139.200 ;
        RECT 377.400 138.600 378.450 142.950 ;
        RECT 385.950 139.950 388.050 142.050 ;
        RECT 371.400 136.350 372.600 137.100 ;
        RECT 377.400 136.350 378.600 138.600 ;
        RECT 334.950 133.950 337.050 136.050 ;
        RECT 337.950 133.950 340.050 136.050 ;
        RECT 340.950 133.950 343.050 136.050 ;
        RECT 352.950 133.950 355.050 136.050 ;
        RECT 355.950 133.950 358.050 136.050 ;
        RECT 358.950 133.950 361.050 136.050 ;
        RECT 364.950 133.950 367.050 136.050 ;
        RECT 370.950 133.950 373.050 136.050 ;
        RECT 373.950 133.950 376.050 136.050 ;
        RECT 376.950 133.950 379.050 136.050 ;
        RECT 379.950 133.950 382.050 136.050 ;
        RECT 338.400 131.400 339.600 133.650 ;
        RECT 338.400 129.450 339.450 131.400 ;
        RECT 349.950 130.950 352.050 133.050 ;
        RECT 356.400 132.900 357.600 133.650 ;
        RECT 335.400 128.400 339.450 129.450 ;
        RECT 328.950 121.950 331.050 124.050 ;
        RECT 331.950 118.950 334.050 121.050 ;
        RECT 325.950 106.950 328.050 109.050 ;
        RECT 319.950 103.950 322.050 106.050 ;
        RECT 326.400 105.600 327.450 106.950 ;
        RECT 332.400 105.600 333.450 118.950 ;
        RECT 335.400 109.050 336.450 128.400 ;
        RECT 340.950 127.950 343.050 130.050 ;
        RECT 337.950 124.950 340.050 127.050 ;
        RECT 334.950 106.950 337.050 109.050 ;
        RECT 338.400 106.050 339.450 124.950 ;
        RECT 326.400 103.350 327.600 105.600 ;
        RECT 332.400 103.350 333.600 105.600 ;
        RECT 337.950 103.950 340.050 106.050 ;
        RECT 322.950 100.950 325.050 103.050 ;
        RECT 325.950 100.950 328.050 103.050 ;
        RECT 328.950 100.950 331.050 103.050 ;
        RECT 331.950 100.950 334.050 103.050 ;
        RECT 334.950 100.950 337.050 103.050 ;
        RECT 319.950 97.950 322.050 100.050 ;
        RECT 323.400 99.000 324.600 100.650 ;
        RECT 320.400 85.050 321.450 97.950 ;
        RECT 322.950 94.950 325.050 99.000 ;
        RECT 329.400 98.400 330.600 100.650 ;
        RECT 335.400 99.900 336.600 100.650 ;
        RECT 329.400 94.050 330.450 98.400 ;
        RECT 334.950 97.800 337.050 99.900 ;
        RECT 341.400 97.050 342.450 127.950 ;
        RECT 350.400 127.050 351.450 130.950 ;
        RECT 355.950 130.800 358.050 132.900 ;
        RECT 349.950 124.950 352.050 127.050 ;
        RECT 343.950 121.950 346.050 124.050 ;
        RECT 344.400 105.450 345.450 121.950 ;
        RECT 356.400 115.050 357.450 130.800 ;
        RECT 364.950 127.950 367.050 132.900 ;
        RECT 374.400 132.000 375.600 133.650 ;
        RECT 380.400 132.900 381.600 133.650 ;
        RECT 386.400 132.900 387.450 139.950 ;
        RECT 389.400 138.450 390.450 166.950 ;
        RECT 392.400 142.050 393.450 187.950 ;
        RECT 398.400 186.450 399.450 208.800 ;
        RECT 413.400 205.050 414.450 209.400 ;
        RECT 412.950 202.950 415.050 205.050 ;
        RECT 403.950 190.950 406.050 193.050 ;
        RECT 404.400 187.050 405.450 190.950 ;
        RECT 422.400 190.050 423.450 232.950 ;
        RECT 427.950 226.950 430.050 229.050 ;
        RECT 428.400 216.600 429.450 226.950 ;
        RECT 449.400 226.050 450.450 250.950 ;
        RECT 430.950 223.950 433.050 226.050 ;
        RECT 448.950 223.950 451.050 226.050 ;
        RECT 431.400 220.050 432.450 223.950 ;
        RECT 439.950 220.950 442.050 223.050 ;
        RECT 430.950 217.950 433.050 220.050 ;
        RECT 428.400 214.350 429.600 216.600 ;
        RECT 427.950 211.950 430.050 214.050 ;
        RECT 430.950 211.950 433.050 214.050 ;
        RECT 433.950 211.950 436.050 214.050 ;
        RECT 431.400 210.900 432.600 211.650 ;
        RECT 430.950 208.800 433.050 210.900 ;
        RECT 421.950 187.950 424.050 190.050 ;
        RECT 395.400 185.400 399.450 186.450 ;
        RECT 395.400 175.050 396.450 185.400 ;
        RECT 403.950 184.950 406.050 187.050 ;
        RECT 427.950 182.100 430.050 184.200 ;
        RECT 401.400 178.950 403.500 181.050 ;
        RECT 406.800 178.950 408.900 181.050 ;
        RECT 419.400 178.950 421.500 181.050 ;
        RECT 424.800 178.950 426.900 181.050 ;
        RECT 407.400 176.400 408.600 178.650 ;
        RECT 425.400 176.400 426.600 178.650 ;
        RECT 428.400 177.450 429.450 182.100 ;
        RECT 431.400 181.050 432.450 208.800 ;
        RECT 440.400 186.450 441.450 220.950 ;
        RECT 449.400 219.450 450.450 223.950 ;
        RECT 452.400 223.050 453.450 254.400 ;
        RECT 457.950 232.950 460.050 235.050 ;
        RECT 454.950 229.950 457.050 232.050 ;
        RECT 455.400 223.050 456.450 229.950 ;
        RECT 458.400 229.050 459.450 232.950 ;
        RECT 457.950 226.950 460.050 229.050 ;
        RECT 451.800 220.950 453.900 223.050 ;
        RECT 454.950 220.950 457.050 223.050 ;
        RECT 449.400 218.400 453.450 219.450 ;
        RECT 445.950 215.100 448.050 217.200 ;
        RECT 452.400 216.600 453.450 218.400 ;
        RECT 446.400 214.350 447.600 215.100 ;
        RECT 452.400 214.350 453.600 216.600 ;
        RECT 445.950 211.950 448.050 214.050 ;
        RECT 448.950 211.950 451.050 214.050 ;
        RECT 451.950 211.950 454.050 214.050 ;
        RECT 454.950 211.950 457.050 214.050 ;
        RECT 449.400 209.400 450.600 211.650 ;
        RECT 455.400 210.900 456.600 211.650 ;
        RECT 449.400 198.450 450.450 209.400 ;
        RECT 454.950 208.800 457.050 210.900 ;
        RECT 451.950 199.950 454.050 202.050 ;
        RECT 446.400 197.400 450.450 198.450 ;
        RECT 446.400 193.050 447.450 197.400 ;
        RECT 448.950 193.950 451.050 196.050 ;
        RECT 445.950 190.950 448.050 193.050 ;
        RECT 440.400 186.000 447.450 186.450 ;
        RECT 440.400 185.400 448.050 186.000 ;
        RECT 439.950 182.100 442.050 184.200 ;
        RECT 440.400 181.350 441.600 182.100 ;
        RECT 445.950 181.950 448.050 185.400 ;
        RECT 430.950 178.950 433.050 181.050 ;
        RECT 436.950 178.950 439.050 181.050 ;
        RECT 439.950 178.950 442.050 181.050 ;
        RECT 442.950 178.950 445.050 181.050 ;
        RECT 428.400 176.400 432.450 177.450 ;
        RECT 394.950 172.950 397.050 175.050 ;
        RECT 403.950 172.950 406.050 175.050 ;
        RECT 404.400 154.050 405.450 172.950 ;
        RECT 403.950 151.950 406.050 154.050 ;
        RECT 407.400 148.050 408.450 176.400 ;
        RECT 425.400 165.450 426.450 176.400 ;
        RECT 425.400 164.400 429.450 165.450 ;
        RECT 424.950 160.950 427.050 163.050 ;
        RECT 409.950 157.950 412.050 160.050 ;
        RECT 410.400 154.050 411.450 157.950 ;
        RECT 409.950 151.950 412.050 154.050 ;
        RECT 406.950 145.950 409.050 148.050 ;
        RECT 391.950 139.950 394.050 142.050 ;
        RECT 410.400 138.600 411.450 151.950 ;
        RECT 425.400 151.050 426.450 160.950 ;
        RECT 428.400 160.050 429.450 164.400 ;
        RECT 431.400 163.050 432.450 176.400 ;
        RECT 437.400 176.400 438.600 178.650 ;
        RECT 443.400 177.900 444.600 178.650 ;
        RECT 449.400 177.900 450.450 193.950 ;
        RECT 433.950 166.950 436.050 169.050 ;
        RECT 430.950 160.950 433.050 163.050 ;
        RECT 427.950 157.950 430.050 160.050 ;
        RECT 424.950 148.950 427.050 151.050 ;
        RECT 421.950 145.950 424.050 148.050 ;
        RECT 392.400 138.450 393.600 138.600 ;
        RECT 389.400 137.400 393.600 138.450 ;
        RECT 373.950 127.950 376.050 132.000 ;
        RECT 379.950 130.800 382.050 132.900 ;
        RECT 385.950 130.800 388.050 132.900 ;
        RECT 389.400 130.050 390.450 137.400 ;
        RECT 392.400 136.350 393.600 137.400 ;
        RECT 410.400 136.350 411.600 138.600 ;
        RECT 392.100 133.950 394.200 136.050 ;
        RECT 397.500 133.950 399.600 136.050 ;
        RECT 409.950 133.950 412.050 136.050 ;
        RECT 412.950 133.950 415.050 136.050 ;
        RECT 413.400 132.000 414.600 133.650 ;
        RECT 388.950 127.950 391.050 130.050 ;
        RECT 412.950 127.950 415.050 132.000 ;
        RECT 422.400 124.050 423.450 145.950 ;
        RECT 425.400 138.600 426.450 148.950 ;
        RECT 434.400 145.050 435.450 166.950 ;
        RECT 437.400 166.050 438.450 176.400 ;
        RECT 442.950 175.800 445.050 177.900 ;
        RECT 448.950 175.800 451.050 177.900 ;
        RECT 452.400 174.450 453.450 199.950 ;
        RECT 455.400 190.050 456.450 208.800 ;
        RECT 461.400 202.050 462.450 260.100 ;
        RECT 467.400 259.350 468.600 260.100 ;
        RECT 473.400 259.350 474.600 261.600 ;
        RECT 478.950 260.100 481.050 262.200 ;
        RECT 466.950 256.950 469.050 259.050 ;
        RECT 469.950 256.950 472.050 259.050 ;
        RECT 472.950 256.950 475.050 259.050 ;
        RECT 475.950 256.950 478.050 259.050 ;
        RECT 463.950 252.300 466.050 256.050 ;
        RECT 470.400 255.900 471.600 256.650 ;
        RECT 469.950 253.800 472.050 255.900 ;
        RECT 476.400 255.000 477.600 256.650 ;
        RECT 469.950 252.300 472.050 252.750 ;
        RECT 463.950 252.000 472.050 252.300 ;
        RECT 464.400 251.250 472.050 252.000 ;
        RECT 469.950 250.650 472.050 251.250 ;
        RECT 475.950 250.950 478.050 255.000 ;
        RECT 478.950 253.800 481.050 255.900 ;
        RECT 479.400 250.050 480.450 253.800 ;
        RECT 478.950 247.950 481.050 250.050 ;
        RECT 463.950 238.950 466.050 241.050 ;
        RECT 464.400 217.050 465.450 238.950 ;
        RECT 466.950 226.950 469.050 229.050 ;
        RECT 467.400 223.050 468.450 226.950 ;
        RECT 466.950 220.950 469.050 223.050 ;
        RECT 472.950 220.950 475.050 223.050 ;
        RECT 463.800 214.950 465.900 217.050 ;
        RECT 466.950 215.100 469.050 217.200 ;
        RECT 473.400 216.600 474.450 220.950 ;
        RECT 467.400 214.350 468.600 215.100 ;
        RECT 473.400 214.350 474.600 216.600 ;
        RECT 466.950 211.950 469.050 214.050 ;
        RECT 469.950 211.950 472.050 214.050 ;
        RECT 472.950 211.950 475.050 214.050 ;
        RECT 475.950 211.950 478.050 214.050 ;
        RECT 463.950 208.950 466.050 211.050 ;
        RECT 470.400 209.400 471.600 211.650 ;
        RECT 476.400 209.400 477.600 211.650 ;
        RECT 460.950 199.950 463.050 202.050 ;
        RECT 460.950 193.950 463.050 196.050 ;
        RECT 454.950 187.950 457.050 190.050 ;
        RECT 461.400 183.600 462.450 193.950 ;
        RECT 464.400 193.050 465.450 208.950 ;
        RECT 470.400 207.450 471.450 209.400 ;
        RECT 470.400 206.400 474.450 207.450 ;
        RECT 469.950 202.950 472.050 205.050 ;
        RECT 463.950 190.950 466.050 193.050 ;
        RECT 466.950 187.950 469.050 190.050 ;
        RECT 461.400 181.350 462.600 183.600 ;
        RECT 455.100 178.950 457.200 181.050 ;
        RECT 460.500 178.950 462.600 181.050 ;
        RECT 463.800 178.950 465.900 181.050 ;
        RECT 455.400 176.400 456.600 178.650 ;
        RECT 464.400 176.400 465.600 178.650 ;
        RECT 467.400 178.050 468.450 187.950 ;
        RECT 455.400 174.450 456.450 176.400 ;
        RECT 452.400 173.400 456.450 174.450 ;
        RECT 457.800 174.000 459.900 175.050 ;
        RECT 442.950 166.950 445.050 169.050 ;
        RECT 436.950 163.950 439.050 166.050 ;
        RECT 439.950 160.950 442.050 163.050 ;
        RECT 434.400 142.950 439.050 145.050 ;
        RECT 434.400 138.600 435.450 142.950 ;
        RECT 425.400 136.350 426.600 138.600 ;
        RECT 434.400 136.350 435.600 138.600 ;
        RECT 436.950 137.100 439.050 139.200 ;
        RECT 425.100 133.950 427.200 136.050 ;
        RECT 428.400 133.950 430.500 136.050 ;
        RECT 433.800 133.950 435.900 136.050 ;
        RECT 428.400 132.000 429.600 133.650 ;
        RECT 427.950 127.950 430.050 132.000 ;
        RECT 421.800 121.950 423.900 124.050 ;
        RECT 424.950 121.950 427.050 124.050 ;
        RECT 376.950 118.950 379.050 121.050 ;
        RECT 355.950 112.950 358.050 115.050 ;
        RECT 361.950 112.950 364.050 115.050 ;
        RECT 373.950 112.950 376.050 115.050 ;
        RECT 346.950 105.450 349.050 106.050 ;
        RECT 344.400 104.400 349.050 105.450 ;
        RECT 346.950 103.950 349.050 104.400 ;
        RECT 362.400 105.600 363.450 112.950 ;
        RECT 347.400 103.350 348.600 103.950 ;
        RECT 362.400 103.350 363.600 105.600 ;
        RECT 367.950 104.100 370.050 106.200 ;
        RECT 374.400 106.050 375.450 112.950 ;
        RECT 368.400 103.350 369.600 104.100 ;
        RECT 373.950 103.950 376.050 106.050 ;
        RECT 346.950 100.950 349.050 103.050 ;
        RECT 349.950 100.950 352.050 103.050 ;
        RECT 361.950 100.950 364.050 103.050 ;
        RECT 364.950 100.950 367.050 103.050 ;
        RECT 367.950 100.950 370.050 103.050 ;
        RECT 370.950 100.950 373.050 103.050 ;
        RECT 350.400 98.400 351.600 100.650 ;
        RECT 365.400 98.400 366.600 100.650 ;
        RECT 371.400 99.000 372.600 100.650 ;
        RECT 325.950 92.400 330.450 94.050 ;
        RECT 325.950 91.950 330.000 92.400 ;
        RECT 331.950 91.950 334.050 97.050 ;
        RECT 340.950 94.950 343.050 97.050 ;
        RECT 319.950 82.950 322.050 85.050 ;
        RECT 322.950 73.950 325.050 76.050 ;
        RECT 316.950 70.950 319.050 73.050 ;
        RECT 301.950 67.950 304.050 70.050 ;
        RECT 284.400 58.350 285.600 60.600 ;
        RECT 289.950 59.100 292.050 61.200 ;
        RECT 290.400 58.350 291.600 59.100 ;
        RECT 283.950 55.950 286.050 58.050 ;
        RECT 286.950 55.950 289.050 58.050 ;
        RECT 289.950 55.950 292.050 58.050 ;
        RECT 292.950 55.950 295.050 58.050 ;
        RECT 287.400 54.900 288.600 55.650 ;
        RECT 275.400 46.050 276.450 52.950 ;
        RECT 277.950 52.800 280.050 54.900 ;
        RECT 286.950 52.800 289.050 54.900 ;
        RECT 293.400 53.400 294.600 55.650 ;
        RECT 268.950 43.950 271.050 46.050 ;
        RECT 274.950 43.950 277.050 46.050 ;
        RECT 248.400 19.050 249.450 26.100 ;
        RECT 254.400 25.350 255.600 26.100 ;
        RECT 260.400 25.350 261.600 27.600 ;
        RECT 269.400 25.050 270.450 43.950 ;
        RECT 293.400 40.050 294.450 53.400 ;
        RECT 295.950 49.950 298.050 52.050 ;
        RECT 292.950 37.950 295.050 40.050 ;
        RECT 277.950 27.000 280.050 31.050 ;
        RECT 296.400 28.200 297.450 49.950 ;
        RECT 302.400 46.050 303.450 67.950 ;
        RECT 310.950 59.100 313.050 61.200 ;
        RECT 316.950 60.000 319.050 64.050 ;
        RECT 311.400 58.350 312.600 59.100 ;
        RECT 317.400 58.350 318.600 60.000 ;
        RECT 307.950 55.950 310.050 58.050 ;
        RECT 310.950 55.950 313.050 58.050 ;
        RECT 313.950 55.950 316.050 58.050 ;
        RECT 316.950 55.950 319.050 58.050 ;
        RECT 308.400 54.000 309.600 55.650 ;
        RECT 314.400 54.900 315.600 55.650 ;
        RECT 323.400 54.900 324.450 73.950 ;
        RECT 328.950 70.950 331.050 73.050 ;
        RECT 346.950 70.950 349.050 73.050 ;
        RECT 329.400 61.200 330.450 70.950 ;
        RECT 334.950 67.950 337.050 70.050 ;
        RECT 335.400 64.050 336.450 67.950 ;
        RECT 328.950 59.100 331.050 61.200 ;
        RECT 334.950 60.000 337.050 64.050 ;
        RECT 329.400 58.350 330.600 59.100 ;
        RECT 335.400 58.350 336.600 60.000 ;
        RECT 343.950 59.100 346.050 61.200 ;
        RECT 347.400 61.050 348.450 70.950 ;
        RECT 350.400 70.050 351.450 98.400 ;
        RECT 365.400 91.050 366.450 98.400 ;
        RECT 370.950 94.950 373.050 99.000 ;
        RECT 373.950 97.950 376.050 100.050 ;
        RECT 364.950 88.950 367.050 91.050 ;
        RECT 358.950 85.950 361.050 88.050 ;
        RECT 355.950 82.950 358.050 85.050 ;
        RECT 352.950 73.950 355.050 76.050 ;
        RECT 356.400 75.450 357.450 82.950 ;
        RECT 359.400 79.050 360.450 85.950 ;
        RECT 364.950 82.950 367.050 85.050 ;
        RECT 358.950 76.950 361.050 79.050 ;
        RECT 356.400 74.400 360.450 75.450 ;
        RECT 349.950 67.950 352.050 70.050 ;
        RECT 353.400 64.050 354.450 73.950 ;
        RECT 355.950 70.950 358.050 73.050 ;
        RECT 352.950 61.950 355.050 64.050 ;
        RECT 328.950 55.950 331.050 58.050 ;
        RECT 331.950 55.950 334.050 58.050 ;
        RECT 334.950 55.950 337.050 58.050 ;
        RECT 337.950 55.950 340.050 58.050 ;
        RECT 307.950 49.950 310.050 54.000 ;
        RECT 313.950 52.800 316.050 54.900 ;
        RECT 322.800 52.800 324.900 54.900 ;
        RECT 332.400 54.000 333.600 55.650 ;
        RECT 331.950 49.950 334.050 54.000 ;
        RECT 338.400 53.400 339.600 55.650 ;
        RECT 301.950 43.950 304.050 46.050 ;
        RECT 319.950 43.950 322.050 46.050 ;
        RECT 307.950 34.950 310.050 37.050 ;
        RECT 301.950 31.950 304.050 34.050 ;
        RECT 278.400 25.350 279.600 27.000 ;
        RECT 286.950 25.950 289.050 28.050 ;
        RECT 295.950 26.100 298.050 28.200 ;
        RECT 302.400 27.600 303.450 31.950 ;
        RECT 253.950 22.950 256.050 25.050 ;
        RECT 256.950 22.950 259.050 25.050 ;
        RECT 259.950 22.950 262.050 25.050 ;
        RECT 262.950 22.950 265.050 25.050 ;
        RECT 268.950 22.950 271.050 25.050 ;
        RECT 274.950 22.950 277.050 25.050 ;
        RECT 277.950 22.950 280.050 25.050 ;
        RECT 280.950 22.950 283.050 25.050 ;
        RECT 257.400 21.900 258.600 22.650 ;
        RECT 263.400 21.900 264.600 22.650 ;
        RECT 256.950 19.800 259.050 21.900 ;
        RECT 262.950 19.800 265.050 21.900 ;
        RECT 275.400 20.400 276.600 22.650 ;
        RECT 281.400 21.900 282.600 22.650 ;
        RECT 287.400 21.900 288.450 25.950 ;
        RECT 296.400 25.350 297.600 26.100 ;
        RECT 302.400 25.350 303.600 27.600 ;
        RECT 292.950 22.950 295.050 25.050 ;
        RECT 295.950 22.950 298.050 25.050 ;
        RECT 298.950 22.950 301.050 25.050 ;
        RECT 301.950 22.950 304.050 25.050 ;
        RECT 293.400 21.900 294.600 22.650 ;
        RECT 247.950 16.950 250.050 19.050 ;
        RECT 244.950 10.950 247.050 13.050 ;
        RECT 248.400 10.050 249.450 16.950 ;
        RECT 275.400 16.050 276.450 20.400 ;
        RECT 280.950 19.800 283.050 21.900 ;
        RECT 286.950 19.800 289.050 21.900 ;
        RECT 292.950 19.800 295.050 21.900 ;
        RECT 299.400 20.400 300.600 22.650 ;
        RECT 308.400 21.900 309.450 34.950 ;
        RECT 313.950 26.100 316.050 28.200 ;
        RECT 320.400 27.600 321.450 43.950 ;
        RECT 328.950 31.950 331.050 34.050 ;
        RECT 338.400 33.450 339.450 53.400 ;
        RECT 344.400 49.050 345.450 59.100 ;
        RECT 346.950 58.950 349.050 61.050 ;
        RECT 349.950 59.100 352.050 61.200 ;
        RECT 356.400 60.600 357.450 70.950 ;
        RECT 359.400 67.050 360.450 74.400 ;
        RECT 358.950 64.950 361.050 67.050 ;
        RECT 350.400 58.350 351.600 59.100 ;
        RECT 356.400 58.350 357.600 60.600 ;
        RECT 349.950 55.950 352.050 58.050 ;
        RECT 352.950 55.950 355.050 58.050 ;
        RECT 355.950 55.950 358.050 58.050 ;
        RECT 358.950 55.950 361.050 58.050 ;
        RECT 346.950 52.950 349.050 55.050 ;
        RECT 353.400 54.900 354.600 55.650 ;
        RECT 343.950 46.950 346.050 49.050 ;
        RECT 347.400 46.050 348.450 52.950 ;
        RECT 352.950 52.800 355.050 54.900 ;
        RECT 359.400 53.400 360.600 55.650 ;
        RECT 365.400 54.450 366.450 82.950 ;
        RECT 374.400 82.050 375.450 97.950 ;
        RECT 377.400 91.050 378.450 118.950 ;
        RECT 385.950 112.950 388.050 115.050 ;
        RECT 403.950 112.950 406.050 115.050 ;
        RECT 409.950 112.950 412.050 115.050 ;
        RECT 418.950 112.950 421.050 115.050 ;
        RECT 386.400 106.200 387.450 112.950 ;
        RECT 385.950 104.100 388.050 106.200 ;
        RECT 404.400 105.600 405.450 112.950 ;
        RECT 410.400 105.600 411.450 112.950 ;
        RECT 392.400 105.450 393.600 105.600 ;
        RECT 392.400 104.400 399.450 105.450 ;
        RECT 386.400 103.350 387.600 104.100 ;
        RECT 392.400 103.350 393.600 104.400 ;
        RECT 382.950 100.950 385.050 103.050 ;
        RECT 385.950 100.950 388.050 103.050 ;
        RECT 388.950 100.950 391.050 103.050 ;
        RECT 391.950 100.950 394.050 103.050 ;
        RECT 379.950 97.950 382.050 100.050 ;
        RECT 383.400 98.400 384.600 100.650 ;
        RECT 389.400 99.900 390.600 100.650 ;
        RECT 376.950 88.950 379.050 91.050 ;
        RECT 373.950 79.950 376.050 82.050 ;
        RECT 367.950 73.950 370.050 76.050 ;
        RECT 368.400 67.050 369.450 73.950 ;
        RECT 380.400 73.050 381.450 97.950 ;
        RECT 383.400 91.050 384.450 98.400 ;
        RECT 388.950 94.950 391.050 99.900 ;
        RECT 382.950 88.950 385.050 91.050 ;
        RECT 382.950 79.950 385.050 82.050 ;
        RECT 373.950 70.950 376.050 73.050 ;
        RECT 379.950 70.950 382.050 73.050 ;
        RECT 367.950 64.950 370.050 67.050 ;
        RECT 374.400 60.600 375.450 70.950 ;
        RECT 379.950 64.950 382.050 67.050 ;
        RECT 380.400 60.600 381.450 64.950 ;
        RECT 383.400 61.050 384.450 79.950 ;
        RECT 385.950 64.950 388.050 67.050 ;
        RECT 394.950 64.950 397.050 67.050 ;
        RECT 374.400 58.350 375.600 60.600 ;
        RECT 380.400 58.350 381.600 60.600 ;
        RECT 382.950 58.950 385.050 61.050 ;
        RECT 370.950 55.950 373.050 58.050 ;
        RECT 373.950 55.950 376.050 58.050 ;
        RECT 376.950 55.950 379.050 58.050 ;
        RECT 379.950 55.950 382.050 58.050 ;
        RECT 371.400 54.450 372.600 55.650 ;
        RECT 365.400 53.400 372.600 54.450 ;
        RECT 377.400 53.400 378.600 55.650 ;
        RECT 359.400 49.050 360.450 53.400 ;
        RECT 365.400 49.050 366.450 53.400 ;
        RECT 370.950 49.950 373.050 52.050 ;
        RECT 358.950 46.950 361.050 49.050 ;
        RECT 364.950 46.950 367.050 49.050 ;
        RECT 371.400 46.050 372.450 49.950 ;
        RECT 346.950 43.950 349.050 46.050 ;
        RECT 370.950 43.950 373.050 46.050 ;
        RECT 377.400 43.050 378.450 53.400 ;
        RECT 386.400 46.050 387.450 64.950 ;
        RECT 395.400 60.600 396.450 64.950 ;
        RECT 398.400 63.450 399.450 104.400 ;
        RECT 404.400 103.350 405.600 105.600 ;
        RECT 410.400 103.350 411.600 105.600 ;
        RECT 419.400 103.050 420.450 112.950 ;
        RECT 425.400 112.050 426.450 121.950 ;
        RECT 437.400 115.050 438.450 137.100 ;
        RECT 440.400 121.050 441.450 160.950 ;
        RECT 443.400 154.050 444.450 166.950 ;
        RECT 452.400 166.050 453.450 173.400 ;
        RECT 457.800 172.950 460.050 174.000 ;
        RECT 460.950 172.950 463.050 175.050 ;
        RECT 457.950 171.450 460.050 172.950 ;
        RECT 455.400 171.000 460.050 171.450 ;
        RECT 455.400 170.400 459.450 171.000 ;
        RECT 451.950 163.950 454.050 166.050 ;
        RECT 455.400 160.050 456.450 170.400 ;
        RECT 457.950 160.950 460.050 163.050 ;
        RECT 454.950 157.950 457.050 160.050 ;
        RECT 454.950 154.800 457.050 156.900 ;
        RECT 442.950 151.950 445.050 154.050 ;
        RECT 451.950 151.950 454.050 154.050 ;
        RECT 448.950 148.950 451.050 151.050 ;
        RECT 449.400 142.050 450.450 148.950 ;
        RECT 448.950 139.950 451.050 142.050 ;
        RECT 445.950 137.100 448.050 139.200 ;
        RECT 452.400 138.600 453.450 151.950 ;
        RECT 455.400 151.050 456.450 154.800 ;
        RECT 454.950 148.950 457.050 151.050 ;
        RECT 458.400 148.050 459.450 160.950 ;
        RECT 457.950 145.950 460.050 148.050 ;
        RECT 446.400 136.350 447.600 137.100 ;
        RECT 452.400 136.350 453.600 138.600 ;
        RECT 445.950 133.950 448.050 136.050 ;
        RECT 448.950 133.950 451.050 136.050 ;
        RECT 451.950 133.950 454.050 136.050 ;
        RECT 454.950 133.950 457.050 136.050 ;
        RECT 449.400 131.400 450.600 133.650 ;
        RECT 455.400 132.900 456.600 133.650 ;
        RECT 449.400 124.050 450.450 131.400 ;
        RECT 454.950 130.800 457.050 132.900 ;
        RECT 457.950 130.950 460.050 133.050 ;
        RECT 448.950 121.950 451.050 124.050 ;
        RECT 439.950 118.950 442.050 121.050 ;
        RECT 446.400 116.400 453.450 117.450 ;
        RECT 436.950 112.950 439.050 115.050 ;
        RECT 446.400 112.050 447.450 116.400 ;
        RECT 448.950 112.950 451.050 115.050 ;
        RECT 424.950 109.950 427.050 112.050 ;
        RECT 445.950 109.950 448.050 112.050 ;
        RECT 449.400 106.200 450.450 112.950 ;
        RECT 452.400 112.050 453.450 116.400 ;
        RECT 451.950 109.950 454.050 112.050 ;
        RECT 427.950 104.100 430.050 106.200 ;
        RECT 435.000 105.600 439.050 106.050 ;
        RECT 428.400 103.350 429.600 104.100 ;
        RECT 434.400 103.950 439.050 105.600 ;
        RECT 439.950 104.100 442.050 106.200 ;
        RECT 448.950 104.100 451.050 106.200 ;
        RECT 454.950 104.100 457.050 106.200 ;
        RECT 458.400 106.050 459.450 130.950 ;
        RECT 434.400 103.350 435.600 103.950 ;
        RECT 403.950 100.950 406.050 103.050 ;
        RECT 406.950 100.950 409.050 103.050 ;
        RECT 409.950 100.950 412.050 103.050 ;
        RECT 412.950 100.950 415.050 103.050 ;
        RECT 418.950 100.950 421.050 103.050 ;
        RECT 424.950 100.950 427.050 103.050 ;
        RECT 427.950 100.950 430.050 103.050 ;
        RECT 430.950 100.950 433.050 103.050 ;
        RECT 433.950 100.950 436.050 103.050 ;
        RECT 407.400 98.400 408.600 100.650 ;
        RECT 413.400 98.400 414.600 100.650 ;
        RECT 425.400 99.900 426.600 100.650 ;
        RECT 431.400 99.900 432.600 100.650 ;
        RECT 407.400 76.050 408.450 98.400 ;
        RECT 413.400 94.050 414.450 98.400 ;
        RECT 424.950 97.800 427.050 99.900 ;
        RECT 430.950 97.800 433.050 99.900 ;
        RECT 436.950 97.800 439.050 99.900 ;
        RECT 412.950 91.950 415.050 94.050 ;
        RECT 437.400 79.050 438.450 97.800 ;
        RECT 440.400 94.050 441.450 104.100 ;
        RECT 449.400 103.350 450.600 104.100 ;
        RECT 455.400 103.350 456.600 104.100 ;
        RECT 457.950 103.950 460.050 106.050 ;
        RECT 445.950 100.950 448.050 103.050 ;
        RECT 448.950 100.950 451.050 103.050 ;
        RECT 451.950 100.950 454.050 103.050 ;
        RECT 454.950 100.950 457.050 103.050 ;
        RECT 446.400 98.400 447.600 100.650 ;
        RECT 452.400 99.900 453.600 100.650 ;
        RECT 442.950 94.950 445.050 97.050 ;
        RECT 439.950 91.950 442.050 94.050 ;
        RECT 436.950 76.950 439.050 79.050 ;
        RECT 443.400 76.050 444.450 94.950 ;
        RECT 446.400 94.050 447.450 98.400 ;
        RECT 451.950 97.800 454.050 99.900 ;
        RECT 451.950 94.650 454.050 96.750 ;
        RECT 457.950 94.950 460.050 100.050 ;
        RECT 445.950 91.950 448.050 94.050 ;
        RECT 452.400 91.050 453.450 94.650 ;
        RECT 451.950 88.950 454.050 91.050 ;
        RECT 454.950 82.950 457.050 85.050 ;
        RECT 406.950 73.950 409.050 76.050 ;
        RECT 442.950 73.950 445.050 76.050 ;
        RECT 445.950 67.950 448.050 70.050 ;
        RECT 398.400 62.400 402.450 63.450 ;
        RECT 401.400 61.200 402.450 62.400 ;
        RECT 395.400 58.350 396.600 60.600 ;
        RECT 400.950 59.100 403.050 61.200 ;
        RECT 415.950 60.000 418.050 64.050 ;
        RECT 401.400 58.350 402.600 59.100 ;
        RECT 416.400 58.350 417.600 60.000 ;
        RECT 421.950 59.100 424.050 61.200 ;
        RECT 427.950 59.100 430.050 61.200 ;
        RECT 436.950 59.100 439.050 61.200 ;
        RECT 442.950 59.100 445.050 64.050 ;
        RECT 446.400 61.050 447.450 67.950 ;
        RECT 455.400 64.050 456.450 82.950 ;
        RECT 457.950 64.950 460.050 67.050 ;
        RECT 454.950 61.950 457.050 64.050 ;
        RECT 422.400 58.350 423.600 59.100 ;
        RECT 391.950 55.950 394.050 58.050 ;
        RECT 394.950 55.950 397.050 58.050 ;
        RECT 397.950 55.950 400.050 58.050 ;
        RECT 400.950 55.950 403.050 58.050 ;
        RECT 412.950 55.950 415.050 58.050 ;
        RECT 415.950 55.950 418.050 58.050 ;
        RECT 418.950 55.950 421.050 58.050 ;
        RECT 421.950 55.950 424.050 58.050 ;
        RECT 388.950 52.950 391.050 55.050 ;
        RECT 392.400 54.000 393.600 55.650 ;
        RECT 379.950 43.950 382.050 46.050 ;
        RECT 385.950 43.950 388.050 46.050 ;
        RECT 343.950 40.950 346.050 43.050 ;
        RECT 376.950 40.950 379.050 43.050 ;
        RECT 344.400 37.050 345.450 40.950 ;
        RECT 373.950 39.450 376.050 40.050 ;
        RECT 380.400 39.450 381.450 43.950 ;
        RECT 373.950 38.400 381.450 39.450 ;
        RECT 373.950 37.950 376.050 38.400 ;
        RECT 344.400 35.400 349.050 37.050 ;
        RECT 345.000 34.950 349.050 35.400 ;
        RECT 352.950 34.950 358.050 37.050 ;
        RECT 370.950 34.950 373.050 37.050 ;
        RECT 382.950 34.950 385.050 37.050 ;
        RECT 338.400 33.000 342.450 33.450 ;
        RECT 338.400 32.400 343.050 33.000 ;
        RECT 314.400 25.350 315.600 26.100 ;
        RECT 320.400 25.350 321.600 27.600 ;
        RECT 313.950 22.950 316.050 25.050 ;
        RECT 316.950 22.950 319.050 25.050 ;
        RECT 319.950 22.950 322.050 25.050 ;
        RECT 322.950 22.950 325.050 25.050 ;
        RECT 293.400 16.050 294.450 19.800 ;
        RECT 274.950 13.950 277.050 16.050 ;
        RECT 292.950 13.950 295.050 16.050 ;
        RECT 247.950 7.950 250.050 10.050 ;
        RECT 299.400 7.050 300.450 20.400 ;
        RECT 307.950 19.800 310.050 21.900 ;
        RECT 317.400 21.000 318.600 22.650 ;
        RECT 323.400 21.900 324.600 22.650 ;
        RECT 329.400 21.900 330.450 31.950 ;
        RECT 331.950 25.950 334.050 31.050 ;
        RECT 337.800 30.000 339.900 31.050 ;
        RECT 337.800 28.950 340.050 30.000 ;
        RECT 340.950 28.950 343.050 32.400 ;
        RECT 337.950 27.000 340.050 28.950 ;
        RECT 338.400 25.350 339.600 27.000 ;
        RECT 343.950 26.100 346.050 28.200 ;
        RECT 355.950 26.100 358.050 28.200 ;
        RECT 361.950 26.100 364.050 28.200 ;
        RECT 344.400 25.350 345.600 26.100 ;
        RECT 356.400 25.350 357.600 26.100 ;
        RECT 362.400 25.350 363.600 26.100 ;
        RECT 334.950 22.950 337.050 25.050 ;
        RECT 337.950 22.950 340.050 25.050 ;
        RECT 340.950 22.950 343.050 25.050 ;
        RECT 343.950 22.950 346.050 25.050 ;
        RECT 355.950 22.950 358.050 25.050 ;
        RECT 358.950 22.950 361.050 25.050 ;
        RECT 361.950 22.950 364.050 25.050 ;
        RECT 364.950 22.950 367.050 25.050 ;
        RECT 316.950 16.950 319.050 21.000 ;
        RECT 322.950 19.800 325.050 21.900 ;
        RECT 328.950 19.800 331.050 21.900 ;
        RECT 335.400 20.400 336.600 22.650 ;
        RECT 341.400 21.900 342.600 22.650 ;
        RECT 319.950 13.950 322.050 16.050 ;
        RECT 320.400 10.050 321.450 13.950 ;
        RECT 329.400 10.050 330.450 19.800 ;
        RECT 335.400 16.050 336.450 20.400 ;
        RECT 340.950 19.800 343.050 21.900 ;
        RECT 359.400 20.400 360.600 22.650 ;
        RECT 365.400 21.900 366.600 22.650 ;
        RECT 359.400 16.050 360.450 20.400 ;
        RECT 364.950 19.800 367.050 21.900 ;
        RECT 371.400 19.050 372.450 34.950 ;
        RECT 376.950 31.950 379.050 34.050 ;
        RECT 377.400 27.600 378.450 31.950 ;
        RECT 383.400 28.200 384.450 34.950 ;
        RECT 377.400 25.350 378.600 27.600 ;
        RECT 382.950 26.100 385.050 28.200 ;
        RECT 389.400 28.050 390.450 52.950 ;
        RECT 391.950 49.950 394.050 54.000 ;
        RECT 398.400 53.400 399.600 55.650 ;
        RECT 398.400 51.450 399.450 53.400 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 413.400 53.400 414.600 55.650 ;
        RECT 419.400 53.400 420.600 55.650 ;
        RECT 395.400 50.400 399.450 51.450 ;
        RECT 391.950 40.950 394.050 43.050 ;
        RECT 383.400 25.350 384.600 26.100 ;
        RECT 388.950 25.950 391.050 28.050 ;
        RECT 376.950 22.950 379.050 25.050 ;
        RECT 379.950 22.950 382.050 25.050 ;
        RECT 382.950 22.950 385.050 25.050 ;
        RECT 385.950 22.950 388.050 25.050 ;
        RECT 380.400 21.900 381.600 22.650 ;
        RECT 386.400 21.900 387.600 22.650 ;
        RECT 370.950 16.950 373.050 19.050 ;
        RECT 376.950 16.050 379.050 19.050 ;
        RECT 379.950 16.950 382.050 21.900 ;
        RECT 385.950 19.800 388.050 21.900 ;
        RECT 386.400 16.050 387.450 19.800 ;
        RECT 392.400 19.050 393.450 40.950 ;
        RECT 395.400 40.050 396.450 50.400 ;
        RECT 410.400 46.050 411.450 52.950 ;
        RECT 409.950 43.950 412.050 46.050 ;
        RECT 400.950 40.950 403.050 43.050 ;
        RECT 394.950 37.950 397.050 40.050 ;
        RECT 401.400 27.600 402.450 40.950 ;
        RECT 413.400 37.050 414.450 53.400 ;
        RECT 419.400 49.050 420.450 53.400 ;
        RECT 428.400 49.050 429.450 59.100 ;
        RECT 437.400 58.350 438.600 59.100 ;
        RECT 443.400 58.350 444.600 59.100 ;
        RECT 445.950 58.950 448.050 61.050 ;
        RECT 458.400 60.600 459.450 64.950 ;
        RECT 461.400 64.050 462.450 172.950 ;
        RECT 464.400 148.050 465.450 176.400 ;
        RECT 466.950 175.950 469.050 178.050 ;
        RECT 470.400 175.050 471.450 202.950 ;
        RECT 473.400 184.050 474.450 206.400 ;
        RECT 476.400 196.050 477.450 209.400 ;
        RECT 482.400 205.050 483.450 274.950 ;
        RECT 484.950 271.950 487.050 274.050 ;
        RECT 485.400 262.050 486.450 271.950 ;
        RECT 491.400 264.450 492.450 280.950 ;
        RECT 494.400 268.050 495.450 286.950 ;
        RECT 493.950 265.950 496.050 268.050 ;
        RECT 497.400 264.450 498.450 313.950 ;
        RECT 500.400 274.050 501.450 316.950 ;
        RECT 503.550 303.300 505.650 305.400 ;
        RECT 503.550 296.700 504.750 303.300 ;
        RECT 503.550 294.600 505.650 296.700 ;
        RECT 503.550 281.700 504.750 294.600 ;
        RECT 508.950 289.950 511.050 292.050 ;
        RECT 509.400 287.400 510.600 289.650 ;
        RECT 509.400 283.050 510.450 287.400 ;
        RECT 503.550 279.600 505.650 281.700 ;
        RECT 508.950 280.950 511.050 283.050 ;
        RECT 515.400 277.050 516.450 332.400 ;
        RECT 520.950 328.950 523.050 333.000 ;
        RECT 526.950 331.800 529.050 333.900 ;
        RECT 527.400 328.050 528.450 331.800 ;
        RECT 526.950 325.950 529.050 328.050 ;
        RECT 533.400 325.050 534.450 340.950 ;
        RECT 542.400 339.600 543.450 340.950 ;
        RECT 542.400 337.350 543.600 339.600 ;
        RECT 548.400 339.450 549.600 339.600 ;
        RECT 551.400 339.450 552.450 343.950 ;
        RECT 563.400 339.600 564.450 349.950 ;
        RECT 548.400 338.400 555.450 339.450 ;
        RECT 548.400 337.350 549.600 338.400 ;
        RECT 538.950 334.950 541.050 337.050 ;
        RECT 541.950 334.950 544.050 337.050 ;
        RECT 544.950 334.950 547.050 337.050 ;
        RECT 547.950 334.950 550.050 337.050 ;
        RECT 539.400 333.900 540.600 334.650 ;
        RECT 538.950 331.800 541.050 333.900 ;
        RECT 545.400 333.000 546.600 334.650 ;
        RECT 554.400 333.900 555.450 338.400 ;
        RECT 563.400 337.350 564.600 339.600 ;
        RECT 559.950 334.950 562.050 337.050 ;
        RECT 562.950 334.950 565.050 337.050 ;
        RECT 565.950 334.950 568.050 337.050 ;
        RECT 560.400 333.900 561.600 334.650 ;
        RECT 544.950 328.950 547.050 333.000 ;
        RECT 553.950 331.800 556.050 333.900 ;
        RECT 559.950 331.800 562.050 333.900 ;
        RECT 568.950 331.950 571.050 334.050 ;
        RECT 565.950 328.650 568.050 330.750 ;
        RECT 559.950 325.950 562.050 328.050 ;
        RECT 562.950 325.950 565.050 328.050 ;
        RECT 532.950 322.950 535.050 325.050 ;
        RECT 553.950 319.950 556.050 322.050 ;
        RECT 523.950 313.950 526.050 316.050 ;
        RECT 517.950 310.950 520.050 313.050 ;
        RECT 518.400 289.050 519.450 310.950 ;
        RECT 520.950 295.950 523.050 298.050 ;
        RECT 517.950 286.950 520.050 289.050 ;
        RECT 514.950 274.950 517.050 277.050 ;
        RECT 499.950 271.950 502.050 274.050 ;
        RECT 502.950 268.950 505.050 271.050 ;
        RECT 491.400 263.400 495.450 264.450 ;
        RECT 497.400 264.000 501.450 264.450 ;
        RECT 497.400 263.400 502.050 264.000 ;
        RECT 484.950 259.950 487.050 262.050 ;
        RECT 487.950 260.100 490.050 262.200 ;
        RECT 494.400 261.600 495.450 263.400 ;
        RECT 488.400 259.350 489.600 260.100 ;
        RECT 494.400 259.350 495.600 261.600 ;
        RECT 499.950 259.950 502.050 263.400 ;
        RECT 487.950 256.950 490.050 259.050 ;
        RECT 490.950 256.950 493.050 259.050 ;
        RECT 493.950 256.950 496.050 259.050 ;
        RECT 496.950 256.950 499.050 259.050 ;
        RECT 484.950 253.950 487.050 256.050 ;
        RECT 491.400 254.400 492.600 256.650 ;
        RECT 497.400 255.900 498.600 256.650 ;
        RECT 485.400 217.050 486.450 253.950 ;
        RECT 491.400 241.050 492.450 254.400 ;
        RECT 496.950 253.800 499.050 255.900 ;
        RECT 499.950 253.950 502.050 256.050 ;
        RECT 500.400 247.050 501.450 253.950 ;
        RECT 503.400 250.050 504.450 268.950 ;
        RECT 505.950 265.950 508.050 268.050 ;
        RECT 502.950 247.950 505.050 250.050 ;
        RECT 499.950 244.950 502.050 247.050 ;
        RECT 490.950 238.950 493.050 241.050 ;
        RECT 506.400 226.050 507.450 265.950 ;
        RECT 509.100 256.950 511.200 259.050 ;
        RECT 512.400 256.950 514.500 259.050 ;
        RECT 517.800 256.950 519.900 259.050 ;
        RECT 521.400 258.450 522.450 295.950 ;
        RECT 524.400 294.600 525.450 313.950 ;
        RECT 541.950 307.950 544.050 310.050 ;
        RECT 524.400 292.350 525.600 294.600 ;
        RECT 532.950 293.100 535.050 295.200 ;
        RECT 542.400 295.050 543.450 307.950 ;
        RECT 554.400 300.450 555.450 319.950 ;
        RECT 560.400 310.050 561.450 325.950 ;
        RECT 556.950 307.950 561.450 310.050 ;
        RECT 560.400 307.050 561.450 307.950 ;
        RECT 559.950 304.950 562.050 307.050 ;
        RECT 545.400 300.000 555.450 300.450 ;
        RECT 544.950 299.400 555.450 300.000 ;
        RECT 544.950 295.950 547.050 299.400 ;
        RECT 533.400 292.350 534.600 293.100 ;
        RECT 538.950 292.950 541.050 295.050 ;
        RECT 541.950 292.950 544.050 295.050 ;
        RECT 547.950 294.000 550.050 298.050 ;
        RECT 555.000 294.600 559.050 295.050 ;
        RECT 524.100 289.950 526.200 292.050 ;
        RECT 529.500 289.950 531.600 292.050 ;
        RECT 532.800 289.950 534.900 292.050 ;
        RECT 539.400 285.450 540.450 292.950 ;
        RECT 548.400 292.350 549.600 294.000 ;
        RECT 554.400 292.950 559.050 294.600 ;
        RECT 559.950 293.100 562.050 295.200 ;
        RECT 554.400 292.350 555.600 292.950 ;
        RECT 544.950 289.950 547.050 292.050 ;
        RECT 547.950 289.950 550.050 292.050 ;
        RECT 550.950 289.950 553.050 292.050 ;
        RECT 553.950 289.950 556.050 292.050 ;
        RECT 545.400 288.900 546.600 289.650 ;
        RECT 551.400 288.900 552.600 289.650 ;
        RECT 544.950 286.800 547.050 288.900 ;
        RECT 550.950 286.800 553.050 288.900 ;
        RECT 556.950 286.950 559.050 289.050 ;
        RECT 539.400 284.400 543.450 285.450 ;
        RECT 535.950 277.950 538.050 282.900 ;
        RECT 538.950 280.950 541.050 283.050 ;
        RECT 536.400 271.050 537.450 277.950 ;
        RECT 532.800 268.950 534.900 271.050 ;
        RECT 535.950 268.950 538.050 271.050 ;
        RECT 533.400 261.600 534.450 268.950 ;
        RECT 539.400 261.600 540.450 280.950 ;
        RECT 542.400 280.050 543.450 284.400 ;
        RECT 544.950 280.950 547.050 283.050 ;
        RECT 541.950 277.950 544.050 280.050 ;
        RECT 533.400 259.350 534.600 261.600 ;
        RECT 539.400 259.350 540.600 261.600 ;
        RECT 521.400 257.400 525.450 258.450 ;
        RECT 509.400 255.900 510.600 256.650 ;
        RECT 508.950 253.800 511.050 255.900 ;
        RECT 518.400 254.400 519.600 256.650 ;
        RECT 505.950 223.950 508.050 226.050 ;
        RECT 493.950 220.950 496.050 223.050 ;
        RECT 502.950 220.950 505.050 223.050 ;
        RECT 484.800 214.950 486.900 217.050 ;
        RECT 487.950 215.100 490.050 217.200 ;
        RECT 494.400 216.600 495.450 220.950 ;
        RECT 488.400 214.350 489.600 215.100 ;
        RECT 494.400 214.350 495.600 216.600 ;
        RECT 487.950 211.950 490.050 214.050 ;
        RECT 490.950 211.950 493.050 214.050 ;
        RECT 493.950 211.950 496.050 214.050 ;
        RECT 491.400 209.400 492.600 211.650 ;
        RECT 487.950 205.950 490.050 208.050 ;
        RECT 481.950 202.950 484.050 205.050 ;
        RECT 475.950 193.950 478.050 196.050 ;
        RECT 472.950 181.950 475.050 184.050 ;
        RECT 478.950 182.100 481.050 184.200 ;
        RECT 479.400 181.350 480.600 182.100 ;
        RECT 475.950 178.950 478.050 181.050 ;
        RECT 478.950 178.950 481.050 181.050 ;
        RECT 481.950 178.950 484.050 181.050 ;
        RECT 476.400 176.400 477.600 178.650 ;
        RECT 482.400 176.400 483.600 178.650 ;
        RECT 469.950 172.950 472.050 175.050 ;
        RECT 466.950 169.950 469.050 172.050 ;
        RECT 467.400 157.050 468.450 169.950 ;
        RECT 476.400 163.050 477.450 176.400 ;
        RECT 482.400 174.450 483.450 176.400 ;
        RECT 479.400 173.400 483.450 174.450 ;
        RECT 475.950 160.950 478.050 163.050 ;
        RECT 466.950 154.950 469.050 157.050 ;
        RECT 472.950 151.950 475.050 154.050 ;
        RECT 463.950 145.950 466.050 148.050 ;
        RECT 463.950 138.600 468.000 139.050 ;
        RECT 473.400 138.600 474.450 151.950 ;
        RECT 479.400 145.050 480.450 173.400 ;
        RECT 484.950 169.950 487.050 172.050 ;
        RECT 485.400 157.050 486.450 169.950 ;
        RECT 488.400 157.050 489.450 205.950 ;
        RECT 491.400 199.050 492.450 209.400 ;
        RECT 496.950 208.950 499.050 211.050 ;
        RECT 503.400 210.900 504.450 220.950 ;
        RECT 509.400 216.600 510.450 253.800 ;
        RECT 518.400 247.050 519.450 254.400 ;
        RECT 524.400 253.050 525.450 257.400 ;
        RECT 529.950 256.950 532.050 259.050 ;
        RECT 532.950 256.950 535.050 259.050 ;
        RECT 535.950 256.950 538.050 259.050 ;
        RECT 538.950 256.950 541.050 259.050 ;
        RECT 530.400 255.450 531.600 256.650 ;
        RECT 527.400 254.400 531.600 255.450 ;
        RECT 536.400 255.000 537.600 256.650 ;
        RECT 523.950 250.950 526.050 253.050 ;
        RECT 517.950 244.950 520.050 247.050 ;
        RECT 527.400 217.200 528.450 254.400 ;
        RECT 535.950 250.950 538.050 255.000 ;
        RECT 532.950 232.950 535.050 235.050 ;
        RECT 533.400 226.050 534.450 232.950 ;
        RECT 535.950 229.950 538.050 232.050 ;
        RECT 541.950 229.950 544.050 232.050 ;
        RECT 532.950 223.950 535.050 226.050 ;
        RECT 536.400 220.050 537.450 229.950 ;
        RECT 509.400 214.350 510.600 216.600 ;
        RECT 514.950 215.100 517.050 217.200 ;
        RECT 526.950 215.100 529.050 217.200 ;
        RECT 535.950 216.000 538.050 220.050 ;
        RECT 515.400 214.350 516.600 215.100 ;
        RECT 527.400 214.350 528.600 215.100 ;
        RECT 536.400 214.350 537.600 216.000 ;
        RECT 508.950 211.950 511.050 214.050 ;
        RECT 511.950 211.950 514.050 214.050 ;
        RECT 514.950 211.950 517.050 214.050 ;
        RECT 527.100 211.950 529.200 214.050 ;
        RECT 530.400 211.950 532.500 214.050 ;
        RECT 535.800 211.950 537.900 214.050 ;
        RECT 512.400 210.900 513.600 211.650 ;
        RECT 490.950 196.950 493.050 199.050 ;
        RECT 497.400 196.050 498.450 208.950 ;
        RECT 502.950 208.800 505.050 210.900 ;
        RECT 511.950 208.800 514.050 210.900 ;
        RECT 542.400 205.050 543.450 229.950 ;
        RECT 511.950 202.950 514.050 205.050 ;
        RECT 541.950 202.950 544.050 205.050 ;
        RECT 499.950 199.950 502.050 202.050 ;
        RECT 496.950 193.950 499.050 196.050 ;
        RECT 500.400 190.050 501.450 199.950 ;
        RECT 499.950 187.950 502.050 190.050 ;
        RECT 505.950 187.950 508.050 190.050 ;
        RECT 490.950 181.950 493.050 184.050 ;
        RECT 499.950 182.100 502.050 184.200 ;
        RECT 506.400 183.600 507.450 187.950 ;
        RECT 491.400 177.900 492.450 181.950 ;
        RECT 500.400 181.350 501.600 182.100 ;
        RECT 506.400 181.350 507.600 183.600 ;
        RECT 496.950 178.950 499.050 181.050 ;
        RECT 499.950 178.950 502.050 181.050 ;
        RECT 502.950 178.950 505.050 181.050 ;
        RECT 505.950 178.950 508.050 181.050 ;
        RECT 497.400 177.900 498.600 178.650 ;
        RECT 490.950 175.800 493.050 177.900 ;
        RECT 496.950 175.800 499.050 177.900 ;
        RECT 503.400 176.400 504.600 178.650 ;
        RECT 491.400 172.050 492.450 175.800 ;
        RECT 499.950 172.050 502.050 175.050 ;
        RECT 490.950 169.950 493.050 172.050 ;
        RECT 496.950 171.000 502.050 172.050 ;
        RECT 496.950 170.400 501.450 171.000 ;
        RECT 496.950 169.950 501.000 170.400 ;
        RECT 503.400 163.050 504.450 176.400 ;
        RECT 508.950 175.950 511.050 178.050 ;
        RECT 499.800 160.950 501.900 163.050 ;
        RECT 502.950 160.950 505.050 163.050 ;
        RECT 509.400 162.450 510.450 175.950 ;
        RECT 506.400 161.400 510.450 162.450 ;
        RECT 484.800 154.950 486.900 157.050 ;
        RECT 487.950 154.950 490.050 157.050 ;
        RECT 481.950 145.950 484.050 148.050 ;
        RECT 478.950 142.950 481.050 145.050 ;
        RECT 482.400 142.050 483.450 145.950 ;
        RECT 481.950 139.950 484.050 142.050 ;
        RECT 463.950 136.950 468.600 138.600 ;
        RECT 467.400 136.350 468.600 136.950 ;
        RECT 473.400 136.350 474.600 138.600 ;
        RECT 485.400 138.450 486.450 154.950 ;
        RECT 488.400 151.050 489.450 154.950 ;
        RECT 493.950 151.950 496.050 154.050 ;
        RECT 487.950 148.950 490.050 151.050 ;
        RECT 494.400 138.600 495.450 151.950 ;
        RECT 500.400 148.050 501.450 160.950 ;
        RECT 502.950 154.950 505.050 157.050 ;
        RECT 499.950 145.950 502.050 148.050 ;
        RECT 488.400 138.450 489.600 138.600 ;
        RECT 482.400 137.400 489.600 138.450 ;
        RECT 466.950 133.950 469.050 136.050 ;
        RECT 469.950 133.950 472.050 136.050 ;
        RECT 472.950 133.950 475.050 136.050 ;
        RECT 475.950 133.950 478.050 136.050 ;
        RECT 470.400 131.400 471.600 133.650 ;
        RECT 476.400 132.900 477.600 133.650 ;
        RECT 470.400 127.050 471.450 131.400 ;
        RECT 475.800 130.800 477.900 132.900 ;
        RECT 478.950 130.950 481.050 133.050 ;
        RECT 476.400 127.050 477.450 130.800 ;
        RECT 463.950 124.950 466.050 127.050 ;
        RECT 469.950 124.950 472.050 127.050 ;
        RECT 475.950 124.950 478.050 127.050 ;
        RECT 460.950 61.950 463.050 64.050 ;
        RECT 464.400 61.200 465.450 124.950 ;
        RECT 469.950 118.950 472.050 121.050 ;
        RECT 470.400 105.600 471.450 118.950 ;
        RECT 479.400 118.050 480.450 130.950 ;
        RECT 478.950 115.950 481.050 118.050 ;
        RECT 470.400 103.350 471.600 105.600 ;
        RECT 475.950 104.100 478.050 106.200 ;
        RECT 482.400 106.050 483.450 137.400 ;
        RECT 488.400 136.350 489.600 137.400 ;
        RECT 494.400 136.350 495.600 138.600 ;
        RECT 499.950 137.100 502.050 139.200 ;
        RECT 503.400 139.050 504.450 154.950 ;
        RECT 500.400 136.350 501.600 137.100 ;
        RECT 502.950 136.950 505.050 139.050 ;
        RECT 487.950 133.950 490.050 136.050 ;
        RECT 490.950 133.950 493.050 136.050 ;
        RECT 493.950 133.950 496.050 136.050 ;
        RECT 496.950 133.950 499.050 136.050 ;
        RECT 499.950 133.950 502.050 136.050 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 497.400 131.400 498.600 133.650 ;
        RECT 476.400 103.350 477.600 104.100 ;
        RECT 481.950 103.950 484.050 106.050 ;
        RECT 469.950 100.950 472.050 103.050 ;
        RECT 472.950 100.950 475.050 103.050 ;
        RECT 475.950 100.950 478.050 103.050 ;
        RECT 478.950 100.950 481.050 103.050 ;
        RECT 473.400 98.400 474.600 100.650 ;
        RECT 479.400 99.900 480.600 100.650 ;
        RECT 473.400 91.050 474.450 98.400 ;
        RECT 478.950 97.800 481.050 99.900 ;
        RECT 481.950 97.950 484.050 100.050 ;
        RECT 472.950 88.950 475.050 91.050 ;
        RECT 479.400 64.050 480.450 97.800 ;
        RECT 482.400 76.050 483.450 97.950 ;
        RECT 485.400 79.050 486.450 130.950 ;
        RECT 497.400 115.050 498.450 131.400 ;
        RECT 502.950 130.950 505.050 133.050 ;
        RECT 496.950 112.950 499.050 115.050 ;
        RECT 490.950 109.800 493.050 111.900 ;
        RECT 491.400 105.600 492.450 109.800 ;
        RECT 503.400 109.050 504.450 130.950 ;
        RECT 506.400 115.050 507.450 161.400 ;
        RECT 508.950 157.950 511.050 160.050 ;
        RECT 509.400 145.050 510.450 157.950 ;
        RECT 508.950 142.950 511.050 145.050 ;
        RECT 512.400 142.050 513.450 202.950 ;
        RECT 526.950 199.950 529.050 202.050 ;
        RECT 514.950 196.950 517.050 199.050 ;
        RECT 515.400 151.050 516.450 196.950 ;
        RECT 517.950 193.950 520.050 196.050 ;
        RECT 518.400 184.050 519.450 193.950 ;
        RECT 527.400 184.200 528.450 199.950 ;
        RECT 545.400 199.050 546.450 280.950 ;
        RECT 557.400 280.050 558.450 286.950 ;
        RECT 556.950 277.950 559.050 280.050 ;
        RECT 557.400 274.050 558.450 277.950 ;
        RECT 556.950 271.950 559.050 274.050 ;
        RECT 547.950 268.950 550.050 271.050 ;
        RECT 548.400 220.050 549.450 268.950 ;
        RECT 556.950 268.800 559.050 270.900 ;
        RECT 557.400 261.600 558.450 268.800 ;
        RECT 560.400 265.050 561.450 293.100 ;
        RECT 563.400 283.050 564.450 325.950 ;
        RECT 566.400 316.050 567.450 328.650 ;
        RECT 565.950 313.950 568.050 316.050 ;
        RECT 569.400 312.450 570.450 331.950 ;
        RECT 572.400 328.050 573.450 362.400 ;
        RECT 580.950 361.950 583.050 366.000 ;
        RECT 587.400 365.400 592.050 366.450 ;
        RECT 589.950 364.950 592.050 365.400 ;
        RECT 574.950 358.950 577.050 361.050 ;
        RECT 575.400 340.050 576.450 358.950 ;
        RECT 586.950 343.950 589.050 346.050 ;
        RECT 582.000 342.450 586.050 343.050 ;
        RECT 581.400 340.950 586.050 342.450 ;
        RECT 574.950 337.950 577.050 340.050 ;
        RECT 581.400 339.600 582.450 340.950 ;
        RECT 581.400 337.350 582.600 339.600 ;
        RECT 587.400 339.450 588.450 343.950 ;
        RECT 590.400 343.050 591.450 364.950 ;
        RECT 597.150 359.700 598.350 378.300 ;
        RECT 601.950 371.100 604.050 373.200 ;
        RECT 602.400 370.350 603.600 371.100 ;
        RECT 607.950 370.950 610.050 373.050 ;
        RECT 602.100 367.950 604.200 370.050 ;
        RECT 608.400 364.050 609.450 370.950 ;
        RECT 607.950 361.950 610.050 364.050 ;
        RECT 596.850 357.600 598.950 359.700 ;
        RECT 611.400 354.450 612.450 397.950 ;
        RECT 614.400 397.050 615.450 403.950 ;
        RECT 635.400 402.450 636.450 418.950 ;
        RECT 643.950 416.100 646.050 418.200 ;
        RECT 644.400 415.350 645.600 416.100 ;
        RECT 640.950 412.950 643.050 415.050 ;
        RECT 643.950 412.950 646.050 415.050 ;
        RECT 650.400 403.050 651.450 418.950 ;
        RECT 655.950 417.000 658.050 421.050 ;
        RECT 656.400 415.350 657.600 417.000 ;
        RECT 664.950 416.100 667.050 418.200 ;
        RECT 673.950 416.100 676.050 418.200 ;
        RECT 655.950 412.950 658.050 415.050 ;
        RECT 658.950 412.950 661.050 415.050 ;
        RECT 659.400 410.400 660.600 412.650 ;
        RECT 659.400 403.050 660.450 410.400 ;
        RECT 637.950 402.450 640.050 403.050 ;
        RECT 635.400 401.400 640.050 402.450 ;
        RECT 637.950 400.950 640.050 401.400 ;
        RECT 649.950 400.950 652.050 403.050 ;
        RECT 658.950 400.950 661.050 403.050 ;
        RECT 613.950 394.950 616.050 397.050 ;
        RECT 614.550 381.300 616.650 383.400 ;
        RECT 614.550 374.700 615.750 381.300 ;
        RECT 625.950 376.950 628.050 379.050 ;
        RECT 614.550 372.600 616.650 374.700 ;
        RECT 614.550 359.700 615.750 372.600 ;
        RECT 619.950 367.950 622.050 370.050 ;
        RECT 620.400 366.450 621.600 367.650 ;
        RECT 620.400 365.400 624.450 366.450 ;
        RECT 614.550 357.600 616.650 359.700 ;
        RECT 623.400 358.050 624.450 365.400 ;
        RECT 622.950 355.950 625.050 358.050 ;
        RECT 626.400 354.450 627.450 376.950 ;
        RECT 638.400 373.200 639.450 400.950 ;
        RECT 652.950 397.950 655.050 400.050 ;
        RECT 643.950 376.950 646.050 379.050 ;
        RECT 637.950 371.100 640.050 373.200 ;
        RECT 644.400 372.600 645.450 376.950 ;
        RECT 653.400 373.050 654.450 397.950 ;
        RECT 665.400 388.050 666.450 416.100 ;
        RECT 674.400 415.350 675.600 416.100 ;
        RECT 670.950 412.950 673.050 415.050 ;
        RECT 673.950 412.950 676.050 415.050 ;
        RECT 676.950 412.950 679.050 415.050 ;
        RECT 667.950 409.950 670.050 412.050 ;
        RECT 677.400 410.400 678.600 412.650 ;
        RECT 683.400 412.050 684.450 442.800 ;
        RECT 692.400 442.050 693.450 445.950 ;
        RECT 691.950 439.950 694.050 442.050 ;
        RECT 695.400 439.050 696.450 470.400 ;
        RECT 700.950 460.950 703.050 463.050 ;
        RECT 742.950 460.950 745.050 463.050 ;
        RECT 701.400 451.200 702.450 460.950 ;
        RECT 736.950 457.950 739.050 460.050 ;
        RECT 706.950 454.950 709.050 457.050 ;
        RECT 707.400 451.200 708.450 454.950 ;
        RECT 700.950 449.100 703.050 451.200 ;
        RECT 706.950 449.100 709.050 451.200 ;
        RECT 712.950 449.100 715.050 451.200 ;
        RECT 718.950 449.100 721.050 451.200 ;
        RECT 737.400 450.600 738.450 457.950 ;
        RECT 743.400 450.600 744.450 460.950 ;
        RECT 725.400 450.450 726.600 450.600 ;
        RECT 725.400 449.400 732.450 450.450 ;
        RECT 701.400 448.350 702.600 449.100 ;
        RECT 707.400 448.350 708.600 449.100 ;
        RECT 700.950 445.950 703.050 448.050 ;
        RECT 703.950 445.950 706.050 448.050 ;
        RECT 706.950 445.950 709.050 448.050 ;
        RECT 704.400 444.000 705.600 445.650 ;
        RECT 703.950 439.950 706.050 444.000 ;
        RECT 694.950 436.950 697.050 439.050 ;
        RECT 713.400 436.050 714.450 449.100 ;
        RECT 719.400 448.350 720.600 449.100 ;
        RECT 725.400 448.350 726.600 449.400 ;
        RECT 718.950 445.950 721.050 448.050 ;
        RECT 721.950 445.950 724.050 448.050 ;
        RECT 724.950 445.950 727.050 448.050 ;
        RECT 722.400 443.400 723.600 445.650 ;
        RECT 731.400 445.050 732.450 449.400 ;
        RECT 737.400 448.350 738.600 450.600 ;
        RECT 743.400 448.350 744.600 450.600 ;
        RECT 736.950 445.950 739.050 448.050 ;
        RECT 739.950 445.950 742.050 448.050 ;
        RECT 742.950 445.950 745.050 448.050 ;
        RECT 722.400 439.050 723.450 443.400 ;
        RECT 730.950 442.950 733.050 445.050 ;
        RECT 740.400 444.900 741.600 445.650 ;
        RECT 739.950 442.800 742.050 444.900 ;
        RECT 749.400 439.050 750.450 494.100 ;
        RECT 752.400 454.050 753.450 506.400 ;
        RECT 760.950 494.100 763.050 496.200 ;
        RECT 761.400 493.350 762.600 494.100 ;
        RECT 755.100 490.950 757.200 493.050 ;
        RECT 760.500 490.950 762.600 493.050 ;
        RECT 763.800 490.950 765.900 493.050 ;
        RECT 755.400 489.900 756.600 490.650 ;
        RECT 754.950 487.800 757.050 489.900 ;
        RECT 764.400 488.400 765.600 490.650 ;
        RECT 767.400 489.900 768.450 518.400 ;
        RECT 773.400 504.450 774.450 559.950 ;
        RECT 778.950 532.950 781.050 535.050 ;
        RECT 779.400 529.200 780.450 532.950 ;
        RECT 778.950 527.100 781.050 529.200 ;
        RECT 784.950 527.100 787.050 529.200 ;
        RECT 779.400 526.350 780.600 527.100 ;
        RECT 785.400 526.350 786.600 527.100 ;
        RECT 778.950 523.950 781.050 526.050 ;
        RECT 781.950 523.950 784.050 526.050 ;
        RECT 784.950 523.950 787.050 526.050 ;
        RECT 775.950 520.950 778.050 523.050 ;
        RECT 782.400 522.900 783.600 523.650 ;
        RECT 770.400 503.400 774.450 504.450 ;
        RECT 764.400 475.050 765.450 488.400 ;
        RECT 766.950 487.800 769.050 489.900 ;
        RECT 763.950 472.950 766.050 475.050 ;
        RECT 760.950 454.950 763.050 457.050 ;
        RECT 751.950 451.950 754.050 454.050 ;
        RECT 754.950 449.100 757.050 451.200 ;
        RECT 761.400 450.600 762.450 454.950 ;
        RECT 767.400 451.050 768.450 487.800 ;
        RECT 770.400 457.050 771.450 503.400 ;
        RECT 776.400 499.050 777.450 520.950 ;
        RECT 781.950 520.800 784.050 522.900 ;
        RECT 787.950 520.950 790.050 523.050 ;
        RECT 788.400 517.050 789.450 520.950 ;
        RECT 787.950 514.950 790.050 517.050 ;
        RECT 791.400 514.050 792.450 566.400 ;
        RECT 800.400 562.050 801.450 566.400 ;
        RECT 805.950 564.450 808.050 568.050 ;
        RECT 809.400 567.450 810.450 599.400 ;
        RECT 814.950 598.800 817.050 600.900 ;
        RECT 825.150 593.700 826.350 612.300 ;
        RECT 829.950 606.000 832.050 610.050 ;
        RECT 833.400 607.050 834.450 644.400 ;
        RECT 835.950 640.950 838.050 643.050 ;
        RECT 830.400 604.350 831.600 606.000 ;
        RECT 832.950 604.950 835.050 607.050 ;
        RECT 830.100 601.950 832.200 604.050 ;
        RECT 836.400 598.050 837.450 640.950 ;
        RECT 829.950 595.950 832.050 598.050 ;
        RECT 835.950 595.950 838.050 598.050 ;
        RECT 824.850 591.600 826.950 593.700 ;
        RECT 826.950 583.950 829.050 586.050 ;
        RECT 814.950 580.950 817.050 583.050 ;
        RECT 811.950 572.100 814.050 577.050 ;
        RECT 815.400 573.600 816.450 580.950 ;
        RECT 815.400 571.350 816.600 573.600 ;
        RECT 820.950 572.100 823.050 574.200 ;
        RECT 821.400 571.350 822.600 572.100 ;
        RECT 814.950 568.950 817.050 571.050 ;
        RECT 817.950 568.950 820.050 571.050 ;
        RECT 820.950 568.950 823.050 571.050 ;
        RECT 818.400 567.900 819.600 568.650 ;
        RECT 809.400 566.400 813.450 567.450 ;
        RECT 808.950 564.450 811.050 565.050 ;
        RECT 805.950 564.000 811.050 564.450 ;
        RECT 806.400 563.400 811.050 564.000 ;
        RECT 808.950 562.950 811.050 563.400 ;
        RECT 799.950 559.950 802.050 562.050 ;
        RECT 796.950 538.950 799.050 541.050 ;
        RECT 797.400 528.600 798.450 538.950 ;
        RECT 802.950 535.950 805.050 538.050 ;
        RECT 803.400 528.600 804.450 535.950 ;
        RECT 809.400 529.050 810.450 562.950 ;
        RECT 797.400 526.350 798.600 528.600 ;
        RECT 803.400 526.350 804.600 528.600 ;
        RECT 808.950 526.950 811.050 529.050 ;
        RECT 796.950 523.950 799.050 526.050 ;
        RECT 799.950 523.950 802.050 526.050 ;
        RECT 802.950 523.950 805.050 526.050 ;
        RECT 805.950 523.950 808.050 526.050 ;
        RECT 800.400 522.900 801.600 523.650 ;
        RECT 806.400 523.050 807.600 523.650 ;
        RECT 812.400 523.050 813.450 566.400 ;
        RECT 817.950 565.800 820.050 567.900 ;
        RECT 827.400 562.050 828.450 583.950 ;
        RECT 814.950 559.950 817.050 562.050 ;
        RECT 826.950 559.950 829.050 562.050 ;
        RECT 799.950 520.800 802.050 522.900 ;
        RECT 806.400 521.400 811.050 523.050 ;
        RECT 807.000 520.950 811.050 521.400 ;
        RECT 811.950 520.950 814.050 523.050 ;
        RECT 815.400 519.450 816.450 559.950 ;
        RECT 830.400 532.050 831.450 595.950 ;
        RECT 839.400 594.450 840.450 676.950 ;
        RECT 842.400 670.050 843.450 688.950 ;
        RECT 845.400 685.050 846.450 722.400 ;
        RECT 854.400 703.050 855.450 722.400 ;
        RECT 856.950 721.950 859.050 724.050 ;
        RECT 853.950 700.950 856.050 703.050 ;
        RECT 853.950 688.950 856.050 691.050 ;
        RECT 844.950 682.950 847.050 685.050 ;
        RECT 847.950 683.100 850.050 685.200 ;
        RECT 854.400 684.600 855.450 688.950 ;
        RECT 857.400 685.050 858.450 721.950 ;
        RECT 848.400 682.350 849.600 683.100 ;
        RECT 854.400 682.350 855.600 684.600 ;
        RECT 856.950 682.950 859.050 685.050 ;
        RECT 847.950 679.950 850.050 682.050 ;
        RECT 850.950 679.950 853.050 682.050 ;
        RECT 853.950 679.950 856.050 682.050 ;
        RECT 851.400 677.400 852.600 679.650 ;
        RECT 851.400 673.050 852.450 677.400 ;
        RECT 856.950 676.950 859.050 679.050 ;
        RECT 850.950 670.950 853.050 673.050 ;
        RECT 841.950 667.950 844.050 670.050 ;
        RECT 850.950 664.950 853.050 667.050 ;
        RECT 847.950 661.950 850.050 664.050 ;
        RECT 842.550 657.300 844.650 659.400 ;
        RECT 842.550 644.400 843.750 657.300 ;
        RECT 848.400 651.600 849.450 661.950 ;
        RECT 851.400 658.050 852.450 664.950 ;
        RECT 850.800 655.950 852.900 658.050 ;
        RECT 853.950 655.950 856.050 661.050 ;
        RECT 857.400 654.450 858.450 676.950 ;
        RECT 854.400 653.400 858.450 654.450 ;
        RECT 848.400 649.350 849.600 651.600 ;
        RECT 847.950 646.950 850.050 649.050 ;
        RECT 842.550 642.300 844.650 644.400 ;
        RECT 850.950 643.950 853.050 646.050 ;
        RECT 842.550 635.700 843.750 642.300 ;
        RECT 842.550 633.600 844.650 635.700 ;
        RECT 836.400 593.400 840.450 594.450 ;
        RECT 842.550 615.300 844.650 617.400 ;
        RECT 842.550 608.700 843.750 615.300 ;
        RECT 842.550 606.600 844.650 608.700 ;
        RECT 851.400 607.050 852.450 643.950 ;
        RECT 842.550 593.700 843.750 606.600 ;
        RECT 850.950 604.950 853.050 607.050 ;
        RECT 847.950 601.950 850.050 604.050 ;
        RECT 848.400 601.050 849.600 601.650 ;
        RECT 844.950 599.400 849.600 601.050 ;
        RECT 844.950 598.950 849.000 599.400 ;
        RECT 850.950 598.950 853.050 601.050 ;
        RECT 847.950 595.950 850.050 598.050 ;
        RECT 836.400 586.050 837.450 593.400 ;
        RECT 842.550 591.600 844.650 593.700 ;
        RECT 838.950 586.950 841.050 589.050 ;
        RECT 835.950 583.950 838.050 586.050 ;
        RECT 839.400 573.600 840.450 586.950 ;
        RECT 839.400 571.350 840.600 573.600 ;
        RECT 835.950 568.950 838.050 571.050 ;
        RECT 838.950 568.950 841.050 571.050 ;
        RECT 841.950 568.950 844.050 571.050 ;
        RECT 836.400 566.400 837.600 568.650 ;
        RECT 842.400 566.400 843.600 568.650 ;
        RECT 836.400 556.050 837.450 566.400 ;
        RECT 835.950 553.950 838.050 556.050 ;
        RECT 842.400 550.050 843.450 566.400 ;
        RECT 841.950 547.950 844.050 550.050 ;
        RECT 838.950 535.950 841.050 538.050 ;
        RECT 832.950 532.950 835.050 535.050 ;
        RECT 829.950 529.950 832.050 532.050 ;
        RECT 817.950 528.600 822.000 529.050 ;
        RECT 817.950 526.950 822.600 528.600 ;
        RECT 821.400 526.350 822.600 526.950 ;
        RECT 820.950 523.950 823.050 526.050 ;
        RECT 823.950 523.950 826.050 526.050 ;
        RECT 824.400 522.900 825.600 523.650 ;
        RECT 823.950 520.800 826.050 522.900 ;
        RECT 812.400 518.400 816.450 519.450 ;
        RECT 778.950 511.950 781.050 514.050 ;
        RECT 790.950 511.950 793.050 514.050 ;
        RECT 775.950 496.950 778.050 499.050 ;
        RECT 779.400 495.600 780.450 511.950 ;
        RECT 802.950 508.950 805.050 511.050 ;
        RECT 790.950 502.950 793.050 505.050 ;
        RECT 784.950 499.950 787.050 502.050 ;
        RECT 785.400 496.200 786.450 499.950 ;
        RECT 779.400 493.350 780.600 495.600 ;
        RECT 784.950 494.100 787.050 496.200 ;
        RECT 785.400 493.350 786.600 494.100 ;
        RECT 775.950 490.950 778.050 493.050 ;
        RECT 778.950 490.950 781.050 493.050 ;
        RECT 781.950 490.950 784.050 493.050 ;
        RECT 784.950 490.950 787.050 493.050 ;
        RECT 776.400 489.450 777.600 490.650 ;
        RECT 782.400 489.900 783.600 490.650 ;
        RECT 773.400 488.400 777.600 489.450 ;
        RECT 773.400 487.050 774.450 488.400 ;
        RECT 781.950 487.800 784.050 489.900 ;
        RECT 772.950 484.950 775.050 487.050 ;
        RECT 769.950 454.950 772.050 457.050 ;
        RECT 769.950 451.800 772.050 453.900 ;
        RECT 755.400 448.350 756.600 449.100 ;
        RECT 761.400 448.350 762.600 450.600 ;
        RECT 766.950 448.950 769.050 451.050 ;
        RECT 754.950 445.950 757.050 448.050 ;
        RECT 757.950 445.950 760.050 448.050 ;
        RECT 760.950 445.950 763.050 448.050 ;
        RECT 763.950 445.950 766.050 448.050 ;
        RECT 751.950 442.950 754.050 445.050 ;
        RECT 758.400 443.400 759.600 445.650 ;
        RECT 764.400 443.400 765.600 445.650 ;
        RECT 721.950 436.950 724.050 439.050 ;
        RECT 748.950 436.950 751.050 439.050 ;
        RECT 712.950 433.950 715.050 436.050 ;
        RECT 721.950 433.800 724.050 435.900 ;
        RECT 688.950 424.950 691.050 427.050 ;
        RECT 694.950 424.950 697.050 427.050 ;
        RECT 712.950 426.450 715.050 427.050 ;
        RECT 718.950 426.450 721.050 427.050 ;
        RECT 712.950 425.400 721.050 426.450 ;
        RECT 712.950 424.950 715.050 425.400 ;
        RECT 718.950 424.950 721.050 425.400 ;
        RECT 689.400 418.200 690.450 424.950 ;
        RECT 688.950 416.100 691.050 418.200 ;
        RECT 695.400 417.600 696.450 424.950 ;
        RECT 715.950 421.950 718.050 424.050 ;
        RECT 689.400 415.350 690.600 416.100 ;
        RECT 695.400 415.350 696.600 417.600 ;
        RECT 709.950 416.100 712.050 418.200 ;
        RECT 716.400 417.600 717.450 421.950 ;
        RECT 722.400 418.050 723.450 433.800 ;
        RECT 724.950 430.950 727.050 433.050 ;
        RECT 710.400 415.350 711.600 416.100 ;
        RECT 716.400 415.350 717.600 417.600 ;
        RECT 721.950 415.950 724.050 418.050 ;
        RECT 688.950 412.950 691.050 415.050 ;
        RECT 691.950 412.950 694.050 415.050 ;
        RECT 694.950 412.950 697.050 415.050 ;
        RECT 697.950 412.950 700.050 415.050 ;
        RECT 703.950 412.950 706.050 415.050 ;
        RECT 709.950 412.950 712.050 415.050 ;
        RECT 712.950 412.950 715.050 415.050 ;
        RECT 715.950 412.950 718.050 415.050 ;
        RECT 718.950 412.950 721.050 415.050 ;
        RECT 664.950 385.950 667.050 388.050 ;
        RECT 638.400 370.350 639.600 371.100 ;
        RECT 644.400 370.350 645.600 372.600 ;
        RECT 652.950 370.950 655.050 373.050 ;
        RECT 658.950 371.100 661.050 373.200 ;
        RECT 665.400 372.450 666.600 372.600 ;
        RECT 668.400 372.450 669.450 409.950 ;
        RECT 677.400 403.050 678.450 410.400 ;
        RECT 682.950 409.950 685.050 412.050 ;
        RECT 692.400 410.400 693.600 412.650 ;
        RECT 698.400 410.400 699.600 412.650 ;
        RECT 679.950 403.950 682.050 406.050 ;
        RECT 676.950 400.950 679.050 403.050 ;
        RECT 670.950 385.950 673.050 388.050 ;
        RECT 665.400 371.400 669.450 372.450 ;
        RECT 659.400 370.350 660.600 371.100 ;
        RECT 665.400 370.350 666.600 371.400 ;
        RECT 634.950 367.950 637.050 370.050 ;
        RECT 637.950 367.950 640.050 370.050 ;
        RECT 640.950 367.950 643.050 370.050 ;
        RECT 643.950 367.950 646.050 370.050 ;
        RECT 655.950 367.950 658.050 370.050 ;
        RECT 658.950 367.950 661.050 370.050 ;
        RECT 661.950 367.950 664.050 370.050 ;
        RECT 664.950 367.950 667.050 370.050 ;
        RECT 611.400 353.400 615.450 354.450 ;
        RECT 607.950 343.950 610.050 346.050 ;
        RECT 589.950 340.950 592.050 343.050 ;
        RECT 592.950 340.950 595.050 343.050 ;
        RECT 587.400 338.400 591.450 339.450 ;
        RECT 577.950 334.950 580.050 337.050 ;
        RECT 580.950 334.950 583.050 337.050 ;
        RECT 583.950 334.950 586.050 337.050 ;
        RECT 578.400 333.000 579.600 334.650 ;
        RECT 584.400 333.450 585.600 334.650 ;
        RECT 590.400 333.450 591.450 338.400 ;
        RECT 593.400 333.900 594.450 340.950 ;
        RECT 601.950 338.100 604.050 340.200 ;
        RECT 608.400 339.600 609.450 343.950 ;
        RECT 602.400 337.350 603.600 338.100 ;
        RECT 608.400 337.350 609.600 339.600 ;
        RECT 598.950 334.950 601.050 337.050 ;
        RECT 601.950 334.950 604.050 337.050 ;
        RECT 604.950 334.950 607.050 337.050 ;
        RECT 607.950 334.950 610.050 337.050 ;
        RECT 599.400 333.900 600.600 334.650 ;
        RECT 605.400 333.900 606.600 334.650 ;
        RECT 577.950 328.950 580.050 333.000 ;
        RECT 584.400 332.400 591.450 333.450 ;
        RECT 592.950 331.800 595.050 333.900 ;
        RECT 598.950 331.800 601.050 333.900 ;
        RECT 604.950 331.800 607.050 333.900 ;
        RECT 605.400 330.450 606.450 331.800 ;
        RECT 602.400 329.400 606.450 330.450 ;
        RECT 571.950 325.950 574.050 328.050 ;
        RECT 580.950 325.950 583.050 328.050 ;
        RECT 598.950 325.950 601.050 328.050 ;
        RECT 571.950 319.950 574.050 322.050 ;
        RECT 572.400 313.050 573.450 319.950 ;
        RECT 566.400 311.400 570.450 312.450 ;
        RECT 566.400 295.200 567.450 311.400 ;
        RECT 571.950 310.950 574.050 313.050 ;
        RECT 565.950 293.100 568.050 295.200 ;
        RECT 574.950 293.100 577.050 295.200 ;
        RECT 566.400 292.350 567.600 293.100 ;
        RECT 575.400 292.350 576.600 293.100 ;
        RECT 566.100 289.950 568.200 292.050 ;
        RECT 571.500 289.950 573.600 292.050 ;
        RECT 574.800 289.950 576.900 292.050 ;
        RECT 581.400 286.050 582.450 325.950 ;
        RECT 599.400 310.050 600.450 325.950 ;
        RECT 598.950 307.950 601.050 310.050 ;
        RECT 583.950 294.600 588.000 295.050 ;
        RECT 583.950 292.950 588.600 294.600 ;
        RECT 592.950 293.100 595.050 295.200 ;
        RECT 587.400 292.350 588.600 292.950 ;
        RECT 593.400 292.350 594.600 293.100 ;
        RECT 598.950 292.950 601.050 295.050 ;
        RECT 586.950 289.950 589.050 292.050 ;
        RECT 589.950 289.950 592.050 292.050 ;
        RECT 592.950 289.950 595.050 292.050 ;
        RECT 590.400 287.400 591.600 289.650 ;
        RECT 580.950 283.950 583.050 286.050 ;
        RECT 586.950 283.950 589.050 286.050 ;
        RECT 562.950 280.950 565.050 283.050 ;
        RECT 583.950 280.950 586.050 283.050 ;
        RECT 580.950 277.950 583.050 280.050 ;
        RECT 568.950 274.950 571.050 277.050 ;
        RECT 565.950 268.950 568.050 271.050 ;
        RECT 559.950 262.950 562.050 265.050 ;
        RECT 557.400 259.350 558.600 261.600 ;
        RECT 553.950 256.950 556.050 259.050 ;
        RECT 556.950 256.950 559.050 259.050 ;
        RECT 559.950 256.950 562.050 259.050 ;
        RECT 560.400 255.900 561.600 256.650 ;
        RECT 559.950 253.800 562.050 255.900 ;
        RECT 562.950 253.950 565.050 256.050 ;
        RECT 566.400 255.900 567.450 268.950 ;
        RECT 569.400 262.050 570.450 274.950 ;
        RECT 568.950 259.950 571.050 262.050 ;
        RECT 574.950 260.100 577.050 262.200 ;
        RECT 581.400 261.600 582.450 277.950 ;
        RECT 584.400 274.050 585.450 280.950 ;
        RECT 583.950 271.950 586.050 274.050 ;
        RECT 575.400 259.350 576.600 260.100 ;
        RECT 581.400 259.350 582.600 261.600 ;
        RECT 571.950 256.950 574.050 259.050 ;
        RECT 574.950 256.950 577.050 259.050 ;
        RECT 577.950 256.950 580.050 259.050 ;
        RECT 580.950 256.950 583.050 259.050 ;
        RECT 572.400 255.900 573.600 256.650 ;
        RECT 550.950 250.950 553.050 253.050 ;
        RECT 551.400 223.050 552.450 250.950 ;
        RECT 556.950 247.950 559.050 250.050 ;
        RECT 550.950 220.950 553.050 223.050 ;
        RECT 547.950 217.950 550.050 220.050 ;
        RECT 553.950 215.100 556.050 217.200 ;
        RECT 554.400 214.350 555.600 215.100 ;
        RECT 548.400 211.950 550.500 214.050 ;
        RECT 553.800 211.950 555.900 214.050 ;
        RECT 535.950 196.950 538.050 199.050 ;
        RECT 544.950 196.950 547.050 199.050 ;
        RECT 550.950 196.950 553.050 199.050 ;
        RECT 517.800 181.950 519.900 184.050 ;
        RECT 520.950 181.950 523.050 184.050 ;
        RECT 526.950 182.100 529.050 184.200 ;
        RECT 521.400 181.350 522.600 181.950 ;
        RECT 527.400 181.350 528.600 182.100 ;
        RECT 520.950 178.950 523.050 181.050 ;
        RECT 523.950 178.950 526.050 181.050 ;
        RECT 526.950 178.950 529.050 181.050 ;
        RECT 529.950 178.950 532.050 181.050 ;
        RECT 524.400 176.400 525.600 178.650 ;
        RECT 530.400 177.900 531.600 178.650 ;
        RECT 520.950 172.950 523.050 175.050 ;
        RECT 514.950 148.950 517.050 151.050 ;
        RECT 511.950 139.950 514.050 142.050 ;
        RECT 521.400 139.200 522.450 172.950 ;
        RECT 524.400 172.050 525.450 176.400 ;
        RECT 529.950 175.800 532.050 177.900 ;
        RECT 536.400 175.050 537.450 196.950 ;
        RECT 541.950 193.950 544.050 196.050 ;
        RECT 542.400 187.050 543.450 193.950 ;
        RECT 541.950 184.950 544.050 187.050 ;
        RECT 544.950 182.100 547.050 184.200 ;
        RECT 551.400 183.600 552.450 196.950 ;
        RECT 557.400 186.450 558.450 247.950 ;
        RECT 560.400 214.050 561.450 253.800 ;
        RECT 563.400 231.450 564.450 253.950 ;
        RECT 565.950 253.800 568.050 255.900 ;
        RECT 571.950 253.800 574.050 255.900 ;
        RECT 578.400 255.000 579.600 256.650 ;
        RECT 577.950 250.950 580.050 255.000 ;
        RECT 583.950 253.950 586.050 256.050 ;
        RECT 578.400 241.050 579.450 250.950 ;
        RECT 577.950 238.950 580.050 241.050 ;
        RECT 584.400 232.050 585.450 253.950 ;
        RECT 587.400 250.050 588.450 283.950 ;
        RECT 590.400 265.050 591.450 287.400 ;
        RECT 599.400 268.050 600.450 292.950 ;
        RECT 602.400 276.450 603.450 329.400 ;
        RECT 607.950 328.950 610.050 331.050 ;
        RECT 604.950 319.950 607.050 322.050 ;
        RECT 605.400 301.050 606.450 319.950 ;
        RECT 608.400 313.050 609.450 328.950 ;
        RECT 614.400 322.050 615.450 353.400 ;
        RECT 623.400 353.400 627.450 354.450 ;
        RECT 635.400 365.400 636.600 367.650 ;
        RECT 641.400 365.400 642.600 367.650 ;
        RECT 656.400 365.400 657.600 367.650 ;
        RECT 662.400 365.400 663.600 367.650 ;
        RECT 623.400 339.600 624.450 353.400 ;
        RECT 635.400 346.050 636.450 365.400 ;
        RECT 637.950 361.950 640.050 364.050 ;
        RECT 628.950 343.950 631.050 346.050 ;
        RECT 634.950 343.950 637.050 346.050 ;
        RECT 629.400 340.050 630.450 343.950 ;
        RECT 638.400 340.050 639.450 361.950 ;
        RECT 641.400 346.050 642.450 365.400 ;
        RECT 656.400 361.050 657.450 365.400 ;
        RECT 655.950 358.950 658.050 361.050 ;
        RECT 652.950 355.950 655.050 358.050 ;
        RECT 640.950 343.950 643.050 346.050 ;
        RECT 623.400 337.350 624.600 339.600 ;
        RECT 628.950 337.950 631.050 340.050 ;
        RECT 634.950 339.600 639.450 340.050 ;
        RECT 634.950 337.950 639.600 339.600 ;
        RECT 643.950 338.100 646.050 340.200 ;
        RECT 638.400 337.350 639.600 337.950 ;
        RECT 644.400 337.350 645.600 338.100 ;
        RECT 649.950 337.950 652.050 343.050 ;
        RECT 619.950 334.950 622.050 337.050 ;
        RECT 622.950 334.950 625.050 337.050 ;
        RECT 625.950 334.950 628.050 337.050 ;
        RECT 637.950 334.950 640.050 337.050 ;
        RECT 640.950 334.950 643.050 337.050 ;
        RECT 643.950 334.950 646.050 337.050 ;
        RECT 646.950 334.950 649.050 337.050 ;
        RECT 616.950 331.950 619.050 334.050 ;
        RECT 620.400 333.000 621.600 334.650 ;
        RECT 626.400 333.900 627.600 334.650 ;
        RECT 613.950 319.950 616.050 322.050 ;
        RECT 607.950 310.950 610.050 313.050 ;
        RECT 604.950 298.950 607.050 301.050 ;
        RECT 608.400 294.600 609.450 310.950 ;
        RECT 617.400 301.050 618.450 331.950 ;
        RECT 619.950 328.950 622.050 333.000 ;
        RECT 625.950 331.800 628.050 333.900 ;
        RECT 634.950 331.950 637.050 334.050 ;
        RECT 641.400 332.400 642.600 334.650 ;
        RECT 647.400 332.400 648.600 334.650 ;
        RECT 622.950 316.950 625.050 319.050 ;
        RECT 619.950 304.950 622.050 307.050 ;
        RECT 616.950 298.950 619.050 301.050 ;
        RECT 608.400 292.350 609.600 294.600 ;
        RECT 607.950 289.950 610.050 292.050 ;
        RECT 610.950 289.950 613.050 292.050 ;
        RECT 613.950 289.950 616.050 292.050 ;
        RECT 604.950 286.950 607.050 289.050 ;
        RECT 611.400 287.400 612.600 289.650 ;
        RECT 605.400 279.450 606.450 286.950 ;
        RECT 605.400 278.400 609.450 279.450 ;
        RECT 602.400 275.400 606.450 276.450 ;
        RECT 598.950 265.950 601.050 268.050 ;
        RECT 589.950 262.950 592.050 265.050 ;
        RECT 591.000 261.900 594.000 262.050 ;
        RECT 589.950 261.600 594.000 261.900 ;
        RECT 589.950 259.950 594.600 261.600 ;
        RECT 598.950 260.100 601.050 262.200 ;
        RECT 605.400 262.050 606.450 275.400 ;
        RECT 589.950 259.800 592.050 259.950 ;
        RECT 593.400 259.350 594.600 259.950 ;
        RECT 599.400 259.350 600.600 260.100 ;
        RECT 604.950 259.950 607.050 262.050 ;
        RECT 592.950 256.950 595.050 259.050 ;
        RECT 595.950 256.950 598.050 259.050 ;
        RECT 598.950 256.950 601.050 259.050 ;
        RECT 601.950 256.950 604.050 259.050 ;
        RECT 596.400 255.900 597.600 256.650 ;
        RECT 595.950 253.800 598.050 255.900 ;
        RECT 602.400 255.000 603.600 256.650 ;
        RECT 589.950 250.950 592.050 253.050 ;
        RECT 586.950 247.950 589.050 250.050 ;
        RECT 590.400 247.050 591.450 250.950 ;
        RECT 589.950 244.950 592.050 247.050 ;
        RECT 565.950 231.450 568.050 232.050 ;
        RECT 563.400 230.400 568.050 231.450 ;
        RECT 565.950 229.950 568.050 230.400 ;
        RECT 574.950 229.950 577.050 232.050 ;
        RECT 577.950 229.950 580.050 232.050 ;
        RECT 583.950 229.950 586.050 232.050 ;
        RECT 566.400 216.600 567.450 229.950 ;
        RECT 575.400 216.600 576.450 229.950 ;
        RECT 566.400 214.350 567.600 216.600 ;
        RECT 575.400 214.350 576.600 216.600 ;
        RECT 559.950 211.950 562.050 214.050 ;
        RECT 566.100 211.950 568.200 214.050 ;
        RECT 569.400 211.950 571.500 214.050 ;
        RECT 574.800 211.950 576.900 214.050 ;
        RECT 560.400 190.050 561.450 211.950 ;
        RECT 569.400 210.900 570.600 211.650 ;
        RECT 568.950 208.800 571.050 210.900 ;
        RECT 569.400 199.050 570.450 208.800 ;
        RECT 568.950 196.950 571.050 199.050 ;
        RECT 559.950 187.950 562.050 190.050 ;
        RECT 568.950 187.950 571.050 190.050 ;
        RECT 557.400 185.400 561.450 186.450 ;
        RECT 545.400 181.350 546.600 182.100 ;
        RECT 551.400 181.350 552.600 183.600 ;
        RECT 560.400 181.050 561.450 185.400 ;
        RECT 569.400 183.600 570.450 187.950 ;
        RECT 569.400 181.350 570.600 183.600 ;
        RECT 541.950 178.950 544.050 181.050 ;
        RECT 544.950 178.950 547.050 181.050 ;
        RECT 547.950 178.950 550.050 181.050 ;
        RECT 550.950 178.950 553.050 181.050 ;
        RECT 553.950 178.950 556.050 181.050 ;
        RECT 559.950 178.950 562.050 181.050 ;
        RECT 565.950 178.950 568.050 181.050 ;
        RECT 568.950 178.950 571.050 181.050 ;
        RECT 571.950 178.950 574.050 181.050 ;
        RECT 542.400 177.900 543.600 178.650 ;
        RECT 541.950 175.800 544.050 177.900 ;
        RECT 548.400 176.400 549.600 178.650 ;
        RECT 554.400 176.400 555.600 178.650 ;
        RECT 526.950 172.950 529.050 175.050 ;
        RECT 535.950 172.950 538.050 175.050 ;
        RECT 523.950 169.950 526.050 172.050 ;
        RECT 514.950 137.100 517.050 139.200 ;
        RECT 520.950 137.100 523.050 139.200 ;
        RECT 515.400 136.350 516.600 137.100 ;
        RECT 521.400 136.350 522.600 137.100 ;
        RECT 511.950 133.950 514.050 136.050 ;
        RECT 514.950 133.950 517.050 136.050 ;
        RECT 517.950 133.950 520.050 136.050 ;
        RECT 520.950 133.950 523.050 136.050 ;
        RECT 508.950 130.950 511.050 133.050 ;
        RECT 512.400 131.400 513.600 133.650 ;
        RECT 518.400 132.000 519.600 133.650 ;
        RECT 509.400 123.450 510.450 130.950 ;
        RECT 512.400 127.050 513.450 131.400 ;
        RECT 514.950 127.950 517.050 130.050 ;
        RECT 517.950 127.950 520.050 132.000 ;
        RECT 511.950 124.950 514.050 127.050 ;
        RECT 515.400 124.050 516.450 127.950 ;
        RECT 527.400 127.050 528.450 172.950 ;
        RECT 541.950 169.950 544.050 172.050 ;
        RECT 542.400 163.050 543.450 169.950 ;
        RECT 541.950 160.950 544.050 163.050 ;
        RECT 548.400 145.050 549.450 176.400 ;
        RECT 554.400 160.050 555.450 176.400 ;
        RECT 559.950 175.800 562.050 177.900 ;
        RECT 562.950 175.950 565.050 178.050 ;
        RECT 566.400 177.900 567.600 178.650 ;
        RECT 560.400 160.050 561.450 175.800 ;
        RECT 563.400 163.050 564.450 175.950 ;
        RECT 565.950 175.800 568.050 177.900 ;
        RECT 572.400 176.400 573.600 178.650 ;
        RECT 568.950 163.950 571.050 166.050 ;
        RECT 562.950 160.950 565.050 163.050 ;
        RECT 553.950 157.950 556.050 160.050 ;
        RECT 559.950 157.950 562.050 160.050 ;
        RECT 554.400 154.050 555.450 157.950 ;
        RECT 553.950 151.950 556.050 154.050 ;
        RECT 565.950 148.950 568.050 151.050 ;
        RECT 547.950 142.950 550.050 145.050 ;
        RECT 559.950 142.950 562.050 145.050 ;
        RECT 529.950 137.100 532.050 142.050 ;
        RECT 535.950 137.100 538.050 142.050 ;
        RECT 547.950 139.800 550.050 141.900 ;
        RECT 541.950 137.100 544.050 139.200 ;
        RECT 536.400 136.350 537.600 137.100 ;
        RECT 542.400 136.350 543.600 137.100 ;
        RECT 532.950 133.950 535.050 136.050 ;
        RECT 535.950 133.950 538.050 136.050 ;
        RECT 538.950 133.950 541.050 136.050 ;
        RECT 541.950 133.950 544.050 136.050 ;
        RECT 533.400 131.400 534.600 133.650 ;
        RECT 539.400 132.900 540.600 133.650 ;
        RECT 526.950 124.950 529.050 127.050 ;
        RECT 509.400 122.400 513.450 123.450 ;
        RECT 505.800 112.950 507.900 115.050 ;
        RECT 508.950 112.950 511.050 115.050 ;
        RECT 502.950 106.950 505.050 109.050 ;
        RECT 491.400 103.350 492.600 105.600 ;
        RECT 496.950 104.100 499.050 106.200 ;
        RECT 497.400 103.350 498.600 104.100 ;
        RECT 490.950 100.950 493.050 103.050 ;
        RECT 493.950 100.950 496.050 103.050 ;
        RECT 496.950 100.950 499.050 103.050 ;
        RECT 499.950 100.950 502.050 103.050 ;
        RECT 487.950 97.950 490.050 100.050 ;
        RECT 494.400 99.900 495.600 100.650 ;
        RECT 484.950 76.950 487.050 79.050 ;
        RECT 481.950 73.950 484.050 76.050 ;
        RECT 472.950 61.950 475.050 64.050 ;
        RECT 478.950 61.950 481.050 64.050 ;
        RECT 481.950 63.450 484.050 67.050 ;
        RECT 485.400 63.450 486.450 76.950 ;
        RECT 488.400 73.050 489.450 97.950 ;
        RECT 493.950 97.800 496.050 99.900 ;
        RECT 500.400 99.000 501.600 100.650 ;
        RECT 499.950 94.950 502.050 99.000 ;
        RECT 502.950 97.950 505.050 100.050 ;
        RECT 503.400 94.050 504.450 97.950 ;
        RECT 506.400 97.050 507.450 112.950 ;
        RECT 509.400 106.050 510.450 112.950 ;
        RECT 512.400 109.050 513.450 122.400 ;
        RECT 514.950 121.950 517.050 124.050 ;
        RECT 511.950 106.950 514.050 109.050 ;
        RECT 508.950 103.950 511.050 106.050 ;
        RECT 515.400 105.600 516.450 121.950 ;
        RECT 520.950 115.950 523.050 118.050 ;
        RECT 515.400 103.350 516.600 105.600 ;
        RECT 517.950 103.950 520.050 109.050 ;
        RECT 511.950 100.950 514.050 103.050 ;
        RECT 514.950 100.950 517.050 103.050 ;
        RECT 512.400 99.900 513.600 100.650 ;
        RECT 511.950 97.800 514.050 99.900 ;
        RECT 517.950 97.950 520.050 100.050 ;
        RECT 505.950 94.950 508.050 97.050 ;
        RECT 518.400 94.050 519.450 97.950 ;
        RECT 502.950 91.950 505.050 94.050 ;
        RECT 508.950 91.950 511.050 94.050 ;
        RECT 517.950 91.950 520.050 94.050 ;
        RECT 487.950 70.950 490.050 73.050 ;
        RECT 481.950 63.000 486.450 63.450 ;
        RECT 482.400 62.400 486.450 63.000 ;
        RECT 458.400 58.350 459.600 60.600 ;
        RECT 463.950 59.100 466.050 61.200 ;
        RECT 464.400 58.350 465.600 59.100 ;
        RECT 469.950 58.950 472.050 61.050 ;
        RECT 433.950 55.950 436.050 58.050 ;
        RECT 436.950 55.950 439.050 58.050 ;
        RECT 439.950 55.950 442.050 58.050 ;
        RECT 442.950 55.950 445.050 58.050 ;
        RECT 454.950 55.950 457.050 58.050 ;
        RECT 457.950 55.950 460.050 58.050 ;
        RECT 460.950 55.950 463.050 58.050 ;
        RECT 463.950 55.950 466.050 58.050 ;
        RECT 434.400 53.400 435.600 55.650 ;
        RECT 440.400 53.400 441.600 55.650 ;
        RECT 418.950 46.950 421.050 49.050 ;
        RECT 427.950 46.950 430.050 49.050 ;
        RECT 412.950 34.950 415.050 37.050 ;
        RECT 434.400 36.450 435.450 53.400 ;
        RECT 440.400 46.050 441.450 53.400 ;
        RECT 445.950 52.950 448.050 55.050 ;
        RECT 451.800 52.950 453.900 55.050 ;
        RECT 455.400 54.900 456.600 55.650 ;
        RECT 461.400 54.900 462.600 55.650 ;
        RECT 439.950 43.950 442.050 46.050 ;
        RECT 431.400 35.400 435.450 36.450 ;
        RECT 413.400 28.050 414.450 34.950 ;
        RECT 408.000 27.600 412.050 28.050 ;
        RECT 401.400 25.350 402.600 27.600 ;
        RECT 407.400 25.950 412.050 27.600 ;
        RECT 412.950 25.950 415.050 28.050 ;
        RECT 421.950 26.100 424.050 31.050 ;
        RECT 431.400 28.050 432.450 35.400 ;
        RECT 439.950 34.950 442.050 37.050 ;
        RECT 433.950 31.950 436.050 34.050 ;
        RECT 407.400 25.350 408.600 25.950 ;
        RECT 422.400 25.350 423.600 26.100 ;
        RECT 430.950 25.950 433.050 28.050 ;
        RECT 434.400 27.600 435.450 31.950 ;
        RECT 440.400 27.600 441.450 34.950 ;
        RECT 446.400 34.050 447.450 52.950 ;
        RECT 452.400 40.050 453.450 52.950 ;
        RECT 454.950 52.800 457.050 54.900 ;
        RECT 460.950 52.800 463.050 54.900 ;
        RECT 463.950 49.950 466.050 52.050 ;
        RECT 451.950 37.950 454.050 40.050 ;
        RECT 445.950 31.950 448.050 34.050 ;
        RECT 434.400 25.350 435.600 27.600 ;
        RECT 440.400 25.350 441.600 27.600 ;
        RECT 457.950 26.100 460.050 28.200 ;
        RECT 464.400 27.600 465.450 49.950 ;
        RECT 470.400 49.050 471.450 58.950 ;
        RECT 473.400 54.900 474.450 61.950 ;
        RECT 482.400 60.600 483.450 62.400 ;
        RECT 482.400 58.350 483.600 60.600 ;
        RECT 487.950 60.000 490.050 64.050 ;
        RECT 493.950 61.950 496.050 64.050 ;
        RECT 488.400 58.350 489.600 60.000 ;
        RECT 478.950 55.950 481.050 58.050 ;
        RECT 481.950 55.950 484.050 58.050 ;
        RECT 484.950 55.950 487.050 58.050 ;
        RECT 487.950 55.950 490.050 58.050 ;
        RECT 472.950 52.800 475.050 54.900 ;
        RECT 479.400 53.400 480.600 55.650 ;
        RECT 485.400 54.900 486.600 55.650 ;
        RECT 469.950 46.950 472.050 49.050 ;
        RECT 474.000 48.900 478.050 49.050 ;
        RECT 472.950 46.950 478.050 48.900 ;
        RECT 472.950 46.800 475.050 46.950 ;
        RECT 479.400 45.450 480.450 53.400 ;
        RECT 484.950 52.800 487.050 54.900 ;
        RECT 485.400 49.050 486.450 52.800 ;
        RECT 484.950 46.950 487.050 49.050 ;
        RECT 476.400 44.400 480.450 45.450 ;
        RECT 476.400 40.050 477.450 44.400 ;
        RECT 494.400 43.050 495.450 61.950 ;
        RECT 502.950 59.100 505.050 61.200 ;
        RECT 503.400 58.350 504.600 59.100 ;
        RECT 499.950 55.950 502.050 58.050 ;
        RECT 502.950 55.950 505.050 58.050 ;
        RECT 500.400 54.000 501.600 55.650 ;
        RECT 499.950 49.950 502.050 54.000 ;
        RECT 509.400 52.050 510.450 91.950 ;
        RECT 521.400 91.050 522.450 115.950 ;
        RECT 533.400 115.050 534.450 131.400 ;
        RECT 538.950 130.800 541.050 132.900 ;
        RECT 544.950 130.950 547.050 133.050 ;
        RECT 538.950 124.950 541.050 127.050 ;
        RECT 535.950 115.950 538.050 118.050 ;
        RECT 532.950 112.950 535.050 115.050 ;
        RECT 536.400 106.200 537.450 115.950 ;
        RECT 539.400 115.050 540.450 124.950 ;
        RECT 545.400 124.050 546.450 130.950 ;
        RECT 548.400 127.050 549.450 139.800 ;
        RECT 553.950 137.100 556.050 139.200 ;
        RECT 560.400 138.600 561.450 142.950 ;
        RECT 566.400 139.050 567.450 148.950 ;
        RECT 554.400 136.350 555.600 137.100 ;
        RECT 560.400 136.350 561.600 138.600 ;
        RECT 565.950 136.950 568.050 139.050 ;
        RECT 553.950 133.950 556.050 136.050 ;
        RECT 556.950 133.950 559.050 136.050 ;
        RECT 559.950 133.950 562.050 136.050 ;
        RECT 562.950 133.950 565.050 136.050 ;
        RECT 550.950 130.950 553.050 133.050 ;
        RECT 557.400 131.400 558.600 133.650 ;
        RECT 563.400 131.400 564.600 133.650 ;
        RECT 547.950 124.950 550.050 127.050 ;
        RECT 544.950 121.950 547.050 124.050 ;
        RECT 538.950 112.950 541.050 115.050 ;
        RECT 544.950 112.950 547.050 115.050 ;
        RECT 529.950 104.100 532.050 106.200 ;
        RECT 535.950 104.100 538.050 106.200 ;
        RECT 530.400 103.350 531.600 104.100 ;
        RECT 536.400 103.350 537.600 104.100 ;
        RECT 526.950 100.950 529.050 103.050 ;
        RECT 529.950 100.950 532.050 103.050 ;
        RECT 532.950 100.950 535.050 103.050 ;
        RECT 535.950 100.950 538.050 103.050 ;
        RECT 538.950 100.950 541.050 103.050 ;
        RECT 527.400 99.000 528.600 100.650 ;
        RECT 526.950 94.950 529.050 99.000 ;
        RECT 533.400 98.400 534.600 100.650 ;
        RECT 539.400 99.900 540.600 100.650 ;
        RECT 520.950 88.950 523.050 91.050 ;
        RECT 529.950 85.950 532.050 88.050 ;
        RECT 514.950 76.950 517.050 79.050 ;
        RECT 515.400 60.600 516.450 76.950 ;
        RECT 515.400 58.350 516.600 60.600 ;
        RECT 520.950 59.100 523.050 61.200 ;
        RECT 521.400 58.350 522.600 59.100 ;
        RECT 514.950 55.950 517.050 58.050 ;
        RECT 517.950 55.950 520.050 58.050 ;
        RECT 520.950 55.950 523.050 58.050 ;
        RECT 523.950 55.950 526.050 58.050 ;
        RECT 518.400 54.900 519.600 55.650 ;
        RECT 517.950 52.800 520.050 54.900 ;
        RECT 524.400 53.400 525.600 55.650 ;
        RECT 530.400 55.050 531.450 85.950 ;
        RECT 533.400 85.050 534.450 98.400 ;
        RECT 538.950 97.800 541.050 99.900 ;
        RECT 539.400 91.050 540.450 97.800 ;
        RECT 538.950 88.950 541.050 91.050 ;
        RECT 545.400 88.050 546.450 112.950 ;
        RECT 551.400 111.450 552.450 130.950 ;
        RECT 553.950 127.950 556.050 130.050 ;
        RECT 554.400 118.050 555.450 127.950 ;
        RECT 553.950 115.950 556.050 118.050 ;
        RECT 557.400 115.050 558.450 131.400 ;
        RECT 563.400 124.050 564.450 131.400 ;
        RECT 565.950 130.950 568.050 133.050 ;
        RECT 562.950 121.950 565.050 124.050 ;
        RECT 556.950 112.950 559.050 115.050 ;
        RECT 553.950 111.450 556.050 112.050 ;
        RECT 551.400 110.400 556.050 111.450 ;
        RECT 553.950 109.950 556.050 110.400 ;
        RECT 554.400 105.600 555.450 109.950 ;
        RECT 554.400 103.350 555.600 105.600 ;
        RECT 566.400 105.450 567.450 130.950 ;
        RECT 569.400 112.050 570.450 163.950 ;
        RECT 572.400 160.050 573.450 176.400 ;
        RECT 574.950 169.950 577.050 175.050 ;
        RECT 578.400 166.050 579.450 229.950 ;
        RECT 580.950 220.950 583.050 223.050 ;
        RECT 581.400 210.900 582.450 220.950 ;
        RECT 586.950 211.950 589.050 214.050 ;
        RECT 589.950 211.950 592.050 214.050 ;
        RECT 590.400 210.900 591.600 211.650 ;
        RECT 580.950 208.800 583.050 210.900 ;
        RECT 589.950 208.800 592.050 210.900 ;
        RECT 592.950 205.950 595.050 208.050 ;
        RECT 583.950 196.950 586.050 199.050 ;
        RECT 580.950 193.950 583.050 196.050 ;
        RECT 581.400 184.050 582.450 193.950 ;
        RECT 580.950 181.950 583.050 184.050 ;
        RECT 584.400 183.600 585.450 196.950 ;
        RECT 593.400 193.050 594.450 205.950 ;
        RECT 596.400 193.050 597.450 253.800 ;
        RECT 601.950 250.950 604.050 255.000 ;
        RECT 608.400 250.050 609.450 278.400 ;
        RECT 611.400 262.200 612.450 287.400 ;
        RECT 616.950 280.950 619.050 283.050 ;
        RECT 617.400 277.050 618.450 280.950 ;
        RECT 620.400 280.050 621.450 304.950 ;
        RECT 623.400 295.050 624.450 316.950 ;
        RECT 622.950 292.950 625.050 295.050 ;
        RECT 625.950 293.100 628.050 295.200 ;
        RECT 635.400 295.050 636.450 331.950 ;
        RECT 641.400 322.050 642.450 332.400 ;
        RECT 647.400 325.050 648.450 332.400 ;
        RECT 649.950 331.950 652.050 334.050 ;
        RECT 650.400 328.050 651.450 331.950 ;
        RECT 649.950 325.950 652.050 328.050 ;
        RECT 646.950 322.950 649.050 325.050 ;
        RECT 640.950 319.950 643.050 322.050 ;
        RECT 647.400 313.050 648.450 322.950 ;
        RECT 640.950 310.950 643.050 313.050 ;
        RECT 646.950 310.950 649.050 313.050 ;
        RECT 641.400 295.050 642.450 310.950 ;
        RECT 650.400 295.050 651.450 325.950 ;
        RECT 626.400 292.350 627.600 293.100 ;
        RECT 634.800 292.950 636.900 295.050 ;
        RECT 640.950 292.950 643.050 295.050 ;
        RECT 649.950 292.950 652.050 295.050 ;
        RECT 625.950 289.950 628.050 292.050 ;
        RECT 628.950 289.950 631.050 292.050 ;
        RECT 631.950 289.950 634.050 292.050 ;
        RECT 643.950 289.950 646.050 292.050 ;
        RECT 646.950 289.950 649.050 292.050 ;
        RECT 622.950 286.950 625.050 289.050 ;
        RECT 629.400 288.900 630.600 289.650 ;
        RECT 619.950 277.950 622.050 280.050 ;
        RECT 616.950 274.950 619.050 277.050 ;
        RECT 620.400 274.050 621.450 277.950 ;
        RECT 619.950 271.950 622.050 274.050 ;
        RECT 619.950 265.950 622.050 268.050 ;
        RECT 610.950 260.100 613.050 262.200 ;
        RECT 616.950 260.100 619.050 265.050 ;
        RECT 620.400 262.050 621.450 265.950 ;
        RECT 617.400 259.350 618.600 260.100 ;
        RECT 619.950 259.950 622.050 262.050 ;
        RECT 613.950 256.950 616.050 259.050 ;
        RECT 616.950 256.950 619.050 259.050 ;
        RECT 610.950 253.950 613.050 256.050 ;
        RECT 614.400 255.900 615.600 256.650 ;
        RECT 607.950 247.950 610.050 250.050 ;
        RECT 604.950 226.950 607.050 229.050 ;
        RECT 605.400 216.600 606.450 226.950 ;
        RECT 611.400 220.050 612.450 253.950 ;
        RECT 613.950 253.800 616.050 255.900 ;
        RECT 619.950 253.950 622.050 256.050 ;
        RECT 616.950 247.950 619.050 250.050 ;
        RECT 613.950 220.950 616.050 223.050 ;
        RECT 610.950 217.950 613.050 220.050 ;
        RECT 605.400 214.350 606.600 216.600 ;
        RECT 611.400 216.450 612.600 216.600 ;
        RECT 614.400 216.450 615.450 220.950 ;
        RECT 611.400 215.400 615.450 216.450 ;
        RECT 611.400 214.350 612.600 215.400 ;
        RECT 601.950 211.950 604.050 214.050 ;
        RECT 604.950 211.950 607.050 214.050 ;
        RECT 607.950 211.950 610.050 214.050 ;
        RECT 610.950 211.950 613.050 214.050 ;
        RECT 602.400 210.000 603.600 211.650 ;
        RECT 601.950 205.950 604.050 210.000 ;
        RECT 608.400 209.400 609.600 211.650 ;
        RECT 592.800 190.950 594.900 193.050 ;
        RECT 595.950 190.950 598.050 193.050 ;
        RECT 598.950 187.950 601.050 190.050 ;
        RECT 584.400 181.350 585.600 183.600 ;
        RECT 589.950 182.100 592.050 184.200 ;
        RECT 590.400 181.350 591.600 182.100 ;
        RECT 583.950 178.950 586.050 181.050 ;
        RECT 586.950 178.950 589.050 181.050 ;
        RECT 589.950 178.950 592.050 181.050 ;
        RECT 592.950 178.950 595.050 181.050 ;
        RECT 580.950 175.800 583.050 177.900 ;
        RECT 587.400 177.000 588.600 178.650 ;
        RECT 593.400 177.900 594.600 178.650 ;
        RECT 577.950 163.950 580.050 166.050 ;
        RECT 571.950 157.950 574.050 160.050 ;
        RECT 577.950 157.950 580.050 160.050 ;
        RECT 572.400 139.050 573.450 157.950 ;
        RECT 571.950 136.950 574.050 139.050 ;
        RECT 578.400 138.600 579.450 157.950 ;
        RECT 581.400 145.050 582.450 175.800 ;
        RECT 586.950 172.950 589.050 177.000 ;
        RECT 592.950 175.800 595.050 177.900 ;
        RECT 593.400 169.050 594.450 175.800 ;
        RECT 592.950 166.950 595.050 169.050 ;
        RECT 595.950 160.950 598.050 163.050 ;
        RECT 596.400 154.050 597.450 160.950 ;
        RECT 599.400 160.050 600.450 187.950 ;
        RECT 608.400 187.200 609.450 209.400 ;
        RECT 617.400 208.050 618.450 247.950 ;
        RECT 620.400 244.050 621.450 253.950 ;
        RECT 619.950 241.950 622.050 244.050 ;
        RECT 623.400 235.050 624.450 286.950 ;
        RECT 628.950 286.800 631.050 288.900 ;
        RECT 625.950 283.950 628.050 286.050 ;
        RECT 634.950 283.950 637.050 289.050 ;
        RECT 640.950 286.950 643.050 289.050 ;
        RECT 647.400 288.900 648.600 289.650 ;
        RECT 626.400 262.050 627.450 283.950 ;
        RECT 637.950 274.800 640.050 276.900 ;
        RECT 625.950 259.950 628.050 262.050 ;
        RECT 631.950 260.100 634.050 262.200 ;
        RECT 638.400 261.600 639.450 274.800 ;
        RECT 641.400 268.050 642.450 286.950 ;
        RECT 646.950 286.800 649.050 288.900 ;
        RECT 653.400 282.450 654.450 355.950 ;
        RECT 662.400 355.050 663.450 365.400 ;
        RECT 661.950 352.950 664.050 355.050 ;
        RECT 671.400 345.450 672.450 385.950 ;
        RECT 677.400 376.050 678.450 400.950 ;
        RECT 676.950 373.950 679.050 376.050 ;
        RECT 680.400 372.600 681.450 403.950 ;
        RECT 688.950 394.950 691.050 397.050 ;
        RECT 680.400 370.350 681.600 372.600 ;
        RECT 685.950 370.950 688.050 376.050 ;
        RECT 676.950 367.950 679.050 370.050 ;
        RECT 679.950 367.950 682.050 370.050 ;
        RECT 682.950 367.950 685.050 370.050 ;
        RECT 677.400 366.000 678.600 367.650 ;
        RECT 683.400 366.900 684.600 367.650 ;
        RECT 676.950 361.950 679.050 366.000 ;
        RECT 682.950 364.800 685.050 366.900 ;
        RECT 685.950 364.950 688.050 367.050 ;
        RECT 689.400 366.450 690.450 394.950 ;
        RECT 692.400 388.050 693.450 410.400 ;
        RECT 698.400 406.050 699.450 410.400 ;
        RECT 700.950 409.950 703.050 412.050 ;
        RECT 697.950 403.950 700.050 406.050 ;
        RECT 701.400 388.050 702.450 409.950 ;
        RECT 704.400 397.050 705.450 412.950 ;
        RECT 713.400 410.400 714.600 412.650 ;
        RECT 719.400 410.400 720.600 412.650 ;
        RECT 703.950 394.950 706.050 397.050 ;
        RECT 691.950 385.950 694.050 388.050 ;
        RECT 700.950 385.950 703.050 388.050 ;
        RECT 713.400 385.050 714.450 410.400 ;
        RECT 719.400 385.050 720.450 410.400 ;
        RECT 721.950 409.950 724.050 412.050 ;
        RECT 712.950 382.950 715.050 385.050 ;
        RECT 718.950 382.950 721.050 385.050 ;
        RECT 691.950 379.950 694.050 382.050 ;
        RECT 709.950 379.950 712.050 382.050 ;
        RECT 692.400 373.050 693.450 379.950 ;
        RECT 691.950 370.950 694.050 373.050 ;
        RECT 697.950 371.100 700.050 373.200 ;
        RECT 710.400 373.050 711.450 379.950 ;
        RECT 698.400 370.350 699.600 371.100 ;
        RECT 706.950 370.950 709.050 373.050 ;
        RECT 709.950 370.950 712.050 373.050 ;
        RECT 712.950 372.000 715.050 376.050 ;
        RECT 722.400 373.050 723.450 409.950 ;
        RECT 694.950 367.950 697.050 370.050 ;
        RECT 697.950 367.950 700.050 370.050 ;
        RECT 700.950 367.950 703.050 370.050 ;
        RECT 695.400 366.900 696.600 367.650 ;
        RECT 689.400 365.400 693.450 366.450 ;
        RECT 683.400 363.450 684.450 364.800 ;
        RECT 680.400 362.400 684.450 363.450 ;
        RECT 671.400 344.400 675.450 345.450 ;
        RECT 658.950 338.100 661.050 340.200 ;
        RECT 664.950 339.000 667.050 343.050 ;
        RECT 670.950 340.950 673.050 343.050 ;
        RECT 659.400 337.350 660.600 338.100 ;
        RECT 665.400 337.350 666.600 339.000 ;
        RECT 658.950 334.950 661.050 337.050 ;
        RECT 661.950 334.950 664.050 337.050 ;
        RECT 664.950 334.950 667.050 337.050 ;
        RECT 655.950 331.950 658.050 334.050 ;
        RECT 662.400 332.400 663.600 334.650 ;
        RECT 656.400 328.050 657.450 331.950 ;
        RECT 655.950 325.950 658.050 328.050 ;
        RECT 662.400 322.050 663.450 332.400 ;
        RECT 671.400 331.050 672.450 340.950 ;
        RECT 664.950 328.950 667.050 331.050 ;
        RECT 670.950 328.950 673.050 331.050 ;
        RECT 661.950 319.950 664.050 322.050 ;
        RECT 658.950 316.950 661.050 319.050 ;
        RECT 655.950 307.950 658.050 310.050 ;
        RECT 656.400 301.050 657.450 307.950 ;
        RECT 659.400 307.050 660.450 316.950 ;
        RECT 658.950 304.950 661.050 307.050 ;
        RECT 655.950 298.950 658.050 301.050 ;
        RECT 665.400 295.200 666.450 328.950 ;
        RECT 670.950 325.800 673.050 327.900 ;
        RECT 671.400 316.050 672.450 325.800 ;
        RECT 670.950 313.950 673.050 316.050 ;
        RECT 670.950 301.950 673.050 304.050 ;
        RECT 655.950 292.950 658.050 295.050 ;
        RECT 664.950 293.100 667.050 295.200 ;
        RECT 671.400 294.600 672.450 301.950 ;
        RECT 674.400 295.050 675.450 344.400 ;
        RECT 680.400 343.050 681.450 362.400 ;
        RECT 686.400 361.050 687.450 364.950 ;
        RECT 688.950 361.950 691.050 364.050 ;
        RECT 685.950 358.950 688.050 361.050 ;
        RECT 685.950 349.950 688.050 352.050 ;
        RECT 686.400 346.050 687.450 349.950 ;
        RECT 689.400 346.050 690.450 361.950 ;
        RECT 692.400 355.050 693.450 365.400 ;
        RECT 694.950 364.800 697.050 366.900 ;
        RECT 701.400 365.400 702.600 367.650 ;
        RECT 701.400 355.050 702.450 365.400 ;
        RECT 703.950 364.950 706.050 367.050 ;
        RECT 704.400 358.050 705.450 364.950 ;
        RECT 707.400 358.050 708.450 370.950 ;
        RECT 713.400 370.350 714.600 372.000 ;
        RECT 721.950 370.950 724.050 373.050 ;
        RECT 712.950 367.950 715.050 370.050 ;
        RECT 715.950 367.950 718.050 370.050 ;
        RECT 718.950 367.950 721.050 370.050 ;
        RECT 716.400 366.900 717.600 367.650 ;
        RECT 715.950 364.800 718.050 366.900 ;
        RECT 725.400 364.050 726.450 430.950 ;
        RECT 733.950 424.950 739.050 427.050 ;
        RECT 752.400 424.050 753.450 442.950 ;
        RECT 758.400 439.050 759.450 443.400 ;
        RECT 760.950 439.950 763.050 442.050 ;
        RECT 757.950 436.950 760.050 439.050 ;
        RECT 757.950 424.950 760.050 427.050 ;
        RECT 736.950 421.050 739.050 423.900 ;
        RECT 742.950 421.950 745.050 424.050 ;
        RECT 736.950 420.000 742.050 421.050 ;
        RECT 737.400 419.400 742.050 420.000 ;
        RECT 738.000 418.950 742.050 419.400 ;
        RECT 730.950 416.100 733.050 418.200 ;
        RECT 731.400 415.350 732.600 416.100 ;
        RECT 730.950 412.950 733.050 415.050 ;
        RECT 733.950 412.950 736.050 415.050 ;
        RECT 734.400 412.050 735.600 412.650 ;
        RECT 727.950 409.950 730.050 412.050 ;
        RECT 734.400 411.900 738.000 412.050 ;
        RECT 734.400 410.400 739.050 411.900 ;
        RECT 743.400 411.450 744.450 421.950 ;
        RECT 745.950 420.450 748.050 424.050 ;
        RECT 751.950 421.950 754.050 424.050 ;
        RECT 745.950 420.000 750.450 420.450 ;
        RECT 746.400 419.400 750.450 420.000 ;
        RECT 749.400 417.600 750.450 419.400 ;
        RECT 749.400 415.350 750.600 417.600 ;
        RECT 746.100 412.950 748.200 415.050 ;
        RECT 749.400 412.950 751.500 415.050 ;
        RECT 754.800 412.950 756.900 415.050 ;
        RECT 746.400 411.450 747.600 412.650 ;
        RECT 743.400 410.400 747.600 411.450 ;
        RECT 755.400 411.000 756.600 412.650 ;
        RECT 735.000 409.950 739.050 410.400 ;
        RECT 728.400 406.050 729.450 409.950 ;
        RECT 736.950 409.800 739.050 409.950 ;
        RECT 754.950 406.950 757.050 411.000 ;
        RECT 727.950 403.950 730.050 406.050 ;
        RECT 745.950 394.950 748.050 397.050 ;
        RECT 742.950 385.950 745.050 388.050 ;
        RECT 736.950 382.950 739.050 385.050 ;
        RECT 730.950 379.950 733.050 382.050 ;
        RECT 731.400 372.600 732.450 379.950 ;
        RECT 737.400 373.200 738.450 382.950 ;
        RECT 731.400 370.350 732.600 372.600 ;
        RECT 736.950 371.100 739.050 373.200 ;
        RECT 743.400 373.050 744.450 385.950 ;
        RECT 737.400 370.350 738.600 371.100 ;
        RECT 742.950 370.950 745.050 373.050 ;
        RECT 730.950 367.950 733.050 370.050 ;
        RECT 733.950 367.950 736.050 370.050 ;
        RECT 736.950 367.950 739.050 370.050 ;
        RECT 739.950 367.950 742.050 370.050 ;
        RECT 709.950 361.950 712.050 364.050 ;
        RECT 724.950 361.950 727.050 364.050 ;
        RECT 727.950 363.450 730.050 367.050 ;
        RECT 734.400 365.400 735.600 367.650 ;
        RECT 740.400 365.400 741.600 367.650 ;
        RECT 727.950 363.000 732.450 363.450 ;
        RECT 728.400 362.400 732.450 363.000 ;
        RECT 703.800 355.950 705.900 358.050 ;
        RECT 706.950 355.950 709.050 358.050 ;
        RECT 691.950 352.950 694.050 355.050 ;
        RECT 700.950 352.950 703.050 355.050 ;
        RECT 682.950 344.400 687.450 346.050 ;
        RECT 682.950 343.950 687.000 344.400 ;
        RECT 688.950 343.950 691.050 346.050 ;
        RECT 679.950 340.950 682.050 343.050 ;
        RECT 682.950 338.100 685.050 340.200 ;
        RECT 683.400 337.350 684.600 338.100 ;
        RECT 679.950 334.950 682.050 337.050 ;
        RECT 682.950 334.950 685.050 337.050 ;
        RECT 685.950 334.950 688.050 337.050 ;
        RECT 680.400 332.400 681.600 334.650 ;
        RECT 680.400 319.050 681.450 332.400 ;
        RECT 688.950 331.950 691.050 334.050 ;
        RECT 685.950 322.800 688.050 324.900 ;
        RECT 679.950 316.950 682.050 319.050 ;
        RECT 680.400 307.050 681.450 316.950 ;
        RECT 679.950 304.950 682.050 307.050 ;
        RECT 686.400 304.050 687.450 322.800 ;
        RECT 689.400 319.050 690.450 331.950 ;
        RECT 688.950 316.950 691.050 319.050 ;
        RECT 688.950 307.950 691.050 310.050 ;
        RECT 689.400 304.050 690.450 307.950 ;
        RECT 685.950 301.950 688.050 304.050 ;
        RECT 688.950 301.950 691.050 304.050 ;
        RECT 656.400 286.050 657.450 292.950 ;
        RECT 665.400 292.350 666.600 293.100 ;
        RECT 671.400 292.350 672.600 294.600 ;
        RECT 673.950 292.950 676.050 295.050 ;
        RECT 682.950 293.100 685.050 295.200 ;
        RECT 688.950 294.000 691.050 298.050 ;
        RECT 692.400 294.450 693.450 352.950 ;
        RECT 700.950 349.800 703.050 351.900 ;
        RECT 694.950 343.950 697.050 346.050 ;
        RECT 695.400 325.050 696.450 343.950 ;
        RECT 701.400 340.200 702.450 349.800 ;
        RECT 700.950 338.100 703.050 340.200 ;
        RECT 701.400 337.350 702.600 338.100 ;
        RECT 698.100 334.950 700.200 337.050 ;
        RECT 701.400 334.950 703.500 337.050 ;
        RECT 706.800 334.950 708.900 337.050 ;
        RECT 698.400 332.400 699.600 334.650 ;
        RECT 707.400 333.900 708.600 334.650 ;
        RECT 698.400 325.050 699.450 332.400 ;
        RECT 706.950 331.800 709.050 333.900 ;
        RECT 694.950 322.950 697.050 325.050 ;
        RECT 697.950 322.950 700.050 325.050 ;
        RECT 710.400 315.450 711.450 361.950 ;
        RECT 712.950 338.100 715.050 340.200 ;
        RECT 721.950 338.100 724.050 340.200 ;
        RECT 727.950 338.100 730.050 340.200 ;
        RECT 731.400 340.050 732.450 362.400 ;
        RECT 734.400 361.050 735.450 365.400 ;
        RECT 733.950 358.950 736.050 361.050 ;
        RECT 740.400 352.050 741.450 365.400 ;
        RECT 746.400 364.050 747.450 394.950 ;
        RECT 758.400 379.050 759.450 424.950 ;
        RECT 761.400 409.050 762.450 439.950 ;
        RECT 764.400 412.050 765.450 443.400 ;
        RECT 770.400 433.050 771.450 451.800 ;
        RECT 773.400 442.050 774.450 484.950 ;
        RECT 782.400 481.050 783.450 487.800 ;
        RECT 787.950 481.950 790.050 484.050 ;
        RECT 781.950 478.950 784.050 481.050 ;
        RECT 781.950 454.950 784.050 457.050 ;
        RECT 782.400 450.600 783.450 454.950 ;
        RECT 782.400 448.350 783.600 450.600 ;
        RECT 778.950 445.950 781.050 448.050 ;
        RECT 781.950 445.950 784.050 448.050 ;
        RECT 779.400 443.400 780.600 445.650 ;
        RECT 788.400 444.450 789.450 481.950 ;
        RECT 791.400 475.050 792.450 502.950 ;
        RECT 796.950 494.100 799.050 496.200 ;
        RECT 803.400 495.600 804.450 508.950 ;
        RECT 797.400 493.350 798.600 494.100 ;
        RECT 803.400 493.350 804.600 495.600 ;
        RECT 796.950 490.950 799.050 493.050 ;
        RECT 799.950 490.950 802.050 493.050 ;
        RECT 802.950 490.950 805.050 493.050 ;
        RECT 805.950 490.950 808.050 493.050 ;
        RECT 800.400 489.000 801.600 490.650 ;
        RECT 799.950 484.950 802.050 489.000 ;
        RECT 806.400 488.400 807.600 490.650 ;
        RECT 790.950 472.950 793.050 475.050 ;
        RECT 806.400 454.050 807.450 488.400 ;
        RECT 808.950 487.800 811.050 489.900 ;
        RECT 796.950 450.000 799.050 454.050 ;
        RECT 805.950 451.950 808.050 454.050 ;
        RECT 797.400 448.350 798.600 450.000 ;
        RECT 802.950 449.100 805.050 451.200 ;
        RECT 803.400 448.350 804.600 449.100 ;
        RECT 793.950 445.950 796.050 448.050 ;
        RECT 796.950 445.950 799.050 448.050 ;
        RECT 799.950 445.950 802.050 448.050 ;
        RECT 802.950 445.950 805.050 448.050 ;
        RECT 785.400 443.400 789.450 444.450 ;
        RECT 794.400 443.400 795.600 445.650 ;
        RECT 800.400 444.000 801.600 445.650 ;
        RECT 772.950 439.950 775.050 442.050 ;
        RECT 769.950 430.950 772.050 433.050 ;
        RECT 766.950 420.450 769.050 421.050 ;
        RECT 772.950 420.450 775.050 421.050 ;
        RECT 766.950 419.400 775.050 420.450 ;
        RECT 766.950 418.950 769.050 419.400 ;
        RECT 772.950 418.950 775.050 419.400 ;
        RECT 769.950 416.100 772.050 418.200 ;
        RECT 770.400 415.350 771.600 416.100 ;
        RECT 767.100 412.950 769.200 415.050 ;
        RECT 770.400 412.950 772.500 415.050 ;
        RECT 775.800 412.950 777.900 415.050 ;
        RECT 763.950 409.950 766.050 412.050 ;
        RECT 767.400 411.900 768.600 412.650 ;
        RECT 776.400 411.900 777.600 412.650 ;
        RECT 779.400 412.050 780.450 443.400 ;
        RECT 781.950 439.950 784.050 442.050 ;
        RECT 766.950 409.800 769.050 411.900 ;
        RECT 775.950 409.800 778.050 411.900 ;
        RECT 778.950 409.950 781.050 412.050 ;
        RECT 760.950 406.950 763.050 409.050 ;
        RECT 769.950 406.950 772.050 409.050 ;
        RECT 760.950 397.950 763.050 400.050 ;
        RECT 748.950 376.950 751.050 379.050 ;
        RECT 757.950 376.950 760.050 379.050 ;
        RECT 745.950 361.950 748.050 364.050 ;
        RECT 739.950 349.950 742.050 352.050 ;
        RECT 733.950 346.950 736.050 349.050 ;
        RECT 713.400 319.050 714.450 338.100 ;
        RECT 722.400 337.350 723.600 338.100 ;
        RECT 728.400 337.350 729.600 338.100 ;
        RECT 730.950 337.950 733.050 340.050 ;
        RECT 718.950 334.950 721.050 337.050 ;
        RECT 721.950 334.950 724.050 337.050 ;
        RECT 724.950 334.950 727.050 337.050 ;
        RECT 727.950 334.950 730.050 337.050 ;
        RECT 719.400 332.400 720.600 334.650 ;
        RECT 725.400 333.900 726.600 334.650 ;
        RECT 719.400 322.050 720.450 332.400 ;
        RECT 724.950 331.800 727.050 333.900 ;
        RECT 730.950 331.950 733.050 334.050 ;
        RECT 718.950 319.950 721.050 322.050 ;
        RECT 712.950 316.950 715.050 319.050 ;
        RECT 710.400 314.400 714.450 315.450 ;
        RECT 703.950 304.950 706.050 307.050 ;
        RECT 694.950 301.950 700.050 304.050 ;
        RECT 700.950 298.950 703.050 301.050 ;
        RECT 701.400 295.200 702.450 298.950 ;
        RECT 704.400 298.050 705.450 304.950 ;
        RECT 703.950 295.950 706.050 298.050 ;
        RECT 683.400 292.350 684.600 293.100 ;
        RECT 689.400 292.350 690.600 294.000 ;
        RECT 692.400 293.400 696.450 294.450 ;
        RECT 661.950 289.950 664.050 292.050 ;
        RECT 664.950 289.950 667.050 292.050 ;
        RECT 667.950 289.950 670.050 292.050 ;
        RECT 670.950 289.950 673.050 292.050 ;
        RECT 676.950 289.800 679.050 291.900 ;
        RECT 682.950 289.950 685.050 292.050 ;
        RECT 685.950 289.950 688.050 292.050 ;
        RECT 688.950 289.950 691.050 292.050 ;
        RECT 662.400 288.000 663.600 289.650 ;
        RECT 668.400 288.000 669.600 289.650 ;
        RECT 655.950 283.950 658.050 286.050 ;
        RECT 661.950 283.950 664.050 288.000 ;
        RECT 667.950 283.950 670.050 288.000 ;
        RECT 673.950 286.950 676.050 289.050 ;
        RECT 653.400 281.400 657.450 282.450 ;
        RECT 643.950 271.950 646.050 274.050 ;
        RECT 640.950 265.950 643.050 268.050 ;
        RECT 632.400 259.350 633.600 260.100 ;
        RECT 638.400 259.350 639.600 261.600 ;
        RECT 640.950 260.100 643.050 264.900 ;
        RECT 628.950 256.950 631.050 259.050 ;
        RECT 631.950 256.950 634.050 259.050 ;
        RECT 634.950 256.950 637.050 259.050 ;
        RECT 637.950 256.950 640.050 259.050 ;
        RECT 625.800 253.950 627.900 256.050 ;
        RECT 629.400 255.900 630.600 256.650 ;
        RECT 622.950 232.950 625.050 235.050 ;
        RECT 626.400 232.050 627.450 253.950 ;
        RECT 628.950 253.800 631.050 255.900 ;
        RECT 635.400 254.400 636.600 256.650 ;
        RECT 631.950 247.950 634.050 253.050 ;
        RECT 635.400 250.050 636.450 254.400 ;
        RECT 644.400 250.050 645.450 271.950 ;
        RECT 656.400 265.050 657.450 281.400 ;
        RECT 670.950 280.950 673.050 283.050 ;
        RECT 661.950 274.950 664.050 277.050 ;
        RECT 646.950 259.950 649.050 265.050 ;
        RECT 655.950 262.950 658.050 265.050 ;
        RECT 652.950 260.100 655.050 262.200 ;
        RECT 658.950 260.100 661.050 262.200 ;
        RECT 662.400 262.050 663.450 274.950 ;
        RECT 671.400 268.050 672.450 280.950 ;
        RECT 670.950 265.950 673.050 268.050 ;
        RECT 674.400 264.450 675.450 286.950 ;
        RECT 677.400 283.050 678.450 289.800 ;
        RECT 686.400 287.400 687.600 289.650 ;
        RECT 676.950 280.950 679.050 283.050 ;
        RECT 682.950 280.950 685.050 283.050 ;
        RECT 671.400 263.400 675.450 264.450 ;
        RECT 653.400 259.350 654.600 260.100 ;
        RECT 659.400 259.350 660.600 260.100 ;
        RECT 661.950 259.950 664.050 262.050 ;
        RECT 671.400 261.600 672.450 263.400 ;
        RECT 671.400 259.350 672.600 261.600 ;
        RECT 676.950 260.100 679.050 262.200 ;
        RECT 677.400 259.350 678.600 260.100 ;
        RECT 649.950 256.950 652.050 259.050 ;
        RECT 652.950 256.950 655.050 259.050 ;
        RECT 655.950 256.950 658.050 259.050 ;
        RECT 658.950 256.950 661.050 259.050 ;
        RECT 670.950 256.950 673.050 259.050 ;
        RECT 673.950 256.950 676.050 259.050 ;
        RECT 676.950 256.950 679.050 259.050 ;
        RECT 650.400 254.400 651.600 256.650 ;
        RECT 656.400 254.400 657.600 256.650 ;
        RECT 634.950 247.950 637.050 250.050 ;
        RECT 643.950 247.950 646.050 250.050 ;
        RECT 650.400 244.050 651.450 254.400 ;
        RECT 656.400 247.050 657.450 254.400 ;
        RECT 661.950 253.950 664.050 256.050 ;
        RECT 667.950 253.950 670.050 256.050 ;
        RECT 674.400 254.400 675.600 256.650 ;
        RECT 655.950 244.950 658.050 247.050 ;
        RECT 649.950 241.950 652.050 244.050 ;
        RECT 637.950 235.950 640.050 238.050 ;
        RECT 625.950 229.950 628.050 232.050 ;
        RECT 631.950 220.950 634.050 223.050 ;
        RECT 625.950 215.100 628.050 217.200 ;
        RECT 626.400 214.350 627.600 215.100 ;
        RECT 622.950 211.950 625.050 214.050 ;
        RECT 625.950 211.950 628.050 214.050 ;
        RECT 623.400 211.050 624.600 211.650 ;
        RECT 619.950 210.900 624.600 211.050 ;
        RECT 619.950 208.950 625.050 210.900 ;
        RECT 616.950 205.950 619.050 208.050 ;
        RECT 616.950 199.950 619.050 202.050 ;
        RECT 607.950 185.100 610.050 187.200 ;
        RECT 617.400 187.050 618.450 199.950 ;
        RECT 620.400 199.050 621.450 208.950 ;
        RECT 622.950 208.800 625.050 208.950 ;
        RECT 632.400 208.050 633.450 220.950 ;
        RECT 634.800 215.100 636.900 217.200 ;
        RECT 638.400 217.050 639.450 235.950 ;
        RECT 649.950 235.800 652.050 237.900 ;
        RECT 643.950 226.950 646.050 229.050 ;
        RECT 622.950 205.650 625.050 207.750 ;
        RECT 631.950 205.950 634.050 208.050 ;
        RECT 619.950 196.950 622.050 199.050 ;
        RECT 619.950 187.950 622.050 190.050 ;
        RECT 616.950 184.950 619.050 187.050 ;
        RECT 607.950 181.950 610.050 184.050 ;
        RECT 613.950 182.100 616.050 184.200 ;
        RECT 608.400 181.350 609.600 181.950 ;
        RECT 614.400 181.350 615.600 182.100 ;
        RECT 604.950 178.950 607.050 181.050 ;
        RECT 607.950 178.950 610.050 181.050 ;
        RECT 610.950 178.950 613.050 181.050 ;
        RECT 613.950 178.950 616.050 181.050 ;
        RECT 605.400 178.050 606.600 178.650 ;
        RECT 601.950 176.400 606.600 178.050 ;
        RECT 611.400 176.400 612.600 178.650 ;
        RECT 601.950 175.950 606.000 176.400 ;
        RECT 607.950 172.950 610.050 175.050 ;
        RECT 598.950 157.950 601.050 160.050 ;
        RECT 583.950 151.950 586.050 154.050 ;
        RECT 595.950 151.950 598.050 154.050 ;
        RECT 580.950 142.950 583.050 145.050 ;
        RECT 584.400 138.600 585.450 151.950 ;
        RECT 589.950 145.950 592.050 148.050 ;
        RECT 578.400 136.350 579.600 138.600 ;
        RECT 584.400 136.350 585.600 138.600 ;
        RECT 574.950 133.950 577.050 136.050 ;
        RECT 577.950 133.950 580.050 136.050 ;
        RECT 580.950 133.950 583.050 136.050 ;
        RECT 583.950 133.950 586.050 136.050 ;
        RECT 575.400 132.000 576.600 133.650 ;
        RECT 581.400 132.900 582.600 133.650 ;
        RECT 590.400 132.900 591.450 145.950 ;
        RECT 592.950 142.950 595.050 145.050 ;
        RECT 593.400 139.050 594.450 142.950 ;
        RECT 592.950 136.950 595.050 139.050 ;
        RECT 596.400 138.600 597.450 151.950 ;
        RECT 596.400 136.350 597.600 138.600 ;
        RECT 595.950 133.950 598.050 136.050 ;
        RECT 598.950 133.950 601.050 136.050 ;
        RECT 601.950 133.950 604.050 136.050 ;
        RECT 599.400 132.900 600.600 133.650 ;
        RECT 574.950 127.950 577.050 132.000 ;
        RECT 580.950 130.800 583.050 132.900 ;
        RECT 589.800 130.800 591.900 132.900 ;
        RECT 598.950 130.800 601.050 132.900 ;
        RECT 571.950 121.950 574.050 124.050 ;
        RECT 568.950 109.950 571.050 112.050 ;
        RECT 563.400 104.400 567.450 105.450 ;
        RECT 572.400 105.600 573.450 121.950 ;
        RECT 580.950 118.950 583.050 121.050 ;
        RECT 550.950 100.950 553.050 103.050 ;
        RECT 553.950 100.950 556.050 103.050 ;
        RECT 556.950 100.950 559.050 103.050 ;
        RECT 551.400 99.900 552.600 100.650 ;
        RECT 557.400 99.900 558.600 100.650 ;
        RECT 550.950 97.800 553.050 99.900 ;
        RECT 556.950 97.800 559.050 99.900 ;
        RECT 544.950 85.950 547.050 88.050 ;
        RECT 532.950 82.950 535.050 85.050 ;
        RECT 535.950 60.000 538.050 64.050 ;
        RECT 563.400 61.200 564.450 104.400 ;
        RECT 572.400 103.350 573.600 105.600 ;
        RECT 568.950 100.950 571.050 103.050 ;
        RECT 571.950 100.950 574.050 103.050 ;
        RECT 574.950 100.950 577.050 103.050 ;
        RECT 569.400 98.400 570.600 100.650 ;
        RECT 581.400 99.900 582.450 118.950 ;
        RECT 601.950 112.950 604.050 115.050 ;
        RECT 598.950 109.950 601.050 112.050 ;
        RECT 589.950 104.100 592.050 106.200 ;
        RECT 590.400 103.350 591.600 104.100 ;
        RECT 586.950 100.950 589.050 103.050 ;
        RECT 589.950 100.950 592.050 103.050 ;
        RECT 592.950 100.950 595.050 103.050 ;
        RECT 587.400 99.900 588.600 100.650 ;
        RECT 569.400 76.050 570.450 98.400 ;
        RECT 580.950 97.800 583.050 99.900 ;
        RECT 586.950 97.800 589.050 99.900 ;
        RECT 593.400 99.000 594.600 100.650 ;
        RECT 592.950 94.950 595.050 99.000 ;
        RECT 595.950 97.950 598.050 100.050 ;
        RECT 596.400 88.050 597.450 97.950 ;
        RECT 599.400 97.050 600.450 109.950 ;
        RECT 602.400 99.900 603.450 112.950 ;
        RECT 608.400 112.050 609.450 172.950 ;
        RECT 611.400 154.050 612.450 176.400 ;
        RECT 610.950 151.950 613.050 154.050 ;
        RECT 611.400 139.050 612.450 151.950 ;
        RECT 610.950 136.950 613.050 139.050 ;
        RECT 616.950 137.100 619.050 139.200 ;
        RECT 620.400 138.450 621.450 187.950 ;
        RECT 623.400 177.450 624.450 205.650 ;
        RECT 628.950 199.950 631.050 202.050 ;
        RECT 629.400 193.050 630.450 199.950 ;
        RECT 635.400 199.050 636.450 215.100 ;
        RECT 637.950 214.950 640.050 217.050 ;
        RECT 644.400 216.600 645.450 226.950 ;
        RECT 650.400 223.050 651.450 235.800 ;
        RECT 656.400 232.050 657.450 244.950 ;
        RECT 662.400 238.050 663.450 253.950 ;
        RECT 668.400 250.050 669.450 253.950 ;
        RECT 670.950 250.950 673.050 253.050 ;
        RECT 667.950 247.950 670.050 250.050 ;
        RECT 661.950 235.950 664.050 238.050 ;
        RECT 658.950 232.950 661.050 235.050 ;
        RECT 652.800 229.950 654.900 232.050 ;
        RECT 655.950 229.950 658.050 232.050 ;
        RECT 649.950 220.950 652.050 223.050 ;
        RECT 644.400 214.350 645.600 216.600 ;
        RECT 649.950 216.000 652.050 219.900 ;
        RECT 653.400 217.050 654.450 229.950 ;
        RECT 655.950 225.450 658.050 226.050 ;
        RECT 659.400 225.450 660.450 232.950 ;
        RECT 661.950 226.950 664.050 229.050 ;
        RECT 655.950 224.400 660.450 225.450 ;
        RECT 655.950 223.950 658.050 224.400 ;
        RECT 650.400 214.350 651.600 216.000 ;
        RECT 652.950 214.950 655.050 217.050 ;
        RECT 640.950 211.950 643.050 214.050 ;
        RECT 643.950 211.950 646.050 214.050 ;
        RECT 646.950 211.950 649.050 214.050 ;
        RECT 649.950 211.950 652.050 214.050 ;
        RECT 641.400 210.900 642.600 211.650 ;
        RECT 640.950 208.800 643.050 210.900 ;
        RECT 647.400 209.400 648.600 211.650 ;
        RECT 637.950 199.950 640.050 205.050 ;
        RECT 640.950 202.950 643.050 205.050 ;
        RECT 634.950 196.950 637.050 199.050 ;
        RECT 628.950 190.950 631.050 193.050 ;
        RECT 629.400 183.600 630.450 190.950 ;
        RECT 629.400 181.350 630.600 183.600 ;
        RECT 626.100 178.950 628.200 181.050 ;
        RECT 629.400 178.950 631.500 181.050 ;
        RECT 634.800 178.950 636.900 181.050 ;
        RECT 626.400 177.900 627.600 178.650 ;
        RECT 625.950 177.450 628.050 177.900 ;
        RECT 623.400 176.400 628.050 177.450 ;
        RECT 635.400 177.000 636.600 178.650 ;
        RECT 625.950 175.800 628.050 176.400 ;
        RECT 634.950 172.950 637.050 177.000 ;
        RECT 641.400 163.050 642.450 202.950 ;
        RECT 643.950 196.950 646.050 199.050 ;
        RECT 644.400 184.050 645.450 196.950 ;
        RECT 647.400 193.050 648.450 209.400 ;
        RECT 656.400 205.050 657.450 223.950 ;
        RECT 662.400 223.050 663.450 226.950 ;
        RECT 671.400 223.050 672.450 250.950 ;
        RECT 674.400 244.050 675.450 254.400 ;
        RECT 673.950 241.950 676.050 244.050 ;
        RECT 673.950 235.950 676.050 238.050 ;
        RECT 661.950 220.950 664.050 223.050 ;
        RECT 670.950 220.950 673.050 223.050 ;
        RECT 661.950 215.100 664.050 217.200 ;
        RECT 662.400 214.350 663.600 215.100 ;
        RECT 661.950 211.950 664.050 214.050 ;
        RECT 664.950 211.950 667.050 214.050 ;
        RECT 667.950 211.950 670.050 214.050 ;
        RECT 658.950 208.950 661.050 211.050 ;
        RECT 665.400 210.900 666.600 211.650 ;
        RECT 655.950 202.950 658.050 205.050 ;
        RECT 646.950 190.950 649.050 193.050 ;
        RECT 643.950 181.950 646.050 184.050 ;
        RECT 649.950 182.100 652.050 184.200 ;
        RECT 650.400 181.350 651.600 182.100 ;
        RECT 646.950 178.950 649.050 181.050 ;
        RECT 649.950 178.950 652.050 181.050 ;
        RECT 652.950 178.950 655.050 181.050 ;
        RECT 647.400 177.900 648.600 178.650 ;
        RECT 646.950 175.800 649.050 177.900 ;
        RECT 653.400 176.400 654.600 178.650 ;
        RECT 653.400 169.050 654.450 176.400 ;
        RECT 655.950 175.950 658.050 178.050 ;
        RECT 656.400 172.050 657.450 175.950 ;
        RECT 655.950 169.950 658.050 172.050 ;
        RECT 652.950 166.950 655.050 169.050 ;
        RECT 643.950 163.950 646.050 166.050 ;
        RECT 640.950 160.950 643.050 163.050 ;
        RECT 631.950 148.950 634.050 151.050 ;
        RECT 632.400 145.050 633.450 148.950 ;
        RECT 631.950 142.950 634.050 145.050 ;
        RECT 620.400 137.400 624.450 138.450 ;
        RECT 617.400 136.350 618.600 137.100 ;
        RECT 613.950 133.950 616.050 136.050 ;
        RECT 616.950 133.950 619.050 136.050 ;
        RECT 614.400 132.900 615.600 133.650 ;
        RECT 613.950 130.800 616.050 132.900 ;
        RECT 623.400 121.050 624.450 137.400 ;
        RECT 631.950 137.100 634.050 139.200 ;
        RECT 637.950 138.000 640.050 142.050 ;
        RECT 632.400 136.350 633.600 137.100 ;
        RECT 638.400 136.350 639.600 138.000 ;
        RECT 628.950 133.950 631.050 136.050 ;
        RECT 631.950 133.950 634.050 136.050 ;
        RECT 634.950 133.950 637.050 136.050 ;
        RECT 637.950 133.950 640.050 136.050 ;
        RECT 629.400 131.400 630.600 133.650 ;
        RECT 635.400 132.900 636.600 133.650 ;
        RECT 622.950 118.950 625.050 121.050 ;
        RECT 607.950 109.950 610.050 112.050 ;
        RECT 622.950 109.950 625.050 112.050 ;
        RECT 610.950 104.100 613.050 106.200 ;
        RECT 616.950 104.100 619.050 106.200 ;
        RECT 611.400 103.350 612.600 104.100 ;
        RECT 617.400 103.350 618.600 104.100 ;
        RECT 607.950 100.950 610.050 103.050 ;
        RECT 610.950 100.950 613.050 103.050 ;
        RECT 613.950 100.950 616.050 103.050 ;
        RECT 616.950 100.950 619.050 103.050 ;
        RECT 608.400 99.900 609.600 100.650 ;
        RECT 601.950 97.800 604.050 99.900 ;
        RECT 607.950 97.800 610.050 99.900 ;
        RECT 614.400 99.000 615.600 100.650 ;
        RECT 598.950 94.950 601.050 97.050 ;
        RECT 613.950 94.950 616.050 99.000 ;
        RECT 619.950 97.950 622.050 100.050 ;
        RECT 599.400 91.050 600.450 94.950 ;
        RECT 598.950 88.950 601.050 91.050 ;
        RECT 595.950 85.950 598.050 88.050 ;
        RECT 568.950 73.950 571.050 76.050 ;
        RECT 620.400 73.050 621.450 97.950 ;
        RECT 623.400 97.050 624.450 109.950 ;
        RECT 629.400 106.200 630.450 131.400 ;
        RECT 634.950 130.800 637.050 132.900 ;
        RECT 644.400 124.050 645.450 163.950 ;
        RECT 656.400 142.050 657.450 169.950 ;
        RECT 659.400 169.050 660.450 208.950 ;
        RECT 664.950 208.800 667.050 210.900 ;
        RECT 667.950 199.950 670.050 202.050 ;
        RECT 668.400 183.600 669.450 199.950 ;
        RECT 674.400 199.050 675.450 235.950 ;
        RECT 683.400 232.050 684.450 280.950 ;
        RECT 686.400 262.050 687.450 287.400 ;
        RECT 695.400 265.050 696.450 293.400 ;
        RECT 700.950 293.100 703.050 295.200 ;
        RECT 706.950 293.100 709.050 295.200 ;
        RECT 713.400 295.050 714.450 314.400 ;
        RECT 731.400 313.050 732.450 331.950 ;
        RECT 734.400 322.050 735.450 346.950 ;
        RECT 749.400 346.050 750.450 376.950 ;
        RECT 761.400 376.050 762.450 397.950 ;
        RECT 770.400 397.050 771.450 406.950 ;
        RECT 782.400 406.050 783.450 439.950 ;
        RECT 772.950 403.950 775.050 406.050 ;
        RECT 781.950 403.950 784.050 406.050 ;
        RECT 769.950 394.950 772.050 397.050 ;
        RECT 760.950 373.950 763.050 376.050 ;
        RECT 757.950 371.100 760.050 373.200 ;
        RECT 763.950 372.000 766.050 379.050 ;
        RECT 758.400 370.350 759.600 371.100 ;
        RECT 764.400 370.350 765.600 372.000 ;
        RECT 754.950 367.950 757.050 370.050 ;
        RECT 757.950 367.950 760.050 370.050 ;
        RECT 760.950 367.950 763.050 370.050 ;
        RECT 763.950 367.950 766.050 370.050 ;
        RECT 766.950 367.950 769.050 370.050 ;
        RECT 751.950 364.950 754.050 367.050 ;
        RECT 755.400 365.400 756.600 367.650 ;
        RECT 761.400 366.900 762.600 367.650 ;
        RECT 767.400 366.900 768.600 367.650 ;
        RECT 742.950 343.950 745.050 346.050 ;
        RECT 748.950 343.950 751.050 346.050 ;
        RECT 743.400 339.600 744.450 343.950 ;
        RECT 743.400 337.350 744.600 339.600 ;
        RECT 748.950 338.100 751.050 340.200 ;
        RECT 752.400 340.050 753.450 364.950 ;
        RECT 755.400 352.050 756.450 365.400 ;
        RECT 760.950 364.800 763.050 366.900 ;
        RECT 766.950 364.800 769.050 366.900 ;
        RECT 769.950 364.950 772.050 367.050 ;
        RECT 757.950 361.950 760.050 364.050 ;
        RECT 754.950 349.950 757.050 352.050 ;
        RECT 754.950 343.950 757.050 346.050 ;
        RECT 749.400 337.350 750.600 338.100 ;
        RECT 751.950 337.950 754.050 340.050 ;
        RECT 739.950 334.950 742.050 337.050 ;
        RECT 742.950 334.950 745.050 337.050 ;
        RECT 745.950 334.950 748.050 337.050 ;
        RECT 748.950 334.950 751.050 337.050 ;
        RECT 736.950 331.950 739.050 334.050 ;
        RECT 740.400 332.400 741.600 334.650 ;
        RECT 746.400 333.900 747.600 334.650 ;
        RECT 733.950 319.950 736.050 322.050 ;
        RECT 737.400 315.450 738.450 331.950 ;
        RECT 740.400 319.050 741.450 332.400 ;
        RECT 745.950 331.800 748.050 333.900 ;
        RECT 751.950 331.950 754.050 334.050 ;
        RECT 739.950 316.950 742.050 319.050 ;
        RECT 737.400 314.400 741.450 315.450 ;
        RECT 730.950 310.950 733.050 313.050 ;
        RECT 731.400 307.050 732.450 310.950 ;
        RECT 715.950 304.950 718.050 307.050 ;
        RECT 721.950 304.950 724.050 307.050 ;
        RECT 730.950 304.950 733.050 307.050 ;
        RECT 701.400 292.350 702.600 293.100 ;
        RECT 707.400 292.350 708.600 293.100 ;
        RECT 712.950 292.950 715.050 295.050 ;
        RECT 700.950 289.950 703.050 292.050 ;
        RECT 703.950 289.950 706.050 292.050 ;
        RECT 706.950 289.950 709.050 292.050 ;
        RECT 709.950 289.950 712.050 292.050 ;
        RECT 704.400 287.400 705.600 289.650 ;
        RECT 710.400 287.400 711.600 289.650 ;
        RECT 704.400 283.050 705.450 287.400 ;
        RECT 703.950 280.950 706.050 283.050 ;
        RECT 710.400 280.050 711.450 287.400 ;
        RECT 716.400 283.050 717.450 304.950 ;
        RECT 718.950 298.950 721.050 301.050 ;
        RECT 719.400 295.200 720.450 298.950 ;
        RECT 718.950 293.100 721.050 295.200 ;
        RECT 722.400 294.600 723.450 304.950 ;
        RECT 722.400 292.350 723.600 294.600 ;
        RECT 727.950 293.100 730.050 295.200 ;
        RECT 728.400 292.350 729.600 293.100 ;
        RECT 721.950 289.950 724.050 292.050 ;
        RECT 724.950 289.950 727.050 292.050 ;
        RECT 727.950 289.950 730.050 292.050 ;
        RECT 730.950 289.950 733.050 292.050 ;
        RECT 718.950 286.950 721.050 289.050 ;
        RECT 725.400 288.900 726.600 289.650 ;
        RECT 731.400 288.900 732.600 289.650 ;
        RECT 715.950 280.950 718.050 283.050 ;
        RECT 709.950 277.950 712.050 280.050 ;
        RECT 712.950 265.950 715.050 268.050 ;
        RECT 694.950 262.950 697.050 265.050 ;
        RECT 700.950 262.950 703.050 265.050 ;
        RECT 685.950 259.950 688.050 262.050 ;
        RECT 691.950 260.100 694.050 262.200 ;
        RECT 692.400 259.350 693.600 260.100 ;
        RECT 688.950 256.950 691.050 259.050 ;
        RECT 691.950 256.950 694.050 259.050 ;
        RECT 694.950 256.950 697.050 259.050 ;
        RECT 685.950 253.950 688.050 256.050 ;
        RECT 689.400 254.400 690.600 256.650 ;
        RECT 686.400 247.050 687.450 253.950 ;
        RECT 685.950 244.950 688.050 247.050 ;
        RECT 689.400 238.050 690.450 254.400 ;
        RECT 688.950 235.950 691.050 238.050 ;
        RECT 682.950 229.950 685.050 232.050 ;
        RECT 697.950 231.450 700.050 232.050 ;
        RECT 692.400 231.000 700.050 231.450 ;
        RECT 691.950 230.400 700.050 231.000 ;
        RECT 691.950 226.950 694.050 230.400 ;
        RECT 697.950 229.950 700.050 230.400 ;
        RECT 701.400 223.050 702.450 262.950 ;
        RECT 706.950 259.950 709.050 262.050 ;
        RECT 713.400 261.600 714.450 265.950 ;
        RECT 707.400 259.350 708.600 259.950 ;
        RECT 713.400 259.350 714.600 261.600 ;
        RECT 706.950 256.950 709.050 259.050 ;
        RECT 709.950 256.950 712.050 259.050 ;
        RECT 712.950 256.950 715.050 259.050 ;
        RECT 710.400 254.400 711.600 256.650 ;
        RECT 719.400 255.450 720.450 286.950 ;
        RECT 724.950 286.800 727.050 288.900 ;
        RECT 730.950 286.800 733.050 288.900 ;
        RECT 725.400 285.450 726.450 286.800 ;
        RECT 722.400 284.400 726.450 285.450 ;
        RECT 722.400 262.050 723.450 284.400 ;
        RECT 740.400 283.050 741.450 314.400 ;
        RECT 742.950 304.950 745.050 307.050 ;
        RECT 743.400 295.050 744.450 304.950 ;
        RECT 742.950 292.950 745.050 295.050 ;
        RECT 748.950 293.100 751.050 295.200 ;
        RECT 752.400 295.050 753.450 331.950 ;
        RECT 749.400 292.350 750.600 293.100 ;
        RECT 751.950 292.950 754.050 295.050 ;
        RECT 745.950 289.950 748.050 292.050 ;
        RECT 748.950 289.950 751.050 292.050 ;
        RECT 746.400 288.900 747.600 289.650 ;
        RECT 745.950 286.800 748.050 288.900 ;
        RECT 739.950 280.950 742.050 283.050 ;
        RECT 745.950 279.450 748.050 283.050 ;
        RECT 745.950 279.000 750.450 279.450 ;
        RECT 746.400 278.400 750.450 279.000 ;
        RECT 730.950 274.950 733.050 277.050 ;
        RECT 724.950 268.950 727.050 271.050 ;
        RECT 721.950 259.950 724.050 262.050 ;
        RECT 725.400 261.600 726.450 268.950 ;
        RECT 731.400 261.600 732.450 274.950 ;
        RECT 742.950 271.950 745.050 274.050 ;
        RECT 739.950 262.950 742.050 265.050 ;
        RECT 725.400 259.350 726.600 261.600 ;
        RECT 731.400 259.350 732.600 261.600 ;
        RECT 724.950 256.950 727.050 259.050 ;
        RECT 727.950 256.950 730.050 259.050 ;
        RECT 730.950 256.950 733.050 259.050 ;
        RECT 733.950 256.950 736.050 259.050 ;
        RECT 716.400 254.400 720.450 255.450 ;
        RECT 728.400 255.000 729.600 256.650 ;
        RECT 710.400 253.050 711.450 254.400 ;
        RECT 703.950 250.950 706.050 253.050 ;
        RECT 710.400 251.400 715.050 253.050 ;
        RECT 711.000 250.950 715.050 251.400 ;
        RECT 694.950 220.950 697.050 223.050 ;
        RECT 700.950 220.950 703.050 223.050 ;
        RECT 691.950 217.950 694.050 220.050 ;
        RECT 676.950 216.600 681.000 217.050 ;
        RECT 676.950 214.950 681.600 216.600 ;
        RECT 685.950 215.100 688.050 217.200 ;
        RECT 680.400 214.350 681.600 214.950 ;
        RECT 686.400 214.350 687.600 215.100 ;
        RECT 679.950 211.950 682.050 214.050 ;
        RECT 682.950 211.950 685.050 214.050 ;
        RECT 685.950 211.950 688.050 214.050 ;
        RECT 683.400 209.400 684.600 211.650 ;
        RECT 683.400 202.050 684.450 209.400 ;
        RECT 688.950 208.950 691.050 211.050 ;
        RECT 689.400 205.050 690.450 208.950 ;
        RECT 688.950 202.950 691.050 205.050 ;
        RECT 682.950 199.950 685.050 202.050 ;
        RECT 673.950 196.950 676.050 199.050 ;
        RECT 679.950 196.950 682.050 199.050 ;
        RECT 668.400 181.350 669.600 183.600 ;
        RECT 673.950 183.000 676.050 187.050 ;
        RECT 680.400 183.450 681.450 196.950 ;
        RECT 689.400 190.050 690.450 202.950 ;
        RECT 692.400 193.050 693.450 217.950 ;
        RECT 695.400 217.050 696.450 220.950 ;
        RECT 704.400 219.450 705.450 250.950 ;
        RECT 709.950 235.950 712.050 238.050 ;
        RECT 710.400 226.050 711.450 235.950 ;
        RECT 709.950 223.950 712.050 226.050 ;
        RECT 701.400 218.400 705.450 219.450 ;
        RECT 694.950 214.950 697.050 217.050 ;
        RECT 701.400 216.600 702.450 218.400 ;
        RECT 701.400 214.350 702.600 216.600 ;
        RECT 706.950 216.000 709.050 220.050 ;
        RECT 710.400 217.050 711.450 223.950 ;
        RECT 712.950 220.950 715.050 223.050 ;
        RECT 707.400 214.350 708.600 216.000 ;
        RECT 709.950 214.950 712.050 217.050 ;
        RECT 697.950 211.950 700.050 214.050 ;
        RECT 700.950 211.950 703.050 214.050 ;
        RECT 703.950 211.950 706.050 214.050 ;
        RECT 706.950 211.950 709.050 214.050 ;
        RECT 694.950 208.950 697.050 211.050 ;
        RECT 698.400 209.400 699.600 211.650 ;
        RECT 704.400 209.400 705.600 211.650 ;
        RECT 691.950 190.950 694.050 193.050 ;
        RECT 695.400 190.050 696.450 208.950 ;
        RECT 698.400 202.050 699.450 209.400 ;
        RECT 697.950 199.950 700.050 202.050 ;
        RECT 688.950 187.950 691.050 190.050 ;
        RECT 694.950 187.950 697.050 190.050 ;
        RECT 700.950 187.950 703.050 190.050 ;
        RECT 674.400 181.350 675.600 183.000 ;
        RECT 680.400 182.400 684.450 183.450 ;
        RECT 664.950 178.950 667.050 181.050 ;
        RECT 667.950 178.950 670.050 181.050 ;
        RECT 670.950 178.950 673.050 181.050 ;
        RECT 673.950 178.950 676.050 181.050 ;
        RECT 676.950 178.950 679.050 181.050 ;
        RECT 665.400 177.900 666.600 178.650 ;
        RECT 664.950 175.800 667.050 177.900 ;
        RECT 671.400 176.400 672.600 178.650 ;
        RECT 677.400 176.400 678.600 178.650 ;
        RECT 683.400 177.900 684.450 182.400 ;
        RECT 688.950 182.100 691.050 184.200 ;
        RECT 694.950 182.100 697.050 184.200 ;
        RECT 701.400 184.050 702.450 187.950 ;
        RECT 689.400 181.350 690.600 182.100 ;
        RECT 695.400 181.350 696.600 182.100 ;
        RECT 700.950 181.950 703.050 184.050 ;
        RECT 688.950 178.950 691.050 181.050 ;
        RECT 691.950 178.950 694.050 181.050 ;
        RECT 694.950 178.950 697.050 181.050 ;
        RECT 697.950 178.950 700.050 181.050 ;
        RECT 658.950 166.950 661.050 169.050 ;
        RECT 659.400 151.050 660.450 166.950 ;
        RECT 671.400 166.050 672.450 176.400 ;
        RECT 677.400 169.050 678.450 176.400 ;
        RECT 682.800 175.800 684.900 177.900 ;
        RECT 685.950 175.950 688.050 178.050 ;
        RECT 692.400 176.400 693.600 178.650 ;
        RECT 698.400 176.400 699.600 178.650 ;
        RECT 683.400 169.050 684.450 175.800 ;
        RECT 676.950 166.950 679.050 169.050 ;
        RECT 682.950 166.950 685.050 169.050 ;
        RECT 670.950 163.950 673.050 166.050 ;
        RECT 686.400 160.050 687.450 175.950 ;
        RECT 692.400 166.050 693.450 176.400 ;
        RECT 698.400 172.050 699.450 176.400 ;
        RECT 700.950 175.950 703.050 178.050 ;
        RECT 697.950 169.950 700.050 172.050 ;
        RECT 691.950 163.950 694.050 166.050 ;
        RECT 670.950 157.950 673.050 160.050 ;
        RECT 685.950 157.950 688.050 160.050 ;
        RECT 671.400 154.050 672.450 157.950 ;
        RECT 692.400 154.050 693.450 163.950 ;
        RECT 670.950 151.950 673.050 154.050 ;
        RECT 685.950 151.950 688.050 154.050 ;
        RECT 691.950 151.950 694.050 154.050 ;
        RECT 658.950 148.950 661.050 151.050 ;
        RECT 649.950 137.100 652.050 142.050 ;
        RECT 655.950 139.950 658.050 142.050 ;
        RECT 656.400 138.600 657.450 139.950 ;
        RECT 671.400 138.600 672.450 151.950 ;
        RECT 676.950 148.950 679.050 151.050 ;
        RECT 677.400 138.600 678.450 148.950 ;
        RECT 650.400 136.350 651.600 137.100 ;
        RECT 656.400 136.350 657.600 138.600 ;
        RECT 671.400 136.350 672.600 138.600 ;
        RECT 677.400 136.350 678.600 138.600 ;
        RECT 649.950 133.950 652.050 136.050 ;
        RECT 652.950 133.950 655.050 136.050 ;
        RECT 655.950 133.950 658.050 136.050 ;
        RECT 658.950 133.950 661.050 136.050 ;
        RECT 670.950 133.950 673.050 136.050 ;
        RECT 673.950 133.950 676.050 136.050 ;
        RECT 676.950 133.950 679.050 136.050 ;
        RECT 679.950 133.950 682.050 136.050 ;
        RECT 653.400 132.900 654.600 133.650 ;
        RECT 652.950 130.800 655.050 132.900 ;
        RECT 659.400 131.400 660.600 133.650 ;
        RECT 674.400 132.000 675.600 133.650 ;
        RECT 680.400 132.900 681.600 133.650 ;
        RECT 686.400 132.900 687.450 151.950 ;
        RECT 701.400 142.050 702.450 175.950 ;
        RECT 704.400 145.050 705.450 209.400 ;
        RECT 709.950 208.950 712.050 211.050 ;
        RECT 710.400 187.050 711.450 208.950 ;
        RECT 713.400 187.200 714.450 220.950 ;
        RECT 709.950 184.950 712.050 187.050 ;
        RECT 712.950 185.100 715.050 187.200 ;
        RECT 716.400 184.050 717.450 254.400 ;
        RECT 727.950 250.950 730.050 255.000 ;
        RECT 734.400 254.400 735.600 256.650 ;
        RECT 734.400 247.050 735.450 254.400 ;
        RECT 736.950 253.950 739.050 256.050 ;
        RECT 733.950 244.950 736.050 247.050 ;
        RECT 721.800 220.500 723.900 222.600 ;
        RECT 719.100 211.950 721.200 214.050 ;
        RECT 722.100 213.300 723.300 220.500 ;
        RECT 725.400 217.350 726.600 219.600 ;
        RECT 731.400 219.300 733.500 221.400 ;
        RECT 725.100 214.950 727.200 217.050 ;
        RECT 728.100 215.700 730.200 217.800 ;
        RECT 728.100 213.300 729.000 215.700 ;
        RECT 722.100 212.100 729.000 213.300 ;
        RECT 719.400 210.900 720.600 211.650 ;
        RECT 718.950 208.800 721.050 210.900 ;
        RECT 722.100 206.700 723.000 212.100 ;
        RECT 723.900 210.300 726.000 211.200 ;
        RECT 731.700 210.300 732.600 219.300 ;
        RECT 733.950 215.100 736.050 217.200 ;
        RECT 734.400 214.350 735.600 215.100 ;
        RECT 733.800 211.950 735.900 214.050 ;
        RECT 723.900 209.100 732.600 210.300 ;
        RECT 721.800 204.600 723.900 206.700 ;
        RECT 725.100 206.100 727.200 208.200 ;
        RECT 729.000 207.300 731.100 209.100 ;
        RECT 737.400 207.450 738.450 253.950 ;
        RECT 734.400 206.400 738.450 207.450 ;
        RECT 725.400 204.000 726.600 205.800 ;
        RECT 721.800 199.950 723.900 202.050 ;
        RECT 724.950 199.950 727.050 204.000 ;
        RECT 718.950 184.950 721.050 187.050 ;
        RECT 712.800 181.950 714.900 184.050 ;
        RECT 715.950 181.950 718.050 184.050 ;
        RECT 713.400 181.350 714.600 181.950 ;
        RECT 709.950 178.950 712.050 181.050 ;
        RECT 712.950 178.950 715.050 181.050 ;
        RECT 706.950 175.950 709.050 178.050 ;
        RECT 710.400 176.400 711.600 178.650 ;
        RECT 707.400 172.050 708.450 175.950 ;
        RECT 706.950 169.950 709.050 172.050 ;
        RECT 710.400 166.050 711.450 176.400 ;
        RECT 719.400 166.050 720.450 184.950 ;
        RECT 722.400 184.050 723.450 199.950 ;
        RECT 727.950 187.950 730.050 190.050 ;
        RECT 721.950 181.950 724.050 184.050 ;
        RECT 728.400 183.600 729.450 187.950 ;
        RECT 734.400 184.050 735.450 206.400 ;
        RECT 740.400 186.450 741.450 262.950 ;
        RECT 743.400 232.050 744.450 271.950 ;
        RECT 749.400 261.600 750.450 278.400 ;
        RECT 755.400 265.200 756.450 343.950 ;
        RECT 758.400 333.900 759.450 361.950 ;
        RECT 770.400 361.050 771.450 364.950 ;
        RECT 769.950 358.950 772.050 361.050 ;
        RECT 773.400 352.050 774.450 403.950 ;
        RECT 785.400 378.450 786.450 443.400 ;
        RECT 794.400 427.050 795.450 443.400 ;
        RECT 799.950 439.950 802.050 444.000 ;
        RECT 809.400 442.050 810.450 487.800 ;
        RECT 812.400 484.050 813.450 518.400 ;
        RECT 820.950 514.950 823.050 517.050 ;
        RECT 821.400 495.600 822.450 514.950 ;
        RECT 824.400 505.050 825.450 520.800 ;
        RECT 823.950 502.950 826.050 505.050 ;
        RECT 821.400 493.350 822.600 495.600 ;
        RECT 817.950 490.950 820.050 493.050 ;
        RECT 820.950 490.950 823.050 493.050 ;
        RECT 823.950 490.950 826.050 493.050 ;
        RECT 818.400 488.400 819.600 490.650 ;
        RECT 824.400 488.400 825.600 490.650 ;
        RECT 818.400 487.050 819.450 488.400 ;
        RECT 811.950 481.950 814.050 484.050 ;
        RECT 817.950 481.950 820.050 487.050 ;
        RECT 824.400 454.050 825.450 488.400 ;
        RECT 830.400 454.050 831.450 529.950 ;
        RECT 833.400 529.050 834.450 532.950 ;
        RECT 832.950 526.950 835.050 529.050 ;
        RECT 839.400 528.600 840.450 535.950 ;
        RECT 841.950 532.950 847.050 535.050 ;
        RECT 839.400 526.350 840.600 528.600 ;
        RECT 844.950 528.000 847.050 531.900 ;
        RECT 848.400 528.450 849.450 595.950 ;
        RECT 851.400 589.050 852.450 598.950 ;
        RECT 850.950 586.950 853.050 589.050 ;
        RECT 854.400 577.050 855.450 653.400 ;
        RECT 860.400 651.450 861.450 734.400 ;
        RECT 865.950 733.950 868.050 736.050 ;
        RECT 866.400 729.600 867.450 733.950 ;
        RECT 866.400 727.350 867.600 729.600 ;
        RECT 865.950 724.950 868.050 727.050 ;
        RECT 868.950 724.950 871.050 727.050 ;
        RECT 869.400 723.900 870.600 724.650 ;
        RECT 868.950 721.800 871.050 723.900 ;
        RECT 869.400 667.050 870.450 721.800 ;
        RECT 868.950 664.950 871.050 667.050 ;
        RECT 862.950 655.950 865.050 658.050 ;
        RECT 857.400 650.400 861.450 651.450 ;
        RECT 863.400 651.600 864.450 655.950 ;
        RECT 857.400 583.050 858.450 650.400 ;
        RECT 863.400 649.350 864.600 651.600 ;
        RECT 868.950 650.100 871.050 652.200 ;
        RECT 875.400 652.050 876.450 736.950 ;
        RECT 869.400 649.350 870.600 650.100 ;
        RECT 874.950 649.950 877.050 652.050 ;
        RECT 862.950 646.950 865.050 649.050 ;
        RECT 865.950 646.950 868.050 649.050 ;
        RECT 868.950 646.950 871.050 649.050 ;
        RECT 871.950 646.950 874.050 649.050 ;
        RECT 859.950 643.950 862.050 646.050 ;
        RECT 866.400 644.400 867.600 646.650 ;
        RECT 872.400 645.000 873.600 646.650 ;
        RECT 860.400 640.050 861.450 643.950 ;
        RECT 866.400 642.450 867.450 644.400 ;
        RECT 866.400 641.400 870.450 642.450 ;
        RECT 859.950 637.950 862.050 640.050 ;
        RECT 865.950 637.950 868.050 640.050 ;
        RECT 859.950 634.800 862.050 636.900 ;
        RECT 860.400 607.050 861.450 634.800 ;
        RECT 862.950 613.950 865.050 616.050 ;
        RECT 863.400 610.050 864.450 613.950 ;
        RECT 862.950 607.950 865.050 610.050 ;
        RECT 859.950 604.950 862.050 607.050 ;
        RECT 866.400 606.600 867.450 637.950 ;
        RECT 869.400 627.450 870.450 641.400 ;
        RECT 871.950 640.950 874.050 645.000 ;
        RECT 874.950 643.950 877.050 646.050 ;
        RECT 869.400 626.400 873.450 627.450 ;
        RECT 866.400 604.350 867.600 606.600 ;
        RECT 862.950 601.950 865.050 604.050 ;
        RECT 865.950 601.950 868.050 604.050 ;
        RECT 859.950 598.950 862.050 601.050 ;
        RECT 863.400 600.000 864.600 601.650 ;
        RECT 860.400 594.450 861.450 598.950 ;
        RECT 862.950 595.950 865.050 600.000 ;
        RECT 868.950 598.950 871.050 601.050 ;
        RECT 860.400 593.400 864.450 594.450 ;
        RECT 856.950 580.950 859.050 583.050 ;
        RECT 853.950 574.950 856.050 577.050 ;
        RECT 856.950 572.100 859.050 574.200 ;
        RECT 863.400 573.600 864.450 593.400 ;
        RECT 865.950 580.950 868.050 583.050 ;
        RECT 866.400 574.050 867.450 580.950 ;
        RECT 857.400 571.350 858.600 572.100 ;
        RECT 863.400 571.350 864.600 573.600 ;
        RECT 865.950 571.950 868.050 574.050 ;
        RECT 853.950 568.950 856.050 571.050 ;
        RECT 856.950 568.950 859.050 571.050 ;
        RECT 859.950 568.950 862.050 571.050 ;
        RECT 862.950 568.950 865.050 571.050 ;
        RECT 850.950 565.950 853.050 568.050 ;
        RECT 854.400 566.400 855.600 568.650 ;
        RECT 860.400 567.900 861.600 568.650 ;
        RECT 851.400 532.050 852.450 565.950 ;
        RECT 854.400 550.050 855.450 566.400 ;
        RECT 859.950 565.800 862.050 567.900 ;
        RECT 865.950 565.950 868.050 568.050 ;
        RECT 869.400 567.900 870.450 598.950 ;
        RECT 853.950 547.950 856.050 550.050 ;
        RECT 856.950 532.950 859.050 535.050 ;
        RECT 850.950 529.950 853.050 532.050 ;
        RECT 850.950 528.450 853.050 528.900 ;
        RECT 845.400 526.350 846.600 528.000 ;
        RECT 848.400 527.400 853.050 528.450 ;
        RECT 850.950 526.800 853.050 527.400 ;
        RECT 857.400 528.600 858.450 532.950 ;
        RECT 835.950 523.950 838.050 526.050 ;
        RECT 838.950 523.950 841.050 526.050 ;
        RECT 841.950 523.950 844.050 526.050 ;
        RECT 844.950 523.950 847.050 526.050 ;
        RECT 836.400 521.400 837.600 523.650 ;
        RECT 842.400 522.900 843.600 523.650 ;
        RECT 836.400 517.050 837.450 521.400 ;
        RECT 841.950 520.800 844.050 522.900 ;
        RECT 851.400 522.450 852.450 526.800 ;
        RECT 857.400 526.350 858.600 528.600 ;
        RECT 862.950 527.100 865.050 529.200 ;
        RECT 866.400 529.050 867.450 565.950 ;
        RECT 868.950 565.800 871.050 567.900 ;
        RECT 868.950 559.950 871.050 562.050 ;
        RECT 863.400 526.350 864.600 527.100 ;
        RECT 865.950 526.950 868.050 529.050 ;
        RECT 856.950 523.950 859.050 526.050 ;
        RECT 859.950 523.950 862.050 526.050 ;
        RECT 862.950 523.950 865.050 526.050 ;
        RECT 848.400 521.400 852.450 522.450 ;
        RECT 835.950 514.950 838.050 517.050 ;
        RECT 848.400 511.050 849.450 521.400 ;
        RECT 853.950 520.950 856.050 523.050 ;
        RECT 860.400 522.900 861.600 523.650 ;
        RECT 869.400 523.050 870.450 559.950 ;
        RECT 872.400 547.050 873.450 626.400 ;
        RECT 871.950 544.950 874.050 547.050 ;
        RECT 871.950 526.950 874.050 529.050 ;
        RECT 847.950 508.950 850.050 511.050 ;
        RECT 848.400 501.450 849.450 508.950 ;
        RECT 854.400 505.050 855.450 520.950 ;
        RECT 859.950 520.800 862.050 522.900 ;
        RECT 868.950 520.950 871.050 523.050 ;
        RECT 853.950 502.950 856.050 505.050 ;
        RECT 859.950 502.950 862.050 505.050 ;
        RECT 848.400 499.200 849.600 501.450 ;
        RECT 832.950 494.100 835.050 496.200 ;
        RECT 843.900 495.900 846.000 497.700 ;
        RECT 847.800 496.800 849.900 498.900 ;
        RECT 851.100 498.300 853.200 500.400 ;
        RECT 842.400 494.700 851.100 495.900 ;
        RECT 823.950 451.950 826.050 454.050 ;
        RECT 829.950 451.950 832.050 454.050 ;
        RECT 811.950 448.950 814.050 451.050 ;
        RECT 820.950 449.100 823.050 451.200 ;
        RECT 808.950 439.950 811.050 442.050 ;
        RECT 812.400 433.050 813.450 448.950 ;
        RECT 821.400 448.350 822.600 449.100 ;
        RECT 817.950 445.950 820.050 448.050 ;
        RECT 820.950 445.950 823.050 448.050 ;
        RECT 823.950 445.950 826.050 448.050 ;
        RECT 818.400 443.400 819.600 445.650 ;
        RECT 824.400 444.900 825.600 445.650 ;
        RECT 818.400 442.050 819.450 443.400 ;
        RECT 823.950 442.800 826.050 444.900 ;
        RECT 817.950 439.950 820.050 442.050 ;
        RECT 799.950 430.950 802.050 433.050 ;
        RECT 811.950 430.950 814.050 433.050 ;
        RECT 793.950 424.950 796.050 427.050 ;
        RECT 793.950 417.000 796.050 421.050 ;
        RECT 794.400 415.350 795.600 417.000 ;
        RECT 788.100 412.950 790.200 415.050 ;
        RECT 793.500 412.950 795.600 415.050 ;
        RECT 796.800 412.950 798.900 415.050 ;
        RECT 788.400 411.900 789.600 412.650 ;
        RECT 787.950 409.800 790.050 411.900 ;
        RECT 797.400 410.400 798.600 412.650 ;
        RECT 797.400 406.050 798.450 410.400 ;
        RECT 796.950 403.950 799.050 406.050 ;
        RECT 800.400 397.050 801.450 430.950 ;
        RECT 818.400 427.050 819.450 439.950 ;
        RECT 824.400 436.050 825.450 442.800 ;
        RECT 830.400 442.050 831.450 451.950 ;
        RECT 829.950 439.950 832.050 442.050 ;
        RECT 833.400 436.050 834.450 494.100 ;
        RECT 839.100 490.950 841.200 493.050 ;
        RECT 839.400 489.900 840.600 490.650 ;
        RECT 838.950 487.800 841.050 489.900 ;
        RECT 842.400 485.700 843.300 494.700 ;
        RECT 849.000 493.800 851.100 494.700 ;
        RECT 852.000 492.900 852.900 498.300 ;
        RECT 853.950 494.100 856.050 496.200 ;
        RECT 854.400 493.350 855.600 494.100 ;
        RECT 846.000 491.700 852.900 492.900 ;
        RECT 846.000 489.300 846.900 491.700 ;
        RECT 844.800 487.200 846.900 489.300 ;
        RECT 847.800 487.950 849.900 490.050 ;
        RECT 835.950 481.950 838.050 484.050 ;
        RECT 841.500 483.600 843.600 485.700 ;
        RECT 848.400 485.400 849.600 487.650 ;
        RECT 851.700 484.500 852.900 491.700 ;
        RECT 853.800 490.950 855.900 493.050 ;
        RECT 851.100 482.400 853.200 484.500 ;
        RECT 836.400 450.600 837.450 481.950 ;
        RECT 853.950 460.950 856.050 463.050 ;
        RECT 844.950 454.950 847.050 457.050 ;
        RECT 845.400 450.600 846.450 454.950 ;
        RECT 836.400 448.350 837.600 450.600 ;
        RECT 845.400 448.350 846.600 450.600 ;
        RECT 847.950 448.950 850.050 451.050 ;
        RECT 836.100 445.950 838.200 448.050 ;
        RECT 841.500 445.950 843.600 448.050 ;
        RECT 844.800 445.950 846.900 448.050 ;
        RECT 842.400 444.900 843.600 445.650 ;
        RECT 848.400 444.900 849.450 448.950 ;
        RECT 841.950 442.800 844.050 444.900 ;
        RECT 847.950 442.800 850.050 444.900 ;
        RECT 823.950 433.950 826.050 436.050 ;
        RECT 832.950 433.950 835.050 436.050 ;
        RECT 850.950 433.950 853.050 436.050 ;
        RECT 820.950 430.950 823.050 433.050 ;
        RECT 817.950 424.950 820.050 427.050 ;
        RECT 811.950 421.950 814.050 424.050 ;
        RECT 812.400 417.600 813.450 421.950 ;
        RECT 812.400 415.350 813.600 417.600 ;
        RECT 808.950 412.950 811.050 415.050 ;
        RECT 811.950 412.950 814.050 415.050 ;
        RECT 814.950 412.950 817.050 415.050 ;
        RECT 809.400 411.900 810.600 412.650 ;
        RECT 808.950 409.800 811.050 411.900 ;
        RECT 815.400 410.400 816.600 412.650 ;
        RECT 809.400 400.050 810.450 409.800 ;
        RECT 815.400 406.050 816.450 410.400 ;
        RECT 814.950 403.950 817.050 406.050 ;
        RECT 808.950 397.950 811.050 400.050 ;
        RECT 799.950 394.950 802.050 397.050 ;
        RECT 817.950 394.950 820.050 397.050 ;
        RECT 785.400 377.400 789.450 378.450 ;
        RECT 781.950 371.100 784.050 373.200 ;
        RECT 782.400 370.350 783.600 371.100 ;
        RECT 778.950 367.950 781.050 370.050 ;
        RECT 781.950 367.950 784.050 370.050 ;
        RECT 779.400 366.900 780.600 367.650 ;
        RECT 778.950 364.800 781.050 366.900 ;
        RECT 779.400 358.050 780.450 364.800 ;
        RECT 788.400 364.050 789.450 377.400 ;
        RECT 790.800 376.950 792.900 379.050 ;
        RECT 791.400 373.200 792.450 376.950 ;
        RECT 799.500 375.300 801.600 377.400 ;
        RECT 809.100 376.500 811.200 378.600 ;
        RECT 790.950 371.100 793.050 373.200 ;
        RECT 796.950 371.100 799.050 373.200 ;
        RECT 797.400 370.350 798.600 371.100 ;
        RECT 797.100 367.950 799.200 370.050 ;
        RECT 800.400 366.300 801.300 375.300 ;
        RECT 802.800 371.700 804.900 373.800 ;
        RECT 806.400 373.350 807.600 375.600 ;
        RECT 804.000 369.300 804.900 371.700 ;
        RECT 805.800 370.950 807.900 373.050 ;
        RECT 809.700 369.300 810.900 376.500 ;
        RECT 814.950 370.950 817.050 373.050 ;
        RECT 804.000 368.100 810.900 369.300 ;
        RECT 807.000 366.300 809.100 367.200 ;
        RECT 800.400 365.100 809.100 366.300 ;
        RECT 787.950 361.950 790.050 364.050 ;
        RECT 793.950 361.800 796.050 363.900 ;
        RECT 801.900 363.300 804.000 365.100 ;
        RECT 805.800 362.100 807.900 364.200 ;
        RECT 810.000 362.700 810.900 368.100 ;
        RECT 811.800 367.950 813.900 370.050 ;
        RECT 812.400 366.900 813.600 367.650 ;
        RECT 811.950 364.800 814.050 366.900 ;
        RECT 778.950 355.950 781.050 358.050 ;
        RECT 787.950 355.950 790.050 358.050 ;
        RECT 772.950 349.950 775.050 352.050 ;
        RECT 778.950 349.950 781.050 352.050 ;
        RECT 766.950 343.950 769.050 346.050 ;
        RECT 767.400 339.600 768.450 343.950 ;
        RECT 767.400 337.350 768.600 339.600 ;
        RECT 772.950 338.100 775.050 340.200 ;
        RECT 773.400 337.350 774.600 338.100 ;
        RECT 763.950 334.950 766.050 337.050 ;
        RECT 766.950 334.950 769.050 337.050 ;
        RECT 769.950 334.950 772.050 337.050 ;
        RECT 772.950 334.950 775.050 337.050 ;
        RECT 757.950 331.800 760.050 333.900 ;
        RECT 764.400 332.400 765.600 334.650 ;
        RECT 770.400 333.900 771.600 334.650 ;
        RECT 760.950 322.950 763.050 325.050 ;
        RECT 761.400 304.050 762.450 322.950 ;
        RECT 764.400 313.050 765.450 332.400 ;
        RECT 769.950 331.800 772.050 333.900 ;
        RECT 779.400 333.450 780.450 349.950 ;
        RECT 788.400 346.050 789.450 355.950 ;
        RECT 787.950 343.950 790.050 346.050 ;
        RECT 787.950 338.100 790.050 340.200 ;
        RECT 794.400 340.050 795.450 361.800 ;
        RECT 806.400 359.550 807.600 361.800 ;
        RECT 809.100 360.600 811.200 362.700 ;
        RECT 815.400 361.050 816.450 370.950 ;
        RECT 818.400 366.450 819.450 394.950 ;
        RECT 821.400 373.050 822.450 430.950 ;
        RECT 832.950 423.000 835.050 427.050 ;
        RECT 851.400 423.450 852.450 433.950 ;
        RECT 854.400 427.050 855.450 460.950 ;
        RECT 860.400 451.200 861.450 502.950 ;
        RECT 872.400 463.050 873.450 526.950 ;
        RECT 871.950 460.950 874.050 463.050 ;
        RECT 865.950 454.950 868.050 457.050 ;
        RECT 866.400 451.200 867.450 454.950 ;
        RECT 859.950 449.100 862.050 451.200 ;
        RECT 865.950 449.100 868.050 451.200 ;
        RECT 871.950 449.100 874.050 451.200 ;
        RECT 860.400 448.350 861.600 449.100 ;
        RECT 866.400 448.350 867.600 449.100 ;
        RECT 859.950 445.950 862.050 448.050 ;
        RECT 862.950 445.950 865.050 448.050 ;
        RECT 865.950 445.950 868.050 448.050 ;
        RECT 863.400 444.000 864.600 445.650 ;
        RECT 862.950 439.950 865.050 444.000 ;
        RECT 853.950 424.950 856.050 427.050 ;
        RECT 868.950 424.950 871.050 427.050 ;
        RECT 833.400 421.200 834.600 423.000 ;
        RECT 851.400 422.400 855.450 423.450 ;
        RECT 829.500 419.100 831.600 421.200 ;
        RECT 827.400 417.450 828.600 417.600 ;
        RECT 824.400 416.400 828.600 417.450 ;
        RECT 824.400 412.050 825.450 416.400 ;
        RECT 827.400 415.350 828.600 416.400 ;
        RECT 827.100 412.950 829.200 415.050 ;
        RECT 830.100 414.000 831.000 419.100 ;
        RECT 832.800 418.800 834.900 420.900 ;
        RECT 839.400 419.400 841.500 421.500 ;
        RECT 837.000 417.000 839.100 417.900 ;
        RECT 831.900 415.800 839.100 417.000 ;
        RECT 831.900 414.900 834.000 415.800 ;
        RECT 837.000 414.000 839.100 414.900 ;
        RECT 830.100 413.100 839.100 414.000 ;
        RECT 823.950 409.950 826.050 412.050 ;
        RECT 826.950 406.950 829.050 409.050 ;
        RECT 827.400 376.050 828.450 406.950 ;
        RECT 830.100 406.500 831.000 413.100 ;
        RECT 837.000 412.800 839.100 413.100 ;
        RECT 832.800 409.950 834.900 412.050 ;
        RECT 833.400 407.400 834.600 409.650 ;
        RECT 840.000 406.800 840.900 419.400 ;
        RECT 847.950 416.100 850.050 418.200 ;
        RECT 854.400 417.600 855.450 422.400 ;
        RECT 841.800 412.950 843.900 415.050 ;
        RECT 842.400 411.450 843.600 412.650 ;
        RECT 842.400 410.400 846.450 411.450 ;
        RECT 830.100 404.400 832.200 406.500 ;
        RECT 839.100 404.700 841.200 406.800 ;
        RECT 845.400 406.050 846.450 410.400 ;
        RECT 844.950 403.950 847.050 406.050 ;
        RECT 848.400 403.050 849.450 416.100 ;
        RECT 854.400 415.350 855.600 417.600 ;
        RECT 859.950 416.100 862.050 418.200 ;
        RECT 860.400 415.350 861.600 416.100 ;
        RECT 853.950 412.950 856.050 415.050 ;
        RECT 856.950 412.950 859.050 415.050 ;
        RECT 859.950 412.950 862.050 415.050 ;
        RECT 862.950 412.950 865.050 415.050 ;
        RECT 857.400 410.400 858.600 412.650 ;
        RECT 863.400 411.000 864.600 412.650 ;
        RECT 857.400 408.450 858.450 410.400 ;
        RECT 854.400 407.400 858.450 408.450 ;
        RECT 832.950 400.950 835.050 403.050 ;
        RECT 847.950 400.950 850.050 403.050 ;
        RECT 833.400 382.050 834.450 400.950 ;
        RECT 832.950 379.950 835.050 382.050 ;
        RECT 826.950 373.950 829.050 376.050 ;
        RECT 829.950 373.050 832.050 373.200 ;
        RECT 820.950 370.950 823.050 373.050 ;
        RECT 828.000 372.600 832.050 373.050 ;
        RECT 827.400 371.100 832.050 372.600 ;
        RECT 827.400 370.950 831.000 371.100 ;
        RECT 827.400 370.350 828.600 370.950 ;
        RECT 833.400 370.050 834.450 379.950 ;
        RECT 838.950 371.100 841.050 373.200 ;
        RECT 844.950 371.100 847.050 373.200 ;
        RECT 839.400 370.350 840.600 371.100 ;
        RECT 845.400 370.350 846.600 371.100 ;
        RECT 823.950 367.950 826.050 370.050 ;
        RECT 826.950 367.950 829.050 370.050 ;
        RECT 832.950 367.950 835.050 370.050 ;
        RECT 838.950 367.950 841.050 370.050 ;
        RECT 841.950 367.950 844.050 370.050 ;
        RECT 844.950 367.950 847.050 370.050 ;
        RECT 847.950 367.950 850.050 370.050 ;
        RECT 824.400 366.900 825.600 367.650 ;
        RECT 818.400 365.400 822.450 366.450 ;
        RECT 799.950 355.950 802.050 358.050 ;
        RECT 800.400 352.050 801.450 355.950 ;
        RECT 799.950 349.950 802.050 352.050 ;
        RECT 806.400 346.050 807.450 359.550 ;
        RECT 814.950 358.950 817.050 361.050 ;
        RECT 814.950 349.950 817.050 352.050 ;
        RECT 811.950 346.950 814.050 349.050 ;
        RECT 799.950 343.950 802.050 346.050 ;
        RECT 805.950 343.950 808.050 346.050 ;
        RECT 800.400 340.050 801.450 343.950 ;
        RECT 788.400 337.350 789.600 338.100 ;
        RECT 793.950 337.950 796.050 340.050 ;
        RECT 799.950 337.950 802.050 340.050 ;
        RECT 805.950 339.000 808.050 342.900 ;
        RECT 812.400 339.600 813.450 346.950 ;
        RECT 815.400 340.050 816.450 349.950 ;
        RECT 821.400 346.050 822.450 365.400 ;
        RECT 823.950 364.800 826.050 366.900 ;
        RECT 829.950 364.950 832.050 367.050 ;
        RECT 824.400 352.050 825.450 364.800 ;
        RECT 826.950 352.950 829.050 355.050 ;
        RECT 823.950 349.950 826.050 352.050 ;
        RECT 827.400 346.050 828.450 352.950 ;
        RECT 830.400 349.050 831.450 364.950 ;
        RECT 832.950 364.800 835.050 366.900 ;
        RECT 842.400 365.400 843.600 367.650 ;
        RECT 848.400 366.900 849.600 367.650 ;
        RECT 854.400 367.050 855.450 407.400 ;
        RECT 862.950 406.950 865.050 411.000 ;
        RECT 865.950 409.950 868.050 412.050 ;
        RECT 862.950 379.950 865.050 382.050 ;
        RECT 863.400 376.050 864.450 379.950 ;
        RECT 862.950 373.950 865.050 376.050 ;
        RECT 859.950 371.100 862.050 373.200 ;
        RECT 866.400 373.050 867.450 409.950 ;
        RECT 860.400 370.350 861.600 371.100 ;
        RECT 865.950 370.950 868.050 373.050 ;
        RECT 859.950 367.950 862.050 370.050 ;
        RECT 862.950 367.950 865.050 370.050 ;
        RECT 863.400 367.050 864.600 367.650 ;
        RECT 829.950 346.950 832.050 349.050 ;
        RECT 820.950 343.950 823.050 346.050 ;
        RECT 826.950 343.950 829.050 346.050 ;
        RECT 830.400 343.050 831.450 346.950 ;
        RECT 817.950 340.950 820.050 343.050 ;
        RECT 806.400 337.350 807.600 339.000 ;
        RECT 812.400 337.350 813.600 339.600 ;
        RECT 814.950 337.950 817.050 340.050 ;
        RECT 784.950 334.950 787.050 337.050 ;
        RECT 787.950 334.950 790.050 337.050 ;
        RECT 790.950 334.950 793.050 337.050 ;
        RECT 802.950 334.950 805.050 337.050 ;
        RECT 805.950 334.950 808.050 337.050 ;
        RECT 808.950 334.950 811.050 337.050 ;
        RECT 811.950 334.950 814.050 337.050 ;
        RECT 776.400 332.400 780.450 333.450 ;
        RECT 791.400 333.450 792.600 334.650 ;
        RECT 791.400 332.400 795.450 333.450 ;
        RECT 772.950 319.050 775.050 322.050 ;
        RECT 769.950 318.000 775.050 319.050 ;
        RECT 769.950 317.400 774.450 318.000 ;
        RECT 769.950 316.950 774.000 317.400 ;
        RECT 763.950 310.950 766.050 313.050 ;
        RECT 763.950 304.950 766.050 307.050 ;
        RECT 769.950 304.950 772.050 307.050 ;
        RECT 760.950 301.950 763.050 304.050 ;
        RECT 757.950 298.950 760.050 301.050 ;
        RECT 758.400 295.050 759.450 298.950 ;
        RECT 764.400 298.050 765.450 304.950 ;
        RECT 764.400 296.400 769.050 298.050 ;
        RECT 765.000 295.950 769.050 296.400 ;
        RECT 757.950 292.950 760.050 295.050 ;
        RECT 763.950 293.100 766.050 295.200 ;
        RECT 770.400 294.600 771.450 304.950 ;
        RECT 772.950 301.950 775.050 304.050 ;
        RECT 773.400 295.050 774.450 301.950 ;
        RECT 764.400 292.350 765.600 293.100 ;
        RECT 770.400 292.350 771.600 294.600 ;
        RECT 772.950 292.950 775.050 295.050 ;
        RECT 760.950 289.950 763.050 292.050 ;
        RECT 763.950 289.950 766.050 292.050 ;
        RECT 766.950 289.950 769.050 292.050 ;
        RECT 769.950 289.950 772.050 292.050 ;
        RECT 757.950 286.950 760.050 289.050 ;
        RECT 761.400 287.400 762.600 289.650 ;
        RECT 767.400 287.400 768.600 289.650 ;
        RECT 758.400 271.050 759.450 286.950 ;
        RECT 761.400 283.050 762.450 287.400 ;
        RECT 760.950 280.950 763.050 283.050 ;
        RECT 763.950 277.950 766.050 280.050 ;
        RECT 757.950 268.950 760.050 271.050 ;
        RECT 754.950 263.100 757.050 265.200 ;
        RECT 749.400 259.350 750.600 261.600 ;
        RECT 754.950 259.950 757.050 262.050 ;
        RECT 755.400 259.350 756.600 259.950 ;
        RECT 748.950 256.950 751.050 259.050 ;
        RECT 751.950 256.950 754.050 259.050 ;
        RECT 754.950 256.950 757.050 259.050 ;
        RECT 757.950 256.950 760.050 259.050 ;
        RECT 752.400 255.900 753.600 256.650 ;
        RECT 751.950 253.800 754.050 255.900 ;
        RECT 758.400 254.400 759.600 256.650 ;
        RECT 754.950 250.950 757.050 253.050 ;
        RECT 742.950 229.950 745.050 232.050 ;
        RECT 742.950 216.450 745.050 217.200 ;
        RECT 755.400 216.600 756.450 250.950 ;
        RECT 746.400 216.450 747.600 216.600 ;
        RECT 742.950 215.400 747.600 216.450 ;
        RECT 742.950 215.100 745.050 215.400 ;
        RECT 743.400 190.050 744.450 215.100 ;
        RECT 746.400 214.350 747.600 215.400 ;
        RECT 755.400 214.350 756.600 216.600 ;
        RECT 746.100 211.950 748.200 214.050 ;
        RECT 749.400 211.950 751.500 214.050 ;
        RECT 754.800 211.950 756.900 214.050 ;
        RECT 749.400 210.900 750.600 211.650 ;
        RECT 748.950 208.800 751.050 210.900 ;
        RECT 754.950 202.950 757.050 205.050 ;
        RECT 742.950 187.950 745.050 190.050 ;
        RECT 751.950 187.950 754.050 190.050 ;
        RECT 737.400 185.400 741.450 186.450 ;
        RECT 728.400 181.350 729.600 183.600 ;
        RECT 733.950 181.950 736.050 184.050 ;
        RECT 724.950 178.950 727.050 181.050 ;
        RECT 727.950 178.950 730.050 181.050 ;
        RECT 730.950 178.950 733.050 181.050 ;
        RECT 721.950 175.950 724.050 178.050 ;
        RECT 725.400 176.400 726.600 178.650 ;
        RECT 731.400 177.900 732.600 178.650 ;
        RECT 709.950 163.950 712.050 166.050 ;
        RECT 718.950 163.950 721.050 166.050 ;
        RECT 712.950 148.950 715.050 151.050 ;
        RECT 703.950 142.950 706.050 145.050 ;
        RECT 691.950 141.450 694.050 142.050 ;
        RECT 691.950 140.400 699.450 141.450 ;
        RECT 691.950 139.950 694.050 140.400 ;
        RECT 694.950 137.100 697.050 139.200 ;
        RECT 698.400 139.050 699.450 140.400 ;
        RECT 700.950 139.950 703.050 142.050 ;
        RECT 698.400 138.900 702.000 139.050 ;
        RECT 698.400 137.400 703.050 138.900 ;
        RECT 695.400 136.350 696.600 137.100 ;
        RECT 699.000 136.950 703.050 137.400 ;
        RECT 706.950 137.100 709.050 139.200 ;
        RECT 713.400 138.600 714.450 148.950 ;
        RECT 700.950 136.800 703.050 136.950 ;
        RECT 707.400 136.350 708.600 137.100 ;
        RECT 713.400 136.350 714.600 138.600 ;
        RECT 691.950 133.950 694.050 136.050 ;
        RECT 694.950 133.950 697.050 136.050 ;
        RECT 700.950 133.800 703.050 135.900 ;
        RECT 706.950 133.950 709.050 136.050 ;
        RECT 709.950 133.950 712.050 136.050 ;
        RECT 712.950 133.950 715.050 136.050 ;
        RECT 715.950 133.950 718.050 136.050 ;
        RECT 692.400 132.900 693.600 133.650 ;
        RECT 643.950 121.950 646.050 124.050 ;
        RECT 640.950 112.950 643.050 115.050 ;
        RECT 628.950 104.100 631.050 106.200 ;
        RECT 634.950 104.100 637.050 106.200 ;
        RECT 641.400 106.050 642.450 112.950 ;
        RECT 659.400 108.450 660.450 131.400 ;
        RECT 664.950 127.950 667.050 130.050 ;
        RECT 673.950 127.950 676.050 132.000 ;
        RECT 679.950 130.800 682.050 132.900 ;
        RECT 685.950 130.800 688.050 132.900 ;
        RECT 691.950 130.800 694.050 132.900 ;
        RECT 656.400 107.400 660.450 108.450 ;
        RECT 656.400 106.200 657.450 107.400 ;
        RECT 629.400 103.350 630.600 104.100 ;
        RECT 635.400 103.350 636.600 104.100 ;
        RECT 640.950 103.950 643.050 106.050 ;
        RECT 650.400 105.450 651.600 105.600 ;
        RECT 644.400 104.400 651.600 105.450 ;
        RECT 628.950 100.950 631.050 103.050 ;
        RECT 631.950 100.950 634.050 103.050 ;
        RECT 634.950 100.950 637.050 103.050 ;
        RECT 637.950 100.950 640.050 103.050 ;
        RECT 632.400 99.000 633.600 100.650 ;
        RECT 622.950 94.950 625.050 97.050 ;
        RECT 631.950 94.950 634.050 99.000 ;
        RECT 638.400 98.400 639.600 100.650 ;
        RECT 638.400 85.050 639.450 98.400 ;
        RECT 637.950 82.950 640.050 85.050 ;
        RECT 644.400 79.050 645.450 104.400 ;
        RECT 650.400 103.350 651.600 104.400 ;
        RECT 655.950 104.100 658.050 106.200 ;
        RECT 656.400 103.350 657.600 104.100 ;
        RECT 649.950 100.950 652.050 103.050 ;
        RECT 652.950 100.950 655.050 103.050 ;
        RECT 655.950 100.950 658.050 103.050 ;
        RECT 658.950 100.950 661.050 103.050 ;
        RECT 646.950 97.950 649.050 100.050 ;
        RECT 653.400 99.900 654.600 100.650 ;
        RECT 659.400 99.900 660.600 100.650 ;
        RECT 643.950 76.950 646.050 79.050 ;
        RECT 613.950 70.950 616.050 73.050 ;
        RECT 619.950 70.950 622.050 73.050 ;
        RECT 595.950 64.950 598.050 67.050 ;
        RECT 607.950 64.950 610.050 67.050 ;
        RECT 536.400 58.350 537.600 60.000 ;
        RECT 541.950 59.100 544.050 61.200 ;
        RECT 547.950 59.100 550.050 61.200 ;
        RECT 556.950 59.100 559.050 61.200 ;
        RECT 562.950 59.100 565.050 61.200 ;
        RECT 542.400 58.350 543.600 59.100 ;
        RECT 535.950 55.950 538.050 58.050 ;
        RECT 538.950 55.950 541.050 58.050 ;
        RECT 541.950 55.950 544.050 58.050 ;
        RECT 508.950 49.950 511.050 52.050 ;
        RECT 517.950 49.650 520.050 51.750 ;
        RECT 478.950 40.950 481.050 43.050 ;
        RECT 493.950 40.950 496.050 43.050 ;
        RECT 475.950 37.950 478.050 40.050 ;
        RECT 479.400 27.600 480.450 40.950 ;
        RECT 496.950 37.950 499.050 40.050 ;
        RECT 508.950 37.950 511.050 40.050 ;
        RECT 487.950 34.950 490.050 37.050 ;
        RECT 488.400 30.450 489.450 34.950 ;
        RECT 488.400 29.400 492.450 30.450 ;
        RECT 458.400 25.350 459.600 26.100 ;
        RECT 464.400 25.350 465.600 27.600 ;
        RECT 479.400 25.350 480.600 27.600 ;
        RECT 487.950 26.100 490.050 28.200 ;
        RECT 397.950 22.950 400.050 25.050 ;
        RECT 400.950 22.950 403.050 25.050 ;
        RECT 403.950 22.950 406.050 25.050 ;
        RECT 406.950 22.950 409.050 25.050 ;
        RECT 412.950 22.800 415.050 24.900 ;
        RECT 418.950 22.950 421.050 25.050 ;
        RECT 421.950 22.950 424.050 25.050 ;
        RECT 433.950 22.950 436.050 25.050 ;
        RECT 436.950 22.950 439.050 25.050 ;
        RECT 439.950 22.950 442.050 25.050 ;
        RECT 442.950 22.950 445.050 25.050 ;
        RECT 454.950 22.950 457.050 25.050 ;
        RECT 457.950 22.950 460.050 25.050 ;
        RECT 460.950 22.950 463.050 25.050 ;
        RECT 463.950 22.950 466.050 25.050 ;
        RECT 475.950 22.950 478.050 25.050 ;
        RECT 478.950 22.950 481.050 25.050 ;
        RECT 481.950 22.950 484.050 25.050 ;
        RECT 398.400 21.900 399.600 22.650 ;
        RECT 397.950 19.800 400.050 21.900 ;
        RECT 404.400 21.000 405.600 22.650 ;
        RECT 391.950 16.950 394.050 19.050 ;
        RECT 403.950 16.950 406.050 21.000 ;
        RECT 413.400 16.050 414.450 22.800 ;
        RECT 419.400 21.000 420.600 22.650 ;
        RECT 437.400 21.900 438.600 22.650 ;
        RECT 443.400 21.900 444.600 22.650 ;
        RECT 418.950 16.950 421.050 21.000 ;
        RECT 436.950 19.800 439.050 21.900 ;
        RECT 442.950 19.800 445.050 21.900 ;
        RECT 455.400 21.450 456.600 22.650 ;
        RECT 452.400 20.400 456.600 21.450 ;
        RECT 461.400 20.400 462.600 22.650 ;
        RECT 476.400 21.000 477.600 22.650 ;
        RECT 482.400 21.900 483.600 22.650 ;
        RECT 488.400 22.050 489.450 26.100 ;
        RECT 334.950 13.950 337.050 16.050 ;
        RECT 358.950 13.950 361.050 16.050 ;
        RECT 376.950 15.900 381.000 16.050 ;
        RECT 376.950 15.000 382.050 15.900 ;
        RECT 377.400 14.400 382.050 15.000 ;
        RECT 378.000 13.950 382.050 14.400 ;
        RECT 385.950 13.950 388.050 16.050 ;
        RECT 393.000 15.900 397.050 16.050 ;
        RECT 391.950 13.950 397.050 15.900 ;
        RECT 400.950 13.950 403.050 16.050 ;
        RECT 412.950 13.950 415.050 16.050 ;
        RECT 379.950 13.800 382.050 13.950 ;
        RECT 391.950 13.800 394.050 13.950 ;
        RECT 319.950 7.950 322.050 10.050 ;
        RECT 328.950 7.950 331.050 10.050 ;
        RECT 401.400 9.450 402.450 13.950 ;
        RECT 401.400 8.400 405.450 9.450 ;
        RECT 79.950 4.950 82.050 7.050 ;
        RECT 214.950 4.950 217.050 7.050 ;
        RECT 220.950 4.950 223.050 7.050 ;
        RECT 298.950 4.950 301.050 7.050 ;
        RECT 404.400 6.450 405.450 8.400 ;
        RECT 452.400 7.050 453.450 20.400 ;
        RECT 457.950 16.950 460.050 19.050 ;
        RECT 454.950 13.950 457.050 16.050 ;
        RECT 404.400 5.400 408.450 6.450 ;
        RECT 407.400 3.450 408.450 5.400 ;
        RECT 412.950 3.450 415.050 7.050 ;
        RECT 451.950 4.950 454.050 7.050 ;
        RECT 455.400 6.450 456.450 13.950 ;
        RECT 458.400 10.050 459.450 16.950 ;
        RECT 461.400 13.050 462.450 20.400 ;
        RECT 475.950 16.950 478.050 21.000 ;
        RECT 481.950 19.800 484.050 21.900 ;
        RECT 487.950 19.950 490.050 22.050 ;
        RECT 491.400 16.050 492.450 29.400 ;
        RECT 497.400 27.600 498.450 37.950 ;
        RECT 497.400 25.350 498.600 27.600 ;
        RECT 494.100 22.950 496.200 25.050 ;
        RECT 497.400 22.950 499.500 25.050 ;
        RECT 502.800 22.950 504.900 25.050 ;
        RECT 494.400 21.900 495.600 22.650 ;
        RECT 493.950 19.800 496.050 21.900 ;
        RECT 503.400 20.400 504.600 22.650 ;
        RECT 509.400 21.900 510.450 37.950 ;
        RECT 518.400 27.600 519.450 49.650 ;
        RECT 524.400 37.050 525.450 53.400 ;
        RECT 529.950 52.950 532.050 55.050 ;
        RECT 539.400 54.900 540.600 55.650 ;
        RECT 538.950 52.800 541.050 54.900 ;
        RECT 544.950 52.950 547.050 55.050 ;
        RECT 532.950 37.950 535.050 40.050 ;
        RECT 523.950 34.950 526.050 37.050 ;
        RECT 518.400 25.350 519.600 27.600 ;
        RECT 526.950 25.950 529.050 28.050 ;
        RECT 533.400 27.600 534.450 37.950 ;
        RECT 538.950 31.950 541.050 34.050 ;
        RECT 539.400 27.600 540.450 31.950 ;
        RECT 545.400 28.050 546.450 52.950 ;
        RECT 514.950 22.950 517.050 25.050 ;
        RECT 517.950 22.950 520.050 25.050 ;
        RECT 520.950 22.950 523.050 25.050 ;
        RECT 515.400 21.900 516.600 22.650 ;
        RECT 490.950 13.950 493.050 16.050 ;
        RECT 503.400 13.050 504.450 20.400 ;
        RECT 508.950 19.800 511.050 21.900 ;
        RECT 514.950 19.800 517.050 21.900 ;
        RECT 521.400 21.000 522.600 22.650 ;
        RECT 520.950 16.950 523.050 21.000 ;
        RECT 527.400 19.050 528.450 25.950 ;
        RECT 533.400 25.350 534.600 27.600 ;
        RECT 539.400 25.350 540.600 27.600 ;
        RECT 544.950 25.950 547.050 28.050 ;
        RECT 532.950 22.950 535.050 25.050 ;
        RECT 535.950 22.950 538.050 25.050 ;
        RECT 538.950 22.950 541.050 25.050 ;
        RECT 541.950 22.950 544.050 25.050 ;
        RECT 536.400 20.400 537.600 22.650 ;
        RECT 542.400 20.400 543.600 22.650 ;
        RECT 526.950 16.950 529.050 19.050 ;
        RECT 521.400 13.050 522.450 16.950 ;
        RECT 536.400 13.050 537.450 20.400 ;
        RECT 542.400 16.050 543.450 20.400 ;
        RECT 548.400 16.050 549.450 59.100 ;
        RECT 557.400 58.350 558.600 59.100 ;
        RECT 563.400 58.350 564.600 59.100 ;
        RECT 568.950 58.950 571.050 61.050 ;
        RECT 577.950 59.100 580.050 61.200 ;
        RECT 553.950 55.950 556.050 58.050 ;
        RECT 556.950 55.950 559.050 58.050 ;
        RECT 559.950 55.950 562.050 58.050 ;
        RECT 562.950 55.950 565.050 58.050 ;
        RECT 554.400 53.400 555.600 55.650 ;
        RECT 560.400 53.400 561.600 55.650 ;
        RECT 569.400 54.900 570.450 58.950 ;
        RECT 578.400 58.350 579.600 59.100 ;
        RECT 586.950 58.950 589.050 61.050 ;
        RECT 596.400 60.600 597.450 64.950 ;
        RECT 574.950 55.950 577.050 58.050 ;
        RECT 577.950 55.950 580.050 58.050 ;
        RECT 575.400 54.900 576.600 55.650 ;
        RECT 587.400 54.900 588.450 58.950 ;
        RECT 596.400 58.350 597.600 60.600 ;
        RECT 601.950 59.100 604.050 61.200 ;
        RECT 602.400 58.350 603.600 59.100 ;
        RECT 592.950 55.950 595.050 58.050 ;
        RECT 595.950 55.950 598.050 58.050 ;
        RECT 598.950 55.950 601.050 58.050 ;
        RECT 601.950 55.950 604.050 58.050 ;
        RECT 593.400 54.900 594.600 55.650 ;
        RECT 554.400 34.050 555.450 53.400 ;
        RECT 560.400 40.050 561.450 53.400 ;
        RECT 568.950 52.800 571.050 54.900 ;
        RECT 574.950 52.800 577.050 54.900 ;
        RECT 586.950 52.800 589.050 54.900 ;
        RECT 592.950 52.800 595.050 54.900 ;
        RECT 599.400 53.400 600.600 55.650 ;
        RECT 608.400 54.450 609.450 64.950 ;
        RECT 614.400 63.450 615.450 70.950 ;
        RECT 616.950 63.450 619.050 67.050 ;
        RECT 643.950 64.950 646.050 67.050 ;
        RECT 614.400 63.000 619.050 63.450 ;
        RECT 614.400 62.400 618.450 63.000 ;
        RECT 617.400 60.600 618.450 62.400 ;
        RECT 617.400 58.350 618.600 60.600 ;
        RECT 622.950 59.100 625.050 61.200 ;
        RECT 637.950 59.100 640.050 61.200 ;
        RECT 644.400 60.600 645.450 64.950 ;
        RECT 623.400 58.350 624.600 59.100 ;
        RECT 638.400 58.350 639.600 59.100 ;
        RECT 644.400 58.350 645.600 60.600 ;
        RECT 647.400 60.450 648.450 97.950 ;
        RECT 652.950 94.950 655.050 99.900 ;
        RECT 658.950 97.800 661.050 99.900 ;
        RECT 661.950 97.950 664.050 100.050 ;
        RECT 665.400 99.900 666.450 127.950 ;
        RECT 685.950 118.950 688.050 121.050 ;
        RECT 694.950 118.950 697.050 121.050 ;
        RECT 679.950 112.950 682.050 115.050 ;
        RECT 667.950 103.950 670.050 109.050 ;
        RECT 673.950 104.100 676.050 106.200 ;
        RECT 680.400 105.600 681.450 112.950 ;
        RECT 674.400 103.350 675.600 104.100 ;
        RECT 680.400 103.350 681.600 105.600 ;
        RECT 670.950 100.950 673.050 103.050 ;
        RECT 673.950 100.950 676.050 103.050 ;
        RECT 676.950 100.950 679.050 103.050 ;
        RECT 679.950 100.950 682.050 103.050 ;
        RECT 655.950 82.950 658.050 85.050 ;
        RECT 652.950 64.950 655.050 67.050 ;
        RECT 647.400 59.400 651.450 60.450 ;
        RECT 613.950 55.950 616.050 58.050 ;
        RECT 616.950 55.950 619.050 58.050 ;
        RECT 619.950 55.950 622.050 58.050 ;
        RECT 622.950 55.950 625.050 58.050 ;
        RECT 634.950 55.950 637.050 58.050 ;
        RECT 637.950 55.950 640.050 58.050 ;
        RECT 640.950 55.950 643.050 58.050 ;
        RECT 643.950 55.950 646.050 58.050 ;
        RECT 614.400 54.450 615.600 55.650 ;
        RECT 608.400 53.400 615.600 54.450 ;
        RECT 620.400 53.400 621.600 55.650 ;
        RECT 635.400 54.900 636.600 55.650 ;
        RECT 559.950 37.950 562.050 40.050 ;
        RECT 553.950 31.950 556.050 34.050 ;
        RECT 559.950 26.100 562.050 28.200 ;
        RECT 565.950 26.100 568.050 28.200 ;
        RECT 575.400 28.050 576.450 52.800 ;
        RECT 583.950 37.950 586.050 40.050 ;
        RECT 560.400 25.350 561.600 26.100 ;
        RECT 566.400 25.350 567.600 26.100 ;
        RECT 574.950 25.950 577.050 28.050 ;
        RECT 577.950 26.100 580.050 28.200 ;
        RECT 584.400 27.600 585.450 37.950 ;
        RECT 593.400 31.050 594.450 52.800 ;
        RECT 592.950 28.950 595.050 31.050 ;
        RECT 599.400 30.450 600.450 53.400 ;
        RECT 620.400 49.050 621.450 53.400 ;
        RECT 634.950 52.800 637.050 54.900 ;
        RECT 641.400 53.400 642.600 55.650 ;
        RECT 619.950 46.950 622.050 49.050 ;
        RECT 635.400 40.050 636.450 52.800 ;
        RECT 641.400 49.050 642.450 53.400 ;
        RECT 646.950 52.950 649.050 55.050 ;
        RECT 640.950 46.950 643.050 49.050 ;
        RECT 647.400 43.050 648.450 52.950 ;
        RECT 646.950 40.950 649.050 43.050 ;
        RECT 634.950 37.950 637.050 40.050 ;
        RECT 643.950 34.950 646.050 37.050 ;
        RECT 644.400 31.050 645.450 34.950 ;
        RECT 596.400 29.400 600.450 30.450 ;
        RECT 578.400 25.350 579.600 26.100 ;
        RECT 584.400 25.350 585.600 27.600 ;
        RECT 596.400 27.450 597.450 29.400 ;
        RECT 643.950 28.950 646.050 31.050 ;
        RECT 593.400 26.400 597.450 27.450 ;
        RECT 556.950 22.950 559.050 25.050 ;
        RECT 559.950 22.950 562.050 25.050 ;
        RECT 562.950 22.950 565.050 25.050 ;
        RECT 565.950 22.950 568.050 25.050 ;
        RECT 577.950 22.950 580.050 25.050 ;
        RECT 580.950 22.950 583.050 25.050 ;
        RECT 583.950 22.950 586.050 25.050 ;
        RECT 586.950 22.950 589.050 25.050 ;
        RECT 557.400 20.400 558.600 22.650 ;
        RECT 563.400 21.900 564.600 22.650 ;
        RECT 581.400 21.900 582.600 22.650 ;
        RECT 587.400 21.900 588.600 22.650 ;
        RECT 541.950 13.950 544.050 16.050 ;
        RECT 547.950 13.950 550.050 16.050 ;
        RECT 460.950 10.950 463.050 13.050 ;
        RECT 502.950 10.950 505.050 13.050 ;
        RECT 520.950 10.950 523.050 13.050 ;
        RECT 535.950 10.950 538.050 13.050 ;
        RECT 457.950 7.950 460.050 10.050 ;
        RECT 557.400 7.050 558.450 20.400 ;
        RECT 562.950 19.800 565.050 21.900 ;
        RECT 574.950 16.950 577.050 21.900 ;
        RECT 580.950 19.800 583.050 21.900 ;
        RECT 586.950 19.800 589.050 21.900 ;
        RECT 587.400 16.050 588.450 19.800 ;
        RECT 586.950 13.950 589.050 16.050 ;
        RECT 593.400 7.050 594.450 26.400 ;
        RECT 598.950 26.100 601.050 28.200 ;
        RECT 604.950 26.100 607.050 28.200 ;
        RECT 613.950 26.100 616.050 28.200 ;
        RECT 616.950 27.600 621.000 28.050 ;
        RECT 599.400 25.350 600.600 26.100 ;
        RECT 605.400 25.350 606.600 26.100 ;
        RECT 598.950 22.950 601.050 25.050 ;
        RECT 601.950 22.950 604.050 25.050 ;
        RECT 604.950 22.950 607.050 25.050 ;
        RECT 607.950 22.950 610.050 25.050 ;
        RECT 602.400 21.900 603.600 22.650 ;
        RECT 608.400 21.900 609.600 22.650 ;
        RECT 595.950 19.800 598.050 21.900 ;
        RECT 601.950 19.800 604.050 21.900 ;
        RECT 607.950 19.800 610.050 21.900 ;
        RECT 610.950 19.950 613.050 22.050 ;
        RECT 460.950 6.450 463.050 7.050 ;
        RECT 455.400 5.400 463.050 6.450 ;
        RECT 460.950 4.950 463.050 5.400 ;
        RECT 556.950 4.950 559.050 7.050 ;
        RECT 592.950 4.950 595.050 7.050 ;
        RECT 596.400 4.050 597.450 19.800 ;
        RECT 611.400 13.050 612.450 19.950 ;
        RECT 614.400 16.050 615.450 26.100 ;
        RECT 616.950 25.950 621.600 27.600 ;
        RECT 625.950 26.100 628.050 28.200 ;
        RECT 620.400 25.350 621.600 25.950 ;
        RECT 626.400 25.350 627.600 26.100 ;
        RECT 634.950 25.950 637.050 28.050 ;
        RECT 640.950 26.100 643.050 28.200 ;
        RECT 647.400 27.600 648.450 40.950 ;
        RECT 650.400 34.050 651.450 59.400 ;
        RECT 653.400 51.450 654.450 64.950 ;
        RECT 656.400 61.050 657.450 82.950 ;
        RECT 662.400 63.450 663.450 97.950 ;
        RECT 664.950 97.800 667.050 99.900 ;
        RECT 671.400 99.000 672.600 100.650 ;
        RECT 677.400 99.900 678.600 100.650 ;
        RECT 659.400 62.400 663.450 63.450 ;
        RECT 655.950 58.950 658.050 61.050 ;
        RECT 659.400 60.600 660.450 62.400 ;
        RECT 665.400 60.600 666.450 97.800 ;
        RECT 670.950 94.950 673.050 99.000 ;
        RECT 676.950 97.800 679.050 99.900 ;
        RECT 686.400 85.050 687.450 118.950 ;
        RECT 695.400 105.600 696.450 118.950 ;
        RECT 701.400 109.200 702.450 133.800 ;
        RECT 710.400 132.900 711.600 133.650 ;
        RECT 716.400 132.900 717.600 133.650 ;
        RECT 709.950 130.800 712.050 132.900 ;
        RECT 715.950 130.800 718.050 132.900 ;
        RECT 722.400 121.050 723.450 175.950 ;
        RECT 725.400 169.050 726.450 176.400 ;
        RECT 730.950 175.800 733.050 177.900 ;
        RECT 724.950 166.950 727.050 169.050 ;
        RECT 733.950 160.950 736.050 163.050 ;
        RECT 734.400 141.450 735.450 160.950 ;
        RECT 737.400 157.050 738.450 185.400 ;
        RECT 739.950 181.950 742.050 184.050 ;
        RECT 745.950 182.100 748.050 184.200 ;
        RECT 752.400 183.600 753.450 187.950 ;
        RECT 736.950 154.950 739.050 157.050 ;
        RECT 740.400 154.050 741.450 181.950 ;
        RECT 746.400 181.350 747.600 182.100 ;
        RECT 752.400 181.350 753.600 183.600 ;
        RECT 755.400 183.450 756.450 202.950 ;
        RECT 758.400 187.050 759.450 254.400 ;
        RECT 760.950 253.950 763.050 256.050 ;
        RECT 761.400 205.050 762.450 253.950 ;
        RECT 764.400 253.050 765.450 277.950 ;
        RECT 767.400 274.050 768.450 287.400 ;
        RECT 772.950 286.950 775.050 289.050 ;
        RECT 773.400 280.050 774.450 286.950 ;
        RECT 772.950 277.950 775.050 280.050 ;
        RECT 766.950 271.950 769.050 274.050 ;
        RECT 776.400 268.050 777.450 332.400 ;
        RECT 778.950 322.950 781.050 325.050 ;
        RECT 779.400 316.050 780.450 322.950 ;
        RECT 778.950 313.950 781.050 316.050 ;
        RECT 778.950 307.950 781.050 310.050 ;
        RECT 779.400 295.050 780.450 307.950 ;
        RECT 784.950 298.950 787.050 301.050 ;
        RECT 778.950 292.950 781.050 295.050 ;
        RECT 785.400 294.600 786.450 298.950 ;
        RECT 785.400 292.350 786.600 294.600 ;
        RECT 790.950 293.100 793.050 295.200 ;
        RECT 794.400 295.050 795.450 332.400 ;
        RECT 796.950 331.950 799.050 334.050 ;
        RECT 803.400 333.450 804.600 334.650 ;
        RECT 809.400 333.900 810.600 334.650 ;
        RECT 800.400 332.400 804.600 333.450 ;
        RECT 797.400 319.050 798.450 331.950 ;
        RECT 800.400 328.050 801.450 332.400 ;
        RECT 808.950 328.950 811.050 333.900 ;
        RECT 814.950 331.950 817.050 334.050 ;
        RECT 799.950 325.950 802.050 328.050 ;
        RECT 796.950 316.950 799.050 319.050 ;
        RECT 796.950 304.950 799.050 307.050 ;
        RECT 797.400 298.050 798.450 304.950 ;
        RECT 800.400 304.050 801.450 325.950 ;
        RECT 802.950 319.950 805.050 322.050 ;
        RECT 799.950 301.950 802.050 304.050 ;
        RECT 796.950 295.950 799.050 298.050 ;
        RECT 791.400 292.350 792.600 293.100 ;
        RECT 793.950 292.950 796.050 295.050 ;
        RECT 781.950 289.950 784.050 292.050 ;
        RECT 784.950 289.950 787.050 292.050 ;
        RECT 787.950 289.950 790.050 292.050 ;
        RECT 790.950 289.950 793.050 292.050 ;
        RECT 782.400 288.000 783.600 289.650 ;
        RECT 788.400 288.900 789.600 289.650 ;
        RECT 781.950 283.950 784.050 288.000 ;
        RECT 787.950 286.800 790.050 288.900 ;
        RECT 793.950 286.950 796.050 289.050 ;
        RECT 784.950 280.950 787.050 283.050 ;
        RECT 766.950 265.950 769.050 268.050 ;
        RECT 775.950 265.950 778.050 268.050 ;
        RECT 767.400 262.050 768.450 265.950 ;
        RECT 766.950 259.950 769.050 262.050 ;
        RECT 772.950 260.100 775.050 262.200 ;
        RECT 785.400 262.050 786.450 280.950 ;
        RECT 794.400 279.450 795.450 286.950 ;
        RECT 797.400 283.050 798.450 295.950 ;
        RECT 799.950 294.450 802.050 298.050 ;
        RECT 803.400 295.200 804.450 319.950 ;
        RECT 815.400 316.050 816.450 331.950 ;
        RECT 818.400 322.050 819.450 340.950 ;
        RECT 826.950 339.000 829.050 342.900 ;
        RECT 829.950 340.950 832.050 343.050 ;
        RECT 833.400 339.600 834.450 364.800 ;
        RECT 838.950 358.950 841.050 361.050 ;
        RECT 835.950 352.950 838.050 355.050 ;
        RECT 836.400 349.050 837.450 352.950 ;
        RECT 835.950 346.950 838.050 349.050 ;
        RECT 835.950 343.800 838.050 345.900 ;
        RECT 836.400 340.050 837.450 343.800 ;
        RECT 827.400 337.350 828.600 339.000 ;
        RECT 833.400 337.350 834.600 339.600 ;
        RECT 835.950 337.950 838.050 340.050 ;
        RECT 823.950 334.950 826.050 337.050 ;
        RECT 826.950 334.950 829.050 337.050 ;
        RECT 829.950 334.950 832.050 337.050 ;
        RECT 832.950 334.950 835.050 337.050 ;
        RECT 824.400 332.400 825.600 334.650 ;
        RECT 830.400 333.900 831.600 334.650 ;
        RECT 824.400 328.050 825.450 332.400 ;
        RECT 829.950 331.800 832.050 333.900 ;
        RECT 835.950 331.950 838.050 334.050 ;
        RECT 829.950 328.650 832.050 330.750 ;
        RECT 823.950 325.950 826.050 328.050 ;
        RECT 817.950 319.950 820.050 322.050 ;
        RECT 817.800 316.800 819.900 318.900 ;
        RECT 820.950 316.950 823.050 319.050 ;
        RECT 814.950 313.950 817.050 316.050 ;
        RECT 802.950 294.450 805.050 295.200 ;
        RECT 799.950 294.000 805.050 294.450 ;
        RECT 808.950 294.000 811.050 298.050 ;
        RECT 800.400 293.400 805.050 294.000 ;
        RECT 802.950 293.100 805.050 293.400 ;
        RECT 803.400 292.350 804.600 293.100 ;
        RECT 809.400 292.350 810.600 294.000 ;
        RECT 802.950 289.950 805.050 292.050 ;
        RECT 805.950 289.950 808.050 292.050 ;
        RECT 808.950 289.950 811.050 292.050 ;
        RECT 811.950 289.950 814.050 292.050 ;
        RECT 806.400 287.400 807.600 289.650 ;
        RECT 812.400 287.400 813.600 289.650 ;
        RECT 802.950 283.950 805.050 286.050 ;
        RECT 796.950 280.950 799.050 283.050 ;
        RECT 794.400 278.400 798.450 279.450 ;
        RECT 787.950 268.950 790.050 271.050 ;
        RECT 793.950 268.950 796.050 271.050 ;
        RECT 773.400 259.350 774.600 260.100 ;
        RECT 781.950 259.950 784.050 262.050 ;
        RECT 784.950 259.950 787.050 262.050 ;
        RECT 788.400 261.600 789.450 268.950 ;
        RECT 794.400 262.200 795.450 268.950 ;
        RECT 797.400 265.050 798.450 278.400 ;
        RECT 799.950 277.950 802.050 280.050 ;
        RECT 800.400 274.050 801.450 277.950 ;
        RECT 799.950 271.950 802.050 274.050 ;
        RECT 796.950 262.950 799.050 265.050 ;
        RECT 769.950 256.950 772.050 259.050 ;
        RECT 772.950 256.950 775.050 259.050 ;
        RECT 775.950 256.950 778.050 259.050 ;
        RECT 770.400 254.400 771.600 256.650 ;
        RECT 776.400 255.900 777.600 256.650 ;
        RECT 782.400 255.900 783.450 259.950 ;
        RECT 788.400 259.350 789.600 261.600 ;
        RECT 793.950 260.100 796.050 262.200 ;
        RECT 794.400 259.350 795.600 260.100 ;
        RECT 787.950 256.950 790.050 259.050 ;
        RECT 790.950 256.950 793.050 259.050 ;
        RECT 793.950 256.950 796.050 259.050 ;
        RECT 796.950 256.950 799.050 259.050 ;
        RECT 763.950 250.950 766.050 253.050 ;
        RECT 770.400 247.050 771.450 254.400 ;
        RECT 775.950 253.800 778.050 255.900 ;
        RECT 781.950 253.800 784.050 255.900 ;
        RECT 784.950 253.950 787.050 256.050 ;
        RECT 791.400 254.400 792.600 256.650 ;
        RECT 797.400 255.450 798.600 256.650 ;
        RECT 797.400 254.400 801.450 255.450 ;
        RECT 778.950 250.950 781.050 253.050 ;
        RECT 769.950 244.950 772.050 247.050 ;
        RECT 763.950 241.950 766.050 244.050 ;
        RECT 764.400 217.050 765.450 241.950 ;
        RECT 779.400 238.050 780.450 250.950 ;
        RECT 785.400 240.450 786.450 253.950 ;
        RECT 785.400 239.400 789.450 240.450 ;
        RECT 778.950 235.950 781.050 238.050 ;
        RECT 784.950 235.950 787.050 238.050 ;
        RECT 766.950 232.950 769.050 235.050 ;
        RECT 763.950 214.950 766.050 217.050 ;
        RECT 767.400 216.600 768.450 232.950 ;
        RECT 772.950 220.950 775.050 223.050 ;
        RECT 773.400 216.600 774.450 220.950 ;
        RECT 779.400 217.200 780.450 235.950 ;
        RECT 767.400 214.350 768.600 216.600 ;
        RECT 773.400 214.350 774.600 216.600 ;
        RECT 778.950 215.100 781.050 217.200 ;
        RECT 779.400 214.350 780.600 215.100 ;
        RECT 766.950 211.950 769.050 214.050 ;
        RECT 769.950 211.950 772.050 214.050 ;
        RECT 772.950 211.950 775.050 214.050 ;
        RECT 775.950 211.950 778.050 214.050 ;
        RECT 778.950 211.950 781.050 214.050 ;
        RECT 763.950 208.950 766.050 211.050 ;
        RECT 760.950 202.950 763.050 205.050 ;
        RECT 764.400 199.050 765.450 208.950 ;
        RECT 785.400 208.050 786.450 235.950 ;
        RECT 778.950 205.950 781.050 208.050 ;
        RECT 784.950 205.950 787.050 208.050 ;
        RECT 766.950 199.950 769.050 202.050 ;
        RECT 763.950 196.950 766.050 199.050 ;
        RECT 767.400 187.050 768.450 199.950 ;
        RECT 769.950 187.950 772.050 190.050 ;
        RECT 757.950 184.950 760.050 187.050 ;
        RECT 766.950 184.950 769.050 187.050 ;
        RECT 755.400 182.400 759.450 183.450 ;
        RECT 745.950 178.950 748.050 181.050 ;
        RECT 748.950 178.950 751.050 181.050 ;
        RECT 751.950 178.950 754.050 181.050 ;
        RECT 742.950 175.950 745.050 178.050 ;
        RECT 749.400 177.900 750.600 178.650 ;
        RECT 739.950 151.950 742.050 154.050 ;
        RECT 734.400 140.400 738.450 141.450 ;
        RECT 724.950 137.100 727.050 139.200 ;
        RECT 730.950 137.100 733.050 139.200 ;
        RECT 737.400 138.600 738.450 140.400 ;
        RECT 725.400 133.050 726.450 137.100 ;
        RECT 731.400 136.350 732.600 137.100 ;
        RECT 737.400 136.350 738.600 138.600 ;
        RECT 730.950 133.950 733.050 136.050 ;
        RECT 733.950 133.950 736.050 136.050 ;
        RECT 736.950 133.950 739.050 136.050 ;
        RECT 724.950 130.950 727.050 133.050 ;
        RECT 734.400 132.000 735.600 133.650 ;
        RECT 725.400 127.050 726.450 130.950 ;
        RECT 733.950 127.950 736.050 132.000 ;
        RECT 724.950 124.950 727.050 127.050 ;
        RECT 721.950 118.950 724.050 121.050 ;
        RECT 727.950 112.950 730.050 115.050 ;
        RECT 736.950 112.950 739.050 115.050 ;
        RECT 700.950 107.100 703.050 109.200 ;
        RECT 706.950 106.950 709.050 109.050 ;
        RECT 695.400 103.350 696.600 105.600 ;
        RECT 700.950 103.950 703.050 106.050 ;
        RECT 701.400 103.350 702.600 103.950 ;
        RECT 691.950 100.950 694.050 103.050 ;
        RECT 694.950 100.950 697.050 103.050 ;
        RECT 697.950 100.950 700.050 103.050 ;
        RECT 700.950 100.950 703.050 103.050 ;
        RECT 692.400 98.400 693.600 100.650 ;
        RECT 698.400 98.400 699.600 100.650 ;
        RECT 673.950 82.950 676.050 85.050 ;
        RECT 685.950 82.950 688.050 85.050 ;
        RECT 659.400 58.350 660.600 60.600 ;
        RECT 665.400 58.350 666.600 60.600 ;
        RECT 658.950 55.950 661.050 58.050 ;
        RECT 661.950 55.950 664.050 58.050 ;
        RECT 664.950 55.950 667.050 58.050 ;
        RECT 667.950 55.950 670.050 58.050 ;
        RECT 662.400 54.900 663.600 55.650 ;
        RECT 661.950 52.800 664.050 54.900 ;
        RECT 668.400 53.400 669.600 55.650 ;
        RECT 653.400 50.400 657.450 51.450 ;
        RECT 652.950 46.950 655.050 49.050 ;
        RECT 649.950 31.950 652.050 34.050 ;
        RECT 653.400 28.050 654.450 46.950 ;
        RECT 656.400 42.450 657.450 50.400 ;
        RECT 668.400 46.050 669.450 53.400 ;
        RECT 674.400 52.050 675.450 82.950 ;
        RECT 692.400 82.050 693.450 98.400 ;
        RECT 698.400 94.050 699.450 98.400 ;
        RECT 697.950 91.950 700.050 94.050 ;
        RECT 691.950 79.950 694.050 82.050 ;
        RECT 682.950 70.950 685.050 73.050 ;
        RECT 683.400 64.050 684.450 70.950 ;
        RECT 707.400 67.050 708.450 106.950 ;
        RECT 712.950 104.100 715.050 106.200 ;
        RECT 718.950 104.100 721.050 106.200 ;
        RECT 713.400 103.350 714.600 104.100 ;
        RECT 719.400 103.350 720.600 104.100 ;
        RECT 712.950 100.950 715.050 103.050 ;
        RECT 715.950 100.950 718.050 103.050 ;
        RECT 718.950 100.950 721.050 103.050 ;
        RECT 721.950 100.950 724.050 103.050 ;
        RECT 716.400 98.400 717.600 100.650 ;
        RECT 722.400 99.900 723.600 100.650 ;
        RECT 712.950 88.950 715.050 91.050 ;
        RECT 694.950 64.950 697.050 67.050 ;
        RECT 706.950 64.950 709.050 67.050 ;
        RECT 682.950 61.950 685.050 64.050 ;
        RECT 683.400 60.600 684.450 61.950 ;
        RECT 683.400 58.350 684.600 60.600 ;
        RECT 688.950 59.100 691.050 61.200 ;
        RECT 689.400 58.350 690.600 59.100 ;
        RECT 679.950 55.950 682.050 58.050 ;
        RECT 682.950 55.950 685.050 58.050 ;
        RECT 685.950 55.950 688.050 58.050 ;
        RECT 688.950 55.950 691.050 58.050 ;
        RECT 676.950 52.800 679.050 54.900 ;
        RECT 680.400 53.400 681.600 55.650 ;
        RECT 686.400 54.900 687.600 55.650 ;
        RECT 673.950 49.950 676.050 52.050 ;
        RECT 677.400 46.050 678.450 52.800 ;
        RECT 680.400 49.050 681.450 53.400 ;
        RECT 685.950 52.800 688.050 54.900 ;
        RECT 679.950 46.950 682.050 49.050 ;
        RECT 667.950 43.950 670.050 46.050 ;
        RECT 676.950 43.950 679.050 46.050 ;
        RECT 656.400 41.400 660.450 42.450 ;
        RECT 655.950 37.950 658.050 40.050 ;
        RECT 619.950 22.950 622.050 25.050 ;
        RECT 622.950 22.950 625.050 25.050 ;
        RECT 625.950 22.950 628.050 25.050 ;
        RECT 628.950 22.950 631.050 25.050 ;
        RECT 623.400 21.900 624.600 22.650 ;
        RECT 629.400 21.900 630.600 22.650 ;
        RECT 622.950 16.950 625.050 21.900 ;
        RECT 628.950 19.800 631.050 21.900 ;
        RECT 635.400 19.050 636.450 25.950 ;
        RECT 641.400 25.350 642.600 26.100 ;
        RECT 647.400 25.350 648.600 27.600 ;
        RECT 652.950 25.950 655.050 28.050 ;
        RECT 640.950 22.950 643.050 25.050 ;
        RECT 643.950 22.950 646.050 25.050 ;
        RECT 646.950 22.950 649.050 25.050 ;
        RECT 649.950 22.950 652.050 25.050 ;
        RECT 644.400 21.900 645.600 22.650 ;
        RECT 650.400 21.900 651.600 22.650 ;
        RECT 643.950 19.800 646.050 21.900 ;
        RECT 649.950 19.800 652.050 21.900 ;
        RECT 634.950 16.950 637.050 19.050 ;
        RECT 656.400 16.050 657.450 37.950 ;
        RECT 659.400 28.050 660.450 41.400 ;
        RECT 664.950 37.950 667.050 40.050 ;
        RECT 658.950 25.950 661.050 28.050 ;
        RECT 665.400 27.600 666.450 37.950 ;
        RECT 676.950 34.950 679.050 37.050 ;
        RECT 665.400 25.350 666.600 27.600 ;
        RECT 670.950 27.000 673.050 31.050 ;
        RECT 671.400 25.350 672.600 27.000 ;
        RECT 661.950 22.950 664.050 25.050 ;
        RECT 664.950 22.950 667.050 25.050 ;
        RECT 667.950 22.950 670.050 25.050 ;
        RECT 670.950 22.950 673.050 25.050 ;
        RECT 662.400 21.900 663.600 22.650 ;
        RECT 661.950 19.800 664.050 21.900 ;
        RECT 668.400 20.400 669.600 22.650 ;
        RECT 668.400 16.050 669.450 20.400 ;
        RECT 673.800 19.950 675.900 22.050 ;
        RECT 677.400 21.900 678.450 34.950 ;
        RECT 685.950 26.100 688.050 28.200 ;
        RECT 691.950 26.100 694.050 31.050 ;
        RECT 695.400 27.450 696.450 64.950 ;
        RECT 700.950 60.000 703.050 64.050 ;
        RECT 713.400 61.200 714.450 88.950 ;
        RECT 716.400 88.050 717.450 98.400 ;
        RECT 721.950 97.800 724.050 99.900 ;
        RECT 728.400 91.050 729.450 112.950 ;
        RECT 737.400 106.200 738.450 112.950 ;
        RECT 743.400 106.200 744.450 175.950 ;
        RECT 748.950 175.800 751.050 177.900 ;
        RECT 749.400 151.050 750.450 175.800 ;
        RECT 758.400 151.050 759.450 182.400 ;
        RECT 763.950 182.100 766.050 184.200 ;
        RECT 770.400 183.600 771.450 187.950 ;
        RECT 764.400 181.350 765.600 182.100 ;
        RECT 770.400 181.350 771.600 183.600 ;
        RECT 763.950 178.950 766.050 181.050 ;
        RECT 766.950 178.950 769.050 181.050 ;
        RECT 769.950 178.950 772.050 181.050 ;
        RECT 772.950 178.950 775.050 181.050 ;
        RECT 760.950 175.950 763.050 178.050 ;
        RECT 767.400 176.400 768.600 178.650 ;
        RECT 773.400 177.900 774.600 178.650 ;
        RECT 748.950 150.450 751.050 151.050 ;
        RECT 746.400 149.400 751.050 150.450 ;
        RECT 746.400 139.050 747.450 149.400 ;
        RECT 748.950 148.950 751.050 149.400 ;
        RECT 757.950 148.950 760.050 151.050 ;
        RECT 757.950 142.950 760.050 145.050 ;
        RECT 745.950 136.950 748.050 139.050 ;
        RECT 751.950 137.100 754.050 139.200 ;
        RECT 758.400 138.600 759.450 142.950 ;
        RECT 761.400 139.050 762.450 175.950 ;
        RECT 752.400 136.350 753.600 137.100 ;
        RECT 758.400 136.350 759.600 138.600 ;
        RECT 760.950 136.950 763.050 139.050 ;
        RECT 763.950 138.450 766.050 139.200 ;
        RECT 767.400 138.450 768.450 176.400 ;
        RECT 772.950 175.800 775.050 177.900 ;
        RECT 773.400 163.050 774.450 175.800 ;
        RECT 772.950 160.950 775.050 163.050 ;
        RECT 775.950 157.950 778.050 160.050 ;
        RECT 763.950 137.400 768.450 138.450 ;
        RECT 763.950 137.100 766.050 137.400 ;
        RECT 769.950 137.100 772.050 139.200 ;
        RECT 776.400 138.600 777.450 157.950 ;
        RECT 779.400 157.050 780.450 205.950 ;
        RECT 788.400 205.050 789.450 239.400 ;
        RECT 787.950 202.950 790.050 205.050 ;
        RECT 791.400 202.050 792.450 254.400 ;
        RECT 800.400 250.050 801.450 254.400 ;
        RECT 799.950 247.950 802.050 250.050 ;
        RECT 803.400 238.050 804.450 283.950 ;
        RECT 806.400 280.050 807.450 287.400 ;
        RECT 805.950 277.950 808.050 280.050 ;
        RECT 806.400 274.050 807.450 277.950 ;
        RECT 812.400 277.050 813.450 287.400 ;
        RECT 814.950 286.950 817.050 289.050 ;
        RECT 811.950 274.950 814.050 277.050 ;
        RECT 805.950 271.950 808.050 274.050 ;
        RECT 811.950 271.800 814.050 273.900 ;
        RECT 812.400 261.600 813.450 271.800 ;
        RECT 815.400 265.050 816.450 286.950 ;
        RECT 818.400 277.050 819.450 316.800 ;
        RECT 821.400 295.050 822.450 316.950 ;
        RECT 826.950 307.950 829.050 310.050 ;
        RECT 820.950 292.950 823.050 295.050 ;
        RECT 827.400 294.600 828.450 307.950 ;
        RECT 830.400 298.050 831.450 328.650 ;
        RECT 836.400 319.050 837.450 331.950 ;
        RECT 835.950 316.950 838.050 319.050 ;
        RECT 829.950 295.950 832.050 298.050 ;
        RECT 827.400 292.350 828.600 294.600 ;
        RECT 832.950 293.100 835.050 295.200 ;
        RECT 833.400 292.350 834.600 293.100 ;
        RECT 839.400 292.050 840.450 358.950 ;
        RECT 842.400 355.050 843.450 365.400 ;
        RECT 847.950 364.800 850.050 366.900 ;
        RECT 853.800 364.950 855.900 367.050 ;
        RECT 856.950 364.950 859.050 367.050 ;
        RECT 863.400 365.400 868.050 367.050 ;
        RECT 864.000 364.950 868.050 365.400 ;
        RECT 841.950 352.950 844.050 355.050 ;
        RECT 850.950 352.950 853.050 355.050 ;
        RECT 841.950 346.950 844.050 349.050 ;
        RECT 842.400 337.050 843.450 346.950 ;
        RECT 844.950 343.950 847.050 346.050 ;
        RECT 845.400 339.600 846.450 343.950 ;
        RECT 851.400 342.450 852.450 352.950 ;
        RECT 854.400 346.050 855.450 364.950 ;
        RECT 853.950 343.950 856.050 346.050 ;
        RECT 851.400 341.400 855.450 342.450 ;
        RECT 845.400 337.350 846.600 339.600 ;
        RECT 841.950 334.950 844.050 337.050 ;
        RECT 845.400 334.950 847.500 337.050 ;
        RECT 850.800 334.950 852.900 337.050 ;
        RECT 841.950 331.800 844.050 333.900 ;
        RECT 823.950 289.950 826.050 292.050 ;
        RECT 826.950 289.950 829.050 292.050 ;
        RECT 829.950 289.950 832.050 292.050 ;
        RECT 832.950 289.950 835.050 292.050 ;
        RECT 838.950 289.950 841.050 292.050 ;
        RECT 824.400 288.900 825.600 289.650 ;
        RECT 823.950 286.800 826.050 288.900 ;
        RECT 830.400 287.400 831.600 289.650 ;
        RECT 817.950 274.950 820.050 277.050 ;
        RECT 814.950 262.950 817.050 265.050 ;
        RECT 812.400 259.350 813.600 261.600 ;
        RECT 817.950 260.100 820.050 262.200 ;
        RECT 818.400 259.350 819.600 260.100 ;
        RECT 808.950 256.950 811.050 259.050 ;
        RECT 811.950 256.950 814.050 259.050 ;
        RECT 814.950 256.950 817.050 259.050 ;
        RECT 817.950 256.950 820.050 259.050 ;
        RECT 809.400 255.900 810.600 256.650 ;
        RECT 808.950 253.800 811.050 255.900 ;
        RECT 815.400 254.400 816.600 256.650 ;
        RECT 815.400 252.450 816.450 254.400 ;
        RECT 812.400 251.400 816.450 252.450 ;
        RECT 812.400 238.050 813.450 251.400 ;
        RECT 824.400 250.050 825.450 286.800 ;
        RECT 830.400 277.050 831.450 287.400 ;
        RECT 835.950 286.950 838.050 289.050 ;
        RECT 829.950 274.950 832.050 277.050 ;
        RECT 836.400 274.050 837.450 286.950 ;
        RECT 835.950 271.950 838.050 274.050 ;
        RECT 829.950 268.950 832.050 271.050 ;
        RECT 830.400 261.600 831.450 268.950 ;
        RECT 842.400 268.050 843.450 331.800 ;
        RECT 854.400 331.050 855.450 341.400 ;
        RECT 857.400 331.050 858.450 364.950 ;
        RECT 859.950 343.950 862.050 346.050 ;
        RECT 844.950 328.950 847.050 331.050 ;
        RECT 853.950 328.950 856.050 331.050 ;
        RECT 856.950 328.950 859.050 331.050 ;
        RECT 845.400 294.600 846.450 328.950 ;
        RECT 853.950 322.950 856.050 325.050 ;
        RECT 854.400 294.600 855.450 322.950 ;
        RECT 856.950 295.950 859.050 298.050 ;
        RECT 845.400 292.350 846.600 294.600 ;
        RECT 854.400 292.350 855.600 294.600 ;
        RECT 845.100 289.950 847.200 292.050 ;
        RECT 848.400 289.950 850.500 292.050 ;
        RECT 853.800 289.950 855.900 292.050 ;
        RECT 848.400 287.400 849.600 289.650 ;
        RECT 848.400 280.050 849.450 287.400 ;
        RECT 847.950 277.950 850.050 280.050 ;
        RECT 847.950 271.950 850.050 274.050 ;
        RECT 841.950 265.950 844.050 268.050 ;
        RECT 830.400 259.350 831.600 261.600 ;
        RECT 835.950 260.100 838.050 262.200 ;
        RECT 844.950 260.100 847.050 262.200 ;
        RECT 848.400 262.050 849.450 271.950 ;
        RECT 836.400 259.350 837.600 260.100 ;
        RECT 829.950 256.950 832.050 259.050 ;
        RECT 832.950 256.950 835.050 259.050 ;
        RECT 835.950 256.950 838.050 259.050 ;
        RECT 838.950 256.950 841.050 259.050 ;
        RECT 833.400 254.400 834.600 256.650 ;
        RECT 839.400 255.450 840.600 256.650 ;
        RECT 845.400 255.450 846.450 260.100 ;
        RECT 847.950 259.950 850.050 262.050 ;
        RECT 850.950 260.100 853.050 262.200 ;
        RECT 857.400 262.050 858.450 295.950 ;
        RECT 851.400 259.350 852.600 260.100 ;
        RECT 856.950 259.950 859.050 262.050 ;
        RECT 850.950 256.950 853.050 259.050 ;
        RECT 853.950 256.950 856.050 259.050 ;
        RECT 839.400 254.400 846.450 255.450 ;
        RECT 833.400 252.450 834.450 254.400 ;
        RECT 830.400 251.400 834.450 252.450 ;
        RECT 823.950 247.950 826.050 250.050 ;
        RECT 814.950 238.950 817.050 241.050 ;
        RECT 802.950 235.950 805.050 238.050 ;
        RECT 811.950 235.950 814.050 238.050 ;
        RECT 808.950 217.950 811.050 220.050 ;
        RECT 793.950 215.100 796.050 217.200 ;
        RECT 803.400 216.450 804.600 216.600 ;
        RECT 803.400 215.400 807.450 216.450 ;
        RECT 794.400 214.350 795.600 215.100 ;
        RECT 803.400 214.350 804.600 215.400 ;
        RECT 794.100 211.950 796.200 214.050 ;
        RECT 799.500 211.950 801.600 214.050 ;
        RECT 802.800 211.950 804.900 214.050 ;
        RECT 806.400 210.900 807.450 215.400 ;
        RECT 805.950 208.800 808.050 210.900 ;
        RECT 809.400 208.050 810.450 217.950 ;
        RECT 815.400 217.200 816.450 238.950 ;
        RECT 830.400 232.050 831.450 251.400 ;
        RECT 832.950 232.950 835.050 235.050 ;
        RECT 829.950 229.950 832.050 232.050 ;
        RECT 829.950 223.950 832.050 226.050 ;
        RECT 820.800 220.950 822.900 223.050 ;
        RECT 814.950 215.100 817.050 217.200 ;
        RECT 821.400 216.600 822.450 220.950 ;
        RECT 815.400 214.350 816.600 215.100 ;
        RECT 821.400 214.350 822.600 216.600 ;
        RECT 814.950 211.950 817.050 214.050 ;
        RECT 817.950 211.950 820.050 214.050 ;
        RECT 820.950 211.950 823.050 214.050 ;
        RECT 823.950 211.950 826.050 214.050 ;
        RECT 818.400 210.900 819.600 211.650 ;
        RECT 817.950 208.800 820.050 210.900 ;
        RECT 824.400 209.400 825.600 211.650 ;
        RECT 808.950 205.950 811.050 208.050 ;
        RECT 817.950 205.650 820.050 207.750 ;
        RECT 805.950 202.950 808.050 205.050 ;
        RECT 814.950 202.950 817.050 205.050 ;
        RECT 790.950 199.950 793.050 202.050 ;
        RECT 796.950 199.950 799.050 202.050 ;
        RECT 781.950 183.450 784.050 187.050 ;
        RECT 785.400 183.450 786.600 183.600 ;
        RECT 781.950 183.000 786.600 183.450 ;
        RECT 782.400 182.400 786.600 183.000 ;
        RECT 785.400 181.350 786.600 182.400 ;
        RECT 790.950 182.100 793.050 184.200 ;
        RECT 791.400 181.350 792.600 182.100 ;
        RECT 784.950 178.950 787.050 181.050 ;
        RECT 787.950 178.950 790.050 181.050 ;
        RECT 790.950 178.950 793.050 181.050 ;
        RECT 781.950 175.950 784.050 178.050 ;
        RECT 788.400 176.400 789.600 178.650 ;
        RECT 782.400 172.050 783.450 175.950 ;
        RECT 788.400 172.050 789.450 176.400 ;
        RECT 781.950 169.950 784.050 172.050 ;
        RECT 787.950 169.950 790.050 172.050 ;
        RECT 797.400 166.050 798.450 199.950 ;
        RECT 799.950 187.950 802.050 190.050 ;
        RECT 800.400 184.050 801.450 187.950 ;
        RECT 799.950 181.950 802.050 184.050 ;
        RECT 806.400 183.600 807.450 202.950 ;
        RECT 806.400 181.350 807.600 183.600 ;
        RECT 811.950 182.100 814.050 184.200 ;
        RECT 815.400 184.050 816.450 202.950 ;
        RECT 812.400 181.350 813.600 182.100 ;
        RECT 814.950 181.950 817.050 184.050 ;
        RECT 802.950 178.950 805.050 181.050 ;
        RECT 805.950 178.950 808.050 181.050 ;
        RECT 808.950 178.950 811.050 181.050 ;
        RECT 811.950 178.950 814.050 181.050 ;
        RECT 803.400 177.900 804.600 178.650 ;
        RECT 802.950 175.800 805.050 177.900 ;
        RECT 809.400 176.400 810.600 178.650 ;
        RECT 796.950 163.950 799.050 166.050 ;
        RECT 803.400 163.050 804.450 175.800 ;
        RECT 787.950 160.950 790.050 163.050 ;
        RECT 802.950 160.950 805.050 163.050 ;
        RECT 778.950 154.950 781.050 157.050 ;
        RECT 784.950 148.950 787.050 151.050 ;
        RECT 748.950 133.950 751.050 136.050 ;
        RECT 751.950 133.950 754.050 136.050 ;
        RECT 754.950 133.950 757.050 136.050 ;
        RECT 757.950 133.950 760.050 136.050 ;
        RECT 749.400 132.900 750.600 133.650 ;
        RECT 755.400 132.900 756.600 133.650 ;
        RECT 748.950 130.800 751.050 132.900 ;
        RECT 754.950 130.800 757.050 132.900 ;
        RECT 764.400 132.450 765.450 137.100 ;
        RECT 770.400 136.350 771.600 137.100 ;
        RECT 776.400 136.350 777.600 138.600 ;
        RECT 769.950 133.950 772.050 136.050 ;
        RECT 772.950 133.950 775.050 136.050 ;
        RECT 775.950 133.950 778.050 136.050 ;
        RECT 778.950 133.950 781.050 136.050 ;
        RECT 761.400 131.400 765.450 132.450 ;
        RECT 745.950 129.450 748.050 130.050 ;
        RECT 751.950 129.450 754.050 130.050 ;
        RECT 745.950 128.400 754.050 129.450 ;
        RECT 745.950 127.950 748.050 128.400 ;
        RECT 751.950 127.950 754.050 128.400 ;
        RECT 761.400 112.050 762.450 131.400 ;
        RECT 766.950 130.950 769.050 133.050 ;
        RECT 773.400 132.000 774.600 133.650 ;
        RECT 767.400 115.050 768.450 130.950 ;
        RECT 772.950 127.950 775.050 132.000 ;
        RECT 779.400 131.400 780.600 133.650 ;
        RECT 772.950 121.950 775.050 124.050 ;
        RECT 766.800 112.950 768.900 115.050 ;
        RECT 769.950 112.950 772.050 115.050 ;
        RECT 760.950 109.950 763.050 112.050 ;
        RECT 736.950 104.100 739.050 106.200 ;
        RECT 742.950 104.100 745.050 106.200 ;
        RECT 737.400 103.350 738.600 104.100 ;
        RECT 743.400 103.350 744.600 104.100 ;
        RECT 748.950 103.950 751.050 106.050 ;
        RECT 757.950 104.100 760.050 106.200 ;
        RECT 763.950 105.000 766.050 109.050 ;
        RECT 733.950 100.950 736.050 103.050 ;
        RECT 736.950 100.950 739.050 103.050 ;
        RECT 739.950 100.950 742.050 103.050 ;
        RECT 742.950 100.950 745.050 103.050 ;
        RECT 734.400 98.400 735.600 100.650 ;
        RECT 740.400 99.900 741.600 100.650 ;
        RECT 727.950 88.950 730.050 91.050 ;
        RECT 734.400 88.050 735.450 98.400 ;
        RECT 739.950 97.800 742.050 99.900 ;
        RECT 736.950 91.950 739.050 94.050 ;
        RECT 715.950 85.950 718.050 88.050 ;
        RECT 733.950 85.950 736.050 88.050 ;
        RECT 737.400 85.050 738.450 91.950 ;
        RECT 736.950 82.950 739.050 85.050 ;
        RECT 742.950 79.950 745.050 82.050 ;
        RECT 721.950 64.950 724.050 67.050 ;
        RECT 701.400 58.350 702.600 60.000 ;
        RECT 706.950 59.100 709.050 61.200 ;
        RECT 712.950 60.450 715.050 61.200 ;
        RECT 722.400 60.600 723.450 64.950 ;
        RECT 712.950 59.400 717.450 60.450 ;
        RECT 712.950 59.100 715.050 59.400 ;
        RECT 707.400 58.350 708.600 59.100 ;
        RECT 700.950 55.950 703.050 58.050 ;
        RECT 703.950 55.950 706.050 58.050 ;
        RECT 706.950 55.950 709.050 58.050 ;
        RECT 709.950 55.950 712.050 58.050 ;
        RECT 704.400 54.900 705.600 55.650 ;
        RECT 703.950 52.800 706.050 54.900 ;
        RECT 710.400 53.400 711.600 55.650 ;
        RECT 703.950 43.950 706.050 46.050 ;
        RECT 700.950 37.950 703.050 40.050 ;
        RECT 701.400 28.050 702.450 37.950 ;
        RECT 704.400 34.050 705.450 43.950 ;
        RECT 710.400 40.050 711.450 53.400 ;
        RECT 716.400 40.050 717.450 59.400 ;
        RECT 722.400 58.350 723.600 60.600 ;
        RECT 727.950 59.100 730.050 61.200 ;
        RECT 733.950 59.100 736.050 61.200 ;
        RECT 743.400 60.600 744.450 79.950 ;
        RECT 728.400 58.350 729.600 59.100 ;
        RECT 721.950 55.950 724.050 58.050 ;
        RECT 724.950 55.950 727.050 58.050 ;
        RECT 727.950 55.950 730.050 58.050 ;
        RECT 725.400 54.900 726.600 55.650 ;
        RECT 734.400 55.050 735.450 59.100 ;
        RECT 743.400 58.350 744.600 60.600 ;
        RECT 739.950 55.950 742.050 58.050 ;
        RECT 742.950 55.950 745.050 58.050 ;
        RECT 724.950 52.800 727.050 54.900 ;
        RECT 733.950 52.950 736.050 55.050 ;
        RECT 740.400 54.900 741.600 55.650 ;
        RECT 749.400 54.900 750.450 103.950 ;
        RECT 758.400 103.350 759.600 104.100 ;
        RECT 764.400 103.350 765.600 105.000 ;
        RECT 754.950 100.950 757.050 103.050 ;
        RECT 757.950 100.950 760.050 103.050 ;
        RECT 760.950 100.950 763.050 103.050 ;
        RECT 763.950 100.950 766.050 103.050 ;
        RECT 755.400 99.450 756.600 100.650 ;
        RECT 761.400 99.900 762.600 100.650 ;
        RECT 770.400 99.900 771.450 112.950 ;
        RECT 773.400 106.050 774.450 121.950 ;
        RECT 779.400 115.050 780.450 131.400 ;
        RECT 785.400 124.050 786.450 148.950 ;
        RECT 788.400 139.050 789.450 160.950 ;
        RECT 809.400 160.050 810.450 176.400 ;
        RECT 814.950 175.950 817.050 178.050 ;
        RECT 815.400 172.050 816.450 175.950 ;
        RECT 814.950 169.950 817.050 172.050 ;
        RECT 808.950 157.950 811.050 160.050 ;
        RECT 815.400 157.050 816.450 169.950 ;
        RECT 818.400 169.050 819.450 205.650 ;
        RECT 824.400 201.450 825.450 209.400 ;
        RECT 826.950 208.950 829.050 211.050 ;
        RECT 827.400 205.050 828.450 208.950 ;
        RECT 826.950 202.950 829.050 205.050 ;
        RECT 824.400 200.400 828.450 201.450 ;
        RECT 823.950 196.950 826.050 199.050 ;
        RECT 820.950 184.950 823.050 187.050 ;
        RECT 817.950 166.950 820.050 169.050 ;
        RECT 802.950 154.950 805.050 157.050 ;
        RECT 814.950 154.950 817.050 157.050 ;
        RECT 796.950 142.950 799.050 145.050 ;
        RECT 797.400 139.200 798.450 142.950 ;
        RECT 787.950 136.950 790.050 139.050 ;
        RECT 790.950 137.100 793.050 139.200 ;
        RECT 796.950 137.100 799.050 139.200 ;
        RECT 791.400 136.350 792.600 137.100 ;
        RECT 797.400 136.350 798.600 137.100 ;
        RECT 790.950 133.950 793.050 136.050 ;
        RECT 793.950 133.950 796.050 136.050 ;
        RECT 796.950 133.950 799.050 136.050 ;
        RECT 787.950 130.950 790.050 133.050 ;
        RECT 794.400 131.400 795.600 133.650 ;
        RECT 784.950 121.950 787.050 124.050 ;
        RECT 778.950 112.950 781.050 115.050 ;
        RECT 772.950 103.950 775.050 106.050 ;
        RECT 775.950 105.000 778.050 109.050 ;
        RECT 776.400 103.350 777.600 105.000 ;
        RECT 781.950 104.100 784.050 106.200 ;
        RECT 788.400 105.450 789.450 130.950 ;
        RECT 794.400 121.050 795.450 131.400 ;
        RECT 799.950 130.950 802.050 133.050 ;
        RECT 793.950 118.950 796.050 121.050 ;
        RECT 791.400 113.400 798.450 114.450 ;
        RECT 791.400 109.050 792.450 113.400 ;
        RECT 793.950 109.950 796.050 112.050 ;
        RECT 790.950 106.950 793.050 109.050 ;
        RECT 794.400 106.050 795.450 109.950 ;
        RECT 788.400 104.400 792.450 105.450 ;
        RECT 782.400 103.350 783.600 104.100 ;
        RECT 775.950 100.950 778.050 103.050 ;
        RECT 778.950 100.950 781.050 103.050 ;
        RECT 781.950 100.950 784.050 103.050 ;
        RECT 784.950 100.950 787.050 103.050 ;
        RECT 752.400 98.400 756.600 99.450 ;
        RECT 739.950 52.800 742.050 54.900 ;
        RECT 748.950 52.800 751.050 54.900 ;
        RECT 718.950 43.950 721.050 46.050 ;
        RECT 709.950 37.950 712.050 40.050 ;
        RECT 715.950 37.950 718.050 40.050 ;
        RECT 719.400 37.050 720.450 43.950 ;
        RECT 730.950 37.950 733.050 40.050 ;
        RECT 718.950 34.950 721.050 37.050 ;
        RECT 703.950 31.950 706.050 34.050 ;
        RECT 709.950 31.950 712.050 34.050 ;
        RECT 695.400 26.400 699.450 27.450 ;
        RECT 686.400 25.350 687.600 26.100 ;
        RECT 692.400 25.350 693.600 26.100 ;
        RECT 682.950 22.950 685.050 25.050 ;
        RECT 685.950 22.950 688.050 25.050 ;
        RECT 688.950 22.950 691.050 25.050 ;
        RECT 691.950 22.950 694.050 25.050 ;
        RECT 683.400 21.900 684.600 22.650 ;
        RECT 613.950 13.950 616.050 16.050 ;
        RECT 655.950 13.950 658.050 16.050 ;
        RECT 667.950 13.950 670.050 16.050 ;
        RECT 610.950 10.950 613.050 13.050 ;
        RECT 674.400 4.050 675.450 19.950 ;
        RECT 676.950 19.800 679.050 21.900 ;
        RECT 682.950 19.800 685.050 21.900 ;
        RECT 689.400 21.000 690.600 22.650 ;
        RECT 688.950 13.950 691.050 21.000 ;
        RECT 698.400 13.050 699.450 26.400 ;
        RECT 700.950 25.950 703.050 28.050 ;
        RECT 703.950 26.100 706.050 28.200 ;
        RECT 710.400 27.600 711.450 31.950 ;
        RECT 704.400 25.350 705.600 26.100 ;
        RECT 710.400 25.350 711.600 27.600 ;
        RECT 703.950 22.950 706.050 25.050 ;
        RECT 706.950 22.950 709.050 25.050 ;
        RECT 709.950 22.950 712.050 25.050 ;
        RECT 712.950 22.950 715.050 25.050 ;
        RECT 707.400 21.000 708.600 22.650 ;
        RECT 713.400 21.900 714.600 22.650 ;
        RECT 719.400 21.900 720.450 34.950 ;
        RECT 731.400 27.600 732.450 37.950 ;
        RECT 740.400 36.450 741.450 52.800 ;
        RECT 752.400 49.050 753.450 98.400 ;
        RECT 760.950 97.800 763.050 99.900 ;
        RECT 769.950 97.800 772.050 99.900 ;
        RECT 772.950 97.950 775.050 100.050 ;
        RECT 779.400 99.900 780.600 100.650 ;
        RECT 757.950 59.100 760.050 61.200 ;
        RECT 763.950 59.100 766.050 61.200 ;
        RECT 769.950 59.100 772.050 64.050 ;
        RECT 758.400 58.350 759.600 59.100 ;
        RECT 764.400 58.350 765.600 59.100 ;
        RECT 757.950 55.950 760.050 58.050 ;
        RECT 760.950 55.950 763.050 58.050 ;
        RECT 763.950 55.950 766.050 58.050 ;
        RECT 766.950 55.950 769.050 58.050 ;
        RECT 761.400 54.900 762.600 55.650 ;
        RECT 760.950 52.800 763.050 54.900 ;
        RECT 767.400 54.000 768.600 55.650 ;
        RECT 766.950 49.950 769.050 54.000 ;
        RECT 769.950 52.950 772.050 55.050 ;
        RECT 751.950 46.950 754.050 49.050 ;
        RECT 745.950 40.950 748.050 43.050 ;
        RECT 737.400 35.400 741.450 36.450 ;
        RECT 731.400 25.350 732.600 27.600 ;
        RECT 725.100 22.950 727.200 25.050 ;
        RECT 730.500 22.950 732.600 25.050 ;
        RECT 733.800 22.950 735.900 25.050 ;
        RECT 706.950 16.950 709.050 21.000 ;
        RECT 712.950 19.800 715.050 21.900 ;
        RECT 718.950 19.800 721.050 21.900 ;
        RECT 725.400 20.400 726.600 22.650 ;
        RECT 734.400 21.000 735.600 22.650 ;
        RECT 725.400 13.050 726.450 20.400 ;
        RECT 733.950 16.950 736.050 21.000 ;
        RECT 697.950 10.950 700.050 13.050 ;
        RECT 724.950 10.950 727.050 13.050 ;
        RECT 737.400 7.050 738.450 35.400 ;
        RECT 746.400 27.600 747.450 40.950 ;
        RECT 770.400 37.050 771.450 52.950 ;
        RECT 757.950 34.950 760.050 37.050 ;
        RECT 769.950 34.950 772.050 37.050 ;
        RECT 758.400 31.050 759.450 34.950 ;
        RECT 760.950 31.950 763.050 34.050 ;
        RECT 746.400 25.350 747.600 27.600 ;
        RECT 751.950 26.100 754.050 28.200 ;
        RECT 752.400 25.350 753.600 26.100 ;
        RECT 757.950 25.950 760.050 31.050 ;
        RECT 739.950 22.950 742.050 25.050 ;
        RECT 745.950 22.950 748.050 25.050 ;
        RECT 748.950 22.950 751.050 25.050 ;
        RECT 751.950 22.950 754.050 25.050 ;
        RECT 754.950 22.950 757.050 25.050 ;
        RECT 740.400 19.050 741.450 22.950 ;
        RECT 749.400 21.900 750.600 22.650 ;
        RECT 748.950 19.800 751.050 21.900 ;
        RECT 755.400 20.400 756.600 22.650 ;
        RECT 739.950 16.950 742.050 19.050 ;
        RECT 747.000 18.750 750.000 19.050 ;
        RECT 745.950 16.950 751.050 18.750 ;
        RECT 745.950 16.650 748.050 16.950 ;
        RECT 748.950 16.650 751.050 16.950 ;
        RECT 755.400 16.050 756.450 20.400 ;
        RECT 761.400 16.050 762.450 31.950 ;
        RECT 773.400 31.050 774.450 97.950 ;
        RECT 778.950 97.800 781.050 99.900 ;
        RECT 785.400 98.400 786.600 100.650 ;
        RECT 781.950 76.950 784.050 79.050 ;
        RECT 782.400 60.600 783.450 76.950 ;
        RECT 785.400 70.050 786.450 98.400 ;
        RECT 791.400 97.050 792.450 104.400 ;
        RECT 793.950 103.950 796.050 106.050 ;
        RECT 797.400 105.600 798.450 113.400 ;
        RECT 800.400 109.050 801.450 130.950 ;
        RECT 803.400 115.050 804.450 154.950 ;
        RECT 805.950 145.950 808.050 148.050 ;
        RECT 806.400 139.050 807.450 145.950 ;
        RECT 821.400 142.050 822.450 184.950 ;
        RECT 824.400 183.450 825.450 196.950 ;
        RECT 827.400 193.050 828.450 200.400 ;
        RECT 830.400 196.050 831.450 223.950 ;
        RECT 833.400 217.050 834.450 232.950 ;
        RECT 832.950 214.950 835.050 217.050 ;
        RECT 835.950 215.100 838.050 217.200 ;
        RECT 842.400 216.600 843.450 254.400 ;
        RECT 847.950 250.950 850.050 256.050 ;
        RECT 854.400 255.000 855.600 256.650 ;
        RECT 853.950 250.950 856.050 255.000 ;
        RECT 856.950 253.950 859.050 256.050 ;
        RECT 853.950 220.950 856.050 223.050 ;
        RECT 836.400 214.350 837.600 215.100 ;
        RECT 842.400 214.350 843.600 216.600 ;
        RECT 847.950 215.100 850.050 217.200 ;
        RECT 848.400 214.350 849.600 215.100 ;
        RECT 835.950 211.950 838.050 214.050 ;
        RECT 838.950 211.950 841.050 214.050 ;
        RECT 841.950 211.950 844.050 214.050 ;
        RECT 844.950 211.950 847.050 214.050 ;
        RECT 847.950 211.950 850.050 214.050 ;
        RECT 839.400 210.900 840.600 211.650 ;
        RECT 838.950 208.800 841.050 210.900 ;
        RECT 845.400 209.400 846.600 211.650 ;
        RECT 854.400 210.900 855.450 220.950 ;
        RECT 857.400 216.450 858.450 253.950 ;
        RECT 860.400 226.050 861.450 343.950 ;
        RECT 869.400 343.050 870.450 424.950 ;
        RECT 872.400 412.050 873.450 449.100 ;
        RECT 871.950 409.950 874.050 412.050 ;
        RECT 875.400 396.450 876.450 643.950 ;
        RECT 872.400 395.400 876.450 396.450 ;
        RECT 868.950 340.950 871.050 343.050 ;
        RECT 862.950 338.100 865.050 340.200 ;
        RECT 863.400 337.350 864.600 338.100 ;
        RECT 863.400 334.950 865.500 337.050 ;
        RECT 868.800 334.950 870.900 337.050 ;
        RECT 862.950 328.950 865.050 331.050 ;
        RECT 863.400 325.050 864.450 328.950 ;
        RECT 862.950 322.950 865.050 325.050 ;
        RECT 872.400 298.050 873.450 395.400 ;
        RECT 874.950 340.950 877.050 343.050 ;
        RECT 862.950 295.950 865.050 298.050 ;
        RECT 871.950 295.950 874.050 298.050 ;
        RECT 859.950 223.950 862.050 226.050 ;
        RECT 863.400 220.050 864.450 295.950 ;
        RECT 868.950 289.950 871.050 292.050 ;
        RECT 865.950 265.950 868.050 268.050 ;
        RECT 866.400 223.050 867.450 265.950 ;
        RECT 869.400 235.050 870.450 289.950 ;
        RECT 871.950 277.950 874.050 280.050 ;
        RECT 868.950 232.950 871.050 235.050 ;
        RECT 865.950 220.950 868.050 223.050 ;
        RECT 862.950 217.950 865.050 220.050 ;
        RECT 860.400 216.450 861.600 216.600 ;
        RECT 857.400 215.400 861.600 216.450 ;
        RECT 860.400 214.350 861.600 215.400 ;
        RECT 865.950 215.100 868.050 217.200 ;
        RECT 872.400 217.050 873.450 277.950 ;
        RECT 866.400 214.350 867.600 215.100 ;
        RECT 871.950 214.950 874.050 217.050 ;
        RECT 859.950 211.950 862.050 214.050 ;
        RECT 862.950 211.950 865.050 214.050 ;
        RECT 865.950 211.950 868.050 214.050 ;
        RECT 868.950 211.950 871.050 214.050 ;
        RECT 845.400 199.050 846.450 209.400 ;
        RECT 853.950 208.800 856.050 210.900 ;
        RECT 856.950 208.950 859.050 211.050 ;
        RECT 863.400 210.900 864.600 211.650 ;
        RECT 869.400 210.900 870.600 211.650 ;
        RECT 847.950 205.950 850.050 208.050 ;
        RECT 844.950 196.950 847.050 199.050 ;
        RECT 829.950 193.950 832.050 196.050 ;
        RECT 841.950 193.950 844.050 196.050 ;
        RECT 826.950 190.950 829.050 193.050 ;
        RECT 829.800 186.300 831.900 188.400 ;
        RECT 832.950 187.950 835.050 190.050 ;
        RECT 833.400 187.200 834.600 187.950 ;
        RECT 842.400 187.050 843.450 193.950 ;
        RECT 844.950 192.450 847.050 193.050 ;
        RECT 848.400 192.450 849.450 205.950 ;
        RECT 850.950 196.950 853.050 199.050 ;
        RECT 844.950 191.400 849.450 192.450 ;
        RECT 844.950 190.950 847.050 191.400 ;
        RECT 827.400 183.450 828.600 183.600 ;
        RECT 824.400 182.400 828.600 183.450 ;
        RECT 827.400 181.350 828.600 182.400 ;
        RECT 823.950 178.950 826.050 181.050 ;
        RECT 827.100 178.950 829.200 181.050 ;
        RECT 830.100 180.900 831.000 186.300 ;
        RECT 833.100 184.800 835.200 186.900 ;
        RECT 837.000 183.900 839.100 185.700 ;
        RECT 841.950 184.950 844.050 187.050 ;
        RECT 831.900 182.700 840.600 183.900 ;
        RECT 831.900 181.800 834.000 182.700 ;
        RECT 830.100 179.700 837.000 180.900 ;
        RECT 824.400 148.050 825.450 178.950 ;
        RECT 830.100 172.500 831.300 179.700 ;
        RECT 833.100 175.950 835.200 178.050 ;
        RECT 836.100 177.300 837.000 179.700 ;
        RECT 833.400 173.400 834.600 175.650 ;
        RECT 836.100 175.200 838.200 177.300 ;
        RECT 839.700 173.700 840.600 182.700 ;
        RECT 841.800 178.950 843.900 181.050 ;
        RECT 842.400 177.450 843.600 178.650 ;
        RECT 845.400 177.450 846.450 190.950 ;
        RECT 847.950 184.950 850.050 187.050 ;
        RECT 842.400 176.400 846.450 177.450 ;
        RECT 829.800 170.400 831.900 172.500 ;
        RECT 839.400 171.600 841.500 173.700 ;
        RECT 838.950 163.950 841.050 166.050 ;
        RECT 823.950 145.950 826.050 148.050 ;
        RECT 813.000 141.450 817.050 142.050 ;
        RECT 812.400 139.950 817.050 141.450 ;
        RECT 820.950 139.950 823.050 142.050 ;
        RECT 805.950 136.950 808.050 139.050 ;
        RECT 812.400 138.600 813.450 139.950 ;
        RECT 812.400 136.350 813.600 138.600 ;
        RECT 808.950 133.950 811.050 136.050 ;
        RECT 811.950 133.950 814.050 136.050 ;
        RECT 814.950 133.950 817.050 136.050 ;
        RECT 809.400 132.900 810.600 133.650 ;
        RECT 815.400 132.900 816.600 133.650 ;
        RECT 808.950 130.800 811.050 132.900 ;
        RECT 814.950 130.800 817.050 132.900 ;
        RECT 809.400 127.050 810.450 130.800 ;
        RECT 808.950 124.950 811.050 127.050 ;
        RECT 805.950 118.950 808.050 121.050 ;
        RECT 802.950 112.950 805.050 115.050 ;
        RECT 799.950 106.950 802.050 109.050 ;
        RECT 806.400 108.450 807.450 118.950 ;
        RECT 808.950 115.950 811.050 118.050 ;
        RECT 803.400 107.400 807.450 108.450 ;
        RECT 803.400 105.600 804.450 107.400 ;
        RECT 809.400 106.050 810.450 115.950 ;
        RECT 811.800 106.950 813.900 109.050 ;
        RECT 797.400 103.350 798.600 105.600 ;
        RECT 803.400 103.350 804.600 105.600 ;
        RECT 808.950 103.950 811.050 106.050 ;
        RECT 796.950 100.950 799.050 103.050 ;
        RECT 799.950 100.950 802.050 103.050 ;
        RECT 802.950 100.950 805.050 103.050 ;
        RECT 805.950 100.950 808.050 103.050 ;
        RECT 800.400 99.000 801.600 100.650 ;
        RECT 806.400 99.000 807.600 100.650 ;
        RECT 790.950 94.950 793.050 97.050 ;
        RECT 799.950 94.950 802.050 99.000 ;
        RECT 805.950 94.950 808.050 99.000 ;
        RECT 806.400 91.050 807.450 94.950 ;
        RECT 787.950 88.950 790.050 91.050 ;
        RECT 805.950 88.950 808.050 91.050 ;
        RECT 784.950 67.950 787.050 70.050 ;
        RECT 785.400 64.050 786.450 67.950 ;
        RECT 784.950 61.950 787.050 64.050 ;
        RECT 788.400 61.200 789.450 88.950 ;
        RECT 793.950 82.950 796.050 85.050 ;
        RECT 782.400 58.350 783.600 60.600 ;
        RECT 787.950 59.100 790.050 61.200 ;
        RECT 788.400 58.350 789.600 59.100 ;
        RECT 778.950 55.950 781.050 58.050 ;
        RECT 781.950 55.950 784.050 58.050 ;
        RECT 784.950 55.950 787.050 58.050 ;
        RECT 787.950 55.950 790.050 58.050 ;
        RECT 779.400 54.900 780.600 55.650 ;
        RECT 785.400 54.900 786.600 55.650 ;
        RECT 778.950 52.800 781.050 54.900 ;
        RECT 784.950 52.800 787.050 54.900 ;
        RECT 790.950 52.950 793.050 55.050 ;
        RECT 775.950 46.950 778.050 49.050 ;
        RECT 769.950 27.000 772.050 31.050 ;
        RECT 772.950 28.950 775.050 31.050 ;
        RECT 776.400 27.600 777.450 46.950 ;
        RECT 791.400 28.200 792.450 52.950 ;
        RECT 794.400 52.050 795.450 82.950 ;
        RECT 796.950 64.950 799.050 67.050 ;
        RECT 797.400 61.050 798.450 64.950 ;
        RECT 796.950 58.950 799.050 61.050 ;
        RECT 802.950 59.100 805.050 61.200 ;
        RECT 808.950 59.100 811.050 61.200 ;
        RECT 812.400 60.450 813.450 106.950 ;
        RECT 814.950 103.950 817.050 109.050 ;
        RECT 821.400 106.200 822.450 139.950 ;
        RECT 823.950 137.100 826.050 142.050 ;
        RECT 829.950 137.100 832.050 142.050 ;
        RECT 835.950 138.000 838.050 142.050 ;
        RECT 839.400 139.050 840.450 163.950 ;
        RECT 844.950 154.950 847.050 157.050 ;
        RECT 841.950 151.950 844.050 154.050 ;
        RECT 830.400 136.350 831.600 137.100 ;
        RECT 836.400 136.350 837.600 138.000 ;
        RECT 838.950 136.950 841.050 139.050 ;
        RECT 826.950 133.950 829.050 136.050 ;
        RECT 829.950 133.950 832.050 136.050 ;
        RECT 832.950 133.950 835.050 136.050 ;
        RECT 835.950 133.950 838.050 136.050 ;
        RECT 827.400 131.400 828.600 133.650 ;
        RECT 833.400 131.400 834.600 133.650 ;
        RECT 823.950 115.950 826.050 118.050 ;
        RECT 824.400 109.050 825.450 115.950 ;
        RECT 827.400 115.050 828.450 131.400 ;
        RECT 833.400 121.050 834.450 131.400 ;
        RECT 838.950 130.950 841.050 133.050 ;
        RECT 839.400 127.050 840.450 130.950 ;
        RECT 838.950 124.950 841.050 127.050 ;
        RECT 832.950 120.450 835.050 121.050 ;
        RECT 830.400 119.400 835.050 120.450 ;
        RECT 826.950 112.950 829.050 115.050 ;
        RECT 823.950 106.950 826.050 109.050 ;
        RECT 820.950 104.100 823.050 106.200 ;
        RECT 826.950 104.100 829.050 106.200 ;
        RECT 830.400 106.050 831.450 119.400 ;
        RECT 832.950 118.950 835.050 119.400 ;
        RECT 842.400 118.050 843.450 151.950 ;
        RECT 845.400 139.050 846.450 154.950 ;
        RECT 848.400 148.050 849.450 184.950 ;
        RECT 851.400 183.450 852.450 196.950 ;
        RECT 857.400 196.050 858.450 208.950 ;
        RECT 862.950 208.800 865.050 210.900 ;
        RECT 868.950 208.800 871.050 210.900 ;
        RECT 856.950 193.950 859.050 196.050 ;
        RECT 862.950 193.950 865.050 196.050 ;
        RECT 859.950 187.950 862.050 190.050 ;
        RECT 860.400 187.200 861.600 187.950 ;
        RECT 856.500 185.100 858.600 187.200 ;
        RECT 863.400 187.050 864.450 193.950 ;
        RECT 871.950 190.950 874.050 193.050 ;
        RECT 854.400 183.450 855.600 183.600 ;
        RECT 851.400 182.400 855.600 183.450 ;
        RECT 854.400 181.350 855.600 182.400 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 854.100 178.950 856.200 181.050 ;
        RECT 857.100 180.000 858.000 185.100 ;
        RECT 859.800 184.800 861.900 186.900 ;
        RECT 862.950 184.950 865.050 187.050 ;
        RECT 866.400 185.400 868.500 187.500 ;
        RECT 864.000 183.000 866.100 183.900 ;
        RECT 858.900 181.800 866.100 183.000 ;
        RECT 858.900 180.900 861.000 181.800 ;
        RECT 864.000 180.000 866.100 180.900 ;
        RECT 857.100 179.100 866.100 180.000 ;
        RECT 851.400 160.050 852.450 178.950 ;
        RECT 857.100 172.500 858.000 179.100 ;
        RECT 864.000 178.800 866.100 179.100 ;
        RECT 859.800 175.950 861.900 178.050 ;
        RECT 860.400 173.400 861.600 175.650 ;
        RECT 867.000 172.800 867.900 185.400 ;
        RECT 868.800 178.950 870.900 181.050 ;
        RECT 869.400 177.450 870.600 178.650 ;
        RECT 872.400 177.450 873.450 190.950 ;
        RECT 869.400 176.400 873.450 177.450 ;
        RECT 875.400 174.450 876.450 340.950 ;
        RECT 872.400 173.400 876.450 174.450 ;
        RECT 857.100 170.400 859.200 172.500 ;
        RECT 866.100 170.700 868.200 172.800 ;
        RECT 868.950 166.950 871.050 169.050 ;
        RECT 850.950 157.950 853.050 160.050 ;
        RECT 847.950 145.950 850.050 148.050 ;
        RECT 851.400 145.050 852.450 157.950 ;
        RECT 862.950 145.950 865.050 148.050 ;
        RECT 850.950 142.950 853.050 145.050 ;
        RECT 856.950 142.950 859.050 145.050 ;
        RECT 844.950 136.950 847.050 139.050 ;
        RECT 850.950 138.000 853.050 141.900 ;
        RECT 857.400 138.600 858.450 142.950 ;
        RECT 851.400 136.350 852.600 138.000 ;
        RECT 857.400 136.350 858.600 138.600 ;
        RECT 847.950 133.950 850.050 136.050 ;
        RECT 850.950 133.950 853.050 136.050 ;
        RECT 853.950 133.950 856.050 136.050 ;
        RECT 856.950 133.950 859.050 136.050 ;
        RECT 848.400 132.900 849.600 133.650 ;
        RECT 847.950 130.800 850.050 132.900 ;
        RECT 854.400 131.400 855.600 133.650 ;
        RECT 850.950 124.950 853.050 127.050 ;
        RECT 844.950 118.950 847.050 121.050 ;
        RECT 835.950 115.950 838.050 118.050 ;
        RECT 841.950 115.950 844.050 118.050 ;
        RECT 821.400 103.350 822.600 104.100 ;
        RECT 827.400 103.350 828.600 104.100 ;
        RECT 829.950 103.950 832.050 106.050 ;
        RECT 836.400 105.450 837.450 115.950 ;
        RECT 833.400 104.400 837.450 105.450 ;
        RECT 838.950 105.000 841.050 109.050 ;
        RECT 845.400 106.200 846.450 118.950 ;
        RECT 851.400 117.450 852.450 124.950 ;
        RECT 854.400 121.050 855.450 131.400 ;
        RECT 853.950 118.950 856.050 121.050 ;
        RECT 851.400 116.400 855.450 117.450 ;
        RECT 817.950 100.950 820.050 103.050 ;
        RECT 820.950 100.950 823.050 103.050 ;
        RECT 823.950 100.950 826.050 103.050 ;
        RECT 826.950 100.950 829.050 103.050 ;
        RECT 814.950 97.950 817.050 100.050 ;
        RECT 818.400 98.400 819.600 100.650 ;
        RECT 824.400 98.400 825.600 100.650 ;
        RECT 815.400 64.050 816.450 97.950 ;
        RECT 818.400 94.050 819.450 98.400 ;
        RECT 820.950 94.950 823.050 97.050 ;
        RECT 817.950 91.950 820.050 94.050 ;
        RECT 814.950 61.950 817.050 64.050 ;
        RECT 821.400 60.600 822.450 94.950 ;
        RECT 824.400 91.050 825.450 98.400 ;
        RECT 829.950 97.950 832.050 100.050 ;
        RECT 830.400 94.050 831.450 97.950 ;
        RECT 829.950 91.950 832.050 94.050 ;
        RECT 823.950 88.950 826.050 91.050 ;
        RECT 833.400 67.050 834.450 104.400 ;
        RECT 839.400 103.350 840.600 105.000 ;
        RECT 844.950 104.100 847.050 106.200 ;
        RECT 845.400 103.350 846.600 104.100 ;
        RECT 838.950 100.950 841.050 103.050 ;
        RECT 841.950 100.950 844.050 103.050 ;
        RECT 844.950 100.950 847.050 103.050 ;
        RECT 847.950 100.950 850.050 103.050 ;
        RECT 842.400 98.400 843.600 100.650 ;
        RECT 848.400 99.000 849.600 100.650 ;
        RECT 835.950 91.950 838.050 94.050 ;
        RECT 832.950 64.950 835.050 67.050 ;
        RECT 812.400 59.400 816.450 60.450 ;
        RECT 803.400 58.350 804.600 59.100 ;
        RECT 809.400 58.350 810.600 59.100 ;
        RECT 799.950 55.950 802.050 58.050 ;
        RECT 802.950 55.950 805.050 58.050 ;
        RECT 805.950 55.950 808.050 58.050 ;
        RECT 808.950 55.950 811.050 58.050 ;
        RECT 796.950 52.950 799.050 55.050 ;
        RECT 800.400 54.000 801.600 55.650 ;
        RECT 806.400 54.000 807.600 55.650 ;
        RECT 793.950 49.950 796.050 52.050 ;
        RECT 797.400 34.050 798.450 52.950 ;
        RECT 799.950 49.950 802.050 54.000 ;
        RECT 805.950 49.950 808.050 54.000 ;
        RECT 811.950 52.950 814.050 55.050 ;
        RECT 806.400 40.050 807.450 49.950 ;
        RECT 805.950 37.950 808.050 40.050 ;
        RECT 812.400 37.050 813.450 52.950 ;
        RECT 811.950 34.950 814.050 37.050 ;
        RECT 796.950 31.950 799.050 34.050 ;
        RECT 802.950 31.950 805.050 34.050 ;
        RECT 796.950 28.800 799.050 30.900 ;
        RECT 770.400 25.350 771.600 27.000 ;
        RECT 776.400 25.350 777.600 27.600 ;
        RECT 781.950 25.950 784.050 28.050 ;
        RECT 790.950 26.100 793.050 28.200 ;
        RECT 766.950 22.950 769.050 25.050 ;
        RECT 769.950 22.950 772.050 25.050 ;
        RECT 772.950 22.950 775.050 25.050 ;
        RECT 775.950 22.950 778.050 25.050 ;
        RECT 767.400 21.000 768.600 22.650 ;
        RECT 773.400 21.900 774.600 22.650 ;
        RECT 766.950 16.950 769.050 21.000 ;
        RECT 772.950 19.800 775.050 21.900 ;
        RECT 782.400 16.050 783.450 25.950 ;
        RECT 791.400 25.350 792.600 26.100 ;
        RECT 787.950 22.950 790.050 25.050 ;
        RECT 790.950 22.950 793.050 25.050 ;
        RECT 788.400 21.900 789.600 22.650 ;
        RECT 797.400 22.050 798.450 28.800 ;
        RECT 803.400 27.600 804.450 31.950 ;
        RECT 815.400 28.200 816.450 59.400 ;
        RECT 821.400 58.350 822.600 60.600 ;
        RECT 826.950 59.100 829.050 61.200 ;
        RECT 827.400 58.350 828.600 59.100 ;
        RECT 820.950 55.950 823.050 58.050 ;
        RECT 823.950 55.950 826.050 58.050 ;
        RECT 826.950 55.950 829.050 58.050 ;
        RECT 829.950 55.950 832.050 58.050 ;
        RECT 817.950 52.950 820.050 55.050 ;
        RECT 824.400 53.400 825.600 55.650 ;
        RECT 830.400 53.400 831.600 55.650 ;
        RECT 818.400 43.050 819.450 52.950 ;
        RECT 824.400 49.050 825.450 53.400 ;
        RECT 823.950 46.950 826.050 49.050 ;
        RECT 817.950 40.950 820.050 43.050 ;
        RECT 826.950 37.950 829.050 40.050 ;
        RECT 820.950 31.950 823.050 34.050 ;
        RECT 803.400 25.350 804.600 27.600 ;
        RECT 808.950 26.100 811.050 28.200 ;
        RECT 814.950 26.100 817.050 28.200 ;
        RECT 821.400 27.600 822.450 31.950 ;
        RECT 827.400 27.600 828.450 37.950 ;
        RECT 830.400 37.050 831.450 53.400 ;
        RECT 836.400 49.050 837.450 91.950 ;
        RECT 842.400 70.050 843.450 98.400 ;
        RECT 847.950 94.950 850.050 99.000 ;
        RECT 850.950 97.950 853.050 100.050 ;
        RECT 841.950 67.950 844.050 70.050 ;
        RECT 844.950 67.950 847.050 70.050 ;
        RECT 845.400 60.600 846.450 67.950 ;
        RECT 848.400 64.050 849.450 94.950 ;
        RECT 847.950 61.950 850.050 64.050 ;
        RECT 851.400 61.200 852.450 97.950 ;
        RECT 854.400 94.050 855.450 116.400 ;
        RECT 863.400 105.600 864.450 145.950 ;
        RECT 863.400 103.350 864.600 105.600 ;
        RECT 859.950 100.950 862.050 103.050 ;
        RECT 862.950 100.950 865.050 103.050 ;
        RECT 860.400 99.900 861.600 100.650 ;
        RECT 869.400 100.050 870.450 166.950 ;
        RECT 859.950 97.800 862.050 99.900 ;
        RECT 868.950 97.950 871.050 100.050 ;
        RECT 853.950 91.950 856.050 94.050 ;
        RECT 856.950 85.950 859.050 88.050 ;
        RECT 845.400 58.350 846.600 60.600 ;
        RECT 850.950 59.100 853.050 61.200 ;
        RECT 851.400 58.350 852.600 59.100 ;
        RECT 841.950 55.950 844.050 58.050 ;
        RECT 844.950 55.950 847.050 58.050 ;
        RECT 847.950 55.950 850.050 58.050 ;
        RECT 850.950 55.950 853.050 58.050 ;
        RECT 842.400 54.900 843.600 55.650 ;
        RECT 848.400 54.900 849.600 55.650 ;
        RECT 841.950 52.800 844.050 54.900 ;
        RECT 847.950 52.800 850.050 54.900 ;
        RECT 835.950 46.950 838.050 49.050 ;
        RECT 838.950 43.950 841.050 46.050 ;
        RECT 835.950 40.950 838.050 43.050 ;
        RECT 829.950 36.450 832.050 37.050 ;
        RECT 829.950 35.400 834.450 36.450 ;
        RECT 829.950 34.950 832.050 35.400 ;
        RECT 833.400 28.050 834.450 35.400 ;
        RECT 809.400 25.350 810.600 26.100 ;
        RECT 821.400 25.350 822.600 27.600 ;
        RECT 827.400 25.350 828.600 27.600 ;
        RECT 832.950 25.950 835.050 28.050 ;
        RECT 836.400 27.450 837.450 40.950 ;
        RECT 839.400 31.050 840.450 43.950 ;
        RECT 838.950 28.950 841.050 31.050 ;
        RECT 848.400 27.600 849.450 52.800 ;
        RECT 850.950 49.950 853.050 52.050 ;
        RECT 851.400 31.050 852.450 49.950 ;
        RECT 853.950 34.950 856.050 37.050 ;
        RECT 850.950 28.950 853.050 31.050 ;
        RECT 842.400 27.450 843.600 27.600 ;
        RECT 836.400 26.400 843.600 27.450 ;
        RECT 802.950 22.950 805.050 25.050 ;
        RECT 805.950 22.950 808.050 25.050 ;
        RECT 808.950 22.950 811.050 25.050 ;
        RECT 820.950 22.950 823.050 25.050 ;
        RECT 823.950 22.950 826.050 25.050 ;
        RECT 826.950 22.950 829.050 25.050 ;
        RECT 829.950 22.950 832.050 25.050 ;
        RECT 787.950 19.800 790.050 21.900 ;
        RECT 796.950 19.950 799.050 22.050 ;
        RECT 806.400 21.900 807.600 22.650 ;
        RECT 805.950 19.800 808.050 21.900 ;
        RECT 824.400 21.000 825.600 22.650 ;
        RECT 830.400 21.900 831.600 22.650 ;
        RECT 823.950 16.950 826.050 21.000 ;
        RECT 829.950 19.800 832.050 21.900 ;
        RECT 836.400 19.050 837.450 26.400 ;
        RECT 842.400 25.350 843.600 26.400 ;
        RECT 848.400 25.350 849.600 27.600 ;
        RECT 854.400 27.450 855.450 34.950 ;
        RECT 857.400 31.050 858.450 85.950 ;
        RECT 872.400 64.050 873.450 173.400 ;
        RECT 874.950 169.950 877.050 172.050 ;
        RECT 862.950 60.000 865.050 64.050 ;
        RECT 871.950 61.950 874.050 64.050 ;
        RECT 863.400 58.350 864.600 60.000 ;
        RECT 862.950 55.950 865.050 58.050 ;
        RECT 865.950 55.950 868.050 58.050 ;
        RECT 866.400 53.400 867.600 55.650 ;
        RECT 866.400 49.050 867.450 53.400 ;
        RECT 875.400 49.050 876.450 169.950 ;
        RECT 865.950 46.950 868.050 49.050 ;
        RECT 874.950 46.950 877.050 49.050 ;
        RECT 856.950 28.950 859.050 31.050 ;
        RECT 854.400 26.400 858.450 27.450 ;
        RECT 865.950 27.000 868.050 31.050 ;
        RECT 841.950 22.950 844.050 25.050 ;
        RECT 844.950 22.950 847.050 25.050 ;
        RECT 847.950 22.950 850.050 25.050 ;
        RECT 850.950 22.950 853.050 25.050 ;
        RECT 845.400 21.900 846.600 22.650 ;
        RECT 851.400 21.900 852.600 22.650 ;
        RECT 857.400 22.050 858.450 26.400 ;
        RECT 866.400 25.350 867.600 27.000 ;
        RECT 862.950 22.950 865.050 25.050 ;
        RECT 865.950 22.950 868.050 25.050 ;
        RECT 844.950 19.800 847.050 21.900 ;
        RECT 850.950 19.800 853.050 21.900 ;
        RECT 856.950 19.950 859.050 22.050 ;
        RECT 863.400 21.900 864.600 22.650 ;
        RECT 862.950 19.800 865.050 21.900 ;
        RECT 835.950 16.950 838.050 19.050 ;
        RECT 754.950 13.950 757.050 16.050 ;
        RECT 760.950 13.950 763.050 16.050 ;
        RECT 781.950 13.950 784.050 16.050 ;
        RECT 736.950 4.950 739.050 7.050 ;
        RECT 407.400 3.000 415.050 3.450 ;
        RECT 407.400 2.400 414.450 3.000 ;
        RECT 595.950 1.950 598.050 4.050 ;
        RECT 673.950 1.950 676.050 4.050 ;
      LAYER metal3 ;
        RECT 454.950 819.600 457.050 820.050 ;
        RECT 484.950 819.600 487.050 820.050 ;
        RECT 454.950 818.400 487.050 819.600 ;
        RECT 454.950 817.950 457.050 818.400 ;
        RECT 484.950 817.950 487.050 818.400 ;
        RECT 394.950 816.600 397.050 817.050 ;
        RECT 409.950 816.600 412.050 817.050 ;
        RECT 394.950 815.400 412.050 816.600 ;
        RECT 394.950 814.950 397.050 815.400 ;
        RECT 409.950 814.950 412.050 815.400 ;
        RECT 205.950 813.600 208.050 814.050 ;
        RECT 217.950 813.600 220.050 814.050 ;
        RECT 205.950 812.400 220.050 813.600 ;
        RECT 205.950 811.950 208.050 812.400 ;
        RECT 217.950 811.950 220.050 812.400 ;
        RECT 277.950 813.600 280.050 814.050 ;
        RECT 313.950 813.600 316.050 814.050 ;
        RECT 385.950 813.600 388.050 814.050 ;
        RECT 277.950 812.400 388.050 813.600 ;
        RECT 277.950 811.950 280.050 812.400 ;
        RECT 313.950 811.950 316.050 812.400 ;
        RECT 385.950 811.950 388.050 812.400 ;
        RECT 391.950 813.600 394.050 814.050 ;
        RECT 406.950 813.600 409.050 814.050 ;
        RECT 391.950 812.400 409.050 813.600 ;
        RECT 391.950 811.950 394.050 812.400 ;
        RECT 406.950 811.950 409.050 812.400 ;
        RECT 421.950 813.600 424.050 814.050 ;
        RECT 469.950 813.600 472.050 814.050 ;
        RECT 421.950 812.400 472.050 813.600 ;
        RECT 421.950 811.950 424.050 812.400 ;
        RECT 469.950 811.950 472.050 812.400 ;
        RECT 481.950 813.600 484.050 814.050 ;
        RECT 565.950 813.600 568.050 814.050 ;
        RECT 481.950 812.400 568.050 813.600 ;
        RECT 481.950 811.950 484.050 812.400 ;
        RECT 565.950 811.950 568.050 812.400 ;
        RECT 574.950 813.600 577.050 814.050 ;
        RECT 595.950 813.600 598.050 814.050 ;
        RECT 574.950 812.400 598.050 813.600 ;
        RECT 574.950 811.950 577.050 812.400 ;
        RECT 595.950 811.950 598.050 812.400 ;
        RECT 817.950 813.600 820.050 814.050 ;
        RECT 853.950 813.600 856.050 814.050 ;
        RECT 817.950 812.400 856.050 813.600 ;
        RECT 817.950 811.950 820.050 812.400 ;
        RECT 853.950 811.950 856.050 812.400 ;
        RECT 97.950 810.600 100.050 811.050 ;
        RECT 112.950 810.600 115.050 811.050 ;
        RECT 97.950 809.400 115.050 810.600 ;
        RECT 97.950 808.950 100.050 809.400 ;
        RECT 112.950 808.950 115.050 809.400 ;
        RECT 388.950 810.600 391.050 811.050 ;
        RECT 394.950 810.600 397.050 811.050 ;
        RECT 388.950 809.400 397.050 810.600 ;
        RECT 388.950 808.950 391.050 809.400 ;
        RECT 394.950 808.950 397.050 809.400 ;
        RECT 418.950 810.600 421.050 811.050 ;
        RECT 478.950 810.600 481.050 811.050 ;
        RECT 418.950 809.400 481.050 810.600 ;
        RECT 418.950 808.950 421.050 809.400 ;
        RECT 478.950 808.950 481.050 809.400 ;
        RECT 31.950 806.100 34.050 808.200 ;
        RECT 49.950 807.600 52.050 808.200 ;
        RECT 55.950 807.600 58.050 808.200 ;
        RECT 49.950 806.400 58.050 807.600 ;
        RECT 49.950 806.100 52.050 806.400 ;
        RECT 55.950 806.100 58.050 806.400 ;
        RECT 91.950 807.750 94.050 808.200 ;
        RECT 103.950 807.750 106.050 808.200 ;
        RECT 91.950 806.550 106.050 807.750 ;
        RECT 121.950 807.600 124.050 808.200 ;
        RECT 91.950 806.100 94.050 806.550 ;
        RECT 103.950 806.100 106.050 806.550 ;
        RECT 107.400 806.400 124.050 807.600 ;
        RECT 32.400 804.600 33.600 806.100 ;
        RECT 40.950 804.600 43.050 805.050 ;
        RECT 32.400 803.400 43.050 804.600 ;
        RECT 40.950 802.950 43.050 803.400 ;
        RECT 56.400 802.050 57.600 806.100 ;
        RECT 52.950 800.400 57.600 802.050 ;
        RECT 73.950 801.600 76.050 801.900 ;
        RECT 91.950 801.600 94.050 802.050 ;
        RECT 107.400 801.900 108.600 806.400 ;
        RECT 121.950 806.100 124.050 806.400 ;
        RECT 196.950 807.600 199.050 808.200 ;
        RECT 211.950 807.600 214.050 808.200 ;
        RECT 220.950 807.750 223.050 808.200 ;
        RECT 226.950 807.750 229.050 808.200 ;
        RECT 196.950 806.400 216.600 807.600 ;
        RECT 196.950 806.100 199.050 806.400 ;
        RECT 211.950 806.100 214.050 806.400 ;
        RECT 215.400 804.600 216.600 806.400 ;
        RECT 220.950 806.550 229.050 807.750 ;
        RECT 220.950 806.100 223.050 806.550 ;
        RECT 226.950 806.100 229.050 806.550 ;
        RECT 241.950 807.600 244.050 808.050 ;
        RECT 250.950 807.600 253.050 808.200 ;
        RECT 241.950 806.400 253.050 807.600 ;
        RECT 241.950 805.950 244.050 806.400 ;
        RECT 250.950 806.100 253.050 806.400 ;
        RECT 268.950 807.600 271.050 808.200 ;
        RECT 289.950 807.600 292.050 808.200 ;
        RECT 301.950 807.600 304.050 808.050 ;
        RECT 268.950 806.400 304.050 807.600 ;
        RECT 268.950 806.100 271.050 806.400 ;
        RECT 289.950 806.100 292.050 806.400 ;
        RECT 301.950 805.950 304.050 806.400 ;
        RECT 322.950 807.600 325.050 808.050 ;
        RECT 328.950 807.600 331.050 808.200 ;
        RECT 367.950 807.600 370.050 808.200 ;
        RECT 382.950 807.600 385.050 808.200 ;
        RECT 403.950 807.600 406.050 808.200 ;
        RECT 322.950 806.400 331.050 807.600 ;
        RECT 322.950 805.950 325.050 806.400 ;
        RECT 328.950 806.100 331.050 806.400 ;
        RECT 332.400 806.400 385.050 807.600 ;
        RECT 259.950 804.600 262.050 805.050 ;
        RECT 332.400 804.600 333.600 806.400 ;
        RECT 367.950 806.100 370.050 806.400 ;
        RECT 382.950 806.100 385.050 806.400 ;
        RECT 386.400 806.400 406.050 807.600 ;
        RECT 386.400 804.600 387.600 806.400 ;
        RECT 403.950 806.100 406.050 806.400 ;
        RECT 463.950 807.750 466.050 808.200 ;
        RECT 469.950 807.750 472.050 808.200 ;
        RECT 463.950 806.550 472.050 807.750 ;
        RECT 463.950 806.100 466.050 806.550 ;
        RECT 469.950 806.100 472.050 806.550 ;
        RECT 478.950 807.600 481.050 808.200 ;
        RECT 496.950 807.600 499.050 811.050 ;
        RECT 646.950 810.600 649.050 811.050 ;
        RECT 670.950 810.600 673.050 811.050 ;
        RECT 646.950 809.400 673.050 810.600 ;
        RECT 646.950 808.950 649.050 809.400 ;
        RECT 670.950 808.950 673.050 809.400 ;
        RECT 502.950 807.600 505.050 808.200 ;
        RECT 478.950 806.400 495.600 807.600 ;
        RECT 496.950 807.000 505.050 807.600 ;
        RECT 497.400 806.400 505.050 807.000 ;
        RECT 478.950 806.100 481.050 806.400 ;
        RECT 472.950 804.600 475.050 805.050 ;
        RECT 215.400 803.400 262.050 804.600 ;
        RECT 259.950 802.950 262.050 803.400 ;
        RECT 311.400 803.400 333.600 804.600 ;
        RECT 350.400 803.400 387.600 804.600 ;
        RECT 413.400 803.400 475.050 804.600 ;
        RECT 494.400 804.600 495.600 806.400 ;
        RECT 502.950 806.100 505.050 806.400 ;
        RECT 511.950 807.600 514.050 808.050 ;
        RECT 559.950 807.600 562.050 808.050 ;
        RECT 511.950 806.400 562.050 807.600 ;
        RECT 511.950 805.950 514.050 806.400 ;
        RECT 559.950 805.950 562.050 806.400 ;
        RECT 565.950 807.750 568.050 808.200 ;
        RECT 583.950 807.750 586.050 808.200 ;
        RECT 565.950 806.550 586.050 807.750 ;
        RECT 565.950 806.100 568.050 806.550 ;
        RECT 583.950 806.100 586.050 806.550 ;
        RECT 628.950 807.600 631.050 808.200 ;
        RECT 634.950 807.600 637.050 808.200 ;
        RECT 628.950 806.400 637.050 807.600 ;
        RECT 628.950 806.100 631.050 806.400 ;
        RECT 634.950 806.100 637.050 806.400 ;
        RECT 700.950 807.750 703.050 808.200 ;
        RECT 709.950 807.750 712.050 808.200 ;
        RECT 700.950 806.550 712.050 807.750 ;
        RECT 700.950 806.100 703.050 806.550 ;
        RECT 709.950 806.100 712.050 806.550 ;
        RECT 715.950 807.600 718.050 808.200 ;
        RECT 730.950 807.600 733.050 808.200 ;
        RECT 715.950 806.400 733.050 807.600 ;
        RECT 715.950 806.100 718.050 806.400 ;
        RECT 730.950 806.100 733.050 806.400 ;
        RECT 736.950 807.750 739.050 808.200 ;
        RECT 745.950 807.750 748.050 808.200 ;
        RECT 736.950 807.600 748.050 807.750 ;
        RECT 757.950 807.600 760.050 808.200 ;
        RECT 736.950 806.550 760.050 807.600 ;
        RECT 736.950 806.100 739.050 806.550 ;
        RECT 745.950 806.400 760.050 806.550 ;
        RECT 745.950 806.100 748.050 806.400 ;
        RECT 757.950 806.100 760.050 806.400 ;
        RECT 769.950 807.750 772.050 808.200 ;
        RECT 775.950 807.750 778.050 808.200 ;
        RECT 769.950 806.550 778.050 807.750 ;
        RECT 781.950 807.600 784.050 808.200 ;
        RECT 769.950 806.100 772.050 806.550 ;
        RECT 775.950 806.100 778.050 806.550 ;
        RECT 779.400 806.400 784.050 807.600 ;
        RECT 592.950 804.600 595.050 805.050 ;
        RECT 667.950 804.600 670.050 805.050 ;
        RECT 779.400 804.600 780.600 806.400 ;
        RECT 781.950 806.100 784.050 806.400 ;
        RECT 826.950 807.750 829.050 808.200 ;
        RECT 832.950 807.750 835.050 808.200 ;
        RECT 826.950 806.550 835.050 807.750 ;
        RECT 826.950 806.100 829.050 806.550 ;
        RECT 832.950 806.100 835.050 806.550 ;
        RECT 838.950 807.750 841.050 808.200 ;
        RECT 844.950 807.750 847.050 808.200 ;
        RECT 838.950 806.550 847.050 807.750 ;
        RECT 838.950 806.100 841.050 806.550 ;
        RECT 844.950 806.100 847.050 806.550 ;
        RECT 494.400 803.400 501.600 804.600 ;
        RECT 73.950 800.400 94.050 801.600 ;
        RECT 52.950 799.950 57.000 800.400 ;
        RECT 73.950 799.800 76.050 800.400 ;
        RECT 91.950 799.950 94.050 800.400 ;
        RECT 106.950 799.800 109.050 801.900 ;
        RECT 178.950 801.600 181.050 801.900 ;
        RECT 205.950 801.600 208.050 802.050 ;
        RECT 178.950 800.400 208.050 801.600 ;
        RECT 178.950 799.800 181.050 800.400 ;
        RECT 205.950 799.950 208.050 800.400 ;
        RECT 214.950 801.600 217.050 801.900 ;
        RECT 229.950 801.600 232.050 801.900 ;
        RECT 214.950 800.400 232.050 801.600 ;
        RECT 214.950 799.800 217.050 800.400 ;
        RECT 229.950 799.800 232.050 800.400 ;
        RECT 235.950 801.450 238.050 801.900 ;
        RECT 241.950 801.450 244.050 801.900 ;
        RECT 235.950 800.250 244.050 801.450 ;
        RECT 235.950 799.800 238.050 800.250 ;
        RECT 241.950 799.800 244.050 800.250 ;
        RECT 271.950 801.450 274.050 801.900 ;
        RECT 277.950 801.450 280.050 801.900 ;
        RECT 271.950 800.250 280.050 801.450 ;
        RECT 271.950 799.800 274.050 800.250 ;
        RECT 277.950 799.800 280.050 800.250 ;
        RECT 295.950 801.600 298.050 801.900 ;
        RECT 307.950 801.600 310.050 801.900 ;
        RECT 295.950 800.400 310.050 801.600 ;
        RECT 295.950 799.800 298.050 800.400 ;
        RECT 307.950 799.800 310.050 800.400 ;
        RECT 46.950 798.600 49.050 799.050 ;
        RECT 100.950 798.600 103.050 799.050 ;
        RECT 46.950 797.400 103.050 798.600 ;
        RECT 46.950 796.950 49.050 797.400 ;
        RECT 100.950 796.950 103.050 797.400 ;
        RECT 142.950 798.600 145.050 799.050 ;
        RECT 169.950 798.600 172.050 799.050 ;
        RECT 142.950 797.400 172.050 798.600 ;
        RECT 142.950 796.950 145.050 797.400 ;
        RECT 169.950 796.950 172.050 797.400 ;
        RECT 274.950 798.600 277.050 799.050 ;
        RECT 311.400 798.600 312.600 803.400 ;
        RECT 350.400 801.900 351.600 803.400 ;
        RECT 413.400 801.900 414.600 803.400 ;
        RECT 472.950 802.950 475.050 803.400 ;
        RECT 500.400 801.900 501.600 803.400 ;
        RECT 592.950 803.400 670.050 804.600 ;
        RECT 592.950 802.950 595.050 803.400 ;
        RECT 349.950 799.800 352.050 801.900 ;
        RECT 385.950 801.600 388.050 801.900 ;
        RECT 406.950 801.600 409.050 801.900 ;
        RECT 385.950 800.400 409.050 801.600 ;
        RECT 385.950 799.800 388.050 800.400 ;
        RECT 406.950 799.800 409.050 800.400 ;
        RECT 412.950 799.800 415.050 801.900 ;
        RECT 499.950 799.800 502.050 801.900 ;
        RECT 505.950 801.450 508.050 801.900 ;
        RECT 511.950 801.450 514.050 801.900 ;
        RECT 505.950 800.250 514.050 801.450 ;
        RECT 505.950 799.800 508.050 800.250 ;
        RECT 511.950 799.800 514.050 800.250 ;
        RECT 565.950 801.600 568.050 802.050 ;
        RECT 626.400 801.900 627.600 803.400 ;
        RECT 667.950 802.950 670.050 803.400 ;
        RECT 755.400 803.400 780.600 804.600 ;
        RECT 571.950 801.600 574.050 801.900 ;
        RECT 565.950 800.400 574.050 801.600 ;
        RECT 565.950 799.950 568.050 800.400 ;
        RECT 571.950 799.800 574.050 800.400 ;
        RECT 625.950 799.800 628.050 801.900 ;
        RECT 646.950 801.450 649.050 801.900 ;
        RECT 652.950 801.450 655.050 801.900 ;
        RECT 646.950 800.250 655.050 801.450 ;
        RECT 646.950 799.800 649.050 800.250 ;
        RECT 652.950 799.800 655.050 800.250 ;
        RECT 670.950 801.600 673.050 802.050 ;
        RECT 755.400 801.900 756.600 803.400 ;
        RECT 712.950 801.600 715.050 801.900 ;
        RECT 670.950 800.400 715.050 801.600 ;
        RECT 670.950 799.950 673.050 800.400 ;
        RECT 712.950 799.800 715.050 800.400 ;
        RECT 739.950 801.600 742.050 801.900 ;
        RECT 754.950 801.600 757.050 801.900 ;
        RECT 739.950 800.400 757.050 801.600 ;
        RECT 739.950 799.800 742.050 800.400 ;
        RECT 754.950 799.800 757.050 800.400 ;
        RECT 784.950 801.600 787.050 801.900 ;
        RECT 796.950 801.600 799.050 801.900 ;
        RECT 784.950 800.400 799.050 801.600 ;
        RECT 784.950 799.800 787.050 800.400 ;
        RECT 796.950 799.800 799.050 800.400 ;
        RECT 805.950 801.600 808.050 802.050 ;
        RECT 835.950 801.600 838.050 801.900 ;
        RECT 805.950 800.400 838.050 801.600 ;
        RECT 805.950 799.950 808.050 800.400 ;
        RECT 835.950 799.800 838.050 800.400 ;
        RECT 844.950 801.450 847.050 801.900 ;
        RECT 850.950 801.450 853.050 801.900 ;
        RECT 844.950 800.250 853.050 801.450 ;
        RECT 844.950 799.800 847.050 800.250 ;
        RECT 850.950 799.800 853.050 800.250 ;
        RECT 274.950 797.400 312.600 798.600 ;
        RECT 466.950 798.600 469.050 799.050 ;
        RECT 481.950 798.600 484.050 799.050 ;
        RECT 466.950 797.400 484.050 798.600 ;
        RECT 274.950 796.950 277.050 797.400 ;
        RECT 466.950 796.950 469.050 797.400 ;
        RECT 481.950 796.950 484.050 797.400 ;
        RECT 556.950 798.600 559.050 799.050 ;
        RECT 610.950 798.600 613.050 799.050 ;
        RECT 661.950 798.600 664.050 799.050 ;
        RECT 556.950 797.400 664.050 798.600 ;
        RECT 556.950 796.950 559.050 797.400 ;
        RECT 610.950 796.950 613.050 797.400 ;
        RECT 661.950 796.950 664.050 797.400 ;
        RECT 259.950 795.600 262.050 796.050 ;
        RECT 265.950 795.600 268.050 796.050 ;
        RECT 316.950 795.600 319.050 796.050 ;
        RECT 259.950 794.400 319.050 795.600 ;
        RECT 259.950 793.950 262.050 794.400 ;
        RECT 265.950 793.950 268.050 794.400 ;
        RECT 316.950 793.950 319.050 794.400 ;
        RECT 373.950 795.600 376.050 796.050 ;
        RECT 394.950 795.600 397.050 796.050 ;
        RECT 373.950 794.400 397.050 795.600 ;
        RECT 373.950 793.950 376.050 794.400 ;
        RECT 394.950 793.950 397.050 794.400 ;
        RECT 400.950 795.600 403.050 796.050 ;
        RECT 454.950 795.600 457.050 796.050 ;
        RECT 400.950 794.400 457.050 795.600 ;
        RECT 400.950 793.950 403.050 794.400 ;
        RECT 454.950 793.950 457.050 794.400 ;
        RECT 559.950 795.600 562.050 796.050 ;
        RECT 592.950 795.600 595.050 796.050 ;
        RECT 559.950 794.400 595.050 795.600 ;
        RECT 559.950 793.950 562.050 794.400 ;
        RECT 592.950 793.950 595.050 794.400 ;
        RECT 667.950 795.600 670.050 796.050 ;
        RECT 706.950 795.600 709.050 796.050 ;
        RECT 667.950 794.400 709.050 795.600 ;
        RECT 667.950 793.950 670.050 794.400 ;
        RECT 706.950 793.950 709.050 794.400 ;
        RECT 100.950 792.600 103.050 793.050 ;
        RECT 106.950 792.600 109.050 793.050 ;
        RECT 100.950 791.400 109.050 792.600 ;
        RECT 100.950 790.950 103.050 791.400 ;
        RECT 106.950 790.950 109.050 791.400 ;
        RECT 112.950 792.600 115.050 793.050 ;
        RECT 118.950 792.600 121.050 793.050 ;
        RECT 220.950 792.600 223.050 793.050 ;
        RECT 112.950 791.400 223.050 792.600 ;
        RECT 112.950 790.950 115.050 791.400 ;
        RECT 118.950 790.950 121.050 791.400 ;
        RECT 220.950 790.950 223.050 791.400 ;
        RECT 268.950 792.600 271.050 792.900 ;
        RECT 274.950 792.600 277.050 793.050 ;
        RECT 268.950 791.400 277.050 792.600 ;
        RECT 268.950 790.800 271.050 791.400 ;
        RECT 274.950 790.950 277.050 791.400 ;
        RECT 571.950 792.600 574.050 793.050 ;
        RECT 598.950 792.600 601.050 793.050 ;
        RECT 571.950 791.400 601.050 792.600 ;
        RECT 571.950 790.950 574.050 791.400 ;
        RECT 598.950 790.950 601.050 791.400 ;
        RECT 718.950 792.600 721.050 793.050 ;
        RECT 763.950 792.600 766.050 793.050 ;
        RECT 718.950 791.400 766.050 792.600 ;
        RECT 718.950 790.950 721.050 791.400 ;
        RECT 763.950 790.950 766.050 791.400 ;
        RECT 169.950 789.600 172.050 790.050 ;
        RECT 442.950 789.600 445.050 790.050 ;
        RECT 448.950 789.600 451.050 790.050 ;
        RECT 169.950 789.000 195.600 789.600 ;
        RECT 169.950 788.400 196.050 789.000 ;
        RECT 169.950 787.950 172.050 788.400 ;
        RECT 4.950 786.600 7.050 787.050 ;
        RECT 82.950 786.600 85.050 787.050 ;
        RECT 88.950 786.600 91.050 787.050 ;
        RECT 103.950 786.600 106.050 787.050 ;
        RECT 142.950 786.600 145.050 787.050 ;
        RECT 4.950 785.400 145.050 786.600 ;
        RECT 4.950 784.950 7.050 785.400 ;
        RECT 82.950 784.950 85.050 785.400 ;
        RECT 88.950 784.950 91.050 785.400 ;
        RECT 103.950 784.950 106.050 785.400 ;
        RECT 142.950 784.950 145.050 785.400 ;
        RECT 193.950 784.950 196.050 788.400 ;
        RECT 442.950 788.400 451.050 789.600 ;
        RECT 442.950 787.950 445.050 788.400 ;
        RECT 448.950 787.950 451.050 788.400 ;
        RECT 220.950 786.600 223.050 787.050 ;
        RECT 247.950 786.600 250.050 787.050 ;
        RECT 268.950 786.600 271.050 787.050 ;
        RECT 220.950 785.400 271.050 786.600 ;
        RECT 220.950 784.950 223.050 785.400 ;
        RECT 247.950 784.950 250.050 785.400 ;
        RECT 268.950 784.950 271.050 785.400 ;
        RECT 472.950 786.600 475.050 787.050 ;
        RECT 640.950 786.600 643.050 787.050 ;
        RECT 691.950 786.600 694.050 787.050 ;
        RECT 472.950 785.400 694.050 786.600 ;
        RECT 472.950 784.950 475.050 785.400 ;
        RECT 640.950 784.950 643.050 785.400 ;
        RECT 691.950 784.950 694.050 785.400 ;
        RECT 727.950 786.600 730.050 787.050 ;
        RECT 769.950 786.600 772.050 787.050 ;
        RECT 727.950 785.400 772.050 786.600 ;
        RECT 727.950 784.950 730.050 785.400 ;
        RECT 769.950 784.950 772.050 785.400 ;
        RECT 154.950 783.600 157.050 784.050 ;
        RECT 328.950 783.600 331.050 784.050 ;
        RECT 154.950 782.400 331.050 783.600 ;
        RECT 154.950 781.950 157.050 782.400 ;
        RECT 328.950 781.950 331.050 782.400 ;
        RECT 523.950 783.600 526.050 784.050 ;
        RECT 532.950 783.600 535.050 784.050 ;
        RECT 523.950 782.400 535.050 783.600 ;
        RECT 523.950 781.950 526.050 782.400 ;
        RECT 532.950 781.950 535.050 782.400 ;
        RECT 193.950 780.600 196.050 781.050 ;
        RECT 307.950 780.600 310.050 781.050 ;
        RECT 340.950 780.600 343.050 781.050 ;
        RECT 193.950 779.400 343.050 780.600 ;
        RECT 193.950 778.950 196.050 779.400 ;
        RECT 307.950 778.950 310.050 779.400 ;
        RECT 340.950 778.950 343.050 779.400 ;
        RECT 403.950 780.600 406.050 781.050 ;
        RECT 421.950 780.600 424.050 781.050 ;
        RECT 403.950 779.400 424.050 780.600 ;
        RECT 403.950 778.950 406.050 779.400 ;
        RECT 421.950 778.950 424.050 779.400 ;
        RECT 436.950 780.600 439.050 781.050 ;
        RECT 514.950 780.600 517.050 781.050 ;
        RECT 556.950 780.600 559.050 781.050 ;
        RECT 565.950 780.600 568.050 781.050 ;
        RECT 436.950 779.400 568.050 780.600 ;
        RECT 436.950 778.950 439.050 779.400 ;
        RECT 514.950 778.950 517.050 779.400 ;
        RECT 556.950 778.950 559.050 779.400 ;
        RECT 565.950 778.950 568.050 779.400 ;
        RECT 577.950 780.600 580.050 781.050 ;
        RECT 700.950 780.600 703.050 781.050 ;
        RECT 733.950 780.600 736.050 781.050 ;
        RECT 577.950 779.400 736.050 780.600 ;
        RECT 577.950 778.950 580.050 779.400 ;
        RECT 700.950 778.950 703.050 779.400 ;
        RECT 733.950 778.950 736.050 779.400 ;
        RECT 10.950 777.600 13.050 778.050 ;
        RECT 16.950 777.600 19.050 778.050 ;
        RECT 10.950 776.400 19.050 777.600 ;
        RECT 10.950 775.950 13.050 776.400 ;
        RECT 16.950 775.950 19.050 776.400 ;
        RECT 181.950 777.600 184.050 778.050 ;
        RECT 388.950 777.600 391.050 778.050 ;
        RECT 181.950 776.400 391.050 777.600 ;
        RECT 181.950 775.950 184.050 776.400 ;
        RECT 388.950 775.950 391.050 776.400 ;
        RECT 487.950 777.600 490.050 778.050 ;
        RECT 526.950 777.600 529.050 778.050 ;
        RECT 487.950 776.400 529.050 777.600 ;
        RECT 487.950 775.950 490.050 776.400 ;
        RECT 526.950 775.950 529.050 776.400 ;
        RECT 772.950 777.600 775.050 778.050 ;
        RECT 805.950 777.600 808.050 778.050 ;
        RECT 772.950 776.400 808.050 777.600 ;
        RECT 772.950 775.950 775.050 776.400 ;
        RECT 805.950 775.950 808.050 776.400 ;
        RECT 421.950 774.600 424.050 775.050 ;
        RECT 601.950 774.600 604.050 775.050 ;
        RECT 421.950 773.400 604.050 774.600 ;
        RECT 421.950 772.950 424.050 773.400 ;
        RECT 601.950 772.950 604.050 773.400 ;
        RECT 721.950 774.600 724.050 775.050 ;
        RECT 736.950 774.600 739.050 775.050 ;
        RECT 820.950 774.600 823.050 775.050 ;
        RECT 721.950 773.400 823.050 774.600 ;
        RECT 721.950 772.950 724.050 773.400 ;
        RECT 736.950 772.950 739.050 773.400 ;
        RECT 820.950 772.950 823.050 773.400 ;
        RECT 40.950 771.600 43.050 772.050 ;
        RECT 145.950 771.600 148.050 772.050 ;
        RECT 40.950 770.400 148.050 771.600 ;
        RECT 40.950 769.950 43.050 770.400 ;
        RECT 145.950 769.950 148.050 770.400 ;
        RECT 169.950 771.600 172.050 772.050 ;
        RECT 187.950 771.600 190.050 772.050 ;
        RECT 169.950 770.400 190.050 771.600 ;
        RECT 169.950 769.950 172.050 770.400 ;
        RECT 187.950 769.950 190.050 770.400 ;
        RECT 211.950 771.600 214.050 772.050 ;
        RECT 262.950 771.600 265.050 772.050 ;
        RECT 298.950 771.600 301.050 772.050 ;
        RECT 211.950 770.400 301.050 771.600 ;
        RECT 211.950 769.950 214.050 770.400 ;
        RECT 262.950 769.950 265.050 770.400 ;
        RECT 298.950 769.950 301.050 770.400 ;
        RECT 364.950 771.600 367.050 772.050 ;
        RECT 412.950 771.600 415.050 772.050 ;
        RECT 364.950 770.400 415.050 771.600 ;
        RECT 364.950 769.950 367.050 770.400 ;
        RECT 412.950 769.950 415.050 770.400 ;
        RECT 439.950 771.600 442.050 772.050 ;
        RECT 445.950 771.600 448.050 772.050 ;
        RECT 439.950 770.400 448.050 771.600 ;
        RECT 439.950 769.950 442.050 770.400 ;
        RECT 445.950 769.950 448.050 770.400 ;
        RECT 451.950 771.600 454.050 772.050 ;
        RECT 493.950 771.600 496.050 772.050 ;
        RECT 451.950 770.400 496.050 771.600 ;
        RECT 451.950 769.950 454.050 770.400 ;
        RECT 493.950 769.950 496.050 770.400 ;
        RECT 616.950 771.600 619.050 772.050 ;
        RECT 676.950 771.600 679.050 772.050 ;
        RECT 616.950 770.400 679.050 771.600 ;
        RECT 616.950 769.950 619.050 770.400 ;
        RECT 676.950 769.950 679.050 770.400 ;
        RECT 691.950 771.600 694.050 772.050 ;
        RECT 712.950 771.600 715.050 772.050 ;
        RECT 691.950 770.400 715.050 771.600 ;
        RECT 691.950 769.950 694.050 770.400 ;
        RECT 712.950 769.950 715.050 770.400 ;
        RECT 724.950 771.600 727.050 772.050 ;
        RECT 778.950 771.600 781.050 772.050 ;
        RECT 724.950 770.400 781.050 771.600 ;
        RECT 724.950 769.950 727.050 770.400 ;
        RECT 778.950 769.950 781.050 770.400 ;
        RECT 148.950 768.600 151.050 769.050 ;
        RECT 175.950 768.600 178.050 769.050 ;
        RECT 208.950 768.600 211.050 769.050 ;
        RECT 148.950 767.400 211.050 768.600 ;
        RECT 148.950 766.950 151.050 767.400 ;
        RECT 175.950 766.950 178.050 767.400 ;
        RECT 208.950 766.950 211.050 767.400 ;
        RECT 229.950 768.600 232.050 769.050 ;
        RECT 241.950 768.600 244.050 769.050 ;
        RECT 229.950 767.400 244.050 768.600 ;
        RECT 229.950 766.950 232.050 767.400 ;
        RECT 241.950 766.950 244.050 767.400 ;
        RECT 301.950 768.600 304.050 769.050 ;
        RECT 352.950 768.600 355.050 769.050 ;
        RECT 301.950 767.400 355.050 768.600 ;
        RECT 301.950 766.950 304.050 767.400 ;
        RECT 352.950 766.950 355.050 767.400 ;
        RECT 358.950 768.600 361.050 769.050 ;
        RECT 448.950 768.600 451.050 769.050 ;
        RECT 358.950 767.400 451.050 768.600 ;
        RECT 358.950 766.950 361.050 767.400 ;
        RECT 448.950 766.950 451.050 767.400 ;
        RECT 460.950 768.600 463.050 769.050 ;
        RECT 475.950 768.600 478.050 769.050 ;
        RECT 460.950 767.400 478.050 768.600 ;
        RECT 460.950 766.950 463.050 767.400 ;
        RECT 475.950 766.950 478.050 767.400 ;
        RECT 574.950 768.600 577.050 769.050 ;
        RECT 595.950 768.600 598.050 769.050 ;
        RECT 574.950 767.400 598.050 768.600 ;
        RECT 574.950 766.950 577.050 767.400 ;
        RECT 595.950 766.950 598.050 767.400 ;
        RECT 682.950 768.600 685.050 769.050 ;
        RECT 721.950 768.600 724.050 769.050 ;
        RECT 682.950 767.400 724.050 768.600 ;
        RECT 682.950 766.950 685.050 767.400 ;
        RECT 721.950 766.950 724.050 767.400 ;
        RECT 817.950 768.600 820.050 769.050 ;
        RECT 826.950 768.600 829.050 769.050 ;
        RECT 856.950 768.600 859.050 769.050 ;
        RECT 862.950 768.600 865.050 769.050 ;
        RECT 817.950 767.400 865.050 768.600 ;
        RECT 817.950 766.950 820.050 767.400 ;
        RECT 826.950 766.950 829.050 767.400 ;
        RECT 856.950 766.950 859.050 767.400 ;
        RECT 862.950 766.950 865.050 767.400 ;
        RECT 82.950 765.600 85.050 766.050 ;
        RECT 121.950 765.600 124.050 766.050 ;
        RECT 82.950 764.400 124.050 765.600 ;
        RECT 82.950 763.950 85.050 764.400 ;
        RECT 121.950 763.950 124.050 764.400 ;
        RECT 298.950 765.600 301.050 766.050 ;
        RECT 355.950 765.600 358.050 766.050 ;
        RECT 298.950 764.400 358.050 765.600 ;
        RECT 298.950 763.950 301.050 764.400 ;
        RECT 355.950 763.950 358.050 764.400 ;
        RECT 634.950 765.600 637.050 766.050 ;
        RECT 643.950 765.600 646.050 766.050 ;
        RECT 634.950 764.400 646.050 765.600 ;
        RECT 634.950 763.950 637.050 764.400 ;
        RECT 643.950 763.950 646.050 764.400 ;
        RECT 751.950 765.600 754.050 766.050 ;
        RECT 766.950 765.600 769.050 766.050 ;
        RECT 751.950 764.400 769.050 765.600 ;
        RECT 751.950 763.950 754.050 764.400 ;
        RECT 766.950 763.950 769.050 764.400 ;
        RECT 7.950 762.750 10.050 763.200 ;
        RECT 16.950 762.750 19.050 763.200 ;
        RECT 7.950 761.550 19.050 762.750 ;
        RECT 7.950 761.100 10.050 761.550 ;
        RECT 16.950 761.100 19.050 761.550 ;
        RECT 22.950 762.750 25.050 763.200 ;
        RECT 28.950 762.750 31.050 763.200 ;
        RECT 22.950 761.550 31.050 762.750 ;
        RECT 22.950 761.100 25.050 761.550 ;
        RECT 28.950 761.100 31.050 761.550 ;
        RECT 34.950 761.100 37.050 763.200 ;
        RECT 46.950 762.600 49.050 763.050 ;
        RECT 58.950 762.600 61.050 763.200 ;
        RECT 46.950 761.400 61.050 762.600 ;
        RECT 35.400 757.050 36.600 761.100 ;
        RECT 46.950 760.950 49.050 761.400 ;
        RECT 58.950 761.100 61.050 761.400 ;
        RECT 67.950 762.750 70.050 763.200 ;
        RECT 76.950 762.750 79.050 763.200 ;
        RECT 67.950 761.550 79.050 762.750 ;
        RECT 67.950 761.100 70.050 761.550 ;
        RECT 76.950 761.100 79.050 761.550 ;
        RECT 97.950 761.100 100.050 763.200 ;
        RECT 130.950 762.600 133.050 763.200 ;
        RECT 116.400 761.400 133.050 762.600 ;
        RECT 19.950 756.600 22.050 756.900 ;
        RECT 11.400 756.000 22.050 756.600 ;
        RECT 10.950 755.400 22.050 756.000 ;
        RECT 10.950 751.950 13.050 755.400 ;
        RECT 19.950 754.800 22.050 755.400 ;
        RECT 31.950 755.400 36.600 757.050 ;
        RECT 49.950 756.600 52.050 757.050 ;
        RECT 55.950 756.600 58.050 756.900 ;
        RECT 49.950 755.400 58.050 756.600 ;
        RECT 31.950 754.950 36.000 755.400 ;
        RECT 49.950 754.950 52.050 755.400 ;
        RECT 55.950 754.800 58.050 755.400 ;
        RECT 79.950 756.600 82.050 756.900 ;
        RECT 98.400 756.600 99.600 761.100 ;
        RECT 116.400 756.900 117.600 761.400 ;
        RECT 130.950 761.100 133.050 761.400 ;
        RECT 145.950 759.600 148.050 763.050 ;
        RECT 160.950 762.750 163.050 763.200 ;
        RECT 169.950 762.750 172.050 763.200 ;
        RECT 160.950 761.550 172.050 762.750 ;
        RECT 160.950 761.100 163.050 761.550 ;
        RECT 169.950 761.100 172.050 761.550 ;
        RECT 202.950 762.750 205.050 763.200 ;
        RECT 226.950 762.750 229.050 763.200 ;
        RECT 202.950 761.550 229.050 762.750 ;
        RECT 202.950 761.100 205.050 761.550 ;
        RECT 226.950 761.100 229.050 761.550 ;
        RECT 235.950 762.750 238.050 763.200 ;
        RECT 247.800 762.750 249.900 763.200 ;
        RECT 235.950 761.550 249.900 762.750 ;
        RECT 235.950 761.100 238.050 761.550 ;
        RECT 247.800 761.100 249.900 761.550 ;
        RECT 250.950 762.750 253.050 763.200 ;
        RECT 256.950 762.750 259.050 763.200 ;
        RECT 250.950 761.550 259.050 762.750 ;
        RECT 277.950 762.600 280.050 763.200 ;
        RECT 295.950 762.600 298.050 763.200 ;
        RECT 250.950 761.100 253.050 761.550 ;
        RECT 256.950 761.100 259.050 761.550 ;
        RECT 260.400 761.400 280.050 762.600 ;
        RECT 260.400 759.600 261.600 761.400 ;
        RECT 277.950 761.100 280.050 761.400 ;
        RECT 290.400 761.400 298.050 762.600 ;
        RECT 290.400 760.050 291.600 761.400 ;
        RECT 295.950 761.100 298.050 761.400 ;
        RECT 334.950 761.100 337.050 763.200 ;
        RECT 343.950 762.750 346.050 763.200 ;
        RECT 349.950 762.750 352.050 763.200 ;
        RECT 343.950 761.550 352.050 762.750 ;
        RECT 343.950 761.100 346.050 761.550 ;
        RECT 349.950 761.100 352.050 761.550 ;
        RECT 373.950 762.600 376.050 763.200 ;
        RECT 382.950 762.600 385.050 763.050 ;
        RECT 373.950 761.400 385.050 762.600 ;
        RECT 373.950 761.100 376.050 761.400 ;
        RECT 288.000 759.900 291.600 760.050 ;
        RECT 145.950 759.000 153.600 759.600 ;
        RECT 146.400 758.400 153.600 759.000 ;
        RECT 79.950 755.400 99.600 756.600 ;
        RECT 115.950 756.600 118.050 756.900 ;
        RECT 139.950 756.600 142.050 757.050 ;
        RECT 152.400 756.900 153.600 758.400 ;
        RECT 245.400 758.400 261.600 759.600 ;
        RECT 286.950 758.400 291.600 759.900 ;
        RECT 115.950 755.400 142.050 756.600 ;
        RECT 79.950 754.800 82.050 755.400 ;
        RECT 115.950 754.800 118.050 755.400 ;
        RECT 139.950 754.950 142.050 755.400 ;
        RECT 151.950 754.800 154.050 756.900 ;
        RECT 211.950 756.450 214.050 756.900 ;
        RECT 220.950 756.450 223.050 756.900 ;
        RECT 211.950 755.250 223.050 756.450 ;
        RECT 211.950 754.800 214.050 755.250 ;
        RECT 220.950 754.800 223.050 755.250 ;
        RECT 226.950 756.600 229.050 757.050 ;
        RECT 245.400 756.900 246.600 758.400 ;
        RECT 286.950 757.950 291.000 758.400 ;
        RECT 286.950 757.800 289.050 757.950 ;
        RECT 238.950 756.600 241.050 756.900 ;
        RECT 226.950 755.400 241.050 756.600 ;
        RECT 226.950 754.950 229.050 755.400 ;
        RECT 238.950 754.800 241.050 755.400 ;
        RECT 244.950 754.800 247.050 756.900 ;
        RECT 253.950 756.600 256.050 757.050 ;
        RECT 259.950 756.600 262.050 756.900 ;
        RECT 253.950 755.400 262.050 756.600 ;
        RECT 253.950 754.950 256.050 755.400 ;
        RECT 259.950 754.800 262.050 755.400 ;
        RECT 316.950 756.600 319.050 756.900 ;
        RECT 331.950 756.600 334.050 756.900 ;
        RECT 316.950 755.400 334.050 756.600 ;
        RECT 335.400 756.600 336.600 761.100 ;
        RECT 382.950 760.950 385.050 761.400 ;
        RECT 394.950 762.750 397.050 763.200 ;
        RECT 400.950 762.750 403.050 763.200 ;
        RECT 394.950 761.550 403.050 762.750 ;
        RECT 394.950 761.100 397.050 761.550 ;
        RECT 400.950 761.100 403.050 761.550 ;
        RECT 418.950 759.600 421.050 763.050 ;
        RECT 442.950 760.950 445.050 763.050 ;
        RECT 454.950 761.100 457.050 763.200 ;
        RECT 472.800 761.100 474.900 763.200 ;
        RECT 475.950 762.600 480.000 763.050 ;
        RECT 505.950 762.600 508.050 763.200 ;
        RECT 514.950 762.600 517.050 763.200 ;
        RECT 389.400 759.000 421.050 759.600 ;
        RECT 389.400 758.400 420.600 759.000 ;
        RECT 352.950 756.600 355.050 756.900 ;
        RECT 335.400 755.400 355.050 756.600 ;
        RECT 316.950 754.800 319.050 755.400 ;
        RECT 331.950 754.800 334.050 755.400 ;
        RECT 352.950 754.800 355.050 755.400 ;
        RECT 358.950 756.600 361.050 756.900 ;
        RECT 376.950 756.600 379.050 756.900 ;
        RECT 389.400 756.600 390.600 758.400 ;
        RECT 358.950 755.400 390.600 756.600 ;
        RECT 391.950 756.450 394.050 756.900 ;
        RECT 403.950 756.450 406.050 756.900 ;
        RECT 358.950 754.800 361.050 755.400 ;
        RECT 376.950 754.800 379.050 755.400 ;
        RECT 391.950 755.250 406.050 756.450 ;
        RECT 391.950 754.800 394.050 755.250 ;
        RECT 403.950 754.800 406.050 755.250 ;
        RECT 415.950 756.450 418.050 756.900 ;
        RECT 421.950 756.450 424.050 756.900 ;
        RECT 415.950 755.250 424.050 756.450 ;
        RECT 443.400 756.600 444.600 760.950 ;
        RECT 451.950 756.600 454.050 756.900 ;
        RECT 443.400 755.400 454.050 756.600 ;
        RECT 455.400 756.600 456.600 761.100 ;
        RECT 473.400 757.050 474.600 761.100 ;
        RECT 475.950 760.950 480.600 762.600 ;
        RECT 505.950 761.400 517.050 762.600 ;
        RECT 505.950 761.100 508.050 761.400 ;
        RECT 514.950 761.100 517.050 761.400 ;
        RECT 550.950 762.750 553.050 763.200 ;
        RECT 556.950 762.750 559.050 763.200 ;
        RECT 550.950 761.550 559.050 762.750 ;
        RECT 550.950 761.100 553.050 761.550 ;
        RECT 556.950 761.100 559.050 761.550 ;
        RECT 571.950 760.950 574.050 763.050 ;
        RECT 580.950 762.750 583.050 763.200 ;
        RECT 589.950 762.750 592.050 763.200 ;
        RECT 580.950 761.550 592.050 762.750 ;
        RECT 580.950 761.100 583.050 761.550 ;
        RECT 589.950 761.100 592.050 761.550 ;
        RECT 595.950 761.100 598.050 763.200 ;
        RECT 601.950 762.600 604.050 763.200 ;
        RECT 619.950 762.750 622.050 763.200 ;
        RECT 625.950 762.750 628.050 763.200 ;
        RECT 601.950 761.400 609.600 762.600 ;
        RECT 601.950 761.100 604.050 761.400 ;
        RECT 469.950 756.600 472.050 756.900 ;
        RECT 455.400 755.400 472.050 756.600 ;
        RECT 473.400 755.400 477.900 757.050 ;
        RECT 479.400 756.900 480.600 760.950 ;
        RECT 415.950 754.800 418.050 755.250 ;
        RECT 421.950 754.800 424.050 755.250 ;
        RECT 451.950 754.800 454.050 755.400 ;
        RECT 469.950 754.800 472.050 755.400 ;
        RECT 474.000 754.950 477.900 755.400 ;
        RECT 478.950 754.800 481.050 756.900 ;
        RECT 508.950 756.600 511.050 757.050 ;
        RECT 568.950 756.600 571.050 757.050 ;
        RECT 508.950 755.400 571.050 756.600 ;
        RECT 572.400 756.600 573.600 760.950 ;
        RECT 577.950 756.600 580.050 756.900 ;
        RECT 572.400 755.400 580.050 756.600 ;
        RECT 508.950 754.950 511.050 755.400 ;
        RECT 568.950 754.950 571.050 755.400 ;
        RECT 577.950 754.800 580.050 755.400 ;
        RECT 586.950 756.600 589.050 757.050 ;
        RECT 596.400 756.600 597.600 761.100 ;
        RECT 608.400 756.900 609.600 761.400 ;
        RECT 619.950 761.550 628.050 762.750 ;
        RECT 619.950 761.100 622.050 761.550 ;
        RECT 625.950 761.100 628.050 761.550 ;
        RECT 649.950 761.100 652.050 763.200 ;
        RECT 655.950 761.100 658.050 763.200 ;
        RECT 664.950 762.600 667.050 763.050 ;
        RECT 673.950 762.600 676.050 763.200 ;
        RECT 664.950 761.400 676.050 762.600 ;
        RECT 586.950 755.400 597.600 756.600 ;
        RECT 586.950 754.950 589.050 755.400 ;
        RECT 607.950 754.800 610.050 756.900 ;
        RECT 121.950 753.600 124.050 754.050 ;
        RECT 133.950 753.600 136.050 754.050 ;
        RECT 121.950 752.400 136.050 753.600 ;
        RECT 121.950 751.950 124.050 752.400 ;
        RECT 133.950 751.950 136.050 752.400 ;
        RECT 148.950 753.600 151.050 754.050 ;
        RECT 157.950 753.600 160.050 754.050 ;
        RECT 148.950 752.400 160.050 753.600 ;
        RECT 148.950 751.950 151.050 752.400 ;
        RECT 157.950 751.950 160.050 752.400 ;
        RECT 169.950 753.600 172.050 754.050 ;
        RECT 181.950 753.600 184.050 754.050 ;
        RECT 169.950 752.400 184.050 753.600 ;
        RECT 169.950 751.950 172.050 752.400 ;
        RECT 181.950 751.950 184.050 752.400 ;
        RECT 247.950 753.600 250.050 754.050 ;
        RECT 274.950 753.600 277.050 754.050 ;
        RECT 247.950 752.400 277.050 753.600 ;
        RECT 247.950 751.950 250.050 752.400 ;
        RECT 274.950 751.950 277.050 752.400 ;
        RECT 430.950 753.600 433.050 754.050 ;
        RECT 439.950 753.600 442.050 754.050 ;
        RECT 430.950 752.400 442.050 753.600 ;
        RECT 430.950 751.950 433.050 752.400 ;
        RECT 439.950 751.950 442.050 752.400 ;
        RECT 598.950 753.600 601.050 754.050 ;
        RECT 604.950 753.600 607.050 754.050 ;
        RECT 598.950 752.400 607.050 753.600 ;
        RECT 598.950 751.950 601.050 752.400 ;
        RECT 604.950 751.950 607.050 752.400 ;
        RECT 610.950 753.600 613.050 754.050 ;
        RECT 650.400 753.600 651.600 761.100 ;
        RECT 610.950 752.400 651.600 753.600 ;
        RECT 610.950 751.950 613.050 752.400 ;
        RECT 28.950 750.600 31.050 751.050 ;
        RECT 37.950 750.600 40.050 751.050 ;
        RECT 28.950 749.400 40.050 750.600 ;
        RECT 28.950 748.950 31.050 749.400 ;
        RECT 37.950 748.950 40.050 749.400 ;
        RECT 103.950 750.600 106.050 751.050 ;
        RECT 118.950 750.600 121.050 751.050 ;
        RECT 103.950 749.400 121.050 750.600 ;
        RECT 103.950 748.950 106.050 749.400 ;
        RECT 118.950 748.950 121.050 749.400 ;
        RECT 211.950 750.600 214.050 751.050 ;
        RECT 250.950 750.600 253.050 751.050 ;
        RECT 211.950 749.400 253.050 750.600 ;
        RECT 211.950 748.950 214.050 749.400 ;
        RECT 250.950 748.950 253.050 749.400 ;
        RECT 337.950 750.600 340.050 751.050 ;
        RECT 364.950 750.600 367.050 751.050 ;
        RECT 337.950 749.400 367.050 750.600 ;
        RECT 337.950 748.950 340.050 749.400 ;
        RECT 364.950 748.950 367.050 749.400 ;
        RECT 370.950 750.600 373.050 751.050 ;
        RECT 397.950 750.600 400.050 751.050 ;
        RECT 370.950 749.400 400.050 750.600 ;
        RECT 370.950 748.950 373.050 749.400 ;
        RECT 397.950 748.950 400.050 749.400 ;
        RECT 409.950 750.600 412.050 751.050 ;
        RECT 418.950 750.600 421.050 751.050 ;
        RECT 409.950 749.400 421.050 750.600 ;
        RECT 409.950 748.950 412.050 749.400 ;
        RECT 418.950 748.950 421.050 749.400 ;
        RECT 493.950 750.600 496.050 751.050 ;
        RECT 541.950 750.600 544.050 751.050 ;
        RECT 493.950 749.400 544.050 750.600 ;
        RECT 493.950 748.950 496.050 749.400 ;
        RECT 541.950 748.950 544.050 749.400 ;
        RECT 589.950 750.600 592.050 751.050 ;
        RECT 607.950 750.600 610.050 751.050 ;
        RECT 589.950 749.400 610.050 750.600 ;
        RECT 589.950 748.950 592.050 749.400 ;
        RECT 607.950 748.950 610.050 749.400 ;
        RECT 619.950 750.600 622.050 751.050 ;
        RECT 652.950 750.600 655.050 751.050 ;
        RECT 619.950 749.400 655.050 750.600 ;
        RECT 656.400 750.600 657.600 761.100 ;
        RECT 664.950 760.950 667.050 761.400 ;
        RECT 673.950 761.100 676.050 761.400 ;
        RECT 697.950 762.750 700.050 763.200 ;
        RECT 706.950 762.750 709.050 763.200 ;
        RECT 697.950 761.550 709.050 762.750 ;
        RECT 697.950 761.100 700.050 761.550 ;
        RECT 706.950 761.100 709.050 761.550 ;
        RECT 721.950 762.600 724.050 763.050 ;
        RECT 727.950 762.600 730.050 763.200 ;
        RECT 742.950 762.600 745.050 763.200 ;
        RECT 721.950 761.400 730.050 762.600 ;
        RECT 721.950 760.950 724.050 761.400 ;
        RECT 727.950 761.100 730.050 761.400 ;
        RECT 740.400 761.400 745.050 762.600 ;
        RECT 740.400 757.050 741.600 761.400 ;
        RECT 742.950 761.100 745.050 761.400 ;
        RECT 760.950 761.100 763.050 763.200 ;
        RECT 766.950 762.600 769.050 763.200 ;
        RECT 781.950 762.600 784.050 763.200 ;
        RECT 766.950 761.400 784.050 762.600 ;
        RECT 766.950 761.100 769.050 761.400 ;
        RECT 781.950 761.100 784.050 761.400 ;
        RECT 790.950 762.600 793.050 763.050 ;
        RECT 799.950 762.600 802.050 763.200 ;
        RECT 790.950 761.400 802.050 762.600 ;
        RECT 761.400 759.600 762.600 761.100 ;
        RECT 790.950 760.950 793.050 761.400 ;
        RECT 799.950 761.100 802.050 761.400 ;
        RECT 808.950 762.750 811.050 763.200 ;
        RECT 823.950 762.750 826.050 763.200 ;
        RECT 808.950 761.550 826.050 762.750 ;
        RECT 808.950 761.100 811.050 761.550 ;
        RECT 823.950 761.100 826.050 761.550 ;
        RECT 829.950 761.100 832.050 763.200 ;
        RECT 838.950 762.600 841.050 763.200 ;
        RECT 847.950 762.600 850.050 763.050 ;
        RECT 838.950 761.400 850.050 762.600 ;
        RECT 838.950 761.100 841.050 761.400 ;
        RECT 761.400 759.000 777.600 759.600 ;
        RECT 761.400 758.400 778.050 759.000 ;
        RECT 685.950 756.600 688.050 757.050 ;
        RECT 700.950 756.600 703.050 757.050 ;
        RECT 685.950 755.400 703.050 756.600 ;
        RECT 685.950 754.950 688.050 755.400 ;
        RECT 700.950 754.950 703.050 755.400 ;
        RECT 715.950 756.450 718.050 756.900 ;
        RECT 721.950 756.450 724.050 756.900 ;
        RECT 715.950 755.250 724.050 756.450 ;
        RECT 715.950 754.800 718.050 755.250 ;
        RECT 721.950 754.800 724.050 755.250 ;
        RECT 730.950 756.450 733.050 756.900 ;
        RECT 736.800 756.450 738.900 756.900 ;
        RECT 730.950 755.250 738.900 756.450 ;
        RECT 730.950 754.800 733.050 755.250 ;
        RECT 736.800 754.800 738.900 755.250 ;
        RECT 739.950 754.950 742.050 757.050 ;
        RECT 745.950 756.450 748.050 756.900 ;
        RECT 751.950 756.450 754.050 756.900 ;
        RECT 745.950 755.250 754.050 756.450 ;
        RECT 745.950 754.800 748.050 755.250 ;
        RECT 751.950 754.800 754.050 755.250 ;
        RECT 763.950 756.450 766.050 756.900 ;
        RECT 772.800 756.450 774.900 756.900 ;
        RECT 763.950 755.250 774.900 756.450 ;
        RECT 763.950 754.800 766.050 755.250 ;
        RECT 772.800 754.800 774.900 755.250 ;
        RECT 775.950 754.950 778.050 758.400 ;
        RECT 784.950 756.450 787.050 756.900 ;
        RECT 790.950 756.450 793.050 756.900 ;
        RECT 784.950 755.250 793.050 756.450 ;
        RECT 784.950 754.800 787.050 755.250 ;
        RECT 790.950 754.800 793.050 755.250 ;
        RECT 823.950 753.600 826.050 754.050 ;
        RECT 830.400 753.600 831.600 761.100 ;
        RECT 847.950 760.950 850.050 761.400 ;
        RECT 823.950 752.400 831.600 753.600 ;
        RECT 823.950 751.950 826.050 752.400 ;
        RECT 709.950 750.600 712.050 751.050 ;
        RECT 656.400 749.400 712.050 750.600 ;
        RECT 619.950 748.950 622.050 749.400 ;
        RECT 652.950 748.950 655.050 749.400 ;
        RECT 709.950 748.950 712.050 749.400 ;
        RECT 736.950 750.600 739.050 751.050 ;
        RECT 814.950 750.600 817.050 751.050 ;
        RECT 736.950 749.400 817.050 750.600 ;
        RECT 736.950 748.950 739.050 749.400 ;
        RECT 814.950 748.950 817.050 749.400 ;
        RECT 820.950 750.600 823.050 751.050 ;
        RECT 847.950 750.600 850.050 751.050 ;
        RECT 820.950 749.400 850.050 750.600 ;
        RECT 820.950 748.950 823.050 749.400 ;
        RECT 847.950 748.950 850.050 749.400 ;
        RECT 61.950 747.600 64.050 748.050 ;
        RECT 97.950 747.600 100.050 748.050 ;
        RECT 127.950 747.600 130.050 748.050 ;
        RECT 61.950 746.400 130.050 747.600 ;
        RECT 61.950 745.950 64.050 746.400 ;
        RECT 97.950 745.950 100.050 746.400 ;
        RECT 127.950 745.950 130.050 746.400 ;
        RECT 139.950 747.600 142.050 748.050 ;
        RECT 184.950 747.600 187.050 748.050 ;
        RECT 139.950 746.400 187.050 747.600 ;
        RECT 139.950 745.950 142.050 746.400 ;
        RECT 184.950 745.950 187.050 746.400 ;
        RECT 478.950 747.600 481.050 748.050 ;
        RECT 487.950 747.600 490.050 748.050 ;
        RECT 478.950 746.400 490.050 747.600 ;
        RECT 478.950 745.950 481.050 746.400 ;
        RECT 487.950 745.950 490.050 746.400 ;
        RECT 784.950 747.600 787.050 748.050 ;
        RECT 790.950 747.600 793.050 748.050 ;
        RECT 802.950 747.600 805.050 748.050 ;
        RECT 784.950 746.400 805.050 747.600 ;
        RECT 784.950 745.950 787.050 746.400 ;
        RECT 790.950 745.950 793.050 746.400 ;
        RECT 802.950 745.950 805.050 746.400 ;
        RECT 106.950 744.600 109.050 745.050 ;
        RECT 112.950 744.600 115.050 745.050 ;
        RECT 106.950 743.400 115.050 744.600 ;
        RECT 106.950 742.950 109.050 743.400 ;
        RECT 112.950 742.950 115.050 743.400 ;
        RECT 145.950 744.600 148.050 745.050 ;
        RECT 178.950 744.600 181.050 745.050 ;
        RECT 145.950 743.400 181.050 744.600 ;
        RECT 145.950 742.950 148.050 743.400 ;
        RECT 178.950 742.950 181.050 743.400 ;
        RECT 214.950 744.600 217.050 745.050 ;
        RECT 247.950 744.600 250.050 745.050 ;
        RECT 214.950 743.400 250.050 744.600 ;
        RECT 214.950 742.950 217.050 743.400 ;
        RECT 247.950 742.950 250.050 743.400 ;
        RECT 376.950 744.600 379.050 745.050 ;
        RECT 394.950 744.600 397.050 745.050 ;
        RECT 376.950 743.400 397.050 744.600 ;
        RECT 376.950 742.950 379.050 743.400 ;
        RECT 394.950 742.950 397.050 743.400 ;
        RECT 412.950 744.600 415.050 745.050 ;
        RECT 460.950 744.600 463.050 745.050 ;
        RECT 412.950 743.400 463.050 744.600 ;
        RECT 412.950 742.950 415.050 743.400 ;
        RECT 460.950 742.950 463.050 743.400 ;
        RECT 541.950 744.600 544.050 745.050 ;
        RECT 559.950 744.600 562.050 745.050 ;
        RECT 541.950 743.400 562.050 744.600 ;
        RECT 541.950 742.950 544.050 743.400 ;
        RECT 559.950 742.950 562.050 743.400 ;
        RECT 676.950 744.600 679.050 745.050 ;
        RECT 757.950 744.600 760.050 745.050 ;
        RECT 676.950 743.400 760.050 744.600 ;
        RECT 676.950 742.950 679.050 743.400 ;
        RECT 757.950 742.950 760.050 743.400 ;
        RECT 808.950 744.600 811.050 745.050 ;
        RECT 820.950 744.600 823.050 745.050 ;
        RECT 808.950 743.400 823.050 744.600 ;
        RECT 808.950 742.950 811.050 743.400 ;
        RECT 820.950 742.950 823.050 743.400 ;
        RECT 13.950 741.600 16.050 742.050 ;
        RECT 31.950 741.600 34.050 742.050 ;
        RECT 73.950 741.600 76.050 742.050 ;
        RECT 142.950 741.600 145.050 742.050 ;
        RECT 211.950 741.600 214.050 742.050 ;
        RECT 13.950 740.400 214.050 741.600 ;
        RECT 13.950 739.950 16.050 740.400 ;
        RECT 31.950 739.950 34.050 740.400 ;
        RECT 73.950 739.950 76.050 740.400 ;
        RECT 142.950 739.950 145.050 740.400 ;
        RECT 211.950 739.950 214.050 740.400 ;
        RECT 250.950 741.600 253.050 742.050 ;
        RECT 445.950 741.600 448.050 742.050 ;
        RECT 250.950 740.400 448.050 741.600 ;
        RECT 250.950 739.950 253.050 740.400 ;
        RECT 445.950 739.950 448.050 740.400 ;
        RECT 697.950 741.600 700.050 742.050 ;
        RECT 736.950 741.600 739.050 742.050 ;
        RECT 697.950 740.400 739.050 741.600 ;
        RECT 697.950 739.950 700.050 740.400 ;
        RECT 736.950 739.950 739.050 740.400 ;
        RECT 106.950 738.600 109.050 739.050 ;
        RECT 169.950 738.600 172.050 739.050 ;
        RECT 106.950 737.400 172.050 738.600 ;
        RECT 106.950 736.950 109.050 737.400 ;
        RECT 169.950 736.950 172.050 737.400 ;
        RECT 289.950 738.600 292.050 739.050 ;
        RECT 304.800 738.600 306.900 739.050 ;
        RECT 289.950 737.400 306.900 738.600 ;
        RECT 289.950 736.950 292.050 737.400 ;
        RECT 304.800 736.950 306.900 737.400 ;
        RECT 307.950 738.600 310.050 739.050 ;
        RECT 313.950 738.600 316.050 739.050 ;
        RECT 307.950 737.400 316.050 738.600 ;
        RECT 307.950 736.950 310.050 737.400 ;
        RECT 313.950 736.950 316.050 737.400 ;
        RECT 328.950 738.600 331.050 739.050 ;
        RECT 334.950 738.600 337.050 739.050 ;
        RECT 370.950 738.600 373.050 739.050 ;
        RECT 328.950 737.400 373.050 738.600 ;
        RECT 328.950 736.950 331.050 737.400 ;
        RECT 334.950 736.950 337.050 737.400 ;
        RECT 370.950 736.950 373.050 737.400 ;
        RECT 469.950 738.600 472.050 739.050 ;
        RECT 481.950 738.600 484.050 739.050 ;
        RECT 469.950 737.400 484.050 738.600 ;
        RECT 469.950 736.950 472.050 737.400 ;
        RECT 481.950 736.950 484.050 737.400 ;
        RECT 670.950 738.600 673.050 739.050 ;
        RECT 682.950 738.600 685.050 739.050 ;
        RECT 688.950 738.600 691.050 739.050 ;
        RECT 670.950 737.400 691.050 738.600 ;
        RECT 670.950 736.950 673.050 737.400 ;
        RECT 682.950 736.950 685.050 737.400 ;
        RECT 688.950 736.950 691.050 737.400 ;
        RECT 748.950 738.600 751.050 739.050 ;
        RECT 796.950 738.600 799.050 739.050 ;
        RECT 748.950 737.400 799.050 738.600 ;
        RECT 748.950 736.950 751.050 737.400 ;
        RECT 796.950 736.950 799.050 737.400 ;
        RECT 856.950 738.600 859.050 739.050 ;
        RECT 874.950 738.600 877.050 739.050 ;
        RECT 856.950 737.400 877.050 738.600 ;
        RECT 856.950 736.950 859.050 737.400 ;
        RECT 874.950 736.950 877.050 737.400 ;
        RECT 34.950 735.600 37.050 736.050 ;
        RECT 40.950 735.600 43.050 736.050 ;
        RECT 46.950 735.600 49.050 736.050 ;
        RECT 34.950 734.400 49.050 735.600 ;
        RECT 34.950 733.950 37.050 734.400 ;
        RECT 40.950 733.950 43.050 734.400 ;
        RECT 46.950 733.950 49.050 734.400 ;
        RECT 172.950 735.600 175.050 736.050 ;
        RECT 193.950 735.600 196.050 736.050 ;
        RECT 172.950 734.400 196.050 735.600 ;
        RECT 172.950 733.950 175.050 734.400 ;
        RECT 193.950 733.950 196.050 734.400 ;
        RECT 199.950 735.600 202.050 736.050 ;
        RECT 223.950 735.600 226.050 736.050 ;
        RECT 199.950 734.400 226.050 735.600 ;
        RECT 199.950 733.950 202.050 734.400 ;
        RECT 223.950 733.950 226.050 734.400 ;
        RECT 238.950 735.600 241.050 736.050 ;
        RECT 250.950 735.600 253.050 736.050 ;
        RECT 349.950 735.600 352.050 736.050 ;
        RECT 361.950 735.600 364.050 736.050 ;
        RECT 238.950 734.400 276.600 735.600 ;
        RECT 238.950 733.950 241.050 734.400 ;
        RECT 250.950 733.950 253.050 734.400 ;
        RECT 275.400 733.050 276.600 734.400 ;
        RECT 349.950 734.400 364.050 735.600 ;
        RECT 349.950 733.950 352.050 734.400 ;
        RECT 361.950 733.950 364.050 734.400 ;
        RECT 403.950 735.600 406.050 736.050 ;
        RECT 433.950 735.600 436.050 736.050 ;
        RECT 403.950 734.400 436.050 735.600 ;
        RECT 403.950 733.950 406.050 734.400 ;
        RECT 433.950 733.950 436.050 734.400 ;
        RECT 442.950 735.600 445.050 736.050 ;
        RECT 460.950 735.600 463.050 736.050 ;
        RECT 442.950 734.400 463.050 735.600 ;
        RECT 442.950 733.950 445.050 734.400 ;
        RECT 460.950 733.950 463.050 734.400 ;
        RECT 466.950 735.600 469.050 736.050 ;
        RECT 487.950 735.600 490.050 736.050 ;
        RECT 466.950 734.400 490.050 735.600 ;
        RECT 466.950 733.950 469.050 734.400 ;
        RECT 487.950 733.950 490.050 734.400 ;
        RECT 529.950 735.600 532.050 736.050 ;
        RECT 559.950 735.600 562.050 736.050 ;
        RECT 529.950 734.400 562.050 735.600 ;
        RECT 529.950 733.950 532.050 734.400 ;
        RECT 559.950 733.950 562.050 734.400 ;
        RECT 691.950 735.600 694.050 736.050 ;
        RECT 703.950 735.600 706.050 736.050 ;
        RECT 691.950 734.400 706.050 735.600 ;
        RECT 691.950 733.950 694.050 734.400 ;
        RECT 703.950 733.950 706.050 734.400 ;
        RECT 715.950 735.600 718.050 736.050 ;
        RECT 739.950 735.600 742.050 736.050 ;
        RECT 715.950 734.400 742.050 735.600 ;
        RECT 715.950 733.950 718.050 734.400 ;
        RECT 739.950 733.950 742.050 734.400 ;
        RECT 757.950 735.600 760.050 736.050 ;
        RECT 769.950 735.600 772.050 736.050 ;
        RECT 757.950 734.400 772.050 735.600 ;
        RECT 757.950 733.950 760.050 734.400 ;
        RECT 769.950 733.950 772.050 734.400 ;
        RECT 832.950 735.600 835.050 736.050 ;
        RECT 853.950 735.600 856.050 736.050 ;
        RECT 832.950 734.400 856.050 735.600 ;
        RECT 832.950 733.950 835.050 734.400 ;
        RECT 853.950 733.950 856.050 734.400 ;
        RECT 85.950 732.600 88.050 733.050 ;
        RECT 112.950 732.600 115.050 733.050 ;
        RECT 85.950 731.400 115.050 732.600 ;
        RECT 85.950 730.950 88.050 731.400 ;
        RECT 112.950 730.950 115.050 731.400 ;
        RECT 124.950 732.600 127.050 733.050 ;
        RECT 133.950 732.600 136.050 733.050 ;
        RECT 166.950 732.600 169.050 733.050 ;
        RECT 124.950 731.400 169.050 732.600 ;
        RECT 124.950 730.950 127.050 731.400 ;
        RECT 133.950 730.950 136.050 731.400 ;
        RECT 166.950 730.950 169.050 731.400 ;
        RECT 274.950 732.600 277.050 733.050 ;
        RECT 286.950 732.600 289.050 733.050 ;
        RECT 274.950 731.400 289.050 732.600 ;
        RECT 274.950 730.950 277.050 731.400 ;
        RECT 286.950 730.950 289.050 731.400 ;
        RECT 382.950 732.600 385.050 733.050 ;
        RECT 388.950 732.600 391.050 733.050 ;
        RECT 382.950 731.400 391.050 732.600 ;
        RECT 382.950 730.950 385.050 731.400 ;
        RECT 388.950 730.950 391.050 731.400 ;
        RECT 493.950 732.600 496.050 733.050 ;
        RECT 499.950 732.600 502.050 733.050 ;
        RECT 493.950 731.400 502.050 732.600 ;
        RECT 493.950 730.950 496.050 731.400 ;
        RECT 499.950 730.950 502.050 731.400 ;
        RECT 532.950 732.600 535.050 733.050 ;
        RECT 538.800 732.600 540.900 733.050 ;
        RECT 532.950 731.400 540.900 732.600 ;
        RECT 532.950 730.950 535.050 731.400 ;
        RECT 538.800 730.950 540.900 731.400 ;
        RECT 7.950 727.950 10.050 730.050 ;
        RECT 13.950 729.600 16.050 730.200 ;
        RECT 22.950 729.600 25.050 730.050 ;
        RECT 13.950 728.400 25.050 729.600 ;
        RECT 13.950 728.100 16.050 728.400 ;
        RECT 22.950 727.950 25.050 728.400 ;
        RECT 28.950 729.600 31.050 730.200 ;
        RECT 46.950 729.600 49.050 730.200 ;
        RECT 28.950 728.400 49.050 729.600 ;
        RECT 28.950 728.100 31.050 728.400 ;
        RECT 46.950 728.100 49.050 728.400 ;
        RECT 52.950 729.600 55.050 730.200 ;
        RECT 61.950 729.600 64.050 730.050 ;
        RECT 52.950 728.400 64.050 729.600 ;
        RECT 52.950 728.100 55.050 728.400 ;
        RECT 8.400 724.050 9.600 727.950 ;
        RECT 47.400 726.600 48.600 728.100 ;
        RECT 61.950 727.950 64.050 728.400 ;
        RECT 91.950 728.100 94.050 730.200 ;
        RECT 181.950 729.750 184.050 730.200 ;
        RECT 187.950 729.750 190.050 730.200 ;
        RECT 181.950 728.550 190.050 729.750 ;
        RECT 181.950 728.100 184.050 728.550 ;
        RECT 187.950 728.100 190.050 728.550 ;
        RECT 214.950 728.100 217.050 730.200 ;
        RECT 256.950 729.600 259.050 730.200 ;
        RECT 265.950 729.600 268.050 730.050 ;
        RECT 256.950 728.400 268.050 729.600 ;
        RECT 256.950 728.100 259.050 728.400 ;
        RECT 47.400 725.400 72.600 726.600 ;
        RECT 7.950 721.950 10.050 724.050 ;
        RECT 40.950 723.450 43.050 723.900 ;
        RECT 49.950 723.450 52.050 723.900 ;
        RECT 40.950 722.250 52.050 723.450 ;
        RECT 40.950 721.800 43.050 722.250 ;
        RECT 49.950 721.800 52.050 722.250 ;
        RECT 61.950 723.450 64.050 723.900 ;
        RECT 67.950 723.450 70.050 723.900 ;
        RECT 61.950 722.250 70.050 723.450 ;
        RECT 71.400 723.600 72.600 725.400 ;
        RECT 88.950 723.600 91.050 723.900 ;
        RECT 71.400 722.400 91.050 723.600 ;
        RECT 92.400 723.600 93.600 728.100 ;
        RECT 109.950 723.600 112.050 723.900 ;
        RECT 124.950 723.600 127.050 723.900 ;
        RECT 92.400 722.400 127.050 723.600 ;
        RECT 61.950 721.800 64.050 722.250 ;
        RECT 67.950 721.800 70.050 722.250 ;
        RECT 88.950 721.800 91.050 722.400 ;
        RECT 109.950 721.800 112.050 722.400 ;
        RECT 124.950 721.800 127.050 722.400 ;
        RECT 178.950 723.600 181.050 723.900 ;
        RECT 196.950 723.600 199.050 723.900 ;
        RECT 178.950 722.400 199.050 723.600 ;
        RECT 215.400 723.600 216.600 728.100 ;
        RECT 265.950 727.950 268.050 728.400 ;
        RECT 343.950 728.100 346.050 730.200 ;
        RECT 355.950 729.750 358.050 730.200 ;
        RECT 370.950 729.750 373.050 730.200 ;
        RECT 355.950 728.550 373.050 729.750 ;
        RECT 379.950 729.600 382.050 730.200 ;
        RECT 424.950 729.600 427.050 730.200 ;
        RECT 355.950 728.100 358.050 728.550 ;
        RECT 370.950 728.100 373.050 728.550 ;
        RECT 374.400 728.400 382.050 729.600 ;
        RECT 288.000 726.600 292.050 727.050 ;
        RECT 287.400 724.950 292.050 726.600 ;
        RECT 220.950 723.600 223.050 724.050 ;
        RECT 215.400 722.400 223.050 723.600 ;
        RECT 178.950 721.800 181.050 722.400 ;
        RECT 196.950 721.800 199.050 722.400 ;
        RECT 220.950 721.950 223.050 722.400 ;
        RECT 259.950 723.600 262.050 723.900 ;
        RECT 287.400 723.600 288.600 724.950 ;
        RECT 259.950 722.400 288.600 723.600 ;
        RECT 334.950 723.450 337.050 723.900 ;
        RECT 340.950 723.450 343.050 723.900 ;
        RECT 259.950 721.800 262.050 722.400 ;
        RECT 334.950 722.250 343.050 723.450 ;
        RECT 344.400 723.600 345.600 728.100 ;
        RECT 374.400 726.600 375.600 728.400 ;
        RECT 379.950 728.100 382.050 728.400 ;
        RECT 410.400 728.400 427.050 729.600 ;
        RECT 365.400 725.400 375.600 726.600 ;
        RECT 365.400 723.900 366.600 725.400 ;
        RECT 410.400 723.900 411.600 728.400 ;
        RECT 424.950 728.100 427.050 728.400 ;
        RECT 436.950 729.600 439.050 730.050 ;
        RECT 451.950 729.600 454.050 730.200 ;
        RECT 436.950 728.400 454.050 729.600 ;
        RECT 436.950 727.950 439.050 728.400 ;
        RECT 451.950 728.100 454.050 728.400 ;
        RECT 457.950 729.600 460.050 730.200 ;
        RECT 463.950 729.600 466.050 730.050 ;
        RECT 469.950 729.600 472.050 730.200 ;
        RECT 457.950 728.400 466.050 729.600 ;
        RECT 457.950 728.100 460.050 728.400 ;
        RECT 463.950 727.950 466.050 728.400 ;
        RECT 467.400 728.400 472.050 729.600 ;
        RECT 344.400 722.400 354.600 723.600 ;
        RECT 334.950 721.800 337.050 722.250 ;
        RECT 340.950 721.800 343.050 722.250 ;
        RECT 22.950 717.600 25.050 718.050 ;
        RECT 73.950 717.600 76.050 718.050 ;
        RECT 103.950 717.600 106.050 718.050 ;
        RECT 22.950 716.400 106.050 717.600 ;
        RECT 151.950 717.600 154.050 721.050 ;
        RECT 217.950 720.600 220.050 721.050 ;
        RECT 235.950 720.600 238.050 721.050 ;
        RECT 253.950 720.600 256.050 721.050 ;
        RECT 217.950 719.400 256.050 720.600 ;
        RECT 217.950 718.950 220.050 719.400 ;
        RECT 235.950 718.950 238.050 719.400 ;
        RECT 253.950 718.950 256.050 719.400 ;
        RECT 265.950 720.600 268.050 721.050 ;
        RECT 289.950 720.600 292.050 721.050 ;
        RECT 265.950 719.400 292.050 720.600 ;
        RECT 353.400 720.600 354.600 722.400 ;
        RECT 364.950 721.800 367.050 723.900 ;
        RECT 409.950 721.800 412.050 723.900 ;
        RECT 433.950 723.450 436.050 723.900 ;
        RECT 442.950 723.450 445.050 723.900 ;
        RECT 433.950 722.250 445.050 723.450 ;
        RECT 433.950 721.800 436.050 722.250 ;
        RECT 442.950 721.800 445.050 722.250 ;
        RECT 454.950 723.600 457.050 723.900 ;
        RECT 467.400 723.600 468.600 728.400 ;
        RECT 469.950 728.100 472.050 728.400 ;
        RECT 475.950 727.950 478.050 730.050 ;
        RECT 487.950 729.600 490.050 730.200 ;
        RECT 514.950 729.600 517.050 730.200 ;
        RECT 541.950 729.600 544.050 733.050 ;
        RECT 565.950 732.600 568.050 733.050 ;
        RECT 583.950 732.600 586.050 733.050 ;
        RECT 565.950 731.400 586.050 732.600 ;
        RECT 565.950 730.950 568.050 731.400 ;
        RECT 583.950 730.950 586.050 731.400 ;
        RECT 667.950 732.600 670.050 733.050 ;
        RECT 685.950 732.600 688.050 733.050 ;
        RECT 667.950 731.400 688.050 732.600 ;
        RECT 667.950 730.950 670.050 731.400 ;
        RECT 685.950 730.950 688.050 731.400 ;
        RECT 709.950 732.600 712.050 733.050 ;
        RECT 721.950 732.600 724.050 733.050 ;
        RECT 709.950 731.400 724.050 732.600 ;
        RECT 709.950 730.950 712.050 731.400 ;
        RECT 721.950 730.950 724.050 731.400 ;
        RECT 547.950 729.600 550.050 730.200 ;
        RECT 487.950 728.400 510.600 729.600 ;
        RECT 487.950 728.100 490.050 728.400 ;
        RECT 476.400 724.050 477.600 727.950 ;
        RECT 509.400 726.600 510.600 728.400 ;
        RECT 514.950 728.400 519.600 729.600 ;
        RECT 541.950 729.000 550.050 729.600 ;
        RECT 542.400 728.400 550.050 729.000 ;
        RECT 514.950 728.100 517.050 728.400 ;
        RECT 509.400 725.400 513.600 726.600 ;
        RECT 454.950 722.400 468.600 723.600 ;
        RECT 454.950 721.800 457.050 722.400 ;
        RECT 475.950 721.950 478.050 724.050 ;
        RECT 481.950 723.600 484.050 724.050 ;
        RECT 512.400 723.900 513.600 725.400 ;
        RECT 490.950 723.600 493.050 723.900 ;
        RECT 481.950 722.400 493.050 723.600 ;
        RECT 481.950 721.950 484.050 722.400 ;
        RECT 490.950 721.800 493.050 722.400 ;
        RECT 511.950 721.800 514.050 723.900 ;
        RECT 394.950 720.600 397.050 721.050 ;
        RECT 353.400 719.400 397.050 720.600 ;
        RECT 265.950 718.950 268.050 719.400 ;
        RECT 289.950 718.950 292.050 719.400 ;
        RECT 394.950 718.950 397.050 719.400 ;
        RECT 427.950 720.600 430.050 721.050 ;
        RECT 448.950 720.600 451.050 721.050 ;
        RECT 427.950 719.400 451.050 720.600 ;
        RECT 427.950 718.950 430.050 719.400 ;
        RECT 448.950 718.950 451.050 719.400 ;
        RECT 466.950 720.600 469.050 721.050 ;
        RECT 472.950 720.600 475.050 721.050 ;
        RECT 466.950 719.400 475.050 720.600 ;
        RECT 518.400 720.600 519.600 728.400 ;
        RECT 547.950 728.100 550.050 728.400 ;
        RECT 553.950 728.100 556.050 730.200 ;
        RECT 568.950 729.600 571.050 730.200 ;
        RECT 574.950 729.600 577.050 730.200 ;
        RECT 568.950 728.400 577.050 729.600 ;
        RECT 568.950 728.100 571.050 728.400 ;
        RECT 574.950 728.100 577.050 728.400 ;
        RECT 622.950 729.600 625.050 730.050 ;
        RECT 652.950 729.600 655.050 730.200 ;
        RECT 622.950 728.400 655.050 729.600 ;
        RECT 520.950 726.600 523.050 727.050 ;
        RECT 554.400 726.600 555.600 728.100 ;
        RECT 622.950 727.950 625.050 728.400 ;
        RECT 652.950 728.100 655.050 728.400 ;
        RECT 658.950 728.100 661.050 730.200 ;
        RECT 739.950 729.600 742.050 730.050 ;
        RECT 763.950 729.600 766.050 730.200 ;
        RECT 850.950 729.600 853.050 730.200 ;
        RECT 856.950 729.600 859.050 732.900 ;
        RECT 739.950 728.400 801.600 729.600 ;
        RECT 520.950 725.400 555.600 726.600 ;
        RECT 583.950 726.600 586.050 727.050 ;
        RECT 659.400 726.600 660.600 728.100 ;
        RECT 739.950 727.950 742.050 728.400 ;
        RECT 763.950 728.100 766.050 728.400 ;
        RECT 583.950 725.400 603.600 726.600 ;
        RECT 659.400 725.400 699.600 726.600 ;
        RECT 520.950 724.950 523.050 725.400 ;
        RECT 583.950 724.950 586.050 725.400 ;
        RECT 544.950 723.600 547.050 723.900 ;
        RECT 562.950 723.600 565.050 724.050 ;
        RECT 602.400 723.900 603.600 725.400 ;
        RECT 698.400 724.050 699.600 725.400 ;
        RECT 544.950 722.400 565.050 723.600 ;
        RECT 544.950 721.800 547.050 722.400 ;
        RECT 562.950 721.950 565.050 722.400 ;
        RECT 601.950 721.800 604.050 723.900 ;
        RECT 637.950 723.600 640.050 723.900 ;
        RECT 643.950 723.600 646.050 724.050 ;
        RECT 637.950 722.400 646.050 723.600 ;
        RECT 698.400 722.400 702.900 724.050 ;
        RECT 637.950 721.800 640.050 722.400 ;
        RECT 643.950 721.950 646.050 722.400 ;
        RECT 699.000 721.950 702.900 722.400 ;
        RECT 703.950 723.600 706.050 724.050 ;
        RECT 730.950 723.600 733.050 723.900 ;
        RECT 703.950 722.400 733.050 723.600 ;
        RECT 703.950 721.950 706.050 722.400 ;
        RECT 730.950 721.800 733.050 722.400 ;
        RECT 766.950 723.600 769.050 723.900 ;
        RECT 775.950 723.600 778.050 724.050 ;
        RECT 800.400 723.900 801.600 728.400 ;
        RECT 850.950 729.000 859.050 729.600 ;
        RECT 850.950 728.400 858.600 729.000 ;
        RECT 850.950 728.100 853.050 728.400 ;
        RECT 766.950 722.400 778.050 723.600 ;
        RECT 766.950 721.800 769.050 722.400 ;
        RECT 775.950 721.950 778.050 722.400 ;
        RECT 799.950 721.800 802.050 723.900 ;
        RECT 805.950 723.600 808.050 723.900 ;
        RECT 823.950 723.600 826.050 724.050 ;
        RECT 805.950 722.400 826.050 723.600 ;
        RECT 805.950 721.800 808.050 722.400 ;
        RECT 823.950 721.950 826.050 722.400 ;
        RECT 841.950 723.600 844.050 724.050 ;
        RECT 868.950 723.600 871.050 723.900 ;
        RECT 841.950 722.400 871.050 723.600 ;
        RECT 841.950 721.950 844.050 722.400 ;
        RECT 868.950 721.800 871.050 722.400 ;
        RECT 526.950 720.600 529.050 721.050 ;
        RECT 518.400 719.400 529.050 720.600 ;
        RECT 466.950 718.950 469.050 719.400 ;
        RECT 472.950 718.950 475.050 719.400 ;
        RECT 526.950 718.950 529.050 719.400 ;
        RECT 571.950 720.600 574.050 721.050 ;
        RECT 592.950 720.600 595.050 721.050 ;
        RECT 571.950 719.400 595.050 720.600 ;
        RECT 571.950 718.950 574.050 719.400 ;
        RECT 592.950 718.950 595.050 719.400 ;
        RECT 655.950 720.600 658.050 721.050 ;
        RECT 673.950 720.600 676.050 721.050 ;
        RECT 655.950 719.400 676.050 720.600 ;
        RECT 655.950 718.950 658.050 719.400 ;
        RECT 673.950 718.950 676.050 719.400 ;
        RECT 694.950 720.600 697.050 721.050 ;
        RECT 739.950 720.600 742.050 721.050 ;
        RECT 694.950 719.400 742.050 720.600 ;
        RECT 694.950 718.950 697.050 719.400 ;
        RECT 739.950 718.950 742.050 719.400 ;
        RECT 166.950 717.600 169.050 718.050 ;
        RECT 151.950 717.000 169.050 717.600 ;
        RECT 152.400 716.400 169.050 717.000 ;
        RECT 22.950 715.950 25.050 716.400 ;
        RECT 73.950 715.950 76.050 716.400 ;
        RECT 103.950 715.950 106.050 716.400 ;
        RECT 166.950 715.950 169.050 716.400 ;
        RECT 325.950 717.600 328.050 718.050 ;
        RECT 349.950 717.600 352.050 718.050 ;
        RECT 325.950 716.400 352.050 717.600 ;
        RECT 325.950 715.950 328.050 716.400 ;
        RECT 349.950 715.950 352.050 716.400 ;
        RECT 382.950 717.600 385.050 718.050 ;
        RECT 409.950 717.600 412.050 718.050 ;
        RECT 382.950 716.400 412.050 717.600 ;
        RECT 382.950 715.950 385.050 716.400 ;
        RECT 409.950 715.950 412.050 716.400 ;
        RECT 454.950 717.600 457.050 718.050 ;
        RECT 550.950 717.600 553.050 718.050 ;
        RECT 622.950 717.600 625.050 718.050 ;
        RECT 454.950 716.400 625.050 717.600 ;
        RECT 454.950 715.950 457.050 716.400 ;
        RECT 550.950 715.950 553.050 716.400 ;
        RECT 622.950 715.950 625.050 716.400 ;
        RECT 700.950 717.600 703.050 718.050 ;
        RECT 712.950 717.600 715.050 718.050 ;
        RECT 700.950 716.400 715.050 717.600 ;
        RECT 700.950 715.950 703.050 716.400 ;
        RECT 712.950 715.950 715.050 716.400 ;
        RECT 751.950 717.600 754.050 718.050 ;
        RECT 757.950 717.600 760.050 718.050 ;
        RECT 781.950 717.600 784.050 718.050 ;
        RECT 751.950 716.400 784.050 717.600 ;
        RECT 751.950 715.950 754.050 716.400 ;
        RECT 757.950 715.950 760.050 716.400 ;
        RECT 781.950 715.950 784.050 716.400 ;
        RECT 118.950 714.600 121.050 715.050 ;
        RECT 160.950 714.600 163.050 715.050 ;
        RECT 118.950 713.400 163.050 714.600 ;
        RECT 118.950 712.950 121.050 713.400 ;
        RECT 160.950 712.950 163.050 713.400 ;
        RECT 208.950 714.600 211.050 715.050 ;
        RECT 244.950 714.600 247.050 715.050 ;
        RECT 208.950 713.400 247.050 714.600 ;
        RECT 208.950 712.950 211.050 713.400 ;
        RECT 244.950 712.950 247.050 713.400 ;
        RECT 253.950 714.600 256.050 715.050 ;
        RECT 286.950 714.600 289.050 715.050 ;
        RECT 310.950 714.600 313.050 715.050 ;
        RECT 253.950 713.400 313.050 714.600 ;
        RECT 253.950 712.950 256.050 713.400 ;
        RECT 286.950 712.950 289.050 713.400 ;
        RECT 310.950 712.950 313.050 713.400 ;
        RECT 319.950 714.600 322.050 715.050 ;
        RECT 337.950 714.600 340.050 715.050 ;
        RECT 319.950 713.400 340.050 714.600 ;
        RECT 319.950 712.950 322.050 713.400 ;
        RECT 337.950 712.950 340.050 713.400 ;
        RECT 397.950 714.600 400.050 715.050 ;
        RECT 418.950 714.600 421.050 715.050 ;
        RECT 397.950 713.400 421.050 714.600 ;
        RECT 397.950 712.950 400.050 713.400 ;
        RECT 418.950 712.950 421.050 713.400 ;
        RECT 661.950 714.600 664.050 715.050 ;
        RECT 682.950 714.600 685.050 715.050 ;
        RECT 661.950 713.400 685.050 714.600 ;
        RECT 661.950 712.950 664.050 713.400 ;
        RECT 682.950 712.950 685.050 713.400 ;
        RECT 367.950 711.600 370.050 712.050 ;
        RECT 445.950 711.600 448.050 712.050 ;
        RECT 475.950 711.600 478.050 712.050 ;
        RECT 508.950 711.600 511.050 712.050 ;
        RECT 586.950 711.600 589.050 712.050 ;
        RECT 367.950 710.400 589.050 711.600 ;
        RECT 367.950 709.950 370.050 710.400 ;
        RECT 445.950 709.950 448.050 710.400 ;
        RECT 475.950 709.950 478.050 710.400 ;
        RECT 508.950 709.950 511.050 710.400 ;
        RECT 586.950 709.950 589.050 710.400 ;
        RECT 643.950 711.600 646.050 712.050 ;
        RECT 694.950 711.600 697.050 712.050 ;
        RECT 721.950 711.600 724.050 712.050 ;
        RECT 772.950 711.600 775.050 712.050 ;
        RECT 805.950 711.600 808.050 712.050 ;
        RECT 643.950 710.400 808.050 711.600 ;
        RECT 643.950 709.950 646.050 710.400 ;
        RECT 694.950 709.950 697.050 710.400 ;
        RECT 721.950 709.950 724.050 710.400 ;
        RECT 772.950 709.950 775.050 710.400 ;
        RECT 805.950 709.950 808.050 710.400 ;
        RECT 97.950 708.600 100.050 709.050 ;
        RECT 133.950 708.600 136.050 709.050 ;
        RECT 97.950 707.400 136.050 708.600 ;
        RECT 97.950 706.950 100.050 707.400 ;
        RECT 133.950 706.950 136.050 707.400 ;
        RECT 187.950 708.600 190.050 709.050 ;
        RECT 202.950 708.600 205.050 709.050 ;
        RECT 208.950 708.600 211.050 709.050 ;
        RECT 187.950 707.400 211.050 708.600 ;
        RECT 187.950 706.950 190.050 707.400 ;
        RECT 202.950 706.950 205.050 707.400 ;
        RECT 208.950 706.950 211.050 707.400 ;
        RECT 226.950 708.600 229.050 709.050 ;
        RECT 268.950 708.600 271.050 709.050 ;
        RECT 226.950 707.400 271.050 708.600 ;
        RECT 226.950 706.950 229.050 707.400 ;
        RECT 268.950 706.950 271.050 707.400 ;
        RECT 370.950 708.600 373.050 709.050 ;
        RECT 376.950 708.600 379.050 709.050 ;
        RECT 415.950 708.600 418.050 709.050 ;
        RECT 370.950 707.400 418.050 708.600 ;
        RECT 370.950 706.950 373.050 707.400 ;
        RECT 376.950 706.950 379.050 707.400 ;
        RECT 415.950 706.950 418.050 707.400 ;
        RECT 667.950 708.600 670.050 709.050 ;
        RECT 673.950 708.600 676.050 709.050 ;
        RECT 667.950 707.400 676.050 708.600 ;
        RECT 667.950 706.950 670.050 707.400 ;
        RECT 673.950 706.950 676.050 707.400 ;
        RECT 808.950 708.600 811.050 709.050 ;
        RECT 817.950 708.600 820.050 709.050 ;
        RECT 808.950 707.400 820.050 708.600 ;
        RECT 808.950 706.950 811.050 707.400 ;
        RECT 817.950 706.950 820.050 707.400 ;
        RECT 307.950 705.600 310.050 706.050 ;
        RECT 424.950 705.600 427.050 706.050 ;
        RECT 307.950 704.400 427.050 705.600 ;
        RECT 307.950 703.950 310.050 704.400 ;
        RECT 424.950 703.950 427.050 704.400 ;
        RECT 463.950 705.600 466.050 706.050 ;
        RECT 520.950 705.600 523.050 706.050 ;
        RECT 463.950 704.400 523.050 705.600 ;
        RECT 463.950 703.950 466.050 704.400 ;
        RECT 520.950 703.950 523.050 704.400 ;
        RECT 565.950 705.600 568.050 706.050 ;
        RECT 574.950 705.600 577.050 706.050 ;
        RECT 565.950 704.400 577.050 705.600 ;
        RECT 565.950 703.950 568.050 704.400 ;
        RECT 574.950 703.950 577.050 704.400 ;
        RECT 730.950 705.600 733.050 706.050 ;
        RECT 736.950 705.600 739.050 706.050 ;
        RECT 730.950 704.400 739.050 705.600 ;
        RECT 730.950 703.950 733.050 704.400 ;
        RECT 736.950 703.950 739.050 704.400 ;
        RECT 820.950 705.600 823.050 706.050 ;
        RECT 826.950 705.600 829.050 706.050 ;
        RECT 820.950 704.400 829.050 705.600 ;
        RECT 820.950 703.950 823.050 704.400 ;
        RECT 826.950 703.950 829.050 704.400 ;
        RECT 220.950 702.600 223.050 703.050 ;
        RECT 256.950 702.600 259.050 703.050 ;
        RECT 220.950 701.400 259.050 702.600 ;
        RECT 220.950 700.950 223.050 701.400 ;
        RECT 256.950 700.950 259.050 701.400 ;
        RECT 397.950 702.600 400.050 703.050 ;
        RECT 433.950 702.600 436.050 703.050 ;
        RECT 397.950 701.400 436.050 702.600 ;
        RECT 397.950 700.950 400.050 701.400 ;
        RECT 433.950 700.950 436.050 701.400 ;
        RECT 496.950 702.600 499.050 703.050 ;
        RECT 553.950 702.600 556.050 703.050 ;
        RECT 496.950 701.400 556.050 702.600 ;
        RECT 496.950 700.950 499.050 701.400 ;
        RECT 553.950 700.950 556.050 701.400 ;
        RECT 769.950 702.600 772.050 703.050 ;
        RECT 853.950 702.600 856.050 703.050 ;
        RECT 769.950 701.400 856.050 702.600 ;
        RECT 769.950 700.950 772.050 701.400 ;
        RECT 853.950 700.950 856.050 701.400 ;
        RECT 103.950 699.600 106.050 700.050 ;
        RECT 151.950 699.600 154.050 700.050 ;
        RECT 103.950 698.400 154.050 699.600 ;
        RECT 103.950 697.950 106.050 698.400 ;
        RECT 151.950 697.950 154.050 698.400 ;
        RECT 373.950 699.600 376.050 700.050 ;
        RECT 388.950 699.600 391.050 700.050 ;
        RECT 442.950 699.600 445.050 700.050 ;
        RECT 373.950 698.400 445.050 699.600 ;
        RECT 373.950 697.950 376.050 698.400 ;
        RECT 388.950 697.950 391.050 698.400 ;
        RECT 442.950 697.950 445.050 698.400 ;
        RECT 538.950 699.600 541.050 700.050 ;
        RECT 550.950 699.600 553.050 700.050 ;
        RECT 538.950 698.400 553.050 699.600 ;
        RECT 538.950 697.950 541.050 698.400 ;
        RECT 550.950 697.950 553.050 698.400 ;
        RECT 568.950 699.600 571.050 700.050 ;
        RECT 670.950 699.600 673.050 700.050 ;
        RECT 568.950 698.400 673.050 699.600 ;
        RECT 568.950 697.950 571.050 698.400 ;
        RECT 670.950 697.950 673.050 698.400 ;
        RECT 109.950 696.600 112.050 697.050 ;
        RECT 142.950 696.600 145.050 697.050 ;
        RECT 109.950 695.400 145.050 696.600 ;
        RECT 109.950 694.950 112.050 695.400 ;
        RECT 142.950 694.950 145.050 695.400 ;
        RECT 313.950 696.600 316.050 697.050 ;
        RECT 319.950 696.600 322.050 697.050 ;
        RECT 313.950 695.400 322.050 696.600 ;
        RECT 313.950 694.950 316.050 695.400 ;
        RECT 319.950 694.950 322.050 695.400 ;
        RECT 403.950 696.600 406.050 697.050 ;
        RECT 421.950 696.600 424.050 697.050 ;
        RECT 403.950 695.400 424.050 696.600 ;
        RECT 403.950 694.950 406.050 695.400 ;
        RECT 421.950 694.950 424.050 695.400 ;
        RECT 490.950 696.600 493.050 697.050 ;
        RECT 517.950 696.600 520.050 697.050 ;
        RECT 490.950 695.400 520.050 696.600 ;
        RECT 490.950 694.950 493.050 695.400 ;
        RECT 517.950 694.950 520.050 695.400 ;
        RECT 529.950 696.600 532.050 697.050 ;
        RECT 559.950 696.600 562.050 697.050 ;
        RECT 529.950 695.400 562.050 696.600 ;
        RECT 529.950 694.950 532.050 695.400 ;
        RECT 559.950 694.950 562.050 695.400 ;
        RECT 676.950 696.600 679.050 697.050 ;
        RECT 727.950 696.600 730.050 697.050 ;
        RECT 676.950 695.400 730.050 696.600 ;
        RECT 676.950 694.950 679.050 695.400 ;
        RECT 727.950 694.950 730.050 695.400 ;
        RECT 424.950 693.600 427.050 694.050 ;
        RECT 538.950 693.600 541.050 694.050 ;
        RECT 424.950 692.400 541.050 693.600 ;
        RECT 424.950 691.950 427.050 692.400 ;
        RECT 538.950 691.950 541.050 692.400 ;
        RECT 592.950 693.600 595.050 694.050 ;
        RECT 643.950 693.600 646.050 694.050 ;
        RECT 592.950 692.400 646.050 693.600 ;
        RECT 592.950 691.950 595.050 692.400 ;
        RECT 643.950 691.950 646.050 692.400 ;
        RECT 667.950 693.600 670.050 694.050 ;
        RECT 685.950 693.600 688.050 694.050 ;
        RECT 667.950 692.400 688.050 693.600 ;
        RECT 667.950 691.950 670.050 692.400 ;
        RECT 685.950 691.950 688.050 692.400 ;
        RECT 16.950 690.600 19.050 691.050 ;
        RECT 55.950 690.600 58.050 691.050 ;
        RECT 64.950 690.600 67.050 691.050 ;
        RECT 16.950 689.400 67.050 690.600 ;
        RECT 16.950 688.950 19.050 689.400 ;
        RECT 55.950 688.950 58.050 689.400 ;
        RECT 64.950 688.950 67.050 689.400 ;
        RECT 148.950 690.600 151.050 691.050 ;
        RECT 163.950 690.600 166.050 691.050 ;
        RECT 148.950 689.400 166.050 690.600 ;
        RECT 148.950 688.950 151.050 689.400 ;
        RECT 163.950 688.950 166.050 689.400 ;
        RECT 301.950 690.600 304.050 691.050 ;
        RECT 313.950 690.600 316.050 691.050 ;
        RECT 301.950 689.400 316.050 690.600 ;
        RECT 301.950 688.950 304.050 689.400 ;
        RECT 313.950 688.950 316.050 689.400 ;
        RECT 355.950 690.600 358.050 691.050 ;
        RECT 397.950 690.600 400.050 691.050 ;
        RECT 406.950 690.600 409.050 691.050 ;
        RECT 355.950 689.400 409.050 690.600 ;
        RECT 355.950 688.950 358.050 689.400 ;
        RECT 397.950 688.950 400.050 689.400 ;
        RECT 406.950 688.950 409.050 689.400 ;
        RECT 433.950 690.600 436.050 691.050 ;
        RECT 514.950 690.600 517.050 691.050 ;
        RECT 547.950 690.600 550.050 691.050 ;
        RECT 433.950 689.400 513.600 690.600 ;
        RECT 433.950 688.950 436.050 689.400 ;
        RECT 184.950 687.600 187.050 688.050 ;
        RECT 190.950 687.600 193.050 688.050 ;
        RECT 184.950 686.400 193.050 687.600 ;
        RECT 184.950 685.950 187.050 686.400 ;
        RECT 190.950 685.950 193.050 686.400 ;
        RECT 211.950 687.600 214.050 688.050 ;
        RECT 274.950 687.600 277.050 688.050 ;
        RECT 298.950 687.600 301.050 688.050 ;
        RECT 211.950 686.400 301.050 687.600 ;
        RECT 211.950 685.950 214.050 686.400 ;
        RECT 274.950 685.950 277.050 686.400 ;
        RECT 298.950 685.950 301.050 686.400 ;
        RECT 409.950 687.600 412.050 688.050 ;
        RECT 424.950 687.600 427.050 688.050 ;
        RECT 409.950 686.400 427.050 687.600 ;
        RECT 409.950 685.950 412.050 686.400 ;
        RECT 424.950 685.950 427.050 686.400 ;
        RECT 448.950 687.600 451.050 688.050 ;
        RECT 454.950 687.600 457.050 688.050 ;
        RECT 478.950 687.600 481.050 688.050 ;
        RECT 448.950 686.400 457.050 687.600 ;
        RECT 448.950 685.950 451.050 686.400 ;
        RECT 454.950 685.950 457.050 686.400 ;
        RECT 473.400 686.400 481.050 687.600 ;
        RECT 512.400 687.600 513.600 689.400 ;
        RECT 514.950 689.400 550.050 690.600 ;
        RECT 514.950 688.950 517.050 689.400 ;
        RECT 547.950 688.950 550.050 689.400 ;
        RECT 565.950 690.600 568.050 691.050 ;
        RECT 661.950 690.600 664.050 691.050 ;
        RECT 688.950 690.600 691.050 691.050 ;
        RECT 733.950 690.600 736.050 691.050 ;
        RECT 565.950 689.400 573.600 690.600 ;
        RECT 565.950 688.950 568.050 689.400 ;
        RECT 538.950 687.600 543.000 688.050 ;
        RECT 572.400 687.600 573.600 689.400 ;
        RECT 661.950 689.400 669.600 690.600 ;
        RECT 661.950 688.950 664.050 689.400 ;
        RECT 580.950 687.600 583.050 688.050 ;
        RECT 512.400 686.400 537.600 687.600 ;
        RECT 10.950 684.600 13.050 685.050 ;
        RECT 22.950 684.600 25.050 685.050 ;
        RECT 31.950 684.600 34.050 685.200 ;
        RECT 10.950 683.400 34.050 684.600 ;
        RECT 10.950 682.950 13.050 683.400 ;
        RECT 22.950 682.950 25.050 683.400 ;
        RECT 31.950 683.100 34.050 683.400 ;
        RECT 40.950 684.750 43.050 685.200 ;
        RECT 46.950 684.750 49.050 685.200 ;
        RECT 40.950 683.550 49.050 684.750 ;
        RECT 40.950 683.100 43.050 683.550 ;
        RECT 46.950 683.100 49.050 683.550 ;
        RECT 52.950 684.750 55.050 685.200 ;
        RECT 58.950 684.750 61.050 685.200 ;
        RECT 52.950 683.550 61.050 684.750 ;
        RECT 52.950 683.100 55.050 683.550 ;
        RECT 58.950 683.100 61.050 683.550 ;
        RECT 70.950 683.100 73.050 685.200 ;
        RECT 76.950 684.750 79.050 685.200 ;
        RECT 85.950 684.750 88.050 685.200 ;
        RECT 76.950 683.550 88.050 684.750 ;
        RECT 76.950 683.100 79.050 683.550 ;
        RECT 85.950 683.100 88.050 683.550 ;
        RECT 91.950 684.750 94.050 685.200 ;
        RECT 97.950 684.750 100.050 685.200 ;
        RECT 91.950 683.550 100.050 684.750 ;
        RECT 91.950 683.100 94.050 683.550 ;
        RECT 97.950 683.100 100.050 683.550 ;
        RECT 109.950 684.600 112.050 685.200 ;
        RECT 109.950 683.400 114.600 684.600 ;
        RECT 109.950 683.100 112.050 683.400 ;
        RECT 71.400 681.600 72.600 683.100 ;
        RECT 65.400 680.400 72.600 681.600 ;
        RECT 13.950 678.450 16.050 678.900 ;
        RECT 22.950 678.450 25.050 678.900 ;
        RECT 13.950 677.250 25.050 678.450 ;
        RECT 13.950 676.800 16.050 677.250 ;
        RECT 22.950 676.800 25.050 677.250 ;
        RECT 34.950 678.600 37.050 678.900 ;
        RECT 40.950 678.600 43.050 679.050 ;
        RECT 34.950 677.400 43.050 678.600 ;
        RECT 34.950 676.800 37.050 677.400 ;
        RECT 40.950 676.950 43.050 677.400 ;
        RECT 49.950 678.600 52.050 678.900 ;
        RECT 65.400 678.600 66.600 680.400 ;
        RECT 113.400 679.050 114.600 683.400 ;
        RECT 124.950 683.100 127.050 685.200 ;
        RECT 151.950 684.750 154.050 685.200 ;
        RECT 157.950 684.750 160.050 685.200 ;
        RECT 151.950 683.550 160.050 684.750 ;
        RECT 151.950 683.100 154.050 683.550 ;
        RECT 157.950 683.100 160.050 683.550 ;
        RECT 217.950 684.600 220.050 685.200 ;
        RECT 235.950 684.600 238.050 685.200 ;
        RECT 241.950 684.600 244.050 685.050 ;
        RECT 217.950 683.400 234.600 684.600 ;
        RECT 217.950 683.100 220.050 683.400 ;
        RECT 49.950 677.400 66.600 678.600 ;
        RECT 67.950 678.600 70.050 678.900 ;
        RECT 76.950 678.600 79.050 679.050 ;
        RECT 67.950 677.400 79.050 678.600 ;
        RECT 49.950 676.800 52.050 677.400 ;
        RECT 67.950 676.800 70.050 677.400 ;
        RECT 76.950 676.950 79.050 677.400 ;
        RECT 112.950 676.950 115.050 679.050 ;
        RECT 125.400 678.600 126.600 683.100 ;
        RECT 233.400 678.900 234.600 683.400 ;
        RECT 235.950 683.400 244.050 684.600 ;
        RECT 235.950 683.100 238.050 683.400 ;
        RECT 241.950 682.950 244.050 683.400 ;
        RECT 262.950 684.600 267.000 685.050 ;
        RECT 268.950 684.600 271.050 685.200 ;
        RECT 289.950 684.600 292.050 685.200 ;
        RECT 307.950 684.600 310.050 685.200 ;
        RECT 262.950 682.950 267.600 684.600 ;
        RECT 268.950 683.400 292.050 684.600 ;
        RECT 268.950 683.100 271.050 683.400 ;
        RECT 289.950 683.100 292.050 683.400 ;
        RECT 293.400 683.400 310.050 684.600 ;
        RECT 259.950 681.600 262.050 682.050 ;
        RECT 242.400 681.000 262.050 681.600 ;
        RECT 241.950 680.400 262.050 681.000 ;
        RECT 122.400 677.400 126.600 678.600 ;
        RECT 142.950 678.450 145.050 678.900 ;
        RECT 148.950 678.450 151.050 678.900 ;
        RECT 88.950 675.600 91.050 676.050 ;
        RECT 122.400 675.600 123.600 677.400 ;
        RECT 142.950 677.250 151.050 678.450 ;
        RECT 142.950 676.800 145.050 677.250 ;
        RECT 148.950 676.800 151.050 677.250 ;
        RECT 211.950 678.450 214.050 678.900 ;
        RECT 220.950 678.450 223.050 678.900 ;
        RECT 211.950 677.250 223.050 678.450 ;
        RECT 211.950 676.800 214.050 677.250 ;
        RECT 220.950 676.800 223.050 677.250 ;
        RECT 232.950 676.800 235.050 678.900 ;
        RECT 241.950 676.950 244.050 680.400 ;
        RECT 259.950 679.950 262.050 680.400 ;
        RECT 266.400 678.900 267.600 682.950 ;
        RECT 293.400 678.900 294.600 683.400 ;
        RECT 307.950 683.100 310.050 683.400 ;
        RECT 328.950 684.750 331.050 685.200 ;
        RECT 334.950 684.750 337.050 685.200 ;
        RECT 328.950 683.550 337.050 684.750 ;
        RECT 328.950 683.100 331.050 683.550 ;
        RECT 334.950 683.100 337.050 683.550 ;
        RECT 379.950 683.100 382.050 685.200 ;
        RECT 265.950 676.800 268.050 678.900 ;
        RECT 292.950 676.800 295.050 678.900 ;
        RECT 298.950 678.600 301.050 679.050 ;
        RECT 310.950 678.600 313.050 678.900 ;
        RECT 298.950 677.400 313.050 678.600 ;
        RECT 298.950 676.950 301.050 677.400 ;
        RECT 310.950 676.800 313.050 677.400 ;
        RECT 346.950 678.450 349.050 678.900 ;
        RECT 352.950 678.450 355.050 678.900 ;
        RECT 346.950 677.250 355.050 678.450 ;
        RECT 346.950 676.800 349.050 677.250 ;
        RECT 352.950 676.800 355.050 677.250 ;
        RECT 364.950 678.600 367.050 678.900 ;
        RECT 380.400 678.600 381.600 683.100 ;
        RECT 400.950 682.950 403.050 685.050 ;
        RECT 463.950 684.750 466.050 685.200 ;
        RECT 469.950 684.750 472.050 685.200 ;
        RECT 463.950 683.550 472.050 684.750 ;
        RECT 463.950 683.100 466.050 683.550 ;
        RECT 469.950 683.100 472.050 683.550 ;
        RECT 401.400 679.050 402.600 682.950 ;
        RECT 364.950 677.400 381.600 678.600 ;
        RECT 397.950 677.400 402.600 679.050 ;
        RECT 473.400 678.900 474.600 686.400 ;
        RECT 478.950 685.950 481.050 686.400 ;
        RECT 502.950 684.600 505.050 685.200 ;
        RECT 500.400 683.400 505.050 684.600 ;
        RECT 500.400 679.050 501.600 683.400 ;
        RECT 502.950 683.100 505.050 683.400 ;
        RECT 508.950 684.600 511.050 685.200 ;
        RECT 536.400 684.600 537.600 686.400 ;
        RECT 538.950 685.950 543.600 687.600 ;
        RECT 572.400 686.400 583.050 687.600 ;
        RECT 580.950 685.950 583.050 686.400 ;
        RECT 542.400 684.600 543.600 685.950 ;
        RECT 568.950 684.600 571.050 685.050 ;
        RECT 508.950 683.400 534.600 684.600 ;
        RECT 536.400 683.400 540.600 684.600 ;
        RECT 542.400 683.400 571.050 684.600 ;
        RECT 508.950 683.100 511.050 683.400 ;
        RECT 409.950 678.600 412.050 678.900 ;
        RECT 427.950 678.600 430.050 678.900 ;
        RECT 409.950 678.450 430.050 678.600 ;
        RECT 457.950 678.450 460.050 678.900 ;
        RECT 409.950 677.400 460.050 678.450 ;
        RECT 364.950 676.800 367.050 677.400 ;
        RECT 397.950 676.950 402.000 677.400 ;
        RECT 409.950 676.800 412.050 677.400 ;
        RECT 427.950 677.250 460.050 677.400 ;
        RECT 427.950 676.800 430.050 677.250 ;
        RECT 457.950 676.800 460.050 677.250 ;
        RECT 472.950 676.800 475.050 678.900 ;
        RECT 499.950 676.950 502.050 679.050 ;
        RECT 533.400 678.900 534.600 683.400 ;
        RECT 539.400 681.600 540.600 683.400 ;
        RECT 568.950 682.950 571.050 683.400 ;
        RECT 583.950 684.600 586.050 685.200 ;
        RECT 589.950 684.600 592.050 688.050 ;
        RECT 601.950 687.600 604.050 688.050 ;
        RECT 601.950 686.400 615.600 687.600 ;
        RECT 601.950 685.950 604.050 686.400 ;
        RECT 583.950 684.000 592.050 684.600 ;
        RECT 583.950 683.400 591.600 684.000 ;
        RECT 583.950 683.100 586.050 683.400 ;
        RECT 607.950 682.950 610.050 685.050 ;
        RECT 614.400 684.600 615.600 686.400 ;
        RECT 616.950 684.600 619.050 685.200 ;
        RECT 614.400 683.400 619.050 684.600 ;
        RECT 616.950 683.100 619.050 683.400 ;
        RECT 652.950 684.750 655.050 685.200 ;
        RECT 658.950 684.750 661.050 685.200 ;
        RECT 652.950 683.550 661.050 684.750 ;
        RECT 664.950 684.600 667.050 685.200 ;
        RECT 652.950 683.100 655.050 683.550 ;
        RECT 658.950 683.100 661.050 683.550 ;
        RECT 662.400 683.400 667.050 684.600 ;
        RECT 539.400 680.400 546.600 681.600 ;
        RECT 505.950 678.600 508.050 678.900 ;
        RECT 505.950 678.000 513.600 678.600 ;
        RECT 505.950 677.400 514.050 678.000 ;
        RECT 505.950 676.800 508.050 677.400 ;
        RECT 88.950 674.400 123.600 675.600 ;
        RECT 169.950 675.600 172.050 676.050 ;
        RECT 199.950 675.600 202.050 676.050 ;
        RECT 355.950 675.600 358.050 676.050 ;
        RECT 169.950 674.400 202.050 675.600 ;
        RECT 88.950 673.950 91.050 674.400 ;
        RECT 169.950 673.950 172.050 674.400 ;
        RECT 199.950 673.950 202.050 674.400 ;
        RECT 332.400 674.400 358.050 675.600 ;
        RECT 28.950 672.600 31.050 673.050 ;
        RECT 58.950 672.600 61.050 673.050 ;
        RECT 28.950 671.400 61.050 672.600 ;
        RECT 28.950 670.950 31.050 671.400 ;
        RECT 58.950 670.950 61.050 671.400 ;
        RECT 229.950 672.600 232.050 673.050 ;
        RECT 253.950 672.600 256.050 673.050 ;
        RECT 229.950 671.400 256.050 672.600 ;
        RECT 229.950 670.950 232.050 671.400 ;
        RECT 253.950 670.950 256.050 671.400 ;
        RECT 289.950 672.600 292.050 673.050 ;
        RECT 332.400 672.600 333.600 674.400 ;
        RECT 355.950 673.950 358.050 674.400 ;
        RECT 511.950 673.950 514.050 677.400 ;
        RECT 532.950 676.800 535.050 678.900 ;
        RECT 545.400 675.600 546.600 680.400 ;
        RECT 608.400 679.050 609.600 682.950 ;
        RECT 662.400 681.600 663.600 683.400 ;
        RECT 664.950 683.100 667.050 683.400 ;
        RECT 632.400 680.400 663.600 681.600 ;
        RECT 668.400 681.600 669.600 689.400 ;
        RECT 688.950 689.400 736.050 690.600 ;
        RECT 688.950 688.950 691.050 689.400 ;
        RECT 733.950 688.950 736.050 689.400 ;
        RECT 739.950 690.600 742.050 691.050 ;
        RECT 754.950 690.600 757.050 691.050 ;
        RECT 835.950 690.600 838.050 691.050 ;
        RECT 739.950 689.400 838.050 690.600 ;
        RECT 739.950 688.950 742.050 689.400 ;
        RECT 754.950 688.950 757.050 689.400 ;
        RECT 835.950 688.950 838.050 689.400 ;
        RECT 841.950 690.600 844.050 691.050 ;
        RECT 853.950 690.600 856.050 691.050 ;
        RECT 841.950 689.400 856.050 690.600 ;
        RECT 841.950 688.950 844.050 689.400 ;
        RECT 853.950 688.950 856.050 689.400 ;
        RECT 703.950 684.600 706.050 685.200 ;
        RECT 692.400 683.400 706.050 684.600 ;
        RECT 668.400 680.400 684.600 681.600 ;
        RECT 547.950 678.600 550.050 679.050 ;
        RECT 586.950 678.600 589.050 678.900 ;
        RECT 547.950 678.450 589.050 678.600 ;
        RECT 592.950 678.450 595.050 678.900 ;
        RECT 547.950 677.400 595.050 678.450 ;
        RECT 547.950 676.950 550.050 677.400 ;
        RECT 586.950 677.250 595.050 677.400 ;
        RECT 586.950 676.800 589.050 677.250 ;
        RECT 592.950 676.800 595.050 677.250 ;
        RECT 607.950 676.950 610.050 679.050 ;
        RECT 632.400 678.900 633.600 680.400 ;
        RECT 631.950 676.800 634.050 678.900 ;
        RECT 661.950 678.600 664.050 678.900 ;
        RECT 679.950 678.600 682.050 678.900 ;
        RECT 661.950 677.400 682.050 678.600 ;
        RECT 683.400 678.600 684.600 680.400 ;
        RECT 692.400 679.050 693.600 683.400 ;
        RECT 703.950 683.100 706.050 683.400 ;
        RECT 712.950 684.600 715.050 685.050 ;
        RECT 721.950 684.600 724.050 685.200 ;
        RECT 712.950 683.400 724.050 684.600 ;
        RECT 712.950 682.950 715.050 683.400 ;
        RECT 721.950 683.100 724.050 683.400 ;
        RECT 727.950 684.600 730.050 685.050 ;
        RECT 745.950 684.600 748.050 685.200 ;
        RECT 763.950 684.600 766.050 685.200 ;
        RECT 727.950 683.400 766.050 684.600 ;
        RECT 727.950 682.950 730.050 683.400 ;
        RECT 745.950 683.100 748.050 683.400 ;
        RECT 763.950 683.100 766.050 683.400 ;
        RECT 769.950 681.600 772.050 685.050 ;
        RECT 781.950 684.750 784.050 685.200 ;
        RECT 787.950 684.750 790.050 685.200 ;
        RECT 781.950 683.550 790.050 684.750 ;
        RECT 817.950 684.600 820.050 685.200 ;
        RECT 781.950 683.100 784.050 683.550 ;
        RECT 787.950 683.100 790.050 683.550 ;
        RECT 809.400 683.400 820.050 684.600 ;
        RECT 809.400 682.050 810.600 683.400 ;
        RECT 817.950 683.100 820.050 683.400 ;
        RECT 847.950 683.100 850.050 685.200 ;
        RECT 749.400 681.000 772.050 681.600 ;
        RECT 748.950 680.400 771.600 681.000 ;
        RECT 805.950 680.400 810.600 682.050 ;
        RECT 848.400 681.600 849.600 683.100 ;
        RECT 856.950 682.950 859.050 685.050 ;
        RECT 833.400 680.400 849.600 681.600 ;
        RECT 685.950 678.600 688.050 678.900 ;
        RECT 683.400 677.400 688.050 678.600 ;
        RECT 661.950 676.800 664.050 677.400 ;
        RECT 679.950 676.800 682.050 677.400 ;
        RECT 685.950 676.800 688.050 677.400 ;
        RECT 691.950 676.950 694.050 679.050 ;
        RECT 706.950 678.450 709.050 678.900 ;
        RECT 712.950 678.450 715.050 678.900 ;
        RECT 706.950 677.250 715.050 678.450 ;
        RECT 706.950 676.800 709.050 677.250 ;
        RECT 712.950 676.800 715.050 677.250 ;
        RECT 748.950 676.950 751.050 680.400 ;
        RECT 805.950 679.950 810.000 680.400 ;
        RECT 754.950 678.450 757.050 678.900 ;
        RECT 766.950 678.450 769.050 678.900 ;
        RECT 754.950 677.250 769.050 678.450 ;
        RECT 754.950 676.800 757.050 677.250 ;
        RECT 766.950 676.800 769.050 677.250 ;
        RECT 790.950 678.450 793.050 678.900 ;
        RECT 799.950 678.450 802.050 678.900 ;
        RECT 790.950 677.250 802.050 678.450 ;
        RECT 790.950 676.800 793.050 677.250 ;
        RECT 799.950 676.800 802.050 677.250 ;
        RECT 814.950 678.600 817.050 678.900 ;
        RECT 833.400 678.600 834.600 680.400 ;
        RECT 857.400 679.050 858.600 682.950 ;
        RECT 814.950 677.400 834.600 678.600 ;
        RECT 814.950 676.800 817.050 677.400 ;
        RECT 856.950 676.950 859.050 679.050 ;
        RECT 700.950 675.600 703.050 676.050 ;
        RECT 742.950 675.600 745.050 676.050 ;
        RECT 545.400 674.400 579.600 675.600 ;
        RECT 578.400 673.050 579.600 674.400 ;
        RECT 700.950 674.400 745.050 675.600 ;
        RECT 700.950 673.950 703.050 674.400 ;
        RECT 742.950 673.950 745.050 674.400 ;
        RECT 289.950 671.400 333.600 672.600 ;
        RECT 334.950 672.600 337.050 673.050 ;
        RECT 352.950 672.600 355.050 673.050 ;
        RECT 334.950 671.400 355.050 672.600 ;
        RECT 289.950 670.950 292.050 671.400 ;
        RECT 334.950 670.950 337.050 671.400 ;
        RECT 352.950 670.950 355.050 671.400 ;
        RECT 361.950 672.600 364.050 673.050 ;
        RECT 382.950 672.600 385.050 673.050 ;
        RECT 361.950 671.400 385.050 672.600 ;
        RECT 361.950 670.950 364.050 671.400 ;
        RECT 382.950 670.950 385.050 671.400 ;
        RECT 388.950 672.600 391.050 673.050 ;
        RECT 403.950 672.600 406.050 673.050 ;
        RECT 388.950 671.400 406.050 672.600 ;
        RECT 388.950 670.950 391.050 671.400 ;
        RECT 403.950 670.950 406.050 671.400 ;
        RECT 496.950 672.600 499.050 673.050 ;
        RECT 526.950 672.600 529.050 673.050 ;
        RECT 496.950 671.400 529.050 672.600 ;
        RECT 578.400 671.400 583.050 673.050 ;
        RECT 496.950 670.950 499.050 671.400 ;
        RECT 526.950 670.950 529.050 671.400 ;
        RECT 579.000 670.950 583.050 671.400 ;
        RECT 601.950 672.600 604.050 673.050 ;
        RECT 610.950 672.600 613.050 673.050 ;
        RECT 601.950 671.400 613.050 672.600 ;
        RECT 601.950 670.950 604.050 671.400 ;
        RECT 610.950 670.950 613.050 671.400 ;
        RECT 646.950 672.600 649.050 673.050 ;
        RECT 652.950 672.600 655.050 673.050 ;
        RECT 685.950 672.600 688.050 673.050 ;
        RECT 646.950 671.400 688.050 672.600 ;
        RECT 646.950 670.950 649.050 671.400 ;
        RECT 652.950 670.950 655.050 671.400 ;
        RECT 685.950 670.950 688.050 671.400 ;
        RECT 781.950 672.600 784.050 673.050 ;
        RECT 814.950 672.600 817.050 673.050 ;
        RECT 781.950 671.400 817.050 672.600 ;
        RECT 781.950 670.950 784.050 671.400 ;
        RECT 814.950 670.950 817.050 671.400 ;
        RECT 832.950 672.600 835.050 673.050 ;
        RECT 850.950 672.600 853.050 673.050 ;
        RECT 832.950 671.400 853.050 672.600 ;
        RECT 832.950 670.950 835.050 671.400 ;
        RECT 850.950 670.950 853.050 671.400 ;
        RECT 97.950 669.600 100.050 670.050 ;
        RECT 160.950 669.600 163.050 670.050 ;
        RECT 97.950 668.400 163.050 669.600 ;
        RECT 97.950 667.950 100.050 668.400 ;
        RECT 160.950 667.950 163.050 668.400 ;
        RECT 172.950 669.600 175.050 670.050 ;
        RECT 178.950 669.600 181.050 670.050 ;
        RECT 220.950 669.600 223.050 670.050 ;
        RECT 226.950 669.600 229.050 670.050 ;
        RECT 172.950 668.400 229.050 669.600 ;
        RECT 172.950 667.950 175.050 668.400 ;
        RECT 178.950 667.950 181.050 668.400 ;
        RECT 220.950 667.950 223.050 668.400 ;
        RECT 226.950 667.950 229.050 668.400 ;
        RECT 388.950 669.600 391.050 669.900 ;
        RECT 394.950 669.600 397.050 670.050 ;
        RECT 388.950 668.400 397.050 669.600 ;
        RECT 388.950 667.800 391.050 668.400 ;
        RECT 394.950 667.950 397.050 668.400 ;
        RECT 424.950 669.600 427.050 670.050 ;
        RECT 499.950 669.600 502.050 670.050 ;
        RECT 538.950 669.600 541.050 670.050 ;
        RECT 424.950 668.400 541.050 669.600 ;
        RECT 424.950 667.950 427.050 668.400 ;
        RECT 499.950 667.950 502.050 668.400 ;
        RECT 538.950 667.950 541.050 668.400 ;
        RECT 655.950 669.600 658.050 670.050 ;
        RECT 670.800 669.600 672.900 670.050 ;
        RECT 655.950 668.400 672.900 669.600 ;
        RECT 655.950 667.950 658.050 668.400 ;
        RECT 670.800 667.950 672.900 668.400 ;
        RECT 673.950 669.600 676.050 670.050 ;
        RECT 688.950 669.600 691.050 670.050 ;
        RECT 673.950 668.400 691.050 669.600 ;
        RECT 673.950 667.950 676.050 668.400 ;
        RECT 688.950 667.950 691.050 668.400 ;
        RECT 730.950 669.600 733.050 670.050 ;
        RECT 745.950 669.600 748.050 670.050 ;
        RECT 730.950 668.400 748.050 669.600 ;
        RECT 730.950 667.950 733.050 668.400 ;
        RECT 745.950 667.950 748.050 668.400 ;
        RECT 820.950 669.600 823.050 670.050 ;
        RECT 835.950 669.600 838.050 670.050 ;
        RECT 841.950 669.600 844.050 670.050 ;
        RECT 820.950 668.400 844.050 669.600 ;
        RECT 820.950 667.950 823.050 668.400 ;
        RECT 835.950 667.950 838.050 668.400 ;
        RECT 841.950 667.950 844.050 668.400 ;
        RECT 40.950 666.600 43.050 667.050 ;
        RECT 55.950 666.600 58.050 667.050 ;
        RECT 40.950 665.400 58.050 666.600 ;
        RECT 40.950 664.950 43.050 665.400 ;
        RECT 55.950 664.950 58.050 665.400 ;
        RECT 190.950 666.600 193.050 667.050 ;
        RECT 205.950 666.600 208.050 667.050 ;
        RECT 232.950 666.600 235.050 667.050 ;
        RECT 190.950 665.400 235.050 666.600 ;
        RECT 190.950 664.950 193.050 665.400 ;
        RECT 205.950 664.950 208.050 665.400 ;
        RECT 232.950 664.950 235.050 665.400 ;
        RECT 364.950 666.600 367.050 667.050 ;
        RECT 397.950 666.600 400.050 667.050 ;
        RECT 454.950 666.600 457.050 667.050 ;
        RECT 466.950 666.600 469.050 667.050 ;
        RECT 559.950 666.600 562.050 667.050 ;
        RECT 364.950 665.400 562.050 666.600 ;
        RECT 364.950 664.950 367.050 665.400 ;
        RECT 397.950 664.950 400.050 665.400 ;
        RECT 454.950 664.950 457.050 665.400 ;
        RECT 466.950 664.950 469.050 665.400 ;
        RECT 559.950 664.950 562.050 665.400 ;
        RECT 589.950 666.600 592.050 667.050 ;
        RECT 601.950 666.600 604.050 667.050 ;
        RECT 613.950 666.600 616.050 667.050 ;
        RECT 589.950 665.400 616.050 666.600 ;
        RECT 589.950 664.950 592.050 665.400 ;
        RECT 601.950 664.950 604.050 665.400 ;
        RECT 613.950 664.950 616.050 665.400 ;
        RECT 778.950 666.600 781.050 667.050 ;
        RECT 787.950 666.600 790.050 667.050 ;
        RECT 778.950 665.400 790.050 666.600 ;
        RECT 778.950 664.950 781.050 665.400 ;
        RECT 787.950 664.950 790.050 665.400 ;
        RECT 826.950 666.600 829.050 667.050 ;
        RECT 832.950 666.600 835.050 667.050 ;
        RECT 826.950 665.400 835.050 666.600 ;
        RECT 826.950 664.950 829.050 665.400 ;
        RECT 832.950 664.950 835.050 665.400 ;
        RECT 850.950 666.600 853.050 667.050 ;
        RECT 868.950 666.600 871.050 667.050 ;
        RECT 850.950 665.400 871.050 666.600 ;
        RECT 850.950 664.950 853.050 665.400 ;
        RECT 868.950 664.950 871.050 665.400 ;
        RECT 82.950 663.600 85.050 664.050 ;
        RECT 142.950 663.600 145.050 664.050 ;
        RECT 82.950 662.400 145.050 663.600 ;
        RECT 82.950 661.950 85.050 662.400 ;
        RECT 142.950 661.950 145.050 662.400 ;
        RECT 457.950 663.600 460.050 664.050 ;
        RECT 514.950 663.600 517.050 664.050 ;
        RECT 547.950 663.600 550.050 664.050 ;
        RECT 457.950 662.400 517.050 663.600 ;
        RECT 457.950 661.950 460.050 662.400 ;
        RECT 514.950 661.950 517.050 662.400 ;
        RECT 533.400 662.400 550.050 663.600 ;
        RECT 58.950 660.600 61.050 661.050 ;
        RECT 73.950 660.600 76.050 661.050 ;
        RECT 58.950 659.400 76.050 660.600 ;
        RECT 58.950 658.950 61.050 659.400 ;
        RECT 73.950 658.950 76.050 659.400 ;
        RECT 208.950 660.600 211.050 661.050 ;
        RECT 238.950 660.600 241.050 661.050 ;
        RECT 208.950 659.400 241.050 660.600 ;
        RECT 208.950 658.950 211.050 659.400 ;
        RECT 238.950 658.950 241.050 659.400 ;
        RECT 349.950 660.600 352.050 661.050 ;
        RECT 379.950 660.600 382.050 661.050 ;
        RECT 349.950 659.400 382.050 660.600 ;
        RECT 349.950 658.950 352.050 659.400 ;
        RECT 379.950 658.950 382.050 659.400 ;
        RECT 397.950 660.600 400.050 661.050 ;
        RECT 421.950 660.600 424.050 661.050 ;
        RECT 397.950 659.400 424.050 660.600 ;
        RECT 397.950 658.950 400.050 659.400 ;
        RECT 421.950 658.950 424.050 659.400 ;
        RECT 442.950 660.600 445.050 661.050 ;
        RECT 484.950 660.600 487.050 661.050 ;
        RECT 493.950 660.600 496.050 661.050 ;
        RECT 533.400 660.600 534.600 662.400 ;
        RECT 547.950 661.950 550.050 662.400 ;
        RECT 604.950 663.600 607.050 664.050 ;
        RECT 700.950 663.600 703.050 664.050 ;
        RECT 604.950 662.400 703.050 663.600 ;
        RECT 604.950 661.950 607.050 662.400 ;
        RECT 700.950 661.950 703.050 662.400 ;
        RECT 724.950 663.600 727.050 664.050 ;
        RECT 754.950 663.600 757.050 664.050 ;
        RECT 724.950 662.400 757.050 663.600 ;
        RECT 724.950 661.950 727.050 662.400 ;
        RECT 754.950 661.950 757.050 662.400 ;
        RECT 763.950 663.600 766.050 664.050 ;
        RECT 805.950 663.600 808.050 664.050 ;
        RECT 763.950 662.400 808.050 663.600 ;
        RECT 763.950 661.950 766.050 662.400 ;
        RECT 805.950 661.950 808.050 662.400 ;
        RECT 814.950 663.600 817.050 664.050 ;
        RECT 847.950 663.600 850.050 664.050 ;
        RECT 814.950 662.400 850.050 663.600 ;
        RECT 814.950 661.950 817.050 662.400 ;
        RECT 847.950 661.950 850.050 662.400 ;
        RECT 442.950 659.400 534.600 660.600 ;
        RECT 580.950 660.600 583.050 661.050 ;
        RECT 586.950 660.600 589.050 661.050 ;
        RECT 580.950 659.400 589.050 660.600 ;
        RECT 442.950 658.950 445.050 659.400 ;
        RECT 484.950 658.950 487.050 659.400 ;
        RECT 493.950 658.950 496.050 659.400 ;
        RECT 580.950 658.950 583.050 659.400 ;
        RECT 586.950 658.950 589.050 659.400 ;
        RECT 592.950 660.600 595.050 661.050 ;
        RECT 616.950 660.600 619.050 661.050 ;
        RECT 673.950 660.600 676.050 661.050 ;
        RECT 592.950 659.400 615.600 660.600 ;
        RECT 592.950 658.950 595.050 659.400 ;
        RECT 7.950 657.600 10.050 658.050 ;
        RECT 46.950 657.600 49.050 658.050 ;
        RECT 7.950 656.400 49.050 657.600 ;
        RECT 7.950 655.950 10.050 656.400 ;
        RECT 46.950 655.950 49.050 656.400 ;
        RECT 82.950 657.600 85.050 658.050 ;
        RECT 91.950 657.600 94.050 658.050 ;
        RECT 82.950 656.400 94.050 657.600 ;
        RECT 82.950 655.950 85.050 656.400 ;
        RECT 91.950 655.950 94.050 656.400 ;
        RECT 175.950 657.600 178.050 658.050 ;
        RECT 208.950 657.600 211.050 657.900 ;
        RECT 175.950 656.400 211.050 657.600 ;
        RECT 175.950 655.950 178.050 656.400 ;
        RECT 208.950 655.800 211.050 656.400 ;
        RECT 319.950 657.600 322.050 658.050 ;
        RECT 337.950 657.600 340.050 658.050 ;
        RECT 319.950 656.400 340.050 657.600 ;
        RECT 614.400 657.600 615.600 659.400 ;
        RECT 616.950 659.400 676.050 660.600 ;
        RECT 616.950 658.950 619.050 659.400 ;
        RECT 673.950 658.950 676.050 659.400 ;
        RECT 700.950 657.600 703.050 658.050 ;
        RECT 724.950 657.600 727.050 658.050 ;
        RECT 614.400 656.400 630.600 657.600 ;
        RECT 319.950 655.950 322.050 656.400 ;
        RECT 337.950 655.950 340.050 656.400 ;
        RECT 70.950 654.600 73.050 655.050 ;
        RECT 94.950 654.600 97.050 655.050 ;
        RECT 103.950 654.600 106.050 655.050 ;
        RECT 70.950 653.400 106.050 654.600 ;
        RECT 70.950 652.950 73.050 653.400 ;
        RECT 94.950 652.950 97.050 653.400 ;
        RECT 103.950 652.950 106.050 653.400 ;
        RECT 136.950 654.600 139.050 655.050 ;
        RECT 145.950 654.600 148.050 655.050 ;
        RECT 163.950 654.600 166.050 655.050 ;
        RECT 136.950 653.400 166.050 654.600 ;
        RECT 136.950 652.950 139.050 653.400 ;
        RECT 145.950 652.950 148.050 653.400 ;
        RECT 163.950 652.950 166.050 653.400 ;
        RECT 286.950 654.600 289.050 655.050 ;
        RECT 301.950 654.600 304.050 655.050 ;
        RECT 310.950 654.600 313.050 655.050 ;
        RECT 286.950 653.400 313.050 654.600 ;
        RECT 286.950 652.950 289.050 653.400 ;
        RECT 301.950 652.950 304.050 653.400 ;
        RECT 310.950 652.950 313.050 653.400 ;
        RECT 439.950 654.600 442.050 655.050 ;
        RECT 445.950 654.600 448.050 655.050 ;
        RECT 439.950 653.400 448.050 654.600 ;
        RECT 439.950 652.950 442.050 653.400 ;
        RECT 445.950 652.950 448.050 653.400 ;
        RECT 538.950 654.600 541.050 655.050 ;
        RECT 550.950 654.600 553.050 655.050 ;
        RECT 574.950 654.600 577.050 655.050 ;
        RECT 615.000 654.600 619.050 655.050 ;
        RECT 538.950 653.400 553.050 654.600 ;
        RECT 538.950 652.950 541.050 653.400 ;
        RECT 550.950 652.950 553.050 653.400 ;
        RECT 569.400 653.400 577.050 654.600 ;
        RECT 13.950 651.600 16.050 652.200 ;
        RECT 37.950 651.600 40.050 652.050 ;
        RECT 13.950 650.400 40.050 651.600 ;
        RECT 13.950 650.100 16.050 650.400 ;
        RECT 37.950 649.950 40.050 650.400 ;
        RECT 61.950 650.100 64.050 652.200 ;
        RECT 88.950 651.600 91.050 652.200 ;
        RECT 106.950 651.600 109.050 652.050 ;
        RECT 68.400 650.400 91.050 651.600 ;
        RECT 10.950 645.600 13.050 645.900 ;
        RECT 28.950 645.600 31.050 645.900 ;
        RECT 10.950 644.400 31.050 645.600 ;
        RECT 10.950 643.800 13.050 644.400 ;
        RECT 28.950 643.800 31.050 644.400 ;
        RECT 37.950 645.450 40.050 645.900 ;
        RECT 43.950 645.450 46.050 645.900 ;
        RECT 37.950 644.250 46.050 645.450 ;
        RECT 37.950 643.800 40.050 644.250 ;
        RECT 43.950 643.800 46.050 644.250 ;
        RECT 52.950 645.600 55.050 646.050 ;
        RECT 62.400 645.600 63.600 650.100 ;
        RECT 52.950 644.400 63.600 645.600 ;
        RECT 64.950 645.600 67.050 645.900 ;
        RECT 68.400 645.600 69.600 650.400 ;
        RECT 88.950 650.100 91.050 650.400 ;
        RECT 98.400 650.400 109.050 651.600 ;
        RECT 98.400 648.600 99.600 650.400 ;
        RECT 106.950 649.950 109.050 650.400 ;
        RECT 154.950 651.600 157.050 652.200 ;
        RECT 196.950 651.600 199.050 652.050 ;
        RECT 154.950 650.400 199.050 651.600 ;
        RECT 154.950 650.100 157.050 650.400 ;
        RECT 196.950 649.950 199.050 650.400 ;
        RECT 214.950 650.100 217.050 652.200 ;
        RECT 346.950 651.750 349.050 652.200 ;
        RECT 358.950 651.750 361.050 652.200 ;
        RECT 346.950 650.550 361.050 651.750 ;
        RECT 346.950 650.100 349.050 650.550 ;
        RECT 358.950 650.100 361.050 650.550 ;
        RECT 364.950 651.600 367.050 652.200 ;
        RECT 364.950 650.400 378.600 651.600 ;
        RECT 364.950 650.100 367.050 650.400 ;
        RECT 80.400 647.400 99.600 648.600 ;
        RECT 80.400 645.900 81.600 647.400 ;
        RECT 64.950 644.400 69.600 645.600 ;
        RECT 52.950 643.950 55.050 644.400 ;
        RECT 64.950 643.800 67.050 644.400 ;
        RECT 79.950 643.800 82.050 645.900 ;
        RECT 145.950 645.450 148.050 645.900 ;
        RECT 151.950 645.450 154.050 645.900 ;
        RECT 145.950 644.250 154.050 645.450 ;
        RECT 145.950 643.800 148.050 644.250 ;
        RECT 151.950 643.800 154.050 644.250 ;
        RECT 175.950 645.600 178.050 646.050 ;
        RECT 181.950 645.600 184.050 645.900 ;
        RECT 175.950 644.400 184.050 645.600 ;
        RECT 175.950 643.950 178.050 644.400 ;
        RECT 181.950 643.800 184.050 644.400 ;
        RECT 193.950 645.600 196.050 646.050 ;
        RECT 215.400 645.600 216.600 650.100 ;
        RECT 226.950 645.600 229.050 645.900 ;
        RECT 193.950 644.400 229.050 645.600 ;
        RECT 193.950 643.950 196.050 644.400 ;
        RECT 226.950 643.800 229.050 644.400 ;
        RECT 328.950 645.600 331.050 645.900 ;
        RECT 346.800 645.600 348.900 646.050 ;
        RECT 377.400 645.900 378.600 650.400 ;
        RECT 403.950 650.100 406.050 652.200 ;
        RECT 409.950 651.750 412.050 652.200 ;
        RECT 418.950 651.750 421.050 652.200 ;
        RECT 409.950 650.550 421.050 651.750 ;
        RECT 409.950 650.100 412.050 650.550 ;
        RECT 418.950 650.100 421.050 650.550 ;
        RECT 499.950 651.600 502.050 652.200 ;
        RECT 499.950 650.400 513.600 651.600 ;
        RECT 499.950 650.100 502.050 650.400 ;
        RECT 404.400 646.050 405.600 650.100 ;
        RECT 328.950 644.400 348.900 645.600 ;
        RECT 328.950 643.800 331.050 644.400 ;
        RECT 346.800 643.950 348.900 644.400 ;
        RECT 349.950 645.450 352.050 645.900 ;
        RECT 355.950 645.450 358.050 645.900 ;
        RECT 349.950 644.250 358.050 645.450 ;
        RECT 349.950 643.800 352.050 644.250 ;
        RECT 355.950 643.800 358.050 644.250 ;
        RECT 376.950 643.800 379.050 645.900 ;
        RECT 404.400 644.400 409.050 646.050 ;
        RECT 512.400 645.600 513.600 650.400 ;
        RECT 532.950 650.100 535.050 652.200 ;
        RECT 553.950 651.600 556.050 652.200 ;
        RECT 542.400 650.400 556.050 651.600 ;
        RECT 533.400 648.600 534.600 650.100 ;
        RECT 542.400 649.050 543.600 650.400 ;
        RECT 553.950 650.100 556.050 650.400 ;
        RECT 559.950 651.750 562.050 652.200 ;
        RECT 565.950 651.750 568.050 652.200 ;
        RECT 559.950 650.550 568.050 651.750 ;
        RECT 559.950 650.100 562.050 650.550 ;
        RECT 565.950 650.100 568.050 650.550 ;
        RECT 541.950 648.600 544.050 649.050 ;
        RECT 533.400 647.400 544.050 648.600 ;
        RECT 541.950 646.950 544.050 647.400 ;
        RECT 569.400 645.900 570.600 653.400 ;
        RECT 574.950 652.950 577.050 653.400 ;
        RECT 614.400 652.950 619.050 654.600 ;
        RECT 629.400 654.600 630.600 656.400 ;
        RECT 700.950 656.400 727.050 657.600 ;
        RECT 700.950 655.950 703.050 656.400 ;
        RECT 724.950 655.950 727.050 656.400 ;
        RECT 814.950 657.600 817.050 658.050 ;
        RECT 850.800 657.600 852.900 658.050 ;
        RECT 814.950 656.400 852.900 657.600 ;
        RECT 853.950 657.600 856.050 661.050 ;
        RECT 862.950 657.600 865.050 658.050 ;
        RECT 853.950 657.000 865.050 657.600 ;
        RECT 854.400 656.400 865.050 657.000 ;
        RECT 814.950 655.950 817.050 656.400 ;
        RECT 850.800 655.950 852.900 656.400 ;
        RECT 862.950 655.950 865.050 656.400 ;
        RECT 629.400 653.400 633.600 654.600 ;
        RECT 583.950 651.600 586.050 652.050 ;
        RECT 614.400 651.600 615.600 652.950 ;
        RECT 583.950 650.400 615.600 651.600 ;
        RECT 583.950 649.950 586.050 650.400 ;
        RECT 619.950 650.100 622.050 652.200 ;
        RECT 514.950 645.600 517.050 645.900 ;
        RECT 512.400 644.400 517.050 645.600 ;
        RECT 405.000 643.950 409.050 644.400 ;
        RECT 514.950 643.800 517.050 644.400 ;
        RECT 568.950 643.800 571.050 645.900 ;
        RECT 580.950 645.450 583.050 645.900 ;
        RECT 595.950 645.450 598.050 645.900 ;
        RECT 580.950 644.250 598.050 645.450 ;
        RECT 580.950 643.800 583.050 644.250 ;
        RECT 595.950 643.800 598.050 644.250 ;
        RECT 613.950 645.600 616.050 645.900 ;
        RECT 620.400 645.600 621.600 650.100 ;
        RECT 613.950 644.400 621.600 645.600 ;
        RECT 632.400 645.600 633.600 653.400 ;
        RECT 718.950 651.600 721.050 652.200 ;
        RECT 724.950 651.600 727.050 652.050 ;
        RECT 730.950 651.600 733.050 652.200 ;
        RECT 742.950 651.600 745.050 655.050 ;
        RECT 718.950 650.400 727.050 651.600 ;
        RECT 718.950 650.100 721.050 650.400 ;
        RECT 724.950 649.950 727.050 650.400 ;
        RECT 728.400 650.400 733.050 651.600 ;
        RECT 728.400 648.600 729.600 650.400 ;
        RECT 730.950 650.100 733.050 650.400 ;
        RECT 740.400 651.000 745.050 651.600 ;
        RECT 769.950 651.600 772.050 652.200 ;
        RECT 775.950 651.600 778.050 655.050 ;
        RECT 769.950 651.000 778.050 651.600 ;
        RECT 740.400 650.400 744.600 651.000 ;
        RECT 769.950 650.400 777.600 651.000 ;
        RECT 740.400 648.600 741.600 650.400 ;
        RECT 769.950 650.100 772.050 650.400 ;
        RECT 781.950 649.950 784.050 652.050 ;
        RECT 787.950 651.600 790.050 652.200 ;
        RECT 796.950 651.600 799.050 652.050 ;
        RECT 787.950 650.400 799.050 651.600 ;
        RECT 787.950 650.100 790.050 650.400 ;
        RECT 796.950 649.950 799.050 650.400 ;
        RECT 802.950 650.100 805.050 652.200 ;
        RECT 719.400 647.400 729.600 648.600 ;
        RECT 734.400 647.400 741.600 648.600 ;
        RECT 637.950 645.600 640.050 645.900 ;
        RECT 632.400 644.400 640.050 645.600 ;
        RECT 613.950 643.800 616.050 644.400 ;
        RECT 637.950 643.800 640.050 644.400 ;
        RECT 673.950 645.450 676.050 645.900 ;
        RECT 691.950 645.450 694.050 645.900 ;
        RECT 673.950 644.250 694.050 645.450 ;
        RECT 673.950 643.800 676.050 644.250 ;
        RECT 691.950 643.800 694.050 644.250 ;
        RECT 715.950 645.600 718.050 645.900 ;
        RECT 719.400 645.600 720.600 647.400 ;
        RECT 734.400 645.900 735.600 647.400 ;
        RECT 715.950 644.400 720.600 645.600 ;
        RECT 715.950 643.800 718.050 644.400 ;
        RECT 733.950 643.800 736.050 645.900 ;
        RECT 742.950 645.600 745.050 646.050 ;
        RECT 751.950 645.600 754.050 645.900 ;
        RECT 742.950 644.400 754.050 645.600 ;
        RECT 742.950 643.950 745.050 644.400 ;
        RECT 751.950 643.800 754.050 644.400 ;
        RECT 772.950 645.600 775.050 645.900 ;
        RECT 782.400 645.600 783.600 649.950 ;
        RECT 772.950 644.400 783.600 645.600 ;
        RECT 803.400 645.600 804.600 650.100 ;
        RECT 832.950 649.950 835.050 652.050 ;
        RECT 868.950 650.100 871.050 652.200 ;
        RECT 817.950 645.600 820.050 646.050 ;
        RECT 803.400 644.400 820.050 645.600 ;
        RECT 833.400 645.600 834.600 649.950 ;
        RECT 850.950 645.600 853.050 646.050 ;
        RECT 833.400 644.400 853.050 645.600 ;
        RECT 772.950 643.800 775.050 644.400 ;
        RECT 817.950 643.950 820.050 644.400 ;
        RECT 850.950 643.950 853.050 644.400 ;
        RECT 859.950 645.600 862.050 646.050 ;
        RECT 869.400 645.600 870.600 650.100 ;
        RECT 874.950 649.950 877.050 652.050 ;
        RECT 875.400 646.050 876.600 649.950 ;
        RECT 859.950 644.400 870.600 645.600 ;
        RECT 859.950 643.950 862.050 644.400 ;
        RECT 874.950 643.950 877.050 646.050 ;
        RECT 238.950 642.600 241.050 643.050 ;
        RECT 283.950 642.600 286.050 643.050 ;
        RECT 238.950 641.400 286.050 642.600 ;
        RECT 238.950 640.950 241.050 641.400 ;
        RECT 283.950 640.950 286.050 641.400 ;
        RECT 409.950 642.600 412.050 643.050 ;
        RECT 418.950 642.600 421.050 643.050 ;
        RECT 409.950 641.400 421.050 642.600 ;
        RECT 409.950 640.950 412.050 641.400 ;
        RECT 418.950 640.950 421.050 641.400 ;
        RECT 430.950 642.600 433.050 643.050 ;
        RECT 445.950 642.600 448.050 643.050 ;
        RECT 505.950 642.600 508.050 643.050 ;
        RECT 430.950 641.400 508.050 642.600 ;
        RECT 430.950 640.950 433.050 641.400 ;
        RECT 445.950 640.950 448.050 641.400 ;
        RECT 505.950 640.950 508.050 641.400 ;
        RECT 592.950 642.600 595.050 643.050 ;
        RECT 607.950 642.600 610.050 643.050 ;
        RECT 592.950 641.400 610.050 642.600 ;
        RECT 592.950 640.950 595.050 641.400 ;
        RECT 607.950 640.950 610.050 641.400 ;
        RECT 646.950 642.600 649.050 643.050 ;
        RECT 673.950 642.600 676.050 643.050 ;
        RECT 703.950 642.600 706.050 643.050 ;
        RECT 646.950 641.400 706.050 642.600 ;
        RECT 646.950 640.950 649.050 641.400 ;
        RECT 673.950 640.950 676.050 641.400 ;
        RECT 703.950 640.950 706.050 641.400 ;
        RECT 802.950 642.600 805.050 643.050 ;
        RECT 811.950 642.600 814.050 643.050 ;
        RECT 802.950 641.400 814.050 642.600 ;
        RECT 802.950 640.950 805.050 641.400 ;
        RECT 811.950 640.950 814.050 641.400 ;
        RECT 97.950 639.600 100.050 640.050 ;
        RECT 124.950 639.600 127.050 640.050 ;
        RECT 97.950 638.400 127.050 639.600 ;
        RECT 97.950 637.950 100.050 638.400 ;
        RECT 124.950 637.950 127.050 638.400 ;
        RECT 142.950 639.600 145.050 640.050 ;
        RECT 148.950 639.600 151.050 640.050 ;
        RECT 157.950 639.600 160.050 640.050 ;
        RECT 193.950 639.600 196.050 640.050 ;
        RECT 142.950 638.400 196.050 639.600 ;
        RECT 142.950 637.950 145.050 638.400 ;
        RECT 148.950 637.950 151.050 638.400 ;
        RECT 157.950 637.950 160.050 638.400 ;
        RECT 193.950 637.950 196.050 638.400 ;
        RECT 220.950 639.600 223.050 640.050 ;
        RECT 226.950 639.600 229.050 640.050 ;
        RECT 220.950 638.400 229.050 639.600 ;
        RECT 220.950 637.950 223.050 638.400 ;
        RECT 226.950 637.950 229.050 638.400 ;
        RECT 295.950 639.600 298.050 640.050 ;
        RECT 394.950 639.600 397.050 640.050 ;
        RECT 295.950 638.400 397.050 639.600 ;
        RECT 295.950 637.950 298.050 638.400 ;
        RECT 394.950 637.950 397.050 638.400 ;
        RECT 589.950 639.600 592.050 640.050 ;
        RECT 598.950 639.600 601.050 640.050 ;
        RECT 589.950 638.400 601.050 639.600 ;
        RECT 589.950 637.950 592.050 638.400 ;
        RECT 598.950 637.950 601.050 638.400 ;
        RECT 613.950 639.600 616.050 640.050 ;
        RECT 661.950 639.600 664.050 640.050 ;
        RECT 613.950 638.400 664.050 639.600 ;
        RECT 613.950 637.950 616.050 638.400 ;
        RECT 661.950 637.950 664.050 638.400 ;
        RECT 796.950 639.600 799.050 640.050 ;
        RECT 808.950 639.600 811.050 640.050 ;
        RECT 796.950 638.400 811.050 639.600 ;
        RECT 796.950 637.950 799.050 638.400 ;
        RECT 808.950 637.950 811.050 638.400 ;
        RECT 814.950 639.600 817.050 640.050 ;
        RECT 829.950 639.600 832.050 643.050 ;
        RECT 835.950 642.600 838.050 643.050 ;
        RECT 871.950 642.600 874.050 643.050 ;
        RECT 835.950 641.400 874.050 642.600 ;
        RECT 835.950 640.950 838.050 641.400 ;
        RECT 871.950 640.950 874.050 641.400 ;
        RECT 814.950 639.000 832.050 639.600 ;
        RECT 859.950 639.600 862.050 640.050 ;
        RECT 865.950 639.600 868.050 640.050 ;
        RECT 814.950 638.400 831.600 639.000 ;
        RECT 859.950 638.400 868.050 639.600 ;
        RECT 814.950 637.950 817.050 638.400 ;
        RECT 859.950 637.950 862.050 638.400 ;
        RECT 865.950 637.950 868.050 638.400 ;
        RECT 235.950 636.600 238.050 637.050 ;
        RECT 361.950 636.600 364.050 637.050 ;
        RECT 448.950 636.600 451.050 637.050 ;
        RECT 235.950 635.400 451.050 636.600 ;
        RECT 235.950 634.950 238.050 635.400 ;
        RECT 361.950 634.950 364.050 635.400 ;
        RECT 448.950 634.950 451.050 635.400 ;
        RECT 490.950 636.600 493.050 637.050 ;
        RECT 499.950 636.600 502.050 637.050 ;
        RECT 538.950 636.600 541.050 637.050 ;
        RECT 490.950 635.400 541.050 636.600 ;
        RECT 490.950 634.950 493.050 635.400 ;
        RECT 499.950 634.950 502.050 635.400 ;
        RECT 538.950 634.950 541.050 635.400 ;
        RECT 604.950 636.600 607.050 637.050 ;
        RECT 655.950 636.600 658.050 637.050 ;
        RECT 604.950 635.400 658.050 636.600 ;
        RECT 604.950 634.950 607.050 635.400 ;
        RECT 655.950 634.950 658.050 635.400 ;
        RECT 205.950 633.600 208.050 634.050 ;
        RECT 211.950 633.600 214.050 634.050 ;
        RECT 205.950 632.400 214.050 633.600 ;
        RECT 205.950 631.950 208.050 632.400 ;
        RECT 211.950 631.950 214.050 632.400 ;
        RECT 259.950 633.600 262.050 634.050 ;
        RECT 265.950 633.600 268.050 634.050 ;
        RECT 280.950 633.600 283.050 634.050 ;
        RECT 259.950 632.400 283.050 633.600 ;
        RECT 259.950 631.950 262.050 632.400 ;
        RECT 265.950 631.950 268.050 632.400 ;
        RECT 280.950 631.950 283.050 632.400 ;
        RECT 304.950 633.600 307.050 634.050 ;
        RECT 358.950 633.600 361.050 634.050 ;
        RECT 304.950 632.400 361.050 633.600 ;
        RECT 304.950 631.950 307.050 632.400 ;
        RECT 358.950 631.950 361.050 632.400 ;
        RECT 406.950 633.600 409.050 634.050 ;
        RECT 421.950 633.600 424.050 634.050 ;
        RECT 406.950 632.400 424.050 633.600 ;
        RECT 406.950 631.950 409.050 632.400 ;
        RECT 421.950 631.950 424.050 632.400 ;
        RECT 667.950 633.600 670.050 634.050 ;
        RECT 745.950 633.600 748.050 634.050 ;
        RECT 802.950 633.600 805.050 634.050 ;
        RECT 667.950 632.400 805.050 633.600 ;
        RECT 667.950 631.950 670.050 632.400 ;
        RECT 745.950 631.950 748.050 632.400 ;
        RECT 802.950 631.950 805.050 632.400 ;
        RECT 85.950 630.600 88.050 631.050 ;
        RECT 97.950 630.600 100.050 631.050 ;
        RECT 85.950 629.400 100.050 630.600 ;
        RECT 85.950 628.950 88.050 629.400 ;
        RECT 97.950 628.950 100.050 629.400 ;
        RECT 244.950 630.600 247.050 631.050 ;
        RECT 301.950 630.600 304.050 631.050 ;
        RECT 244.950 629.400 304.050 630.600 ;
        RECT 244.950 628.950 247.050 629.400 ;
        RECT 301.950 628.950 304.050 629.400 ;
        RECT 403.950 630.600 406.050 631.050 ;
        RECT 436.950 630.600 439.050 631.050 ;
        RECT 403.950 629.400 439.050 630.600 ;
        RECT 403.950 628.950 406.050 629.400 ;
        RECT 436.950 628.950 439.050 629.400 ;
        RECT 448.950 630.600 451.050 631.050 ;
        RECT 496.950 630.600 499.050 631.050 ;
        RECT 538.950 630.600 541.050 631.050 ;
        RECT 448.950 629.400 541.050 630.600 ;
        RECT 448.950 628.950 451.050 629.400 ;
        RECT 496.950 628.950 499.050 629.400 ;
        RECT 538.950 628.950 541.050 629.400 ;
        RECT 547.950 630.600 550.050 631.050 ;
        RECT 586.950 630.600 589.050 631.050 ;
        RECT 547.950 629.400 618.600 630.600 ;
        RECT 547.950 628.950 550.050 629.400 ;
        RECT 586.950 628.950 589.050 629.400 ;
        RECT 334.950 627.600 337.050 628.050 ;
        RECT 400.950 627.600 403.050 628.050 ;
        RECT 334.950 626.400 403.050 627.600 ;
        RECT 334.950 625.950 337.050 626.400 ;
        RECT 400.950 625.950 403.050 626.400 ;
        RECT 463.950 627.600 466.050 628.050 ;
        RECT 478.950 627.600 481.050 628.050 ;
        RECT 505.950 627.600 508.050 628.050 ;
        RECT 463.950 626.400 508.050 627.600 ;
        RECT 463.950 625.950 466.050 626.400 ;
        RECT 478.950 625.950 481.050 626.400 ;
        RECT 505.950 625.950 508.050 626.400 ;
        RECT 541.950 627.600 544.050 628.050 ;
        RECT 598.950 627.600 601.050 628.050 ;
        RECT 541.950 626.400 601.050 627.600 ;
        RECT 617.400 627.600 618.600 629.400 ;
        RECT 688.950 627.600 691.050 628.050 ;
        RECT 766.950 627.600 769.050 628.050 ;
        RECT 775.950 627.600 778.050 628.050 ;
        RECT 617.400 626.400 778.050 627.600 ;
        RECT 541.950 625.950 544.050 626.400 ;
        RECT 598.950 625.950 601.050 626.400 ;
        RECT 688.950 625.950 691.050 626.400 ;
        RECT 766.950 625.950 769.050 626.400 ;
        RECT 775.950 625.950 778.050 626.400 ;
        RECT 55.950 624.600 58.050 625.050 ;
        RECT 61.950 624.600 64.050 625.050 ;
        RECT 55.950 623.400 64.050 624.600 ;
        RECT 55.950 622.950 58.050 623.400 ;
        RECT 61.950 622.950 64.050 623.400 ;
        RECT 253.950 624.600 256.050 625.050 ;
        RECT 385.950 624.600 388.050 625.050 ;
        RECT 535.950 624.600 538.050 625.050 ;
        RECT 601.950 624.600 604.050 625.050 ;
        RECT 253.950 623.400 604.050 624.600 ;
        RECT 253.950 622.950 256.050 623.400 ;
        RECT 385.950 622.950 388.050 623.400 ;
        RECT 535.950 622.950 538.050 623.400 ;
        RECT 601.950 622.950 604.050 623.400 ;
        RECT 694.950 624.600 697.050 625.050 ;
        RECT 715.950 624.600 718.050 625.050 ;
        RECT 694.950 623.400 718.050 624.600 ;
        RECT 694.950 622.950 697.050 623.400 ;
        RECT 715.950 622.950 718.050 623.400 ;
        RECT 412.950 621.600 415.050 622.050 ;
        RECT 475.950 621.600 478.050 622.050 ;
        RECT 412.950 620.400 478.050 621.600 ;
        RECT 412.950 619.950 415.050 620.400 ;
        RECT 475.950 619.950 478.050 620.400 ;
        RECT 493.950 621.600 496.050 622.050 ;
        RECT 550.950 621.600 553.050 622.050 ;
        RECT 493.950 620.400 553.050 621.600 ;
        RECT 493.950 619.950 496.050 620.400 ;
        RECT 550.950 619.950 553.050 620.400 ;
        RECT 577.950 621.600 580.050 622.050 ;
        RECT 595.950 621.600 598.050 622.050 ;
        RECT 577.950 620.400 598.050 621.600 ;
        RECT 577.950 619.950 580.050 620.400 ;
        RECT 595.950 619.950 598.050 620.400 ;
        RECT 631.950 621.600 634.050 622.050 ;
        RECT 646.950 621.600 649.050 622.050 ;
        RECT 631.950 620.400 649.050 621.600 ;
        RECT 631.950 619.950 634.050 620.400 ;
        RECT 646.950 619.950 649.050 620.400 ;
        RECT 703.950 621.600 706.050 622.050 ;
        RECT 820.950 621.600 823.050 622.050 ;
        RECT 703.950 620.400 823.050 621.600 ;
        RECT 703.950 619.950 706.050 620.400 ;
        RECT 820.950 619.950 823.050 620.400 ;
        RECT 16.950 618.600 19.050 619.050 ;
        RECT 55.950 618.600 58.050 619.050 ;
        RECT 16.950 617.400 58.050 618.600 ;
        RECT 16.950 616.950 19.050 617.400 ;
        RECT 55.950 616.950 58.050 617.400 ;
        RECT 136.950 618.600 139.050 619.050 ;
        RECT 166.950 618.600 169.050 619.050 ;
        RECT 190.950 618.600 193.050 619.050 ;
        RECT 217.950 618.600 220.050 619.050 ;
        RECT 247.950 618.600 250.050 619.050 ;
        RECT 334.950 618.600 337.050 619.050 ;
        RECT 136.950 617.400 337.050 618.600 ;
        RECT 136.950 616.950 139.050 617.400 ;
        RECT 166.950 616.950 169.050 617.400 ;
        RECT 190.950 616.950 193.050 617.400 ;
        RECT 217.950 616.950 220.050 617.400 ;
        RECT 247.950 616.950 250.050 617.400 ;
        RECT 334.950 616.950 337.050 617.400 ;
        RECT 607.950 618.600 610.050 619.050 ;
        RECT 622.950 618.600 625.050 619.050 ;
        RECT 607.950 617.400 625.050 618.600 ;
        RECT 607.950 616.950 610.050 617.400 ;
        RECT 622.950 616.950 625.050 617.400 ;
        RECT 673.950 618.600 676.050 619.050 ;
        RECT 787.950 618.600 790.050 619.050 ;
        RECT 673.950 617.400 790.050 618.600 ;
        RECT 673.950 616.950 676.050 617.400 ;
        RECT 787.950 616.950 790.050 617.400 ;
        RECT 340.950 615.600 343.050 616.050 ;
        RECT 370.950 615.600 373.050 616.050 ;
        RECT 340.950 614.400 373.050 615.600 ;
        RECT 340.950 613.950 343.050 614.400 ;
        RECT 370.950 613.950 373.050 614.400 ;
        RECT 442.950 615.600 445.050 616.050 ;
        RECT 478.950 615.600 481.050 616.050 ;
        RECT 442.950 614.400 481.050 615.600 ;
        RECT 442.950 613.950 445.050 614.400 ;
        RECT 478.950 613.950 481.050 614.400 ;
        RECT 487.950 615.600 490.050 616.050 ;
        RECT 511.950 615.600 514.050 616.050 ;
        RECT 487.950 614.400 514.050 615.600 ;
        RECT 487.950 613.950 490.050 614.400 ;
        RECT 511.950 613.950 514.050 614.400 ;
        RECT 598.950 615.600 601.050 616.050 ;
        RECT 670.950 615.600 673.050 616.050 ;
        RECT 598.950 614.400 673.050 615.600 ;
        RECT 598.950 613.950 601.050 614.400 ;
        RECT 670.950 613.950 673.050 614.400 ;
        RECT 685.950 615.600 688.050 616.050 ;
        RECT 718.950 615.600 721.050 616.050 ;
        RECT 685.950 614.400 721.050 615.600 ;
        RECT 685.950 613.950 688.050 614.400 ;
        RECT 718.950 613.950 721.050 614.400 ;
        RECT 790.950 615.600 793.050 616.050 ;
        RECT 862.950 615.600 865.050 616.050 ;
        RECT 790.950 614.400 865.050 615.600 ;
        RECT 790.950 613.950 793.050 614.400 ;
        RECT 862.950 613.950 865.050 614.400 ;
        RECT 70.950 612.600 73.050 613.050 ;
        RECT 100.950 612.600 103.050 613.050 ;
        RECT 70.950 611.400 103.050 612.600 ;
        RECT 70.950 610.950 73.050 611.400 ;
        RECT 100.950 610.950 103.050 611.400 ;
        RECT 184.950 612.600 187.050 613.050 ;
        RECT 235.950 612.600 238.050 613.050 ;
        RECT 184.950 611.400 238.050 612.600 ;
        RECT 184.950 610.950 187.050 611.400 ;
        RECT 235.950 610.950 238.050 611.400 ;
        RECT 412.950 612.600 415.050 613.050 ;
        RECT 433.950 612.600 436.050 613.050 ;
        RECT 412.950 611.400 436.050 612.600 ;
        RECT 412.950 610.950 415.050 611.400 ;
        RECT 433.950 610.950 436.050 611.400 ;
        RECT 520.950 612.600 523.050 613.050 ;
        RECT 532.950 612.600 535.050 613.050 ;
        RECT 556.950 612.600 559.050 613.050 ;
        RECT 520.950 611.400 559.050 612.600 ;
        RECT 520.950 610.950 523.050 611.400 ;
        RECT 532.950 610.950 535.050 611.400 ;
        RECT 556.950 610.950 559.050 611.400 ;
        RECT 595.950 612.600 598.050 613.050 ;
        RECT 643.950 612.600 646.050 613.050 ;
        RECT 652.950 612.600 655.050 613.050 ;
        RECT 595.950 611.400 655.050 612.600 ;
        RECT 595.950 610.950 598.050 611.400 ;
        RECT 643.950 610.950 646.050 611.400 ;
        RECT 652.950 610.950 655.050 611.400 ;
        RECT 676.950 612.600 679.050 613.050 ;
        RECT 748.950 612.600 751.050 613.050 ;
        RECT 676.950 611.400 751.050 612.600 ;
        RECT 676.950 610.950 679.050 611.400 ;
        RECT 748.950 610.950 751.050 611.400 ;
        RECT 204.000 609.600 208.050 610.050 ;
        RECT 203.400 607.950 208.050 609.600 ;
        RECT 22.950 606.600 25.050 607.200 ;
        RECT 28.950 606.600 31.050 607.050 ;
        RECT 34.950 606.600 37.050 607.200 ;
        RECT 22.950 605.400 37.050 606.600 ;
        RECT 22.950 605.100 25.050 605.400 ;
        RECT 28.950 604.950 31.050 605.400 ;
        RECT 34.950 605.100 37.050 605.400 ;
        RECT 40.950 605.100 43.050 607.200 ;
        RECT 85.950 606.600 88.050 607.200 ;
        RECT 106.950 606.600 109.050 607.200 ;
        RECT 85.950 605.400 109.050 606.600 ;
        RECT 85.950 605.100 88.050 605.400 ;
        RECT 106.950 605.100 109.050 605.400 ;
        RECT 115.950 606.600 118.050 607.200 ;
        RECT 121.950 606.750 124.050 607.200 ;
        RECT 127.950 606.750 130.050 607.200 ;
        RECT 115.950 605.400 120.600 606.600 ;
        RECT 115.950 605.100 118.050 605.400 ;
        RECT 41.400 603.600 42.600 605.100 ;
        RECT 119.400 603.600 120.600 605.400 ;
        RECT 121.950 605.550 130.050 606.750 ;
        RECT 121.950 605.100 124.050 605.550 ;
        RECT 127.950 605.100 130.050 605.550 ;
        RECT 133.950 605.100 136.050 607.200 ;
        RECT 157.950 606.600 160.050 607.200 ;
        RECT 203.400 607.050 204.600 607.950 ;
        RECT 155.400 605.400 160.050 606.600 ;
        RECT 134.400 603.600 135.600 605.100 ;
        RECT 151.950 603.600 154.050 604.050 ;
        RECT 41.400 602.400 57.600 603.600 ;
        RECT 119.400 602.400 154.050 603.600 ;
        RECT 28.950 600.450 31.050 600.900 ;
        RECT 52.950 600.450 55.050 600.900 ;
        RECT 28.950 599.250 55.050 600.450 ;
        RECT 56.400 600.600 57.600 602.400 ;
        RECT 151.950 601.950 154.050 602.400 ;
        RECT 155.400 601.050 156.600 605.400 ;
        RECT 157.950 605.100 160.050 605.400 ;
        RECT 199.950 605.400 204.600 607.050 ;
        RECT 208.950 606.600 211.050 607.200 ;
        RECT 208.950 605.400 240.600 606.600 ;
        RECT 199.950 604.950 204.000 605.400 ;
        RECT 208.950 605.100 211.050 605.400 ;
        RECT 64.950 600.600 67.050 601.050 ;
        RECT 56.400 599.400 67.050 600.600 ;
        RECT 28.950 598.800 31.050 599.250 ;
        RECT 52.950 598.800 55.050 599.250 ;
        RECT 64.950 598.950 67.050 599.400 ;
        RECT 154.950 598.950 157.050 601.050 ;
        RECT 226.950 600.600 229.050 601.050 ;
        RECT 239.400 600.900 240.600 605.400 ;
        RECT 241.950 605.100 244.050 607.200 ;
        RECT 256.950 606.750 259.050 607.200 ;
        RECT 262.950 606.750 265.050 607.200 ;
        RECT 256.950 605.550 265.050 606.750 ;
        RECT 256.950 605.100 259.050 605.550 ;
        RECT 262.950 605.100 265.050 605.550 ;
        RECT 283.950 606.750 286.050 607.200 ;
        RECT 289.950 606.750 292.050 607.200 ;
        RECT 283.950 605.550 292.050 606.750 ;
        RECT 283.950 605.100 286.050 605.550 ;
        RECT 289.950 605.100 292.050 605.550 ;
        RECT 301.950 605.100 304.050 607.200 ;
        RECT 325.950 605.100 328.050 607.200 ;
        RECT 352.950 606.600 355.050 607.200 ;
        RECT 388.950 606.600 391.050 610.050 ;
        RECT 442.950 609.600 445.050 610.050 ;
        RECT 469.950 609.600 472.050 610.050 ;
        RECT 442.950 608.400 472.050 609.600 ;
        RECT 442.950 607.950 445.050 608.400 ;
        RECT 469.950 607.950 472.050 608.400 ;
        RECT 484.950 609.600 487.050 610.050 ;
        RECT 517.950 609.600 520.050 610.050 ;
        RECT 484.950 608.400 520.050 609.600 ;
        RECT 484.950 607.950 487.050 608.400 ;
        RECT 517.950 607.950 520.050 608.400 ;
        RECT 529.950 609.600 532.050 610.050 ;
        RECT 559.950 609.600 562.050 610.050 ;
        RECT 529.950 608.400 562.050 609.600 ;
        RECT 529.950 607.950 532.050 608.400 ;
        RECT 559.950 607.950 562.050 608.400 ;
        RECT 565.950 609.600 568.050 610.050 ;
        RECT 583.950 609.600 586.050 610.050 ;
        RECT 565.950 608.400 586.050 609.600 ;
        RECT 565.950 607.950 568.050 608.400 ;
        RECT 583.950 607.950 586.050 608.400 ;
        RECT 664.950 609.600 667.050 610.050 ;
        RECT 673.950 609.600 676.050 610.050 ;
        RECT 775.950 609.600 778.050 610.050 ;
        RECT 829.950 609.600 832.050 610.050 ;
        RECT 664.950 608.400 676.050 609.600 ;
        RECT 664.950 607.950 667.050 608.400 ;
        RECT 673.950 607.950 676.050 608.400 ;
        RECT 770.400 608.400 778.050 609.600 ;
        RECT 352.950 606.000 391.050 606.600 ;
        RECT 400.950 606.600 403.050 607.200 ;
        RECT 415.950 606.600 418.050 607.050 ;
        RECT 442.950 606.600 445.050 607.200 ;
        RECT 352.950 605.400 390.600 606.000 ;
        RECT 400.950 605.400 418.050 606.600 ;
        RECT 352.950 605.100 355.050 605.400 ;
        RECT 232.950 600.600 235.050 600.900 ;
        RECT 226.950 599.400 235.050 600.600 ;
        RECT 226.950 598.950 229.050 599.400 ;
        RECT 232.950 598.800 235.050 599.400 ;
        RECT 238.950 598.800 241.050 600.900 ;
        RECT 242.400 600.600 243.600 605.100 ;
        RECT 302.400 601.050 303.600 605.100 ;
        RECT 277.950 600.600 280.050 601.050 ;
        RECT 242.400 599.400 280.050 600.600 ;
        RECT 302.400 599.400 307.050 601.050 ;
        RECT 277.950 598.950 280.050 599.400 ;
        RECT 303.000 598.950 307.050 599.400 ;
        RECT 37.950 597.600 40.050 598.050 ;
        RECT 46.950 597.600 49.050 598.050 ;
        RECT 37.950 596.400 49.050 597.600 ;
        RECT 37.950 595.950 40.050 596.400 ;
        RECT 46.950 595.950 49.050 596.400 ;
        RECT 112.950 597.600 115.050 598.050 ;
        RECT 121.950 597.600 124.050 598.050 ;
        RECT 139.950 597.600 142.050 598.050 ;
        RECT 112.950 596.400 142.050 597.600 ;
        RECT 326.400 597.600 327.600 605.100 ;
        RECT 371.400 603.600 372.600 605.400 ;
        RECT 400.950 605.100 403.050 605.400 ;
        RECT 415.950 604.950 418.050 605.400 ;
        RECT 419.400 605.400 445.050 606.600 ;
        RECT 419.400 603.600 420.600 605.400 ;
        RECT 442.950 605.100 445.050 605.400 ;
        RECT 448.950 606.750 451.050 607.200 ;
        RECT 457.950 606.750 460.050 607.200 ;
        RECT 448.950 605.550 460.050 606.750 ;
        RECT 448.950 605.100 451.050 605.550 ;
        RECT 457.950 605.100 460.050 605.550 ;
        RECT 475.950 604.950 478.050 607.050 ;
        RECT 495.000 606.600 499.050 607.050 ;
        RECT 494.400 604.950 499.050 606.600 ;
        RECT 502.950 604.950 505.050 607.050 ;
        RECT 577.950 604.950 580.050 607.050 ;
        RECT 595.950 604.950 598.050 607.050 ;
        RECT 604.950 605.100 607.050 607.200 ;
        RECT 610.950 605.100 613.050 607.200 ;
        RECT 658.950 606.600 661.050 607.200 ;
        RECT 676.950 606.600 679.050 607.200 ;
        RECT 658.950 605.400 679.050 606.600 ;
        RECT 658.950 605.100 661.050 605.400 ;
        RECT 676.950 605.100 679.050 605.400 ;
        RECT 682.950 606.750 685.050 607.200 ;
        RECT 688.950 606.750 691.050 607.200 ;
        RECT 682.950 605.550 691.050 606.750 ;
        RECT 712.950 606.600 715.050 607.200 ;
        RECT 682.950 605.100 685.050 605.550 ;
        RECT 688.950 605.100 691.050 605.550 ;
        RECT 692.400 605.400 715.050 606.600 ;
        RECT 371.400 602.400 420.600 603.600 ;
        RECT 340.950 600.450 343.050 600.900 ;
        RECT 367.950 600.450 370.050 600.900 ;
        RECT 340.950 599.250 370.050 600.450 ;
        RECT 340.950 598.800 343.050 599.250 ;
        RECT 367.950 598.800 370.050 599.250 ;
        RECT 418.950 600.600 421.050 601.050 ;
        RECT 427.950 600.600 430.050 600.900 ;
        RECT 418.950 599.400 430.050 600.600 ;
        RECT 418.950 598.950 421.050 599.400 ;
        RECT 427.950 598.800 430.050 599.400 ;
        RECT 436.950 600.600 439.050 601.050 ;
        RECT 445.950 600.600 448.050 600.900 ;
        RECT 436.950 599.400 448.050 600.600 ;
        RECT 436.950 598.950 439.050 599.400 ;
        RECT 445.950 598.800 448.050 599.400 ;
        RECT 451.950 600.600 454.050 600.900 ;
        RECT 466.950 600.600 469.050 600.900 ;
        RECT 476.400 600.600 477.600 604.950 ;
        RECT 451.950 599.400 477.600 600.600 ;
        RECT 478.950 600.600 481.050 601.050 ;
        RECT 490.950 600.600 493.050 600.900 ;
        RECT 478.950 599.400 493.050 600.600 ;
        RECT 451.950 598.800 454.050 599.400 ;
        RECT 466.950 598.800 469.050 599.400 ;
        RECT 478.950 598.950 481.050 599.400 ;
        RECT 490.950 598.800 493.050 599.400 ;
        RECT 494.400 598.050 495.600 604.950 ;
        RECT 503.400 600.600 504.600 604.950 ;
        RECT 508.950 600.600 511.050 600.900 ;
        RECT 503.400 599.400 511.050 600.600 ;
        RECT 508.950 598.800 511.050 599.400 ;
        RECT 517.950 600.450 520.050 600.900 ;
        RECT 562.950 600.450 565.050 600.900 ;
        RECT 517.950 599.250 565.050 600.450 ;
        RECT 517.950 598.800 520.050 599.250 ;
        RECT 562.950 598.800 565.050 599.250 ;
        RECT 568.950 600.600 571.050 600.900 ;
        RECT 578.400 600.600 579.600 604.950 ;
        RECT 568.950 599.400 579.600 600.600 ;
        RECT 586.950 600.600 589.050 600.900 ;
        RECT 596.400 600.600 597.600 604.950 ;
        RECT 605.400 603.600 606.600 605.100 ;
        RECT 611.400 603.600 612.600 605.100 ;
        RECT 628.950 603.600 631.050 604.050 ;
        RECT 605.400 603.000 609.600 603.600 ;
        RECT 605.400 602.400 610.050 603.000 ;
        RECT 611.400 602.400 631.050 603.600 ;
        RECT 586.950 599.400 597.600 600.600 ;
        RECT 568.950 598.800 571.050 599.400 ;
        RECT 586.950 598.800 589.050 599.400 ;
        RECT 607.950 598.950 610.050 602.400 ;
        RECT 628.950 601.950 631.050 602.400 ;
        RECT 637.950 600.450 640.050 600.900 ;
        RECT 643.950 600.450 646.050 600.900 ;
        RECT 637.950 599.250 646.050 600.450 ;
        RECT 637.950 598.800 640.050 599.250 ;
        RECT 643.950 598.800 646.050 599.250 ;
        RECT 655.950 600.600 658.050 600.900 ;
        RECT 664.950 600.600 667.050 601.050 ;
        RECT 655.950 599.400 667.050 600.600 ;
        RECT 655.950 598.800 658.050 599.400 ;
        RECT 664.950 598.950 667.050 599.400 ;
        RECT 334.950 597.600 337.050 598.050 ;
        RECT 326.400 596.400 337.050 597.600 ;
        RECT 112.950 595.950 115.050 596.400 ;
        RECT 121.950 595.950 124.050 596.400 ;
        RECT 139.950 595.950 142.050 596.400 ;
        RECT 334.950 595.950 337.050 596.400 ;
        RECT 367.950 597.600 370.050 598.050 ;
        RECT 388.950 597.600 391.050 598.050 ;
        RECT 367.950 596.400 391.050 597.600 ;
        RECT 367.950 595.950 370.050 596.400 ;
        RECT 388.950 595.950 391.050 596.400 ;
        RECT 493.950 595.950 496.050 598.050 ;
        RECT 562.950 597.600 565.050 598.050 ;
        RECT 580.950 597.600 583.050 598.050 ;
        RECT 562.950 596.400 583.050 597.600 ;
        RECT 677.400 597.600 678.600 605.100 ;
        RECT 692.400 600.900 693.600 605.400 ;
        RECT 712.950 605.100 715.050 605.400 ;
        RECT 754.950 606.750 757.050 607.200 ;
        RECT 760.950 606.750 763.050 606.900 ;
        RECT 754.950 605.550 763.050 606.750 ;
        RECT 754.950 605.100 757.050 605.550 ;
        RECT 760.950 604.800 763.050 605.550 ;
        RECT 770.400 600.900 771.600 608.400 ;
        RECT 775.950 607.950 778.050 608.400 ;
        RECT 794.400 608.400 832.050 609.600 ;
        RECT 794.400 600.900 795.600 608.400 ;
        RECT 829.950 607.950 832.050 608.400 ;
        RECT 796.950 606.750 799.050 607.200 ;
        RECT 808.950 606.750 811.050 607.200 ;
        RECT 796.950 605.550 811.050 606.750 ;
        RECT 817.950 606.600 820.050 607.050 ;
        RECT 796.950 605.100 799.050 605.550 ;
        RECT 808.950 605.100 811.050 605.550 ;
        RECT 812.400 605.400 820.050 606.600 ;
        RECT 691.950 598.800 694.050 600.900 ;
        RECT 721.950 600.450 724.050 600.900 ;
        RECT 730.950 600.450 733.050 600.900 ;
        RECT 721.950 599.250 733.050 600.450 ;
        RECT 721.950 598.800 724.050 599.250 ;
        RECT 730.950 598.800 733.050 599.250 ;
        RECT 739.950 600.450 742.050 600.900 ;
        RECT 745.950 600.450 748.050 600.900 ;
        RECT 739.950 599.250 748.050 600.450 ;
        RECT 739.950 598.800 742.050 599.250 ;
        RECT 745.950 598.800 748.050 599.250 ;
        RECT 769.950 598.800 772.050 600.900 ;
        RECT 793.950 598.800 796.050 600.900 ;
        RECT 688.950 597.600 691.050 598.050 ;
        RECT 697.950 597.600 700.050 598.050 ;
        RECT 677.400 596.400 700.050 597.600 ;
        RECT 562.950 595.950 565.050 596.400 ;
        RECT 580.950 595.950 583.050 596.400 ;
        RECT 688.950 595.950 691.050 596.400 ;
        RECT 697.950 595.950 700.050 596.400 ;
        RECT 766.950 597.600 769.050 598.050 ;
        RECT 799.950 597.600 802.050 598.050 ;
        RECT 766.950 596.400 802.050 597.600 ;
        RECT 766.950 595.950 769.050 596.400 ;
        RECT 799.950 595.950 802.050 596.400 ;
        RECT 805.950 597.600 808.050 598.050 ;
        RECT 812.400 597.600 813.600 605.400 ;
        RECT 817.950 604.950 820.050 605.400 ;
        RECT 832.950 603.600 835.050 607.050 ;
        RECT 850.950 604.950 853.050 607.050 ;
        RECT 859.950 606.600 862.050 607.050 ;
        RECT 859.950 605.400 870.600 606.600 ;
        RECT 859.950 604.950 862.050 605.400 ;
        RECT 815.400 603.000 846.600 603.600 ;
        RECT 815.400 602.400 847.050 603.000 ;
        RECT 815.400 600.900 816.600 602.400 ;
        RECT 814.950 598.800 817.050 600.900 ;
        RECT 844.950 598.950 847.050 602.400 ;
        RECT 851.400 601.050 852.600 604.950 ;
        RECT 869.400 601.050 870.600 605.400 ;
        RECT 850.950 598.950 853.050 601.050 ;
        RECT 868.950 598.950 871.050 601.050 ;
        RECT 805.950 596.400 813.600 597.600 ;
        RECT 829.950 597.600 832.050 598.050 ;
        RECT 835.950 597.600 838.050 598.050 ;
        RECT 829.950 596.400 838.050 597.600 ;
        RECT 805.950 595.950 808.050 596.400 ;
        RECT 829.950 595.950 832.050 596.400 ;
        RECT 835.950 595.950 838.050 596.400 ;
        RECT 847.950 597.600 850.050 598.050 ;
        RECT 862.950 597.600 865.050 598.050 ;
        RECT 847.950 596.400 865.050 597.600 ;
        RECT 847.950 595.950 850.050 596.400 ;
        RECT 862.950 595.950 865.050 596.400 ;
        RECT 19.950 594.600 22.050 595.050 ;
        RECT 46.950 594.600 49.050 594.900 ;
        RECT 19.950 593.400 49.050 594.600 ;
        RECT 19.950 592.950 22.050 593.400 ;
        RECT 46.950 592.800 49.050 593.400 ;
        RECT 151.950 594.600 154.050 595.050 ;
        RECT 181.950 594.600 184.050 595.050 ;
        RECT 190.950 594.600 193.050 595.050 ;
        RECT 151.950 593.400 193.050 594.600 ;
        RECT 151.950 592.950 154.050 593.400 ;
        RECT 181.950 592.950 184.050 593.400 ;
        RECT 190.950 592.950 193.050 593.400 ;
        RECT 298.950 594.600 301.050 595.050 ;
        RECT 307.950 594.600 310.050 595.050 ;
        RECT 346.950 594.600 349.050 595.050 ;
        RECT 298.950 593.400 349.050 594.600 ;
        RECT 298.950 592.950 301.050 593.400 ;
        RECT 307.950 592.950 310.050 593.400 ;
        RECT 346.950 592.950 349.050 593.400 ;
        RECT 472.950 594.600 475.050 595.050 ;
        RECT 520.950 594.600 523.050 595.050 ;
        RECT 592.950 594.600 595.050 595.050 ;
        RECT 472.950 593.400 595.050 594.600 ;
        RECT 472.950 592.950 475.050 593.400 ;
        RECT 520.950 592.950 523.050 593.400 ;
        RECT 592.950 592.950 595.050 593.400 ;
        RECT 673.950 594.600 676.050 595.050 ;
        RECT 682.950 594.600 685.050 595.050 ;
        RECT 673.950 593.400 685.050 594.600 ;
        RECT 673.950 592.950 676.050 593.400 ;
        RECT 682.950 592.950 685.050 593.400 ;
        RECT 718.950 594.600 721.050 595.050 ;
        RECT 751.950 594.600 754.050 595.050 ;
        RECT 718.950 593.400 754.050 594.600 ;
        RECT 718.950 592.950 721.050 593.400 ;
        RECT 751.950 592.950 754.050 593.400 ;
        RECT 484.950 591.600 487.050 592.050 ;
        RECT 499.950 591.600 502.050 592.050 ;
        RECT 484.950 590.400 502.050 591.600 ;
        RECT 484.950 589.950 487.050 590.400 ;
        RECT 499.950 589.950 502.050 590.400 ;
        RECT 583.950 591.600 586.050 592.050 ;
        RECT 589.950 591.600 592.050 592.050 ;
        RECT 583.950 590.400 592.050 591.600 ;
        RECT 583.950 589.950 586.050 590.400 ;
        RECT 589.950 589.950 592.050 590.400 ;
        RECT 595.950 591.600 598.050 592.050 ;
        RECT 619.950 591.600 622.050 592.050 ;
        RECT 595.950 590.400 622.050 591.600 ;
        RECT 595.950 589.950 598.050 590.400 ;
        RECT 619.950 589.950 622.050 590.400 ;
        RECT 625.950 591.600 628.050 592.050 ;
        RECT 637.950 591.600 640.050 592.050 ;
        RECT 625.950 590.400 640.050 591.600 ;
        RECT 625.950 589.950 628.050 590.400 ;
        RECT 637.950 589.950 640.050 590.400 ;
        RECT 73.950 588.600 76.050 589.050 ;
        RECT 85.950 588.600 88.050 589.050 ;
        RECT 97.950 588.600 100.050 589.050 ;
        RECT 103.950 588.600 106.050 589.050 ;
        RECT 109.950 588.600 112.050 589.050 ;
        RECT 73.950 587.400 112.050 588.600 ;
        RECT 73.950 586.950 76.050 587.400 ;
        RECT 85.950 586.950 88.050 587.400 ;
        RECT 97.950 586.950 100.050 587.400 ;
        RECT 103.950 586.950 106.050 587.400 ;
        RECT 109.950 586.950 112.050 587.400 ;
        RECT 181.950 588.600 184.050 589.050 ;
        RECT 199.950 588.600 202.050 589.050 ;
        RECT 181.950 587.400 202.050 588.600 ;
        RECT 181.950 586.950 184.050 587.400 ;
        RECT 199.950 586.950 202.050 587.400 ;
        RECT 262.950 588.600 265.050 589.050 ;
        RECT 271.950 588.600 274.050 589.050 ;
        RECT 262.950 587.400 274.050 588.600 ;
        RECT 262.950 586.950 265.050 587.400 ;
        RECT 271.950 586.950 274.050 587.400 ;
        RECT 283.950 588.600 286.050 589.050 ;
        RECT 349.950 588.600 352.050 589.050 ;
        RECT 364.950 588.600 367.050 589.050 ;
        RECT 283.950 587.400 367.050 588.600 ;
        RECT 283.950 586.950 286.050 587.400 ;
        RECT 349.950 586.950 352.050 587.400 ;
        RECT 364.950 586.950 367.050 587.400 ;
        RECT 505.950 588.600 508.050 589.050 ;
        RECT 523.950 588.600 526.050 589.050 ;
        RECT 559.950 588.600 562.050 589.050 ;
        RECT 505.950 587.400 562.050 588.600 ;
        RECT 505.950 586.950 508.050 587.400 ;
        RECT 523.950 586.950 526.050 587.400 ;
        RECT 559.950 586.950 562.050 587.400 ;
        RECT 592.950 588.600 595.050 589.050 ;
        RECT 634.950 588.600 637.050 589.050 ;
        RECT 592.950 587.400 637.050 588.600 ;
        RECT 592.950 586.950 595.050 587.400 ;
        RECT 634.950 586.950 637.050 587.400 ;
        RECT 727.950 588.600 730.050 589.050 ;
        RECT 736.950 588.600 739.050 589.050 ;
        RECT 727.950 587.400 739.050 588.600 ;
        RECT 727.950 586.950 730.050 587.400 ;
        RECT 736.950 586.950 739.050 587.400 ;
        RECT 784.950 588.600 787.050 589.050 ;
        RECT 802.950 588.600 805.050 589.050 ;
        RECT 784.950 587.400 805.050 588.600 ;
        RECT 784.950 586.950 787.050 587.400 ;
        RECT 802.950 586.950 805.050 587.400 ;
        RECT 838.950 588.600 841.050 589.050 ;
        RECT 850.950 588.600 853.050 589.050 ;
        RECT 838.950 587.400 853.050 588.600 ;
        RECT 838.950 586.950 841.050 587.400 ;
        RECT 850.950 586.950 853.050 587.400 ;
        RECT 34.950 585.600 37.050 586.050 ;
        RECT 43.950 585.600 46.050 586.050 ;
        RECT 52.950 585.600 55.050 586.050 ;
        RECT 34.950 584.400 55.050 585.600 ;
        RECT 34.950 583.950 37.050 584.400 ;
        RECT 43.950 583.950 46.050 584.400 ;
        RECT 52.950 583.950 55.050 584.400 ;
        RECT 238.950 585.600 241.050 586.050 ;
        RECT 292.950 585.600 295.050 586.050 ;
        RECT 238.950 584.400 295.050 585.600 ;
        RECT 238.950 583.950 241.050 584.400 ;
        RECT 292.950 583.950 295.050 584.400 ;
        RECT 307.950 585.600 310.050 586.050 ;
        RECT 319.950 585.600 322.050 586.050 ;
        RECT 307.950 584.400 322.050 585.600 ;
        RECT 307.950 583.950 310.050 584.400 ;
        RECT 319.950 583.950 322.050 584.400 ;
        RECT 457.950 585.600 460.050 586.050 ;
        RECT 520.950 585.600 523.050 586.050 ;
        RECT 457.950 584.400 523.050 585.600 ;
        RECT 457.950 583.950 460.050 584.400 ;
        RECT 520.950 583.950 523.050 584.400 ;
        RECT 601.950 585.600 604.050 586.050 ;
        RECT 607.950 585.600 610.050 586.050 ;
        RECT 601.950 584.400 610.050 585.600 ;
        RECT 601.950 583.950 604.050 584.400 ;
        RECT 607.950 583.950 610.050 584.400 ;
        RECT 748.950 585.600 751.050 586.050 ;
        RECT 760.950 585.600 763.050 586.050 ;
        RECT 748.950 584.400 763.050 585.600 ;
        RECT 748.950 583.950 751.050 584.400 ;
        RECT 760.950 583.950 763.050 584.400 ;
        RECT 826.950 585.600 829.050 586.050 ;
        RECT 835.950 585.600 838.050 586.050 ;
        RECT 826.950 584.400 838.050 585.600 ;
        RECT 826.950 583.950 829.050 584.400 ;
        RECT 835.950 583.950 838.050 584.400 ;
        RECT 58.950 582.600 61.050 583.050 ;
        RECT 73.950 582.600 76.050 583.050 ;
        RECT 58.950 581.400 76.050 582.600 ;
        RECT 58.950 580.950 61.050 581.400 ;
        RECT 73.950 580.950 76.050 581.400 ;
        RECT 79.950 582.600 82.050 583.050 ;
        RECT 91.950 582.600 94.050 583.050 ;
        RECT 103.950 582.600 106.050 583.050 ;
        RECT 130.950 582.600 133.050 583.050 ;
        RECT 79.950 581.400 133.050 582.600 ;
        RECT 79.950 580.950 82.050 581.400 ;
        RECT 91.950 580.950 94.050 581.400 ;
        RECT 103.950 580.950 106.050 581.400 ;
        RECT 130.950 580.950 133.050 581.400 ;
        RECT 193.950 582.600 196.050 583.050 ;
        RECT 211.950 582.600 214.050 583.050 ;
        RECT 193.950 581.400 214.050 582.600 ;
        RECT 193.950 580.950 196.050 581.400 ;
        RECT 211.950 580.950 214.050 581.400 ;
        RECT 241.950 582.600 244.050 583.050 ;
        RECT 265.950 582.600 268.050 583.050 ;
        RECT 241.950 581.400 268.050 582.600 ;
        RECT 241.950 580.950 244.050 581.400 ;
        RECT 265.950 580.950 268.050 581.400 ;
        RECT 355.950 582.600 358.050 583.050 ;
        RECT 433.950 582.600 436.050 583.050 ;
        RECT 355.950 581.400 436.050 582.600 ;
        RECT 355.950 580.950 358.050 581.400 ;
        RECT 433.950 580.950 436.050 581.400 ;
        RECT 451.950 582.600 454.050 583.050 ;
        RECT 463.950 582.600 466.050 583.050 ;
        RECT 505.950 582.600 508.050 583.050 ;
        RECT 451.950 581.400 508.050 582.600 ;
        RECT 451.950 580.950 454.050 581.400 ;
        RECT 463.950 580.950 466.050 581.400 ;
        RECT 505.950 580.950 508.050 581.400 ;
        RECT 574.950 582.600 577.050 583.050 ;
        RECT 586.950 582.600 589.050 583.050 ;
        RECT 574.950 581.400 589.050 582.600 ;
        RECT 574.950 580.950 577.050 581.400 ;
        RECT 586.950 580.950 589.050 581.400 ;
        RECT 787.950 582.600 790.050 583.050 ;
        RECT 814.950 582.600 817.050 583.050 ;
        RECT 787.950 581.400 817.050 582.600 ;
        RECT 787.950 580.950 790.050 581.400 ;
        RECT 814.950 580.950 817.050 581.400 ;
        RECT 856.950 582.600 859.050 583.050 ;
        RECT 865.950 582.600 868.050 583.050 ;
        RECT 856.950 581.400 868.050 582.600 ;
        RECT 856.950 580.950 859.050 581.400 ;
        RECT 865.950 580.950 868.050 581.400 ;
        RECT 37.950 579.600 40.050 580.050 ;
        RECT 43.950 579.600 46.050 580.050 ;
        RECT 37.950 578.400 46.050 579.600 ;
        RECT 37.950 577.950 40.050 578.400 ;
        RECT 43.950 577.950 46.050 578.400 ;
        RECT 106.950 579.600 109.050 580.050 ;
        RECT 115.950 579.600 118.050 580.050 ;
        RECT 106.950 578.400 118.050 579.600 ;
        RECT 106.950 577.950 109.050 578.400 ;
        RECT 115.950 577.950 118.050 578.400 ;
        RECT 124.950 579.600 127.050 580.050 ;
        RECT 148.950 579.600 151.050 580.050 ;
        RECT 157.950 579.600 160.050 580.050 ;
        RECT 124.950 578.400 160.050 579.600 ;
        RECT 124.950 577.950 127.050 578.400 ;
        RECT 148.950 577.950 151.050 578.400 ;
        RECT 157.950 577.950 160.050 578.400 ;
        RECT 190.950 579.600 193.050 580.050 ;
        RECT 238.950 579.600 241.050 580.050 ;
        RECT 190.950 578.400 241.050 579.600 ;
        RECT 190.950 577.950 193.050 578.400 ;
        RECT 238.950 577.950 241.050 578.400 ;
        RECT 274.950 579.600 277.050 580.050 ;
        RECT 295.950 579.600 298.050 580.050 ;
        RECT 274.950 578.400 298.050 579.600 ;
        RECT 274.950 577.950 277.050 578.400 ;
        RECT 295.950 577.950 298.050 578.400 ;
        RECT 610.950 579.600 613.050 580.050 ;
        RECT 775.950 579.600 778.050 580.050 ;
        RECT 784.950 579.600 787.050 580.050 ;
        RECT 610.950 578.400 648.600 579.600 ;
        RECT 610.950 577.950 613.050 578.400 ;
        RECT 647.400 577.050 648.600 578.400 ;
        RECT 775.950 578.400 787.050 579.600 ;
        RECT 775.950 577.950 778.050 578.400 ;
        RECT 784.950 577.950 787.050 578.400 ;
        RECT 46.950 576.600 49.050 577.050 ;
        RECT 67.950 576.600 70.050 577.050 ;
        RECT 172.950 576.600 175.050 577.050 ;
        RECT 46.950 575.400 70.050 576.600 ;
        RECT 46.950 574.950 49.050 575.400 ;
        RECT 67.950 574.950 70.050 575.400 ;
        RECT 92.400 575.400 175.050 576.600 ;
        RECT 22.950 573.750 25.050 574.200 ;
        RECT 28.950 573.750 31.050 574.200 ;
        RECT 22.950 572.550 31.050 573.750 ;
        RECT 22.950 572.100 25.050 572.550 ;
        RECT 28.950 572.100 31.050 572.550 ;
        RECT 58.950 571.950 61.050 574.050 ;
        RECT 64.950 571.950 67.050 574.050 ;
        RECT 85.950 573.600 88.050 574.050 ;
        RECT 92.400 573.600 93.600 575.400 ;
        RECT 172.950 574.950 175.050 575.400 ;
        RECT 71.400 572.400 88.050 573.600 ;
        RECT 59.400 568.050 60.600 571.950 ;
        RECT 65.400 568.050 66.600 571.950 ;
        RECT 16.950 567.600 19.050 567.900 ;
        RECT 22.950 567.600 25.050 568.050 ;
        RECT 16.950 566.400 25.050 567.600 ;
        RECT 16.950 565.800 19.050 566.400 ;
        RECT 22.950 565.950 25.050 566.400 ;
        RECT 37.950 567.450 40.050 567.900 ;
        RECT 43.950 567.450 46.050 567.900 ;
        RECT 37.950 566.250 46.050 567.450 ;
        RECT 37.950 565.800 40.050 566.250 ;
        RECT 43.950 565.800 46.050 566.250 ;
        RECT 58.950 565.950 61.050 568.050 ;
        RECT 64.950 565.950 67.050 568.050 ;
        RECT 71.400 567.900 72.600 572.400 ;
        RECT 85.950 571.950 88.050 572.400 ;
        RECT 89.400 572.400 93.600 573.600 ;
        RECT 100.950 573.600 103.050 574.050 ;
        RECT 133.950 573.600 136.050 574.200 ;
        RECT 142.950 573.600 145.050 574.050 ;
        RECT 100.950 572.400 132.600 573.600 ;
        RECT 89.400 567.900 90.600 572.400 ;
        RECT 100.950 571.950 103.050 572.400 ;
        RECT 131.400 570.600 132.600 572.400 ;
        RECT 133.950 572.400 145.050 573.600 ;
        RECT 133.950 572.100 136.050 572.400 ;
        RECT 142.950 571.950 145.050 572.400 ;
        RECT 178.950 573.600 181.050 574.050 ;
        RECT 193.950 573.600 196.050 574.050 ;
        RECT 178.950 572.400 196.050 573.600 ;
        RECT 178.950 571.950 181.050 572.400 ;
        RECT 193.950 571.950 196.050 572.400 ;
        RECT 199.950 573.750 202.050 574.200 ;
        RECT 205.950 573.750 208.050 574.200 ;
        RECT 199.950 572.550 208.050 573.750 ;
        RECT 217.950 573.600 220.050 577.050 ;
        RECT 373.950 576.600 376.050 577.050 ;
        RECT 379.950 576.600 382.050 577.050 ;
        RECT 373.950 575.400 382.050 576.600 ;
        RECT 373.950 574.950 376.050 575.400 ;
        RECT 379.950 574.950 382.050 575.400 ;
        RECT 415.950 574.950 418.050 577.050 ;
        RECT 592.950 576.600 595.050 577.050 ;
        RECT 613.950 576.600 616.050 577.050 ;
        RECT 592.950 575.400 616.050 576.600 ;
        RECT 592.950 574.950 595.050 575.400 ;
        RECT 613.950 574.950 616.050 575.400 ;
        RECT 229.950 573.600 232.050 574.200 ;
        RECT 217.950 573.000 232.050 573.600 ;
        RECT 199.950 572.100 202.050 572.550 ;
        RECT 205.950 572.100 208.050 572.550 ;
        RECT 218.400 572.400 232.050 573.000 ;
        RECT 229.950 572.100 232.050 572.400 ;
        RECT 280.950 573.750 283.050 574.200 ;
        RECT 289.950 573.750 292.050 574.200 ;
        RECT 280.950 572.550 292.050 573.750 ;
        RECT 280.950 572.100 283.050 572.550 ;
        RECT 289.950 572.100 292.050 572.550 ;
        RECT 295.950 572.100 298.050 574.200 ;
        RECT 313.950 573.600 316.050 574.200 ;
        RECT 322.950 573.750 325.050 574.200 ;
        RECT 328.950 573.750 331.050 574.200 ;
        RECT 313.950 572.400 321.600 573.600 ;
        RECT 313.950 572.100 316.050 572.400 ;
        RECT 296.400 570.600 297.600 572.100 ;
        RECT 131.400 569.400 135.600 570.600 ;
        RECT 296.400 569.400 309.600 570.600 ;
        RECT 70.950 565.800 73.050 567.900 ;
        RECT 88.950 565.800 91.050 567.900 ;
        RECT 124.950 567.450 127.050 567.900 ;
        RECT 130.950 567.450 133.050 567.900 ;
        RECT 124.950 566.250 133.050 567.450 ;
        RECT 124.950 565.800 127.050 566.250 ;
        RECT 130.950 565.800 133.050 566.250 ;
        RECT 134.400 565.050 135.600 569.400 ;
        RECT 142.950 567.450 145.050 567.900 ;
        RECT 148.950 567.450 151.050 567.900 ;
        RECT 142.950 566.250 151.050 567.450 ;
        RECT 142.950 565.800 145.050 566.250 ;
        RECT 148.950 565.800 151.050 566.250 ;
        RECT 172.950 567.450 175.050 567.900 ;
        RECT 178.950 567.450 181.050 567.900 ;
        RECT 172.950 566.250 181.050 567.450 ;
        RECT 172.950 565.800 175.050 566.250 ;
        RECT 178.950 565.800 181.050 566.250 ;
        RECT 199.950 567.600 202.050 568.050 ;
        RECT 226.950 567.600 229.050 567.900 ;
        RECT 199.950 566.400 229.050 567.600 ;
        RECT 199.950 565.950 202.050 566.400 ;
        RECT 226.950 565.800 229.050 566.400 ;
        RECT 232.950 567.600 235.050 567.900 ;
        RECT 238.950 567.600 241.050 568.050 ;
        RECT 232.950 566.400 241.050 567.600 ;
        RECT 232.950 565.800 235.050 566.400 ;
        RECT 238.950 565.950 241.050 566.400 ;
        RECT 292.950 567.600 295.050 567.900 ;
        RECT 301.950 567.600 304.050 568.050 ;
        RECT 292.950 566.400 304.050 567.600 ;
        RECT 308.400 567.600 309.600 569.400 ;
        RECT 320.400 568.050 321.600 572.400 ;
        RECT 322.950 572.550 331.050 573.750 ;
        RECT 339.000 573.600 343.050 574.050 ;
        RECT 322.950 572.100 325.050 572.550 ;
        RECT 328.950 572.100 331.050 572.550 ;
        RECT 338.400 571.950 343.050 573.600 ;
        RECT 346.950 571.950 349.050 574.050 ;
        RECT 361.950 573.750 364.050 574.200 ;
        RECT 367.950 573.750 370.050 574.200 ;
        RECT 361.950 572.550 370.050 573.750 ;
        RECT 361.950 572.100 364.050 572.550 ;
        RECT 367.950 572.100 370.050 572.550 ;
        RECT 310.950 567.600 313.050 567.900 ;
        RECT 308.400 566.400 313.050 567.600 ;
        RECT 292.950 565.800 295.050 566.400 ;
        RECT 301.950 565.950 304.050 566.400 ;
        RECT 310.950 565.800 313.050 566.400 ;
        RECT 319.950 565.950 322.050 568.050 ;
        RECT 338.400 567.900 339.600 571.950 ;
        RECT 337.950 565.800 340.050 567.900 ;
        RECT 347.400 567.600 348.600 571.950 ;
        RECT 416.400 567.900 417.600 574.950 ;
        RECT 442.950 573.750 445.050 574.200 ;
        RECT 460.950 573.750 463.050 574.200 ;
        RECT 442.950 572.550 463.050 573.750 ;
        RECT 442.950 572.100 445.050 572.550 ;
        RECT 460.950 572.100 463.050 572.550 ;
        RECT 505.950 573.600 508.050 574.050 ;
        RECT 514.950 573.600 517.050 574.200 ;
        RECT 505.950 572.400 517.050 573.600 ;
        RECT 505.950 571.950 508.050 572.400 ;
        RECT 514.950 572.100 517.050 572.400 ;
        RECT 523.950 572.100 526.050 574.200 ;
        RECT 556.950 573.600 559.050 574.050 ;
        RECT 568.950 573.600 571.050 574.200 ;
        RECT 556.950 572.400 571.050 573.600 ;
        RECT 349.950 567.600 352.050 567.900 ;
        RECT 347.400 566.400 352.050 567.600 ;
        RECT 349.950 565.800 352.050 566.400 ;
        RECT 391.950 567.450 394.050 567.900 ;
        RECT 397.950 567.450 400.050 567.900 ;
        RECT 391.950 566.250 400.050 567.450 ;
        RECT 391.950 565.800 394.050 566.250 ;
        RECT 397.950 565.800 400.050 566.250 ;
        RECT 406.950 567.600 409.050 567.900 ;
        RECT 415.950 567.600 418.050 567.900 ;
        RECT 406.950 566.400 418.050 567.600 ;
        RECT 406.950 565.800 409.050 566.400 ;
        RECT 415.950 565.800 418.050 566.400 ;
        RECT 424.950 567.450 427.050 567.900 ;
        RECT 430.950 567.450 433.050 567.900 ;
        RECT 424.950 566.250 433.050 567.450 ;
        RECT 424.950 565.800 427.050 566.250 ;
        RECT 430.950 565.800 433.050 566.250 ;
        RECT 460.950 567.450 463.050 567.900 ;
        RECT 469.950 567.450 472.050 567.900 ;
        RECT 460.950 566.250 472.050 567.450 ;
        RECT 460.950 565.800 463.050 566.250 ;
        RECT 469.950 565.800 472.050 566.250 ;
        RECT 499.950 567.600 502.050 567.900 ;
        RECT 511.950 567.600 514.050 567.900 ;
        RECT 499.950 566.400 514.050 567.600 ;
        RECT 499.950 565.800 502.050 566.400 ;
        RECT 511.950 565.800 514.050 566.400 ;
        RECT 517.950 567.600 520.050 567.900 ;
        RECT 524.400 567.600 525.600 572.100 ;
        RECT 556.950 571.950 559.050 572.400 ;
        RECT 568.950 572.100 571.050 572.400 ;
        RECT 574.950 573.600 577.050 574.200 ;
        RECT 580.950 573.750 583.050 574.200 ;
        RECT 586.950 573.750 589.050 574.200 ;
        RECT 580.950 573.600 589.050 573.750 ;
        RECT 597.000 573.600 601.050 574.050 ;
        RECT 574.950 572.550 589.050 573.600 ;
        RECT 574.950 572.400 583.050 572.550 ;
        RECT 574.950 572.100 577.050 572.400 ;
        RECT 580.950 572.100 583.050 572.400 ;
        RECT 586.950 572.100 589.050 572.550 ;
        RECT 596.400 571.950 601.050 573.600 ;
        RECT 619.950 573.600 622.050 577.050 ;
        RECT 628.950 576.600 631.050 577.050 ;
        RECT 640.950 576.600 643.050 577.050 ;
        RECT 628.950 575.400 643.050 576.600 ;
        RECT 628.950 574.950 631.050 575.400 ;
        RECT 640.950 574.950 643.050 575.400 ;
        RECT 646.950 576.600 649.050 577.050 ;
        RECT 697.950 576.600 700.050 577.050 ;
        RECT 852.000 576.600 856.050 577.050 ;
        RECT 646.950 575.400 700.050 576.600 ;
        RECT 646.950 574.950 649.050 575.400 ;
        RECT 697.950 574.950 700.050 575.400 ;
        RECT 851.400 574.950 856.050 576.600 ;
        RECT 649.950 573.600 652.050 574.050 ;
        RECT 619.950 573.000 652.050 573.600 ;
        RECT 620.400 572.400 652.050 573.000 ;
        RECT 649.950 571.950 652.050 572.400 ;
        RECT 691.950 573.600 694.050 574.050 ;
        RECT 703.950 573.600 706.050 574.200 ;
        RECT 691.950 572.400 706.050 573.600 ;
        RECT 691.950 571.950 694.050 572.400 ;
        RECT 703.950 572.100 706.050 572.400 ;
        RECT 712.950 573.600 715.050 574.050 ;
        RECT 721.950 573.600 724.050 574.200 ;
        RECT 712.950 572.400 724.050 573.600 ;
        RECT 712.950 571.950 715.050 572.400 ;
        RECT 721.950 572.100 724.050 572.400 ;
        RECT 727.950 571.950 730.050 574.050 ;
        RECT 745.950 573.750 748.050 574.200 ;
        RECT 757.950 573.750 760.050 574.200 ;
        RECT 745.950 572.550 760.050 573.750 ;
        RECT 745.950 572.100 748.050 572.550 ;
        RECT 757.950 572.100 760.050 572.550 ;
        RECT 769.950 573.750 772.050 574.200 ;
        RECT 778.950 573.750 781.050 574.200 ;
        RECT 769.950 572.550 781.050 573.750 ;
        RECT 769.950 572.100 772.050 572.550 ;
        RECT 778.950 572.100 781.050 572.550 ;
        RECT 796.950 572.100 799.050 574.200 ;
        RECT 596.400 567.900 597.600 571.950 ;
        RECT 728.400 568.050 729.600 571.950 ;
        RECT 517.950 566.400 525.600 567.600 ;
        RECT 541.950 567.450 544.050 567.900 ;
        RECT 556.950 567.450 559.050 567.900 ;
        RECT 517.950 565.800 520.050 566.400 ;
        RECT 541.950 566.250 559.050 567.450 ;
        RECT 541.950 565.800 544.050 566.250 ;
        RECT 556.950 565.800 559.050 566.250 ;
        RECT 595.950 565.800 598.050 567.900 ;
        RECT 613.950 567.450 616.050 567.900 ;
        RECT 619.950 567.450 622.050 567.900 ;
        RECT 613.950 566.250 622.050 567.450 ;
        RECT 613.950 565.800 616.050 566.250 ;
        RECT 619.950 565.800 622.050 566.250 ;
        RECT 628.950 567.600 631.050 567.900 ;
        RECT 640.950 567.600 643.050 568.050 ;
        RECT 664.950 567.600 667.050 567.900 ;
        RECT 673.950 567.600 676.050 568.050 ;
        RECT 628.950 566.400 676.050 567.600 ;
        RECT 628.950 565.800 631.050 566.400 ;
        RECT 640.950 565.950 643.050 566.400 ;
        RECT 664.950 565.800 667.050 566.400 ;
        RECT 673.950 565.950 676.050 566.400 ;
        RECT 691.950 567.450 694.050 567.900 ;
        RECT 700.950 567.450 703.050 567.900 ;
        RECT 691.950 566.250 703.050 567.450 ;
        RECT 691.950 565.800 694.050 566.250 ;
        RECT 700.950 565.800 703.050 566.250 ;
        RECT 706.950 567.450 709.050 567.900 ;
        RECT 712.950 567.450 715.050 567.900 ;
        RECT 706.950 566.250 715.050 567.450 ;
        RECT 706.950 565.800 709.050 566.250 ;
        RECT 712.950 565.800 715.050 566.250 ;
        RECT 727.950 565.950 730.050 568.050 ;
        RECT 763.950 567.450 766.050 567.900 ;
        RECT 772.950 567.450 775.050 567.900 ;
        RECT 763.950 566.250 775.050 567.450 ;
        RECT 763.950 565.800 766.050 566.250 ;
        RECT 772.950 565.800 775.050 566.250 ;
        RECT 103.950 564.600 106.050 565.050 ;
        RECT 118.950 564.600 121.050 565.050 ;
        RECT 103.950 563.400 121.050 564.600 ;
        RECT 103.950 562.950 106.050 563.400 ;
        RECT 118.950 562.950 121.050 563.400 ;
        RECT 133.950 562.950 136.050 565.050 ;
        RECT 286.950 564.600 289.050 565.050 ;
        RECT 307.950 564.600 310.050 565.050 ;
        RECT 286.950 563.400 310.050 564.600 ;
        RECT 286.950 562.950 289.050 563.400 ;
        RECT 307.950 562.950 310.050 563.400 ;
        RECT 358.950 564.600 361.050 565.050 ;
        RECT 373.950 564.600 376.050 565.050 ;
        RECT 358.950 563.400 376.050 564.600 ;
        RECT 358.950 562.950 361.050 563.400 ;
        RECT 373.950 562.950 376.050 563.400 ;
        RECT 643.950 564.600 646.050 565.050 ;
        RECT 649.950 564.600 652.050 565.050 ;
        RECT 643.950 563.400 652.050 564.600 ;
        RECT 643.950 562.950 646.050 563.400 ;
        RECT 649.950 562.950 652.050 563.400 ;
        RECT 700.950 564.600 703.050 565.050 ;
        RECT 718.950 564.600 721.050 565.050 ;
        RECT 700.950 563.400 721.050 564.600 ;
        RECT 700.950 562.950 703.050 563.400 ;
        RECT 718.950 562.950 721.050 563.400 ;
        RECT 724.950 564.600 727.050 565.050 ;
        RECT 745.950 564.600 748.050 565.050 ;
        RECT 760.950 564.600 763.050 565.050 ;
        RECT 724.950 563.400 763.050 564.600 ;
        RECT 797.400 564.600 798.600 572.100 ;
        RECT 805.950 571.950 808.050 574.050 ;
        RECT 811.950 573.750 814.050 574.200 ;
        RECT 820.950 573.750 823.050 574.200 ;
        RECT 811.950 572.550 823.050 573.750 ;
        RECT 811.950 572.100 814.050 572.550 ;
        RECT 820.950 572.100 823.050 572.550 ;
        RECT 806.400 567.600 807.600 571.950 ;
        RECT 851.400 568.050 852.600 574.950 ;
        RECT 856.950 572.100 859.050 574.200 ;
        RECT 817.950 567.600 820.050 567.900 ;
        RECT 806.400 566.400 820.050 567.600 ;
        RECT 817.950 565.800 820.050 566.400 ;
        RECT 850.950 565.950 853.050 568.050 ;
        RECT 808.950 564.600 811.050 565.050 ;
        RECT 797.400 563.400 811.050 564.600 ;
        RECT 724.950 562.950 727.050 563.400 ;
        RECT 745.950 562.950 748.050 563.400 ;
        RECT 760.950 562.950 763.050 563.400 ;
        RECT 808.950 562.950 811.050 563.400 ;
        RECT 28.950 561.600 31.050 562.050 ;
        RECT 46.950 561.600 49.050 562.050 ;
        RECT 28.950 560.400 49.050 561.600 ;
        RECT 28.950 559.950 31.050 560.400 ;
        RECT 46.950 559.950 49.050 560.400 ;
        RECT 55.950 561.600 58.050 562.050 ;
        RECT 94.950 561.600 97.050 562.050 ;
        RECT 55.950 560.400 97.050 561.600 ;
        RECT 55.950 559.950 58.050 560.400 ;
        RECT 94.950 559.950 97.050 560.400 ;
        RECT 127.950 561.600 130.050 562.050 ;
        RECT 136.950 561.600 139.050 562.050 ;
        RECT 127.950 560.400 139.050 561.600 ;
        RECT 127.950 559.950 130.050 560.400 ;
        RECT 136.950 559.950 139.050 560.400 ;
        RECT 289.950 561.600 292.050 562.050 ;
        RECT 298.950 561.600 301.050 562.050 ;
        RECT 289.950 560.400 301.050 561.600 ;
        RECT 289.950 559.950 292.050 560.400 ;
        RECT 298.950 559.950 301.050 560.400 ;
        RECT 316.950 561.600 319.050 562.050 ;
        RECT 322.950 561.600 325.050 562.050 ;
        RECT 355.950 561.600 358.050 562.050 ;
        RECT 511.950 561.600 514.050 562.050 ;
        RECT 580.950 561.600 583.050 562.050 ;
        RECT 316.950 560.400 583.050 561.600 ;
        RECT 316.950 559.950 319.050 560.400 ;
        RECT 322.950 559.950 325.050 560.400 ;
        RECT 355.950 559.950 358.050 560.400 ;
        RECT 511.950 559.950 514.050 560.400 ;
        RECT 580.950 559.950 583.050 560.400 ;
        RECT 685.950 561.600 688.050 562.050 ;
        RECT 766.950 561.600 769.050 562.050 ;
        RECT 685.950 560.400 769.050 561.600 ;
        RECT 685.950 559.950 688.050 560.400 ;
        RECT 766.950 559.950 769.050 560.400 ;
        RECT 772.950 561.600 775.050 562.050 ;
        RECT 799.950 561.600 802.050 562.050 ;
        RECT 772.950 560.400 802.050 561.600 ;
        RECT 772.950 559.950 775.050 560.400 ;
        RECT 799.950 559.950 802.050 560.400 ;
        RECT 814.950 561.600 817.050 562.050 ;
        RECT 826.950 561.600 829.050 562.050 ;
        RECT 814.950 560.400 829.050 561.600 ;
        RECT 857.400 561.600 858.600 572.100 ;
        RECT 859.950 567.450 862.050 567.900 ;
        RECT 868.950 567.450 871.050 567.900 ;
        RECT 859.950 566.250 871.050 567.450 ;
        RECT 859.950 565.800 862.050 566.250 ;
        RECT 868.950 565.800 871.050 566.250 ;
        RECT 868.950 561.600 871.050 562.050 ;
        RECT 857.400 560.400 871.050 561.600 ;
        RECT 814.950 559.950 817.050 560.400 ;
        RECT 826.950 559.950 829.050 560.400 ;
        RECT 868.950 559.950 871.050 560.400 ;
        RECT 235.950 558.600 238.050 559.050 ;
        RECT 280.950 558.600 283.050 559.050 ;
        RECT 235.950 557.400 283.050 558.600 ;
        RECT 235.950 556.950 238.050 557.400 ;
        RECT 280.950 556.950 283.050 557.400 ;
        RECT 517.950 558.600 520.050 559.050 ;
        RECT 550.950 558.600 553.050 559.050 ;
        RECT 571.950 558.600 574.050 559.050 ;
        RECT 517.950 557.400 574.050 558.600 ;
        RECT 517.950 556.950 520.050 557.400 ;
        RECT 550.950 556.950 553.050 557.400 ;
        RECT 571.950 556.950 574.050 557.400 ;
        RECT 613.950 558.600 616.050 559.050 ;
        RECT 634.950 558.600 637.050 559.050 ;
        RECT 613.950 557.400 637.050 558.600 ;
        RECT 613.950 556.950 616.050 557.400 ;
        RECT 634.950 556.950 637.050 557.400 ;
        RECT 673.950 558.600 676.050 559.050 ;
        RECT 730.950 558.600 733.050 559.050 ;
        RECT 673.950 557.400 733.050 558.600 ;
        RECT 673.950 556.950 676.050 557.400 ;
        RECT 730.950 556.950 733.050 557.400 ;
        RECT 10.950 555.600 13.050 556.050 ;
        RECT 31.950 555.600 34.050 556.050 ;
        RECT 10.950 554.400 34.050 555.600 ;
        RECT 10.950 553.950 13.050 554.400 ;
        RECT 31.950 553.950 34.050 554.400 ;
        RECT 79.950 555.600 82.050 556.050 ;
        RECT 154.950 555.600 157.050 556.050 ;
        RECT 79.950 554.400 157.050 555.600 ;
        RECT 79.950 553.950 82.050 554.400 ;
        RECT 154.950 553.950 157.050 554.400 ;
        RECT 226.950 555.600 229.050 556.050 ;
        RECT 229.950 555.600 232.050 556.050 ;
        RECT 259.950 555.600 262.050 556.050 ;
        RECT 226.950 554.400 262.050 555.600 ;
        RECT 226.950 553.950 229.050 554.400 ;
        RECT 229.950 553.950 232.050 554.400 ;
        RECT 259.950 553.950 262.050 554.400 ;
        RECT 274.950 555.600 277.050 556.050 ;
        RECT 319.950 555.600 322.050 556.050 ;
        RECT 274.950 554.400 322.050 555.600 ;
        RECT 274.950 553.950 277.050 554.400 ;
        RECT 319.950 553.950 322.050 554.400 ;
        RECT 505.950 555.600 508.050 556.050 ;
        RECT 565.950 555.600 568.050 556.050 ;
        RECT 505.950 554.400 568.050 555.600 ;
        RECT 505.950 553.950 508.050 554.400 ;
        RECT 565.950 553.950 568.050 554.400 ;
        RECT 574.950 555.600 577.050 556.050 ;
        RECT 637.950 555.600 640.050 556.050 ;
        RECT 574.950 554.400 640.050 555.600 ;
        RECT 574.950 553.950 577.050 554.400 ;
        RECT 637.950 553.950 640.050 554.400 ;
        RECT 694.950 555.600 697.050 556.050 ;
        RECT 742.950 555.600 745.050 556.050 ;
        RECT 694.950 554.400 745.050 555.600 ;
        RECT 694.950 553.950 697.050 554.400 ;
        RECT 742.950 553.950 745.050 554.400 ;
        RECT 760.950 555.600 763.050 556.050 ;
        RECT 835.950 555.600 838.050 556.050 ;
        RECT 760.950 554.400 838.050 555.600 ;
        RECT 760.950 553.950 763.050 554.400 ;
        RECT 835.950 553.950 838.050 554.400 ;
        RECT 181.950 552.600 184.050 553.050 ;
        RECT 187.950 552.600 190.050 553.050 ;
        RECT 181.950 551.400 190.050 552.600 ;
        RECT 181.950 550.950 184.050 551.400 ;
        RECT 187.950 550.950 190.050 551.400 ;
        RECT 283.950 552.600 286.050 553.050 ;
        RECT 310.950 552.600 313.050 553.050 ;
        RECT 283.950 551.400 313.050 552.600 ;
        RECT 283.950 550.950 286.050 551.400 ;
        RECT 310.950 550.950 313.050 551.400 ;
        RECT 361.950 552.600 364.050 553.050 ;
        RECT 463.950 552.600 466.050 553.050 ;
        RECT 361.950 551.400 466.050 552.600 ;
        RECT 361.950 550.950 364.050 551.400 ;
        RECT 463.950 550.950 466.050 551.400 ;
        RECT 571.950 552.600 574.050 553.050 ;
        RECT 628.800 552.600 630.900 553.050 ;
        RECT 571.950 551.400 630.900 552.600 ;
        RECT 571.950 550.950 574.050 551.400 ;
        RECT 628.800 550.950 630.900 551.400 ;
        RECT 58.950 549.600 61.050 550.050 ;
        RECT 154.950 549.600 157.050 550.050 ;
        RECT 58.950 548.400 157.050 549.600 ;
        RECT 58.950 547.950 61.050 548.400 ;
        RECT 154.950 547.950 157.050 548.400 ;
        RECT 457.950 549.600 460.050 550.050 ;
        RECT 535.950 549.600 538.050 550.050 ;
        RECT 457.950 548.400 538.050 549.600 ;
        RECT 457.950 547.950 460.050 548.400 ;
        RECT 535.950 547.950 538.050 548.400 ;
        RECT 727.950 549.600 730.050 550.050 ;
        RECT 748.950 549.600 751.050 550.050 ;
        RECT 727.950 548.400 751.050 549.600 ;
        RECT 727.950 547.950 730.050 548.400 ;
        RECT 748.950 547.950 751.050 548.400 ;
        RECT 766.950 549.600 769.050 550.050 ;
        RECT 841.950 549.600 844.050 550.050 ;
        RECT 853.950 549.600 856.050 550.050 ;
        RECT 766.950 548.400 856.050 549.600 ;
        RECT 766.950 547.950 769.050 548.400 ;
        RECT 841.950 547.950 844.050 548.400 ;
        RECT 853.950 547.950 856.050 548.400 ;
        RECT 223.950 546.600 226.050 547.050 ;
        RECT 256.950 546.600 259.050 547.050 ;
        RECT 223.950 545.400 259.050 546.600 ;
        RECT 223.950 544.950 226.050 545.400 ;
        RECT 256.950 544.950 259.050 545.400 ;
        RECT 298.950 546.600 301.050 547.050 ;
        RECT 364.950 546.600 367.050 547.050 ;
        RECT 298.950 545.400 367.050 546.600 ;
        RECT 298.950 544.950 301.050 545.400 ;
        RECT 364.950 544.950 367.050 545.400 ;
        RECT 472.950 546.600 475.050 547.050 ;
        RECT 478.950 546.600 481.050 547.050 ;
        RECT 517.950 546.600 520.050 547.050 ;
        RECT 472.950 545.400 520.050 546.600 ;
        RECT 472.950 544.950 475.050 545.400 ;
        RECT 478.950 544.950 481.050 545.400 ;
        RECT 517.950 544.950 520.050 545.400 ;
        RECT 589.950 546.600 592.050 547.050 ;
        RECT 607.950 546.600 610.050 547.050 ;
        RECT 589.950 545.400 610.050 546.600 ;
        RECT 589.950 544.950 592.050 545.400 ;
        RECT 607.950 544.950 610.050 545.400 ;
        RECT 625.950 546.600 628.050 547.050 ;
        RECT 676.950 546.600 679.050 547.050 ;
        RECT 700.950 546.600 703.050 547.050 ;
        RECT 625.950 545.400 703.050 546.600 ;
        RECT 625.950 544.950 628.050 545.400 ;
        RECT 676.950 544.950 679.050 545.400 ;
        RECT 700.950 544.950 703.050 545.400 ;
        RECT 760.950 546.600 763.050 547.050 ;
        RECT 871.950 546.600 874.050 547.050 ;
        RECT 760.950 545.400 874.050 546.600 ;
        RECT 760.950 544.950 763.050 545.400 ;
        RECT 871.950 544.950 874.050 545.400 ;
        RECT 1.950 543.600 4.050 544.050 ;
        RECT 79.950 543.600 82.050 544.050 ;
        RECT 1.950 542.400 82.050 543.600 ;
        RECT 1.950 541.950 4.050 542.400 ;
        RECT 79.950 541.950 82.050 542.400 ;
        RECT 259.950 543.600 262.050 544.050 ;
        RECT 265.950 543.600 268.050 544.050 ;
        RECT 358.950 543.600 361.050 544.050 ;
        RECT 259.950 542.400 361.050 543.600 ;
        RECT 259.950 541.950 262.050 542.400 ;
        RECT 265.950 541.950 268.050 542.400 ;
        RECT 358.950 541.950 361.050 542.400 ;
        RECT 85.950 540.600 88.050 541.050 ;
        RECT 103.950 540.600 106.050 541.050 ;
        RECT 85.950 539.400 106.050 540.600 ;
        RECT 85.950 538.950 88.050 539.400 ;
        RECT 103.950 538.950 106.050 539.400 ;
        RECT 151.950 540.600 154.050 541.050 ;
        RECT 181.950 540.600 184.050 541.050 ;
        RECT 151.950 539.400 184.050 540.600 ;
        RECT 151.950 538.950 154.050 539.400 ;
        RECT 181.950 538.950 184.050 539.400 ;
        RECT 244.950 540.600 247.050 541.050 ;
        RECT 331.950 540.600 334.050 541.050 ;
        RECT 244.950 539.400 334.050 540.600 ;
        RECT 244.950 538.950 247.050 539.400 ;
        RECT 331.950 538.950 334.050 539.400 ;
        RECT 502.950 540.600 505.050 541.050 ;
        RECT 604.950 540.600 607.050 541.050 ;
        RECT 502.950 539.400 607.050 540.600 ;
        RECT 502.950 538.950 505.050 539.400 ;
        RECT 604.950 538.950 607.050 539.400 ;
        RECT 622.950 540.600 625.050 541.050 ;
        RECT 628.950 540.600 631.050 541.050 ;
        RECT 622.950 539.400 631.050 540.600 ;
        RECT 622.950 538.950 625.050 539.400 ;
        RECT 628.950 538.950 631.050 539.400 ;
        RECT 634.950 540.600 637.050 541.050 ;
        RECT 691.950 540.600 694.050 541.050 ;
        RECT 634.950 539.400 694.050 540.600 ;
        RECT 634.950 538.950 637.050 539.400 ;
        RECT 691.950 538.950 694.050 539.400 ;
        RECT 709.950 540.600 712.050 541.050 ;
        RECT 766.950 540.600 769.050 541.050 ;
        RECT 796.950 540.600 799.050 541.050 ;
        RECT 709.950 539.400 799.050 540.600 ;
        RECT 709.950 538.950 712.050 539.400 ;
        RECT 766.950 538.950 769.050 539.400 ;
        RECT 796.950 538.950 799.050 539.400 ;
        RECT 106.950 537.600 109.050 538.050 ;
        RECT 148.950 537.600 151.050 538.050 ;
        RECT 106.950 536.400 151.050 537.600 ;
        RECT 106.950 535.950 109.050 536.400 ;
        RECT 148.950 535.950 151.050 536.400 ;
        RECT 160.950 537.600 163.050 538.050 ;
        RECT 169.950 537.600 172.050 538.050 ;
        RECT 160.950 536.400 172.050 537.600 ;
        RECT 160.950 535.950 163.050 536.400 ;
        RECT 169.950 535.950 172.050 536.400 ;
        RECT 196.950 537.600 199.050 538.050 ;
        RECT 238.950 537.600 241.050 538.050 ;
        RECT 196.950 536.400 241.050 537.600 ;
        RECT 196.950 535.950 199.050 536.400 ;
        RECT 238.950 535.950 241.050 536.400 ;
        RECT 256.950 537.600 259.050 538.050 ;
        RECT 361.950 537.600 364.050 538.050 ;
        RECT 256.950 536.400 364.050 537.600 ;
        RECT 256.950 535.950 259.050 536.400 ;
        RECT 361.950 535.950 364.050 536.400 ;
        RECT 433.950 537.600 436.050 538.050 ;
        RECT 454.950 537.600 457.050 538.050 ;
        RECT 433.950 536.400 457.050 537.600 ;
        RECT 433.950 535.950 436.050 536.400 ;
        RECT 454.950 535.950 457.050 536.400 ;
        RECT 559.950 537.600 562.050 538.050 ;
        RECT 625.950 537.600 628.050 538.050 ;
        RECT 559.950 536.400 628.050 537.600 ;
        RECT 559.950 535.950 562.050 536.400 ;
        RECT 625.950 535.950 628.050 536.400 ;
        RECT 712.950 537.600 715.050 538.050 ;
        RECT 802.950 537.600 805.050 538.050 ;
        RECT 838.950 537.600 841.050 538.050 ;
        RECT 712.950 536.400 805.050 537.600 ;
        RECT 712.950 535.950 715.050 536.400 ;
        RECT 802.950 535.950 805.050 536.400 ;
        RECT 830.400 536.400 841.050 537.600 ;
        RECT 64.950 534.600 67.050 535.050 ;
        RECT 79.950 534.600 82.050 535.050 ;
        RECT 139.950 534.600 142.050 535.050 ;
        RECT 64.950 533.400 142.050 534.600 ;
        RECT 64.950 532.950 67.050 533.400 ;
        RECT 79.950 532.950 82.050 533.400 ;
        RECT 139.950 532.950 142.050 533.400 ;
        RECT 481.950 534.600 484.050 535.050 ;
        RECT 535.950 534.600 538.050 535.050 ;
        RECT 481.950 533.400 538.050 534.600 ;
        RECT 481.950 532.950 484.050 533.400 ;
        RECT 535.950 532.950 538.050 533.400 ;
        RECT 547.950 534.600 550.050 535.050 ;
        RECT 556.950 534.600 559.050 535.050 ;
        RECT 547.950 533.400 559.050 534.600 ;
        RECT 547.950 532.950 550.050 533.400 ;
        RECT 556.950 532.950 559.050 533.400 ;
        RECT 565.950 534.600 568.050 535.050 ;
        RECT 610.950 534.600 613.050 535.050 ;
        RECT 565.950 533.400 613.050 534.600 ;
        RECT 565.950 532.950 568.050 533.400 ;
        RECT 610.950 532.950 613.050 533.400 ;
        RECT 673.950 534.600 676.050 535.050 ;
        RECT 688.950 534.600 691.050 535.050 ;
        RECT 709.950 534.600 712.050 535.050 ;
        RECT 673.950 533.400 712.050 534.600 ;
        RECT 673.950 532.950 676.050 533.400 ;
        RECT 688.950 532.950 691.050 533.400 ;
        RECT 709.950 532.950 712.050 533.400 ;
        RECT 736.950 534.600 739.050 535.050 ;
        RECT 760.950 534.600 763.050 535.050 ;
        RECT 736.950 533.400 763.050 534.600 ;
        RECT 736.950 532.950 739.050 533.400 ;
        RECT 760.950 532.950 763.050 533.400 ;
        RECT 778.950 534.600 781.050 535.050 ;
        RECT 830.400 534.600 831.600 536.400 ;
        RECT 838.950 535.950 841.050 536.400 ;
        RECT 778.950 533.400 831.600 534.600 ;
        RECT 832.950 534.600 835.050 535.050 ;
        RECT 841.950 534.600 844.050 535.050 ;
        RECT 832.950 533.400 844.050 534.600 ;
        RECT 778.950 532.950 781.050 533.400 ;
        RECT 832.950 532.950 835.050 533.400 ;
        RECT 841.950 532.950 844.050 533.400 ;
        RECT 46.950 531.600 49.050 532.050 ;
        RECT 52.950 531.600 55.050 532.050 ;
        RECT 97.950 531.600 100.050 532.050 ;
        RECT 163.950 531.600 166.050 532.050 ;
        RECT 190.950 531.600 193.050 532.050 ;
        RECT 196.950 531.600 199.050 532.050 ;
        RECT 46.950 530.400 199.050 531.600 ;
        RECT 46.950 529.950 49.050 530.400 ;
        RECT 52.950 529.950 55.050 530.400 ;
        RECT 97.950 529.950 100.050 530.400 ;
        RECT 163.950 529.950 166.050 530.400 ;
        RECT 190.950 529.950 193.050 530.400 ;
        RECT 196.950 529.950 199.050 530.400 ;
        RECT 370.950 531.600 373.050 532.050 ;
        RECT 388.950 531.600 391.050 532.050 ;
        RECT 406.950 531.600 409.050 532.050 ;
        RECT 370.950 530.400 409.050 531.600 ;
        RECT 370.950 529.950 373.050 530.400 ;
        RECT 388.950 529.950 391.050 530.400 ;
        RECT 406.950 529.950 409.050 530.400 ;
        RECT 523.950 531.600 526.050 532.050 ;
        RECT 532.950 531.600 535.050 532.050 ;
        RECT 523.950 530.400 535.050 531.600 ;
        RECT 523.950 529.950 526.050 530.400 ;
        RECT 532.950 529.950 535.050 530.400 ;
        RECT 574.950 531.600 577.050 532.050 ;
        RECT 592.950 531.600 595.050 532.050 ;
        RECT 574.950 530.400 595.050 531.600 ;
        RECT 574.950 529.950 577.050 530.400 ;
        RECT 592.950 529.950 595.050 530.400 ;
        RECT 634.950 531.600 637.050 532.050 ;
        RECT 640.950 531.600 643.050 532.050 ;
        RECT 829.950 531.600 832.050 532.050 ;
        RECT 844.950 531.600 847.050 531.900 ;
        RECT 634.950 530.400 643.050 531.600 ;
        RECT 634.950 529.950 637.050 530.400 ;
        RECT 640.950 529.950 643.050 530.400 ;
        RECT 764.400 530.400 783.600 531.600 ;
        RECT 7.950 526.950 10.050 529.050 ;
        RECT 16.950 528.600 19.050 529.050 ;
        RECT 31.950 528.600 34.050 529.050 ;
        RECT 16.950 527.400 34.050 528.600 ;
        RECT 16.950 526.950 19.050 527.400 ;
        RECT 31.950 526.950 34.050 527.400 ;
        RECT 37.950 527.100 40.050 529.200 ;
        RECT 64.950 528.600 67.050 529.200 ;
        RECT 115.950 528.600 118.050 529.200 ;
        RECT 64.950 527.400 118.050 528.600 ;
        RECT 64.950 527.100 67.050 527.400 ;
        RECT 115.950 527.100 118.050 527.400 ;
        RECT 121.950 528.750 124.050 529.200 ;
        RECT 127.950 528.750 130.050 529.200 ;
        RECT 121.950 527.550 130.050 528.750 ;
        RECT 121.950 527.100 124.050 527.550 ;
        RECT 127.950 527.100 130.050 527.550 ;
        RECT 8.400 523.050 9.600 526.950 ;
        RECT 7.950 520.950 10.050 523.050 ;
        RECT 38.400 520.050 39.600 527.100 ;
        RECT 151.950 526.950 154.050 529.050 ;
        RECT 175.950 528.600 178.050 529.200 ;
        RECT 170.400 527.400 178.050 528.600 ;
        RECT 61.950 522.450 64.050 522.900 ;
        RECT 67.950 522.450 70.050 522.900 ;
        RECT 61.950 521.250 70.050 522.450 ;
        RECT 61.950 520.800 64.050 521.250 ;
        RECT 67.950 520.800 70.050 521.250 ;
        RECT 103.950 522.450 106.050 522.900 ;
        RECT 118.950 522.450 121.050 522.900 ;
        RECT 103.950 521.250 121.050 522.450 ;
        RECT 103.950 520.800 106.050 521.250 ;
        RECT 118.950 520.800 121.050 521.250 ;
        RECT 142.950 522.600 145.050 522.900 ;
        RECT 152.400 522.600 153.600 526.950 ;
        RECT 142.950 521.400 153.600 522.600 ;
        RECT 163.950 522.600 166.050 522.900 ;
        RECT 170.400 522.600 171.600 527.400 ;
        RECT 175.950 527.100 178.050 527.400 ;
        RECT 238.950 528.750 241.050 529.200 ;
        RECT 247.950 528.750 250.050 529.200 ;
        RECT 238.950 528.600 250.050 528.750 ;
        RECT 274.950 528.600 277.050 529.200 ;
        RECT 238.950 527.550 277.050 528.600 ;
        RECT 238.950 527.100 241.050 527.550 ;
        RECT 247.950 527.400 277.050 527.550 ;
        RECT 247.950 527.100 250.050 527.400 ;
        RECT 274.950 527.100 277.050 527.400 ;
        RECT 280.950 528.600 283.050 529.200 ;
        RECT 298.950 528.600 301.050 529.200 ;
        RECT 280.950 527.400 301.050 528.600 ;
        RECT 280.950 527.100 283.050 527.400 ;
        RECT 298.950 527.100 301.050 527.400 ;
        RECT 319.950 528.750 322.050 529.200 ;
        RECT 325.950 528.750 328.050 529.200 ;
        RECT 319.950 528.600 328.050 528.750 ;
        RECT 334.950 528.600 337.050 529.200 ;
        RECT 319.950 527.550 337.050 528.600 ;
        RECT 319.950 527.100 322.050 527.550 ;
        RECT 325.950 527.400 337.050 527.550 ;
        RECT 325.950 527.100 328.050 527.400 ;
        RECT 334.950 527.100 337.050 527.400 ;
        RECT 340.950 528.750 343.050 529.200 ;
        RECT 346.950 528.750 349.050 529.200 ;
        RECT 340.950 527.550 349.050 528.750 ;
        RECT 340.950 527.100 343.050 527.550 ;
        RECT 346.950 527.100 349.050 527.550 ;
        RECT 358.950 528.600 361.050 529.200 ;
        RECT 364.950 528.600 367.050 529.050 ;
        RECT 370.950 528.600 373.050 529.200 ;
        RECT 358.950 527.400 373.050 528.600 ;
        RECT 358.950 527.100 361.050 527.400 ;
        RECT 364.950 526.950 367.050 527.400 ;
        RECT 370.950 527.100 373.050 527.400 ;
        RECT 376.950 528.750 379.050 529.200 ;
        RECT 382.950 528.750 385.050 529.200 ;
        RECT 376.950 527.550 385.050 528.750 ;
        RECT 376.950 527.100 379.050 527.550 ;
        RECT 382.950 527.100 385.050 527.550 ;
        RECT 394.950 528.750 397.050 529.200 ;
        RECT 400.950 528.750 403.050 529.200 ;
        RECT 394.950 527.550 403.050 528.750 ;
        RECT 394.950 527.100 397.050 527.550 ;
        RECT 400.950 527.100 403.050 527.550 ;
        RECT 412.950 527.100 415.050 529.200 ;
        RECT 418.950 527.100 421.050 529.200 ;
        RECT 427.950 528.750 430.050 529.200 ;
        RECT 433.950 528.750 436.050 529.200 ;
        RECT 427.950 527.550 436.050 528.750 ;
        RECT 427.950 527.100 430.050 527.550 ;
        RECT 433.950 527.100 436.050 527.550 ;
        RECT 454.950 528.750 457.050 529.200 ;
        RECT 463.950 528.750 466.050 529.200 ;
        RECT 454.950 527.550 466.050 528.750 ;
        RECT 454.950 527.100 457.050 527.550 ;
        RECT 463.950 527.100 466.050 527.550 ;
        RECT 508.950 527.100 511.050 529.200 ;
        RECT 541.950 527.100 544.050 529.200 ;
        RECT 598.950 527.100 601.050 529.200 ;
        RECT 413.400 523.050 414.600 527.100 ;
        RECT 163.950 521.400 171.600 522.600 ;
        RECT 262.950 522.600 265.050 522.900 ;
        RECT 262.950 521.400 267.600 522.600 ;
        RECT 142.950 520.800 145.050 521.400 ;
        RECT 163.950 520.800 166.050 521.400 ;
        RECT 262.950 520.800 265.050 521.400 ;
        RECT 10.950 519.600 13.050 520.050 ;
        RECT 19.950 519.600 22.050 520.050 ;
        RECT 10.950 518.400 22.050 519.600 ;
        RECT 10.950 517.950 13.050 518.400 ;
        RECT 19.950 517.950 22.050 518.400 ;
        RECT 37.950 517.950 40.050 520.050 ;
        RECT 178.950 519.600 181.050 520.050 ;
        RECT 241.950 519.600 244.050 520.050 ;
        RECT 178.950 518.400 244.050 519.600 ;
        RECT 266.400 519.600 267.600 521.400 ;
        RECT 277.950 522.450 280.050 522.900 ;
        RECT 286.950 522.450 289.050 522.900 ;
        RECT 277.950 521.250 289.050 522.450 ;
        RECT 277.950 520.800 280.050 521.250 ;
        RECT 286.950 520.800 289.050 521.250 ;
        RECT 301.950 522.600 304.050 522.900 ;
        RECT 325.950 522.600 328.050 523.050 ;
        RECT 301.950 521.400 328.050 522.600 ;
        RECT 301.950 520.800 304.050 521.400 ;
        RECT 325.950 520.950 328.050 521.400 ;
        RECT 352.950 522.450 355.050 522.900 ;
        RECT 361.950 522.450 364.050 522.900 ;
        RECT 352.950 521.250 364.050 522.450 ;
        RECT 413.400 521.400 418.050 523.050 ;
        RECT 352.950 520.800 355.050 521.250 ;
        RECT 361.950 520.800 364.050 521.250 ;
        RECT 414.000 520.950 418.050 521.400 ;
        RECT 277.950 519.600 280.050 520.050 ;
        RECT 266.400 518.400 280.050 519.600 ;
        RECT 178.950 517.950 181.050 518.400 ;
        RECT 241.950 517.950 244.050 518.400 ;
        RECT 277.950 517.950 280.050 518.400 ;
        RECT 385.950 519.600 388.050 520.050 ;
        RECT 419.400 519.600 420.600 527.100 ;
        RECT 445.950 522.600 448.050 522.900 ;
        RECT 454.950 522.600 457.050 523.050 ;
        RECT 445.950 521.400 457.050 522.600 ;
        RECT 445.950 520.800 448.050 521.400 ;
        RECT 454.950 520.950 457.050 521.400 ;
        RECT 484.950 522.600 487.050 522.900 ;
        RECT 490.950 522.600 493.050 522.900 ;
        RECT 484.950 521.400 493.050 522.600 ;
        RECT 509.400 522.600 510.600 527.100 ;
        RECT 542.400 525.600 543.600 527.100 ;
        RECT 542.400 524.400 558.600 525.600 ;
        RECT 532.950 522.600 535.050 522.900 ;
        RECT 509.400 521.400 535.050 522.600 ;
        RECT 557.400 522.600 558.600 524.400 ;
        RECT 599.400 523.050 600.600 527.100 ;
        RECT 607.950 526.950 610.050 529.050 ;
        RECT 619.950 528.750 622.050 529.200 ;
        RECT 658.950 528.750 661.050 529.200 ;
        RECT 619.950 527.550 661.050 528.750 ;
        RECT 667.950 528.600 670.050 529.200 ;
        RECT 685.950 528.600 688.050 529.200 ;
        RECT 619.950 527.100 622.050 527.550 ;
        RECT 658.950 527.100 661.050 527.550 ;
        RECT 662.400 527.400 688.050 528.600 ;
        RECT 559.950 522.600 562.050 522.900 ;
        RECT 577.950 522.600 580.050 522.900 ;
        RECT 557.400 521.400 580.050 522.600 ;
        RECT 599.400 521.400 604.050 523.050 ;
        RECT 484.950 520.800 487.050 521.400 ;
        RECT 490.950 520.800 493.050 521.400 ;
        RECT 532.950 520.800 535.050 521.400 ;
        RECT 559.950 520.800 562.050 521.400 ;
        RECT 577.950 520.800 580.050 521.400 ;
        RECT 600.000 520.950 604.050 521.400 ;
        RECT 385.950 518.400 420.600 519.600 ;
        RECT 433.950 519.600 436.050 520.050 ;
        RECT 478.950 519.600 481.050 520.050 ;
        RECT 433.950 518.400 481.050 519.600 ;
        RECT 608.400 519.600 609.600 526.950 ;
        RECT 662.400 525.600 663.600 527.400 ;
        RECT 667.950 527.100 670.050 527.400 ;
        RECT 685.950 527.100 688.050 527.400 ;
        RECT 715.950 528.750 718.050 529.200 ;
        RECT 724.950 528.750 727.050 529.200 ;
        RECT 715.950 527.550 727.050 528.750 ;
        RECT 715.950 527.100 718.050 527.550 ;
        RECT 724.950 527.100 727.050 527.550 ;
        RECT 730.950 528.600 733.050 529.200 ;
        RECT 742.950 528.600 745.050 529.200 ;
        RECT 730.950 527.400 745.050 528.600 ;
        RECT 730.950 527.100 733.050 527.400 ;
        RECT 742.950 527.100 745.050 527.400 ;
        RECT 748.950 526.950 751.050 529.050 ;
        RECT 653.400 524.400 663.600 525.600 ;
        RECT 616.950 522.600 619.050 522.900 ;
        RECT 640.950 522.600 643.050 523.050 ;
        RECT 653.400 522.900 654.600 524.400 ;
        RECT 749.400 523.050 750.600 526.950 ;
        RECT 616.950 521.400 643.050 522.600 ;
        RECT 616.950 520.800 619.050 521.400 ;
        RECT 640.950 520.950 643.050 521.400 ;
        RECT 652.950 520.800 655.050 522.900 ;
        RECT 658.950 522.600 661.050 523.050 ;
        RECT 688.950 522.600 691.050 522.900 ;
        RECT 658.950 521.400 691.050 522.600 ;
        RECT 658.950 520.950 661.050 521.400 ;
        RECT 688.950 520.800 691.050 521.400 ;
        RECT 727.950 522.600 730.050 522.900 ;
        RECT 736.950 522.600 739.050 523.050 ;
        RECT 727.950 521.400 739.050 522.600 ;
        RECT 727.950 520.800 730.050 521.400 ;
        RECT 736.950 520.950 739.050 521.400 ;
        RECT 748.950 520.950 751.050 523.050 ;
        RECT 764.400 522.900 765.600 530.400 ;
        RECT 778.950 528.600 781.050 529.200 ;
        RECT 776.400 527.400 781.050 528.600 ;
        RECT 776.400 523.050 777.600 527.400 ;
        RECT 778.950 527.100 781.050 527.400 ;
        RECT 763.950 520.800 766.050 522.900 ;
        RECT 775.950 520.950 778.050 523.050 ;
        RECT 782.400 522.900 783.600 530.400 ;
        RECT 829.950 530.400 847.050 531.600 ;
        RECT 829.950 529.950 832.050 530.400 ;
        RECT 844.950 529.800 847.050 530.400 ;
        RECT 784.950 527.100 787.050 529.200 ;
        RECT 785.400 523.050 786.600 527.100 ;
        RECT 808.950 525.600 811.050 529.050 ;
        RECT 832.950 526.950 835.050 529.050 ;
        RECT 850.950 528.750 853.050 528.900 ;
        RECT 862.950 528.750 865.050 529.200 ;
        RECT 850.950 527.550 865.050 528.750 ;
        RECT 808.950 525.000 816.600 525.600 ;
        RECT 809.400 524.400 816.600 525.000 ;
        RECT 781.950 520.800 784.050 522.900 ;
        RECT 785.400 521.400 790.050 523.050 ;
        RECT 786.000 520.950 790.050 521.400 ;
        RECT 799.950 522.600 802.050 522.900 ;
        RECT 811.950 522.600 814.050 523.050 ;
        RECT 799.950 521.400 814.050 522.600 ;
        RECT 815.400 522.600 816.600 524.400 ;
        RECT 823.950 522.600 826.050 522.900 ;
        RECT 815.400 521.400 826.050 522.600 ;
        RECT 833.400 522.600 834.600 526.950 ;
        RECT 850.950 526.800 853.050 527.550 ;
        RECT 862.950 527.100 865.050 527.550 ;
        RECT 841.950 522.600 844.050 522.900 ;
        RECT 833.400 521.400 844.050 522.600 ;
        RECT 799.950 520.800 802.050 521.400 ;
        RECT 811.950 520.950 814.050 521.400 ;
        RECT 823.950 520.800 826.050 521.400 ;
        RECT 841.950 520.800 844.050 521.400 ;
        RECT 859.950 522.600 862.050 522.900 ;
        RECT 868.950 522.600 871.050 523.050 ;
        RECT 859.950 521.400 871.050 522.600 ;
        RECT 859.950 520.800 862.050 521.400 ;
        RECT 868.950 520.950 871.050 521.400 ;
        RECT 613.950 519.600 616.050 520.050 ;
        RECT 608.400 518.400 616.050 519.600 ;
        RECT 385.950 517.950 388.050 518.400 ;
        RECT 433.950 517.950 436.050 518.400 ;
        RECT 478.950 517.950 481.050 518.400 ;
        RECT 613.950 517.950 616.050 518.400 ;
        RECT 751.950 519.600 754.050 520.050 ;
        RECT 757.950 519.600 760.050 520.050 ;
        RECT 751.950 518.400 760.050 519.600 ;
        RECT 751.950 517.950 754.050 518.400 ;
        RECT 757.950 517.950 760.050 518.400 ;
        RECT 112.950 516.600 115.050 517.050 ;
        RECT 118.950 516.600 121.050 517.050 ;
        RECT 112.950 515.400 121.050 516.600 ;
        RECT 112.950 514.950 115.050 515.400 ;
        RECT 118.950 514.950 121.050 515.400 ;
        RECT 136.950 516.600 139.050 517.050 ;
        RECT 157.950 516.600 160.050 517.050 ;
        RECT 136.950 515.400 160.050 516.600 ;
        RECT 136.950 514.950 139.050 515.400 ;
        RECT 157.950 514.950 160.050 515.400 ;
        RECT 181.950 516.600 184.050 517.050 ;
        RECT 409.950 516.600 412.050 517.050 ;
        RECT 181.950 515.400 412.050 516.600 ;
        RECT 181.950 514.950 184.050 515.400 ;
        RECT 409.950 514.950 412.050 515.400 ;
        RECT 577.950 516.600 580.050 517.050 ;
        RECT 589.950 516.600 592.050 517.050 ;
        RECT 577.950 515.400 592.050 516.600 ;
        RECT 577.950 514.950 580.050 515.400 ;
        RECT 589.950 514.950 592.050 515.400 ;
        RECT 643.950 516.600 646.050 517.050 ;
        RECT 670.950 516.600 673.050 517.050 ;
        RECT 643.950 515.400 673.050 516.600 ;
        RECT 643.950 514.950 646.050 515.400 ;
        RECT 670.950 514.950 673.050 515.400 ;
        RECT 715.950 516.600 718.050 517.050 ;
        RECT 727.950 516.600 730.050 517.050 ;
        RECT 715.950 515.400 730.050 516.600 ;
        RECT 715.950 514.950 718.050 515.400 ;
        RECT 727.950 514.950 730.050 515.400 ;
        RECT 745.950 516.600 748.050 517.050 ;
        RECT 787.950 516.600 790.050 517.050 ;
        RECT 820.950 516.600 823.050 517.050 ;
        RECT 835.950 516.600 838.050 517.050 ;
        RECT 745.950 515.400 838.050 516.600 ;
        RECT 745.950 514.950 748.050 515.400 ;
        RECT 787.950 514.950 790.050 515.400 ;
        RECT 820.950 514.950 823.050 515.400 ;
        RECT 835.950 514.950 838.050 515.400 ;
        RECT 289.950 513.600 292.050 514.050 ;
        RECT 307.950 513.600 310.050 514.050 ;
        RECT 289.950 512.400 310.050 513.600 ;
        RECT 289.950 511.950 292.050 512.400 ;
        RECT 307.950 511.950 310.050 512.400 ;
        RECT 346.950 513.600 349.050 514.050 ;
        RECT 391.950 513.600 394.050 514.050 ;
        RECT 346.950 512.400 394.050 513.600 ;
        RECT 346.950 511.950 349.050 512.400 ;
        RECT 391.950 511.950 394.050 512.400 ;
        RECT 415.950 513.600 418.050 514.050 ;
        RECT 484.950 513.600 487.050 514.050 ;
        RECT 415.950 512.400 487.050 513.600 ;
        RECT 415.950 511.950 418.050 512.400 ;
        RECT 484.950 511.950 487.050 512.400 ;
        RECT 532.950 513.600 535.050 514.050 ;
        RECT 547.950 513.600 550.050 514.050 ;
        RECT 532.950 512.400 550.050 513.600 ;
        RECT 532.950 511.950 535.050 512.400 ;
        RECT 547.950 511.950 550.050 512.400 ;
        RECT 556.950 513.600 559.050 514.050 ;
        RECT 610.950 513.600 613.050 514.050 ;
        RECT 556.950 512.400 613.050 513.600 ;
        RECT 556.950 511.950 559.050 512.400 ;
        RECT 610.950 511.950 613.050 512.400 ;
        RECT 706.950 513.600 709.050 514.050 ;
        RECT 721.950 513.600 724.050 514.050 ;
        RECT 706.950 512.400 724.050 513.600 ;
        RECT 706.950 511.950 709.050 512.400 ;
        RECT 721.950 511.950 724.050 512.400 ;
        RECT 778.950 513.600 781.050 514.050 ;
        RECT 790.950 513.600 793.050 514.050 ;
        RECT 778.950 512.400 793.050 513.600 ;
        RECT 778.950 511.950 781.050 512.400 ;
        RECT 790.950 511.950 793.050 512.400 ;
        RECT 25.950 510.600 28.050 511.050 ;
        RECT 52.950 510.600 55.050 511.050 ;
        RECT 25.950 509.400 55.050 510.600 ;
        RECT 25.950 508.950 28.050 509.400 ;
        RECT 52.950 508.950 55.050 509.400 ;
        RECT 130.950 510.600 133.050 511.050 ;
        RECT 208.950 510.600 211.050 511.050 ;
        RECT 130.950 509.400 211.050 510.600 ;
        RECT 130.950 508.950 133.050 509.400 ;
        RECT 208.950 508.950 211.050 509.400 ;
        RECT 226.950 510.600 229.050 511.050 ;
        RECT 232.950 510.600 235.050 511.050 ;
        RECT 226.950 509.400 235.050 510.600 ;
        RECT 226.950 508.950 229.050 509.400 ;
        RECT 232.950 508.950 235.050 509.400 ;
        RECT 265.950 510.600 268.050 511.050 ;
        RECT 271.950 510.600 274.050 511.050 ;
        RECT 265.950 509.400 274.050 510.600 ;
        RECT 265.950 508.950 268.050 509.400 ;
        RECT 271.950 508.950 274.050 509.400 ;
        RECT 310.950 510.600 313.050 511.050 ;
        RECT 373.950 510.600 376.050 511.050 ;
        RECT 310.950 509.400 376.050 510.600 ;
        RECT 310.950 508.950 313.050 509.400 ;
        RECT 373.950 508.950 376.050 509.400 ;
        RECT 445.950 510.600 448.050 511.050 ;
        RECT 457.950 510.600 460.050 511.050 ;
        RECT 445.950 509.400 460.050 510.600 ;
        RECT 445.950 508.950 448.050 509.400 ;
        RECT 457.950 508.950 460.050 509.400 ;
        RECT 472.950 510.600 475.050 511.050 ;
        RECT 484.950 510.600 487.050 510.900 ;
        RECT 562.950 510.600 565.050 511.050 ;
        RECT 571.950 510.600 574.050 511.050 ;
        RECT 472.950 509.400 487.050 510.600 ;
        RECT 472.950 508.950 475.050 509.400 ;
        RECT 484.950 508.800 487.050 509.400 ;
        RECT 536.400 509.400 574.050 510.600 ;
        RECT 70.950 507.600 73.050 508.050 ;
        RECT 106.950 507.600 109.050 508.050 ;
        RECT 70.950 506.400 109.050 507.600 ;
        RECT 70.950 505.950 73.050 506.400 ;
        RECT 106.950 505.950 109.050 506.400 ;
        RECT 127.950 507.600 130.050 508.050 ;
        RECT 181.950 507.600 184.050 508.050 ;
        RECT 127.950 506.400 184.050 507.600 ;
        RECT 127.950 505.950 130.050 506.400 ;
        RECT 181.950 505.950 184.050 506.400 ;
        RECT 256.950 507.600 259.050 508.050 ;
        RECT 268.950 507.600 271.050 508.050 ;
        RECT 256.950 506.400 271.050 507.600 ;
        RECT 256.950 505.950 259.050 506.400 ;
        RECT 268.950 505.950 271.050 506.400 ;
        RECT 277.950 507.600 280.050 508.050 ;
        RECT 295.950 507.600 298.050 508.050 ;
        RECT 277.950 506.400 298.050 507.600 ;
        RECT 277.950 505.950 280.050 506.400 ;
        RECT 295.950 505.950 298.050 506.400 ;
        RECT 400.950 507.600 403.050 508.050 ;
        RECT 536.400 507.600 537.600 509.400 ;
        RECT 562.950 508.950 565.050 509.400 ;
        RECT 571.950 508.950 574.050 509.400 ;
        RECT 583.950 510.600 586.050 511.050 ;
        RECT 643.950 510.600 646.050 511.050 ;
        RECT 583.950 509.400 646.050 510.600 ;
        RECT 583.950 508.950 586.050 509.400 ;
        RECT 643.950 508.950 646.050 509.400 ;
        RECT 691.950 510.600 694.050 511.050 ;
        RECT 733.950 510.600 736.050 511.050 ;
        RECT 691.950 509.400 736.050 510.600 ;
        RECT 691.950 508.950 694.050 509.400 ;
        RECT 733.950 508.950 736.050 509.400 ;
        RECT 802.950 510.600 805.050 511.050 ;
        RECT 847.950 510.600 850.050 511.050 ;
        RECT 802.950 509.400 850.050 510.600 ;
        RECT 802.950 508.950 805.050 509.400 ;
        RECT 847.950 508.950 850.050 509.400 ;
        RECT 400.950 506.400 537.600 507.600 ;
        RECT 712.950 507.600 715.050 508.050 ;
        RECT 721.950 507.600 724.050 508.050 ;
        RECT 712.950 506.400 724.050 507.600 ;
        RECT 400.950 505.950 403.050 506.400 ;
        RECT 712.950 505.950 715.050 506.400 ;
        RECT 721.950 505.950 724.050 506.400 ;
        RECT 13.950 504.600 16.050 505.050 ;
        RECT 28.950 504.600 31.050 505.050 ;
        RECT 13.950 503.400 31.050 504.600 ;
        RECT 13.950 502.950 16.050 503.400 ;
        RECT 28.950 502.950 31.050 503.400 ;
        RECT 88.950 504.600 91.050 505.050 ;
        RECT 142.950 504.600 145.050 505.050 ;
        RECT 283.950 504.600 286.050 505.050 ;
        RECT 88.950 503.400 286.050 504.600 ;
        RECT 88.950 502.950 91.050 503.400 ;
        RECT 142.950 502.950 145.050 503.400 ;
        RECT 283.950 502.950 286.050 503.400 ;
        RECT 301.950 504.600 304.050 505.050 ;
        RECT 316.950 504.600 319.050 505.050 ;
        RECT 301.950 503.400 319.050 504.600 ;
        RECT 301.950 502.950 304.050 503.400 ;
        RECT 316.950 502.950 319.050 503.400 ;
        RECT 493.950 504.600 496.050 505.050 ;
        RECT 538.950 504.600 541.050 505.050 ;
        RECT 565.950 504.600 568.050 505.050 ;
        RECT 493.950 503.400 568.050 504.600 ;
        RECT 493.950 502.950 496.050 503.400 ;
        RECT 538.950 502.950 541.050 503.400 ;
        RECT 565.950 502.950 568.050 503.400 ;
        RECT 790.950 504.600 793.050 505.050 ;
        RECT 823.950 504.600 826.050 505.050 ;
        RECT 790.950 503.400 826.050 504.600 ;
        RECT 790.950 502.950 793.050 503.400 ;
        RECT 823.950 502.950 826.050 503.400 ;
        RECT 853.950 504.600 856.050 505.050 ;
        RECT 859.950 504.600 862.050 505.050 ;
        RECT 853.950 503.400 862.050 504.600 ;
        RECT 853.950 502.950 856.050 503.400 ;
        RECT 859.950 502.950 862.050 503.400 ;
        RECT 145.950 501.600 148.050 502.050 ;
        RECT 193.950 501.600 196.050 502.050 ;
        RECT 145.950 500.400 196.050 501.600 ;
        RECT 145.950 499.950 148.050 500.400 ;
        RECT 193.950 499.950 196.050 500.400 ;
        RECT 244.950 501.600 247.050 502.050 ;
        RECT 259.950 501.600 262.050 502.050 ;
        RECT 244.950 500.400 262.050 501.600 ;
        RECT 244.950 499.950 247.050 500.400 ;
        RECT 259.950 499.950 262.050 500.400 ;
        RECT 406.950 501.600 409.050 502.050 ;
        RECT 439.950 501.600 442.050 502.050 ;
        RECT 406.950 500.400 442.050 501.600 ;
        RECT 406.950 499.950 409.050 500.400 ;
        RECT 439.950 499.950 442.050 500.400 ;
        RECT 523.950 501.600 526.050 502.050 ;
        RECT 535.950 501.600 538.050 502.050 ;
        RECT 556.950 501.600 559.050 502.050 ;
        RECT 523.950 500.400 559.050 501.600 ;
        RECT 523.950 499.950 526.050 500.400 ;
        RECT 535.950 499.950 538.050 500.400 ;
        RECT 556.950 499.950 559.050 500.400 ;
        RECT 628.950 501.600 631.050 502.050 ;
        RECT 661.950 501.600 664.050 502.050 ;
        RECT 628.950 500.400 664.050 501.600 ;
        RECT 628.950 499.950 631.050 500.400 ;
        RECT 661.950 499.950 664.050 500.400 ;
        RECT 700.950 501.600 703.050 502.050 ;
        RECT 784.950 501.600 787.050 502.050 ;
        RECT 700.950 500.400 787.050 501.600 ;
        RECT 700.950 499.950 703.050 500.400 ;
        RECT 784.950 499.950 787.050 500.400 ;
        RECT 10.950 498.600 15.000 499.050 ;
        RECT 373.950 498.600 376.050 499.050 ;
        RECT 382.950 498.600 385.050 499.050 ;
        RECT 409.950 498.600 412.050 499.050 ;
        RECT 10.950 496.950 15.600 498.600 ;
        RECT 373.950 497.400 412.050 498.600 ;
        RECT 373.950 496.950 376.050 497.400 ;
        RECT 382.950 496.950 385.050 497.400 ;
        RECT 409.950 496.950 412.050 497.400 ;
        RECT 502.950 498.600 505.050 499.050 ;
        RECT 508.950 498.600 511.050 499.050 ;
        RECT 502.950 497.400 511.050 498.600 ;
        RECT 502.950 496.950 505.050 497.400 ;
        RECT 508.950 496.950 511.050 497.400 ;
        RECT 730.950 498.600 733.050 499.050 ;
        RECT 739.950 498.600 742.050 499.050 ;
        RECT 730.950 497.400 742.050 498.600 ;
        RECT 730.950 496.950 733.050 497.400 ;
        RECT 739.950 496.950 742.050 497.400 ;
        RECT 775.950 496.950 778.050 499.050 ;
        RECT 7.950 493.950 10.050 496.050 ;
        RECT 8.400 490.050 9.600 493.950 ;
        RECT 7.950 487.950 10.050 490.050 ;
        RECT 14.400 487.050 15.600 496.950 ;
        RECT 31.950 494.100 34.050 496.200 ;
        RECT 46.950 495.600 49.050 496.050 ;
        RECT 55.950 495.600 58.050 496.200 ;
        RECT 46.950 494.400 58.050 495.600 ;
        RECT 32.400 492.600 33.600 494.100 ;
        RECT 46.950 493.950 49.050 494.400 ;
        RECT 55.950 494.100 58.050 494.400 ;
        RECT 64.950 495.750 67.050 496.200 ;
        RECT 70.950 495.750 73.050 496.200 ;
        RECT 64.950 494.550 73.050 495.750 ;
        RECT 88.950 495.600 91.050 496.050 ;
        RECT 64.950 494.100 67.050 494.550 ;
        RECT 70.950 494.100 73.050 494.550 ;
        RECT 74.400 494.400 91.050 495.600 ;
        RECT 32.400 491.400 39.600 492.600 ;
        RECT 22.950 489.450 25.050 489.900 ;
        RECT 34.950 489.450 37.050 489.900 ;
        RECT 22.950 488.250 37.050 489.450 ;
        RECT 38.400 489.600 39.600 491.400 ;
        RECT 74.400 489.900 75.600 494.400 ;
        RECT 88.950 493.950 91.050 494.400 ;
        RECT 100.950 495.750 103.050 496.200 ;
        RECT 112.950 495.750 115.050 496.200 ;
        RECT 100.950 494.550 115.050 495.750 ;
        RECT 100.950 494.100 103.050 494.550 ;
        RECT 112.950 494.100 115.050 494.550 ;
        RECT 157.950 495.750 160.050 496.200 ;
        RECT 163.950 495.750 166.050 496.200 ;
        RECT 157.950 495.600 166.050 495.750 ;
        RECT 175.950 495.600 178.050 496.200 ;
        RECT 157.950 494.550 178.050 495.600 ;
        RECT 157.950 494.100 160.050 494.550 ;
        RECT 163.950 494.400 178.050 494.550 ;
        RECT 163.950 494.100 166.050 494.400 ;
        RECT 175.950 494.100 178.050 494.400 ;
        RECT 199.950 495.600 202.050 496.200 ;
        RECT 274.950 495.600 277.050 496.050 ;
        RECT 280.950 495.600 283.050 496.200 ;
        RECT 199.950 494.400 219.600 495.600 ;
        RECT 199.950 494.100 202.050 494.400 ;
        RECT 184.950 492.600 187.050 493.050 ;
        RECT 184.950 491.400 210.600 492.600 ;
        RECT 184.950 490.950 187.050 491.400 ;
        RECT 52.950 489.600 55.050 489.900 ;
        RECT 38.400 488.400 55.050 489.600 ;
        RECT 22.950 487.800 25.050 488.250 ;
        RECT 34.950 487.800 37.050 488.250 ;
        RECT 52.950 487.800 55.050 488.400 ;
        RECT 73.950 487.800 76.050 489.900 ;
        RECT 79.950 489.600 82.050 489.900 ;
        RECT 91.950 489.600 94.050 489.900 ;
        RECT 79.950 488.400 94.050 489.600 ;
        RECT 79.950 487.800 82.050 488.400 ;
        RECT 91.950 487.800 94.050 488.400 ;
        RECT 145.950 489.600 148.050 490.050 ;
        RECT 209.400 489.900 210.600 491.400 ;
        RECT 218.400 489.900 219.600 494.400 ;
        RECT 274.950 494.400 283.050 495.600 ;
        RECT 274.950 493.950 277.050 494.400 ;
        RECT 280.950 494.100 283.050 494.400 ;
        RECT 301.950 494.100 304.050 496.200 ;
        RECT 418.950 495.600 421.050 496.200 ;
        RECT 424.950 495.750 427.050 496.200 ;
        RECT 430.950 495.750 433.050 496.200 ;
        RECT 418.950 494.400 423.600 495.600 ;
        RECT 418.950 494.100 421.050 494.400 ;
        RECT 154.950 489.600 157.050 489.900 ;
        RECT 196.950 489.600 199.050 489.900 ;
        RECT 145.950 488.400 157.050 489.600 ;
        RECT 145.950 487.950 148.050 488.400 ;
        RECT 154.950 487.800 157.050 488.400 ;
        RECT 194.400 488.400 199.050 489.600 ;
        RECT 10.950 485.400 15.600 487.050 ;
        RECT 109.950 486.600 112.050 487.050 ;
        RECT 121.950 486.600 124.050 487.050 ;
        RECT 109.950 485.400 124.050 486.600 ;
        RECT 10.950 484.950 15.000 485.400 ;
        RECT 109.950 484.950 112.050 485.400 ;
        RECT 121.950 484.950 124.050 485.400 ;
        RECT 172.950 486.600 175.050 487.050 ;
        RECT 194.400 486.600 195.600 488.400 ;
        RECT 196.950 487.800 199.050 488.400 ;
        RECT 208.950 487.800 211.050 489.900 ;
        RECT 217.950 487.800 220.050 489.900 ;
        RECT 241.950 489.450 244.050 489.900 ;
        RECT 250.950 489.450 253.050 489.900 ;
        RECT 241.950 488.250 253.050 489.450 ;
        RECT 241.950 487.800 244.050 488.250 ;
        RECT 250.950 487.800 253.050 488.250 ;
        RECT 295.950 489.600 298.050 489.900 ;
        RECT 302.400 489.600 303.600 494.100 ;
        RECT 337.950 492.600 340.050 493.050 ;
        RECT 406.950 492.600 409.050 493.050 ;
        RECT 326.400 491.400 340.050 492.600 ;
        RECT 295.950 488.400 303.600 489.600 ;
        RECT 319.950 489.600 322.050 489.900 ;
        RECT 326.400 489.600 327.600 491.400 ;
        RECT 337.950 490.950 340.050 491.400 ;
        RECT 392.400 491.400 409.050 492.600 ;
        RECT 422.400 492.600 423.600 494.400 ;
        RECT 424.950 494.550 433.050 495.750 ;
        RECT 424.950 494.100 427.050 494.550 ;
        RECT 430.950 494.100 433.050 494.550 ;
        RECT 451.950 495.750 454.050 496.200 ;
        RECT 460.950 495.750 463.050 496.200 ;
        RECT 451.950 494.550 463.050 495.750 ;
        RECT 499.950 495.600 502.050 496.200 ;
        RECT 517.950 495.600 520.050 496.200 ;
        RECT 451.950 494.100 454.050 494.550 ;
        RECT 460.950 494.100 463.050 494.550 ;
        RECT 488.400 494.400 502.050 495.600 ;
        RECT 488.400 492.600 489.600 494.400 ;
        RECT 499.950 494.100 502.050 494.400 ;
        RECT 506.400 494.400 520.050 495.600 ;
        RECT 506.400 492.600 507.600 494.400 ;
        RECT 517.950 494.100 520.050 494.400 ;
        RECT 523.950 495.750 526.050 496.200 ;
        RECT 544.950 495.750 547.050 496.200 ;
        RECT 523.950 495.600 547.050 495.750 ;
        RECT 559.950 495.600 562.050 496.050 ;
        RECT 601.950 495.600 604.050 496.050 ;
        RECT 523.950 494.550 604.050 495.600 ;
        RECT 523.950 494.100 526.050 494.550 ;
        RECT 544.950 494.400 604.050 494.550 ;
        RECT 544.950 494.100 547.050 494.400 ;
        RECT 559.950 493.950 562.050 494.400 ;
        RECT 601.950 493.950 604.050 494.400 ;
        RECT 649.950 495.750 652.050 496.200 ;
        RECT 655.950 495.750 658.050 496.200 ;
        RECT 649.950 494.550 658.050 495.750 ;
        RECT 649.950 494.100 652.050 494.550 ;
        RECT 655.950 494.100 658.050 494.550 ;
        RECT 664.950 494.100 667.050 496.200 ;
        RECT 670.950 495.600 673.050 496.200 ;
        RECT 676.950 495.600 679.050 496.050 ;
        RECT 670.950 494.400 679.050 495.600 ;
        RECT 670.950 494.100 673.050 494.400 ;
        RECT 422.400 491.400 435.600 492.600 ;
        RECT 392.400 489.900 393.600 491.400 ;
        RECT 406.950 490.950 409.050 491.400 ;
        RECT 319.950 488.400 327.600 489.600 ;
        RECT 295.950 487.800 298.050 488.400 ;
        RECT 319.950 487.800 322.050 488.400 ;
        RECT 391.950 487.800 394.050 489.900 ;
        RECT 409.950 489.600 412.050 490.050 ;
        RECT 415.950 489.600 418.050 489.900 ;
        RECT 409.950 488.400 418.050 489.600 ;
        RECT 434.400 489.600 435.600 491.400 ;
        RECT 470.400 491.400 489.600 492.600 ;
        RECT 503.400 491.400 507.600 492.600 ;
        RECT 470.400 489.900 471.600 491.400 ;
        RECT 503.400 489.900 504.600 491.400 ;
        RECT 436.950 489.600 439.050 489.900 ;
        RECT 434.400 488.400 439.050 489.600 ;
        RECT 409.950 487.950 412.050 488.400 ;
        RECT 415.950 487.800 418.050 488.400 ;
        RECT 436.950 487.800 439.050 488.400 ;
        RECT 469.950 487.800 472.050 489.900 ;
        RECT 502.950 487.800 505.050 489.900 ;
        RECT 577.950 489.450 580.050 489.900 ;
        RECT 583.950 489.450 586.050 489.900 ;
        RECT 577.950 488.250 586.050 489.450 ;
        RECT 577.950 487.800 580.050 488.250 ;
        RECT 583.950 487.800 586.050 488.250 ;
        RECT 592.950 489.450 595.050 489.900 ;
        RECT 628.950 489.450 631.050 489.900 ;
        RECT 592.950 488.250 631.050 489.450 ;
        RECT 592.950 487.800 595.050 488.250 ;
        RECT 628.950 487.800 631.050 488.250 ;
        RECT 665.400 487.050 666.600 494.100 ;
        RECT 676.950 493.950 679.050 494.400 ;
        RECT 685.950 495.750 688.050 496.200 ;
        RECT 691.950 495.750 694.050 496.200 ;
        RECT 685.950 494.550 694.050 495.750 ;
        RECT 685.950 494.100 688.050 494.550 ;
        RECT 691.950 494.100 694.050 494.550 ;
        RECT 700.950 495.600 703.050 496.200 ;
        RECT 748.950 495.750 751.050 496.200 ;
        RECT 760.950 495.750 763.050 496.200 ;
        RECT 700.950 494.400 738.600 495.600 ;
        RECT 700.950 494.100 703.050 494.400 ;
        RECT 667.950 489.600 670.050 489.900 ;
        RECT 682.950 489.600 685.050 489.900 ;
        RECT 706.950 489.600 709.050 490.050 ;
        RECT 737.400 489.900 738.600 494.400 ;
        RECT 748.950 494.550 763.050 495.750 ;
        RECT 748.950 494.100 751.050 494.550 ;
        RECT 760.950 494.100 763.050 494.550 ;
        RECT 667.950 488.400 709.050 489.600 ;
        RECT 667.950 487.800 670.050 488.400 ;
        RECT 682.950 487.800 685.050 488.400 ;
        RECT 706.950 487.950 709.050 488.400 ;
        RECT 718.950 489.450 721.050 489.900 ;
        RECT 724.950 489.450 727.050 489.900 ;
        RECT 718.950 488.250 727.050 489.450 ;
        RECT 718.950 487.800 721.050 488.250 ;
        RECT 724.950 487.800 727.050 488.250 ;
        RECT 736.950 487.800 739.050 489.900 ;
        RECT 754.950 489.450 757.050 489.900 ;
        RECT 766.950 489.450 769.050 489.900 ;
        RECT 754.950 488.250 769.050 489.450 ;
        RECT 776.400 489.600 777.600 496.950 ;
        RECT 784.950 495.600 787.050 496.200 ;
        RECT 796.950 495.600 799.050 496.200 ;
        RECT 784.950 494.400 799.050 495.600 ;
        RECT 784.950 494.100 787.050 494.400 ;
        RECT 796.950 494.100 799.050 494.400 ;
        RECT 832.950 495.750 835.050 496.200 ;
        RECT 853.950 495.750 856.050 496.200 ;
        RECT 832.950 494.550 856.050 495.750 ;
        RECT 832.950 494.100 835.050 494.550 ;
        RECT 853.950 494.100 856.050 494.550 ;
        RECT 781.950 489.600 784.050 489.900 ;
        RECT 776.400 488.400 784.050 489.600 ;
        RECT 754.950 487.800 757.050 488.250 ;
        RECT 766.950 487.800 769.050 488.250 ;
        RECT 781.950 487.800 784.050 488.400 ;
        RECT 808.950 489.450 811.050 489.900 ;
        RECT 838.950 489.450 841.050 489.900 ;
        RECT 808.950 488.250 841.050 489.450 ;
        RECT 808.950 487.800 811.050 488.250 ;
        RECT 838.950 487.800 841.050 488.250 ;
        RECT 172.950 485.400 195.600 486.600 ;
        RECT 328.950 486.600 331.050 487.050 ;
        RECT 364.950 486.600 367.050 487.050 ;
        RECT 385.950 486.600 388.050 487.050 ;
        RECT 400.950 486.600 403.050 487.050 ;
        RECT 328.950 485.400 403.050 486.600 ;
        RECT 172.950 484.950 175.050 485.400 ;
        RECT 328.950 484.950 331.050 485.400 ;
        RECT 364.950 484.950 367.050 485.400 ;
        RECT 385.950 484.950 388.050 485.400 ;
        RECT 400.950 484.950 403.050 485.400 ;
        RECT 664.950 484.950 667.050 487.050 ;
        RECT 697.950 486.600 700.050 487.050 ;
        RECT 703.950 486.600 706.050 487.050 ;
        RECT 697.950 485.400 706.050 486.600 ;
        RECT 697.950 484.950 700.050 485.400 ;
        RECT 703.950 484.950 706.050 485.400 ;
        RECT 742.950 486.600 745.050 487.050 ;
        RECT 772.950 486.600 775.050 487.050 ;
        RECT 742.950 485.400 775.050 486.600 ;
        RECT 742.950 484.950 745.050 485.400 ;
        RECT 772.950 484.950 775.050 485.400 ;
        RECT 181.950 483.600 184.050 484.050 ;
        RECT 268.950 483.600 271.050 484.050 ;
        RECT 181.950 482.400 271.050 483.600 ;
        RECT 181.950 481.950 184.050 482.400 ;
        RECT 268.950 481.950 271.050 482.400 ;
        RECT 460.950 483.600 463.050 484.050 ;
        RECT 514.950 483.600 517.050 484.050 ;
        RECT 460.950 482.400 517.050 483.600 ;
        RECT 460.950 481.950 463.050 482.400 ;
        RECT 514.950 481.950 517.050 482.400 ;
        RECT 580.950 483.600 583.050 484.050 ;
        RECT 712.950 483.600 715.050 484.050 ;
        RECT 727.950 483.600 730.050 484.050 ;
        RECT 580.950 482.400 730.050 483.600 ;
        RECT 580.950 481.950 583.050 482.400 ;
        RECT 712.950 481.950 715.050 482.400 ;
        RECT 727.950 481.950 730.050 482.400 ;
        RECT 787.950 483.600 790.050 484.050 ;
        RECT 811.950 483.600 814.050 484.050 ;
        RECT 787.950 482.400 814.050 483.600 ;
        RECT 787.950 481.950 790.050 482.400 ;
        RECT 811.950 481.950 814.050 482.400 ;
        RECT 817.950 483.600 820.050 484.050 ;
        RECT 835.950 483.600 838.050 484.050 ;
        RECT 817.950 482.400 838.050 483.600 ;
        RECT 817.950 481.950 820.050 482.400 ;
        RECT 835.950 481.950 838.050 482.400 ;
        RECT 19.950 480.600 22.050 481.050 ;
        RECT 52.950 480.600 55.050 481.050 ;
        RECT 118.950 480.600 121.050 481.050 ;
        RECT 127.950 480.600 130.050 481.050 ;
        RECT 19.950 479.400 130.050 480.600 ;
        RECT 19.950 478.950 22.050 479.400 ;
        RECT 52.950 478.950 55.050 479.400 ;
        RECT 118.950 478.950 121.050 479.400 ;
        RECT 127.950 478.950 130.050 479.400 ;
        RECT 148.950 480.600 151.050 481.050 ;
        RECT 163.950 480.600 166.050 481.050 ;
        RECT 148.950 479.400 166.050 480.600 ;
        RECT 148.950 478.950 151.050 479.400 ;
        RECT 163.950 478.950 166.050 479.400 ;
        RECT 187.950 480.600 190.050 481.050 ;
        RECT 193.950 480.600 196.050 481.050 ;
        RECT 187.950 479.400 196.050 480.600 ;
        RECT 187.950 478.950 190.050 479.400 ;
        RECT 193.950 478.950 196.050 479.400 ;
        RECT 202.950 480.600 205.050 481.050 ;
        RECT 226.950 480.600 229.050 481.050 ;
        RECT 202.950 479.400 229.050 480.600 ;
        RECT 202.950 478.950 205.050 479.400 ;
        RECT 226.950 478.950 229.050 479.400 ;
        RECT 493.950 480.600 496.050 481.050 ;
        RECT 538.950 480.600 541.050 481.050 ;
        RECT 493.950 479.400 541.050 480.600 ;
        RECT 493.950 478.950 496.050 479.400 ;
        RECT 538.950 478.950 541.050 479.400 ;
        RECT 676.950 480.600 679.050 481.050 ;
        RECT 781.950 480.600 784.050 481.050 ;
        RECT 676.950 479.400 784.050 480.600 ;
        RECT 676.950 478.950 679.050 479.400 ;
        RECT 781.950 478.950 784.050 479.400 ;
        RECT 154.950 477.600 157.050 478.050 ;
        RECT 181.950 477.600 184.050 478.050 ;
        RECT 154.950 476.400 184.050 477.600 ;
        RECT 154.950 475.950 157.050 476.400 ;
        RECT 181.950 475.950 184.050 476.400 ;
        RECT 235.950 477.600 238.050 478.050 ;
        RECT 328.950 477.600 331.050 478.050 ;
        RECT 235.950 476.400 331.050 477.600 ;
        RECT 235.950 475.950 238.050 476.400 ;
        RECT 328.950 475.950 331.050 476.400 ;
        RECT 514.950 477.600 517.050 478.050 ;
        RECT 532.950 477.600 535.050 478.050 ;
        RECT 514.950 476.400 535.050 477.600 ;
        RECT 514.950 475.950 517.050 476.400 ;
        RECT 532.950 475.950 535.050 476.400 ;
        RECT 58.950 474.600 61.050 475.050 ;
        RECT 460.950 474.600 463.050 475.050 ;
        RECT 58.950 473.400 463.050 474.600 ;
        RECT 58.950 472.950 61.050 473.400 ;
        RECT 460.950 472.950 463.050 473.400 ;
        RECT 538.950 474.600 541.050 475.050 ;
        RECT 631.950 474.600 634.050 475.050 ;
        RECT 661.950 474.600 664.050 475.050 ;
        RECT 538.950 473.400 664.050 474.600 ;
        RECT 538.950 472.950 541.050 473.400 ;
        RECT 631.950 472.950 634.050 473.400 ;
        RECT 661.950 472.950 664.050 473.400 ;
        RECT 763.950 474.600 766.050 475.050 ;
        RECT 790.950 474.600 793.050 475.050 ;
        RECT 763.950 473.400 793.050 474.600 ;
        RECT 763.950 472.950 766.050 473.400 ;
        RECT 790.950 472.950 793.050 473.400 ;
        RECT 304.950 471.600 307.050 472.050 ;
        RECT 310.950 471.600 313.050 472.050 ;
        RECT 304.950 470.400 313.050 471.600 ;
        RECT 304.950 469.950 307.050 470.400 ;
        RECT 310.950 469.950 313.050 470.400 ;
        RECT 55.950 468.600 58.050 469.050 ;
        RECT 64.950 468.600 67.050 469.050 ;
        RECT 55.950 467.400 67.050 468.600 ;
        RECT 55.950 466.950 58.050 467.400 ;
        RECT 64.950 466.950 67.050 467.400 ;
        RECT 199.950 468.600 202.050 469.050 ;
        RECT 253.950 468.600 256.050 469.050 ;
        RECT 199.950 467.400 256.050 468.600 ;
        RECT 199.950 466.950 202.050 467.400 ;
        RECT 253.950 466.950 256.050 467.400 ;
        RECT 346.950 468.600 349.050 469.050 ;
        RECT 496.950 468.600 499.050 469.050 ;
        RECT 346.950 467.400 499.050 468.600 ;
        RECT 346.950 466.950 349.050 467.400 ;
        RECT 496.950 466.950 499.050 467.400 ;
        RECT 520.950 468.600 523.050 469.050 ;
        RECT 553.950 468.600 556.050 469.050 ;
        RECT 520.950 467.400 556.050 468.600 ;
        RECT 520.950 466.950 523.050 467.400 ;
        RECT 553.950 466.950 556.050 467.400 ;
        RECT 616.950 468.600 619.050 469.050 ;
        RECT 625.950 468.600 628.050 469.050 ;
        RECT 616.950 467.400 628.050 468.600 ;
        RECT 616.950 466.950 619.050 467.400 ;
        RECT 625.950 466.950 628.050 467.400 ;
        RECT 118.950 465.600 121.050 466.050 ;
        RECT 223.950 465.600 226.050 466.050 ;
        RECT 118.950 464.400 226.050 465.600 ;
        RECT 118.950 463.950 121.050 464.400 ;
        RECT 223.950 463.950 226.050 464.400 ;
        RECT 160.950 462.600 163.050 463.050 ;
        RECT 244.950 462.600 247.050 463.050 ;
        RECT 334.950 462.600 337.050 463.050 ;
        RECT 160.950 461.400 337.050 462.600 ;
        RECT 160.950 460.950 163.050 461.400 ;
        RECT 244.950 460.950 247.050 461.400 ;
        RECT 334.950 460.950 337.050 461.400 ;
        RECT 400.950 462.600 403.050 463.050 ;
        RECT 421.950 462.600 424.050 463.050 ;
        RECT 460.950 462.600 463.050 463.050 ;
        RECT 520.950 462.600 523.050 463.050 ;
        RECT 400.950 461.400 523.050 462.600 ;
        RECT 400.950 460.950 403.050 461.400 ;
        RECT 421.950 460.950 424.050 461.400 ;
        RECT 460.950 460.950 463.050 461.400 ;
        RECT 520.950 460.950 523.050 461.400 ;
        RECT 589.950 462.600 592.050 463.050 ;
        RECT 604.950 462.600 607.050 463.050 ;
        RECT 679.950 462.600 682.050 463.050 ;
        RECT 589.950 461.400 682.050 462.600 ;
        RECT 589.950 460.950 592.050 461.400 ;
        RECT 604.950 460.950 607.050 461.400 ;
        RECT 679.950 460.950 682.050 461.400 ;
        RECT 700.950 462.600 703.050 463.050 ;
        RECT 742.950 462.600 745.050 463.050 ;
        RECT 700.950 461.400 745.050 462.600 ;
        RECT 700.950 460.950 703.050 461.400 ;
        RECT 742.950 460.950 745.050 461.400 ;
        RECT 853.950 462.600 856.050 463.050 ;
        RECT 871.950 462.600 874.050 463.050 ;
        RECT 853.950 461.400 874.050 462.600 ;
        RECT 853.950 460.950 856.050 461.400 ;
        RECT 871.950 460.950 874.050 461.400 ;
        RECT 73.950 459.600 76.050 460.050 ;
        RECT 85.950 459.600 88.050 460.050 ;
        RECT 73.950 458.400 88.050 459.600 ;
        RECT 73.950 457.950 76.050 458.400 ;
        RECT 85.950 457.950 88.050 458.400 ;
        RECT 166.950 459.600 169.050 460.050 ;
        RECT 190.950 459.600 193.050 460.050 ;
        RECT 166.950 458.400 193.050 459.600 ;
        RECT 166.950 457.950 169.050 458.400 ;
        RECT 190.950 457.950 193.050 458.400 ;
        RECT 271.950 459.600 274.050 460.050 ;
        RECT 301.950 459.600 304.050 460.050 ;
        RECT 736.950 459.600 739.050 460.050 ;
        RECT 271.950 458.400 304.050 459.600 ;
        RECT 271.950 457.950 274.050 458.400 ;
        RECT 301.950 457.950 304.050 458.400 ;
        RECT 689.400 458.400 739.050 459.600 ;
        RECT 85.950 456.600 88.050 456.900 ;
        RECT 100.950 456.600 103.050 457.050 ;
        RECT 85.950 455.400 103.050 456.600 ;
        RECT 85.950 454.800 88.050 455.400 ;
        RECT 100.950 454.950 103.050 455.400 ;
        RECT 274.950 456.600 277.050 457.050 ;
        RECT 283.950 456.600 286.050 457.050 ;
        RECT 274.950 455.400 286.050 456.600 ;
        RECT 274.950 454.950 277.050 455.400 ;
        RECT 283.950 454.950 286.050 455.400 ;
        RECT 328.950 456.600 331.050 457.050 ;
        RECT 334.950 456.600 337.050 457.050 ;
        RECT 394.950 456.600 397.050 457.050 ;
        RECT 328.950 455.400 397.050 456.600 ;
        RECT 328.950 454.950 331.050 455.400 ;
        RECT 334.950 454.950 337.050 455.400 ;
        RECT 394.950 454.950 397.050 455.400 ;
        RECT 433.950 456.600 436.050 457.050 ;
        RECT 508.950 456.600 511.050 457.050 ;
        RECT 433.950 455.400 511.050 456.600 ;
        RECT 433.950 454.950 436.050 455.400 ;
        RECT 508.950 454.950 511.050 455.400 ;
        RECT 541.950 456.600 544.050 457.050 ;
        RECT 565.950 456.600 568.050 457.050 ;
        RECT 541.950 455.400 568.050 456.600 ;
        RECT 541.950 454.950 544.050 455.400 ;
        RECT 565.950 454.950 568.050 455.400 ;
        RECT 601.950 456.600 604.050 457.050 ;
        RECT 649.950 456.600 652.050 457.050 ;
        RECT 689.400 456.600 690.600 458.400 ;
        RECT 736.950 457.950 739.050 458.400 ;
        RECT 601.950 455.400 690.600 456.600 ;
        RECT 691.950 456.600 694.050 457.050 ;
        RECT 706.950 456.600 709.050 457.050 ;
        RECT 691.950 455.400 709.050 456.600 ;
        RECT 601.950 454.950 604.050 455.400 ;
        RECT 649.950 454.950 652.050 455.400 ;
        RECT 691.950 454.950 694.050 455.400 ;
        RECT 706.950 454.950 709.050 455.400 ;
        RECT 760.950 456.600 763.050 457.050 ;
        RECT 769.950 456.600 772.050 457.050 ;
        RECT 781.950 456.600 784.050 457.050 ;
        RECT 760.950 455.400 784.050 456.600 ;
        RECT 760.950 454.950 763.050 455.400 ;
        RECT 769.950 454.950 772.050 455.400 ;
        RECT 781.950 454.950 784.050 455.400 ;
        RECT 844.950 456.600 847.050 457.050 ;
        RECT 865.950 456.600 868.050 457.050 ;
        RECT 844.950 455.400 868.050 456.600 ;
        RECT 844.950 454.950 847.050 455.400 ;
        RECT 865.950 454.950 868.050 455.400 ;
        RECT 4.950 453.600 7.050 454.050 ;
        RECT 16.950 453.600 19.050 454.050 ;
        RECT 4.950 452.400 19.050 453.600 ;
        RECT 4.950 451.950 7.050 452.400 ;
        RECT 16.950 451.950 19.050 452.400 ;
        RECT 22.950 453.600 25.050 454.050 ;
        RECT 40.950 453.600 43.050 454.050 ;
        RECT 22.950 452.400 43.050 453.600 ;
        RECT 22.950 451.950 25.050 452.400 ;
        RECT 40.950 451.950 43.050 452.400 ;
        RECT 136.950 453.600 139.050 454.050 ;
        RECT 148.950 453.600 151.050 454.050 ;
        RECT 136.950 452.400 151.050 453.600 ;
        RECT 136.950 451.950 139.050 452.400 ;
        RECT 148.950 451.950 151.050 452.400 ;
        RECT 322.950 453.600 325.050 454.050 ;
        RECT 340.950 453.600 343.050 454.050 ;
        RECT 361.950 453.600 364.050 454.050 ;
        RECT 367.950 453.600 370.050 454.050 ;
        RECT 484.950 453.600 487.050 454.050 ;
        RECT 322.950 452.400 370.050 453.600 ;
        RECT 322.950 451.950 325.050 452.400 ;
        RECT 340.950 451.950 343.050 452.400 ;
        RECT 361.950 451.950 364.050 452.400 ;
        RECT 367.950 451.950 370.050 452.400 ;
        RECT 440.400 452.400 487.050 453.600 ;
        RECT 440.400 451.200 441.600 452.400 ;
        RECT 484.950 451.950 487.050 452.400 ;
        RECT 751.950 453.600 754.050 454.050 ;
        RECT 769.950 453.600 772.050 453.900 ;
        RECT 751.950 452.400 772.050 453.600 ;
        RECT 751.950 451.950 754.050 452.400 ;
        RECT 769.950 451.800 772.050 452.400 ;
        RECT 796.950 453.600 799.050 454.050 ;
        RECT 805.950 453.600 808.050 454.050 ;
        RECT 823.950 453.600 826.050 454.050 ;
        RECT 829.950 453.600 832.050 454.050 ;
        RECT 796.950 452.400 832.050 453.600 ;
        RECT 796.950 451.950 799.050 452.400 ;
        RECT 805.950 451.950 808.050 452.400 ;
        RECT 823.950 451.950 826.050 452.400 ;
        RECT 829.950 451.950 832.050 452.400 ;
        RECT 18.000 450.600 22.050 451.050 ;
        RECT 17.400 448.950 22.050 450.600 ;
        RECT 31.950 450.600 34.050 451.200 ;
        RECT 58.950 450.600 61.050 451.050 ;
        RECT 31.950 449.400 61.050 450.600 ;
        RECT 31.950 449.100 34.050 449.400 ;
        RECT 58.950 448.950 61.050 449.400 ;
        RECT 67.950 450.600 70.050 451.200 ;
        RECT 94.950 450.750 97.050 451.200 ;
        RECT 103.950 450.750 106.050 451.200 ;
        RECT 94.950 450.600 106.050 450.750 ;
        RECT 67.950 449.550 106.050 450.600 ;
        RECT 67.950 449.400 97.050 449.550 ;
        RECT 67.950 449.100 70.050 449.400 ;
        RECT 94.950 449.100 97.050 449.400 ;
        RECT 103.950 449.100 106.050 449.550 ;
        RECT 109.950 450.750 112.050 451.200 ;
        RECT 115.950 450.750 118.050 451.200 ;
        RECT 109.950 449.550 118.050 450.750 ;
        RECT 109.950 449.100 112.050 449.550 ;
        RECT 115.950 449.100 118.050 449.550 ;
        RECT 127.950 450.600 130.050 451.200 ;
        RECT 160.950 450.600 163.050 451.200 ;
        RECT 166.950 450.600 169.050 451.200 ;
        RECT 178.950 450.600 181.050 451.200 ;
        RECT 127.950 449.400 163.050 450.600 ;
        RECT 127.950 449.100 130.050 449.400 ;
        RECT 160.950 449.100 163.050 449.400 ;
        RECT 164.400 449.400 181.050 450.600 ;
        RECT 17.400 444.900 18.600 448.950 ;
        RECT 164.400 447.600 165.600 449.400 ;
        RECT 166.950 449.100 169.050 449.400 ;
        RECT 178.950 449.100 181.050 449.400 ;
        RECT 184.950 449.100 187.050 451.200 ;
        RECT 199.950 449.100 202.050 451.200 ;
        RECT 220.950 450.600 223.050 451.050 ;
        RECT 226.950 450.600 229.050 451.200 ;
        RECT 220.950 449.400 229.050 450.600 ;
        RECT 101.400 446.400 108.600 447.600 ;
        RECT 16.950 442.800 19.050 444.900 ;
        RECT 49.950 444.600 52.050 444.900 ;
        RECT 64.950 444.600 67.050 444.900 ;
        RECT 49.950 443.400 67.050 444.600 ;
        RECT 49.950 442.800 52.050 443.400 ;
        RECT 64.950 442.800 67.050 443.400 ;
        RECT 88.950 444.600 91.050 444.900 ;
        RECT 94.950 444.600 97.050 445.050 ;
        RECT 101.400 444.900 102.600 446.400 ;
        RECT 88.950 443.400 97.050 444.600 ;
        RECT 88.950 442.800 91.050 443.400 ;
        RECT 94.950 442.950 97.050 443.400 ;
        RECT 100.950 442.800 103.050 444.900 ;
        RECT 107.400 444.600 108.600 446.400 ;
        RECT 161.400 446.400 165.600 447.600 ;
        RECT 130.950 444.600 133.050 445.050 ;
        RECT 107.400 443.400 133.050 444.600 ;
        RECT 130.950 442.950 133.050 443.400 ;
        RECT 145.950 444.600 148.050 444.900 ;
        RECT 161.400 444.600 162.600 446.400 ;
        RECT 145.950 443.400 162.600 444.600 ;
        RECT 175.950 444.600 178.050 445.050 ;
        RECT 185.400 444.600 186.600 449.100 ;
        RECT 175.950 443.400 186.600 444.600 ;
        RECT 187.950 444.600 190.050 444.900 ;
        RECT 200.400 444.600 201.600 449.100 ;
        RECT 220.950 448.950 223.050 449.400 ;
        RECT 226.950 449.100 229.050 449.400 ;
        RECT 277.950 450.600 280.050 451.200 ;
        RECT 292.950 450.600 295.050 451.200 ;
        RECT 277.950 449.400 295.050 450.600 ;
        RECT 277.950 449.100 280.050 449.400 ;
        RECT 292.950 449.100 295.050 449.400 ;
        RECT 370.950 450.750 373.050 451.200 ;
        RECT 409.950 450.750 412.050 451.200 ;
        RECT 370.950 449.550 412.050 450.750 ;
        RECT 370.950 449.100 373.050 449.550 ;
        RECT 409.950 449.100 412.050 449.550 ;
        RECT 415.950 449.100 418.050 451.200 ;
        RECT 421.950 450.600 424.050 451.200 ;
        RECT 439.950 450.600 442.050 451.200 ;
        RECT 421.950 449.400 442.050 450.600 ;
        RECT 421.950 449.100 424.050 449.400 ;
        RECT 439.950 449.100 442.050 449.400 ;
        RECT 448.950 450.600 451.050 451.050 ;
        RECT 454.950 450.600 457.050 451.200 ;
        RECT 448.950 449.400 457.050 450.600 ;
        RECT 416.400 447.600 417.600 449.100 ;
        RECT 448.950 448.950 451.050 449.400 ;
        RECT 454.950 449.100 457.050 449.400 ;
        RECT 472.950 450.750 475.050 451.200 ;
        RECT 478.950 450.750 481.050 451.200 ;
        RECT 472.950 449.550 481.050 450.750 ;
        RECT 520.950 450.600 523.050 451.200 ;
        RECT 544.950 450.600 547.050 451.200 ;
        RECT 472.950 449.100 475.050 449.550 ;
        RECT 478.950 449.100 481.050 449.550 ;
        RECT 509.400 449.400 547.050 450.600 ;
        RECT 407.400 446.400 417.600 447.600 ;
        RECT 187.950 443.400 201.600 444.600 ;
        RECT 244.950 444.450 247.050 444.900 ;
        RECT 250.950 444.450 253.050 444.900 ;
        RECT 145.950 442.800 148.050 443.400 ;
        RECT 175.950 442.950 178.050 443.400 ;
        RECT 187.950 442.800 190.050 443.400 ;
        RECT 244.950 443.250 253.050 444.450 ;
        RECT 244.950 442.800 247.050 443.250 ;
        RECT 250.950 442.800 253.050 443.250 ;
        RECT 283.950 444.450 286.050 444.900 ;
        RECT 289.950 444.450 292.050 444.900 ;
        RECT 283.950 443.250 292.050 444.450 ;
        RECT 283.950 442.800 286.050 443.250 ;
        RECT 289.950 442.800 292.050 443.250 ;
        RECT 295.950 444.600 298.050 445.050 ;
        RECT 325.950 444.600 328.050 444.900 ;
        RECT 295.950 443.400 328.050 444.600 ;
        RECT 295.950 442.950 298.050 443.400 ;
        RECT 325.950 442.800 328.050 443.400 ;
        RECT 334.950 444.450 337.050 444.900 ;
        RECT 352.950 444.450 355.050 444.900 ;
        RECT 334.950 443.250 355.050 444.450 ;
        RECT 334.950 442.800 337.050 443.250 ;
        RECT 352.950 442.800 355.050 443.250 ;
        RECT 397.950 444.600 400.050 444.900 ;
        RECT 407.400 444.600 408.600 446.400 ;
        RECT 397.950 443.400 408.600 444.600 ;
        RECT 409.950 444.600 412.050 445.050 ;
        RECT 418.950 444.600 421.050 444.900 ;
        RECT 409.950 443.400 421.050 444.600 ;
        RECT 397.950 442.800 400.050 443.400 ;
        RECT 409.950 442.950 412.050 443.400 ;
        RECT 418.950 442.800 421.050 443.400 ;
        RECT 424.950 444.450 427.050 444.900 ;
        RECT 433.950 444.450 436.050 444.900 ;
        RECT 424.950 443.250 436.050 444.450 ;
        RECT 424.950 442.800 427.050 443.250 ;
        RECT 433.950 442.800 436.050 443.250 ;
        RECT 457.950 444.600 460.050 444.900 ;
        RECT 472.950 444.600 475.050 445.050 ;
        RECT 509.400 444.900 510.600 449.400 ;
        RECT 520.950 449.100 523.050 449.400 ;
        RECT 544.950 449.100 547.050 449.400 ;
        RECT 571.950 449.100 574.050 451.200 ;
        RECT 595.950 450.750 598.050 451.200 ;
        RECT 601.950 450.750 604.050 451.200 ;
        RECT 595.950 449.550 604.050 450.750 ;
        RECT 595.950 449.100 598.050 449.550 ;
        RECT 601.950 449.100 604.050 449.550 ;
        RECT 610.950 450.600 613.050 451.200 ;
        RECT 625.950 450.600 628.050 451.200 ;
        RECT 610.950 449.400 628.050 450.600 ;
        RECT 610.950 449.100 613.050 449.400 ;
        RECT 625.950 449.100 628.050 449.400 ;
        RECT 637.950 450.750 640.050 451.200 ;
        RECT 643.950 450.750 646.050 451.200 ;
        RECT 637.950 449.550 646.050 450.750 ;
        RECT 637.950 449.100 640.050 449.550 ;
        RECT 643.950 449.100 646.050 449.550 ;
        RECT 700.950 449.100 703.050 451.200 ;
        RECT 706.950 450.600 709.050 451.200 ;
        RECT 712.950 450.750 715.050 451.200 ;
        RECT 718.950 450.750 721.050 451.200 ;
        RECT 712.950 450.600 721.050 450.750 ;
        RECT 706.950 449.550 721.050 450.600 ;
        RECT 706.950 449.400 715.050 449.550 ;
        RECT 706.950 449.100 709.050 449.400 ;
        RECT 712.950 449.100 715.050 449.400 ;
        RECT 718.950 449.100 721.050 449.550 ;
        RECT 754.950 449.100 757.050 451.200 ;
        RECT 766.950 450.600 769.050 451.050 ;
        RECT 761.400 449.400 769.050 450.600 ;
        RECT 457.950 443.400 475.050 444.600 ;
        RECT 457.950 442.800 460.050 443.400 ;
        RECT 472.950 442.950 475.050 443.400 ;
        RECT 508.950 442.800 511.050 444.900 ;
        RECT 136.950 441.600 139.050 442.050 ;
        RECT 142.950 441.600 145.050 442.050 ;
        RECT 136.950 440.400 145.050 441.600 ;
        RECT 136.950 439.950 139.050 440.400 ;
        RECT 142.950 439.950 145.050 440.400 ;
        RECT 163.950 441.600 166.050 442.050 ;
        RECT 172.950 441.600 175.050 442.050 ;
        RECT 223.950 441.600 226.050 442.050 ;
        RECT 163.950 440.400 175.050 441.600 ;
        RECT 163.950 439.950 166.050 440.400 ;
        RECT 172.950 439.950 175.050 440.400 ;
        RECT 191.400 440.400 226.050 441.600 ;
        RECT 58.950 438.600 61.050 439.050 ;
        RECT 106.950 438.600 109.050 439.050 ;
        RECT 58.950 437.400 109.050 438.600 ;
        RECT 58.950 436.950 61.050 437.400 ;
        RECT 106.950 436.950 109.050 437.400 ;
        RECT 115.950 438.600 118.050 439.050 ;
        RECT 191.400 438.600 192.600 440.400 ;
        RECT 223.950 439.950 226.050 440.400 ;
        RECT 253.950 441.600 256.050 442.050 ;
        RECT 496.950 441.600 499.050 442.050 ;
        RECT 502.950 441.600 505.050 442.050 ;
        RECT 253.950 440.400 264.600 441.600 ;
        RECT 253.950 439.950 256.050 440.400 ;
        RECT 115.950 437.400 192.600 438.600 ;
        RECT 220.950 438.600 223.050 439.050 ;
        RECT 256.950 438.600 259.050 439.050 ;
        RECT 220.950 437.400 259.050 438.600 ;
        RECT 263.400 438.600 264.600 440.400 ;
        RECT 496.950 440.400 505.050 441.600 ;
        RECT 496.950 439.950 499.050 440.400 ;
        RECT 502.950 439.950 505.050 440.400 ;
        RECT 523.950 441.600 526.050 442.050 ;
        RECT 535.950 441.600 538.050 442.050 ;
        RECT 523.950 440.400 538.050 441.600 ;
        RECT 523.950 439.950 526.050 440.400 ;
        RECT 535.950 439.950 538.050 440.400 ;
        RECT 343.950 438.600 346.050 439.050 ;
        RECT 263.400 437.400 346.050 438.600 ;
        RECT 115.950 436.950 118.050 437.400 ;
        RECT 220.950 436.950 223.050 437.400 ;
        RECT 256.950 436.950 259.050 437.400 ;
        RECT 343.950 436.950 346.050 437.400 ;
        RECT 403.950 438.600 406.050 439.050 ;
        RECT 412.950 438.600 415.050 439.050 ;
        RECT 430.950 438.600 433.050 439.050 ;
        RECT 463.950 438.600 466.050 439.050 ;
        RECT 403.950 437.400 466.050 438.600 ;
        RECT 403.950 436.950 406.050 437.400 ;
        RECT 412.950 436.950 415.050 437.400 ;
        RECT 430.950 436.950 433.050 437.400 ;
        RECT 463.950 436.950 466.050 437.400 ;
        RECT 487.950 438.600 490.050 439.050 ;
        RECT 524.400 438.600 525.600 439.950 ;
        RECT 487.950 437.400 525.600 438.600 ;
        RECT 572.400 438.600 573.600 449.100 ;
        RECT 691.950 447.600 694.050 448.050 ;
        RECT 677.400 446.400 694.050 447.600 ;
        RECT 574.950 444.600 577.050 444.900 ;
        RECT 580.950 444.600 583.050 445.050 ;
        RECT 574.950 443.400 583.050 444.600 ;
        RECT 574.950 442.800 577.050 443.400 ;
        RECT 580.950 442.950 583.050 443.400 ;
        RECT 616.950 444.600 619.050 445.050 ;
        RECT 622.950 444.600 625.050 444.900 ;
        RECT 616.950 443.400 625.050 444.600 ;
        RECT 616.950 442.950 619.050 443.400 ;
        RECT 622.950 442.800 625.050 443.400 ;
        RECT 646.950 444.600 649.050 444.900 ;
        RECT 655.950 444.600 658.050 445.050 ;
        RECT 661.950 444.600 664.050 444.900 ;
        RECT 646.950 443.400 664.050 444.600 ;
        RECT 646.950 442.800 649.050 443.400 ;
        RECT 655.950 442.950 658.050 443.400 ;
        RECT 661.950 442.800 664.050 443.400 ;
        RECT 667.950 444.600 670.050 444.900 ;
        RECT 677.400 444.600 678.600 446.400 ;
        RECT 691.950 445.950 694.050 446.400 ;
        RECT 667.950 443.400 678.600 444.600 ;
        RECT 682.950 444.600 685.050 444.900 ;
        RECT 701.400 444.600 702.600 449.100 ;
        RECT 755.400 445.050 756.600 449.100 ;
        RECT 682.950 443.400 702.600 444.600 ;
        RECT 730.950 444.600 733.050 445.050 ;
        RECT 739.950 444.600 742.050 444.900 ;
        RECT 730.950 443.400 742.050 444.600 ;
        RECT 667.950 442.800 670.050 443.400 ;
        RECT 682.950 442.800 685.050 443.400 ;
        RECT 730.950 442.950 733.050 443.400 ;
        RECT 739.950 442.800 742.050 443.400 ;
        RECT 751.950 443.400 756.600 445.050 ;
        RECT 751.950 442.950 756.000 443.400 ;
        RECT 761.400 442.050 762.600 449.400 ;
        RECT 766.950 448.950 769.050 449.400 ;
        RECT 802.950 449.100 805.050 451.200 ;
        RECT 811.950 450.600 814.050 451.050 ;
        RECT 820.950 450.600 823.050 451.200 ;
        RECT 811.950 449.400 823.050 450.600 ;
        RECT 803.400 444.600 804.600 449.100 ;
        RECT 811.950 448.950 814.050 449.400 ;
        RECT 820.950 449.100 823.050 449.400 ;
        RECT 847.950 450.600 850.050 451.050 ;
        RECT 859.950 450.600 862.050 451.200 ;
        RECT 847.950 449.400 862.050 450.600 ;
        RECT 847.950 448.950 850.050 449.400 ;
        RECT 859.950 449.100 862.050 449.400 ;
        RECT 865.950 450.750 868.050 451.200 ;
        RECT 871.950 450.750 874.050 451.200 ;
        RECT 865.950 449.550 874.050 450.750 ;
        RECT 865.950 449.100 868.050 449.550 ;
        RECT 871.950 449.100 874.050 449.550 ;
        RECT 823.950 444.600 826.050 444.900 ;
        RECT 803.400 443.400 826.050 444.600 ;
        RECT 823.950 442.800 826.050 443.400 ;
        RECT 841.950 444.450 844.050 444.900 ;
        RECT 847.950 444.450 850.050 444.900 ;
        RECT 841.950 443.250 850.050 444.450 ;
        RECT 841.950 442.800 844.050 443.250 ;
        RECT 847.950 442.800 850.050 443.250 ;
        RECT 691.950 441.600 694.050 442.050 ;
        RECT 703.950 441.600 706.050 442.050 ;
        RECT 691.950 440.400 706.050 441.600 ;
        RECT 691.950 439.950 694.050 440.400 ;
        RECT 703.950 439.950 706.050 440.400 ;
        RECT 760.950 439.950 763.050 442.050 ;
        RECT 772.950 441.600 775.050 442.050 ;
        RECT 781.950 441.600 784.050 442.050 ;
        RECT 772.950 440.400 784.050 441.600 ;
        RECT 772.950 439.950 775.050 440.400 ;
        RECT 781.950 439.950 784.050 440.400 ;
        RECT 829.950 441.600 832.050 442.050 ;
        RECT 862.950 441.600 865.050 442.050 ;
        RECT 829.950 440.400 865.050 441.600 ;
        RECT 829.950 439.950 832.050 440.400 ;
        RECT 862.950 439.950 865.050 440.400 ;
        RECT 586.950 438.600 589.050 439.050 ;
        RECT 572.400 437.400 589.050 438.600 ;
        RECT 487.950 436.950 490.050 437.400 ;
        RECT 586.950 436.950 589.050 437.400 ;
        RECT 595.950 438.600 598.050 439.050 ;
        RECT 601.950 438.600 604.050 439.050 ;
        RECT 607.950 438.600 610.050 439.050 ;
        RECT 595.950 437.400 610.050 438.600 ;
        RECT 595.950 436.950 598.050 437.400 ;
        RECT 601.950 436.950 604.050 437.400 ;
        RECT 607.950 436.950 610.050 437.400 ;
        RECT 694.950 438.600 697.050 439.050 ;
        RECT 721.950 438.600 724.050 439.050 ;
        RECT 694.950 437.400 724.050 438.600 ;
        RECT 694.950 436.950 697.050 437.400 ;
        RECT 721.950 436.950 724.050 437.400 ;
        RECT 748.950 438.600 751.050 439.050 ;
        RECT 757.950 438.600 760.050 439.050 ;
        RECT 748.950 437.400 760.050 438.600 ;
        RECT 748.950 436.950 751.050 437.400 ;
        RECT 757.950 436.950 760.050 437.400 ;
        RECT 133.950 435.600 136.050 436.050 ;
        RECT 169.950 435.600 172.050 436.050 ;
        RECT 202.950 435.600 205.050 436.050 ;
        RECT 208.950 435.600 211.050 436.050 ;
        RECT 133.950 434.400 211.050 435.600 ;
        RECT 133.950 433.950 136.050 434.400 ;
        RECT 169.950 433.950 172.050 434.400 ;
        RECT 202.950 433.950 205.050 434.400 ;
        RECT 208.950 433.950 211.050 434.400 ;
        RECT 223.950 435.600 226.050 436.050 ;
        RECT 253.950 435.600 256.050 436.050 ;
        RECT 223.950 434.400 256.050 435.600 ;
        RECT 223.950 433.950 226.050 434.400 ;
        RECT 253.950 433.950 256.050 434.400 ;
        RECT 265.950 435.600 268.050 436.050 ;
        RECT 295.950 435.600 298.050 436.050 ;
        RECT 265.950 434.400 298.050 435.600 ;
        RECT 265.950 433.950 268.050 434.400 ;
        RECT 295.950 433.950 298.050 434.400 ;
        RECT 301.950 435.600 304.050 436.050 ;
        RECT 307.950 435.600 310.050 436.050 ;
        RECT 301.950 434.400 310.050 435.600 ;
        RECT 301.950 433.950 304.050 434.400 ;
        RECT 307.950 433.950 310.050 434.400 ;
        RECT 313.950 435.600 316.050 436.050 ;
        RECT 712.950 435.600 715.050 436.050 ;
        RECT 721.950 435.600 724.050 435.900 ;
        RECT 313.950 434.400 420.600 435.600 ;
        RECT 313.950 433.950 316.050 434.400 ;
        RECT 31.950 432.600 34.050 433.050 ;
        RECT 419.400 432.600 420.600 434.400 ;
        RECT 712.950 434.400 724.050 435.600 ;
        RECT 712.950 433.950 715.050 434.400 ;
        RECT 721.950 433.800 724.050 434.400 ;
        RECT 823.950 435.600 826.050 436.050 ;
        RECT 832.950 435.600 835.050 436.050 ;
        RECT 850.950 435.600 853.050 436.050 ;
        RECT 823.950 434.400 853.050 435.600 ;
        RECT 823.950 433.950 826.050 434.400 ;
        RECT 832.950 433.950 835.050 434.400 ;
        RECT 850.950 433.950 853.050 434.400 ;
        RECT 442.950 432.600 445.050 433.050 ;
        RECT 31.950 431.400 312.600 432.600 ;
        RECT 419.400 431.400 445.050 432.600 ;
        RECT 31.950 430.950 34.050 431.400 ;
        RECT 311.400 430.050 312.600 431.400 ;
        RECT 442.950 430.950 445.050 431.400 ;
        RECT 592.950 432.600 595.050 433.050 ;
        RECT 628.950 432.600 631.050 433.050 ;
        RECT 637.950 432.600 640.050 433.050 ;
        RECT 724.950 432.600 727.050 433.050 ;
        RECT 592.950 431.400 727.050 432.600 ;
        RECT 592.950 430.950 595.050 431.400 ;
        RECT 628.950 430.950 631.050 431.400 ;
        RECT 637.950 430.950 640.050 431.400 ;
        RECT 724.950 430.950 727.050 431.400 ;
        RECT 769.950 432.600 772.050 433.050 ;
        RECT 799.950 432.600 802.050 433.050 ;
        RECT 769.950 431.400 802.050 432.600 ;
        RECT 769.950 430.950 772.050 431.400 ;
        RECT 799.950 430.950 802.050 431.400 ;
        RECT 811.950 432.600 814.050 433.050 ;
        RECT 820.950 432.600 823.050 433.050 ;
        RECT 811.950 431.400 823.050 432.600 ;
        RECT 811.950 430.950 814.050 431.400 ;
        RECT 820.950 430.950 823.050 431.400 ;
        RECT 7.950 429.600 10.050 430.050 ;
        RECT 19.950 429.600 22.050 430.050 ;
        RECT 7.950 428.400 22.050 429.600 ;
        RECT 7.950 427.950 10.050 428.400 ;
        RECT 19.950 427.950 22.050 428.400 ;
        RECT 181.950 429.600 184.050 430.050 ;
        RECT 241.950 429.600 244.050 430.050 ;
        RECT 181.950 428.400 244.050 429.600 ;
        RECT 181.950 427.950 184.050 428.400 ;
        RECT 241.950 427.950 244.050 428.400 ;
        RECT 310.950 429.600 313.050 430.050 ;
        RECT 355.950 429.600 358.050 430.050 ;
        RECT 310.950 428.400 358.050 429.600 ;
        RECT 310.950 427.950 313.050 428.400 ;
        RECT 355.950 427.950 358.050 428.400 ;
        RECT 361.950 429.600 364.050 430.050 ;
        RECT 370.950 429.600 373.050 430.050 ;
        RECT 361.950 428.400 373.050 429.600 ;
        RECT 361.950 427.950 364.050 428.400 ;
        RECT 370.950 427.950 373.050 428.400 ;
        RECT 517.950 429.600 520.050 430.050 ;
        RECT 529.950 429.600 532.050 430.050 ;
        RECT 517.950 428.400 532.050 429.600 ;
        RECT 517.950 427.950 520.050 428.400 ;
        RECT 529.950 427.950 532.050 428.400 ;
        RECT 184.950 426.600 187.050 427.050 ;
        RECT 190.950 426.600 193.050 427.050 ;
        RECT 184.950 425.400 193.050 426.600 ;
        RECT 184.950 424.950 187.050 425.400 ;
        RECT 190.950 424.950 193.050 425.400 ;
        RECT 304.950 426.600 307.050 427.050 ;
        RECT 313.950 426.600 316.050 427.050 ;
        RECT 304.950 425.400 316.050 426.600 ;
        RECT 304.950 424.950 307.050 425.400 ;
        RECT 313.950 424.950 316.050 425.400 ;
        RECT 655.950 426.600 658.050 427.050 ;
        RECT 688.950 426.600 691.050 427.050 ;
        RECT 655.950 425.400 691.050 426.600 ;
        RECT 655.950 424.950 658.050 425.400 ;
        RECT 688.950 424.950 691.050 425.400 ;
        RECT 694.950 426.600 697.050 427.050 ;
        RECT 712.950 426.600 715.050 427.050 ;
        RECT 694.950 425.400 715.050 426.600 ;
        RECT 694.950 424.950 697.050 425.400 ;
        RECT 712.950 424.950 715.050 425.400 ;
        RECT 718.950 426.600 721.050 427.050 ;
        RECT 733.950 426.600 736.050 427.050 ;
        RECT 718.950 425.400 736.050 426.600 ;
        RECT 718.950 424.950 721.050 425.400 ;
        RECT 733.950 424.950 736.050 425.400 ;
        RECT 757.950 426.600 760.050 427.050 ;
        RECT 793.950 426.600 796.050 427.050 ;
        RECT 757.950 425.400 796.050 426.600 ;
        RECT 757.950 424.950 760.050 425.400 ;
        RECT 793.950 424.950 796.050 425.400 ;
        RECT 817.950 426.600 820.050 427.050 ;
        RECT 832.950 426.600 835.050 427.050 ;
        RECT 817.950 425.400 835.050 426.600 ;
        RECT 817.950 424.950 820.050 425.400 ;
        RECT 832.950 424.950 835.050 425.400 ;
        RECT 853.950 426.600 856.050 427.050 ;
        RECT 868.950 426.600 871.050 427.050 ;
        RECT 853.950 425.400 871.050 426.600 ;
        RECT 853.950 424.950 856.050 425.400 ;
        RECT 868.950 424.950 871.050 425.400 ;
        RECT 355.950 423.600 358.050 424.050 ;
        RECT 445.950 423.600 448.050 424.050 ;
        RECT 499.950 423.600 502.050 424.050 ;
        RECT 550.950 423.600 553.050 424.050 ;
        RECT 553.950 423.600 556.050 424.050 ;
        RECT 355.950 422.400 556.050 423.600 ;
        RECT 355.950 421.950 358.050 422.400 ;
        RECT 445.950 421.950 448.050 422.400 ;
        RECT 499.950 421.950 502.050 422.400 ;
        RECT 550.950 421.950 553.050 422.400 ;
        RECT 553.950 421.950 556.050 422.400 ;
        RECT 571.950 423.600 574.050 424.050 ;
        RECT 598.950 423.600 601.050 424.050 ;
        RECT 571.950 422.400 601.050 423.600 ;
        RECT 571.950 421.950 574.050 422.400 ;
        RECT 598.950 421.950 601.050 422.400 ;
        RECT 715.950 423.600 718.050 424.050 ;
        RECT 736.950 423.600 739.050 423.900 ;
        RECT 715.950 422.400 739.050 423.600 ;
        RECT 715.950 421.950 718.050 422.400 ;
        RECT 736.950 421.800 739.050 422.400 ;
        RECT 742.950 423.600 745.050 424.050 ;
        RECT 751.950 423.600 754.050 424.050 ;
        RECT 811.950 423.600 814.050 424.050 ;
        RECT 742.950 422.400 814.050 423.600 ;
        RECT 742.950 421.950 745.050 422.400 ;
        RECT 751.950 421.950 754.050 422.400 ;
        RECT 811.950 421.950 814.050 422.400 ;
        RECT 4.950 420.600 7.050 421.050 ;
        RECT 22.950 420.600 25.050 421.050 ;
        RECT 4.950 419.400 25.050 420.600 ;
        RECT 4.950 418.950 7.050 419.400 ;
        RECT 22.950 418.950 25.050 419.400 ;
        RECT 73.950 420.600 76.050 421.050 ;
        RECT 82.950 420.600 85.050 421.050 ;
        RECT 73.950 419.400 85.050 420.600 ;
        RECT 73.950 418.950 76.050 419.400 ;
        RECT 82.950 418.950 85.050 419.400 ;
        RECT 133.950 418.950 136.050 421.050 ;
        RECT 163.950 420.600 166.050 421.050 ;
        RECT 178.950 420.600 181.050 421.050 ;
        RECT 163.950 419.400 181.050 420.600 ;
        RECT 163.950 418.950 166.050 419.400 ;
        RECT 178.950 418.950 181.050 419.400 ;
        RECT 211.950 420.600 214.050 421.050 ;
        RECT 223.950 420.600 226.050 421.050 ;
        RECT 244.950 420.600 247.050 421.050 ;
        RECT 211.950 419.400 247.050 420.600 ;
        RECT 211.950 418.950 214.050 419.400 ;
        RECT 223.950 418.950 226.050 419.400 ;
        RECT 244.950 418.950 247.050 419.400 ;
        RECT 283.950 420.600 286.050 421.050 ;
        RECT 301.950 420.600 304.050 421.050 ;
        RECT 283.950 419.400 304.050 420.600 ;
        RECT 283.950 418.950 286.050 419.400 ;
        RECT 301.950 418.950 304.050 419.400 ;
        RECT 307.950 420.600 310.050 421.050 ;
        RECT 322.950 420.600 325.050 421.050 ;
        RECT 307.950 419.400 325.050 420.600 ;
        RECT 307.950 418.950 310.050 419.400 ;
        RECT 322.950 418.950 325.050 419.400 ;
        RECT 436.950 420.600 439.050 421.050 ;
        RECT 442.950 420.600 445.050 421.050 ;
        RECT 436.950 419.400 445.050 420.600 ;
        RECT 436.950 418.950 439.050 419.400 ;
        RECT 442.950 418.950 445.050 419.400 ;
        RECT 601.950 420.600 604.050 421.050 ;
        RECT 634.950 420.600 637.050 421.050 ;
        RECT 601.950 419.400 637.050 420.600 ;
        RECT 601.950 418.950 604.050 419.400 ;
        RECT 634.950 418.950 637.050 419.400 ;
        RECT 649.950 420.600 652.050 421.050 ;
        RECT 655.950 420.600 658.050 421.050 ;
        RECT 649.950 419.400 658.050 420.600 ;
        RECT 649.950 418.950 652.050 419.400 ;
        RECT 655.950 418.950 658.050 419.400 ;
        RECT 739.950 420.600 742.050 421.050 ;
        RECT 766.950 420.600 769.050 421.050 ;
        RECT 739.950 419.400 769.050 420.600 ;
        RECT 739.950 418.950 742.050 419.400 ;
        RECT 766.950 418.950 769.050 419.400 ;
        RECT 772.950 420.600 775.050 421.050 ;
        RECT 793.950 420.600 796.050 421.050 ;
        RECT 772.950 419.400 796.050 420.600 ;
        RECT 772.950 418.950 775.050 419.400 ;
        RECT 793.950 418.950 796.050 419.400 ;
        RECT 1.950 415.950 4.050 418.050 ;
        RECT 52.950 417.600 55.050 418.200 ;
        RECT 64.950 417.600 67.050 418.200 ;
        RECT 70.950 417.600 73.050 418.050 ;
        RECT 52.950 416.400 73.050 417.600 ;
        RECT 52.950 416.100 55.050 416.400 ;
        RECT 64.950 416.100 67.050 416.400 ;
        RECT 70.950 415.950 73.050 416.400 ;
        RECT 2.400 412.050 3.600 415.950 ;
        RECT 1.950 409.950 4.050 412.050 ;
        RECT 49.950 411.600 52.050 411.900 ;
        RECT 58.950 411.600 61.050 412.050 ;
        RECT 134.400 411.900 135.600 418.950 ;
        RECT 148.950 417.600 151.050 418.200 ;
        RECT 154.950 417.600 157.050 418.050 ;
        RECT 168.000 417.600 172.050 418.050 ;
        RECT 148.950 416.400 157.050 417.600 ;
        RECT 148.950 416.100 151.050 416.400 ;
        RECT 154.950 415.950 157.050 416.400 ;
        RECT 167.400 415.950 172.050 417.600 ;
        RECT 175.950 415.950 178.050 418.050 ;
        RECT 199.950 417.750 202.050 418.200 ;
        RECT 208.950 417.750 211.050 418.200 ;
        RECT 199.950 416.550 211.050 417.750 ;
        RECT 199.950 416.100 202.050 416.550 ;
        RECT 208.950 416.100 211.050 416.550 ;
        RECT 229.950 417.600 232.050 418.050 ;
        RECT 238.950 417.600 241.050 418.200 ;
        RECT 229.950 416.400 241.050 417.600 ;
        RECT 229.950 415.950 232.050 416.400 ;
        RECT 238.950 416.100 241.050 416.400 ;
        RECT 247.950 417.600 250.050 418.050 ;
        RECT 253.950 417.600 256.050 418.200 ;
        RECT 247.950 416.400 256.050 417.600 ;
        RECT 247.950 415.950 250.050 416.400 ;
        RECT 253.950 416.100 256.050 416.400 ;
        RECT 259.950 417.600 262.050 418.200 ;
        RECT 265.950 417.750 268.050 418.200 ;
        RECT 277.950 417.750 280.050 418.200 ;
        RECT 265.950 417.600 280.050 417.750 ;
        RECT 304.950 417.600 307.050 418.050 ;
        RECT 259.950 416.550 280.050 417.600 ;
        RECT 259.950 416.400 268.050 416.550 ;
        RECT 259.950 416.100 262.050 416.400 ;
        RECT 265.950 416.100 268.050 416.400 ;
        RECT 277.950 416.100 280.050 416.550 ;
        RECT 284.400 416.400 307.050 417.600 ;
        RECT 167.400 411.900 168.600 415.950 ;
        RECT 176.400 412.050 177.600 415.950 ;
        RECT 49.950 410.400 61.050 411.600 ;
        RECT 49.950 409.800 52.050 410.400 ;
        RECT 58.950 409.950 61.050 410.400 ;
        RECT 67.950 411.450 70.050 411.900 ;
        RECT 85.950 411.450 88.050 411.900 ;
        RECT 67.950 410.250 88.050 411.450 ;
        RECT 67.950 409.800 70.050 410.250 ;
        RECT 85.950 409.800 88.050 410.250 ;
        RECT 133.950 409.800 136.050 411.900 ;
        RECT 154.950 411.450 157.050 411.900 ;
        RECT 160.950 411.450 163.050 411.900 ;
        RECT 154.950 410.250 163.050 411.450 ;
        RECT 154.950 409.800 157.050 410.250 ;
        RECT 160.950 409.800 163.050 410.250 ;
        RECT 166.950 409.800 169.050 411.900 ;
        RECT 175.950 409.950 178.050 412.050 ;
        RECT 284.400 411.900 285.600 416.400 ;
        RECT 304.950 415.950 307.050 416.400 ;
        RECT 325.950 417.600 328.050 418.050 ;
        RECT 331.950 417.600 334.050 418.200 ;
        RECT 325.950 416.400 334.050 417.600 ;
        RECT 325.950 415.950 328.050 416.400 ;
        RECT 331.950 416.100 334.050 416.400 ;
        RECT 340.950 417.750 343.050 418.200 ;
        RECT 346.950 417.750 349.050 418.200 ;
        RECT 340.950 417.600 349.050 417.750 ;
        RECT 355.950 417.600 358.050 418.200 ;
        RECT 340.950 416.550 358.050 417.600 ;
        RECT 340.950 416.100 343.050 416.550 ;
        RECT 346.950 416.400 358.050 416.550 ;
        RECT 346.950 416.100 349.050 416.400 ;
        RECT 355.950 416.100 358.050 416.400 ;
        RECT 370.950 417.750 373.050 418.200 ;
        RECT 391.950 417.750 394.050 418.050 ;
        RECT 397.950 417.750 400.050 418.200 ;
        RECT 370.950 416.550 400.050 417.750 ;
        RECT 370.950 416.100 373.050 416.550 ;
        RECT 391.950 415.950 394.050 416.550 ;
        RECT 397.950 416.100 400.050 416.550 ;
        RECT 415.950 417.600 418.050 418.050 ;
        RECT 424.950 417.600 427.050 418.200 ;
        RECT 415.950 416.400 427.050 417.600 ;
        RECT 415.950 415.950 418.050 416.400 ;
        RECT 424.950 416.100 427.050 416.400 ;
        RECT 433.950 417.600 436.050 418.050 ;
        RECT 448.950 417.600 451.050 418.050 ;
        RECT 481.950 417.600 484.050 418.050 ;
        RECT 433.950 416.400 451.050 417.600 ;
        RECT 433.950 415.950 436.050 416.400 ;
        RECT 448.950 415.950 451.050 416.400 ;
        RECT 470.400 416.400 484.050 417.600 ;
        RECT 388.950 414.600 391.050 415.050 ;
        RECT 380.400 413.400 391.050 414.600 ;
        RECT 181.950 411.450 184.050 411.900 ;
        RECT 211.950 411.450 214.050 411.900 ;
        RECT 181.950 410.250 214.050 411.450 ;
        RECT 181.950 409.800 184.050 410.250 ;
        RECT 211.950 409.800 214.050 410.250 ;
        RECT 241.950 411.450 244.050 411.900 ;
        RECT 247.800 411.450 249.900 411.900 ;
        RECT 256.950 411.600 259.050 411.900 ;
        RECT 241.950 410.250 249.900 411.450 ;
        RECT 251.400 411.000 259.050 411.600 ;
        RECT 241.950 409.800 244.050 410.250 ;
        RECT 247.800 409.800 249.900 410.250 ;
        RECT 250.950 410.400 259.050 411.000 ;
        RECT 187.950 408.600 190.050 409.050 ;
        RECT 208.950 408.600 211.050 409.050 ;
        RECT 229.950 408.600 232.050 409.050 ;
        RECT 187.950 407.400 232.050 408.600 ;
        RECT 187.950 406.950 190.050 407.400 ;
        RECT 208.950 406.950 211.050 407.400 ;
        RECT 229.950 406.950 232.050 407.400 ;
        RECT 250.950 406.950 253.050 410.400 ;
        RECT 256.950 409.800 259.050 410.400 ;
        RECT 283.950 409.800 286.050 411.900 ;
        RECT 304.950 411.450 307.050 411.900 ;
        RECT 310.950 411.450 313.050 411.900 ;
        RECT 304.950 410.250 313.050 411.450 ;
        RECT 304.950 409.800 307.050 410.250 ;
        RECT 310.950 409.800 313.050 410.250 ;
        RECT 322.950 411.450 325.050 411.900 ;
        RECT 334.950 411.450 337.050 411.900 ;
        RECT 322.950 410.250 337.050 411.450 ;
        RECT 322.950 409.800 325.050 410.250 ;
        RECT 334.950 409.800 337.050 410.250 ;
        RECT 373.950 411.600 376.050 411.900 ;
        RECT 380.400 411.600 381.600 413.400 ;
        RECT 388.950 412.950 391.050 413.400 ;
        RECT 470.400 411.900 471.600 416.400 ;
        RECT 481.950 415.950 484.050 416.400 ;
        RECT 559.950 417.750 562.050 418.200 ;
        RECT 592.950 417.750 595.050 418.200 ;
        RECT 559.950 416.550 595.050 417.750 ;
        RECT 559.950 416.100 562.050 416.550 ;
        RECT 592.950 416.100 595.050 416.550 ;
        RECT 616.950 417.600 619.050 418.050 ;
        RECT 625.950 417.600 628.050 418.200 ;
        RECT 616.950 416.400 628.050 417.600 ;
        RECT 616.950 415.950 619.050 416.400 ;
        RECT 625.950 416.100 628.050 416.400 ;
        RECT 643.950 417.750 646.050 418.200 ;
        RECT 664.950 417.750 667.050 418.200 ;
        RECT 643.950 416.550 667.050 417.750 ;
        RECT 673.950 417.600 676.050 418.200 ;
        RECT 643.950 416.100 646.050 416.550 ;
        RECT 664.950 416.100 667.050 416.550 ;
        RECT 668.400 416.400 676.050 417.600 ;
        RECT 668.400 414.600 669.600 416.400 ;
        RECT 673.950 416.100 676.050 416.400 ;
        RECT 688.950 417.600 691.050 418.200 ;
        RECT 709.950 417.600 712.050 418.200 ;
        RECT 688.950 416.400 712.050 417.600 ;
        RECT 688.950 416.100 691.050 416.400 ;
        RECT 709.950 416.100 712.050 416.400 ;
        RECT 721.950 415.950 724.050 418.050 ;
        RECT 730.950 416.100 733.050 418.200 ;
        RECT 769.950 416.100 772.050 418.200 ;
        RECT 847.950 417.750 850.050 418.200 ;
        RECT 859.950 417.750 862.050 418.200 ;
        RECT 847.950 416.550 862.050 417.750 ;
        RECT 847.950 416.100 850.050 416.550 ;
        RECT 859.950 416.100 862.050 416.550 ;
        RECT 703.950 414.600 706.050 415.050 ;
        RECT 491.400 413.400 588.600 414.600 ;
        RECT 491.400 411.900 492.600 413.400 ;
        RECT 533.400 411.900 534.600 413.400 ;
        RECT 373.950 410.400 381.600 411.600 ;
        RECT 406.950 411.450 409.050 411.900 ;
        RECT 415.950 411.450 418.050 411.900 ;
        RECT 373.950 409.800 376.050 410.400 ;
        RECT 406.950 410.250 418.050 411.450 ;
        RECT 406.950 409.800 409.050 410.250 ;
        RECT 415.950 409.800 418.050 410.250 ;
        RECT 427.950 411.450 430.050 411.900 ;
        RECT 433.950 411.450 436.050 411.900 ;
        RECT 427.950 410.250 436.050 411.450 ;
        RECT 427.950 409.800 430.050 410.250 ;
        RECT 433.950 409.800 436.050 410.250 ;
        RECT 469.950 409.800 472.050 411.900 ;
        RECT 478.950 411.450 481.050 411.900 ;
        RECT 490.950 411.450 493.050 411.900 ;
        RECT 478.950 410.250 493.050 411.450 ;
        RECT 478.950 409.800 481.050 410.250 ;
        RECT 490.950 409.800 493.050 410.250 ;
        RECT 517.950 411.450 520.050 411.900 ;
        RECT 523.950 411.450 526.050 411.900 ;
        RECT 517.950 410.250 526.050 411.450 ;
        RECT 517.950 409.800 520.050 410.250 ;
        RECT 523.950 409.800 526.050 410.250 ;
        RECT 532.950 409.800 535.050 411.900 ;
        RECT 571.950 411.600 574.050 412.050 ;
        RECT 587.400 411.900 588.600 413.400 ;
        RECT 668.400 413.400 706.050 414.600 ;
        RECT 668.400 412.050 669.600 413.400 ;
        RECT 703.950 412.950 706.050 413.400 ;
        RECT 722.400 412.050 723.600 415.950 ;
        RECT 731.400 412.050 732.600 416.100 ;
        RECT 577.950 411.600 580.050 411.900 ;
        RECT 571.950 410.400 580.050 411.600 ;
        RECT 571.950 409.950 574.050 410.400 ;
        RECT 577.950 409.800 580.050 410.400 ;
        RECT 586.950 409.800 589.050 411.900 ;
        RECT 604.950 411.600 607.050 411.900 ;
        RECT 622.950 411.600 625.050 411.900 ;
        RECT 604.950 410.400 625.050 411.600 ;
        RECT 604.950 409.800 607.050 410.400 ;
        RECT 622.950 409.800 625.050 410.400 ;
        RECT 667.950 409.950 670.050 412.050 ;
        RECT 682.950 411.600 685.050 412.050 ;
        RECT 700.950 411.600 703.050 412.050 ;
        RECT 682.950 410.400 703.050 411.600 ;
        RECT 682.950 409.950 685.050 410.400 ;
        RECT 700.950 409.950 703.050 410.400 ;
        RECT 721.950 409.950 724.050 412.050 ;
        RECT 727.950 410.400 732.600 412.050 ;
        RECT 736.950 411.450 739.050 411.900 ;
        RECT 763.950 411.450 766.050 412.050 ;
        RECT 766.950 411.450 769.050 411.900 ;
        RECT 727.950 409.950 732.000 410.400 ;
        RECT 736.950 410.250 769.050 411.450 ;
        RECT 736.950 409.800 739.050 410.250 ;
        RECT 763.950 409.950 766.050 410.250 ;
        RECT 766.950 409.800 769.050 410.250 ;
        RECT 770.400 409.050 771.600 416.100 ;
        RECT 775.950 411.600 778.050 411.900 ;
        RECT 778.950 411.600 781.050 412.050 ;
        RECT 787.950 411.600 790.050 411.900 ;
        RECT 775.950 410.400 790.050 411.600 ;
        RECT 775.950 409.800 778.050 410.400 ;
        RECT 778.950 409.950 781.050 410.400 ;
        RECT 787.950 409.800 790.050 410.400 ;
        RECT 808.950 411.600 811.050 411.900 ;
        RECT 823.950 411.600 826.050 412.050 ;
        RECT 808.950 410.400 826.050 411.600 ;
        RECT 808.950 409.800 811.050 410.400 ;
        RECT 823.950 409.950 826.050 410.400 ;
        RECT 364.950 408.600 367.050 409.050 ;
        RECT 367.950 408.600 370.050 409.050 ;
        RECT 382.950 408.600 385.050 409.050 ;
        RECT 364.950 407.400 385.050 408.600 ;
        RECT 364.950 406.950 367.050 407.400 ;
        RECT 367.950 406.950 370.050 407.400 ;
        RECT 382.950 406.950 385.050 407.400 ;
        RECT 391.950 408.600 394.050 409.050 ;
        RECT 421.950 408.600 424.050 409.050 ;
        RECT 391.950 407.400 424.050 408.600 ;
        RECT 391.950 406.950 394.050 407.400 ;
        RECT 421.950 406.950 424.050 407.400 ;
        RECT 589.950 408.600 592.050 409.050 ;
        RECT 595.950 408.600 598.050 409.050 ;
        RECT 589.950 407.400 598.050 408.600 ;
        RECT 589.950 406.950 592.050 407.400 ;
        RECT 595.950 406.950 598.050 407.400 ;
        RECT 607.950 408.600 610.050 409.050 ;
        RECT 754.950 408.600 757.050 409.050 ;
        RECT 760.950 408.600 763.050 409.050 ;
        RECT 607.950 407.400 621.600 408.600 ;
        RECT 607.950 406.950 610.050 407.400 ;
        RECT 193.950 405.600 196.050 406.050 ;
        RECT 202.950 405.600 205.050 406.050 ;
        RECT 193.950 404.400 205.050 405.600 ;
        RECT 193.950 403.950 196.050 404.400 ;
        RECT 202.950 403.950 205.050 404.400 ;
        RECT 247.950 405.600 250.050 406.050 ;
        RECT 340.950 405.600 343.050 406.050 ;
        RECT 247.950 404.400 343.050 405.600 ;
        RECT 247.950 403.950 250.050 404.400 ;
        RECT 340.950 403.950 343.050 404.400 ;
        RECT 349.950 405.600 352.050 406.050 ;
        RECT 400.950 405.600 403.050 406.050 ;
        RECT 349.950 404.400 403.050 405.600 ;
        RECT 349.950 403.950 352.050 404.400 ;
        RECT 400.950 403.950 403.050 404.400 ;
        RECT 463.950 405.600 466.050 406.050 ;
        RECT 493.950 405.600 496.050 406.050 ;
        RECT 463.950 404.400 496.050 405.600 ;
        RECT 463.950 403.950 466.050 404.400 ;
        RECT 493.950 403.950 496.050 404.400 ;
        RECT 514.950 405.600 517.050 406.050 ;
        RECT 520.950 405.600 523.050 406.050 ;
        RECT 514.950 404.400 523.050 405.600 ;
        RECT 514.950 403.950 517.050 404.400 ;
        RECT 520.950 403.950 523.050 404.400 ;
        RECT 532.950 405.600 535.050 406.050 ;
        RECT 541.950 405.600 544.050 406.050 ;
        RECT 532.950 404.400 544.050 405.600 ;
        RECT 532.950 403.950 535.050 404.400 ;
        RECT 541.950 403.950 544.050 404.400 ;
        RECT 550.950 405.600 553.050 406.050 ;
        RECT 613.950 405.600 616.050 406.050 ;
        RECT 550.950 404.400 616.050 405.600 ;
        RECT 620.400 405.600 621.600 407.400 ;
        RECT 754.950 407.400 763.050 408.600 ;
        RECT 754.950 406.950 757.050 407.400 ;
        RECT 760.950 406.950 763.050 407.400 ;
        RECT 769.950 406.950 772.050 409.050 ;
        RECT 826.950 408.600 829.050 409.050 ;
        RECT 862.950 408.600 865.050 409.050 ;
        RECT 826.950 407.400 865.050 408.600 ;
        RECT 826.950 406.950 829.050 407.400 ;
        RECT 862.950 406.950 865.050 407.400 ;
        RECT 679.950 405.600 682.050 406.050 ;
        RECT 697.950 405.600 700.050 406.050 ;
        RECT 727.950 405.600 730.050 406.050 ;
        RECT 620.400 404.400 660.600 405.600 ;
        RECT 550.950 403.950 553.050 404.400 ;
        RECT 613.950 403.950 616.050 404.400 ;
        RECT 659.400 403.050 660.600 404.400 ;
        RECT 679.950 404.400 730.050 405.600 ;
        RECT 679.950 403.950 682.050 404.400 ;
        RECT 697.950 403.950 700.050 404.400 ;
        RECT 727.950 403.950 730.050 404.400 ;
        RECT 772.950 405.600 775.050 406.050 ;
        RECT 781.950 405.600 784.050 406.050 ;
        RECT 772.950 404.400 784.050 405.600 ;
        RECT 772.950 403.950 775.050 404.400 ;
        RECT 781.950 403.950 784.050 404.400 ;
        RECT 796.950 405.600 799.050 406.050 ;
        RECT 814.950 405.600 817.050 406.050 ;
        RECT 844.950 405.600 847.050 406.050 ;
        RECT 796.950 404.400 847.050 405.600 ;
        RECT 796.950 403.950 799.050 404.400 ;
        RECT 814.950 403.950 817.050 404.400 ;
        RECT 844.950 403.950 847.050 404.400 ;
        RECT 4.950 402.600 7.050 403.050 ;
        RECT 40.950 402.600 43.050 403.050 ;
        RECT 100.950 402.600 103.050 403.050 ;
        RECT 127.950 402.600 130.050 403.050 ;
        RECT 4.950 401.400 130.050 402.600 ;
        RECT 4.950 400.950 7.050 401.400 ;
        RECT 40.950 400.950 43.050 401.400 ;
        RECT 100.950 400.950 103.050 401.400 ;
        RECT 127.950 400.950 130.050 401.400 ;
        RECT 235.950 402.600 238.050 403.050 ;
        RECT 277.950 402.600 280.050 403.050 ;
        RECT 328.950 402.600 331.050 403.050 ;
        RECT 235.950 401.400 331.050 402.600 ;
        RECT 235.950 400.950 238.050 401.400 ;
        RECT 277.950 400.950 280.050 401.400 ;
        RECT 328.950 400.950 331.050 401.400 ;
        RECT 637.950 402.600 640.050 403.050 ;
        RECT 649.950 402.600 652.050 403.050 ;
        RECT 637.950 401.400 652.050 402.600 ;
        RECT 637.950 400.950 640.050 401.400 ;
        RECT 649.950 400.950 652.050 401.400 ;
        RECT 658.950 402.600 661.050 403.050 ;
        RECT 676.950 402.600 679.050 403.050 ;
        RECT 658.950 401.400 679.050 402.600 ;
        RECT 658.950 400.950 661.050 401.400 ;
        RECT 676.950 400.950 679.050 401.400 ;
        RECT 832.950 402.600 835.050 403.050 ;
        RECT 847.950 402.600 850.050 403.050 ;
        RECT 832.950 401.400 850.050 402.600 ;
        RECT 832.950 400.950 835.050 401.400 ;
        RECT 847.950 400.950 850.050 401.400 ;
        RECT 151.950 399.600 154.050 400.050 ;
        RECT 220.950 399.600 223.050 400.050 ;
        RECT 151.950 398.400 223.050 399.600 ;
        RECT 151.950 397.950 154.050 398.400 ;
        RECT 220.950 397.950 223.050 398.400 ;
        RECT 292.950 399.600 295.050 400.050 ;
        RECT 367.950 399.600 370.050 400.050 ;
        RECT 292.950 398.400 370.050 399.600 ;
        RECT 292.950 397.950 295.050 398.400 ;
        RECT 367.950 397.950 370.050 398.400 ;
        RECT 529.950 399.600 532.050 400.050 ;
        RECT 568.950 399.600 571.050 400.050 ;
        RECT 529.950 398.400 571.050 399.600 ;
        RECT 529.950 397.950 532.050 398.400 ;
        RECT 568.950 397.950 571.050 398.400 ;
        RECT 592.950 399.600 595.050 400.050 ;
        RECT 607.800 399.600 609.900 400.050 ;
        RECT 592.950 398.400 609.900 399.600 ;
        RECT 592.950 397.950 595.050 398.400 ;
        RECT 607.800 397.950 609.900 398.400 ;
        RECT 610.950 399.600 613.050 400.050 ;
        RECT 652.950 399.600 655.050 400.050 ;
        RECT 610.950 398.400 655.050 399.600 ;
        RECT 610.950 397.950 613.050 398.400 ;
        RECT 652.950 397.950 655.050 398.400 ;
        RECT 760.950 399.600 763.050 400.050 ;
        RECT 808.950 399.600 811.050 400.050 ;
        RECT 760.950 398.400 811.050 399.600 ;
        RECT 760.950 397.950 763.050 398.400 ;
        RECT 808.950 397.950 811.050 398.400 ;
        RECT 454.950 396.600 457.050 397.050 ;
        RECT 478.950 396.600 481.050 397.050 ;
        RECT 454.950 395.400 481.050 396.600 ;
        RECT 454.950 394.950 457.050 395.400 ;
        RECT 478.950 394.950 481.050 395.400 ;
        RECT 613.950 396.600 616.050 397.050 ;
        RECT 688.950 396.600 691.050 397.050 ;
        RECT 613.950 395.400 691.050 396.600 ;
        RECT 613.950 394.950 616.050 395.400 ;
        RECT 688.950 394.950 691.050 395.400 ;
        RECT 703.950 396.600 706.050 397.050 ;
        RECT 745.950 396.600 748.050 397.050 ;
        RECT 769.950 396.600 772.050 397.050 ;
        RECT 703.950 395.400 772.050 396.600 ;
        RECT 703.950 394.950 706.050 395.400 ;
        RECT 745.950 394.950 748.050 395.400 ;
        RECT 769.950 394.950 772.050 395.400 ;
        RECT 799.950 396.600 802.050 397.050 ;
        RECT 817.950 396.600 820.050 397.050 ;
        RECT 799.950 395.400 820.050 396.600 ;
        RECT 799.950 394.950 802.050 395.400 ;
        RECT 817.950 394.950 820.050 395.400 ;
        RECT 349.950 393.600 352.050 394.050 ;
        RECT 439.950 393.600 442.050 394.050 ;
        RECT 349.950 392.400 442.050 393.600 ;
        RECT 349.950 391.950 352.050 392.400 ;
        RECT 439.950 391.950 442.050 392.400 ;
        RECT 583.950 393.600 586.050 394.050 ;
        RECT 604.950 393.600 607.050 394.050 ;
        RECT 583.950 392.400 607.050 393.600 ;
        RECT 583.950 391.950 586.050 392.400 ;
        RECT 604.950 391.950 607.050 392.400 ;
        RECT 268.950 390.600 271.050 391.050 ;
        RECT 292.950 390.600 295.050 391.050 ;
        RECT 472.950 390.600 475.050 391.050 ;
        RECT 268.950 389.400 295.050 390.600 ;
        RECT 268.950 388.950 271.050 389.400 ;
        RECT 292.950 388.950 295.050 389.400 ;
        RECT 371.400 389.400 475.050 390.600 ;
        RECT 22.950 387.600 25.050 388.050 ;
        RECT 28.950 387.600 31.050 388.050 ;
        RECT 22.950 386.400 31.050 387.600 ;
        RECT 22.950 385.950 25.050 386.400 ;
        RECT 28.950 385.950 31.050 386.400 ;
        RECT 283.950 387.600 286.050 388.050 ;
        RECT 371.400 387.600 372.600 389.400 ;
        RECT 472.950 388.950 475.050 389.400 ;
        RECT 520.950 390.600 523.050 391.050 ;
        RECT 562.950 390.600 565.050 391.050 ;
        RECT 520.950 389.400 565.050 390.600 ;
        RECT 520.950 388.950 523.050 389.400 ;
        RECT 562.950 388.950 565.050 389.400 ;
        RECT 283.950 386.400 372.600 387.600 ;
        RECT 664.950 387.600 667.050 388.050 ;
        RECT 670.950 387.600 673.050 388.050 ;
        RECT 691.950 387.600 694.050 388.050 ;
        RECT 664.950 386.400 694.050 387.600 ;
        RECT 283.950 385.950 286.050 386.400 ;
        RECT 664.950 385.950 667.050 386.400 ;
        RECT 670.950 385.950 673.050 386.400 ;
        RECT 691.950 385.950 694.050 386.400 ;
        RECT 700.950 387.600 703.050 388.050 ;
        RECT 742.950 387.600 745.050 388.050 ;
        RECT 700.950 386.400 745.050 387.600 ;
        RECT 700.950 385.950 703.050 386.400 ;
        RECT 742.950 385.950 745.050 386.400 ;
        RECT 40.950 384.600 43.050 385.050 ;
        RECT 46.950 384.600 49.050 385.050 ;
        RECT 55.950 384.600 58.050 385.050 ;
        RECT 40.950 383.400 58.050 384.600 ;
        RECT 40.950 382.950 43.050 383.400 ;
        RECT 46.950 382.950 49.050 383.400 ;
        RECT 55.950 382.950 58.050 383.400 ;
        RECT 259.950 384.600 262.050 385.050 ;
        RECT 274.950 384.600 277.050 385.050 ;
        RECT 712.950 384.600 715.050 385.050 ;
        RECT 259.950 383.400 277.050 384.600 ;
        RECT 259.950 382.950 262.050 383.400 ;
        RECT 274.950 382.950 277.050 383.400 ;
        RECT 707.400 383.400 715.050 384.600 ;
        RECT 115.950 381.600 118.050 382.050 ;
        RECT 163.950 381.600 166.050 382.050 ;
        RECT 187.950 381.600 190.050 382.050 ;
        RECT 208.950 381.600 211.050 382.050 ;
        RECT 115.950 380.400 211.050 381.600 ;
        RECT 115.950 379.950 118.050 380.400 ;
        RECT 163.950 379.950 166.050 380.400 ;
        RECT 187.950 379.950 190.050 380.400 ;
        RECT 208.950 379.950 211.050 380.400 ;
        RECT 436.950 381.600 439.050 382.050 ;
        RECT 445.950 381.600 448.050 382.050 ;
        RECT 436.950 380.400 448.050 381.600 ;
        RECT 436.950 379.950 439.050 380.400 ;
        RECT 445.950 379.950 448.050 380.400 ;
        RECT 538.950 381.600 541.050 382.050 ;
        RECT 547.950 381.600 550.050 382.050 ;
        RECT 538.950 380.400 550.050 381.600 ;
        RECT 538.950 379.950 541.050 380.400 ;
        RECT 547.950 379.950 550.050 380.400 ;
        RECT 586.950 381.600 589.050 382.050 ;
        RECT 592.950 381.600 595.050 382.050 ;
        RECT 586.950 380.400 595.050 381.600 ;
        RECT 586.950 379.950 589.050 380.400 ;
        RECT 592.950 379.950 595.050 380.400 ;
        RECT 691.950 381.600 694.050 382.050 ;
        RECT 707.400 381.600 708.600 383.400 ;
        RECT 712.950 382.950 715.050 383.400 ;
        RECT 718.950 384.600 721.050 385.050 ;
        RECT 736.950 384.600 739.050 385.050 ;
        RECT 718.950 383.400 739.050 384.600 ;
        RECT 718.950 382.950 721.050 383.400 ;
        RECT 736.950 382.950 739.050 383.400 ;
        RECT 691.950 380.400 708.600 381.600 ;
        RECT 709.950 381.600 712.050 382.050 ;
        RECT 730.950 381.600 733.050 382.050 ;
        RECT 709.950 380.400 733.050 381.600 ;
        RECT 691.950 379.950 694.050 380.400 ;
        RECT 709.950 379.950 712.050 380.400 ;
        RECT 730.950 379.950 733.050 380.400 ;
        RECT 832.950 381.600 835.050 382.050 ;
        RECT 862.950 381.600 865.050 382.050 ;
        RECT 832.950 380.400 865.050 381.600 ;
        RECT 832.950 379.950 835.050 380.400 ;
        RECT 862.950 379.950 865.050 380.400 ;
        RECT 313.950 378.600 316.050 379.050 ;
        RECT 391.950 378.600 394.050 379.050 ;
        RECT 313.950 377.400 394.050 378.600 ;
        RECT 313.950 376.950 316.050 377.400 ;
        RECT 391.950 376.950 394.050 377.400 ;
        RECT 397.950 378.600 400.050 379.050 ;
        RECT 403.950 378.600 406.050 379.050 ;
        RECT 412.950 378.600 415.050 379.050 ;
        RECT 397.950 377.400 415.050 378.600 ;
        RECT 397.950 376.950 400.050 377.400 ;
        RECT 403.950 376.950 406.050 377.400 ;
        RECT 412.950 376.950 415.050 377.400 ;
        RECT 526.950 378.600 529.050 379.050 ;
        RECT 550.950 378.600 553.050 379.050 ;
        RECT 526.950 377.400 553.050 378.600 ;
        RECT 526.950 376.950 529.050 377.400 ;
        RECT 550.950 376.950 553.050 377.400 ;
        RECT 625.950 378.600 628.050 379.050 ;
        RECT 643.950 378.600 646.050 379.050 ;
        RECT 625.950 377.400 646.050 378.600 ;
        RECT 625.950 376.950 628.050 377.400 ;
        RECT 643.950 376.950 646.050 377.400 ;
        RECT 748.950 378.600 751.050 379.050 ;
        RECT 757.950 378.600 760.050 379.050 ;
        RECT 748.950 377.400 760.050 378.600 ;
        RECT 748.950 376.950 751.050 377.400 ;
        RECT 757.950 376.950 760.050 377.400 ;
        RECT 763.950 378.600 766.050 379.050 ;
        RECT 790.800 378.600 792.900 379.050 ;
        RECT 763.950 377.400 792.900 378.600 ;
        RECT 763.950 376.950 766.050 377.400 ;
        RECT 790.800 376.950 792.900 377.400 ;
        RECT 10.950 375.600 13.050 376.050 ;
        RECT 19.950 375.600 22.050 376.050 ;
        RECT 10.950 374.400 22.050 375.600 ;
        RECT 10.950 373.950 13.050 374.400 ;
        RECT 19.950 373.950 22.050 374.400 ;
        RECT 67.950 375.600 70.050 376.050 ;
        RECT 73.950 375.600 76.050 376.050 ;
        RECT 67.950 374.400 76.050 375.600 ;
        RECT 67.950 373.950 70.050 374.400 ;
        RECT 73.950 373.950 76.050 374.400 ;
        RECT 82.950 375.600 85.050 376.050 ;
        RECT 100.950 375.600 103.050 376.050 ;
        RECT 106.950 375.600 109.050 376.050 ;
        RECT 82.950 374.400 109.050 375.600 ;
        RECT 82.950 373.950 85.050 374.400 ;
        RECT 100.950 373.950 103.050 374.400 ;
        RECT 106.950 373.950 109.050 374.400 ;
        RECT 259.950 373.950 262.050 376.050 ;
        RECT 445.950 375.600 448.050 376.050 ;
        RECT 502.950 375.600 505.050 376.050 ;
        RECT 520.950 375.600 523.050 376.050 ;
        RECT 445.950 374.400 523.050 375.600 ;
        RECT 445.950 373.950 448.050 374.400 ;
        RECT 502.950 373.950 505.050 374.400 ;
        RECT 520.950 373.950 523.050 374.400 ;
        RECT 562.950 375.600 565.050 376.050 ;
        RECT 583.950 375.600 586.050 376.050 ;
        RECT 562.950 374.400 586.050 375.600 ;
        RECT 562.950 373.950 565.050 374.400 ;
        RECT 583.950 373.950 586.050 374.400 ;
        RECT 676.950 375.600 681.000 376.050 ;
        RECT 685.950 375.600 688.050 376.050 ;
        RECT 712.950 375.600 715.050 376.050 ;
        RECT 676.950 373.950 681.600 375.600 ;
        RECT 685.950 374.400 715.050 375.600 ;
        RECT 685.950 373.950 688.050 374.400 ;
        RECT 712.950 373.950 715.050 374.400 ;
        RECT 760.950 373.950 763.050 376.050 ;
        RECT 826.950 373.950 829.050 376.050 ;
        RECT 10.950 371.100 13.050 373.200 ;
        RECT 31.950 372.600 34.050 373.050 ;
        RECT 37.950 372.600 40.050 373.200 ;
        RECT 31.950 371.400 40.050 372.600 ;
        RECT 11.400 364.050 12.600 371.100 ;
        RECT 31.950 370.950 34.050 371.400 ;
        RECT 37.950 371.100 40.050 371.400 ;
        RECT 64.950 372.600 67.050 373.200 ;
        RECT 91.950 372.600 94.050 373.050 ;
        RECT 64.950 371.400 94.050 372.600 ;
        RECT 64.950 371.100 67.050 371.400 ;
        RECT 91.950 370.950 94.050 371.400 ;
        RECT 121.950 371.100 124.050 373.200 ;
        RECT 136.950 372.750 139.050 373.200 ;
        RECT 142.950 372.750 145.050 373.200 ;
        RECT 136.950 371.550 145.050 372.750 ;
        RECT 136.950 371.100 139.050 371.550 ;
        RECT 142.950 371.100 145.050 371.550 ;
        RECT 172.950 372.750 175.050 373.200 ;
        RECT 178.950 372.750 181.050 373.200 ;
        RECT 172.950 371.550 181.050 372.750 ;
        RECT 172.950 371.100 175.050 371.550 ;
        RECT 178.950 371.100 181.050 371.550 ;
        RECT 193.950 371.100 196.050 373.200 ;
        RECT 214.950 372.750 217.050 373.200 ;
        RECT 223.800 372.750 225.900 373.200 ;
        RECT 214.950 371.550 225.900 372.750 ;
        RECT 214.950 371.100 217.050 371.550 ;
        RECT 223.800 371.100 225.900 371.550 ;
        RECT 226.950 371.100 229.050 373.200 ;
        RECT 13.950 366.600 16.050 366.900 ;
        RECT 19.950 366.600 22.050 366.900 ;
        RECT 13.950 366.450 22.050 366.600 ;
        RECT 28.950 366.450 31.050 366.900 ;
        RECT 13.950 365.400 31.050 366.450 ;
        RECT 13.950 364.800 16.050 365.400 ;
        RECT 19.950 365.250 31.050 365.400 ;
        RECT 19.950 364.800 22.050 365.250 ;
        RECT 28.950 364.800 31.050 365.250 ;
        RECT 82.950 366.600 85.050 366.900 ;
        RECT 97.950 366.600 100.050 366.900 ;
        RECT 82.950 365.400 100.050 366.600 ;
        RECT 82.950 364.800 85.050 365.400 ;
        RECT 97.950 364.800 100.050 365.400 ;
        RECT 106.950 366.450 109.050 366.900 ;
        RECT 112.950 366.450 115.050 366.900 ;
        RECT 106.950 365.250 115.050 366.450 ;
        RECT 122.400 366.600 123.600 371.100 ;
        RECT 194.400 369.600 195.600 371.100 ;
        RECT 220.950 369.600 223.050 370.050 ;
        RECT 194.400 368.400 223.050 369.600 ;
        RECT 220.950 367.950 223.050 368.400 ;
        RECT 145.950 366.600 148.050 367.050 ;
        RECT 122.400 365.400 148.050 366.600 ;
        RECT 106.950 364.800 109.050 365.250 ;
        RECT 112.950 364.800 115.050 365.250 ;
        RECT 145.950 364.950 148.050 365.400 ;
        RECT 154.950 366.450 157.050 366.900 ;
        RECT 160.950 366.600 163.050 366.900 ;
        RECT 169.950 366.600 172.050 366.900 ;
        RECT 160.950 366.450 172.050 366.600 ;
        RECT 154.950 365.400 172.050 366.450 ;
        RECT 154.950 365.250 163.050 365.400 ;
        RECT 154.950 364.800 157.050 365.250 ;
        RECT 160.950 364.800 163.050 365.250 ;
        RECT 169.950 364.800 172.050 365.400 ;
        RECT 178.950 366.600 181.050 367.050 ;
        RECT 184.950 366.600 187.050 366.900 ;
        RECT 178.950 365.400 187.050 366.600 ;
        RECT 178.950 364.950 181.050 365.400 ;
        RECT 184.950 364.800 187.050 365.400 ;
        RECT 196.950 366.600 199.050 366.900 ;
        RECT 211.950 366.600 214.050 366.900 ;
        RECT 196.950 365.400 214.050 366.600 ;
        RECT 196.950 364.800 199.050 365.400 ;
        RECT 211.950 364.800 214.050 365.400 ;
        RECT 10.950 361.950 13.050 364.050 ;
        RECT 214.950 363.600 217.050 364.050 ;
        RECT 220.950 363.600 223.050 364.050 ;
        RECT 214.950 362.400 223.050 363.600 ;
        RECT 227.400 363.600 228.600 371.100 ;
        RECT 260.400 366.900 261.600 373.950 ;
        RECT 262.950 372.600 265.050 373.200 ;
        RECT 277.950 372.600 280.050 373.200 ;
        RECT 262.950 371.400 280.050 372.600 ;
        RECT 262.950 371.100 265.050 371.400 ;
        RECT 277.950 371.100 280.050 371.400 ;
        RECT 319.950 372.750 322.050 373.200 ;
        RECT 325.950 372.750 328.050 373.200 ;
        RECT 319.950 371.550 328.050 372.750 ;
        RECT 319.950 371.100 322.050 371.550 ;
        RECT 325.950 371.100 328.050 371.550 ;
        RECT 334.950 371.100 337.050 373.200 ;
        RECT 352.950 372.750 355.050 373.200 ;
        RECT 358.950 372.750 361.050 373.200 ;
        RECT 352.950 371.550 361.050 372.750 ;
        RECT 352.950 371.100 355.050 371.550 ;
        RECT 358.950 371.100 361.050 371.550 ;
        RECT 376.950 372.750 379.050 373.200 ;
        RECT 382.950 372.750 385.050 373.200 ;
        RECT 376.950 371.550 385.050 372.750 ;
        RECT 388.950 372.600 391.050 373.200 ;
        RECT 376.950 371.100 379.050 371.550 ;
        RECT 382.950 371.100 385.050 371.550 ;
        RECT 386.400 371.400 391.050 372.600 ;
        RECT 335.400 369.600 336.600 371.100 ;
        RECT 386.400 369.600 387.600 371.400 ;
        RECT 388.950 371.100 391.050 371.400 ;
        RECT 439.950 371.100 442.050 373.200 ;
        RECT 463.950 372.600 466.050 373.200 ;
        RECT 469.950 372.600 472.050 373.050 ;
        RECT 463.950 371.400 472.050 372.600 ;
        RECT 463.950 371.100 466.050 371.400 ;
        RECT 440.400 369.600 441.600 371.100 ;
        RECT 469.950 370.950 472.050 371.400 ;
        RECT 508.950 372.750 511.050 373.200 ;
        RECT 514.950 372.750 517.050 373.200 ;
        RECT 508.950 371.550 517.050 372.750 ;
        RECT 508.950 371.100 511.050 371.550 ;
        RECT 514.950 371.100 517.050 371.550 ;
        RECT 526.950 370.950 529.050 373.050 ;
        RECT 571.950 372.750 574.050 373.200 ;
        RECT 577.950 372.750 580.050 373.200 ;
        RECT 571.950 371.550 580.050 372.750 ;
        RECT 588.000 372.600 592.050 373.050 ;
        RECT 571.950 371.100 574.050 371.550 ;
        RECT 577.950 371.100 580.050 371.550 ;
        RECT 587.400 370.950 592.050 372.600 ;
        RECT 601.950 372.600 604.050 373.200 ;
        RECT 607.950 372.600 610.050 373.050 ;
        RECT 601.950 371.400 610.050 372.600 ;
        RECT 601.950 371.100 604.050 371.400 ;
        RECT 607.950 370.950 610.050 371.400 ;
        RECT 637.950 371.100 640.050 373.200 ;
        RECT 335.400 368.400 387.600 369.600 ;
        RECT 431.400 368.400 441.600 369.600 ;
        RECT 452.400 368.400 495.600 369.600 ;
        RECT 259.950 364.800 262.050 366.900 ;
        RECT 295.950 366.450 298.050 366.900 ;
        RECT 301.950 366.450 304.050 366.900 ;
        RECT 295.950 365.250 304.050 366.450 ;
        RECT 295.950 364.800 298.050 365.250 ;
        RECT 301.950 364.800 304.050 365.250 ;
        RECT 325.950 366.600 328.050 367.050 ;
        RECT 331.950 366.600 334.050 366.900 ;
        RECT 340.950 366.600 343.050 366.900 ;
        RECT 325.950 365.400 343.050 366.600 ;
        RECT 325.950 364.950 328.050 365.400 ;
        RECT 331.950 364.800 334.050 365.400 ;
        RECT 340.950 364.800 343.050 365.400 ;
        RECT 232.950 363.600 235.050 364.050 ;
        RECT 227.400 362.400 235.050 363.600 ;
        RECT 214.950 361.950 217.050 362.400 ;
        RECT 220.950 361.950 223.050 362.400 ;
        RECT 232.950 361.950 235.050 362.400 ;
        RECT 286.950 363.600 289.050 364.050 ;
        RECT 316.950 363.600 319.050 364.050 ;
        RECT 286.950 362.400 319.050 363.600 ;
        RECT 286.950 361.950 289.050 362.400 ;
        RECT 316.950 361.950 319.050 362.400 ;
        RECT 334.950 363.600 337.050 364.050 ;
        RECT 344.400 363.600 345.600 368.400 ;
        RECT 352.950 366.600 355.050 367.050 ;
        RECT 385.950 366.600 388.050 366.900 ;
        RECT 352.950 365.400 388.050 366.600 ;
        RECT 352.950 364.950 355.050 365.400 ;
        RECT 385.950 364.800 388.050 365.400 ;
        RECT 391.950 366.450 394.050 366.900 ;
        RECT 397.950 366.450 400.050 366.900 ;
        RECT 391.950 365.250 400.050 366.450 ;
        RECT 391.950 364.800 394.050 365.250 ;
        RECT 397.950 364.800 400.050 365.250 ;
        RECT 424.950 366.600 427.050 366.900 ;
        RECT 431.400 366.600 432.600 368.400 ;
        RECT 424.950 365.400 432.600 366.600 ;
        RECT 433.950 366.600 436.050 367.050 ;
        RECT 452.400 366.600 453.600 368.400 ;
        RECT 433.950 365.400 453.600 366.600 ;
        RECT 484.950 366.600 487.050 367.050 ;
        RECT 490.950 366.600 493.050 367.050 ;
        RECT 484.950 365.400 493.050 366.600 ;
        RECT 494.400 366.600 495.600 368.400 ;
        RECT 523.950 366.600 526.050 366.900 ;
        RECT 527.400 366.600 528.600 370.950 ;
        RECT 587.400 369.600 588.600 370.950 ;
        RECT 584.400 368.400 588.600 369.600 ;
        RECT 494.400 365.400 528.600 366.600 ;
        RECT 559.950 366.600 562.050 366.900 ;
        RECT 571.800 366.600 573.900 367.050 ;
        RECT 559.950 365.400 573.900 366.600 ;
        RECT 424.950 364.800 427.050 365.400 ;
        RECT 433.950 364.950 436.050 365.400 ;
        RECT 484.950 364.950 487.050 365.400 ;
        RECT 490.950 364.950 493.050 365.400 ;
        RECT 523.950 364.800 526.050 365.400 ;
        RECT 559.950 364.800 562.050 365.400 ;
        RECT 571.800 364.950 573.900 365.400 ;
        RECT 574.950 366.600 577.050 367.050 ;
        RECT 584.400 366.600 585.600 368.400 ;
        RECT 574.950 365.400 585.600 366.600 ;
        RECT 589.950 366.600 592.050 367.050 ;
        RECT 589.950 365.400 630.600 366.600 ;
        RECT 574.950 364.950 577.050 365.400 ;
        RECT 589.950 364.950 592.050 365.400 ;
        RECT 334.950 362.400 345.600 363.600 ;
        RECT 442.950 363.600 445.050 364.050 ;
        RECT 469.950 363.600 472.050 364.050 ;
        RECT 442.950 362.400 472.050 363.600 ;
        RECT 334.950 361.950 337.050 362.400 ;
        RECT 442.950 361.950 445.050 362.400 ;
        RECT 469.950 361.950 472.050 362.400 ;
        RECT 499.950 363.600 502.050 364.050 ;
        RECT 508.950 363.600 511.050 364.050 ;
        RECT 499.950 362.400 511.050 363.600 ;
        RECT 499.950 361.950 502.050 362.400 ;
        RECT 508.950 361.950 511.050 362.400 ;
        RECT 580.950 363.600 583.050 364.050 ;
        RECT 607.950 363.600 610.050 364.050 ;
        RECT 580.950 362.400 610.050 363.600 ;
        RECT 629.400 363.600 630.600 365.400 ;
        RECT 638.400 364.050 639.600 371.100 ;
        RECT 652.950 369.600 655.050 373.050 ;
        RECT 658.950 371.100 661.050 373.200 ;
        RECT 659.400 369.600 660.600 371.100 ;
        RECT 652.950 369.000 660.600 369.600 ;
        RECT 653.400 368.400 660.600 369.000 ;
        RECT 629.400 362.400 636.600 363.600 ;
        RECT 580.950 361.950 583.050 362.400 ;
        RECT 607.950 361.950 610.050 362.400 ;
        RECT 142.950 360.600 145.050 361.050 ;
        RECT 190.950 360.600 193.050 361.050 ;
        RECT 142.950 359.400 193.050 360.600 ;
        RECT 142.950 358.950 145.050 359.400 ;
        RECT 190.950 358.950 193.050 359.400 ;
        RECT 202.950 360.600 205.050 361.050 ;
        RECT 235.950 360.600 238.050 361.050 ;
        RECT 202.950 359.400 238.050 360.600 ;
        RECT 202.950 358.950 205.050 359.400 ;
        RECT 235.950 358.950 238.050 359.400 ;
        RECT 376.950 360.600 379.050 361.050 ;
        RECT 406.950 360.600 409.050 361.050 ;
        RECT 376.950 359.400 409.050 360.600 ;
        RECT 376.950 358.950 379.050 359.400 ;
        RECT 406.950 358.950 409.050 359.400 ;
        RECT 505.950 360.600 508.050 361.050 ;
        RECT 517.950 360.600 520.050 361.050 ;
        RECT 505.950 359.400 520.050 360.600 ;
        RECT 505.950 358.950 508.050 359.400 ;
        RECT 517.950 358.950 520.050 359.400 ;
        RECT 526.950 360.600 529.050 361.050 ;
        RECT 574.950 360.600 577.050 361.050 ;
        RECT 526.950 359.400 577.050 360.600 ;
        RECT 635.400 360.600 636.600 362.400 ;
        RECT 637.950 361.950 640.050 364.050 ;
        RECT 676.950 363.600 679.050 364.050 ;
        RECT 671.400 362.400 679.050 363.600 ;
        RECT 680.400 363.600 681.600 373.950 ;
        RECT 691.950 370.950 694.050 373.050 ;
        RECT 697.950 372.600 700.050 373.200 ;
        RECT 706.950 372.600 709.050 373.050 ;
        RECT 736.950 372.600 739.050 373.200 ;
        RECT 757.950 372.600 760.050 373.200 ;
        RECT 697.950 371.400 709.050 372.600 ;
        RECT 697.950 371.100 700.050 371.400 ;
        RECT 706.950 370.950 709.050 371.400 ;
        RECT 728.400 371.400 760.050 372.600 ;
        RECT 682.950 366.600 685.050 366.900 ;
        RECT 692.400 366.600 693.600 370.950 ;
        RECT 694.950 366.600 697.050 366.900 ;
        RECT 682.950 365.400 697.050 366.600 ;
        RECT 682.950 364.800 685.050 365.400 ;
        RECT 694.950 364.800 697.050 365.400 ;
        RECT 715.950 366.600 718.050 366.900 ;
        RECT 728.400 366.600 729.600 371.400 ;
        RECT 736.950 371.100 739.050 371.400 ;
        RECT 757.950 371.100 760.050 371.400 ;
        RECT 761.400 366.900 762.600 373.950 ;
        RECT 781.950 372.600 784.050 373.200 ;
        RECT 767.400 371.400 784.050 372.600 ;
        RECT 767.400 366.900 768.600 371.400 ;
        RECT 781.950 371.100 784.050 371.400 ;
        RECT 790.950 372.750 793.050 373.200 ;
        RECT 796.950 372.750 799.050 373.200 ;
        RECT 790.950 371.550 799.050 372.750 ;
        RECT 790.950 371.100 793.050 371.550 ;
        RECT 796.950 371.100 799.050 371.550 ;
        RECT 814.950 372.600 817.050 373.050 ;
        RECT 820.950 372.600 823.050 373.050 ;
        RECT 814.950 371.400 823.050 372.600 ;
        RECT 814.950 370.950 817.050 371.400 ;
        RECT 820.950 370.950 823.050 371.400 ;
        RECT 827.400 369.600 828.600 373.950 ;
        RECT 829.950 372.750 832.050 373.200 ;
        RECT 838.950 372.750 841.050 373.200 ;
        RECT 829.950 371.550 841.050 372.750 ;
        RECT 829.950 371.100 832.050 371.550 ;
        RECT 838.950 371.100 841.050 371.550 ;
        RECT 844.950 372.600 847.050 373.200 ;
        RECT 859.950 372.600 862.050 373.200 ;
        RECT 844.950 371.400 862.050 372.600 ;
        RECT 844.950 371.100 847.050 371.400 ;
        RECT 859.950 371.100 862.050 371.400 ;
        RECT 865.950 370.950 868.050 373.050 ;
        RECT 824.400 368.400 828.600 369.600 ;
        RECT 824.400 366.900 825.600 368.400 ;
        RECT 715.950 365.400 729.600 366.600 ;
        RECT 715.950 364.800 718.050 365.400 ;
        RECT 760.950 364.800 763.050 366.900 ;
        RECT 766.950 364.800 769.050 366.900 ;
        RECT 778.950 366.600 781.050 366.900 ;
        RECT 811.950 366.600 814.050 366.900 ;
        RECT 778.950 365.400 814.050 366.600 ;
        RECT 778.950 364.800 781.050 365.400 ;
        RECT 811.950 364.800 814.050 365.400 ;
        RECT 823.950 364.800 826.050 366.900 ;
        RECT 832.950 366.450 835.050 366.900 ;
        RECT 847.950 366.600 850.050 366.900 ;
        RECT 853.800 366.600 855.900 367.050 ;
        RECT 847.950 366.450 855.900 366.600 ;
        RECT 832.950 365.400 855.900 366.450 ;
        RECT 832.950 365.250 850.050 365.400 ;
        RECT 832.950 364.800 835.050 365.250 ;
        RECT 847.950 364.800 850.050 365.250 ;
        RECT 853.800 364.950 855.900 365.400 ;
        RECT 856.950 366.600 859.050 367.050 ;
        RECT 866.400 366.600 867.600 370.950 ;
        RECT 856.950 365.400 867.600 366.600 ;
        RECT 856.950 364.950 859.050 365.400 ;
        RECT 688.950 363.600 691.050 364.050 ;
        RECT 680.400 362.400 691.050 363.600 ;
        RECT 655.950 360.600 658.050 361.050 ;
        RECT 671.400 360.600 672.600 362.400 ;
        RECT 676.950 361.950 679.050 362.400 ;
        RECT 688.950 361.950 691.050 362.400 ;
        RECT 709.950 363.600 712.050 364.050 ;
        RECT 724.950 363.600 727.050 364.050 ;
        RECT 709.950 362.400 727.050 363.600 ;
        RECT 709.950 361.950 712.050 362.400 ;
        RECT 724.950 361.950 727.050 362.400 ;
        RECT 745.950 363.600 748.050 364.050 ;
        RECT 757.950 363.600 760.050 364.050 ;
        RECT 745.950 362.400 760.050 363.600 ;
        RECT 745.950 361.950 748.050 362.400 ;
        RECT 757.950 361.950 760.050 362.400 ;
        RECT 787.950 363.600 790.050 364.050 ;
        RECT 793.950 363.600 796.050 363.900 ;
        RECT 787.950 362.400 796.050 363.600 ;
        RECT 787.950 361.950 790.050 362.400 ;
        RECT 793.950 361.800 796.050 362.400 ;
        RECT 685.950 360.600 688.050 361.050 ;
        RECT 635.400 359.400 672.600 360.600 ;
        RECT 674.400 359.400 688.050 360.600 ;
        RECT 526.950 358.950 529.050 359.400 ;
        RECT 574.950 358.950 577.050 359.400 ;
        RECT 655.950 358.950 658.050 359.400 ;
        RECT 91.950 357.600 94.050 358.050 ;
        RECT 118.950 357.600 121.050 358.050 ;
        RECT 91.950 356.400 121.050 357.600 ;
        RECT 91.950 355.950 94.050 356.400 ;
        RECT 118.950 355.950 121.050 356.400 ;
        RECT 145.950 357.600 148.050 358.050 ;
        RECT 187.950 357.600 190.050 358.050 ;
        RECT 145.950 356.400 190.050 357.600 ;
        RECT 145.950 355.950 148.050 356.400 ;
        RECT 187.950 355.950 190.050 356.400 ;
        RECT 193.950 357.600 196.050 358.050 ;
        RECT 310.950 357.600 313.050 358.050 ;
        RECT 193.950 356.400 313.050 357.600 ;
        RECT 193.950 355.950 196.050 356.400 ;
        RECT 310.950 355.950 313.050 356.400 ;
        RECT 325.950 357.600 328.050 358.050 ;
        RECT 349.950 357.600 352.050 358.050 ;
        RECT 355.950 357.600 358.050 358.050 ;
        RECT 325.950 356.400 358.050 357.600 ;
        RECT 325.950 355.950 328.050 356.400 ;
        RECT 349.950 355.950 352.050 356.400 ;
        RECT 355.950 355.950 358.050 356.400 ;
        RECT 511.950 357.600 514.050 358.050 ;
        RECT 532.950 357.600 535.050 358.050 ;
        RECT 511.950 356.400 535.050 357.600 ;
        RECT 511.950 355.950 514.050 356.400 ;
        RECT 532.950 355.950 535.050 356.400 ;
        RECT 622.950 357.600 625.050 358.050 ;
        RECT 652.950 357.600 655.050 358.050 ;
        RECT 674.400 357.600 675.600 359.400 ;
        RECT 685.950 358.950 688.050 359.400 ;
        RECT 733.950 360.600 736.050 361.050 ;
        RECT 769.950 360.600 772.050 361.050 ;
        RECT 733.950 359.400 772.050 360.600 ;
        RECT 733.950 358.950 736.050 359.400 ;
        RECT 769.950 358.950 772.050 359.400 ;
        RECT 814.950 360.600 817.050 361.050 ;
        RECT 838.950 360.600 841.050 361.050 ;
        RECT 814.950 359.400 841.050 360.600 ;
        RECT 814.950 358.950 817.050 359.400 ;
        RECT 838.950 358.950 841.050 359.400 ;
        RECT 703.800 357.600 705.900 358.050 ;
        RECT 622.950 356.400 675.600 357.600 ;
        RECT 683.400 356.400 705.900 357.600 ;
        RECT 622.950 355.950 625.050 356.400 ;
        RECT 652.950 355.950 655.050 356.400 ;
        RECT 223.950 354.600 226.050 355.050 ;
        RECT 274.950 354.600 277.050 355.050 ;
        RECT 283.950 354.600 286.050 355.050 ;
        RECT 223.950 353.400 286.050 354.600 ;
        RECT 223.950 352.950 226.050 353.400 ;
        RECT 274.950 352.950 277.050 353.400 ;
        RECT 283.950 352.950 286.050 353.400 ;
        RECT 313.950 354.600 316.050 355.050 ;
        RECT 388.950 354.600 391.050 355.050 ;
        RECT 313.950 353.400 391.050 354.600 ;
        RECT 313.950 352.950 316.050 353.400 ;
        RECT 388.950 352.950 391.050 353.400 ;
        RECT 661.950 354.600 664.050 355.050 ;
        RECT 683.400 354.600 684.600 356.400 ;
        RECT 703.800 355.950 705.900 356.400 ;
        RECT 706.950 357.600 709.050 358.050 ;
        RECT 778.950 357.600 781.050 358.050 ;
        RECT 706.950 356.400 781.050 357.600 ;
        RECT 706.950 355.950 709.050 356.400 ;
        RECT 778.950 355.950 781.050 356.400 ;
        RECT 787.950 357.600 790.050 358.050 ;
        RECT 799.950 357.600 802.050 358.050 ;
        RECT 787.950 356.400 802.050 357.600 ;
        RECT 787.950 355.950 790.050 356.400 ;
        RECT 799.950 355.950 802.050 356.400 ;
        RECT 661.950 353.400 684.600 354.600 ;
        RECT 691.950 354.600 694.050 355.050 ;
        RECT 700.950 354.600 703.050 355.050 ;
        RECT 691.950 353.400 703.050 354.600 ;
        RECT 661.950 352.950 664.050 353.400 ;
        RECT 691.950 352.950 694.050 353.400 ;
        RECT 700.950 352.950 703.050 353.400 ;
        RECT 826.950 354.600 829.050 355.050 ;
        RECT 835.950 354.600 838.050 355.050 ;
        RECT 826.950 353.400 838.050 354.600 ;
        RECT 826.950 352.950 829.050 353.400 ;
        RECT 835.950 352.950 838.050 353.400 ;
        RECT 841.950 354.600 844.050 355.050 ;
        RECT 850.950 354.600 853.050 355.050 ;
        RECT 841.950 353.400 853.050 354.600 ;
        RECT 841.950 352.950 844.050 353.400 ;
        RECT 850.950 352.950 853.050 353.400 ;
        RECT 160.950 351.600 163.050 352.050 ;
        RECT 250.950 351.600 253.050 352.050 ;
        RECT 160.950 350.400 253.050 351.600 ;
        RECT 160.950 349.950 163.050 350.400 ;
        RECT 250.950 349.950 253.050 350.400 ;
        RECT 349.950 351.600 352.050 352.050 ;
        RECT 430.950 351.600 433.050 352.050 ;
        RECT 448.950 351.600 451.050 352.050 ;
        RECT 349.950 350.400 451.050 351.600 ;
        RECT 349.950 349.950 352.050 350.400 ;
        RECT 430.950 349.950 433.050 350.400 ;
        RECT 448.950 349.950 451.050 350.400 ;
        RECT 469.950 351.600 472.050 352.050 ;
        RECT 481.950 351.600 484.050 352.050 ;
        RECT 469.950 350.400 484.050 351.600 ;
        RECT 469.950 349.950 472.050 350.400 ;
        RECT 310.950 348.600 313.050 349.050 ;
        RECT 340.950 348.600 343.050 349.050 ;
        RECT 310.950 347.400 343.050 348.600 ;
        RECT 481.950 348.600 484.050 350.400 ;
        RECT 487.950 351.600 490.050 352.050 ;
        RECT 562.950 351.600 565.050 352.050 ;
        RECT 487.950 350.400 565.050 351.600 ;
        RECT 487.950 349.950 490.050 350.400 ;
        RECT 562.950 349.950 565.050 350.400 ;
        RECT 685.950 351.600 690.000 352.050 ;
        RECT 700.950 351.600 703.050 351.900 ;
        RECT 739.950 351.600 742.050 352.050 ;
        RECT 754.950 351.600 757.050 352.050 ;
        RECT 685.950 349.950 690.600 351.600 ;
        RECT 526.950 348.600 529.050 349.050 ;
        RECT 481.950 348.000 529.050 348.600 ;
        RECT 482.400 347.400 529.050 348.000 ;
        RECT 689.400 348.600 690.600 349.950 ;
        RECT 700.950 350.400 757.050 351.600 ;
        RECT 700.950 349.800 703.050 350.400 ;
        RECT 739.950 349.950 742.050 350.400 ;
        RECT 754.950 349.950 757.050 350.400 ;
        RECT 772.950 351.600 775.050 352.050 ;
        RECT 778.950 351.600 781.050 352.050 ;
        RECT 772.950 350.400 781.050 351.600 ;
        RECT 772.950 349.950 775.050 350.400 ;
        RECT 778.950 349.950 781.050 350.400 ;
        RECT 799.950 351.600 802.050 352.050 ;
        RECT 814.950 351.600 817.050 352.050 ;
        RECT 823.950 351.600 826.050 352.050 ;
        RECT 799.950 350.400 826.050 351.600 ;
        RECT 799.950 349.950 802.050 350.400 ;
        RECT 814.950 349.950 817.050 350.400 ;
        RECT 823.950 349.950 826.050 350.400 ;
        RECT 733.950 348.600 736.050 349.050 ;
        RECT 689.400 347.400 736.050 348.600 ;
        RECT 310.950 346.950 313.050 347.400 ;
        RECT 340.950 346.950 343.050 347.400 ;
        RECT 526.950 346.950 529.050 347.400 ;
        RECT 733.950 346.950 736.050 347.400 ;
        RECT 811.950 348.600 814.050 349.050 ;
        RECT 829.950 348.600 832.050 349.050 ;
        RECT 811.950 347.400 832.050 348.600 ;
        RECT 811.950 346.950 814.050 347.400 ;
        RECT 829.950 346.950 832.050 347.400 ;
        RECT 835.950 348.600 838.050 349.050 ;
        RECT 841.950 348.600 844.050 349.050 ;
        RECT 835.950 347.400 844.050 348.600 ;
        RECT 835.950 346.950 838.050 347.400 ;
        RECT 841.950 346.950 844.050 347.400 ;
        RECT 16.950 345.600 19.050 346.050 ;
        RECT 31.950 345.600 34.050 346.050 ;
        RECT 16.950 344.400 34.050 345.600 ;
        RECT 16.950 343.950 19.050 344.400 ;
        RECT 31.950 343.950 34.050 344.400 ;
        RECT 91.950 345.600 94.050 346.050 ;
        RECT 151.950 345.600 154.050 346.050 ;
        RECT 163.950 345.600 166.050 346.050 ;
        RECT 91.950 344.400 166.050 345.600 ;
        RECT 91.950 343.950 94.050 344.400 ;
        RECT 151.950 343.950 154.050 344.400 ;
        RECT 163.950 343.950 166.050 344.400 ;
        RECT 220.950 345.600 223.050 346.050 ;
        RECT 235.950 345.600 238.050 346.050 ;
        RECT 244.950 345.600 247.050 346.050 ;
        RECT 262.950 345.600 265.050 346.050 ;
        RECT 220.950 344.400 265.050 345.600 ;
        RECT 220.950 343.950 223.050 344.400 ;
        RECT 235.950 343.950 238.050 344.400 ;
        RECT 244.950 343.950 247.050 344.400 ;
        RECT 262.950 343.950 265.050 344.400 ;
        RECT 271.950 345.600 274.050 346.050 ;
        RECT 280.950 345.600 283.050 346.050 ;
        RECT 361.950 345.600 364.050 346.050 ;
        RECT 400.950 345.600 403.050 346.050 ;
        RECT 271.950 344.400 303.600 345.600 ;
        RECT 271.950 343.950 274.050 344.400 ;
        RECT 280.950 343.950 283.050 344.400 ;
        RECT 178.950 343.050 181.050 343.200 ;
        RECT 79.950 342.600 82.050 343.050 ;
        RECT 88.950 342.600 91.050 343.050 ;
        RECT 79.950 341.400 91.050 342.600 ;
        RECT 79.950 340.950 82.050 341.400 ;
        RECT 88.950 340.950 91.050 341.400 ;
        RECT 142.950 342.600 145.050 343.050 ;
        RECT 178.950 342.600 183.000 343.050 ;
        RECT 302.400 342.600 303.600 344.400 ;
        RECT 361.950 344.400 403.050 345.600 ;
        RECT 361.950 343.950 364.050 344.400 ;
        RECT 400.950 343.950 403.050 344.400 ;
        RECT 472.950 345.600 475.050 346.050 ;
        RECT 508.950 345.600 511.050 346.050 ;
        RECT 472.950 344.400 511.050 345.600 ;
        RECT 472.950 343.950 475.050 344.400 ;
        RECT 508.950 343.950 511.050 344.400 ;
        RECT 541.950 343.950 544.050 346.050 ;
        RECT 550.950 345.600 553.050 346.050 ;
        RECT 586.950 345.600 589.050 346.050 ;
        RECT 607.950 345.600 610.050 346.050 ;
        RECT 628.950 345.600 631.050 346.050 ;
        RECT 634.950 345.600 637.050 346.050 ;
        RECT 550.950 344.400 637.050 345.600 ;
        RECT 550.950 343.950 553.050 344.400 ;
        RECT 586.950 343.950 589.050 344.400 ;
        RECT 607.950 343.950 610.050 344.400 ;
        RECT 628.950 343.950 631.050 344.400 ;
        RECT 634.950 343.950 637.050 344.400 ;
        RECT 640.950 345.600 643.050 346.050 ;
        RECT 682.950 345.600 685.050 346.050 ;
        RECT 640.950 344.400 685.050 345.600 ;
        RECT 640.950 343.950 643.050 344.400 ;
        RECT 682.950 343.950 685.050 344.400 ;
        RECT 694.950 345.600 697.050 346.050 ;
        RECT 742.950 345.600 745.050 346.050 ;
        RECT 694.950 344.400 745.050 345.600 ;
        RECT 694.950 343.950 697.050 344.400 ;
        RECT 742.950 343.950 745.050 344.400 ;
        RECT 748.950 345.600 751.050 346.050 ;
        RECT 754.950 345.600 757.050 346.050 ;
        RECT 748.950 344.400 757.050 345.600 ;
        RECT 748.950 343.950 751.050 344.400 ;
        RECT 754.950 343.950 757.050 344.400 ;
        RECT 766.950 345.600 769.050 346.050 ;
        RECT 787.950 345.600 790.050 346.050 ;
        RECT 766.950 344.400 790.050 345.600 ;
        RECT 766.950 343.950 769.050 344.400 ;
        RECT 787.950 343.950 790.050 344.400 ;
        RECT 799.950 345.600 802.050 346.050 ;
        RECT 805.950 345.600 808.050 346.050 ;
        RECT 799.950 344.400 808.050 345.600 ;
        RECT 799.950 343.950 802.050 344.400 ;
        RECT 805.950 343.950 808.050 344.400 ;
        RECT 820.950 345.600 823.050 346.050 ;
        RECT 826.950 345.600 829.050 346.050 ;
        RECT 820.950 344.400 829.050 345.600 ;
        RECT 820.950 343.950 823.050 344.400 ;
        RECT 826.950 343.950 829.050 344.400 ;
        RECT 835.950 345.600 838.050 345.900 ;
        RECT 844.950 345.600 847.050 346.050 ;
        RECT 835.950 344.400 847.050 345.600 ;
        RECT 313.950 342.600 316.050 343.050 ;
        RECT 142.950 341.400 183.600 342.600 ;
        RECT 302.400 341.400 316.050 342.600 ;
        RECT 142.950 340.950 145.050 341.400 ;
        RECT 178.950 341.100 183.000 341.400 ;
        RECT 180.000 340.950 183.000 341.100 ;
        RECT 313.950 340.950 316.050 341.400 ;
        RECT 421.950 342.600 424.050 343.050 ;
        RECT 433.950 342.600 436.050 343.050 ;
        RECT 421.950 341.400 436.050 342.600 ;
        RECT 421.950 340.950 424.050 341.400 ;
        RECT 433.950 340.950 436.050 341.400 ;
        RECT 532.950 342.600 535.050 343.050 ;
        RECT 538.950 342.600 541.050 343.050 ;
        RECT 532.950 341.400 541.050 342.600 ;
        RECT 532.950 340.950 535.050 341.400 ;
        RECT 538.950 340.950 541.050 341.400 ;
        RECT 22.950 339.750 25.050 340.200 ;
        RECT 28.800 339.750 30.900 340.200 ;
        RECT 22.950 338.550 30.900 339.750 ;
        RECT 22.950 338.100 25.050 338.550 ;
        RECT 28.800 338.100 30.900 338.550 ;
        RECT 31.950 339.600 34.050 340.050 ;
        RECT 40.950 339.600 43.050 340.200 ;
        RECT 31.950 338.400 43.050 339.600 ;
        RECT 31.950 337.950 34.050 338.400 ;
        RECT 40.950 338.100 43.050 338.400 ;
        RECT 58.950 339.600 61.050 340.200 ;
        RECT 67.950 339.600 70.050 340.050 ;
        RECT 58.950 338.400 70.050 339.600 ;
        RECT 58.950 338.100 61.050 338.400 ;
        RECT 67.950 337.950 70.050 338.400 ;
        RECT 85.950 339.600 88.050 340.200 ;
        RECT 97.950 339.600 100.050 340.200 ;
        RECT 85.950 338.400 100.050 339.600 ;
        RECT 85.950 338.100 88.050 338.400 ;
        RECT 97.950 338.100 100.050 338.400 ;
        RECT 103.950 338.100 106.050 340.200 ;
        RECT 112.950 339.600 115.050 340.050 ;
        RECT 118.950 339.600 121.050 340.200 ;
        RECT 112.950 338.400 121.050 339.600 ;
        RECT 19.950 333.450 22.050 333.900 ;
        RECT 31.950 333.450 34.050 333.900 ;
        RECT 19.950 332.250 34.050 333.450 ;
        RECT 104.400 333.600 105.600 338.100 ;
        RECT 112.950 337.950 115.050 338.400 ;
        RECT 118.950 338.100 121.050 338.400 ;
        RECT 124.950 339.750 127.050 340.200 ;
        RECT 133.950 339.750 136.050 340.200 ;
        RECT 124.950 338.550 136.050 339.750 ;
        RECT 124.950 338.100 127.050 338.550 ;
        RECT 133.950 338.100 136.050 338.550 ;
        RECT 166.950 339.600 169.050 340.200 ;
        RECT 178.950 339.600 181.050 340.050 ;
        RECT 166.950 338.400 181.050 339.600 ;
        RECT 166.950 338.100 169.050 338.400 ;
        RECT 178.950 337.950 181.050 338.400 ;
        RECT 184.950 339.750 187.050 340.200 ;
        RECT 193.950 339.750 196.050 340.200 ;
        RECT 184.950 339.600 196.050 339.750 ;
        RECT 205.950 339.600 208.050 340.200 ;
        RECT 184.950 338.550 208.050 339.600 ;
        RECT 184.950 338.100 187.050 338.550 ;
        RECT 193.950 338.400 208.050 338.550 ;
        RECT 193.950 338.100 196.050 338.400 ;
        RECT 205.950 338.100 208.050 338.400 ;
        RECT 226.950 339.600 229.050 340.200 ;
        RECT 232.950 339.600 235.050 340.050 ;
        RECT 244.950 339.600 247.050 340.200 ;
        RECT 226.950 338.400 247.050 339.600 ;
        RECT 226.950 338.100 229.050 338.400 ;
        RECT 232.950 337.950 235.050 338.400 ;
        RECT 244.950 338.100 247.050 338.400 ;
        RECT 298.950 338.100 301.050 340.200 ;
        RECT 316.950 339.600 319.050 340.200 ;
        RECT 370.950 339.600 373.050 340.050 ;
        RECT 379.950 339.600 382.050 340.200 ;
        RECT 316.950 338.400 348.600 339.600 ;
        RECT 316.950 338.100 319.050 338.400 ;
        RECT 121.950 333.600 124.050 333.900 ;
        RECT 104.400 332.400 124.050 333.600 ;
        RECT 19.950 331.800 22.050 332.250 ;
        RECT 31.950 331.800 34.050 332.250 ;
        RECT 121.950 331.800 124.050 332.400 ;
        RECT 127.950 333.600 130.050 333.900 ;
        RECT 139.950 333.600 142.050 333.900 ;
        RECT 127.950 332.400 142.050 333.600 ;
        RECT 127.950 331.800 130.050 332.400 ;
        RECT 139.950 331.800 142.050 332.400 ;
        RECT 151.950 333.450 154.050 333.900 ;
        RECT 157.950 333.450 160.050 333.900 ;
        RECT 151.950 332.250 160.050 333.450 ;
        RECT 151.950 331.800 154.050 332.250 ;
        RECT 157.950 331.800 160.050 332.250 ;
        RECT 187.950 333.600 190.050 333.900 ;
        RECT 202.950 333.600 205.050 333.900 ;
        RECT 187.950 332.400 205.050 333.600 ;
        RECT 187.950 331.800 190.050 332.400 ;
        RECT 202.950 331.800 205.050 332.400 ;
        RECT 208.950 333.600 211.050 333.900 ;
        RECT 223.950 333.600 226.050 333.900 ;
        RECT 208.950 332.400 226.050 333.600 ;
        RECT 208.950 331.800 211.050 332.400 ;
        RECT 223.950 331.800 226.050 332.400 ;
        RECT 265.950 333.450 268.050 333.900 ;
        RECT 271.950 333.450 274.050 333.900 ;
        RECT 265.950 332.250 274.050 333.450 ;
        RECT 265.950 331.800 268.050 332.250 ;
        RECT 271.950 331.800 274.050 332.250 ;
        RECT 299.400 331.050 300.600 338.100 ;
        RECT 347.400 334.050 348.600 338.400 ;
        RECT 370.950 338.400 382.050 339.600 ;
        RECT 370.950 337.950 373.050 338.400 ;
        RECT 379.950 338.100 382.050 338.400 ;
        RECT 388.950 339.600 391.050 340.200 ;
        RECT 397.950 339.600 400.050 340.050 ;
        RECT 388.950 338.400 400.050 339.600 ;
        RECT 388.950 338.100 391.050 338.400 ;
        RECT 397.950 337.950 400.050 338.400 ;
        RECT 439.950 338.100 442.050 340.200 ;
        RECT 451.950 339.600 454.050 340.050 ;
        RECT 469.950 339.600 472.050 340.050 ;
        RECT 451.950 338.400 472.050 339.600 ;
        RECT 440.400 334.050 441.600 338.100 ;
        RECT 451.950 337.950 454.050 338.400 ;
        RECT 469.950 337.950 472.050 338.400 ;
        RECT 475.950 338.100 478.050 340.200 ;
        RECT 504.000 339.600 508.050 340.050 ;
        RECT 313.950 333.450 316.050 333.900 ;
        RECT 328.950 333.450 331.050 333.900 ;
        RECT 313.950 332.250 331.050 333.450 ;
        RECT 313.950 331.800 316.050 332.250 ;
        RECT 328.950 331.800 331.050 332.250 ;
        RECT 346.950 331.950 349.050 334.050 ;
        RECT 364.950 333.450 367.050 333.900 ;
        RECT 370.950 333.450 373.050 333.900 ;
        RECT 364.950 332.250 373.050 333.450 ;
        RECT 364.950 331.800 367.050 332.250 ;
        RECT 370.950 331.800 373.050 332.250 ;
        RECT 400.950 333.450 403.050 333.900 ;
        RECT 406.950 333.450 409.050 333.900 ;
        RECT 400.950 332.250 409.050 333.450 ;
        RECT 400.950 331.800 403.050 332.250 ;
        RECT 406.950 331.800 409.050 332.250 ;
        RECT 436.950 332.400 441.600 334.050 ;
        RECT 448.950 333.600 451.050 334.050 ;
        RECT 469.950 333.600 472.050 334.050 ;
        RECT 448.950 332.400 472.050 333.600 ;
        RECT 476.400 333.600 477.600 338.100 ;
        RECT 503.400 337.950 508.050 339.600 ;
        RECT 517.950 338.100 520.050 340.200 ;
        RECT 490.800 333.600 492.900 334.050 ;
        RECT 476.400 332.400 492.900 333.600 ;
        RECT 436.950 331.950 441.000 332.400 ;
        RECT 448.950 331.950 451.050 332.400 ;
        RECT 469.950 331.950 472.050 332.400 ;
        RECT 490.800 331.950 492.900 332.400 ;
        RECT 493.950 333.600 496.050 333.900 ;
        RECT 503.400 333.600 504.600 337.950 ;
        RECT 518.400 333.600 519.600 338.100 ;
        RECT 529.950 337.950 532.050 340.050 ;
        RECT 542.400 339.600 543.600 343.950 ;
        RECT 835.950 343.800 838.050 344.400 ;
        RECT 844.950 343.950 847.050 344.400 ;
        RECT 853.950 345.600 856.050 346.050 ;
        RECT 859.950 345.600 862.050 346.050 ;
        RECT 853.950 344.400 862.050 345.600 ;
        RECT 853.950 343.950 856.050 344.400 ;
        RECT 859.950 343.950 862.050 344.400 ;
        RECT 589.950 340.950 592.050 343.050 ;
        RECT 539.400 338.400 543.600 339.600 ;
        RECT 493.950 332.400 504.600 333.600 ;
        RECT 512.400 333.000 519.600 333.600 ;
        RECT 511.950 332.400 519.600 333.000 ;
        RECT 526.950 333.600 529.050 333.900 ;
        RECT 530.400 333.600 531.600 337.950 ;
        RECT 539.400 333.900 540.600 338.400 ;
        RECT 590.400 336.600 591.600 340.950 ;
        RECT 601.950 339.600 604.050 340.200 ;
        RECT 627.000 339.600 631.050 340.050 ;
        RECT 601.950 338.400 606.600 339.600 ;
        RECT 601.950 338.100 604.050 338.400 ;
        RECT 605.400 336.600 606.600 338.400 ;
        RECT 626.400 337.950 631.050 339.600 ;
        RECT 643.950 339.600 646.050 340.200 ;
        RECT 649.950 339.600 652.050 343.050 ;
        RECT 805.950 342.600 808.050 342.900 ;
        RECT 817.950 342.600 820.050 343.050 ;
        RECT 805.950 341.400 820.050 342.600 ;
        RECT 805.950 340.800 808.050 341.400 ;
        RECT 817.950 340.950 820.050 341.400 ;
        RECT 829.950 342.600 832.050 343.050 ;
        RECT 868.950 342.600 871.050 343.050 ;
        RECT 874.950 342.600 877.050 343.050 ;
        RECT 829.950 341.400 843.600 342.600 ;
        RECT 829.950 340.950 832.050 341.400 ;
        RECT 643.950 339.000 652.050 339.600 ;
        RECT 643.950 338.400 651.600 339.000 ;
        RECT 643.950 338.100 646.050 338.400 ;
        RECT 658.950 338.100 661.050 340.200 ;
        RECT 682.950 339.600 685.050 340.200 ;
        RECT 700.950 339.600 703.050 340.200 ;
        RECT 682.950 338.400 703.050 339.600 ;
        RECT 682.950 338.100 685.050 338.400 ;
        RECT 700.950 338.100 703.050 338.400 ;
        RECT 712.950 339.750 715.050 340.200 ;
        RECT 721.950 339.750 724.050 340.200 ;
        RECT 712.950 338.550 724.050 339.750 ;
        RECT 712.950 338.100 715.050 338.550 ;
        RECT 721.950 338.100 724.050 338.550 ;
        RECT 727.950 339.600 730.050 340.200 ;
        RECT 748.950 339.600 751.050 340.200 ;
        RECT 772.950 339.600 775.050 340.200 ;
        RECT 787.950 339.600 790.050 340.200 ;
        RECT 727.950 338.400 732.600 339.600 ;
        RECT 727.950 338.100 730.050 338.400 ;
        RECT 590.400 335.400 603.600 336.600 ;
        RECT 605.400 335.400 609.600 336.600 ;
        RECT 526.950 332.400 531.600 333.600 ;
        RECT 493.950 331.800 496.050 332.400 ;
        RECT 100.950 330.600 103.050 331.050 ;
        RECT 127.950 330.600 130.050 331.050 ;
        RECT 100.950 329.400 130.050 330.600 ;
        RECT 100.950 328.950 103.050 329.400 ;
        RECT 127.950 328.950 130.050 329.400 ;
        RECT 181.950 330.600 184.050 331.050 ;
        RECT 208.950 330.600 211.050 331.050 ;
        RECT 181.950 329.400 211.050 330.600 ;
        RECT 181.950 328.950 184.050 329.400 ;
        RECT 208.950 328.950 211.050 329.400 ;
        RECT 274.950 330.600 277.050 331.050 ;
        RECT 286.950 330.600 289.050 331.050 ;
        RECT 274.950 329.400 289.050 330.600 ;
        RECT 274.950 328.950 277.050 329.400 ;
        RECT 286.950 328.950 289.050 329.400 ;
        RECT 298.950 328.950 301.050 331.050 ;
        RECT 319.950 330.600 322.050 331.050 ;
        RECT 325.950 330.600 328.050 331.050 ;
        RECT 319.950 329.400 328.050 330.600 ;
        RECT 319.950 328.950 322.050 329.400 ;
        RECT 325.950 328.950 328.050 329.400 ;
        RECT 466.950 330.600 469.050 331.050 ;
        RECT 484.950 330.600 487.050 331.050 ;
        RECT 466.950 329.400 487.050 330.600 ;
        RECT 466.950 328.950 469.050 329.400 ;
        RECT 484.950 328.950 487.050 329.400 ;
        RECT 511.950 328.950 514.050 332.400 ;
        RECT 526.950 331.800 529.050 332.400 ;
        RECT 538.950 331.800 541.050 333.900 ;
        RECT 553.950 333.450 556.050 333.900 ;
        RECT 559.950 333.450 562.050 333.900 ;
        RECT 553.950 332.250 562.050 333.450 ;
        RECT 553.950 331.800 556.050 332.250 ;
        RECT 559.950 331.800 562.050 332.250 ;
        RECT 592.950 333.450 595.050 333.900 ;
        RECT 598.950 333.450 601.050 333.900 ;
        RECT 592.950 332.250 601.050 333.450 ;
        RECT 602.400 333.600 603.600 335.400 ;
        RECT 604.950 333.600 607.050 333.900 ;
        RECT 602.400 332.400 607.050 333.600 ;
        RECT 608.400 333.600 609.600 335.400 ;
        RECT 616.950 333.600 619.050 334.050 ;
        RECT 626.400 333.900 627.600 337.950 ;
        RECT 659.400 336.600 660.600 338.100 ;
        RECT 656.400 335.400 660.600 336.600 ;
        RECT 608.400 332.400 619.050 333.600 ;
        RECT 592.950 331.800 595.050 332.250 ;
        RECT 598.950 331.800 601.050 332.250 ;
        RECT 604.950 331.800 607.050 332.400 ;
        RECT 616.950 331.950 619.050 332.400 ;
        RECT 625.950 331.800 628.050 333.900 ;
        RECT 649.950 333.600 652.050 334.050 ;
        RECT 656.400 333.600 657.600 335.400 ;
        RECT 731.400 334.050 732.600 338.400 ;
        RECT 748.950 338.400 790.050 339.600 ;
        RECT 748.950 338.100 751.050 338.400 ;
        RECT 772.950 338.100 775.050 338.400 ;
        RECT 787.950 338.100 790.050 338.400 ;
        RECT 793.950 337.950 796.050 340.050 ;
        RECT 799.950 339.600 804.000 340.050 ;
        RECT 835.950 339.600 838.050 340.050 ;
        RECT 799.950 337.950 804.600 339.600 ;
        RECT 794.400 334.050 795.600 337.950 ;
        RECT 803.400 336.600 804.600 337.950 ;
        RECT 815.400 338.400 838.050 339.600 ;
        RECT 803.400 335.400 810.600 336.600 ;
        RECT 649.950 332.400 657.600 333.600 ;
        RECT 706.950 333.600 709.050 333.900 ;
        RECT 724.950 333.600 727.050 333.900 ;
        RECT 706.950 332.400 727.050 333.600 ;
        RECT 649.950 331.950 652.050 332.400 ;
        RECT 706.950 331.800 709.050 332.400 ;
        RECT 724.950 331.800 727.050 332.400 ;
        RECT 730.950 331.950 733.050 334.050 ;
        RECT 745.950 333.600 748.050 333.900 ;
        RECT 757.950 333.600 760.050 333.900 ;
        RECT 745.950 333.450 760.050 333.600 ;
        RECT 769.950 333.450 772.050 333.900 ;
        RECT 745.950 332.400 772.050 333.450 ;
        RECT 794.400 332.400 799.050 334.050 ;
        RECT 809.400 333.900 810.600 335.400 ;
        RECT 815.400 334.050 816.600 338.400 ;
        RECT 835.950 337.950 838.050 338.400 ;
        RECT 745.950 331.800 748.050 332.400 ;
        RECT 757.950 332.250 772.050 332.400 ;
        RECT 757.950 331.800 760.050 332.250 ;
        RECT 769.950 331.800 772.050 332.250 ;
        RECT 795.000 331.950 799.050 332.400 ;
        RECT 808.950 331.800 811.050 333.900 ;
        RECT 814.950 331.950 817.050 334.050 ;
        RECT 842.400 333.900 843.600 341.400 ;
        RECT 868.950 341.400 877.050 342.600 ;
        RECT 868.950 340.950 871.050 341.400 ;
        RECT 874.950 340.950 877.050 341.400 ;
        RECT 862.950 338.100 865.050 340.200 ;
        RECT 829.950 331.800 832.050 333.900 ;
        RECT 841.950 331.800 844.050 333.900 ;
        RECT 607.950 330.600 610.050 331.050 ;
        RECT 619.950 330.600 622.050 331.050 ;
        RECT 607.950 329.400 622.050 330.600 ;
        RECT 607.950 328.950 610.050 329.400 ;
        RECT 619.950 328.950 622.050 329.400 ;
        RECT 808.950 330.600 811.050 331.050 ;
        RECT 830.400 330.600 831.600 331.800 ;
        RECT 863.400 331.050 864.600 338.100 ;
        RECT 808.950 329.400 831.600 330.600 ;
        RECT 844.950 330.600 847.050 331.050 ;
        RECT 856.950 330.600 859.050 331.050 ;
        RECT 844.950 329.400 859.050 330.600 ;
        RECT 808.950 328.950 811.050 329.400 ;
        RECT 844.950 328.950 847.050 329.400 ;
        RECT 856.950 328.950 859.050 329.400 ;
        RECT 862.950 328.950 865.050 331.050 ;
        RECT 67.950 327.600 70.050 328.050 ;
        RECT 82.950 327.600 85.050 328.050 ;
        RECT 67.950 326.400 85.050 327.600 ;
        RECT 67.950 325.950 70.050 326.400 ;
        RECT 82.950 325.950 85.050 326.400 ;
        RECT 103.950 327.600 106.050 328.050 ;
        RECT 121.950 327.600 124.050 328.050 ;
        RECT 103.950 326.400 124.050 327.600 ;
        RECT 103.950 325.950 106.050 326.400 ;
        RECT 121.950 325.950 124.050 326.400 ;
        RECT 139.950 327.600 142.050 328.050 ;
        RECT 163.950 327.600 166.050 328.050 ;
        RECT 139.950 326.400 166.050 327.600 ;
        RECT 139.950 325.950 142.050 326.400 ;
        RECT 163.950 325.950 166.050 326.400 ;
        RECT 193.950 327.600 196.050 328.050 ;
        RECT 199.950 327.600 202.050 328.050 ;
        RECT 193.950 326.400 202.050 327.600 ;
        RECT 193.950 325.950 196.050 326.400 ;
        RECT 199.950 325.950 202.050 326.400 ;
        RECT 229.950 327.600 232.050 328.050 ;
        RECT 241.950 327.600 244.050 328.050 ;
        RECT 313.950 327.600 316.050 328.050 ;
        RECT 229.950 326.400 316.050 327.600 ;
        RECT 229.950 325.950 232.050 326.400 ;
        RECT 241.950 325.950 244.050 326.400 ;
        RECT 313.950 325.950 316.050 326.400 ;
        RECT 388.950 327.600 391.050 328.050 ;
        RECT 421.950 327.600 424.050 328.050 ;
        RECT 388.950 326.400 424.050 327.600 ;
        RECT 485.400 327.600 486.600 328.950 ;
        RECT 502.950 327.600 505.050 328.050 ;
        RECT 485.400 326.400 505.050 327.600 ;
        RECT 388.950 325.950 391.050 326.400 ;
        RECT 421.950 325.950 424.050 326.400 ;
        RECT 502.950 325.950 505.050 326.400 ;
        RECT 526.950 327.600 529.050 328.050 ;
        RECT 562.950 327.600 565.050 328.050 ;
        RECT 526.950 326.400 565.050 327.600 ;
        RECT 526.950 325.950 529.050 326.400 ;
        RECT 562.950 325.950 565.050 326.400 ;
        RECT 571.950 327.600 574.050 328.050 ;
        RECT 580.950 327.600 583.050 328.050 ;
        RECT 571.950 326.400 583.050 327.600 ;
        RECT 571.950 325.950 574.050 326.400 ;
        RECT 580.950 325.950 583.050 326.400 ;
        RECT 598.950 327.600 601.050 328.050 ;
        RECT 649.950 327.600 652.050 328.050 ;
        RECT 598.950 326.400 652.050 327.600 ;
        RECT 598.950 325.950 601.050 326.400 ;
        RECT 649.950 325.950 652.050 326.400 ;
        RECT 655.950 327.600 658.050 328.050 ;
        RECT 670.950 327.600 673.050 327.900 ;
        RECT 655.950 326.400 673.050 327.600 ;
        RECT 655.950 325.950 658.050 326.400 ;
        RECT 670.950 325.800 673.050 326.400 ;
        RECT 799.950 327.600 802.050 328.050 ;
        RECT 823.950 327.600 826.050 328.050 ;
        RECT 799.950 326.400 826.050 327.600 ;
        RECT 799.950 325.950 802.050 326.400 ;
        RECT 823.950 325.950 826.050 326.400 ;
        RECT 61.950 324.600 64.050 325.050 ;
        RECT 112.950 324.600 115.050 325.050 ;
        RECT 61.950 323.400 115.050 324.600 ;
        RECT 61.950 322.950 64.050 323.400 ;
        RECT 112.950 322.950 115.050 323.400 ;
        RECT 259.950 324.600 262.050 325.050 ;
        RECT 289.950 324.600 292.050 325.050 ;
        RECT 295.950 324.600 298.050 325.050 ;
        RECT 259.950 323.400 298.050 324.600 ;
        RECT 259.950 322.950 262.050 323.400 ;
        RECT 289.950 322.950 292.050 323.400 ;
        RECT 295.950 322.950 298.050 323.400 ;
        RECT 337.950 324.600 340.050 325.050 ;
        RECT 400.950 324.600 403.050 325.050 ;
        RECT 337.950 323.400 403.050 324.600 ;
        RECT 337.950 322.950 340.050 323.400 ;
        RECT 400.950 322.950 403.050 323.400 ;
        RECT 433.950 324.600 436.050 325.050 ;
        RECT 451.800 324.600 453.900 325.050 ;
        RECT 433.950 323.400 453.900 324.600 ;
        RECT 433.950 322.950 436.050 323.400 ;
        RECT 451.800 322.950 453.900 323.400 ;
        RECT 454.950 324.600 457.050 325.050 ;
        RECT 532.950 324.600 535.050 325.050 ;
        RECT 454.950 323.400 535.050 324.600 ;
        RECT 454.950 322.950 457.050 323.400 ;
        RECT 532.950 322.950 535.050 323.400 ;
        RECT 646.950 324.600 649.050 325.050 ;
        RECT 697.950 324.600 700.050 325.050 ;
        RECT 646.950 323.400 700.050 324.600 ;
        RECT 646.950 322.950 649.050 323.400 ;
        RECT 697.950 322.950 700.050 323.400 ;
        RECT 760.950 324.600 763.050 325.050 ;
        RECT 778.950 324.600 781.050 325.050 ;
        RECT 862.950 324.600 865.050 325.050 ;
        RECT 760.950 323.400 781.050 324.600 ;
        RECT 760.950 322.950 763.050 323.400 ;
        RECT 778.950 322.950 781.050 323.400 ;
        RECT 785.400 323.400 865.050 324.600 ;
        RECT 76.950 321.600 79.050 322.050 ;
        RECT 91.950 321.600 94.050 322.050 ;
        RECT 76.950 320.400 94.050 321.600 ;
        RECT 76.950 319.950 79.050 320.400 ;
        RECT 91.950 319.950 94.050 320.400 ;
        RECT 121.950 321.600 124.050 322.050 ;
        RECT 133.950 321.600 136.050 322.050 ;
        RECT 121.950 320.400 136.050 321.600 ;
        RECT 121.950 319.950 124.050 320.400 ;
        RECT 133.950 319.950 136.050 320.400 ;
        RECT 325.950 321.600 328.050 322.050 ;
        RECT 361.950 321.600 364.050 322.050 ;
        RECT 376.950 321.600 379.050 322.050 ;
        RECT 409.950 321.600 412.050 322.050 ;
        RECT 325.950 320.400 412.050 321.600 ;
        RECT 325.950 319.950 328.050 320.400 ;
        RECT 361.950 319.950 364.050 320.400 ;
        RECT 376.950 319.950 379.050 320.400 ;
        RECT 409.950 319.950 412.050 320.400 ;
        RECT 553.950 321.600 556.050 322.050 ;
        RECT 571.950 321.600 574.050 322.050 ;
        RECT 553.950 320.400 574.050 321.600 ;
        RECT 553.950 319.950 556.050 320.400 ;
        RECT 571.950 319.950 574.050 320.400 ;
        RECT 604.950 321.600 607.050 322.050 ;
        RECT 613.950 321.600 616.050 322.050 ;
        RECT 640.950 321.600 643.050 322.050 ;
        RECT 604.950 320.400 643.050 321.600 ;
        RECT 604.950 319.950 607.050 320.400 ;
        RECT 613.950 319.950 616.050 320.400 ;
        RECT 640.950 319.950 643.050 320.400 ;
        RECT 661.950 321.600 664.050 322.050 ;
        RECT 718.950 321.600 721.050 322.050 ;
        RECT 661.950 320.400 721.050 321.600 ;
        RECT 661.950 319.950 664.050 320.400 ;
        RECT 718.950 319.950 721.050 320.400 ;
        RECT 733.950 321.600 736.050 322.050 ;
        RECT 772.950 321.600 775.050 322.050 ;
        RECT 785.400 321.600 786.600 323.400 ;
        RECT 862.950 322.950 865.050 323.400 ;
        RECT 733.950 320.400 744.600 321.600 ;
        RECT 733.950 319.950 736.050 320.400 ;
        RECT 247.950 318.600 250.050 319.050 ;
        RECT 265.950 318.600 268.050 319.050 ;
        RECT 247.950 317.400 268.050 318.600 ;
        RECT 247.950 316.950 250.050 317.400 ;
        RECT 265.950 316.950 268.050 317.400 ;
        RECT 316.950 318.600 319.050 319.050 ;
        RECT 382.950 318.600 385.050 319.050 ;
        RECT 316.950 317.400 385.050 318.600 ;
        RECT 316.950 316.950 319.050 317.400 ;
        RECT 382.950 316.950 385.050 317.400 ;
        RECT 499.950 318.600 502.050 319.050 ;
        RECT 511.950 318.600 514.050 319.050 ;
        RECT 499.950 317.400 514.050 318.600 ;
        RECT 499.950 316.950 502.050 317.400 ;
        RECT 511.950 316.950 514.050 317.400 ;
        RECT 622.950 318.600 625.050 319.050 ;
        RECT 658.950 318.600 661.050 319.050 ;
        RECT 622.950 317.400 661.050 318.600 ;
        RECT 622.950 316.950 625.050 317.400 ;
        RECT 658.950 316.950 661.050 317.400 ;
        RECT 679.950 318.600 682.050 319.050 ;
        RECT 688.950 318.600 691.050 319.050 ;
        RECT 679.950 317.400 691.050 318.600 ;
        RECT 679.950 316.950 682.050 317.400 ;
        RECT 688.950 316.950 691.050 317.400 ;
        RECT 712.950 318.600 715.050 319.050 ;
        RECT 739.950 318.600 742.050 319.050 ;
        RECT 712.950 317.400 742.050 318.600 ;
        RECT 743.400 318.600 744.600 320.400 ;
        RECT 772.950 320.400 786.600 321.600 ;
        RECT 802.950 321.600 805.050 322.050 ;
        RECT 817.950 321.600 820.050 322.050 ;
        RECT 802.950 320.400 820.050 321.600 ;
        RECT 772.950 319.950 775.050 320.400 ;
        RECT 802.950 319.950 805.050 320.400 ;
        RECT 817.950 319.950 820.050 320.400 ;
        RECT 769.950 318.600 772.050 319.050 ;
        RECT 743.400 317.400 772.050 318.600 ;
        RECT 712.950 316.950 715.050 317.400 ;
        RECT 13.950 315.600 16.050 316.050 ;
        RECT 37.950 315.600 40.050 316.050 ;
        RECT 55.950 315.600 58.050 316.050 ;
        RECT 76.950 315.600 79.050 316.050 ;
        RECT 13.950 314.400 79.050 315.600 ;
        RECT 13.950 313.950 16.050 314.400 ;
        RECT 37.950 313.950 40.050 314.400 ;
        RECT 55.950 313.950 58.050 314.400 ;
        RECT 76.950 313.950 79.050 314.400 ;
        RECT 127.950 315.600 130.050 316.050 ;
        RECT 274.950 315.600 277.050 316.050 ;
        RECT 127.950 314.400 277.050 315.600 ;
        RECT 127.950 313.950 130.050 314.400 ;
        RECT 274.950 313.950 277.050 314.400 ;
        RECT 415.950 315.600 418.050 316.050 ;
        RECT 466.950 315.600 469.050 316.050 ;
        RECT 415.950 314.400 469.050 315.600 ;
        RECT 415.950 313.950 418.050 314.400 ;
        RECT 466.950 313.950 469.050 314.400 ;
        RECT 472.950 315.600 475.050 316.050 ;
        RECT 496.950 315.600 499.050 316.050 ;
        RECT 523.950 315.600 526.050 316.050 ;
        RECT 565.950 315.600 568.050 316.050 ;
        RECT 472.950 314.400 568.050 315.600 ;
        RECT 472.950 313.950 475.050 314.400 ;
        RECT 496.950 313.950 499.050 314.400 ;
        RECT 523.950 313.950 526.050 314.400 ;
        RECT 565.950 313.950 568.050 314.400 ;
        RECT 670.950 315.600 673.050 316.050 ;
        RECT 739.950 315.600 742.050 317.400 ;
        RECT 769.950 316.950 772.050 317.400 ;
        RECT 796.950 318.600 799.050 319.050 ;
        RECT 817.800 318.600 819.900 318.900 ;
        RECT 796.950 317.400 819.900 318.600 ;
        RECT 796.950 316.950 799.050 317.400 ;
        RECT 817.800 316.800 819.900 317.400 ;
        RECT 820.950 318.600 823.050 319.050 ;
        RECT 835.950 318.600 838.050 319.050 ;
        RECT 820.950 317.400 838.050 318.600 ;
        RECT 820.950 316.950 823.050 317.400 ;
        RECT 835.950 316.950 838.050 317.400 ;
        RECT 670.950 315.000 742.050 315.600 ;
        RECT 778.950 315.600 781.050 316.050 ;
        RECT 814.950 315.600 817.050 316.050 ;
        RECT 670.950 314.400 741.600 315.000 ;
        RECT 778.950 314.400 817.050 315.600 ;
        RECT 670.950 313.950 673.050 314.400 ;
        RECT 778.950 313.950 781.050 314.400 ;
        RECT 814.950 313.950 817.050 314.400 ;
        RECT 319.950 312.600 322.050 313.050 ;
        RECT 358.950 312.600 361.050 313.050 ;
        RECT 319.950 311.400 361.050 312.600 ;
        RECT 319.950 310.950 322.050 311.400 ;
        RECT 358.950 310.950 361.050 311.400 ;
        RECT 382.950 312.600 385.050 313.050 ;
        RECT 436.950 312.600 439.050 313.050 ;
        RECT 382.950 311.400 439.050 312.600 ;
        RECT 382.950 310.950 385.050 311.400 ;
        RECT 436.950 310.950 439.050 311.400 ;
        RECT 469.950 312.600 472.050 313.050 ;
        RECT 517.950 312.600 520.050 313.050 ;
        RECT 571.950 312.600 574.050 313.050 ;
        RECT 607.950 312.600 610.050 313.050 ;
        RECT 469.950 311.400 570.600 312.600 ;
        RECT 469.950 310.950 472.050 311.400 ;
        RECT 517.950 310.950 520.050 311.400 ;
        RECT 133.950 309.600 136.050 310.050 ;
        RECT 160.950 309.600 163.050 310.050 ;
        RECT 133.950 308.400 163.050 309.600 ;
        RECT 133.950 307.950 136.050 308.400 ;
        RECT 160.950 307.950 163.050 308.400 ;
        RECT 181.950 309.600 184.050 310.050 ;
        RECT 235.950 309.600 238.050 310.050 ;
        RECT 181.950 308.400 238.050 309.600 ;
        RECT 181.950 307.950 184.050 308.400 ;
        RECT 235.950 307.950 238.050 308.400 ;
        RECT 262.950 309.600 265.050 310.050 ;
        RECT 304.950 309.600 307.050 310.050 ;
        RECT 262.950 308.400 307.050 309.600 ;
        RECT 262.950 307.950 265.050 308.400 ;
        RECT 304.950 307.950 307.050 308.400 ;
        RECT 457.950 309.600 460.050 310.050 ;
        RECT 541.950 309.600 544.050 310.050 ;
        RECT 556.950 309.600 559.050 310.050 ;
        RECT 457.950 308.400 559.050 309.600 ;
        RECT 569.400 309.600 570.600 311.400 ;
        RECT 571.950 311.400 610.050 312.600 ;
        RECT 571.950 310.950 574.050 311.400 ;
        RECT 607.950 310.950 610.050 311.400 ;
        RECT 640.950 312.600 643.050 313.050 ;
        RECT 646.950 312.600 649.050 313.050 ;
        RECT 640.950 311.400 649.050 312.600 ;
        RECT 640.950 310.950 643.050 311.400 ;
        RECT 646.950 310.950 649.050 311.400 ;
        RECT 730.950 312.600 733.050 313.050 ;
        RECT 763.950 312.600 766.050 313.050 ;
        RECT 730.950 311.400 766.050 312.600 ;
        RECT 730.950 310.950 733.050 311.400 ;
        RECT 763.950 310.950 766.050 311.400 ;
        RECT 598.950 309.600 601.050 310.050 ;
        RECT 569.400 308.400 601.050 309.600 ;
        RECT 457.950 307.950 460.050 308.400 ;
        RECT 541.950 307.950 544.050 308.400 ;
        RECT 556.950 307.950 559.050 308.400 ;
        RECT 598.950 307.950 601.050 308.400 ;
        RECT 655.950 309.600 658.050 310.050 ;
        RECT 688.950 309.600 691.050 310.050 ;
        RECT 655.950 308.400 691.050 309.600 ;
        RECT 655.950 307.950 658.050 308.400 ;
        RECT 688.950 307.950 691.050 308.400 ;
        RECT 778.950 309.600 781.050 310.050 ;
        RECT 826.950 309.600 829.050 310.050 ;
        RECT 778.950 308.400 829.050 309.600 ;
        RECT 778.950 307.950 781.050 308.400 ;
        RECT 826.950 307.950 829.050 308.400 ;
        RECT 79.950 306.600 82.050 307.050 ;
        RECT 127.950 306.600 130.050 307.050 ;
        RECT 79.950 305.400 130.050 306.600 ;
        RECT 79.950 304.950 82.050 305.400 ;
        RECT 127.950 304.950 130.050 305.400 ;
        RECT 274.950 306.600 277.050 307.050 ;
        RECT 304.950 306.600 307.050 306.900 ;
        RECT 319.950 306.600 322.050 307.050 ;
        RECT 274.950 305.400 307.050 306.600 ;
        RECT 274.950 304.950 277.050 305.400 ;
        RECT 304.950 304.800 307.050 305.400 ;
        RECT 308.400 305.400 322.050 306.600 ;
        RECT 106.950 303.600 109.050 304.050 ;
        RECT 121.950 303.600 124.050 304.050 ;
        RECT 106.950 302.400 124.050 303.600 ;
        RECT 106.950 301.950 109.050 302.400 ;
        RECT 121.950 301.950 124.050 302.400 ;
        RECT 142.950 303.600 145.050 304.050 ;
        RECT 217.950 303.600 220.050 304.050 ;
        RECT 142.950 302.400 220.050 303.600 ;
        RECT 142.950 301.950 145.050 302.400 ;
        RECT 217.950 301.950 220.050 302.400 ;
        RECT 244.950 303.600 247.050 304.050 ;
        RECT 253.950 303.600 256.050 304.050 ;
        RECT 244.950 302.400 256.050 303.600 ;
        RECT 244.950 301.950 247.050 302.400 ;
        RECT 253.950 301.950 256.050 302.400 ;
        RECT 283.950 303.600 286.050 304.050 ;
        RECT 308.400 303.600 309.600 305.400 ;
        RECT 319.950 304.950 322.050 305.400 ;
        RECT 328.950 306.600 331.050 307.050 ;
        RECT 334.950 306.600 337.050 307.050 ;
        RECT 367.950 306.600 370.050 307.050 ;
        RECT 328.950 305.400 370.050 306.600 ;
        RECT 328.950 304.950 331.050 305.400 ;
        RECT 334.950 304.950 337.050 305.400 ;
        RECT 367.950 304.950 370.050 305.400 ;
        RECT 433.950 306.600 436.050 307.050 ;
        RECT 472.800 306.600 474.900 307.050 ;
        RECT 433.950 305.400 474.900 306.600 ;
        RECT 433.950 304.950 436.050 305.400 ;
        RECT 472.800 304.950 474.900 305.400 ;
        RECT 475.950 306.600 478.050 307.050 ;
        RECT 487.950 306.600 490.050 307.050 ;
        RECT 475.950 305.400 490.050 306.600 ;
        RECT 475.950 304.950 478.050 305.400 ;
        RECT 487.950 304.950 490.050 305.400 ;
        RECT 559.950 306.600 562.050 307.050 ;
        RECT 619.950 306.600 622.050 307.050 ;
        RECT 559.950 305.400 622.050 306.600 ;
        RECT 559.950 304.950 562.050 305.400 ;
        RECT 619.950 304.950 622.050 305.400 ;
        RECT 658.950 306.600 661.050 307.050 ;
        RECT 679.950 306.600 682.050 307.050 ;
        RECT 658.950 305.400 682.050 306.600 ;
        RECT 658.950 304.950 661.050 305.400 ;
        RECT 679.950 304.950 682.050 305.400 ;
        RECT 703.950 306.600 706.050 307.050 ;
        RECT 715.950 306.600 718.050 307.050 ;
        RECT 721.950 306.600 724.050 307.050 ;
        RECT 730.950 306.600 733.050 307.050 ;
        RECT 703.950 305.400 733.050 306.600 ;
        RECT 703.950 304.950 706.050 305.400 ;
        RECT 715.950 304.950 718.050 305.400 ;
        RECT 721.950 304.950 724.050 305.400 ;
        RECT 730.950 304.950 733.050 305.400 ;
        RECT 742.950 306.600 745.050 307.050 ;
        RECT 763.950 306.600 766.050 307.050 ;
        RECT 742.950 305.400 766.050 306.600 ;
        RECT 742.950 304.950 745.050 305.400 ;
        RECT 763.950 304.950 766.050 305.400 ;
        RECT 769.950 306.600 772.050 307.050 ;
        RECT 796.950 306.600 799.050 307.050 ;
        RECT 769.950 305.400 799.050 306.600 ;
        RECT 769.950 304.950 772.050 305.400 ;
        RECT 796.950 304.950 799.050 305.400 ;
        RECT 283.950 302.400 309.600 303.600 ;
        RECT 415.950 303.600 418.050 304.050 ;
        RECT 445.950 303.600 448.050 304.050 ;
        RECT 415.950 302.400 448.050 303.600 ;
        RECT 283.950 301.950 286.050 302.400 ;
        RECT 415.950 301.950 418.050 302.400 ;
        RECT 445.950 301.950 448.050 302.400 ;
        RECT 670.950 303.600 673.050 304.050 ;
        RECT 685.950 303.600 688.050 304.050 ;
        RECT 670.950 302.400 688.050 303.600 ;
        RECT 670.950 301.950 673.050 302.400 ;
        RECT 685.950 301.950 688.050 302.400 ;
        RECT 697.950 303.600 700.050 304.050 ;
        RECT 760.950 303.600 763.050 304.050 ;
        RECT 697.950 302.400 763.050 303.600 ;
        RECT 697.950 301.950 700.050 302.400 ;
        RECT 760.950 301.950 763.050 302.400 ;
        RECT 772.950 303.600 775.050 304.050 ;
        RECT 799.950 303.600 802.050 304.050 ;
        RECT 772.950 302.400 802.050 303.600 ;
        RECT 772.950 301.950 775.050 302.400 ;
        RECT 799.950 301.950 802.050 302.400 ;
        RECT 187.950 300.600 190.050 301.050 ;
        RECT 295.950 300.600 298.050 301.050 ;
        RECT 310.950 300.600 313.050 301.050 ;
        RECT 187.950 299.400 195.600 300.600 ;
        RECT 187.950 298.950 190.050 299.400 ;
        RECT 16.950 297.600 19.050 298.050 ;
        RECT 22.950 297.600 25.050 298.050 ;
        RECT 16.950 296.400 25.050 297.600 ;
        RECT 16.950 295.950 19.050 296.400 ;
        RECT 22.950 295.950 25.050 296.400 ;
        RECT 151.950 297.600 154.050 298.050 ;
        RECT 172.950 297.600 175.050 298.050 ;
        RECT 151.950 296.400 175.050 297.600 ;
        RECT 151.950 295.950 154.050 296.400 ;
        RECT 172.950 295.950 175.050 296.400 ;
        RECT 4.950 294.750 7.050 295.200 ;
        RECT 10.950 294.750 13.050 295.200 ;
        RECT 4.950 294.600 13.050 294.750 ;
        RECT 31.950 294.600 34.050 295.200 ;
        RECT 4.950 293.550 34.050 294.600 ;
        RECT 4.950 293.100 7.050 293.550 ;
        RECT 10.950 293.400 34.050 293.550 ;
        RECT 10.950 293.100 13.050 293.400 ;
        RECT 31.950 293.100 34.050 293.400 ;
        RECT 37.950 294.600 40.050 295.200 ;
        RECT 55.950 294.600 58.050 295.200 ;
        RECT 60.000 294.600 63.900 295.050 ;
        RECT 37.950 293.400 58.050 294.600 ;
        RECT 37.950 293.100 40.050 293.400 ;
        RECT 55.950 293.100 58.050 293.400 ;
        RECT 59.400 292.950 63.900 294.600 ;
        RECT 64.950 294.600 67.050 295.050 ;
        RECT 70.950 294.600 73.050 295.200 ;
        RECT 85.950 294.600 88.050 295.200 ;
        RECT 64.950 293.400 88.050 294.600 ;
        RECT 64.950 292.950 67.050 293.400 ;
        RECT 70.950 293.100 73.050 293.400 ;
        RECT 85.950 293.100 88.050 293.400 ;
        RECT 91.950 294.750 94.050 295.200 ;
        RECT 100.950 294.750 103.050 295.200 ;
        RECT 91.950 293.550 103.050 294.750 ;
        RECT 91.950 293.100 94.050 293.550 ;
        RECT 100.950 293.100 103.050 293.550 ;
        RECT 106.950 293.100 109.050 295.200 ;
        RECT 112.950 293.100 115.050 295.200 ;
        RECT 157.950 294.750 160.050 295.200 ;
        RECT 163.950 294.750 166.050 295.200 ;
        RECT 157.950 293.550 166.050 294.750 ;
        RECT 157.950 293.100 160.050 293.550 ;
        RECT 163.950 293.100 166.050 293.550 ;
        RECT 172.950 294.600 175.050 295.200 ;
        RECT 190.950 294.600 193.050 295.200 ;
        RECT 172.950 293.400 193.050 294.600 ;
        RECT 172.950 293.100 175.050 293.400 ;
        RECT 190.950 293.100 193.050 293.400 ;
        RECT 59.400 288.900 60.600 292.950 ;
        RECT 107.400 289.050 108.600 293.100 ;
        RECT 113.400 291.600 114.600 293.100 ;
        RECT 113.400 290.400 141.600 291.600 ;
        RECT 58.950 286.800 61.050 288.900 ;
        RECT 73.950 288.450 76.050 288.900 ;
        RECT 79.950 288.450 82.050 288.900 ;
        RECT 73.950 287.250 82.050 288.450 ;
        RECT 73.950 286.800 76.050 287.250 ;
        RECT 79.950 286.800 82.050 287.250 ;
        RECT 103.950 287.400 108.600 289.050 ;
        RECT 121.950 288.600 124.050 289.050 ;
        RECT 136.950 288.600 139.050 288.900 ;
        RECT 121.950 287.400 139.050 288.600 ;
        RECT 140.400 288.600 141.600 290.400 ;
        RECT 194.400 288.900 195.600 299.400 ;
        RECT 295.950 299.400 313.050 300.600 ;
        RECT 295.950 298.950 298.050 299.400 ;
        RECT 310.950 298.950 313.050 299.400 ;
        RECT 409.950 300.600 412.050 301.050 ;
        RECT 460.950 300.600 463.050 301.050 ;
        RECT 604.950 300.600 607.050 301.050 ;
        RECT 409.950 299.400 463.050 300.600 ;
        RECT 409.950 298.950 412.050 299.400 ;
        RECT 460.950 298.950 463.050 299.400 ;
        RECT 563.400 299.400 607.050 300.600 ;
        RECT 250.950 297.600 255.000 298.050 ;
        RECT 258.000 297.600 262.050 298.050 ;
        RECT 250.950 295.950 255.600 297.600 ;
        RECT 196.950 293.100 199.050 295.200 ;
        RECT 211.950 293.100 214.050 295.200 ;
        RECT 217.950 294.750 220.050 295.200 ;
        RECT 223.950 294.750 226.050 295.200 ;
        RECT 217.950 293.550 226.050 294.750 ;
        RECT 247.950 294.600 250.050 295.200 ;
        RECT 217.950 293.100 220.050 293.550 ;
        RECT 223.950 293.100 226.050 293.550 ;
        RECT 239.400 293.400 250.050 294.600 ;
        RECT 197.400 291.600 198.600 293.100 ;
        RECT 202.950 291.600 205.050 292.050 ;
        RECT 197.400 290.400 205.050 291.600 ;
        RECT 202.950 289.950 205.050 290.400 ;
        RECT 148.950 288.600 151.050 288.900 ;
        RECT 140.400 287.400 151.050 288.600 ;
        RECT 103.950 286.950 108.000 287.400 ;
        RECT 121.950 286.950 124.050 287.400 ;
        RECT 136.950 286.800 139.050 287.400 ;
        RECT 148.950 286.800 151.050 287.400 ;
        RECT 193.950 286.800 196.050 288.900 ;
        RECT 1.950 285.600 4.050 286.050 ;
        RECT 19.950 285.600 22.050 286.050 ;
        RECT 1.950 284.400 22.050 285.600 ;
        RECT 1.950 283.950 4.050 284.400 ;
        RECT 19.950 283.950 22.050 284.400 ;
        RECT 28.950 285.600 31.050 286.050 ;
        RECT 40.950 285.600 43.050 286.050 ;
        RECT 46.950 285.600 49.050 286.050 ;
        RECT 28.950 284.400 49.050 285.600 ;
        RECT 28.950 283.950 31.050 284.400 ;
        RECT 40.950 283.950 43.050 284.400 ;
        RECT 46.950 283.950 49.050 284.400 ;
        RECT 115.950 285.600 118.050 286.050 ;
        RECT 130.950 285.600 133.050 286.050 ;
        RECT 115.950 284.400 133.050 285.600 ;
        RECT 115.950 283.950 118.050 284.400 ;
        RECT 130.950 283.950 133.050 284.400 ;
        RECT 142.950 285.600 145.050 286.050 ;
        RECT 154.950 285.600 157.050 286.050 ;
        RECT 142.950 284.400 157.050 285.600 ;
        RECT 142.950 283.950 145.050 284.400 ;
        RECT 154.950 283.950 157.050 284.400 ;
        RECT 196.950 285.600 199.050 286.050 ;
        RECT 212.400 285.600 213.600 293.100 ;
        RECT 239.400 289.050 240.600 293.400 ;
        RECT 247.950 293.100 250.050 293.400 ;
        RECT 238.950 286.950 241.050 289.050 ;
        RECT 250.950 288.600 253.050 288.900 ;
        RECT 254.400 288.600 255.600 295.950 ;
        RECT 257.400 295.950 262.050 297.600 ;
        RECT 286.950 295.950 289.050 298.050 ;
        RECT 397.950 297.600 400.050 298.050 ;
        RECT 520.950 297.600 523.050 298.050 ;
        RECT 547.950 297.600 550.050 298.050 ;
        RECT 563.400 297.600 564.600 299.400 ;
        RECT 604.950 298.950 607.050 299.400 ;
        RECT 616.950 300.600 619.050 301.050 ;
        RECT 655.950 300.600 658.050 301.050 ;
        RECT 616.950 299.400 658.050 300.600 ;
        RECT 616.950 298.950 619.050 299.400 ;
        RECT 655.950 298.950 658.050 299.400 ;
        RECT 700.950 300.600 703.050 301.050 ;
        RECT 718.950 300.600 721.050 301.050 ;
        RECT 700.950 299.400 721.050 300.600 ;
        RECT 700.950 298.950 703.050 299.400 ;
        RECT 718.950 298.950 721.050 299.400 ;
        RECT 757.950 300.600 760.050 301.050 ;
        RECT 784.950 300.600 787.050 301.050 ;
        RECT 757.950 299.400 787.050 300.600 ;
        RECT 757.950 298.950 760.050 299.400 ;
        RECT 784.950 298.950 787.050 299.400 ;
        RECT 397.950 296.400 414.600 297.600 ;
        RECT 397.950 295.950 400.050 296.400 ;
        RECT 257.400 288.900 258.600 295.950 ;
        RECT 274.950 294.750 277.050 295.200 ;
        RECT 280.950 294.750 283.050 295.200 ;
        RECT 274.950 293.550 283.050 294.750 ;
        RECT 274.950 293.100 277.050 293.550 ;
        RECT 280.950 293.100 283.050 293.550 ;
        RECT 250.950 287.400 255.600 288.600 ;
        RECT 250.950 286.800 253.050 287.400 ;
        RECT 256.950 286.800 259.050 288.900 ;
        RECT 262.950 288.450 265.050 288.900 ;
        RECT 271.950 288.450 274.050 288.900 ;
        RECT 262.950 287.250 274.050 288.450 ;
        RECT 262.950 286.800 265.050 287.250 ;
        RECT 271.950 286.800 274.050 287.250 ;
        RECT 287.400 286.050 288.600 295.950 ;
        RECT 343.950 292.950 346.050 295.050 ;
        RECT 394.950 293.100 397.050 295.200 ;
        RECT 413.400 294.600 414.600 296.400 ;
        RECT 520.950 296.400 564.600 297.600 ;
        RECT 766.950 297.600 769.050 298.050 ;
        RECT 799.950 297.600 802.050 298.050 ;
        RECT 766.950 296.400 802.050 297.600 ;
        RECT 520.950 295.950 523.050 296.400 ;
        RECT 547.950 295.950 550.050 296.400 ;
        RECT 766.950 295.950 769.050 296.400 ;
        RECT 799.950 295.950 802.050 296.400 ;
        RECT 829.950 297.600 832.050 298.050 ;
        RECT 856.950 297.600 859.050 298.050 ;
        RECT 829.950 296.400 859.050 297.600 ;
        RECT 829.950 295.950 832.050 296.400 ;
        RECT 856.950 295.950 859.050 296.400 ;
        RECT 415.950 294.600 418.050 295.200 ;
        RECT 413.400 293.400 418.050 294.600 ;
        RECT 415.950 293.100 418.050 293.400 ;
        RECT 304.950 288.600 307.050 289.050 ;
        RECT 331.950 288.600 334.050 288.900 ;
        RECT 304.950 287.400 334.050 288.600 ;
        RECT 304.950 286.950 307.050 287.400 ;
        RECT 331.950 286.800 334.050 287.400 ;
        RECT 344.400 286.050 345.600 292.950 ;
        RECT 355.950 288.450 358.050 288.900 ;
        RECT 361.950 288.600 364.050 288.900 ;
        RECT 385.950 288.600 388.050 288.900 ;
        RECT 361.950 288.450 388.050 288.600 ;
        RECT 355.950 287.400 388.050 288.450 ;
        RECT 395.400 288.600 396.600 293.100 ;
        RECT 457.950 291.600 460.050 295.050 ;
        RECT 469.950 294.600 472.050 295.200 ;
        RECT 469.950 293.400 480.600 294.600 ;
        RECT 469.950 293.100 472.050 293.400 ;
        RECT 443.400 291.000 460.050 291.600 ;
        RECT 443.400 290.400 459.600 291.000 ;
        RECT 443.400 289.050 444.600 290.400 ;
        RECT 479.400 289.050 480.600 293.400 ;
        RECT 490.800 293.100 492.900 295.200 ;
        RECT 412.950 288.600 415.050 288.900 ;
        RECT 395.400 287.400 415.050 288.600 ;
        RECT 355.950 287.250 364.050 287.400 ;
        RECT 355.950 286.800 358.050 287.250 ;
        RECT 361.950 286.800 364.050 287.250 ;
        RECT 385.950 286.800 388.050 287.400 ;
        RECT 412.950 286.800 415.050 287.400 ;
        RECT 430.950 288.600 433.050 288.900 ;
        RECT 443.400 288.600 448.050 289.050 ;
        RECT 430.950 287.400 448.050 288.600 ;
        RECT 430.950 286.800 433.050 287.400 ;
        RECT 444.000 286.950 448.050 287.400 ;
        RECT 460.950 288.450 463.050 288.900 ;
        RECT 466.950 288.450 469.050 288.900 ;
        RECT 460.950 287.250 469.050 288.450 ;
        RECT 460.950 286.800 463.050 287.250 ;
        RECT 466.950 286.800 469.050 287.250 ;
        RECT 478.950 286.950 481.050 289.050 ;
        RECT 196.950 284.400 213.600 285.600 ;
        RECT 274.950 285.600 277.050 286.050 ;
        RECT 280.950 285.600 283.050 286.050 ;
        RECT 274.950 284.400 283.050 285.600 ;
        RECT 196.950 283.950 199.050 284.400 ;
        RECT 274.950 283.950 277.050 284.400 ;
        RECT 280.950 283.950 283.050 284.400 ;
        RECT 286.950 283.950 289.050 286.050 ;
        RECT 344.400 284.400 349.050 286.050 ;
        RECT 345.000 283.950 349.050 284.400 ;
        RECT 472.950 285.600 475.050 286.050 ;
        RECT 491.400 285.600 492.600 293.100 ;
        RECT 493.950 292.950 496.050 295.050 ;
        RECT 532.950 294.600 535.050 295.200 ;
        RECT 538.950 294.600 541.050 295.050 ;
        RECT 532.950 293.400 541.050 294.600 ;
        RECT 532.950 293.100 535.050 293.400 ;
        RECT 538.950 292.950 541.050 293.400 ;
        RECT 559.950 294.750 562.050 295.200 ;
        RECT 565.950 294.750 568.050 295.200 ;
        RECT 559.950 293.550 568.050 294.750 ;
        RECT 559.950 293.100 562.050 293.550 ;
        RECT 565.950 293.100 568.050 293.550 ;
        RECT 574.950 294.600 577.050 295.200 ;
        RECT 592.950 294.600 595.050 295.200 ;
        RECT 598.950 294.600 601.050 295.050 ;
        RECT 574.950 293.400 601.050 294.600 ;
        RECT 574.950 293.100 577.050 293.400 ;
        RECT 592.950 293.100 595.050 293.400 ;
        RECT 598.950 292.950 601.050 293.400 ;
        RECT 625.950 293.100 628.050 295.200 ;
        RECT 634.800 294.000 636.900 295.050 ;
        RECT 649.950 294.600 652.050 295.050 ;
        RECT 655.950 294.600 658.050 295.050 ;
        RECT 494.400 289.050 495.600 292.950 ;
        RECT 626.400 291.600 627.600 293.100 ;
        RECT 634.800 292.950 637.050 294.000 ;
        RECT 649.950 293.400 658.050 294.600 ;
        RECT 649.950 292.950 652.050 293.400 ;
        RECT 655.950 292.950 658.050 293.400 ;
        RECT 664.950 293.100 667.050 295.200 ;
        RECT 623.400 291.000 627.600 291.600 ;
        RECT 634.950 291.600 637.050 292.950 ;
        RECT 634.950 291.000 639.600 291.600 ;
        RECT 622.950 290.400 627.600 291.000 ;
        RECT 635.250 290.400 639.600 291.000 ;
        RECT 493.950 286.950 496.050 289.050 ;
        RECT 517.950 288.600 520.050 289.050 ;
        RECT 544.950 288.600 547.050 288.900 ;
        RECT 517.950 287.400 547.050 288.600 ;
        RECT 517.950 286.950 520.050 287.400 ;
        RECT 544.950 286.800 547.050 287.400 ;
        RECT 550.950 288.600 553.050 288.900 ;
        RECT 604.950 288.600 607.050 289.050 ;
        RECT 550.950 287.400 607.050 288.600 ;
        RECT 550.950 286.800 553.050 287.400 ;
        RECT 604.950 286.950 607.050 287.400 ;
        RECT 622.950 286.950 625.050 290.400 ;
        RECT 638.400 289.050 639.600 290.400 ;
        RECT 628.950 288.600 631.050 288.900 ;
        RECT 628.950 288.000 636.600 288.600 ;
        RECT 628.950 287.400 637.050 288.000 ;
        RECT 638.400 287.400 643.050 289.050 ;
        RECT 628.950 286.800 631.050 287.400 ;
        RECT 472.950 284.400 492.600 285.600 ;
        RECT 580.950 285.600 583.050 286.050 ;
        RECT 586.950 285.600 589.050 286.050 ;
        RECT 580.950 284.400 589.050 285.600 ;
        RECT 472.950 283.950 475.050 284.400 ;
        RECT 580.950 283.950 583.050 284.400 ;
        RECT 586.950 283.950 589.050 284.400 ;
        RECT 634.950 283.950 637.050 287.400 ;
        RECT 639.000 286.950 643.050 287.400 ;
        RECT 646.950 288.600 649.050 288.900 ;
        RECT 665.400 288.600 666.600 293.100 ;
        RECT 673.950 292.050 676.050 295.050 ;
        RECT 682.950 294.600 685.050 295.200 ;
        RECT 700.950 294.600 703.050 295.200 ;
        RECT 682.950 293.400 703.050 294.600 ;
        RECT 682.950 293.100 685.050 293.400 ;
        RECT 700.950 293.100 703.050 293.400 ;
        RECT 706.950 293.100 709.050 295.200 ;
        RECT 718.950 294.750 721.050 295.200 ;
        RECT 727.950 294.750 730.050 295.200 ;
        RECT 718.950 293.550 730.050 294.750 ;
        RECT 718.950 293.100 721.050 293.550 ;
        RECT 727.950 293.100 730.050 293.550 ;
        RECT 673.950 291.900 678.000 292.050 ;
        RECT 673.950 291.000 679.050 291.900 ;
        RECT 674.400 290.400 679.050 291.000 ;
        RECT 675.000 289.950 679.050 290.400 ;
        RECT 676.950 289.800 679.050 289.950 ;
        RECT 673.950 288.600 676.050 289.050 ;
        RECT 646.950 287.400 676.050 288.600 ;
        RECT 646.950 286.800 649.050 287.400 ;
        RECT 673.950 286.950 676.050 287.400 ;
        RECT 655.950 285.600 658.050 286.050 ;
        RECT 661.950 285.600 664.050 286.050 ;
        RECT 655.950 284.400 664.050 285.600 ;
        RECT 655.950 283.950 658.050 284.400 ;
        RECT 661.950 283.950 664.050 284.400 ;
        RECT 667.950 285.600 670.050 286.050 ;
        RECT 683.400 285.600 684.600 293.100 ;
        RECT 707.400 288.600 708.600 293.100 ;
        RECT 742.950 292.950 745.050 295.050 ;
        RECT 748.950 294.600 751.050 295.200 ;
        RECT 757.950 294.600 760.050 295.050 ;
        RECT 763.950 294.600 766.050 295.200 ;
        RECT 748.950 293.400 766.050 294.600 ;
        RECT 748.950 293.100 751.050 293.400 ;
        RECT 757.950 292.950 760.050 293.400 ;
        RECT 763.950 293.100 766.050 293.400 ;
        RECT 772.950 292.950 775.050 295.050 ;
        RECT 724.950 288.600 727.050 288.900 ;
        RECT 707.400 287.400 727.050 288.600 ;
        RECT 724.950 286.800 727.050 287.400 ;
        RECT 730.950 288.600 733.050 288.900 ;
        RECT 743.400 288.600 744.600 292.950 ;
        RECT 773.400 289.050 774.600 292.950 ;
        RECT 778.950 291.600 781.050 295.050 ;
        RECT 790.950 293.100 793.050 295.200 ;
        RECT 802.950 294.600 805.050 295.200 ;
        RECT 802.950 293.400 816.600 294.600 ;
        RECT 802.950 293.100 805.050 293.400 ;
        RECT 778.950 291.000 786.600 291.600 ;
        RECT 779.400 290.400 786.600 291.000 ;
        RECT 745.950 288.600 748.050 288.900 ;
        RECT 730.950 287.400 748.050 288.600 ;
        RECT 730.950 286.800 733.050 287.400 ;
        RECT 745.950 286.800 748.050 287.400 ;
        RECT 772.950 286.950 775.050 289.050 ;
        RECT 785.400 288.600 786.600 290.400 ;
        RECT 787.950 288.600 790.050 288.900 ;
        RECT 785.400 287.400 790.050 288.600 ;
        RECT 791.400 288.600 792.600 293.100 ;
        RECT 815.400 289.050 816.600 293.400 ;
        RECT 820.950 292.950 823.050 295.050 ;
        RECT 832.950 293.100 835.050 295.200 ;
        RECT 791.400 287.400 801.600 288.600 ;
        RECT 787.950 286.800 790.050 287.400 ;
        RECT 800.400 286.050 801.600 287.400 ;
        RECT 814.950 286.950 817.050 289.050 ;
        RECT 821.400 288.600 822.600 292.950 ;
        RECT 833.400 289.050 834.600 293.100 ;
        RECT 838.950 291.600 841.050 292.050 ;
        RECT 868.950 291.600 871.050 292.050 ;
        RECT 838.950 290.400 871.050 291.600 ;
        RECT 838.950 289.950 841.050 290.400 ;
        RECT 868.950 289.950 871.050 290.400 ;
        RECT 823.950 288.600 826.050 288.900 ;
        RECT 821.400 287.400 826.050 288.600 ;
        RECT 833.400 287.400 838.050 289.050 ;
        RECT 823.950 286.800 826.050 287.400 ;
        RECT 834.000 286.950 838.050 287.400 ;
        RECT 781.950 285.600 784.050 286.050 ;
        RECT 667.950 284.400 684.600 285.600 ;
        RECT 761.400 284.400 784.050 285.600 ;
        RECT 800.400 284.400 805.050 286.050 ;
        RECT 667.950 283.950 670.050 284.400 ;
        RECT 761.400 283.050 762.600 284.400 ;
        RECT 781.950 283.950 784.050 284.400 ;
        RECT 801.000 283.950 805.050 284.400 ;
        RECT 169.950 282.600 172.050 283.050 ;
        RECT 175.950 282.600 178.050 283.050 ;
        RECT 169.950 281.400 178.050 282.600 ;
        RECT 169.950 280.950 172.050 281.400 ;
        RECT 175.950 280.950 178.050 281.400 ;
        RECT 181.950 282.600 184.050 283.050 ;
        RECT 214.950 282.600 217.050 283.050 ;
        RECT 181.950 281.400 217.050 282.600 ;
        RECT 181.950 280.950 184.050 281.400 ;
        RECT 214.950 280.950 217.050 281.400 ;
        RECT 250.950 282.600 253.050 283.050 ;
        RECT 262.950 282.600 265.050 283.050 ;
        RECT 250.950 281.400 265.050 282.600 ;
        RECT 250.950 280.950 253.050 281.400 ;
        RECT 262.950 280.950 265.050 281.400 ;
        RECT 385.950 282.600 388.050 283.050 ;
        RECT 391.950 282.600 394.050 283.050 ;
        RECT 385.950 281.400 394.050 282.600 ;
        RECT 385.950 280.950 388.050 281.400 ;
        RECT 391.950 280.950 394.050 281.400 ;
        RECT 472.950 282.600 475.050 282.900 ;
        RECT 490.950 282.600 493.050 283.050 ;
        RECT 472.950 281.400 493.050 282.600 ;
        RECT 472.950 280.800 475.050 281.400 ;
        RECT 490.950 280.950 493.050 281.400 ;
        RECT 508.950 282.600 511.050 283.050 ;
        RECT 535.950 282.600 538.050 282.900 ;
        RECT 508.950 281.400 538.050 282.600 ;
        RECT 508.950 280.950 511.050 281.400 ;
        RECT 535.950 280.800 538.050 281.400 ;
        RECT 544.950 282.600 547.050 283.050 ;
        RECT 562.950 282.600 565.050 283.050 ;
        RECT 544.950 281.400 565.050 282.600 ;
        RECT 544.950 280.950 547.050 281.400 ;
        RECT 562.950 280.950 565.050 281.400 ;
        RECT 616.950 282.600 619.050 283.050 ;
        RECT 670.950 282.600 673.050 283.050 ;
        RECT 616.950 281.400 673.050 282.600 ;
        RECT 616.950 280.950 619.050 281.400 ;
        RECT 670.950 280.950 673.050 281.400 ;
        RECT 676.950 282.600 679.050 283.050 ;
        RECT 682.950 282.600 685.050 283.050 ;
        RECT 676.950 281.400 685.050 282.600 ;
        RECT 676.950 280.950 679.050 281.400 ;
        RECT 682.950 280.950 685.050 281.400 ;
        RECT 703.950 282.600 706.050 283.050 ;
        RECT 715.950 282.600 718.050 283.050 ;
        RECT 760.950 282.600 763.050 283.050 ;
        RECT 703.950 281.400 718.050 282.600 ;
        RECT 703.950 280.950 706.050 281.400 ;
        RECT 715.950 280.950 718.050 281.400 ;
        RECT 722.400 281.400 763.050 282.600 ;
        RECT 13.950 279.600 16.050 280.050 ;
        RECT 31.950 279.600 34.050 280.050 ;
        RECT 13.950 278.400 34.050 279.600 ;
        RECT 13.950 277.950 16.050 278.400 ;
        RECT 31.950 277.950 34.050 278.400 ;
        RECT 43.950 279.600 46.050 280.050 ;
        RECT 100.950 279.600 103.050 280.050 ;
        RECT 142.950 279.600 145.050 280.050 ;
        RECT 43.950 278.400 145.050 279.600 ;
        RECT 43.950 277.950 46.050 278.400 ;
        RECT 100.950 277.950 103.050 278.400 ;
        RECT 142.950 277.950 145.050 278.400 ;
        RECT 211.950 279.600 214.050 280.050 ;
        RECT 220.950 279.600 223.050 280.050 ;
        RECT 211.950 278.400 223.050 279.600 ;
        RECT 211.950 277.950 214.050 278.400 ;
        RECT 220.950 277.950 223.050 278.400 ;
        RECT 283.950 279.600 286.050 280.050 ;
        RECT 334.950 279.600 337.050 280.050 ;
        RECT 283.950 278.400 337.050 279.600 ;
        RECT 283.950 277.950 286.050 278.400 ;
        RECT 334.950 277.950 337.050 278.400 ;
        RECT 349.950 279.600 352.050 280.050 ;
        RECT 364.950 279.600 367.050 280.050 ;
        RECT 349.950 278.400 367.050 279.600 ;
        RECT 349.950 277.950 352.050 278.400 ;
        RECT 364.950 277.950 367.050 278.400 ;
        RECT 418.950 279.600 421.050 280.050 ;
        RECT 457.950 279.600 460.050 280.050 ;
        RECT 418.950 278.400 460.050 279.600 ;
        RECT 418.950 277.950 421.050 278.400 ;
        RECT 457.950 277.950 460.050 278.400 ;
        RECT 541.950 279.600 544.050 280.050 ;
        RECT 556.950 279.600 559.050 280.050 ;
        RECT 541.950 278.400 559.050 279.600 ;
        RECT 541.950 277.950 544.050 278.400 ;
        RECT 556.950 277.950 559.050 278.400 ;
        RECT 580.950 279.600 583.050 280.050 ;
        RECT 619.950 279.600 622.050 280.050 ;
        RECT 580.950 278.400 622.050 279.600 ;
        RECT 580.950 277.950 583.050 278.400 ;
        RECT 619.950 277.950 622.050 278.400 ;
        RECT 709.950 279.600 712.050 280.050 ;
        RECT 722.400 279.600 723.600 281.400 ;
        RECT 760.950 280.950 763.050 281.400 ;
        RECT 784.950 282.600 787.050 283.050 ;
        RECT 796.950 282.600 799.050 283.050 ;
        RECT 784.950 281.400 799.050 282.600 ;
        RECT 784.950 280.950 787.050 281.400 ;
        RECT 796.950 280.950 799.050 281.400 ;
        RECT 709.950 278.400 723.600 279.600 ;
        RECT 763.950 279.600 766.050 280.050 ;
        RECT 772.950 279.600 775.050 280.050 ;
        RECT 763.950 278.400 775.050 279.600 ;
        RECT 709.950 277.950 712.050 278.400 ;
        RECT 763.950 277.950 766.050 278.400 ;
        RECT 772.950 277.950 775.050 278.400 ;
        RECT 799.950 279.600 802.050 280.050 ;
        RECT 805.950 279.600 808.050 280.050 ;
        RECT 799.950 278.400 808.050 279.600 ;
        RECT 799.950 277.950 802.050 278.400 ;
        RECT 805.950 277.950 808.050 278.400 ;
        RECT 847.950 279.600 850.050 280.050 ;
        RECT 871.950 279.600 874.050 280.050 ;
        RECT 847.950 278.400 874.050 279.600 ;
        RECT 847.950 277.950 850.050 278.400 ;
        RECT 871.950 277.950 874.050 278.400 ;
        RECT 55.950 276.600 58.050 277.050 ;
        RECT 73.950 276.600 76.050 277.050 ;
        RECT 55.950 275.400 76.050 276.600 ;
        RECT 55.950 274.950 58.050 275.400 ;
        RECT 73.950 274.950 76.050 275.400 ;
        RECT 163.950 276.600 166.050 277.050 ;
        RECT 181.950 276.600 184.050 277.050 ;
        RECT 163.950 275.400 184.050 276.600 ;
        RECT 163.950 274.950 166.050 275.400 ;
        RECT 181.950 274.950 184.050 275.400 ;
        RECT 190.950 276.600 193.050 277.050 ;
        RECT 202.950 276.600 205.050 277.050 ;
        RECT 232.950 276.600 235.050 277.050 ;
        RECT 190.950 275.400 235.050 276.600 ;
        RECT 190.950 274.950 193.050 275.400 ;
        RECT 202.950 274.950 205.050 275.400 ;
        RECT 232.950 274.950 235.050 275.400 ;
        RECT 238.950 276.600 241.050 277.050 ;
        RECT 247.950 276.600 250.050 277.050 ;
        RECT 238.950 275.400 250.050 276.600 ;
        RECT 238.950 274.950 241.050 275.400 ;
        RECT 247.950 274.950 250.050 275.400 ;
        RECT 427.950 276.600 430.050 277.050 ;
        RECT 442.950 276.600 445.050 277.050 ;
        RECT 427.950 275.400 445.050 276.600 ;
        RECT 427.950 274.950 430.050 275.400 ;
        RECT 442.950 274.950 445.050 275.400 ;
        RECT 481.950 276.600 484.050 277.050 ;
        RECT 514.950 276.600 517.050 277.050 ;
        RECT 481.950 275.400 517.050 276.600 ;
        RECT 481.950 274.950 484.050 275.400 ;
        RECT 514.950 274.950 517.050 275.400 ;
        RECT 568.950 276.600 571.050 277.050 ;
        RECT 616.950 276.600 619.050 277.050 ;
        RECT 568.950 275.400 619.050 276.600 ;
        RECT 568.950 274.950 571.050 275.400 ;
        RECT 616.950 274.950 619.050 275.400 ;
        RECT 637.950 276.600 640.050 276.900 ;
        RECT 661.950 276.600 664.050 277.050 ;
        RECT 637.950 275.400 664.050 276.600 ;
        RECT 637.950 274.800 640.050 275.400 ;
        RECT 661.950 274.950 664.050 275.400 ;
        RECT 730.950 276.600 733.050 277.050 ;
        RECT 811.950 276.600 814.050 277.050 ;
        RECT 817.950 276.600 820.050 277.050 ;
        RECT 829.950 276.600 832.050 277.050 ;
        RECT 730.950 275.400 780.600 276.600 ;
        RECT 730.950 274.950 733.050 275.400 ;
        RECT 61.950 273.600 64.050 274.050 ;
        RECT 70.950 273.600 73.050 274.050 ;
        RECT 88.800 273.600 90.900 274.050 ;
        RECT 61.950 272.400 90.900 273.600 ;
        RECT 61.950 271.950 64.050 272.400 ;
        RECT 70.950 271.950 73.050 272.400 ;
        RECT 88.800 271.950 90.900 272.400 ;
        RECT 91.950 273.600 94.050 274.050 ;
        RECT 103.950 273.600 106.050 274.050 ;
        RECT 91.950 272.400 106.050 273.600 ;
        RECT 91.950 271.950 94.050 272.400 ;
        RECT 103.950 271.950 106.050 272.400 ;
        RECT 223.950 273.600 226.050 274.050 ;
        RECT 292.950 273.600 295.050 274.050 ;
        RECT 223.950 272.400 295.050 273.600 ;
        RECT 223.950 271.950 226.050 272.400 ;
        RECT 292.950 271.950 295.050 272.400 ;
        RECT 370.950 273.600 373.050 274.050 ;
        RECT 376.950 273.600 379.050 274.050 ;
        RECT 370.950 272.400 379.050 273.600 ;
        RECT 370.950 271.950 373.050 272.400 ;
        RECT 376.950 271.950 379.050 272.400 ;
        RECT 457.950 273.600 460.050 274.050 ;
        RECT 478.950 273.600 481.050 274.050 ;
        RECT 457.950 272.400 481.050 273.600 ;
        RECT 457.950 271.950 460.050 272.400 ;
        RECT 478.950 271.950 481.050 272.400 ;
        RECT 484.950 273.600 487.050 274.050 ;
        RECT 499.950 273.600 502.050 274.050 ;
        RECT 484.950 272.400 502.050 273.600 ;
        RECT 484.950 271.950 487.050 272.400 ;
        RECT 499.950 271.950 502.050 272.400 ;
        RECT 556.950 273.600 559.050 274.050 ;
        RECT 583.950 273.600 586.050 274.050 ;
        RECT 556.950 272.400 586.050 273.600 ;
        RECT 556.950 271.950 559.050 272.400 ;
        RECT 583.950 271.950 586.050 272.400 ;
        RECT 619.950 273.600 622.050 274.050 ;
        RECT 643.950 273.600 646.050 274.050 ;
        RECT 619.950 272.400 646.050 273.600 ;
        RECT 619.950 271.950 622.050 272.400 ;
        RECT 643.950 271.950 646.050 272.400 ;
        RECT 742.950 273.600 745.050 274.050 ;
        RECT 766.950 273.600 769.050 274.050 ;
        RECT 742.950 272.400 769.050 273.600 ;
        RECT 779.400 273.600 780.600 275.400 ;
        RECT 811.950 275.400 832.050 276.600 ;
        RECT 811.950 274.950 814.050 275.400 ;
        RECT 817.950 274.950 820.050 275.400 ;
        RECT 829.950 274.950 832.050 275.400 ;
        RECT 799.950 273.600 802.050 274.050 ;
        RECT 779.400 272.400 802.050 273.600 ;
        RECT 742.950 271.950 745.050 272.400 ;
        RECT 766.950 271.950 769.050 272.400 ;
        RECT 799.950 271.950 802.050 272.400 ;
        RECT 805.950 273.600 808.050 274.050 ;
        RECT 811.950 273.600 814.050 273.900 ;
        RECT 805.950 272.400 814.050 273.600 ;
        RECT 805.950 271.950 808.050 272.400 ;
        RECT 811.950 271.800 814.050 272.400 ;
        RECT 835.950 273.600 838.050 274.050 ;
        RECT 847.950 273.600 850.050 274.050 ;
        RECT 835.950 272.400 850.050 273.600 ;
        RECT 835.950 271.950 838.050 272.400 ;
        RECT 847.950 271.950 850.050 272.400 ;
        RECT 64.950 270.600 67.050 271.050 ;
        RECT 127.950 270.600 130.050 271.050 ;
        RECT 64.950 269.400 130.050 270.600 ;
        RECT 64.950 268.950 67.050 269.400 ;
        RECT 127.950 268.950 130.050 269.400 ;
        RECT 187.950 270.600 190.050 271.050 ;
        RECT 193.950 270.600 196.050 271.050 ;
        RECT 244.950 270.600 247.050 271.050 ;
        RECT 352.950 270.600 355.050 271.050 ;
        RECT 187.950 269.400 247.050 270.600 ;
        RECT 187.950 268.950 190.050 269.400 ;
        RECT 193.950 268.950 196.050 269.400 ;
        RECT 244.950 268.950 247.050 269.400 ;
        RECT 338.400 269.400 355.050 270.600 ;
        RECT 88.950 267.600 91.050 268.050 ;
        RECT 97.950 267.600 100.050 268.050 ;
        RECT 88.950 266.400 100.050 267.600 ;
        RECT 88.950 265.950 91.050 266.400 ;
        RECT 97.950 265.950 100.050 266.400 ;
        RECT 133.950 267.600 136.050 268.050 ;
        RECT 148.950 267.600 151.050 268.050 ;
        RECT 319.950 267.600 322.050 268.050 ;
        RECT 133.950 266.400 151.050 267.600 ;
        RECT 133.950 265.950 136.050 266.400 ;
        RECT 148.950 265.950 151.050 266.400 ;
        RECT 266.400 266.400 322.050 267.600 ;
        RECT 52.950 264.600 55.050 265.050 ;
        RECT 64.950 264.600 67.050 265.050 ;
        RECT 52.950 263.400 67.050 264.600 ;
        RECT 52.950 262.950 55.050 263.400 ;
        RECT 64.950 262.950 67.050 263.400 ;
        RECT 196.950 264.600 199.050 265.050 ;
        RECT 220.950 264.600 223.050 265.050 ;
        RECT 196.950 263.400 223.050 264.600 ;
        RECT 196.950 262.950 199.050 263.400 ;
        RECT 220.950 262.950 223.050 263.400 ;
        RECT 253.950 264.600 256.050 265.050 ;
        RECT 266.400 264.600 267.600 266.400 ;
        RECT 319.950 265.950 322.050 266.400 ;
        RECT 325.950 267.600 328.050 268.050 ;
        RECT 338.400 267.600 339.600 269.400 ;
        RECT 352.950 268.950 355.050 269.400 ;
        RECT 421.950 270.600 424.050 271.050 ;
        RECT 442.950 270.600 445.050 271.050 ;
        RECT 421.950 269.400 445.050 270.600 ;
        RECT 421.950 268.950 424.050 269.400 ;
        RECT 442.950 268.950 445.050 269.400 ;
        RECT 502.950 270.600 505.050 271.050 ;
        RECT 532.800 270.600 534.900 271.050 ;
        RECT 502.950 269.400 534.900 270.600 ;
        RECT 502.950 268.950 505.050 269.400 ;
        RECT 532.800 268.950 534.900 269.400 ;
        RECT 535.950 270.600 538.050 271.050 ;
        RECT 547.950 270.600 550.050 271.050 ;
        RECT 535.950 269.400 550.050 270.600 ;
        RECT 535.950 268.950 538.050 269.400 ;
        RECT 547.950 268.950 550.050 269.400 ;
        RECT 556.950 270.600 559.050 270.900 ;
        RECT 565.950 270.600 568.050 271.050 ;
        RECT 724.950 270.600 727.050 271.050 ;
        RECT 556.950 269.400 568.050 270.600 ;
        RECT 556.950 268.800 559.050 269.400 ;
        RECT 565.950 268.950 568.050 269.400 ;
        RECT 713.400 269.400 727.050 270.600 ;
        RECT 713.400 268.050 714.600 269.400 ;
        RECT 724.950 268.950 727.050 269.400 ;
        RECT 757.950 270.600 760.050 271.050 ;
        RECT 787.950 270.600 790.050 271.050 ;
        RECT 757.950 269.400 790.050 270.600 ;
        RECT 757.950 268.950 760.050 269.400 ;
        RECT 787.950 268.950 790.050 269.400 ;
        RECT 793.950 270.600 796.050 271.050 ;
        RECT 829.950 270.600 832.050 271.050 ;
        RECT 793.950 269.400 832.050 270.600 ;
        RECT 793.950 268.950 796.050 269.400 ;
        RECT 829.950 268.950 832.050 269.400 ;
        RECT 325.950 266.400 339.600 267.600 ;
        RECT 340.950 267.600 343.050 268.050 ;
        RECT 391.950 267.600 394.050 268.050 ;
        RECT 340.950 266.400 394.050 267.600 ;
        RECT 325.950 265.950 328.050 266.400 ;
        RECT 340.950 265.950 343.050 266.400 ;
        RECT 391.950 265.950 394.050 266.400 ;
        RECT 493.950 267.600 496.050 268.050 ;
        RECT 505.950 267.600 508.050 268.050 ;
        RECT 493.950 266.400 508.050 267.600 ;
        RECT 493.950 265.950 496.050 266.400 ;
        RECT 505.950 265.950 508.050 266.400 ;
        RECT 598.950 267.600 601.050 268.050 ;
        RECT 619.950 267.600 622.050 268.050 ;
        RECT 598.950 266.400 622.050 267.600 ;
        RECT 598.950 265.950 601.050 266.400 ;
        RECT 619.950 265.950 622.050 266.400 ;
        RECT 253.950 263.400 267.600 264.600 ;
        RECT 253.950 262.950 256.050 263.400 ;
        RECT 337.950 262.950 340.050 265.050 ;
        RECT 400.950 264.600 403.050 265.050 ;
        RECT 400.950 263.400 417.600 264.600 ;
        RECT 400.950 262.950 403.050 263.400 ;
        RECT 7.950 261.750 10.050 262.200 ;
        RECT 25.950 261.750 28.050 262.200 ;
        RECT 7.950 260.550 28.050 261.750 ;
        RECT 7.950 260.100 10.050 260.550 ;
        RECT 25.950 260.100 28.050 260.550 ;
        RECT 37.950 260.100 40.050 262.200 ;
        RECT 76.950 261.600 79.050 262.200 ;
        RECT 74.400 260.400 79.050 261.600 ;
        RECT 1.950 255.450 4.050 255.900 ;
        RECT 10.950 255.450 13.050 255.900 ;
        RECT 1.950 254.250 13.050 255.450 ;
        RECT 1.950 253.800 4.050 254.250 ;
        RECT 10.950 253.800 13.050 254.250 ;
        RECT 38.400 253.050 39.600 260.100 ;
        RECT 74.400 256.050 75.600 260.400 ;
        RECT 76.950 260.100 79.050 260.400 ;
        RECT 82.950 261.750 85.050 262.200 ;
        RECT 91.950 261.750 94.050 262.200 ;
        RECT 82.950 260.550 94.050 261.750 ;
        RECT 82.950 260.100 85.050 260.550 ;
        RECT 91.950 260.100 94.050 260.550 ;
        RECT 109.800 259.950 111.900 262.050 ;
        RECT 112.950 261.600 115.050 262.050 ;
        RECT 121.950 261.600 124.050 262.200 ;
        RECT 126.000 261.600 130.050 262.050 ;
        RECT 112.950 260.400 124.050 261.600 ;
        RECT 112.950 259.950 115.050 260.400 ;
        RECT 121.950 260.100 124.050 260.400 ;
        RECT 125.400 259.950 130.050 261.600 ;
        RECT 148.950 261.600 151.050 262.200 ;
        RECT 154.950 261.750 157.050 262.200 ;
        RECT 160.950 261.750 163.050 262.200 ;
        RECT 154.950 261.600 163.050 261.750 ;
        RECT 184.950 261.600 187.050 262.200 ;
        RECT 193.950 261.600 196.050 262.050 ;
        RECT 148.950 260.550 163.050 261.600 ;
        RECT 148.950 260.400 157.050 260.550 ;
        RECT 148.950 260.100 151.050 260.400 ;
        RECT 154.950 260.100 157.050 260.400 ;
        RECT 160.950 260.100 163.050 260.550 ;
        RECT 170.400 260.400 187.050 261.600 ;
        RECT 73.950 253.950 76.050 256.050 ;
        RECT 85.950 255.600 88.050 255.900 ;
        RECT 100.950 255.600 103.050 255.900 ;
        RECT 110.250 255.600 111.450 259.950 ;
        RECT 125.400 255.900 126.600 259.950 ;
        RECT 170.400 255.900 171.600 260.400 ;
        RECT 184.950 260.100 187.050 260.400 ;
        RECT 188.400 260.400 196.050 261.600 ;
        RECT 188.400 255.900 189.600 260.400 ;
        RECT 193.950 259.950 196.050 260.400 ;
        RECT 214.950 259.950 217.050 262.050 ;
        RECT 238.950 261.750 241.050 262.200 ;
        RECT 250.950 261.750 253.050 262.200 ;
        RECT 238.950 260.550 253.050 261.750 ;
        RECT 238.950 260.100 241.050 260.550 ;
        RECT 250.950 260.100 253.050 260.550 ;
        RECT 262.950 261.750 265.050 262.200 ;
        RECT 268.950 261.750 271.050 262.200 ;
        RECT 262.950 260.550 271.050 261.750 ;
        RECT 262.950 260.100 265.050 260.550 ;
        RECT 268.950 260.100 271.050 260.550 ;
        RECT 289.950 261.750 292.050 262.200 ;
        RECT 298.950 261.750 301.050 262.200 ;
        RECT 289.950 260.550 301.050 261.750 ;
        RECT 289.950 260.100 292.050 260.550 ;
        RECT 298.950 260.100 301.050 260.550 ;
        RECT 85.950 254.400 111.450 255.600 ;
        RECT 85.950 253.800 88.050 254.400 ;
        RECT 100.950 253.800 103.050 254.400 ;
        RECT 124.950 253.800 127.050 255.900 ;
        RECT 133.950 255.450 136.050 255.900 ;
        RECT 139.950 255.450 142.050 255.900 ;
        RECT 133.950 254.250 142.050 255.450 ;
        RECT 133.950 253.800 136.050 254.250 ;
        RECT 139.950 253.800 142.050 254.250 ;
        RECT 169.950 253.800 172.050 255.900 ;
        RECT 187.950 253.800 190.050 255.900 ;
        RECT 208.950 255.600 211.050 256.050 ;
        RECT 215.400 255.600 216.600 259.950 ;
        RECT 208.950 254.400 216.600 255.600 ;
        RECT 223.950 255.600 226.050 255.900 ;
        RECT 235.950 255.600 238.050 255.900 ;
        RECT 223.950 254.400 238.050 255.600 ;
        RECT 208.950 253.950 211.050 254.400 ;
        RECT 223.950 253.800 226.050 254.400 ;
        RECT 235.950 253.800 238.050 254.400 ;
        RECT 319.950 255.600 322.050 255.900 ;
        RECT 325.950 255.600 328.050 256.050 ;
        RECT 338.400 255.900 339.600 262.950 ;
        RECT 352.950 261.600 357.000 262.050 ;
        RECT 358.950 261.600 361.050 262.200 ;
        RECT 367.950 261.600 370.050 262.050 ;
        RECT 352.950 259.950 357.600 261.600 ;
        RECT 358.950 260.400 370.050 261.600 ;
        RECT 358.950 260.100 361.050 260.400 ;
        RECT 367.950 259.950 370.050 260.400 ;
        RECT 376.950 261.600 379.050 262.200 ;
        RECT 382.950 261.600 385.050 262.050 ;
        RECT 397.950 261.600 400.050 262.200 ;
        RECT 376.950 260.400 381.600 261.600 ;
        RECT 376.950 260.100 379.050 260.400 ;
        RECT 356.400 258.600 357.600 259.950 ;
        RECT 380.400 258.600 381.600 260.400 ;
        RECT 382.950 260.400 400.050 261.600 ;
        RECT 382.950 259.950 385.050 260.400 ;
        RECT 397.950 260.100 400.050 260.400 ;
        RECT 403.950 261.600 406.050 262.050 ;
        RECT 412.950 261.600 415.050 262.200 ;
        RECT 403.950 260.400 415.050 261.600 ;
        RECT 403.950 259.950 406.050 260.400 ;
        RECT 412.950 260.100 415.050 260.400 ;
        RECT 356.400 257.400 363.600 258.600 ;
        RECT 380.400 257.400 390.600 258.600 ;
        RECT 362.400 255.900 363.600 257.400 ;
        RECT 389.400 255.900 390.600 257.400 ;
        RECT 319.950 254.400 328.050 255.600 ;
        RECT 319.950 253.800 322.050 254.400 ;
        RECT 325.950 253.950 328.050 254.400 ;
        RECT 337.950 253.800 340.050 255.900 ;
        RECT 343.950 255.600 346.050 255.900 ;
        RECT 361.950 255.600 364.050 255.900 ;
        RECT 343.950 254.400 364.050 255.600 ;
        RECT 343.950 253.800 346.050 254.400 ;
        RECT 361.950 253.800 364.050 254.400 ;
        RECT 388.950 253.800 391.050 255.900 ;
        RECT 416.400 255.600 417.600 263.400 ;
        RECT 559.950 262.950 562.050 265.050 ;
        RECT 589.950 264.600 592.050 265.050 ;
        RECT 616.950 264.600 619.050 265.050 ;
        RECT 640.950 264.600 643.050 268.050 ;
        RECT 670.950 267.600 673.050 268.050 ;
        RECT 712.950 267.600 715.050 268.050 ;
        RECT 670.950 266.400 715.050 267.600 ;
        RECT 670.950 265.950 673.050 266.400 ;
        RECT 712.950 265.950 715.050 266.400 ;
        RECT 766.950 267.600 769.050 268.050 ;
        RECT 775.950 267.600 778.050 268.050 ;
        RECT 766.950 266.400 778.050 267.600 ;
        RECT 766.950 265.950 769.050 266.400 ;
        RECT 775.950 265.950 778.050 266.400 ;
        RECT 841.950 267.600 844.050 268.050 ;
        RECT 865.950 267.600 868.050 268.050 ;
        RECT 841.950 266.400 868.050 267.600 ;
        RECT 841.950 265.950 844.050 266.400 ;
        RECT 865.950 265.950 868.050 266.400 ;
        RECT 589.950 263.400 597.600 264.600 ;
        RECT 589.950 262.950 592.050 263.400 ;
        RECT 454.950 260.100 457.050 262.200 ;
        RECT 460.950 261.750 463.050 262.200 ;
        RECT 466.950 261.750 469.050 262.200 ;
        RECT 460.950 260.550 469.050 261.750 ;
        RECT 460.950 260.100 463.050 260.550 ;
        RECT 466.950 260.100 469.050 260.550 ;
        RECT 478.950 261.750 481.050 262.200 ;
        RECT 487.950 261.750 490.050 262.200 ;
        RECT 478.950 260.550 490.050 261.750 ;
        RECT 478.950 260.100 481.050 260.550 ;
        RECT 487.950 260.100 490.050 260.550 ;
        RECT 455.400 258.600 456.600 260.100 ;
        RECT 455.400 257.400 459.600 258.600 ;
        RECT 421.950 255.600 424.050 256.050 ;
        RECT 416.400 254.400 424.050 255.600 ;
        RECT 458.400 255.600 459.600 257.400 ;
        RECT 463.950 255.600 466.050 256.050 ;
        RECT 560.400 255.900 561.600 262.950 ;
        RECT 574.950 261.600 577.050 262.200 ;
        RECT 574.950 260.400 585.600 261.600 ;
        RECT 574.950 260.100 577.050 260.400 ;
        RECT 458.400 254.400 466.050 255.600 ;
        RECT 421.950 253.950 424.050 254.400 ;
        RECT 463.950 253.950 466.050 254.400 ;
        RECT 469.950 255.450 472.050 255.900 ;
        RECT 478.950 255.450 481.050 255.900 ;
        RECT 469.950 254.250 481.050 255.450 ;
        RECT 469.950 253.800 472.050 254.250 ;
        RECT 478.950 253.800 481.050 254.250 ;
        RECT 496.950 255.600 499.050 255.900 ;
        RECT 508.950 255.600 511.050 255.900 ;
        RECT 496.950 254.400 511.050 255.600 ;
        RECT 496.950 253.800 499.050 254.400 ;
        RECT 508.950 253.800 511.050 254.400 ;
        RECT 559.950 253.800 562.050 255.900 ;
        RECT 565.950 255.450 568.050 255.900 ;
        RECT 571.950 255.450 574.050 255.900 ;
        RECT 565.950 254.250 574.050 255.450 ;
        RECT 584.400 255.600 585.600 260.400 ;
        RECT 596.400 255.900 597.600 263.400 ;
        RECT 616.950 263.400 630.600 264.600 ;
        RECT 640.950 264.000 645.600 264.600 ;
        RECT 641.400 263.400 645.600 264.000 ;
        RECT 616.950 262.950 619.050 263.400 ;
        RECT 598.950 260.100 601.050 262.200 ;
        RECT 610.950 261.750 613.050 262.200 ;
        RECT 616.950 261.750 619.050 262.200 ;
        RECT 610.950 260.550 619.050 261.750 ;
        RECT 610.950 260.100 613.050 260.550 ;
        RECT 616.950 260.100 619.050 260.550 ;
        RECT 584.400 254.400 594.600 255.600 ;
        RECT 565.950 253.800 568.050 254.250 ;
        RECT 571.950 253.800 574.050 254.250 ;
        RECT 37.950 250.950 40.050 253.050 ;
        RECT 106.950 252.600 109.050 253.050 ;
        RECT 169.950 252.600 172.050 253.050 ;
        RECT 106.950 251.400 172.050 252.600 ;
        RECT 106.950 250.950 109.050 251.400 ;
        RECT 169.950 250.950 172.050 251.400 ;
        RECT 229.950 252.600 232.050 253.050 ;
        RECT 256.950 252.600 259.050 253.050 ;
        RECT 271.950 252.600 274.050 253.050 ;
        RECT 295.950 252.600 298.050 253.050 ;
        RECT 229.950 251.400 298.050 252.600 ;
        RECT 229.950 250.950 232.050 251.400 ;
        RECT 256.950 250.950 259.050 251.400 ;
        RECT 271.950 250.950 274.050 251.400 ;
        RECT 295.950 250.950 298.050 251.400 ;
        RECT 355.950 252.600 358.050 253.050 ;
        RECT 397.950 252.600 400.050 253.050 ;
        RECT 355.950 251.400 400.050 252.600 ;
        RECT 355.950 250.950 358.050 251.400 ;
        RECT 397.950 250.950 400.050 251.400 ;
        RECT 448.950 252.600 451.050 253.050 ;
        RECT 523.950 252.600 526.050 253.050 ;
        RECT 535.950 252.600 538.050 253.050 ;
        RECT 550.950 252.600 553.050 253.050 ;
        RECT 448.950 251.400 553.050 252.600 ;
        RECT 593.400 252.600 594.600 254.400 ;
        RECT 595.950 253.800 598.050 255.900 ;
        RECT 599.400 255.600 600.600 260.100 ;
        RECT 625.950 259.950 628.050 262.050 ;
        RECT 626.400 256.050 627.600 259.950 ;
        RECT 613.950 255.600 616.050 255.900 ;
        RECT 599.400 254.400 616.050 255.600 ;
        RECT 613.950 253.800 616.050 254.400 ;
        RECT 625.800 253.950 627.900 256.050 ;
        RECT 629.400 255.900 630.600 263.400 ;
        RECT 631.950 261.750 634.050 262.200 ;
        RECT 640.950 261.750 643.050 262.200 ;
        RECT 631.950 260.550 643.050 261.750 ;
        RECT 631.950 260.100 634.050 260.550 ;
        RECT 640.950 260.100 643.050 260.550 ;
        RECT 628.950 253.800 631.050 255.900 ;
        RECT 601.950 252.600 604.050 253.050 ;
        RECT 593.400 251.400 604.050 252.600 ;
        RECT 448.950 250.950 451.050 251.400 ;
        RECT 523.950 250.950 526.050 251.400 ;
        RECT 535.950 250.950 538.050 251.400 ;
        RECT 550.950 250.950 553.050 251.400 ;
        RECT 601.950 250.950 604.050 251.400 ;
        RECT 631.950 252.600 634.050 253.050 ;
        RECT 644.400 252.600 645.600 263.400 ;
        RECT 646.950 261.600 649.050 265.050 ;
        RECT 655.950 262.950 658.050 265.050 ;
        RECT 694.950 264.600 697.050 265.050 ;
        RECT 700.950 264.600 703.050 265.050 ;
        RECT 694.950 263.400 703.050 264.600 ;
        RECT 694.950 262.950 697.050 263.400 ;
        RECT 700.950 262.950 703.050 263.400 ;
        RECT 739.950 264.600 742.050 265.050 ;
        RECT 754.950 264.600 757.050 265.200 ;
        RECT 739.950 263.400 757.050 264.600 ;
        RECT 739.950 262.950 742.050 263.400 ;
        RECT 754.950 263.100 757.050 263.400 ;
        RECT 796.950 262.950 799.050 265.050 ;
        RECT 814.950 264.600 817.050 265.050 ;
        RECT 809.400 263.400 817.050 264.600 ;
        RECT 652.950 261.600 655.050 262.200 ;
        RECT 646.950 261.000 655.050 261.600 ;
        RECT 647.400 260.400 655.050 261.000 ;
        RECT 652.950 260.100 655.050 260.400 ;
        RECT 656.400 255.600 657.600 262.950 ;
        RECT 658.950 261.600 661.050 262.200 ;
        RECT 676.950 261.600 679.050 262.200 ;
        RECT 658.950 260.400 679.050 261.600 ;
        RECT 658.950 260.100 661.050 260.400 ;
        RECT 668.400 256.050 669.600 260.400 ;
        RECT 676.950 260.100 679.050 260.400 ;
        RECT 691.950 261.600 694.050 262.200 ;
        RECT 706.950 261.600 709.050 262.050 ;
        RECT 691.950 260.400 717.600 261.600 ;
        RECT 691.950 260.100 694.050 260.400 ;
        RECT 706.950 259.950 709.050 260.400 ;
        RECT 716.400 258.600 717.600 260.400 ;
        RECT 754.950 259.950 757.050 262.050 ;
        RECT 772.950 261.600 775.050 262.200 ;
        RECT 758.400 260.400 775.050 261.600 ;
        RECT 755.400 258.600 756.600 259.950 ;
        RECT 716.400 257.400 720.600 258.600 ;
        RECT 737.400 258.000 756.600 258.600 ;
        RECT 661.950 255.600 664.050 256.050 ;
        RECT 656.400 254.400 664.050 255.600 ;
        RECT 661.950 253.950 664.050 254.400 ;
        RECT 667.950 253.950 670.050 256.050 ;
        RECT 631.950 251.400 645.600 252.600 ;
        RECT 703.950 252.600 706.050 253.050 ;
        RECT 719.400 252.600 720.600 257.400 ;
        RECT 736.950 257.400 756.600 258.000 ;
        RECT 736.950 253.950 739.050 257.400 ;
        RECT 751.950 255.600 754.050 255.900 ;
        RECT 758.400 255.600 759.600 260.400 ;
        RECT 772.950 260.100 775.050 260.400 ;
        RECT 781.950 261.600 784.050 262.050 ;
        RECT 793.950 261.600 796.050 262.200 ;
        RECT 781.950 260.400 796.050 261.600 ;
        RECT 781.950 259.950 784.050 260.400 ;
        RECT 793.950 260.100 796.050 260.400 ;
        RECT 751.950 254.400 759.600 255.600 ;
        RECT 775.950 255.450 778.050 255.900 ;
        RECT 781.950 255.450 784.050 255.900 ;
        RECT 797.400 255.600 798.600 262.950 ;
        RECT 809.400 255.900 810.600 263.400 ;
        RECT 814.950 262.950 817.050 263.400 ;
        RECT 817.950 261.600 820.050 262.200 ;
        RECT 835.950 261.600 838.050 262.200 ;
        RECT 817.950 260.400 838.050 261.600 ;
        RECT 817.950 260.100 820.050 260.400 ;
        RECT 835.950 260.100 838.050 260.400 ;
        RECT 844.950 261.750 847.050 262.200 ;
        RECT 850.950 261.750 853.050 262.200 ;
        RECT 844.950 260.550 853.050 261.750 ;
        RECT 844.950 260.100 847.050 260.550 ;
        RECT 850.950 260.100 853.050 260.550 ;
        RECT 856.950 259.950 859.050 262.050 ;
        RECT 857.400 256.050 858.600 259.950 ;
        RECT 751.950 253.800 754.050 254.400 ;
        RECT 775.950 254.250 784.050 255.450 ;
        RECT 775.950 253.800 778.050 254.250 ;
        RECT 781.950 253.800 784.050 254.250 ;
        RECT 794.400 254.400 798.600 255.600 ;
        RECT 727.950 252.600 730.050 253.050 ;
        RECT 703.950 251.400 730.050 252.600 ;
        RECT 631.950 250.950 634.050 251.400 ;
        RECT 703.950 250.950 706.050 251.400 ;
        RECT 727.950 250.950 730.050 251.400 ;
        RECT 754.950 252.600 757.050 253.050 ;
        RECT 763.950 252.600 766.050 253.050 ;
        RECT 754.950 251.400 766.050 252.600 ;
        RECT 754.950 250.950 757.050 251.400 ;
        RECT 763.950 250.950 766.050 251.400 ;
        RECT 778.950 252.600 781.050 253.050 ;
        RECT 794.400 252.600 795.600 254.400 ;
        RECT 808.950 253.800 811.050 255.900 ;
        RECT 856.950 253.950 859.050 256.050 ;
        RECT 778.950 251.400 795.600 252.600 ;
        RECT 847.950 252.600 850.050 253.050 ;
        RECT 853.950 252.600 856.050 253.050 ;
        RECT 847.950 251.400 856.050 252.600 ;
        RECT 778.950 250.950 781.050 251.400 ;
        RECT 847.950 250.950 850.050 251.400 ;
        RECT 853.950 250.950 856.050 251.400 ;
        RECT 79.950 249.600 82.050 250.050 ;
        RECT 107.400 249.600 108.600 250.950 ;
        RECT 79.950 248.400 108.600 249.600 ;
        RECT 181.950 249.600 184.050 250.050 ;
        RECT 196.950 249.600 199.050 250.050 ;
        RECT 181.950 248.400 199.050 249.600 ;
        RECT 79.950 247.950 82.050 248.400 ;
        RECT 181.950 247.950 184.050 248.400 ;
        RECT 196.950 247.950 199.050 248.400 ;
        RECT 280.950 249.600 283.050 250.050 ;
        RECT 286.950 249.600 289.050 250.050 ;
        RECT 280.950 248.400 289.050 249.600 ;
        RECT 280.950 247.950 283.050 248.400 ;
        RECT 286.950 247.950 289.050 248.400 ;
        RECT 298.950 249.600 301.050 250.050 ;
        RECT 307.950 249.600 310.050 250.050 ;
        RECT 298.950 248.400 310.050 249.600 ;
        RECT 298.950 247.950 301.050 248.400 ;
        RECT 307.950 247.950 310.050 248.400 ;
        RECT 394.950 249.600 397.050 250.050 ;
        RECT 403.950 249.600 406.050 250.050 ;
        RECT 394.950 248.400 406.050 249.600 ;
        RECT 394.950 247.950 397.050 248.400 ;
        RECT 403.950 247.950 406.050 248.400 ;
        RECT 409.950 249.600 412.050 250.050 ;
        RECT 439.950 249.600 442.050 250.050 ;
        RECT 409.950 248.400 442.050 249.600 ;
        RECT 409.950 247.950 412.050 248.400 ;
        RECT 439.950 247.950 442.050 248.400 ;
        RECT 478.950 249.600 481.050 250.050 ;
        RECT 502.950 249.600 505.050 250.050 ;
        RECT 478.950 248.400 505.050 249.600 ;
        RECT 478.950 247.950 481.050 248.400 ;
        RECT 502.950 247.950 505.050 248.400 ;
        RECT 556.950 249.600 559.050 250.050 ;
        RECT 586.950 249.600 589.050 250.050 ;
        RECT 556.950 248.400 589.050 249.600 ;
        RECT 556.950 247.950 559.050 248.400 ;
        RECT 586.950 247.950 589.050 248.400 ;
        RECT 607.950 249.600 610.050 250.050 ;
        RECT 634.950 249.600 637.050 250.050 ;
        RECT 607.950 248.400 637.050 249.600 ;
        RECT 607.950 247.950 610.050 248.400 ;
        RECT 634.950 247.950 637.050 248.400 ;
        RECT 643.950 249.600 646.050 250.050 ;
        RECT 667.950 249.600 670.050 250.050 ;
        RECT 643.950 248.400 670.050 249.600 ;
        RECT 643.950 247.950 646.050 248.400 ;
        RECT 667.950 247.950 670.050 248.400 ;
        RECT 799.950 249.600 802.050 250.050 ;
        RECT 823.950 249.600 826.050 250.050 ;
        RECT 799.950 248.400 826.050 249.600 ;
        RECT 799.950 247.950 802.050 248.400 ;
        RECT 823.950 247.950 826.050 248.400 ;
        RECT 4.950 246.600 7.050 247.050 ;
        RECT 10.950 246.600 13.050 247.050 ;
        RECT 4.950 245.400 13.050 246.600 ;
        RECT 4.950 244.950 7.050 245.400 ;
        RECT 10.950 244.950 13.050 245.400 ;
        RECT 22.950 246.600 25.050 247.050 ;
        RECT 31.950 246.600 34.050 247.050 ;
        RECT 22.950 245.400 34.050 246.600 ;
        RECT 22.950 244.950 25.050 245.400 ;
        RECT 31.950 244.950 34.050 245.400 ;
        RECT 124.950 246.600 127.050 247.050 ;
        RECT 154.950 246.600 157.050 247.050 ;
        RECT 124.950 245.400 157.050 246.600 ;
        RECT 124.950 244.950 127.050 245.400 ;
        RECT 154.950 244.950 157.050 245.400 ;
        RECT 199.950 246.600 202.050 247.050 ;
        RECT 211.950 246.600 214.050 247.050 ;
        RECT 199.950 245.400 214.050 246.600 ;
        RECT 199.950 244.950 202.050 245.400 ;
        RECT 211.950 244.950 214.050 245.400 ;
        RECT 352.950 246.600 355.050 247.050 ;
        RECT 410.400 246.600 411.600 247.950 ;
        RECT 352.950 245.400 411.600 246.600 ;
        RECT 412.950 246.600 415.050 247.050 ;
        RECT 430.950 246.600 433.050 247.050 ;
        RECT 412.950 245.400 433.050 246.600 ;
        RECT 352.950 244.950 355.050 245.400 ;
        RECT 412.950 244.950 415.050 245.400 ;
        RECT 430.950 244.950 433.050 245.400 ;
        RECT 499.950 246.600 502.050 247.050 ;
        RECT 517.950 246.600 520.050 247.050 ;
        RECT 499.950 245.400 520.050 246.600 ;
        RECT 499.950 244.950 502.050 245.400 ;
        RECT 517.950 244.950 520.050 245.400 ;
        RECT 589.950 246.600 592.050 247.050 ;
        RECT 655.950 246.600 658.050 247.050 ;
        RECT 589.950 245.400 658.050 246.600 ;
        RECT 589.950 244.950 592.050 245.400 ;
        RECT 655.950 244.950 658.050 245.400 ;
        RECT 685.950 246.600 688.050 247.050 ;
        RECT 733.950 246.600 736.050 247.050 ;
        RECT 685.950 245.400 736.050 246.600 ;
        RECT 685.950 244.950 688.050 245.400 ;
        RECT 733.950 244.950 736.050 245.400 ;
        RECT 769.950 246.600 772.050 247.050 ;
        RECT 800.400 246.600 801.600 247.950 ;
        RECT 769.950 245.400 801.600 246.600 ;
        RECT 769.950 244.950 772.050 245.400 ;
        RECT 79.950 243.600 82.050 244.050 ;
        RECT 91.950 243.600 94.050 244.050 ;
        RECT 79.950 242.400 94.050 243.600 ;
        RECT 79.950 241.950 82.050 242.400 ;
        RECT 91.950 241.950 94.050 242.400 ;
        RECT 145.950 243.600 148.050 244.050 ;
        RECT 163.950 243.600 166.050 244.050 ;
        RECT 235.950 243.600 238.050 244.050 ;
        RECT 145.950 242.400 238.050 243.600 ;
        RECT 145.950 241.950 148.050 242.400 ;
        RECT 163.950 241.950 166.050 242.400 ;
        RECT 235.950 241.950 238.050 242.400 ;
        RECT 250.950 243.600 253.050 244.050 ;
        RECT 283.950 243.600 286.050 244.050 ;
        RECT 250.950 242.400 286.050 243.600 ;
        RECT 250.950 241.950 253.050 242.400 ;
        RECT 283.950 241.950 286.050 242.400 ;
        RECT 301.950 243.600 304.050 244.050 ;
        RECT 325.950 243.600 328.050 244.050 ;
        RECT 301.950 242.400 328.050 243.600 ;
        RECT 301.950 241.950 304.050 242.400 ;
        RECT 325.950 241.950 328.050 242.400 ;
        RECT 421.950 243.600 424.050 244.050 ;
        RECT 619.950 243.600 622.050 244.050 ;
        RECT 649.950 243.600 652.050 244.050 ;
        RECT 421.950 242.400 492.600 243.600 ;
        RECT 421.950 241.950 424.050 242.400 ;
        RECT 491.400 241.050 492.600 242.400 ;
        RECT 619.950 242.400 652.050 243.600 ;
        RECT 619.950 241.950 622.050 242.400 ;
        RECT 649.950 241.950 652.050 242.400 ;
        RECT 673.950 243.600 676.050 244.050 ;
        RECT 763.950 243.600 766.050 244.050 ;
        RECT 673.950 242.400 766.050 243.600 ;
        RECT 673.950 241.950 676.050 242.400 ;
        RECT 763.950 241.950 766.050 242.400 ;
        RECT 247.950 240.600 250.050 241.050 ;
        RECT 352.950 240.600 355.050 241.050 ;
        RECT 247.950 239.400 355.050 240.600 ;
        RECT 247.950 238.950 250.050 239.400 ;
        RECT 352.950 238.950 355.050 239.400 ;
        RECT 445.950 240.600 448.050 241.050 ;
        RECT 463.950 240.600 466.050 241.050 ;
        RECT 445.950 239.400 466.050 240.600 ;
        RECT 445.950 238.950 448.050 239.400 ;
        RECT 463.950 238.950 466.050 239.400 ;
        RECT 490.950 240.600 493.050 241.050 ;
        RECT 577.950 240.600 580.050 241.050 ;
        RECT 490.950 239.400 580.050 240.600 ;
        RECT 650.400 240.600 651.600 241.950 ;
        RECT 814.950 240.600 817.050 241.050 ;
        RECT 650.400 239.400 817.050 240.600 ;
        RECT 490.950 238.950 493.050 239.400 ;
        RECT 577.950 238.950 580.050 239.400 ;
        RECT 814.950 238.950 817.050 239.400 ;
        RECT 112.950 237.600 115.050 238.050 ;
        RECT 142.950 237.600 145.050 238.050 ;
        RECT 112.950 236.400 145.050 237.600 ;
        RECT 112.950 235.950 115.050 236.400 ;
        RECT 142.950 235.950 145.050 236.400 ;
        RECT 166.950 237.600 169.050 238.050 ;
        RECT 238.950 237.600 241.050 238.050 ;
        RECT 253.950 237.600 256.050 238.050 ;
        RECT 166.950 236.400 256.050 237.600 ;
        RECT 166.950 235.950 169.050 236.400 ;
        RECT 238.950 235.950 241.050 236.400 ;
        RECT 253.950 235.950 256.050 236.400 ;
        RECT 295.950 237.600 298.050 238.050 ;
        RECT 310.950 237.600 313.050 238.050 ;
        RECT 406.950 237.600 409.050 238.050 ;
        RECT 295.950 236.400 409.050 237.600 ;
        RECT 295.950 235.950 298.050 236.400 ;
        RECT 310.950 235.950 313.050 236.400 ;
        RECT 406.950 235.950 409.050 236.400 ;
        RECT 637.950 237.600 640.050 238.050 ;
        RECT 649.950 237.600 652.050 237.900 ;
        RECT 637.950 236.400 652.050 237.600 ;
        RECT 637.950 235.950 640.050 236.400 ;
        RECT 649.950 235.800 652.050 236.400 ;
        RECT 661.950 237.600 664.050 238.050 ;
        RECT 673.950 237.600 676.050 238.050 ;
        RECT 688.950 237.600 691.050 238.050 ;
        RECT 661.950 236.400 691.050 237.600 ;
        RECT 661.950 235.950 664.050 236.400 ;
        RECT 673.950 235.950 676.050 236.400 ;
        RECT 688.950 235.950 691.050 236.400 ;
        RECT 709.950 237.600 712.050 238.050 ;
        RECT 778.950 237.600 781.050 238.050 ;
        RECT 709.950 236.400 781.050 237.600 ;
        RECT 709.950 235.950 712.050 236.400 ;
        RECT 778.950 235.950 781.050 236.400 ;
        RECT 784.950 237.600 787.050 238.050 ;
        RECT 802.950 237.600 805.050 238.050 ;
        RECT 811.950 237.600 814.050 238.050 ;
        RECT 784.950 236.400 814.050 237.600 ;
        RECT 784.950 235.950 787.050 236.400 ;
        RECT 802.950 235.950 805.050 236.400 ;
        RECT 811.950 235.950 814.050 236.400 ;
        RECT 118.950 234.600 121.050 235.050 ;
        RECT 247.950 234.600 250.050 235.050 ;
        RECT 118.950 233.400 250.050 234.600 ;
        RECT 118.950 232.950 121.050 233.400 ;
        RECT 247.950 232.950 250.050 233.400 ;
        RECT 277.950 234.600 280.050 235.050 ;
        RECT 316.950 234.600 319.050 235.050 ;
        RECT 382.950 234.600 385.050 235.050 ;
        RECT 277.950 233.400 315.600 234.600 ;
        RECT 277.950 232.950 280.050 233.400 ;
        RECT 205.950 231.600 208.050 232.050 ;
        RECT 229.950 231.600 232.050 232.050 ;
        RECT 205.950 230.400 232.050 231.600 ;
        RECT 314.400 231.600 315.600 233.400 ;
        RECT 316.950 233.400 385.050 234.600 ;
        RECT 316.950 232.950 319.050 233.400 ;
        RECT 382.950 232.950 385.050 233.400 ;
        RECT 421.950 234.600 424.050 235.050 ;
        RECT 442.950 234.600 445.050 235.050 ;
        RECT 421.950 233.400 445.050 234.600 ;
        RECT 421.950 232.950 424.050 233.400 ;
        RECT 442.950 232.950 445.050 233.400 ;
        RECT 457.950 234.600 462.000 235.050 ;
        RECT 532.950 234.600 535.050 235.050 ;
        RECT 622.950 234.600 625.050 235.050 ;
        RECT 658.950 234.600 661.050 235.050 ;
        RECT 766.950 234.600 769.050 235.050 ;
        RECT 457.950 232.950 462.600 234.600 ;
        RECT 532.950 233.400 661.050 234.600 ;
        RECT 532.950 232.950 535.050 233.400 ;
        RECT 622.950 232.950 625.050 233.400 ;
        RECT 658.950 232.950 661.050 233.400 ;
        RECT 737.400 233.400 769.050 234.600 ;
        RECT 454.950 231.600 457.050 232.050 ;
        RECT 314.400 230.400 457.050 231.600 ;
        RECT 461.400 231.600 462.600 232.950 ;
        RECT 535.950 231.600 538.050 232.050 ;
        RECT 461.400 230.400 538.050 231.600 ;
        RECT 205.950 229.950 208.050 230.400 ;
        RECT 229.950 229.950 232.050 230.400 ;
        RECT 454.950 229.950 457.050 230.400 ;
        RECT 535.950 229.950 538.050 230.400 ;
        RECT 541.950 231.600 544.050 232.050 ;
        RECT 565.950 231.600 568.050 232.050 ;
        RECT 541.950 230.400 568.050 231.600 ;
        RECT 541.950 229.950 544.050 230.400 ;
        RECT 565.950 229.950 568.050 230.400 ;
        RECT 574.950 231.600 577.050 232.050 ;
        RECT 625.950 231.600 628.050 232.050 ;
        RECT 652.800 231.600 654.900 232.050 ;
        RECT 574.950 230.400 654.900 231.600 ;
        RECT 574.950 229.950 577.050 230.400 ;
        RECT 625.950 229.950 628.050 230.400 ;
        RECT 652.800 229.950 654.900 230.400 ;
        RECT 655.950 231.600 658.050 232.050 ;
        RECT 682.950 231.600 685.050 232.050 ;
        RECT 655.950 230.400 685.050 231.600 ;
        RECT 655.950 229.950 658.050 230.400 ;
        RECT 682.950 229.950 685.050 230.400 ;
        RECT 697.950 231.600 700.050 232.050 ;
        RECT 737.400 231.600 738.600 233.400 ;
        RECT 766.950 232.950 769.050 233.400 ;
        RECT 832.950 234.600 835.050 235.050 ;
        RECT 868.950 234.600 871.050 235.050 ;
        RECT 832.950 233.400 871.050 234.600 ;
        RECT 832.950 232.950 835.050 233.400 ;
        RECT 868.950 232.950 871.050 233.400 ;
        RECT 697.950 230.400 738.600 231.600 ;
        RECT 742.950 231.600 745.050 232.050 ;
        RECT 829.950 231.600 832.050 232.050 ;
        RECT 742.950 230.400 832.050 231.600 ;
        RECT 697.950 229.950 700.050 230.400 ;
        RECT 742.950 229.950 745.050 230.400 ;
        RECT 829.950 229.950 832.050 230.400 ;
        RECT 88.950 228.600 91.050 229.050 ;
        RECT 190.950 228.600 193.050 229.050 ;
        RECT 406.950 228.600 409.050 229.050 ;
        RECT 427.950 228.600 430.050 229.050 ;
        RECT 457.950 228.600 460.050 229.050 ;
        RECT 88.950 227.400 138.600 228.600 ;
        RECT 88.950 226.950 91.050 227.400 ;
        RECT 137.400 226.050 138.600 227.400 ;
        RECT 190.950 227.400 219.600 228.600 ;
        RECT 190.950 226.950 193.050 227.400 ;
        RECT 218.400 226.050 219.600 227.400 ;
        RECT 406.950 227.400 460.050 228.600 ;
        RECT 406.950 226.950 409.050 227.400 ;
        RECT 427.950 226.950 430.050 227.400 ;
        RECT 457.950 226.950 460.050 227.400 ;
        RECT 466.950 228.600 469.050 229.050 ;
        RECT 604.950 228.600 607.050 229.050 ;
        RECT 643.950 228.600 646.050 229.050 ;
        RECT 466.950 227.400 646.050 228.600 ;
        RECT 466.950 226.950 469.050 227.400 ;
        RECT 604.950 226.950 607.050 227.400 ;
        RECT 643.950 226.950 646.050 227.400 ;
        RECT 661.950 228.600 664.050 229.050 ;
        RECT 691.950 228.600 694.050 229.050 ;
        RECT 661.950 227.400 694.050 228.600 ;
        RECT 661.950 226.950 664.050 227.400 ;
        RECT 691.950 226.950 694.050 227.400 ;
        RECT 10.950 225.600 13.050 226.050 ;
        RECT 43.950 225.600 46.050 226.050 ;
        RECT 10.950 224.400 46.050 225.600 ;
        RECT 10.950 223.950 13.050 224.400 ;
        RECT 43.950 223.950 46.050 224.400 ;
        RECT 136.950 225.600 139.050 226.050 ;
        RECT 160.950 225.600 163.050 226.050 ;
        RECT 136.950 224.400 163.050 225.600 ;
        RECT 136.950 223.950 139.050 224.400 ;
        RECT 160.950 223.950 163.050 224.400 ;
        RECT 217.950 225.600 220.050 226.050 ;
        RECT 265.950 225.600 268.050 226.050 ;
        RECT 304.950 225.600 307.050 225.900 ;
        RECT 217.950 224.400 307.050 225.600 ;
        RECT 217.950 223.950 220.050 224.400 ;
        RECT 265.950 223.950 268.050 224.400 ;
        RECT 304.950 223.800 307.050 224.400 ;
        RECT 400.950 225.600 403.050 226.050 ;
        RECT 418.950 225.600 421.050 226.050 ;
        RECT 400.950 224.400 421.050 225.600 ;
        RECT 400.950 223.950 403.050 224.400 ;
        RECT 418.950 223.950 421.050 224.400 ;
        RECT 430.950 225.600 433.050 226.050 ;
        RECT 448.950 225.600 451.050 226.050 ;
        RECT 430.950 224.400 451.050 225.600 ;
        RECT 430.950 223.950 433.050 224.400 ;
        RECT 448.950 223.950 451.050 224.400 ;
        RECT 505.950 225.600 508.050 226.050 ;
        RECT 532.950 225.600 535.050 226.050 ;
        RECT 505.950 224.400 535.050 225.600 ;
        RECT 505.950 223.950 508.050 224.400 ;
        RECT 532.950 223.950 535.050 224.400 ;
        RECT 655.950 225.600 658.050 226.050 ;
        RECT 709.950 225.600 712.050 226.050 ;
        RECT 655.950 224.400 712.050 225.600 ;
        RECT 655.950 223.950 658.050 224.400 ;
        RECT 709.950 223.950 712.050 224.400 ;
        RECT 829.950 225.600 832.050 226.050 ;
        RECT 859.950 225.600 862.050 226.050 ;
        RECT 829.950 224.400 862.050 225.600 ;
        RECT 829.950 223.950 832.050 224.400 ;
        RECT 859.950 223.950 862.050 224.400 ;
        RECT 64.950 222.600 67.050 223.050 ;
        RECT 70.950 222.600 73.050 223.050 ;
        RECT 64.950 221.400 73.050 222.600 ;
        RECT 64.950 220.950 67.050 221.400 ;
        RECT 70.950 220.950 73.050 221.400 ;
        RECT 112.950 222.600 115.050 223.050 ;
        RECT 121.950 222.600 124.050 223.050 ;
        RECT 151.950 222.600 154.050 223.050 ;
        RECT 112.950 221.400 154.050 222.600 ;
        RECT 112.950 220.950 115.050 221.400 ;
        RECT 121.950 220.950 124.050 221.400 ;
        RECT 151.950 220.950 154.050 221.400 ;
        RECT 172.950 222.600 175.050 223.050 ;
        RECT 196.950 222.600 199.050 223.050 ;
        RECT 172.950 221.400 199.050 222.600 ;
        RECT 172.950 220.950 175.050 221.400 ;
        RECT 196.950 220.950 199.050 221.400 ;
        RECT 211.950 222.600 214.050 223.050 ;
        RECT 232.950 222.600 235.050 223.050 ;
        RECT 244.950 222.600 247.050 223.050 ;
        RECT 268.950 222.600 271.050 223.050 ;
        RECT 286.950 222.600 289.050 223.050 ;
        RECT 211.950 221.400 231.600 222.600 ;
        RECT 211.950 220.950 214.050 221.400 ;
        RECT 230.400 219.600 231.600 221.400 ;
        RECT 232.950 221.400 247.050 222.600 ;
        RECT 232.950 220.950 235.050 221.400 ;
        RECT 244.950 220.950 247.050 221.400 ;
        RECT 254.400 221.400 289.050 222.600 ;
        RECT 254.400 219.600 255.600 221.400 ;
        RECT 268.950 220.950 271.050 221.400 ;
        RECT 286.950 220.950 289.050 221.400 ;
        RECT 295.950 222.600 298.050 223.050 ;
        RECT 358.950 222.600 361.050 223.050 ;
        RECT 295.950 221.400 361.050 222.600 ;
        RECT 295.950 220.950 298.050 221.400 ;
        RECT 358.950 220.950 361.050 221.400 ;
        RECT 439.950 222.600 442.050 223.050 ;
        RECT 451.800 222.600 453.900 223.050 ;
        RECT 439.950 221.400 453.900 222.600 ;
        RECT 439.950 220.950 442.050 221.400 ;
        RECT 451.800 220.950 453.900 221.400 ;
        RECT 454.950 222.600 457.050 223.050 ;
        RECT 466.950 222.600 469.050 223.050 ;
        RECT 454.950 221.400 469.050 222.600 ;
        RECT 454.950 220.950 457.050 221.400 ;
        RECT 466.950 220.950 469.050 221.400 ;
        RECT 472.950 222.600 475.050 223.050 ;
        RECT 493.950 222.600 496.050 223.050 ;
        RECT 502.950 222.600 505.050 223.050 ;
        RECT 472.950 221.400 505.050 222.600 ;
        RECT 472.950 220.950 475.050 221.400 ;
        RECT 493.950 220.950 496.050 221.400 ;
        RECT 502.950 220.950 505.050 221.400 ;
        RECT 550.950 222.600 553.050 223.050 ;
        RECT 580.950 222.600 583.050 223.050 ;
        RECT 550.950 221.400 583.050 222.600 ;
        RECT 550.950 220.950 553.050 221.400 ;
        RECT 580.950 220.950 583.050 221.400 ;
        RECT 613.950 222.600 616.050 223.050 ;
        RECT 631.950 222.600 634.050 223.050 ;
        RECT 613.950 221.400 634.050 222.600 ;
        RECT 613.950 220.950 616.050 221.400 ;
        RECT 631.950 220.950 634.050 221.400 ;
        RECT 670.950 222.600 673.050 223.050 ;
        RECT 694.950 222.600 697.050 223.050 ;
        RECT 670.950 221.400 697.050 222.600 ;
        RECT 670.950 220.950 673.050 221.400 ;
        RECT 694.950 220.950 697.050 221.400 ;
        RECT 700.950 222.600 703.050 223.050 ;
        RECT 712.950 222.600 715.050 223.050 ;
        RECT 700.950 221.400 715.050 222.600 ;
        RECT 700.950 220.950 703.050 221.400 ;
        RECT 712.950 220.950 715.050 221.400 ;
        RECT 772.950 222.600 775.050 223.050 ;
        RECT 820.800 222.600 822.900 223.050 ;
        RECT 772.950 221.400 822.900 222.600 ;
        RECT 772.950 220.950 775.050 221.400 ;
        RECT 820.800 220.950 822.900 221.400 ;
        RECT 230.400 218.400 255.600 219.600 ;
        RECT 289.950 217.950 292.050 220.050 ;
        RECT 319.950 219.600 322.050 220.050 ;
        RECT 328.950 219.600 331.050 220.050 ;
        RECT 319.950 218.400 331.050 219.600 ;
        RECT 319.950 217.950 322.050 218.400 ;
        RECT 328.950 217.950 331.050 218.400 ;
        RECT 373.950 217.950 376.050 220.050 ;
        RECT 394.950 219.600 397.050 220.050 ;
        RECT 415.950 219.600 418.050 220.050 ;
        RECT 430.950 219.600 433.050 220.050 ;
        RECT 394.950 218.400 433.050 219.600 ;
        RECT 394.950 217.950 397.050 218.400 ;
        RECT 415.950 217.950 418.050 218.400 ;
        RECT 430.950 217.950 433.050 218.400 ;
        RECT 535.950 219.600 538.050 220.050 ;
        RECT 547.950 219.600 550.050 220.050 ;
        RECT 535.950 218.400 550.050 219.600 ;
        RECT 535.950 217.950 538.050 218.400 ;
        RECT 547.950 217.950 550.050 218.400 ;
        RECT 649.950 219.600 652.050 219.900 ;
        RECT 691.950 219.600 694.050 220.050 ;
        RECT 706.950 219.600 709.050 220.050 ;
        RECT 649.950 218.400 681.600 219.600 ;
        RECT 16.950 216.600 19.050 217.200 ;
        RECT 31.950 216.600 34.050 217.200 ;
        RECT 49.950 216.600 52.050 217.200 ;
        RECT 16.950 215.400 27.600 216.600 ;
        RECT 16.950 215.100 19.050 215.400 ;
        RECT 26.400 211.050 27.600 215.400 ;
        RECT 31.950 215.400 52.050 216.600 ;
        RECT 31.950 215.100 34.050 215.400 ;
        RECT 49.950 215.100 52.050 215.400 ;
        RECT 94.950 215.100 97.050 217.200 ;
        RECT 106.950 215.100 109.050 217.200 ;
        RECT 95.400 211.050 96.600 215.100 ;
        RECT 107.400 211.050 108.600 215.100 ;
        RECT 124.950 214.950 127.050 217.050 ;
        RECT 130.950 215.100 133.050 217.200 ;
        RECT 184.950 215.100 187.050 217.200 ;
        RECT 247.950 215.100 250.050 217.200 ;
        RECT 253.950 215.100 256.050 217.200 ;
        RECT 259.950 216.750 262.050 217.200 ;
        RECT 265.950 216.750 268.050 217.200 ;
        RECT 259.950 215.550 268.050 216.750 ;
        RECT 259.950 215.100 262.050 215.550 ;
        RECT 265.950 215.100 268.050 215.550 ;
        RECT 271.950 216.750 274.050 217.200 ;
        RECT 277.950 216.750 280.050 217.200 ;
        RECT 271.950 215.550 280.050 216.750 ;
        RECT 271.950 215.100 274.050 215.550 ;
        RECT 277.950 215.100 280.050 215.550 ;
        RECT 125.400 211.050 126.600 214.950 ;
        RECT 1.950 210.600 4.050 211.050 ;
        RECT 13.950 210.600 16.050 210.900 ;
        RECT 1.950 209.400 16.050 210.600 ;
        RECT 1.950 208.950 4.050 209.400 ;
        RECT 13.950 208.800 16.050 209.400 ;
        RECT 25.950 208.950 28.050 211.050 ;
        RECT 58.950 210.450 61.050 210.900 ;
        RECT 73.950 210.450 76.050 210.900 ;
        RECT 58.950 209.250 76.050 210.450 ;
        RECT 58.950 208.800 61.050 209.250 ;
        RECT 73.950 208.800 76.050 209.250 ;
        RECT 79.950 210.600 82.050 211.050 ;
        RECT 85.950 210.600 88.050 210.900 ;
        RECT 79.950 209.400 88.050 210.600 ;
        RECT 95.400 209.400 100.050 211.050 ;
        RECT 79.950 208.950 82.050 209.400 ;
        RECT 85.950 208.800 88.050 209.400 ;
        RECT 96.000 208.950 100.050 209.400 ;
        RECT 103.950 209.400 108.600 211.050 ;
        RECT 103.950 208.950 108.000 209.400 ;
        RECT 124.950 208.950 127.050 211.050 ;
        RECT 131.400 208.050 132.600 215.100 ;
        RECT 185.400 211.050 186.600 215.100 ;
        RECT 181.950 209.400 186.600 211.050 ;
        RECT 208.950 210.600 211.050 210.900 ;
        RECT 188.400 209.400 211.050 210.600 ;
        RECT 181.950 208.950 186.000 209.400 ;
        RECT 127.950 206.400 132.600 208.050 ;
        RECT 148.950 207.600 151.050 208.050 ;
        RECT 163.950 207.600 166.050 208.050 ;
        RECT 169.950 207.600 172.050 208.050 ;
        RECT 148.950 206.400 172.050 207.600 ;
        RECT 127.950 205.950 132.000 206.400 ;
        RECT 148.950 205.950 151.050 206.400 ;
        RECT 163.950 205.950 166.050 206.400 ;
        RECT 169.950 205.950 172.050 206.400 ;
        RECT 178.950 207.600 181.050 208.050 ;
        RECT 188.400 207.600 189.600 209.400 ;
        RECT 208.950 208.800 211.050 209.400 ;
        RECT 229.950 210.600 232.050 210.900 ;
        RECT 248.400 210.600 249.600 215.100 ;
        RECT 229.950 209.400 249.600 210.600 ;
        RECT 254.400 210.600 255.600 215.100 ;
        RECT 290.400 213.600 291.600 217.950 ;
        RECT 310.950 215.100 313.050 217.200 ;
        RECT 331.950 216.600 334.050 217.200 ;
        RECT 331.950 215.400 336.600 216.600 ;
        RECT 331.950 215.100 334.050 215.400 ;
        RECT 284.400 212.400 291.600 213.600 ;
        RECT 268.950 210.600 271.050 210.900 ;
        RECT 254.400 209.400 271.050 210.600 ;
        RECT 229.950 208.800 232.050 209.400 ;
        RECT 268.950 208.800 271.050 209.400 ;
        RECT 274.950 210.600 277.050 210.900 ;
        RECT 284.400 210.600 285.600 212.400 ;
        RECT 274.950 209.400 285.600 210.600 ;
        RECT 301.950 210.600 304.050 211.050 ;
        RECT 311.400 210.600 312.600 215.100 ;
        RECT 301.950 209.400 312.600 210.600 ;
        RECT 335.400 210.600 336.600 215.400 ;
        RECT 343.950 214.950 346.050 217.050 ;
        RECT 364.950 214.950 367.050 217.050 ;
        RECT 344.400 210.600 345.600 214.950 ;
        RECT 365.400 211.050 366.600 214.950 ;
        RECT 349.950 210.600 352.050 210.900 ;
        RECT 335.400 209.400 339.600 210.600 ;
        RECT 344.400 209.400 352.050 210.600 ;
        RECT 274.950 208.800 277.050 209.400 ;
        RECT 301.950 208.950 304.050 209.400 ;
        RECT 178.950 206.400 189.600 207.600 ;
        RECT 199.950 207.600 202.050 208.050 ;
        RECT 205.950 207.600 208.050 208.050 ;
        RECT 199.950 206.400 208.050 207.600 ;
        RECT 178.950 205.950 181.050 206.400 ;
        RECT 199.950 205.950 202.050 206.400 ;
        RECT 205.950 205.950 208.050 206.400 ;
        RECT 286.950 207.600 289.050 208.050 ;
        RECT 298.950 207.600 301.050 208.050 ;
        RECT 286.950 206.400 301.050 207.600 ;
        RECT 338.400 207.600 339.600 209.400 ;
        RECT 349.950 208.800 352.050 209.400 ;
        RECT 364.950 208.950 367.050 211.050 ;
        RECT 374.400 210.900 375.600 217.950 ;
        RECT 649.950 217.800 652.050 218.400 ;
        RECT 376.950 215.100 379.050 217.200 ;
        RECT 382.950 216.750 385.050 217.200 ;
        RECT 388.950 216.750 391.050 217.200 ;
        RECT 382.950 215.550 391.050 216.750 ;
        RECT 382.950 215.100 385.050 215.550 ;
        RECT 388.950 215.100 391.050 215.550 ;
        RECT 377.400 211.050 378.600 215.100 ;
        RECT 400.950 214.950 403.050 217.050 ;
        RECT 445.950 215.100 448.050 217.200 ;
        RECT 463.800 216.600 465.900 217.050 ;
        RECT 455.400 215.400 465.900 216.600 ;
        RECT 373.950 208.800 376.050 210.900 ;
        RECT 377.400 209.400 382.050 211.050 ;
        RECT 378.000 208.950 382.050 209.400 ;
        RECT 397.950 210.600 400.050 210.900 ;
        RECT 401.400 210.600 402.600 214.950 ;
        RECT 397.950 209.400 402.600 210.600 ;
        RECT 430.950 210.600 433.050 210.900 ;
        RECT 446.400 210.600 447.600 215.100 ;
        RECT 455.400 210.900 456.600 215.400 ;
        RECT 463.800 214.950 465.900 215.400 ;
        RECT 466.950 215.100 469.050 217.200 ;
        RECT 467.400 211.050 468.600 215.100 ;
        RECT 484.800 214.950 486.900 217.050 ;
        RECT 487.950 215.100 490.050 217.200 ;
        RECT 514.950 216.600 517.050 217.200 ;
        RECT 526.950 216.600 529.050 217.200 ;
        RECT 514.950 215.400 529.050 216.600 ;
        RECT 514.950 215.100 517.050 215.400 ;
        RECT 526.950 215.100 529.050 215.400 ;
        RECT 553.950 215.100 556.050 217.200 ;
        RECT 625.950 216.750 628.050 217.200 ;
        RECT 634.800 216.750 636.900 217.200 ;
        RECT 625.950 215.550 636.900 216.750 ;
        RECT 625.950 215.100 628.050 215.550 ;
        RECT 634.800 215.100 636.900 215.550 ;
        RECT 430.950 209.400 447.600 210.600 ;
        RECT 397.950 208.800 400.050 209.400 ;
        RECT 430.950 208.800 433.050 209.400 ;
        RECT 454.950 208.800 457.050 210.900 ;
        RECT 463.950 209.400 468.600 211.050 ;
        RECT 463.950 208.950 468.000 209.400 ;
        RECT 485.250 208.050 486.450 214.950 ;
        RECT 488.400 213.600 489.600 215.100 ;
        RECT 554.400 213.600 555.600 215.100 ;
        RECT 559.950 213.600 562.050 214.050 ;
        RECT 637.950 213.600 640.050 217.050 ;
        RECT 652.950 216.600 655.050 217.050 ;
        RECT 661.950 216.600 664.050 217.200 ;
        RECT 676.950 216.600 679.050 217.050 ;
        RECT 652.950 215.400 679.050 216.600 ;
        RECT 652.950 214.950 655.050 215.400 ;
        RECT 661.950 215.100 664.050 215.400 ;
        RECT 662.400 213.600 663.600 215.100 ;
        RECT 676.950 214.950 679.050 215.400 ;
        RECT 488.400 212.400 492.600 213.600 ;
        RECT 554.400 212.400 558.600 213.600 ;
        RECT 491.400 210.600 492.600 212.400 ;
        RECT 496.950 210.600 499.050 211.050 ;
        RECT 491.400 209.400 499.050 210.600 ;
        RECT 496.950 208.950 499.050 209.400 ;
        RECT 502.950 210.450 505.050 210.900 ;
        RECT 511.950 210.450 514.050 210.900 ;
        RECT 502.950 209.250 514.050 210.450 ;
        RECT 557.400 210.600 558.600 212.400 ;
        RECT 559.950 213.000 640.050 213.600 ;
        RECT 659.400 213.000 663.600 213.600 ;
        RECT 559.950 212.400 639.600 213.000 ;
        RECT 658.950 212.400 663.600 213.000 ;
        RECT 559.950 211.950 562.050 212.400 ;
        RECT 568.950 210.600 571.050 210.900 ;
        RECT 557.400 209.400 571.050 210.600 ;
        RECT 502.950 208.800 505.050 209.250 ;
        RECT 511.950 208.800 514.050 209.250 ;
        RECT 568.950 208.800 571.050 209.400 ;
        RECT 580.950 210.450 583.050 210.900 ;
        RECT 589.950 210.450 592.050 210.900 ;
        RECT 580.950 209.250 592.050 210.450 ;
        RECT 580.950 208.800 583.050 209.250 ;
        RECT 589.950 208.800 592.050 209.250 ;
        RECT 622.950 210.600 625.050 210.900 ;
        RECT 640.950 210.600 643.050 210.900 ;
        RECT 622.950 209.400 643.050 210.600 ;
        RECT 622.950 208.800 625.050 209.400 ;
        RECT 640.950 208.800 643.050 209.400 ;
        RECT 658.950 208.950 661.050 212.400 ;
        RECT 664.950 210.600 667.050 210.900 ;
        RECT 680.400 210.600 681.600 218.400 ;
        RECT 691.950 218.400 709.050 219.600 ;
        RECT 691.950 217.950 694.050 218.400 ;
        RECT 706.950 217.950 709.050 218.400 ;
        RECT 808.950 219.600 811.050 220.050 ;
        RECT 808.950 218.400 864.600 219.600 ;
        RECT 808.950 217.950 811.050 218.400 ;
        RECT 685.950 215.100 688.050 217.200 ;
        RECT 686.400 211.050 687.600 215.100 ;
        RECT 694.950 214.950 697.050 217.050 ;
        RECT 709.950 214.950 712.050 217.050 ;
        RECT 733.950 216.750 736.050 217.200 ;
        RECT 742.950 216.750 745.050 217.200 ;
        RECT 733.950 215.550 745.050 216.750 ;
        RECT 733.950 215.100 736.050 215.550 ;
        RECT 742.950 215.100 745.050 215.550 ;
        RECT 778.950 216.600 781.050 217.200 ;
        RECT 793.950 216.600 796.050 217.200 ;
        RECT 778.950 215.400 796.050 216.600 ;
        RECT 778.950 215.100 781.050 215.400 ;
        RECT 793.950 215.100 796.050 215.400 ;
        RECT 814.950 216.600 817.050 217.200 ;
        RECT 835.950 216.600 838.050 217.200 ;
        RECT 814.950 215.400 838.050 216.600 ;
        RECT 814.950 215.100 817.050 215.400 ;
        RECT 835.950 215.100 838.050 215.400 ;
        RECT 847.950 215.100 850.050 217.200 ;
        RECT 863.400 216.600 864.600 218.400 ;
        RECT 865.950 216.600 868.050 217.200 ;
        RECT 863.400 215.400 868.050 216.600 ;
        RECT 865.950 215.100 868.050 215.400 ;
        RECT 695.400 211.050 696.600 214.950 ;
        RECT 710.400 211.050 711.600 214.950 ;
        RECT 664.950 209.400 684.600 210.600 ;
        RECT 686.400 209.400 691.050 211.050 ;
        RECT 664.950 208.800 667.050 209.400 ;
        RECT 338.400 206.400 384.600 207.600 ;
        RECT 485.250 206.400 490.050 208.050 ;
        RECT 286.950 205.950 289.050 206.400 ;
        RECT 298.950 205.950 301.050 206.400 ;
        RECT 383.400 205.050 384.600 206.400 ;
        RECT 486.000 205.950 490.050 206.400 ;
        RECT 592.950 207.600 595.050 208.050 ;
        RECT 601.950 207.600 604.050 208.050 ;
        RECT 616.950 207.600 619.050 208.050 ;
        RECT 592.950 206.400 619.050 207.600 ;
        RECT 592.950 205.950 595.050 206.400 ;
        RECT 601.950 205.950 604.050 206.400 ;
        RECT 616.950 205.950 619.050 206.400 ;
        RECT 622.950 207.600 625.050 207.750 ;
        RECT 631.950 207.600 634.050 208.050 ;
        RECT 622.950 206.400 634.050 207.600 ;
        RECT 683.400 207.600 684.600 209.400 ;
        RECT 687.000 208.950 691.050 209.400 ;
        RECT 694.950 208.950 697.050 211.050 ;
        RECT 709.950 208.950 712.050 211.050 ;
        RECT 718.950 210.600 721.050 210.900 ;
        RECT 748.950 210.600 751.050 210.900 ;
        RECT 718.950 209.400 751.050 210.600 ;
        RECT 718.950 208.800 721.050 209.400 ;
        RECT 748.950 208.800 751.050 209.400 ;
        RECT 805.950 210.450 808.050 210.900 ;
        RECT 817.950 210.600 820.050 210.900 ;
        RECT 838.950 210.600 841.050 210.900 ;
        RECT 817.950 210.450 841.050 210.600 ;
        RECT 805.950 209.400 841.050 210.450 ;
        RECT 805.950 209.250 820.050 209.400 ;
        RECT 805.950 208.800 808.050 209.250 ;
        RECT 817.950 208.800 820.050 209.250 ;
        RECT 838.950 208.800 841.050 209.400 ;
        RECT 719.400 207.600 720.600 208.800 ;
        RECT 848.400 208.050 849.600 215.100 ;
        RECT 871.950 214.950 874.050 217.050 ;
        RECT 853.950 210.450 856.050 210.900 ;
        RECT 862.950 210.450 865.050 210.900 ;
        RECT 853.950 209.250 865.050 210.450 ;
        RECT 853.950 208.800 856.050 209.250 ;
        RECT 862.950 208.800 865.050 209.250 ;
        RECT 868.950 210.600 871.050 210.900 ;
        RECT 872.400 210.600 873.600 214.950 ;
        RECT 868.950 209.400 873.600 210.600 ;
        RECT 868.950 208.800 871.050 209.400 ;
        RECT 683.400 206.400 720.600 207.600 ;
        RECT 622.950 205.650 625.050 206.400 ;
        RECT 631.950 205.950 634.050 206.400 ;
        RECT 847.950 205.950 850.050 208.050 ;
        RECT 4.950 204.600 7.050 205.050 ;
        RECT 13.950 204.600 16.050 205.050 ;
        RECT 4.950 203.400 16.050 204.600 ;
        RECT 4.950 202.950 7.050 203.400 ;
        RECT 13.950 202.950 16.050 203.400 ;
        RECT 103.950 204.600 106.050 205.050 ;
        RECT 139.950 204.600 142.050 205.050 ;
        RECT 103.950 203.400 142.050 204.600 ;
        RECT 103.950 202.950 106.050 203.400 ;
        RECT 139.950 202.950 142.050 203.400 ;
        RECT 160.950 204.600 163.050 205.050 ;
        RECT 187.950 204.600 190.050 205.050 ;
        RECT 160.950 203.400 190.050 204.600 ;
        RECT 160.950 202.950 163.050 203.400 ;
        RECT 187.950 202.950 190.050 203.400 ;
        RECT 271.950 204.600 274.050 205.050 ;
        RECT 280.950 204.600 283.050 205.050 ;
        RECT 271.950 203.400 283.050 204.600 ;
        RECT 271.950 202.950 274.050 203.400 ;
        RECT 280.950 202.950 283.050 203.400 ;
        RECT 382.950 204.600 385.050 205.050 ;
        RECT 412.950 204.600 415.050 205.050 ;
        RECT 382.950 203.400 415.050 204.600 ;
        RECT 382.950 202.950 385.050 203.400 ;
        RECT 412.950 202.950 415.050 203.400 ;
        RECT 469.950 204.600 472.050 205.050 ;
        RECT 481.950 204.600 484.050 205.050 ;
        RECT 469.950 203.400 484.050 204.600 ;
        RECT 469.950 202.950 472.050 203.400 ;
        RECT 481.950 202.950 484.050 203.400 ;
        RECT 511.950 204.600 514.050 205.050 ;
        RECT 541.950 204.600 544.050 205.050 ;
        RECT 511.950 203.400 544.050 204.600 ;
        RECT 511.950 202.950 514.050 203.400 ;
        RECT 541.950 202.950 544.050 203.400 ;
        RECT 640.950 204.600 643.050 205.050 ;
        RECT 655.950 204.600 658.050 205.050 ;
        RECT 640.950 203.400 658.050 204.600 ;
        RECT 640.950 202.950 643.050 203.400 ;
        RECT 655.950 202.950 658.050 203.400 ;
        RECT 688.950 204.600 691.050 205.050 ;
        RECT 754.950 204.600 757.050 205.050 ;
        RECT 760.950 204.600 763.050 205.050 ;
        RECT 688.950 203.400 717.600 204.600 ;
        RECT 688.950 202.950 691.050 203.400 ;
        RECT 22.950 201.600 25.050 202.050 ;
        RECT 34.950 201.600 37.050 202.050 ;
        RECT 22.950 200.400 37.050 201.600 ;
        RECT 22.950 199.950 25.050 200.400 ;
        RECT 34.950 199.950 37.050 200.400 ;
        RECT 190.950 201.600 193.050 202.050 ;
        RECT 196.950 201.600 199.050 202.050 ;
        RECT 214.950 201.600 217.050 202.050 ;
        RECT 283.950 201.600 286.050 202.050 ;
        RECT 190.950 200.400 286.050 201.600 ;
        RECT 190.950 199.950 193.050 200.400 ;
        RECT 196.950 199.950 199.050 200.400 ;
        RECT 214.950 199.950 217.050 200.400 ;
        RECT 283.950 199.950 286.050 200.400 ;
        RECT 319.950 201.600 322.050 202.050 ;
        RECT 334.950 201.600 337.050 202.050 ;
        RECT 319.950 200.400 337.050 201.600 ;
        RECT 319.950 199.950 322.050 200.400 ;
        RECT 334.950 199.950 337.050 200.400 ;
        RECT 379.950 201.600 382.050 202.050 ;
        RECT 391.950 201.600 394.050 202.050 ;
        RECT 379.950 200.400 394.050 201.600 ;
        RECT 379.950 199.950 382.050 200.400 ;
        RECT 391.950 199.950 394.050 200.400 ;
        RECT 451.950 201.600 454.050 202.050 ;
        RECT 460.950 201.600 463.050 202.050 ;
        RECT 451.950 200.400 463.050 201.600 ;
        RECT 451.950 199.950 454.050 200.400 ;
        RECT 460.950 199.950 463.050 200.400 ;
        RECT 499.950 201.600 502.050 202.050 ;
        RECT 526.950 201.600 529.050 202.050 ;
        RECT 616.950 201.600 619.050 202.050 ;
        RECT 499.950 200.400 529.050 201.600 ;
        RECT 499.950 199.950 502.050 200.400 ;
        RECT 526.950 199.950 529.050 200.400 ;
        RECT 569.400 200.400 619.050 201.600 ;
        RECT 569.400 199.050 570.600 200.400 ;
        RECT 616.950 199.950 619.050 200.400 ;
        RECT 637.950 201.600 640.050 202.050 ;
        RECT 667.950 201.600 670.050 202.050 ;
        RECT 637.950 200.400 670.050 201.600 ;
        RECT 637.950 199.950 640.050 200.400 ;
        RECT 667.950 199.950 670.050 200.400 ;
        RECT 682.950 201.600 685.050 202.050 ;
        RECT 697.950 201.600 700.050 202.050 ;
        RECT 682.950 200.400 700.050 201.600 ;
        RECT 716.400 201.600 717.600 203.400 ;
        RECT 754.950 203.400 763.050 204.600 ;
        RECT 754.950 202.950 757.050 203.400 ;
        RECT 760.950 202.950 763.050 203.400 ;
        RECT 787.950 204.600 790.050 205.050 ;
        RECT 805.950 204.600 808.050 205.050 ;
        RECT 787.950 203.400 808.050 204.600 ;
        RECT 787.950 202.950 790.050 203.400 ;
        RECT 805.950 202.950 808.050 203.400 ;
        RECT 814.950 204.600 817.050 205.050 ;
        RECT 826.950 204.600 829.050 205.050 ;
        RECT 814.950 203.400 829.050 204.600 ;
        RECT 814.950 202.950 817.050 203.400 ;
        RECT 826.950 202.950 829.050 203.400 ;
        RECT 721.800 201.600 723.900 202.050 ;
        RECT 716.400 200.400 723.900 201.600 ;
        RECT 682.950 199.950 685.050 200.400 ;
        RECT 697.950 199.950 700.050 200.400 ;
        RECT 721.800 199.950 723.900 200.400 ;
        RECT 724.950 201.600 727.050 202.050 ;
        RECT 766.950 201.600 769.050 202.050 ;
        RECT 724.950 200.400 769.050 201.600 ;
        RECT 724.950 199.950 727.050 200.400 ;
        RECT 766.950 199.950 769.050 200.400 ;
        RECT 790.950 201.600 793.050 202.050 ;
        RECT 796.950 201.600 799.050 202.050 ;
        RECT 790.950 200.400 799.050 201.600 ;
        RECT 790.950 199.950 793.050 200.400 ;
        RECT 796.950 199.950 799.050 200.400 ;
        RECT 97.950 198.600 100.050 199.050 ;
        RECT 127.950 198.600 130.050 199.050 ;
        RECT 97.950 197.400 130.050 198.600 ;
        RECT 97.950 196.950 100.050 197.400 ;
        RECT 127.950 196.950 130.050 197.400 ;
        RECT 139.950 198.600 142.050 199.050 ;
        RECT 229.950 198.600 232.050 199.050 ;
        RECT 139.950 197.400 232.050 198.600 ;
        RECT 139.950 196.950 142.050 197.400 ;
        RECT 229.950 196.950 232.050 197.400 ;
        RECT 250.950 198.600 253.050 199.050 ;
        RECT 307.950 198.600 310.050 199.050 ;
        RECT 250.950 197.400 310.050 198.600 ;
        RECT 250.950 196.950 253.050 197.400 ;
        RECT 307.950 196.950 310.050 197.400 ;
        RECT 313.950 198.600 316.050 199.050 ;
        RECT 334.950 198.600 337.050 198.900 ;
        RECT 313.950 197.400 337.050 198.600 ;
        RECT 313.950 196.950 316.050 197.400 ;
        RECT 334.950 196.800 337.050 197.400 ;
        RECT 490.950 198.600 493.050 199.050 ;
        RECT 514.950 198.600 517.050 199.050 ;
        RECT 490.950 197.400 517.050 198.600 ;
        RECT 490.950 196.950 493.050 197.400 ;
        RECT 514.950 196.950 517.050 197.400 ;
        RECT 535.950 198.600 538.050 199.050 ;
        RECT 544.950 198.600 547.050 199.050 ;
        RECT 535.950 197.400 547.050 198.600 ;
        RECT 535.950 196.950 538.050 197.400 ;
        RECT 544.950 196.950 547.050 197.400 ;
        RECT 550.950 198.600 553.050 199.050 ;
        RECT 568.950 198.600 571.050 199.050 ;
        RECT 550.950 197.400 571.050 198.600 ;
        RECT 550.950 196.950 553.050 197.400 ;
        RECT 568.950 196.950 571.050 197.400 ;
        RECT 583.950 198.600 586.050 199.050 ;
        RECT 619.950 198.600 622.050 199.050 ;
        RECT 583.950 197.400 622.050 198.600 ;
        RECT 583.950 196.950 586.050 197.400 ;
        RECT 619.950 196.950 622.050 197.400 ;
        RECT 634.950 198.600 637.050 199.050 ;
        RECT 643.950 198.600 646.050 199.050 ;
        RECT 673.950 198.600 676.050 199.050 ;
        RECT 679.950 198.600 682.050 199.050 ;
        RECT 634.950 197.400 682.050 198.600 ;
        RECT 634.950 196.950 637.050 197.400 ;
        RECT 643.950 196.950 646.050 197.400 ;
        RECT 673.950 196.950 676.050 197.400 ;
        RECT 679.950 196.950 682.050 197.400 ;
        RECT 763.950 198.600 766.050 199.050 ;
        RECT 823.950 198.600 826.050 199.050 ;
        RECT 844.950 198.600 847.050 199.050 ;
        RECT 850.950 198.600 853.050 199.050 ;
        RECT 763.950 197.400 853.050 198.600 ;
        RECT 763.950 196.950 766.050 197.400 ;
        RECT 823.950 196.950 826.050 197.400 ;
        RECT 844.950 196.950 847.050 197.400 ;
        RECT 850.950 196.950 853.050 197.400 ;
        RECT 1.950 195.600 4.050 196.050 ;
        RECT 28.950 195.600 31.050 196.050 ;
        RECT 1.950 194.400 31.050 195.600 ;
        RECT 1.950 193.950 4.050 194.400 ;
        RECT 28.950 193.950 31.050 194.400 ;
        RECT 100.950 195.600 103.050 196.050 ;
        RECT 109.950 195.600 112.050 196.050 ;
        RECT 100.950 194.400 112.050 195.600 ;
        RECT 100.950 193.950 103.050 194.400 ;
        RECT 109.950 193.950 112.050 194.400 ;
        RECT 154.950 195.600 157.050 196.050 ;
        RECT 178.950 195.600 181.050 196.050 ;
        RECT 154.950 194.400 181.050 195.600 ;
        RECT 154.950 193.950 157.050 194.400 ;
        RECT 178.950 193.950 181.050 194.400 ;
        RECT 232.950 195.600 235.050 196.050 ;
        RECT 238.950 195.600 241.050 196.050 ;
        RECT 232.950 194.400 241.050 195.600 ;
        RECT 232.950 193.950 235.050 194.400 ;
        RECT 238.950 193.950 241.050 194.400 ;
        RECT 316.950 195.600 319.050 196.050 ;
        RECT 352.950 195.600 355.050 196.050 ;
        RECT 316.950 194.400 355.050 195.600 ;
        RECT 316.950 193.950 319.050 194.400 ;
        RECT 352.950 193.950 355.050 194.400 ;
        RECT 358.950 195.600 361.050 196.050 ;
        RECT 373.950 195.600 376.050 196.050 ;
        RECT 358.950 194.400 376.050 195.600 ;
        RECT 358.950 193.950 361.050 194.400 ;
        RECT 373.950 193.950 376.050 194.400 ;
        RECT 448.950 195.600 451.050 196.050 ;
        RECT 460.950 195.600 463.050 196.050 ;
        RECT 475.950 195.600 478.050 196.050 ;
        RECT 496.950 195.600 499.050 196.050 ;
        RECT 448.950 194.400 499.050 195.600 ;
        RECT 448.950 193.950 451.050 194.400 ;
        RECT 460.950 193.950 463.050 194.400 ;
        RECT 475.950 193.950 478.050 194.400 ;
        RECT 496.950 193.950 499.050 194.400 ;
        RECT 517.950 195.600 520.050 196.050 ;
        RECT 541.950 195.600 544.050 196.050 ;
        RECT 580.950 195.600 583.050 196.050 ;
        RECT 829.950 195.600 832.050 196.050 ;
        RECT 841.950 195.600 844.050 196.050 ;
        RECT 517.950 194.400 544.050 195.600 ;
        RECT 517.950 193.950 520.050 194.400 ;
        RECT 541.950 193.950 544.050 194.400 ;
        RECT 557.400 194.400 573.600 195.600 ;
        RECT 91.950 192.600 94.050 193.050 ;
        RECT 121.950 192.600 124.050 193.050 ;
        RECT 133.950 192.600 136.050 193.050 ;
        RECT 91.950 191.400 136.050 192.600 ;
        RECT 91.950 190.950 94.050 191.400 ;
        RECT 121.950 190.950 124.050 191.400 ;
        RECT 133.950 190.950 136.050 191.400 ;
        RECT 181.950 192.600 184.050 193.050 ;
        RECT 259.950 192.600 262.050 193.050 ;
        RECT 181.950 191.400 262.050 192.600 ;
        RECT 181.950 190.950 184.050 191.400 ;
        RECT 259.950 190.950 262.050 191.400 ;
        RECT 361.950 192.600 364.050 193.050 ;
        RECT 367.950 192.600 370.050 193.050 ;
        RECT 361.950 191.400 370.050 192.600 ;
        RECT 361.950 190.950 364.050 191.400 ;
        RECT 367.950 190.950 370.050 191.400 ;
        RECT 403.950 192.600 406.050 193.050 ;
        RECT 445.950 192.600 448.050 193.050 ;
        RECT 463.950 192.600 466.050 193.050 ;
        RECT 557.400 192.600 558.600 194.400 ;
        RECT 403.950 191.400 429.600 192.600 ;
        RECT 403.950 190.950 406.050 191.400 ;
        RECT 79.950 189.600 82.050 190.050 ;
        RECT 115.950 189.600 118.050 190.050 ;
        RECT 79.950 188.400 118.050 189.600 ;
        RECT 79.950 187.950 82.050 188.400 ;
        RECT 115.950 187.950 118.050 188.400 ;
        RECT 316.950 189.600 319.050 190.050 ;
        RECT 328.950 189.600 331.050 190.050 ;
        RECT 316.950 188.400 331.050 189.600 ;
        RECT 316.950 187.950 319.050 188.400 ;
        RECT 328.950 187.950 331.050 188.400 ;
        RECT 343.950 189.600 346.050 190.050 ;
        RECT 349.950 189.600 352.050 190.050 ;
        RECT 343.950 188.400 352.050 189.600 ;
        RECT 343.950 187.950 346.050 188.400 ;
        RECT 349.950 187.950 352.050 188.400 ;
        RECT 391.950 189.600 394.050 190.050 ;
        RECT 421.950 189.600 424.050 190.050 ;
        RECT 391.950 188.400 424.050 189.600 ;
        RECT 428.400 189.600 429.600 191.400 ;
        RECT 445.950 191.400 466.050 192.600 ;
        RECT 445.950 190.950 448.050 191.400 ;
        RECT 463.950 190.950 466.050 191.400 ;
        RECT 551.400 191.400 558.600 192.600 ;
        RECT 572.400 192.600 573.600 194.400 ;
        RECT 580.950 194.400 615.600 195.600 ;
        RECT 580.950 193.950 583.050 194.400 ;
        RECT 592.800 192.600 594.900 193.050 ;
        RECT 572.400 191.400 594.900 192.600 ;
        RECT 454.950 189.600 457.050 190.050 ;
        RECT 428.400 188.400 457.050 189.600 ;
        RECT 391.950 187.950 394.050 188.400 ;
        RECT 421.950 187.950 424.050 188.400 ;
        RECT 454.950 187.950 457.050 188.400 ;
        RECT 466.950 189.600 469.050 190.050 ;
        RECT 499.950 189.600 502.050 190.050 ;
        RECT 466.950 188.400 502.050 189.600 ;
        RECT 466.950 187.950 469.050 188.400 ;
        RECT 499.950 187.950 502.050 188.400 ;
        RECT 505.950 189.600 508.050 190.050 ;
        RECT 551.400 189.600 552.600 191.400 ;
        RECT 592.800 190.950 594.900 191.400 ;
        RECT 595.950 192.600 598.050 193.050 ;
        RECT 614.400 192.600 615.600 194.400 ;
        RECT 829.950 194.400 844.050 195.600 ;
        RECT 829.950 193.950 832.050 194.400 ;
        RECT 841.950 193.950 844.050 194.400 ;
        RECT 856.950 195.600 859.050 196.050 ;
        RECT 862.950 195.600 865.050 196.050 ;
        RECT 856.950 194.400 865.050 195.600 ;
        RECT 856.950 193.950 859.050 194.400 ;
        RECT 862.950 193.950 865.050 194.400 ;
        RECT 628.950 192.600 631.050 193.050 ;
        RECT 595.950 191.400 612.600 192.600 ;
        RECT 614.400 191.400 631.050 192.600 ;
        RECT 595.950 190.950 598.050 191.400 ;
        RECT 505.950 188.400 552.600 189.600 ;
        RECT 505.950 187.950 508.050 188.400 ;
        RECT 4.950 186.600 7.050 187.050 ;
        RECT 19.950 186.600 22.050 187.050 ;
        RECT 4.950 185.400 22.050 186.600 ;
        RECT 4.950 184.950 7.050 185.400 ;
        RECT 19.950 184.950 22.050 185.400 ;
        RECT 88.950 186.600 91.050 187.050 ;
        RECT 97.950 186.600 100.050 187.050 ;
        RECT 88.950 185.400 100.050 186.600 ;
        RECT 88.950 184.950 91.050 185.400 ;
        RECT 97.950 184.950 100.050 185.400 ;
        RECT 154.950 186.600 157.050 187.050 ;
        RECT 160.950 186.600 163.050 187.050 ;
        RECT 154.950 185.400 163.050 186.600 ;
        RECT 154.950 184.950 157.050 185.400 ;
        RECT 160.950 184.950 163.050 185.400 ;
        RECT 178.950 186.600 181.050 187.050 ;
        RECT 187.950 186.600 190.050 187.050 ;
        RECT 178.950 185.400 190.050 186.600 ;
        RECT 178.950 184.950 181.050 185.400 ;
        RECT 187.950 184.950 190.050 185.400 ;
        RECT 307.950 186.600 310.050 187.050 ;
        RECT 313.950 186.600 316.050 187.050 ;
        RECT 307.950 185.400 316.050 186.600 ;
        RECT 307.950 184.950 310.050 185.400 ;
        RECT 313.950 184.950 316.050 185.400 ;
        RECT 352.950 186.600 355.050 187.050 ;
        RECT 403.950 186.600 406.050 187.050 ;
        RECT 352.950 185.400 406.050 186.600 ;
        RECT 352.950 184.950 355.050 185.400 ;
        RECT 403.950 184.950 406.050 185.400 ;
        RECT 541.950 186.600 544.050 187.050 ;
        RECT 559.950 186.600 562.050 190.050 ;
        RECT 568.950 189.600 571.050 190.050 ;
        RECT 598.950 189.600 601.050 190.050 ;
        RECT 568.950 188.400 601.050 189.600 ;
        RECT 611.400 189.600 612.600 191.400 ;
        RECT 628.950 190.950 631.050 191.400 ;
        RECT 646.950 192.600 649.050 193.050 ;
        RECT 691.950 192.600 694.050 193.050 ;
        RECT 646.950 191.400 694.050 192.600 ;
        RECT 646.950 190.950 649.050 191.400 ;
        RECT 691.950 190.950 694.050 191.400 ;
        RECT 826.950 192.600 829.050 193.050 ;
        RECT 844.950 192.600 847.050 193.050 ;
        RECT 871.950 192.600 874.050 193.050 ;
        RECT 826.950 191.400 874.050 192.600 ;
        RECT 826.950 190.950 829.050 191.400 ;
        RECT 844.950 190.950 847.050 191.400 ;
        RECT 871.950 190.950 874.050 191.400 ;
        RECT 619.950 189.600 622.050 190.050 ;
        RECT 687.000 189.600 691.050 190.050 ;
        RECT 611.400 188.400 622.050 189.600 ;
        RECT 568.950 187.950 571.050 188.400 ;
        RECT 598.950 187.950 601.050 188.400 ;
        RECT 619.950 187.950 622.050 188.400 ;
        RECT 686.400 187.950 691.050 189.600 ;
        RECT 694.950 189.600 697.050 190.050 ;
        RECT 700.950 189.600 703.050 190.050 ;
        RECT 694.950 188.400 703.050 189.600 ;
        RECT 694.950 187.950 697.050 188.400 ;
        RECT 700.950 187.950 703.050 188.400 ;
        RECT 727.950 189.600 730.050 190.050 ;
        RECT 742.950 189.600 745.050 190.050 ;
        RECT 751.950 189.600 754.050 190.050 ;
        RECT 727.950 188.400 754.050 189.600 ;
        RECT 727.950 187.950 730.050 188.400 ;
        RECT 742.950 187.950 745.050 188.400 ;
        RECT 751.950 187.950 754.050 188.400 ;
        RECT 769.950 189.600 772.050 190.050 ;
        RECT 799.950 189.600 802.050 190.050 ;
        RECT 832.950 189.600 835.050 190.050 ;
        RECT 859.950 189.600 862.050 190.050 ;
        RECT 769.950 188.400 802.050 189.600 ;
        RECT 769.950 187.950 772.050 188.400 ;
        RECT 799.950 187.950 802.050 188.400 ;
        RECT 824.400 188.400 835.050 189.600 ;
        RECT 541.950 186.000 562.050 186.600 ;
        RECT 616.950 186.600 619.050 187.050 ;
        RECT 673.950 186.600 676.050 187.050 ;
        RECT 686.400 186.600 687.600 187.950 ;
        RECT 824.400 187.050 825.600 188.400 ;
        RECT 832.950 187.950 835.050 188.400 ;
        RECT 851.400 188.400 862.050 189.600 ;
        RECT 541.950 185.400 561.600 186.000 ;
        RECT 616.950 185.400 687.600 186.600 ;
        RECT 541.950 184.950 544.050 185.400 ;
        RECT 616.950 184.950 619.050 185.400 ;
        RECT 673.950 184.950 676.050 185.400 ;
        RECT 25.950 183.600 28.050 184.050 ;
        RECT 40.950 183.600 43.050 184.200 ;
        RECT 55.950 183.600 58.050 184.200 ;
        RECT 25.950 182.400 39.600 183.600 ;
        RECT 25.950 181.950 28.050 182.400 ;
        RECT 38.400 180.600 39.600 182.400 ;
        RECT 40.950 182.400 58.050 183.600 ;
        RECT 40.950 182.100 43.050 182.400 ;
        RECT 55.950 182.100 58.050 182.400 ;
        RECT 61.950 183.750 64.050 184.200 ;
        RECT 67.950 183.750 70.050 184.200 ;
        RECT 61.950 182.550 70.050 183.750 ;
        RECT 61.950 182.100 64.050 182.550 ;
        RECT 67.950 182.100 70.050 182.550 ;
        RECT 73.950 183.750 76.050 184.200 ;
        RECT 79.950 183.750 82.050 184.200 ;
        RECT 73.950 182.550 82.050 183.750 ;
        RECT 73.950 182.100 76.050 182.550 ;
        RECT 79.950 182.100 82.050 182.550 ;
        RECT 91.950 181.950 94.050 184.050 ;
        RECT 109.950 183.600 112.050 184.050 ;
        RECT 115.950 183.600 118.050 184.200 ;
        RECT 109.950 182.400 118.050 183.600 ;
        RECT 109.950 181.950 112.050 182.400 ;
        RECT 115.950 182.100 118.050 182.400 ;
        RECT 127.950 181.950 130.050 184.050 ;
        RECT 172.950 183.600 175.050 184.200 ;
        RECT 190.950 183.600 193.050 184.200 ;
        RECT 202.950 183.600 205.050 184.050 ;
        RECT 172.950 182.400 193.050 183.600 ;
        RECT 172.950 182.100 175.050 182.400 ;
        RECT 190.950 182.100 193.050 182.400 ;
        RECT 197.400 182.400 205.050 183.600 ;
        RECT 38.400 179.400 45.600 180.600 ;
        RECT 44.400 177.900 45.600 179.400 ;
        RECT 4.950 177.450 7.050 177.900 ;
        RECT 10.950 177.450 13.050 177.900 ;
        RECT 4.950 176.250 13.050 177.450 ;
        RECT 4.950 175.800 7.050 176.250 ;
        RECT 10.950 175.800 13.050 176.250 ;
        RECT 16.950 177.600 19.050 177.900 ;
        RECT 25.950 177.600 28.050 177.900 ;
        RECT 16.950 177.450 28.050 177.600 ;
        RECT 31.950 177.450 34.050 177.900 ;
        RECT 16.950 176.400 34.050 177.450 ;
        RECT 16.950 175.800 19.050 176.400 ;
        RECT 25.950 176.250 34.050 176.400 ;
        RECT 25.950 175.800 28.050 176.250 ;
        RECT 31.950 175.800 34.050 176.250 ;
        RECT 43.950 175.800 46.050 177.900 ;
        RECT 82.950 177.600 85.050 177.900 ;
        RECT 92.400 177.600 93.600 181.950 ;
        RECT 82.950 176.400 93.600 177.600 ;
        RECT 124.950 177.600 127.050 177.900 ;
        RECT 128.400 177.600 129.600 181.950 ;
        RECT 136.950 177.600 139.050 177.900 ;
        RECT 124.950 176.400 139.050 177.600 ;
        RECT 82.950 175.800 85.050 176.400 ;
        RECT 124.950 175.800 127.050 176.400 ;
        RECT 136.950 175.800 139.050 176.400 ;
        RECT 166.950 177.600 169.050 177.900 ;
        RECT 187.950 177.600 190.050 177.900 ;
        RECT 166.950 176.400 190.050 177.600 ;
        RECT 197.400 177.600 198.600 182.400 ;
        RECT 202.950 181.950 205.050 182.400 ;
        RECT 208.950 183.600 211.050 184.050 ;
        RECT 220.950 183.600 223.050 184.200 ;
        RECT 208.950 182.400 223.050 183.600 ;
        RECT 208.950 181.950 211.050 182.400 ;
        RECT 220.950 182.100 223.050 182.400 ;
        RECT 232.950 180.600 235.050 184.050 ;
        RECT 238.950 183.750 241.050 184.200 ;
        RECT 247.950 183.750 250.050 184.200 ;
        RECT 238.950 182.550 250.050 183.750 ;
        RECT 238.950 182.100 241.050 182.550 ;
        RECT 247.950 182.100 250.050 182.550 ;
        RECT 319.950 183.750 322.050 184.200 ;
        RECT 328.950 183.750 331.050 184.200 ;
        RECT 319.950 182.550 331.050 183.750 ;
        RECT 319.950 182.100 322.050 182.550 ;
        RECT 328.950 182.100 331.050 182.550 ;
        RECT 334.950 181.950 337.050 184.050 ;
        RECT 340.950 183.750 343.050 184.200 ;
        RECT 349.950 183.750 352.050 184.200 ;
        RECT 340.950 182.550 352.050 183.750 ;
        RECT 340.950 182.100 343.050 182.550 ;
        RECT 349.950 182.100 352.050 182.550 ;
        RECT 427.950 183.750 430.050 184.200 ;
        RECT 439.950 183.750 442.050 184.200 ;
        RECT 427.950 182.550 442.050 183.750 ;
        RECT 427.950 182.100 430.050 182.550 ;
        RECT 439.950 182.100 442.050 182.550 ;
        RECT 445.950 183.600 448.050 184.050 ;
        RECT 472.950 183.600 475.050 184.050 ;
        RECT 445.950 182.400 475.050 183.600 ;
        RECT 445.950 181.950 448.050 182.400 ;
        RECT 472.950 181.950 475.050 182.400 ;
        RECT 478.950 183.600 481.050 184.200 ;
        RECT 490.950 183.600 493.050 184.050 ;
        RECT 478.950 182.400 493.050 183.600 ;
        RECT 478.950 182.100 481.050 182.400 ;
        RECT 490.950 181.950 493.050 182.400 ;
        RECT 499.950 182.100 502.050 184.200 ;
        RECT 232.950 180.000 237.600 180.600 ;
        RECT 233.400 179.400 237.600 180.000 ;
        RECT 236.400 177.900 237.600 179.400 ;
        RECT 199.950 177.600 202.050 177.900 ;
        RECT 197.400 176.400 202.050 177.600 ;
        RECT 166.950 175.800 169.050 176.400 ;
        RECT 187.950 175.800 190.050 176.400 ;
        RECT 199.950 175.800 202.050 176.400 ;
        RECT 235.950 175.800 238.050 177.900 ;
        RECT 253.950 177.450 256.050 177.900 ;
        RECT 277.950 177.450 280.050 177.900 ;
        RECT 253.950 176.250 280.050 177.450 ;
        RECT 253.950 175.800 256.050 176.250 ;
        RECT 277.950 175.800 280.050 176.250 ;
        RECT 331.950 177.600 334.050 177.900 ;
        RECT 335.400 177.600 336.600 181.950 ;
        RECT 430.950 180.600 433.050 181.050 ;
        RECT 347.400 179.400 433.050 180.600 ;
        RECT 347.400 177.900 348.600 179.400 ;
        RECT 430.950 178.950 433.050 179.400 ;
        RECT 331.950 176.400 336.600 177.600 ;
        RECT 331.950 175.800 334.050 176.400 ;
        RECT 346.950 175.800 349.050 177.900 ;
        RECT 442.950 177.450 445.050 177.900 ;
        RECT 448.950 177.450 451.050 177.900 ;
        RECT 466.950 177.600 469.050 178.050 ;
        RECT 442.950 176.250 451.050 177.450 ;
        RECT 458.400 177.000 469.050 177.600 ;
        RECT 442.950 175.800 445.050 176.250 ;
        RECT 448.950 175.800 451.050 176.250 ;
        RECT 457.950 176.400 469.050 177.000 ;
        RECT 457.950 175.050 460.050 176.400 ;
        RECT 466.950 175.950 469.050 176.400 ;
        RECT 490.950 177.450 493.050 177.900 ;
        RECT 496.950 177.450 499.050 177.900 ;
        RECT 490.950 176.250 499.050 177.450 ;
        RECT 500.400 177.600 501.600 182.100 ;
        RECT 517.800 181.950 519.900 184.050 ;
        RECT 520.950 181.950 523.050 184.050 ;
        RECT 526.950 183.600 529.050 184.200 ;
        RECT 544.950 183.600 547.050 184.200 ;
        RECT 580.950 183.600 583.050 184.050 ;
        RECT 526.950 182.400 583.050 183.600 ;
        RECT 526.950 182.100 529.050 182.400 ;
        RECT 544.950 182.100 547.050 182.400 ;
        RECT 508.950 177.600 511.050 178.050 ;
        RECT 500.400 176.400 511.050 177.600 ;
        RECT 490.950 175.800 493.050 176.250 ;
        RECT 496.950 175.800 499.050 176.250 ;
        RECT 508.950 175.950 511.050 176.400 ;
        RECT 49.950 174.600 52.050 175.050 ;
        RECT 64.950 174.600 67.050 175.050 ;
        RECT 49.950 173.400 67.050 174.600 ;
        RECT 49.950 172.950 52.050 173.400 ;
        RECT 64.950 172.950 67.050 173.400 ;
        RECT 205.950 174.600 208.050 175.050 ;
        RECT 214.950 174.600 217.050 175.050 ;
        RECT 205.950 173.400 217.050 174.600 ;
        RECT 205.950 172.950 208.050 173.400 ;
        RECT 214.950 172.950 217.050 173.400 ;
        RECT 274.950 174.600 277.050 175.050 ;
        RECT 394.950 174.600 397.050 175.050 ;
        RECT 274.950 173.400 397.050 174.600 ;
        RECT 274.950 172.950 277.050 173.400 ;
        RECT 394.950 172.950 397.050 173.400 ;
        RECT 403.950 174.600 406.050 175.050 ;
        RECT 403.950 173.400 456.600 174.600 ;
        RECT 403.950 172.950 406.050 173.400 ;
        RECT 160.950 171.600 163.050 172.050 ;
        RECT 196.950 171.600 199.050 172.050 ;
        RECT 217.950 171.600 220.050 172.050 ;
        RECT 160.950 170.400 220.050 171.600 ;
        RECT 160.950 169.950 163.050 170.400 ;
        RECT 196.950 169.950 199.050 170.400 ;
        RECT 217.950 169.950 220.050 170.400 ;
        RECT 223.950 171.600 226.050 171.900 ;
        RECT 244.950 171.600 247.050 172.050 ;
        RECT 325.950 171.600 328.050 171.900 ;
        RECT 223.950 170.400 328.050 171.600 ;
        RECT 223.950 169.800 226.050 170.400 ;
        RECT 244.950 169.950 247.050 170.400 ;
        RECT 325.950 169.800 328.050 170.400 ;
        RECT 331.950 171.600 334.050 172.050 ;
        RECT 352.950 171.600 355.050 172.050 ;
        RECT 331.950 170.400 355.050 171.600 ;
        RECT 455.400 171.600 456.600 173.400 ;
        RECT 457.800 174.000 460.050 175.050 ;
        RECT 460.950 174.600 463.050 175.050 ;
        RECT 469.950 174.600 472.050 175.050 ;
        RECT 457.800 172.950 459.900 174.000 ;
        RECT 460.950 173.400 472.050 174.600 ;
        RECT 460.950 172.950 463.050 173.400 ;
        RECT 469.950 172.950 472.050 173.400 ;
        RECT 499.950 174.600 502.050 175.050 ;
        RECT 518.250 174.600 519.450 181.950 ;
        RECT 521.400 175.050 522.600 181.950 ;
        RECT 566.400 177.900 567.600 182.400 ;
        RECT 580.950 181.950 583.050 182.400 ;
        RECT 589.950 183.600 592.050 184.200 ;
        RECT 607.950 183.600 610.050 184.050 ;
        RECT 613.950 183.600 616.050 184.200 ;
        RECT 589.950 182.400 610.050 183.600 ;
        RECT 589.950 182.100 592.050 182.400 ;
        RECT 607.950 181.950 610.050 182.400 ;
        RECT 611.400 182.400 616.050 183.600 ;
        RECT 611.400 180.600 612.600 182.400 ;
        RECT 613.950 182.100 616.050 182.400 ;
        RECT 649.950 183.600 652.050 184.200 ;
        RECT 649.950 182.400 654.600 183.600 ;
        RECT 649.950 182.100 652.050 182.400 ;
        RECT 608.400 179.400 612.600 180.600 ;
        RECT 529.950 177.600 532.050 177.900 ;
        RECT 541.950 177.600 544.050 177.900 ;
        RECT 529.950 177.450 544.050 177.600 ;
        RECT 559.950 177.450 562.050 177.900 ;
        RECT 529.950 176.400 562.050 177.450 ;
        RECT 529.950 175.800 532.050 176.400 ;
        RECT 541.950 176.250 562.050 176.400 ;
        RECT 541.950 175.800 544.050 176.250 ;
        RECT 559.950 175.800 562.050 176.250 ;
        RECT 565.950 175.800 568.050 177.900 ;
        RECT 580.950 177.450 583.050 177.900 ;
        RECT 592.950 177.450 595.050 177.900 ;
        RECT 580.950 176.250 595.050 177.450 ;
        RECT 580.950 175.800 583.050 176.250 ;
        RECT 592.950 175.800 595.050 176.250 ;
        RECT 608.400 175.050 609.600 179.400 ;
        RECT 653.400 178.050 654.600 182.400 ;
        RECT 688.950 182.100 691.050 184.200 ;
        RECT 694.950 183.600 697.050 184.200 ;
        RECT 709.950 183.600 712.050 187.050 ;
        RECT 766.950 186.600 769.050 187.050 ;
        RECT 781.950 186.600 784.050 187.050 ;
        RECT 766.950 185.400 784.050 186.600 ;
        RECT 766.950 184.950 769.050 185.400 ;
        RECT 781.950 184.950 784.050 185.400 ;
        RECT 820.950 185.400 825.600 187.050 ;
        RECT 841.950 186.600 844.050 187.050 ;
        RECT 847.950 186.600 850.050 187.050 ;
        RECT 841.950 185.400 850.050 186.600 ;
        RECT 820.950 184.950 825.000 185.400 ;
        RECT 841.950 184.950 844.050 185.400 ;
        RECT 847.950 184.950 850.050 185.400 ;
        RECT 712.800 183.600 714.900 184.050 ;
        RECT 694.950 182.400 708.600 183.600 ;
        RECT 709.950 183.000 714.900 183.600 ;
        RECT 710.400 182.400 714.900 183.000 ;
        RECT 694.950 182.100 697.050 182.400 ;
        RECT 689.400 178.050 690.600 182.100 ;
        RECT 707.400 178.050 708.600 182.400 ;
        RECT 712.800 181.950 714.900 182.400 ;
        RECT 715.950 181.950 718.050 184.050 ;
        RECT 625.950 177.600 628.050 177.900 ;
        RECT 646.950 177.600 649.050 177.900 ;
        RECT 625.950 176.400 649.050 177.600 ;
        RECT 653.400 176.400 658.050 178.050 ;
        RECT 625.950 175.800 628.050 176.400 ;
        RECT 646.950 175.800 649.050 176.400 ;
        RECT 654.000 175.950 658.050 176.400 ;
        RECT 664.950 177.450 667.050 177.900 ;
        RECT 682.800 177.450 684.900 177.900 ;
        RECT 664.950 176.250 684.900 177.450 ;
        RECT 664.950 175.800 667.050 176.250 ;
        RECT 682.800 175.800 684.900 176.250 ;
        RECT 685.950 176.400 690.600 178.050 ;
        RECT 685.950 175.950 690.000 176.400 ;
        RECT 706.950 175.950 709.050 178.050 ;
        RECT 716.400 177.600 717.600 181.950 ;
        RECT 721.950 180.600 724.050 184.050 ;
        RECT 739.950 183.600 742.050 184.050 ;
        RECT 745.950 183.600 748.050 184.200 ;
        RECT 739.950 182.400 748.050 183.600 ;
        RECT 739.950 181.950 742.050 182.400 ;
        RECT 745.950 182.100 748.050 182.400 ;
        RECT 763.950 182.100 766.050 184.200 ;
        RECT 782.400 183.600 783.600 184.950 ;
        RECT 773.400 182.400 783.600 183.600 ;
        RECT 721.950 180.000 732.600 180.600 ;
        RECT 722.400 179.400 732.600 180.000 ;
        RECT 721.950 177.600 724.050 178.050 ;
        RECT 731.400 177.900 732.600 179.400 ;
        RECT 716.400 176.400 724.050 177.600 ;
        RECT 721.950 175.950 724.050 176.400 ;
        RECT 730.950 175.800 733.050 177.900 ;
        RECT 748.950 177.600 751.050 177.900 ;
        RECT 764.400 177.600 765.600 182.100 ;
        RECT 773.400 177.900 774.600 182.400 ;
        RECT 790.950 182.100 793.050 184.200 ;
        RECT 799.950 183.600 804.000 184.050 ;
        RECT 748.950 176.400 765.600 177.600 ;
        RECT 748.950 175.800 751.050 176.400 ;
        RECT 772.950 175.800 775.050 177.900 ;
        RECT 781.950 177.600 784.050 178.050 ;
        RECT 791.400 177.600 792.600 182.100 ;
        RECT 799.950 181.950 804.600 183.600 ;
        RECT 811.950 182.100 814.050 184.200 ;
        RECT 803.400 177.900 804.600 181.950 ;
        RECT 812.400 178.050 813.600 182.100 ;
        RECT 851.400 181.050 852.600 188.400 ;
        RECT 859.950 187.950 862.050 188.400 ;
        RECT 862.950 186.600 865.050 187.050 ;
        RECT 862.950 185.400 876.600 186.600 ;
        RECT 862.950 184.950 865.050 185.400 ;
        RECT 850.950 178.950 853.050 181.050 ;
        RECT 781.950 176.400 792.600 177.600 ;
        RECT 781.950 175.950 784.050 176.400 ;
        RECT 802.950 175.800 805.050 177.900 ;
        RECT 812.400 176.400 817.050 178.050 ;
        RECT 813.000 175.950 817.050 176.400 ;
        RECT 499.950 173.400 519.450 174.600 ;
        RECT 499.950 172.950 502.050 173.400 ;
        RECT 520.950 172.950 523.050 175.050 ;
        RECT 607.950 172.950 610.050 175.050 ;
        RECT 875.400 172.050 876.600 185.400 ;
        RECT 466.950 171.600 469.050 172.050 ;
        RECT 455.400 170.400 469.050 171.600 ;
        RECT 331.950 169.950 334.050 170.400 ;
        RECT 352.950 169.950 355.050 170.400 ;
        RECT 466.950 169.950 469.050 170.400 ;
        RECT 490.950 171.600 493.050 172.050 ;
        RECT 523.950 171.600 526.050 172.050 ;
        RECT 490.950 170.400 526.050 171.600 ;
        RECT 490.950 169.950 493.050 170.400 ;
        RECT 523.950 169.950 526.050 170.400 ;
        RECT 541.950 171.600 544.050 172.050 ;
        RECT 574.950 171.600 577.050 172.050 ;
        RECT 541.950 170.400 577.050 171.600 ;
        RECT 541.950 169.950 544.050 170.400 ;
        RECT 574.950 169.950 577.050 170.400 ;
        RECT 655.950 171.600 658.050 172.050 ;
        RECT 697.950 171.600 700.050 172.050 ;
        RECT 655.950 170.400 700.050 171.600 ;
        RECT 655.950 169.950 658.050 170.400 ;
        RECT 697.950 169.950 700.050 170.400 ;
        RECT 706.950 171.600 709.050 172.050 ;
        RECT 781.950 171.600 784.050 172.050 ;
        RECT 706.950 170.400 784.050 171.600 ;
        RECT 706.950 169.950 709.050 170.400 ;
        RECT 781.950 169.950 784.050 170.400 ;
        RECT 787.950 171.600 790.050 172.050 ;
        RECT 814.950 171.600 817.050 172.050 ;
        RECT 787.950 170.400 817.050 171.600 ;
        RECT 787.950 169.950 790.050 170.400 ;
        RECT 814.950 169.950 817.050 170.400 ;
        RECT 874.950 169.950 877.050 172.050 ;
        RECT 37.950 168.600 40.050 169.050 ;
        RECT 67.950 168.600 70.050 169.050 ;
        RECT 37.950 167.400 70.050 168.600 ;
        RECT 37.950 166.950 40.050 167.400 ;
        RECT 67.950 166.950 70.050 167.400 ;
        RECT 73.950 168.600 76.050 169.050 ;
        RECT 100.950 168.600 103.050 169.050 ;
        RECT 193.950 168.600 196.050 169.050 ;
        RECT 73.950 167.400 196.050 168.600 ;
        RECT 73.950 166.950 76.050 167.400 ;
        RECT 100.950 166.950 103.050 167.400 ;
        RECT 193.950 166.950 196.050 167.400 ;
        RECT 235.950 168.600 238.050 169.050 ;
        RECT 247.950 168.600 250.050 169.050 ;
        RECT 235.950 167.400 250.050 168.600 ;
        RECT 235.950 166.950 238.050 167.400 ;
        RECT 247.950 166.950 250.050 167.400 ;
        RECT 283.950 168.600 286.050 169.050 ;
        RECT 319.950 168.600 322.050 169.050 ;
        RECT 283.950 167.400 322.050 168.600 ;
        RECT 283.950 166.950 286.050 167.400 ;
        RECT 319.950 166.950 322.050 167.400 ;
        RECT 328.950 168.600 331.050 169.050 ;
        RECT 334.950 168.600 337.050 169.050 ;
        RECT 328.950 167.400 337.050 168.600 ;
        RECT 328.950 166.950 331.050 167.400 ;
        RECT 334.950 166.950 337.050 167.400 ;
        RECT 352.950 168.600 355.050 168.900 ;
        RECT 388.950 168.600 391.050 169.050 ;
        RECT 433.950 168.600 436.050 169.050 ;
        RECT 352.950 167.400 391.050 168.600 ;
        RECT 352.950 166.800 355.050 167.400 ;
        RECT 388.950 166.950 391.050 167.400 ;
        RECT 416.400 167.400 436.050 168.600 ;
        RECT 94.950 165.600 97.050 166.050 ;
        RECT 178.950 165.600 181.050 166.050 ;
        RECT 94.950 164.400 181.050 165.600 ;
        RECT 94.950 163.950 97.050 164.400 ;
        RECT 178.950 163.950 181.050 164.400 ;
        RECT 211.950 165.600 214.050 166.050 ;
        RECT 223.950 165.600 226.050 166.050 ;
        RECT 211.950 164.400 226.050 165.600 ;
        RECT 211.950 163.950 214.050 164.400 ;
        RECT 223.950 163.950 226.050 164.400 ;
        RECT 346.950 165.600 349.050 166.050 ;
        RECT 416.400 165.600 417.600 167.400 ;
        RECT 433.950 166.950 436.050 167.400 ;
        RECT 442.950 168.600 445.050 169.050 ;
        RECT 592.950 168.600 595.050 169.050 ;
        RECT 652.950 168.600 655.050 169.050 ;
        RECT 442.950 167.400 489.600 168.600 ;
        RECT 442.950 166.950 445.050 167.400 ;
        RECT 346.950 164.400 417.600 165.600 ;
        RECT 436.950 165.600 439.050 166.050 ;
        RECT 451.950 165.600 454.050 166.050 ;
        RECT 436.950 164.400 454.050 165.600 ;
        RECT 488.400 165.600 489.600 167.400 ;
        RECT 592.950 167.400 655.050 168.600 ;
        RECT 592.950 166.950 595.050 167.400 ;
        RECT 652.950 166.950 655.050 167.400 ;
        RECT 658.950 168.600 661.050 169.050 ;
        RECT 676.950 168.600 679.050 169.050 ;
        RECT 658.950 167.400 679.050 168.600 ;
        RECT 658.950 166.950 661.050 167.400 ;
        RECT 676.950 166.950 679.050 167.400 ;
        RECT 682.950 168.600 685.050 169.050 ;
        RECT 724.950 168.600 727.050 169.050 ;
        RECT 682.950 167.400 727.050 168.600 ;
        RECT 682.950 166.950 685.050 167.400 ;
        RECT 724.950 166.950 727.050 167.400 ;
        RECT 817.950 168.600 820.050 169.050 ;
        RECT 868.950 168.600 871.050 169.050 ;
        RECT 817.950 167.400 871.050 168.600 ;
        RECT 817.950 166.950 820.050 167.400 ;
        RECT 868.950 166.950 871.050 167.400 ;
        RECT 568.950 165.600 571.050 166.050 ;
        RECT 577.950 165.600 580.050 166.050 ;
        RECT 643.950 165.600 646.050 166.050 ;
        RECT 488.400 164.400 504.600 165.600 ;
        RECT 346.950 163.950 349.050 164.400 ;
        RECT 436.950 163.950 439.050 164.400 ;
        RECT 451.950 163.950 454.050 164.400 ;
        RECT 503.400 163.050 504.600 164.400 ;
        RECT 568.950 164.400 580.050 165.600 ;
        RECT 568.950 163.950 571.050 164.400 ;
        RECT 577.950 163.950 580.050 164.400 ;
        RECT 581.400 164.400 646.050 165.600 ;
        RECT 301.950 162.600 304.050 163.050 ;
        RECT 310.950 162.600 313.050 163.050 ;
        RECT 301.950 161.400 313.050 162.600 ;
        RECT 301.950 160.950 304.050 161.400 ;
        RECT 310.950 160.950 313.050 161.400 ;
        RECT 349.950 162.600 352.050 163.050 ;
        RECT 424.950 162.600 427.050 163.050 ;
        RECT 349.950 161.400 427.050 162.600 ;
        RECT 349.950 160.950 352.050 161.400 ;
        RECT 424.950 160.950 427.050 161.400 ;
        RECT 430.950 162.600 433.050 163.050 ;
        RECT 439.950 162.600 442.050 163.050 ;
        RECT 430.950 161.400 442.050 162.600 ;
        RECT 430.950 160.950 433.050 161.400 ;
        RECT 439.950 160.950 442.050 161.400 ;
        RECT 457.950 162.600 460.050 163.050 ;
        RECT 475.950 162.600 478.050 163.050 ;
        RECT 499.800 162.600 501.900 163.050 ;
        RECT 457.950 161.400 501.900 162.600 ;
        RECT 457.950 160.950 460.050 161.400 ;
        RECT 475.950 160.950 478.050 161.400 ;
        RECT 499.800 160.950 501.900 161.400 ;
        RECT 502.950 162.600 505.050 163.050 ;
        RECT 541.950 162.600 544.050 163.050 ;
        RECT 502.950 161.400 544.050 162.600 ;
        RECT 502.950 160.950 505.050 161.400 ;
        RECT 541.950 160.950 544.050 161.400 ;
        RECT 562.950 162.600 565.050 163.050 ;
        RECT 581.400 162.600 582.600 164.400 ;
        RECT 643.950 163.950 646.050 164.400 ;
        RECT 670.950 165.600 673.050 166.050 ;
        RECT 691.950 165.600 694.050 166.050 ;
        RECT 670.950 164.400 694.050 165.600 ;
        RECT 670.950 163.950 673.050 164.400 ;
        RECT 691.950 163.950 694.050 164.400 ;
        RECT 709.950 165.600 712.050 166.050 ;
        RECT 718.950 165.600 721.050 166.050 ;
        RECT 709.950 164.400 721.050 165.600 ;
        RECT 709.950 163.950 712.050 164.400 ;
        RECT 718.950 163.950 721.050 164.400 ;
        RECT 796.950 165.600 799.050 166.050 ;
        RECT 838.950 165.600 841.050 166.050 ;
        RECT 796.950 164.400 841.050 165.600 ;
        RECT 796.950 163.950 799.050 164.400 ;
        RECT 838.950 163.950 841.050 164.400 ;
        RECT 562.950 161.400 582.600 162.600 ;
        RECT 595.950 162.600 598.050 163.050 ;
        RECT 640.950 162.600 643.050 163.050 ;
        RECT 595.950 161.400 643.050 162.600 ;
        RECT 562.950 160.950 565.050 161.400 ;
        RECT 595.950 160.950 598.050 161.400 ;
        RECT 640.950 160.950 643.050 161.400 ;
        RECT 733.950 162.600 736.050 163.050 ;
        RECT 772.950 162.600 775.050 163.050 ;
        RECT 733.950 161.400 775.050 162.600 ;
        RECT 733.950 160.950 736.050 161.400 ;
        RECT 772.950 160.950 775.050 161.400 ;
        RECT 787.950 162.600 790.050 163.050 ;
        RECT 802.950 162.600 805.050 163.050 ;
        RECT 787.950 161.400 805.050 162.600 ;
        RECT 787.950 160.950 790.050 161.400 ;
        RECT 802.950 160.950 805.050 161.400 ;
        RECT 229.950 159.600 232.050 160.050 ;
        RECT 256.950 159.600 259.050 160.050 ;
        RECT 229.950 158.400 259.050 159.600 ;
        RECT 229.950 157.950 232.050 158.400 ;
        RECT 256.950 157.950 259.050 158.400 ;
        RECT 376.950 159.600 379.050 160.050 ;
        RECT 409.950 159.600 412.050 160.050 ;
        RECT 376.950 158.400 412.050 159.600 ;
        RECT 376.950 157.950 379.050 158.400 ;
        RECT 409.950 157.950 412.050 158.400 ;
        RECT 427.950 159.600 430.050 160.050 ;
        RECT 454.950 159.600 457.050 160.050 ;
        RECT 427.950 158.400 457.050 159.600 ;
        RECT 427.950 157.950 430.050 158.400 ;
        RECT 454.950 157.950 457.050 158.400 ;
        RECT 508.950 159.600 511.050 160.050 ;
        RECT 553.950 159.600 556.050 160.050 ;
        RECT 508.950 158.400 556.050 159.600 ;
        RECT 508.950 157.950 511.050 158.400 ;
        RECT 553.950 157.950 556.050 158.400 ;
        RECT 559.950 159.600 562.050 160.050 ;
        RECT 571.950 159.600 574.050 160.050 ;
        RECT 559.950 158.400 574.050 159.600 ;
        RECT 559.950 157.950 562.050 158.400 ;
        RECT 571.950 157.950 574.050 158.400 ;
        RECT 577.950 159.600 580.050 160.050 ;
        RECT 598.950 159.600 601.050 160.050 ;
        RECT 670.950 159.600 673.050 160.050 ;
        RECT 685.950 159.600 688.050 160.050 ;
        RECT 577.950 158.400 633.600 159.600 ;
        RECT 577.950 157.950 580.050 158.400 ;
        RECT 598.950 157.950 601.050 158.400 ;
        RECT 223.950 156.600 226.050 157.050 ;
        RECT 310.950 156.600 313.050 157.050 ;
        RECT 223.950 155.400 313.050 156.600 ;
        RECT 223.950 154.950 226.050 155.400 ;
        RECT 310.950 154.950 313.050 155.400 ;
        RECT 334.950 156.600 337.050 157.050 ;
        RECT 352.950 156.600 355.050 157.050 ;
        RECT 334.950 155.400 355.050 156.600 ;
        RECT 334.950 154.950 337.050 155.400 ;
        RECT 352.950 154.950 355.050 155.400 ;
        RECT 373.950 156.600 376.050 157.050 ;
        RECT 454.950 156.600 457.050 156.900 ;
        RECT 373.950 155.400 457.050 156.600 ;
        RECT 373.950 154.950 376.050 155.400 ;
        RECT 454.950 154.800 457.050 155.400 ;
        RECT 466.950 156.600 469.050 157.050 ;
        RECT 484.800 156.600 486.900 157.050 ;
        RECT 466.950 155.400 486.900 156.600 ;
        RECT 466.950 154.950 469.050 155.400 ;
        RECT 484.800 154.950 486.900 155.400 ;
        RECT 487.950 156.600 490.050 157.050 ;
        RECT 502.950 156.600 505.050 157.050 ;
        RECT 487.950 155.400 505.050 156.600 ;
        RECT 632.400 156.600 633.600 158.400 ;
        RECT 670.950 158.400 688.050 159.600 ;
        RECT 670.950 157.950 673.050 158.400 ;
        RECT 685.950 157.950 688.050 158.400 ;
        RECT 775.950 159.600 778.050 160.050 ;
        RECT 808.950 159.600 811.050 160.050 ;
        RECT 850.950 159.600 853.050 160.050 ;
        RECT 775.950 158.400 853.050 159.600 ;
        RECT 775.950 157.950 778.050 158.400 ;
        RECT 808.950 157.950 811.050 158.400 ;
        RECT 850.950 157.950 853.050 158.400 ;
        RECT 736.950 156.600 739.050 157.050 ;
        RECT 778.950 156.600 781.050 157.050 ;
        RECT 802.950 156.600 805.050 157.050 ;
        RECT 632.400 155.400 717.600 156.600 ;
        RECT 487.950 154.950 490.050 155.400 ;
        RECT 502.950 154.950 505.050 155.400 ;
        RECT 61.950 153.600 64.050 154.050 ;
        RECT 316.800 153.600 318.900 154.050 ;
        RECT 61.950 152.400 318.900 153.600 ;
        RECT 61.950 151.950 64.050 152.400 ;
        RECT 316.800 151.950 318.900 152.400 ;
        RECT 319.950 153.600 322.050 154.050 ;
        RECT 349.800 153.600 351.900 154.050 ;
        RECT 319.950 152.400 351.900 153.600 ;
        RECT 319.950 151.950 322.050 152.400 ;
        RECT 349.800 151.950 351.900 152.400 ;
        RECT 352.950 153.600 355.050 153.900 ;
        RECT 367.800 153.600 369.900 154.050 ;
        RECT 352.950 152.400 369.900 153.600 ;
        RECT 352.950 151.800 355.050 152.400 ;
        RECT 367.800 151.950 369.900 152.400 ;
        RECT 370.950 153.600 373.050 154.050 ;
        RECT 403.950 153.600 406.050 154.050 ;
        RECT 370.950 152.400 406.050 153.600 ;
        RECT 370.950 151.950 373.050 152.400 ;
        RECT 403.950 151.950 406.050 152.400 ;
        RECT 409.950 153.600 412.050 154.050 ;
        RECT 442.950 153.600 445.050 154.050 ;
        RECT 409.950 152.400 445.050 153.600 ;
        RECT 409.950 151.950 412.050 152.400 ;
        RECT 442.950 151.950 445.050 152.400 ;
        RECT 451.950 153.600 454.050 154.050 ;
        RECT 472.950 153.600 475.050 154.050 ;
        RECT 493.950 153.600 496.050 154.050 ;
        RECT 451.950 152.400 496.050 153.600 ;
        RECT 451.950 151.950 454.050 152.400 ;
        RECT 472.950 151.950 475.050 152.400 ;
        RECT 493.950 151.950 496.050 152.400 ;
        RECT 553.950 153.600 556.050 154.050 ;
        RECT 583.950 153.600 586.050 154.050 ;
        RECT 595.950 153.600 598.050 154.050 ;
        RECT 553.950 152.400 598.050 153.600 ;
        RECT 553.950 151.950 556.050 152.400 ;
        RECT 583.950 151.950 586.050 152.400 ;
        RECT 595.950 151.950 598.050 152.400 ;
        RECT 610.950 153.600 613.050 154.050 ;
        RECT 670.950 153.600 673.050 154.050 ;
        RECT 610.950 152.400 673.050 153.600 ;
        RECT 610.950 151.950 613.050 152.400 ;
        RECT 670.950 151.950 673.050 152.400 ;
        RECT 685.950 153.600 688.050 154.050 ;
        RECT 691.950 153.600 694.050 154.050 ;
        RECT 685.950 152.400 694.050 153.600 ;
        RECT 716.400 153.600 717.600 155.400 ;
        RECT 736.950 155.400 777.600 156.600 ;
        RECT 736.950 154.950 739.050 155.400 ;
        RECT 739.950 153.600 742.050 154.050 ;
        RECT 716.400 152.400 742.050 153.600 ;
        RECT 776.400 153.600 777.600 155.400 ;
        RECT 778.950 155.400 805.050 156.600 ;
        RECT 778.950 154.950 781.050 155.400 ;
        RECT 802.950 154.950 805.050 155.400 ;
        RECT 814.950 156.600 817.050 157.050 ;
        RECT 844.950 156.600 847.050 157.050 ;
        RECT 814.950 155.400 847.050 156.600 ;
        RECT 814.950 154.950 817.050 155.400 ;
        RECT 844.950 154.950 847.050 155.400 ;
        RECT 841.950 153.600 844.050 154.050 ;
        RECT 776.400 152.400 844.050 153.600 ;
        RECT 685.950 151.950 688.050 152.400 ;
        RECT 691.950 151.950 694.050 152.400 ;
        RECT 739.950 151.950 742.050 152.400 ;
        RECT 841.950 151.950 844.050 152.400 ;
        RECT 94.950 150.600 97.050 151.050 ;
        RECT 109.950 150.600 112.050 151.050 ;
        RECT 94.950 149.400 112.050 150.600 ;
        RECT 94.950 148.950 97.050 149.400 ;
        RECT 109.950 148.950 112.050 149.400 ;
        RECT 190.950 150.600 193.050 151.050 ;
        RECT 325.950 150.600 328.050 151.050 ;
        RECT 349.950 150.600 352.050 150.900 ;
        RECT 190.950 149.400 252.600 150.600 ;
        RECT 190.950 148.950 193.050 149.400 ;
        RECT 251.400 148.050 252.600 149.400 ;
        RECT 325.950 149.400 352.050 150.600 ;
        RECT 325.950 148.950 328.050 149.400 ;
        RECT 349.950 148.800 352.050 149.400 ;
        RECT 424.950 150.600 427.050 151.050 ;
        RECT 448.950 150.600 451.050 151.050 ;
        RECT 424.950 149.400 451.050 150.600 ;
        RECT 424.950 148.950 427.050 149.400 ;
        RECT 448.950 148.950 451.050 149.400 ;
        RECT 454.950 150.600 457.050 151.050 ;
        RECT 487.950 150.600 490.050 151.050 ;
        RECT 454.950 149.400 490.050 150.600 ;
        RECT 454.950 148.950 457.050 149.400 ;
        RECT 487.950 148.950 490.050 149.400 ;
        RECT 514.950 150.600 517.050 151.050 ;
        RECT 565.950 150.600 568.050 151.050 ;
        RECT 514.950 149.400 568.050 150.600 ;
        RECT 514.950 148.950 517.050 149.400 ;
        RECT 565.950 148.950 568.050 149.400 ;
        RECT 631.950 150.600 634.050 151.050 ;
        RECT 658.950 150.600 661.050 151.050 ;
        RECT 631.950 149.400 661.050 150.600 ;
        RECT 631.950 148.950 634.050 149.400 ;
        RECT 658.950 148.950 661.050 149.400 ;
        RECT 676.950 150.600 679.050 151.050 ;
        RECT 712.950 150.600 715.050 151.050 ;
        RECT 748.950 150.600 751.050 151.050 ;
        RECT 676.950 149.400 751.050 150.600 ;
        RECT 676.950 148.950 679.050 149.400 ;
        RECT 712.950 148.950 715.050 149.400 ;
        RECT 748.950 148.950 751.050 149.400 ;
        RECT 757.950 150.600 760.050 151.050 ;
        RECT 784.950 150.600 787.050 151.050 ;
        RECT 757.950 149.400 787.050 150.600 ;
        RECT 757.950 148.950 760.050 149.400 ;
        RECT 784.950 148.950 787.050 149.400 ;
        RECT 187.950 147.600 190.050 148.050 ;
        RECT 220.950 147.600 223.050 148.050 ;
        RECT 187.950 146.400 223.050 147.600 ;
        RECT 187.950 145.950 190.050 146.400 ;
        RECT 220.950 145.950 223.050 146.400 ;
        RECT 250.950 147.600 253.050 148.050 ;
        RECT 277.950 147.600 280.050 148.050 ;
        RECT 250.950 146.400 280.050 147.600 ;
        RECT 250.950 145.950 253.050 146.400 ;
        RECT 277.950 145.950 280.050 146.400 ;
        RECT 289.950 147.600 292.050 148.050 ;
        RECT 361.950 147.600 364.050 148.050 ;
        RECT 289.950 146.400 364.050 147.600 ;
        RECT 289.950 145.950 292.050 146.400 ;
        RECT 361.950 145.950 364.050 146.400 ;
        RECT 367.950 147.600 370.050 148.050 ;
        RECT 406.950 147.600 409.050 148.050 ;
        RECT 421.950 147.600 424.050 148.050 ;
        RECT 457.950 147.600 460.050 148.050 ;
        RECT 367.950 146.400 460.050 147.600 ;
        RECT 367.950 145.950 370.050 146.400 ;
        RECT 406.950 145.950 409.050 146.400 ;
        RECT 421.950 145.950 424.050 146.400 ;
        RECT 457.950 145.950 460.050 146.400 ;
        RECT 463.950 147.600 466.050 148.050 ;
        RECT 481.950 147.600 484.050 148.050 ;
        RECT 463.950 146.400 484.050 147.600 ;
        RECT 463.950 145.950 466.050 146.400 ;
        RECT 481.950 145.950 484.050 146.400 ;
        RECT 499.950 147.600 502.050 148.050 ;
        RECT 589.950 147.600 592.050 148.050 ;
        RECT 499.950 146.400 592.050 147.600 ;
        RECT 499.950 145.950 502.050 146.400 ;
        RECT 589.950 145.950 592.050 146.400 ;
        RECT 805.950 147.600 808.050 148.050 ;
        RECT 823.950 147.600 826.050 148.050 ;
        RECT 805.950 146.400 826.050 147.600 ;
        RECT 805.950 145.950 808.050 146.400 ;
        RECT 823.950 145.950 826.050 146.400 ;
        RECT 847.950 147.600 850.050 148.050 ;
        RECT 862.950 147.600 865.050 148.050 ;
        RECT 847.950 146.400 865.050 147.600 ;
        RECT 847.950 145.950 850.050 146.400 ;
        RECT 862.950 145.950 865.050 146.400 ;
        RECT 76.950 144.600 79.050 145.050 ;
        RECT 103.950 144.600 106.050 145.050 ;
        RECT 76.950 143.400 106.050 144.600 ;
        RECT 76.950 142.950 79.050 143.400 ;
        RECT 103.950 142.950 106.050 143.400 ;
        RECT 130.950 144.600 133.050 145.050 ;
        RECT 145.950 144.600 148.050 144.900 ;
        RECT 130.950 143.400 148.050 144.600 ;
        RECT 130.950 142.950 133.050 143.400 ;
        RECT 145.950 142.800 148.050 143.400 ;
        RECT 256.950 144.600 259.050 145.050 ;
        RECT 304.950 144.600 307.050 145.050 ;
        RECT 256.950 143.400 307.050 144.600 ;
        RECT 256.950 142.950 259.050 143.400 ;
        RECT 304.950 142.950 307.050 143.400 ;
        RECT 313.950 144.600 316.050 145.050 ;
        RECT 358.950 144.600 361.050 145.050 ;
        RECT 313.950 143.400 361.050 144.600 ;
        RECT 313.950 142.950 316.050 143.400 ;
        RECT 358.950 142.950 361.050 143.400 ;
        RECT 373.950 142.950 379.050 145.050 ;
        RECT 436.950 144.600 439.050 145.050 ;
        RECT 478.950 144.600 481.050 145.050 ;
        RECT 508.950 144.600 511.050 145.050 ;
        RECT 436.950 143.400 511.050 144.600 ;
        RECT 436.950 142.950 439.050 143.400 ;
        RECT 478.950 142.950 481.050 143.400 ;
        RECT 508.950 142.950 511.050 143.400 ;
        RECT 547.950 144.600 550.050 145.050 ;
        RECT 559.950 144.600 562.050 145.050 ;
        RECT 580.950 144.600 583.050 145.050 ;
        RECT 547.950 143.400 562.050 144.600 ;
        RECT 547.950 142.950 550.050 143.400 ;
        RECT 559.950 142.950 562.050 143.400 ;
        RECT 566.400 143.400 583.050 144.600 ;
        RECT 22.950 141.600 25.050 142.050 ;
        RECT 37.950 141.600 40.050 142.050 ;
        RECT 22.950 140.400 40.050 141.600 ;
        RECT 22.950 139.950 25.050 140.400 ;
        RECT 37.950 139.950 40.050 140.400 ;
        RECT 88.950 141.600 91.050 141.900 ;
        RECT 94.950 141.600 97.050 142.050 ;
        RECT 88.950 140.400 97.050 141.600 ;
        RECT 88.950 139.800 91.050 140.400 ;
        RECT 94.950 139.950 97.050 140.400 ;
        RECT 322.950 139.950 325.050 142.050 ;
        RECT 385.950 141.600 388.050 142.050 ;
        RECT 391.950 141.600 394.050 142.050 ;
        RECT 385.950 140.400 394.050 141.600 ;
        RECT 385.950 139.950 388.050 140.400 ;
        RECT 391.950 139.950 394.050 140.400 ;
        RECT 448.950 141.600 451.050 142.050 ;
        RECT 481.950 141.600 486.000 142.050 ;
        RECT 511.950 141.600 514.050 142.050 ;
        RECT 566.400 141.600 567.600 143.400 ;
        RECT 580.950 142.950 583.050 143.400 ;
        RECT 592.950 144.600 595.050 145.050 ;
        RECT 631.950 144.600 634.050 145.050 ;
        RECT 592.950 143.400 634.050 144.600 ;
        RECT 592.950 142.950 595.050 143.400 ;
        RECT 631.950 142.950 634.050 143.400 ;
        RECT 703.950 144.600 706.050 145.050 ;
        RECT 757.950 144.600 760.050 145.050 ;
        RECT 796.950 144.600 799.050 145.050 ;
        RECT 703.950 143.400 799.050 144.600 ;
        RECT 703.950 142.950 706.050 143.400 ;
        RECT 757.950 142.950 760.050 143.400 ;
        RECT 796.950 142.950 799.050 143.400 ;
        RECT 850.950 144.600 853.050 145.050 ;
        RECT 856.950 144.600 859.050 145.050 ;
        RECT 850.950 143.400 859.050 144.600 ;
        RECT 850.950 142.950 853.050 143.400 ;
        RECT 856.950 142.950 859.050 143.400 ;
        RECT 448.950 140.400 477.600 141.600 ;
        RECT 448.950 139.950 451.050 140.400 ;
        RECT 13.950 137.100 16.050 139.200 ;
        RECT 37.950 137.100 40.050 139.200 ;
        RECT 46.950 138.750 49.050 139.200 ;
        RECT 55.950 138.750 58.050 139.200 ;
        RECT 46.950 137.550 58.050 138.750 ;
        RECT 61.800 138.600 63.900 139.200 ;
        RECT 46.950 137.100 49.050 137.550 ;
        RECT 55.950 137.100 58.050 137.550 ;
        RECT 59.400 137.400 63.900 138.600 ;
        RECT 1.950 132.600 4.050 133.050 ;
        RECT 10.950 132.600 13.050 132.900 ;
        RECT 1.950 131.400 13.050 132.600 ;
        RECT 1.950 130.950 4.050 131.400 ;
        RECT 10.950 130.800 13.050 131.400 ;
        RECT 14.400 129.600 15.600 137.100 ;
        RECT 38.400 132.600 39.600 137.100 ;
        RECT 59.400 135.600 60.600 137.400 ;
        RECT 61.800 137.100 63.900 137.400 ;
        RECT 64.950 136.950 67.050 139.050 ;
        RECT 82.950 138.600 85.050 139.200 ;
        RECT 97.950 138.600 100.050 139.200 ;
        RECT 82.950 137.400 100.050 138.600 ;
        RECT 82.950 137.100 85.050 137.400 ;
        RECT 97.950 137.100 100.050 137.400 ;
        RECT 103.950 138.750 106.050 139.200 ;
        RECT 109.950 138.750 112.050 139.200 ;
        RECT 103.950 137.550 112.050 138.750 ;
        RECT 103.950 137.100 106.050 137.550 ;
        RECT 109.950 137.100 112.050 137.550 ;
        RECT 118.950 137.100 121.050 139.200 ;
        RECT 124.950 137.100 127.050 139.200 ;
        RECT 139.950 138.600 142.050 139.200 ;
        RECT 163.950 138.600 166.050 139.050 ;
        RECT 139.950 137.400 166.050 138.600 ;
        RECT 139.950 137.100 142.050 137.400 ;
        RECT 56.400 134.400 60.600 135.600 ;
        RECT 49.950 132.600 52.050 133.050 ;
        RECT 38.400 131.400 52.050 132.600 ;
        RECT 49.950 130.950 52.050 131.400 ;
        RECT 56.400 130.050 57.600 134.400 ;
        RECT 58.950 132.600 61.050 132.900 ;
        RECT 65.400 132.600 66.600 136.950 ;
        RECT 58.950 131.400 66.600 132.600 ;
        RECT 79.950 132.600 82.050 132.900 ;
        RECT 100.950 132.600 103.050 132.900 ;
        RECT 79.950 131.400 103.050 132.600 ;
        RECT 58.950 130.800 61.050 131.400 ;
        RECT 79.950 130.800 82.050 131.400 ;
        RECT 100.950 130.800 103.050 131.400 ;
        RECT 112.950 132.600 115.050 133.050 ;
        RECT 119.400 132.600 120.600 137.100 ;
        RECT 112.950 131.400 120.600 132.600 ;
        RECT 125.400 132.600 126.600 137.100 ;
        RECT 163.950 136.950 166.050 137.400 ;
        RECT 169.950 137.100 172.050 139.200 ;
        RECT 232.950 138.600 235.050 139.050 ;
        RECT 238.950 138.600 241.050 139.050 ;
        RECT 232.950 137.400 241.050 138.600 ;
        RECT 133.950 132.600 136.050 133.050 ;
        RECT 125.400 131.400 136.050 132.600 ;
        RECT 112.950 130.950 115.050 131.400 ;
        RECT 133.950 130.950 136.050 131.400 ;
        RECT 142.950 132.450 145.050 132.900 ;
        RECT 151.950 132.450 154.050 132.900 ;
        RECT 142.950 131.250 154.050 132.450 ;
        RECT 164.400 132.600 165.600 136.950 ;
        RECT 170.400 135.600 171.600 137.100 ;
        RECT 232.950 136.950 235.050 137.400 ;
        RECT 238.950 136.950 241.050 137.400 ;
        RECT 193.950 135.600 196.050 136.050 ;
        RECT 170.400 134.400 196.050 135.600 ;
        RECT 259.950 135.600 262.050 139.050 ;
        RECT 295.950 137.100 298.050 139.200 ;
        RECT 301.950 138.600 304.050 139.200 ;
        RECT 319.950 138.600 322.050 139.200 ;
        RECT 301.950 137.400 322.050 138.600 ;
        RECT 301.950 137.100 304.050 137.400 ;
        RECT 319.950 137.100 322.050 137.400 ;
        RECT 296.400 135.600 297.600 137.100 ;
        RECT 259.950 135.000 297.600 135.600 ;
        RECT 260.400 134.400 297.600 135.000 ;
        RECT 193.950 133.950 196.050 134.400 ;
        RECT 226.950 132.600 229.050 132.900 ;
        RECT 238.950 132.600 241.050 132.900 ;
        RECT 164.400 131.400 171.600 132.600 ;
        RECT 142.950 130.800 145.050 131.250 ;
        RECT 151.950 130.800 154.050 131.250 ;
        RECT 19.950 129.600 22.050 130.050 ;
        RECT 14.400 128.400 22.050 129.600 ;
        RECT 19.950 127.950 22.050 128.400 ;
        RECT 31.950 129.600 34.050 130.050 ;
        RECT 55.950 129.600 58.050 130.050 ;
        RECT 31.950 128.400 58.050 129.600 ;
        RECT 31.950 127.950 34.050 128.400 ;
        RECT 55.950 127.950 58.050 128.400 ;
        RECT 61.950 129.600 64.050 130.050 ;
        RECT 67.950 129.600 70.050 130.050 ;
        RECT 61.950 128.400 70.050 129.600 ;
        RECT 61.950 127.950 64.050 128.400 ;
        RECT 67.950 127.950 70.050 128.400 ;
        RECT 82.950 129.600 85.050 130.050 ;
        RECT 88.950 129.600 91.050 130.050 ;
        RECT 82.950 128.400 91.050 129.600 ;
        RECT 152.400 129.600 153.600 130.800 ;
        RECT 166.950 129.600 169.050 130.050 ;
        RECT 152.400 128.400 169.050 129.600 ;
        RECT 170.400 129.600 171.600 131.400 ;
        RECT 226.950 132.450 241.050 132.600 ;
        RECT 247.950 132.450 250.050 132.900 ;
        RECT 226.950 131.400 250.050 132.450 ;
        RECT 226.950 130.800 229.050 131.400 ;
        RECT 238.950 131.250 250.050 131.400 ;
        RECT 238.950 130.800 241.050 131.250 ;
        RECT 247.950 130.800 250.050 131.250 ;
        RECT 278.400 130.050 279.600 134.400 ;
        RECT 289.950 132.450 292.050 132.900 ;
        RECT 298.950 132.450 301.050 132.900 ;
        RECT 289.950 131.250 301.050 132.450 ;
        RECT 289.950 130.800 292.050 131.250 ;
        RECT 298.950 130.800 301.050 131.250 ;
        RECT 184.950 129.600 187.050 130.050 ;
        RECT 170.400 128.400 187.050 129.600 ;
        RECT 82.950 127.950 85.050 128.400 ;
        RECT 88.950 127.950 91.050 128.400 ;
        RECT 166.950 127.950 169.050 128.400 ;
        RECT 184.950 127.950 187.050 128.400 ;
        RECT 202.950 129.600 205.050 130.050 ;
        RECT 220.950 129.600 223.050 130.050 ;
        RECT 202.950 128.400 223.050 129.600 ;
        RECT 202.950 127.950 205.050 128.400 ;
        RECT 220.950 127.950 223.050 128.400 ;
        RECT 277.950 127.950 280.050 130.050 ;
        RECT 316.950 129.600 319.050 130.050 ;
        RECT 323.400 129.600 324.600 139.950 ;
        RECT 334.950 138.600 337.050 139.200 ;
        RECT 326.400 137.400 337.050 138.600 ;
        RECT 326.400 133.050 327.600 137.400 ;
        RECT 334.950 137.100 337.050 137.400 ;
        RECT 349.950 138.600 352.050 139.050 ;
        RECT 358.950 138.600 361.050 139.200 ;
        RECT 349.950 137.400 361.050 138.600 ;
        RECT 349.950 136.950 352.050 137.400 ;
        RECT 358.950 137.100 361.050 137.400 ;
        RECT 370.950 137.100 373.050 139.200 ;
        RECT 436.950 138.750 439.050 139.200 ;
        RECT 445.950 138.750 448.050 139.200 ;
        RECT 436.950 137.550 448.050 138.750 ;
        RECT 436.950 137.100 439.050 137.550 ;
        RECT 445.950 137.100 448.050 137.550 ;
        RECT 359.400 135.600 360.600 137.100 ;
        RECT 364.950 135.600 367.050 136.050 ;
        RECT 350.400 135.000 367.050 135.600 ;
        RECT 349.950 134.400 367.050 135.000 ;
        RECT 325.950 130.950 328.050 133.050 ;
        RECT 349.950 130.950 352.050 134.400 ;
        RECT 364.950 133.950 367.050 134.400 ;
        RECT 355.950 132.600 358.050 132.900 ;
        RECT 371.400 132.600 372.600 137.100 ;
        RECT 476.400 135.600 477.600 140.400 ;
        RECT 481.950 139.950 486.600 141.600 ;
        RECT 511.950 140.400 567.600 141.600 ;
        RECT 649.950 141.600 652.050 142.050 ;
        RECT 691.950 141.600 694.050 142.050 ;
        RECT 649.950 140.400 694.050 141.600 ;
        RECT 511.950 139.950 514.050 140.400 ;
        RECT 476.400 135.000 480.600 135.600 ;
        RECT 476.400 134.400 481.050 135.000 ;
        RECT 355.950 131.400 372.600 132.600 ;
        RECT 379.950 132.450 382.050 132.900 ;
        RECT 385.950 132.450 388.050 132.900 ;
        RECT 355.950 130.800 358.050 131.400 ;
        RECT 379.950 131.250 388.050 132.450 ;
        RECT 379.950 130.800 382.050 131.250 ;
        RECT 385.950 130.800 388.050 131.250 ;
        RECT 454.950 132.600 457.050 132.900 ;
        RECT 475.800 132.600 477.900 132.900 ;
        RECT 454.950 131.400 477.900 132.600 ;
        RECT 454.950 130.800 457.050 131.400 ;
        RECT 475.800 130.800 477.900 131.400 ;
        RECT 478.950 130.950 481.050 134.400 ;
        RECT 485.400 133.050 486.600 139.950 ;
        RECT 499.950 137.100 502.050 139.200 ;
        RECT 514.950 137.100 517.050 139.200 ;
        RECT 520.950 138.600 523.050 139.200 ;
        RECT 529.950 138.750 532.050 139.200 ;
        RECT 535.950 138.750 538.050 139.200 ;
        RECT 520.950 137.400 525.600 138.600 ;
        RECT 520.950 137.100 523.050 137.400 ;
        RECT 500.400 133.050 501.600 137.100 ;
        RECT 484.950 130.950 487.050 133.050 ;
        RECT 500.400 131.400 505.050 133.050 ;
        RECT 501.000 130.950 505.050 131.400 ;
        RECT 515.400 130.050 516.600 137.100 ;
        RECT 524.400 132.600 525.600 137.400 ;
        RECT 529.950 137.550 538.050 138.750 ;
        RECT 529.950 137.100 532.050 137.550 ;
        RECT 535.950 137.100 538.050 137.550 ;
        RECT 541.950 137.100 544.050 139.200 ;
        RECT 553.950 137.100 556.050 139.200 ;
        RECT 542.400 133.050 543.600 137.100 ;
        RECT 554.400 133.050 555.600 137.100 ;
        RECT 538.950 132.600 541.050 132.900 ;
        RECT 524.400 131.400 541.050 132.600 ;
        RECT 542.400 131.400 547.050 133.050 ;
        RECT 538.950 130.800 541.050 131.400 ;
        RECT 543.000 130.950 547.050 131.400 ;
        RECT 550.950 131.400 555.600 133.050 ;
        RECT 550.950 130.950 555.000 131.400 ;
        RECT 316.950 128.400 324.600 129.600 ;
        RECT 364.950 129.600 367.050 130.050 ;
        RECT 373.950 129.600 376.050 130.050 ;
        RECT 364.950 128.400 376.050 129.600 ;
        RECT 316.950 127.950 319.050 128.400 ;
        RECT 364.950 127.950 367.050 128.400 ;
        RECT 373.950 127.950 376.050 128.400 ;
        RECT 388.950 129.600 391.050 130.050 ;
        RECT 412.950 129.600 415.050 130.050 ;
        RECT 427.950 129.600 430.050 130.050 ;
        RECT 388.950 128.400 430.050 129.600 ;
        RECT 388.950 127.950 391.050 128.400 ;
        RECT 412.950 127.950 415.050 128.400 ;
        RECT 427.950 127.950 430.050 128.400 ;
        RECT 514.950 127.950 517.050 130.050 ;
        RECT 553.950 129.600 556.050 130.050 ;
        RECT 563.400 129.600 564.600 140.400 ;
        RECT 649.950 139.950 652.050 140.400 ;
        RECT 691.950 139.950 694.050 140.400 ;
        RECT 820.950 141.600 823.050 142.050 ;
        RECT 835.950 141.600 838.050 142.050 ;
        RECT 820.950 140.400 838.050 141.600 ;
        RECT 820.950 139.950 823.050 140.400 ;
        RECT 835.950 139.950 838.050 140.400 ;
        RECT 565.950 136.950 568.050 139.050 ;
        RECT 571.950 138.600 574.050 139.050 ;
        RECT 592.950 138.600 595.050 139.050 ;
        RECT 571.950 137.400 595.050 138.600 ;
        RECT 571.950 136.950 574.050 137.400 ;
        RECT 592.950 136.950 595.050 137.400 ;
        RECT 610.950 136.950 613.050 139.050 ;
        RECT 616.950 138.600 619.050 139.200 ;
        RECT 631.950 138.600 634.050 139.200 ;
        RECT 649.950 138.600 652.050 139.200 ;
        RECT 694.950 138.600 697.050 139.200 ;
        RECT 700.950 138.750 703.050 138.900 ;
        RECT 706.950 138.750 709.050 139.200 ;
        RECT 616.950 137.400 652.050 138.600 ;
        RECT 616.950 137.100 619.050 137.400 ;
        RECT 631.950 137.100 634.050 137.400 ;
        RECT 649.950 137.100 652.050 137.400 ;
        RECT 668.400 137.400 699.600 138.600 ;
        RECT 566.400 133.050 567.600 136.950 ;
        RECT 565.950 130.950 568.050 133.050 ;
        RECT 580.950 132.450 583.050 132.900 ;
        RECT 589.800 132.450 591.900 132.900 ;
        RECT 580.950 131.250 591.900 132.450 ;
        RECT 580.950 130.800 583.050 131.250 ;
        RECT 589.800 130.800 591.900 131.250 ;
        RECT 598.950 132.600 601.050 132.900 ;
        RECT 611.400 132.600 612.600 136.950 ;
        RECT 668.400 135.600 669.600 137.400 ;
        RECT 694.950 137.100 697.050 137.400 ;
        RECT 656.400 134.400 669.600 135.600 ;
        RECT 613.950 132.600 616.050 132.900 ;
        RECT 598.950 131.400 616.050 132.600 ;
        RECT 598.950 130.800 601.050 131.400 ;
        RECT 613.950 130.800 616.050 131.400 ;
        RECT 634.950 132.600 637.050 132.900 ;
        RECT 652.950 132.600 655.050 132.900 ;
        RECT 656.400 132.600 657.600 134.400 ;
        RECT 634.950 131.400 657.600 132.600 ;
        RECT 679.950 132.600 682.050 132.900 ;
        RECT 685.950 132.600 688.050 132.900 ;
        RECT 679.950 132.450 688.050 132.600 ;
        RECT 691.950 132.450 694.050 132.900 ;
        RECT 679.950 131.400 694.050 132.450 ;
        RECT 698.400 132.600 699.600 137.400 ;
        RECT 700.950 137.550 709.050 138.750 ;
        RECT 700.950 136.800 703.050 137.550 ;
        RECT 706.950 137.100 709.050 137.550 ;
        RECT 724.950 138.750 727.050 139.200 ;
        RECT 730.950 138.750 733.050 139.200 ;
        RECT 724.950 137.550 733.050 138.750 ;
        RECT 724.950 137.100 727.050 137.550 ;
        RECT 730.950 137.100 733.050 137.550 ;
        RECT 745.950 138.600 750.000 139.050 ;
        RECT 751.950 138.750 754.050 139.200 ;
        RECT 763.950 138.750 766.050 139.200 ;
        RECT 745.950 136.950 750.600 138.600 ;
        RECT 751.950 137.550 766.050 138.750 ;
        RECT 751.950 137.100 754.050 137.550 ;
        RECT 763.950 137.100 766.050 137.550 ;
        RECT 769.950 137.100 772.050 139.200 ;
        RECT 790.950 137.100 793.050 139.200 ;
        RECT 796.950 138.600 799.050 139.200 ;
        RECT 823.950 138.750 826.050 139.200 ;
        RECT 829.950 138.750 832.050 139.200 ;
        RECT 796.950 137.400 816.600 138.600 ;
        RECT 796.950 137.100 799.050 137.400 ;
        RECT 709.950 132.600 712.050 132.900 ;
        RECT 698.400 131.400 712.050 132.600 ;
        RECT 634.950 130.800 637.050 131.400 ;
        RECT 652.950 130.800 655.050 131.400 ;
        RECT 679.950 130.800 682.050 131.400 ;
        RECT 685.950 131.250 694.050 131.400 ;
        RECT 685.950 130.800 688.050 131.250 ;
        RECT 691.950 130.800 694.050 131.250 ;
        RECT 709.950 130.800 712.050 131.400 ;
        RECT 715.950 132.600 718.050 132.900 ;
        RECT 724.950 132.600 727.050 133.050 ;
        RECT 749.400 132.900 750.600 136.950 ;
        RECT 715.950 131.400 727.050 132.600 ;
        RECT 715.950 130.800 718.050 131.400 ;
        RECT 724.950 130.950 727.050 131.400 ;
        RECT 748.950 130.800 751.050 132.900 ;
        RECT 754.950 132.600 757.050 132.900 ;
        RECT 770.400 132.600 771.600 137.100 ;
        RECT 754.950 131.400 771.600 132.600 ;
        RECT 791.400 132.600 792.600 137.100 ;
        RECT 815.400 132.900 816.600 137.400 ;
        RECT 823.950 137.550 832.050 138.750 ;
        RECT 823.950 137.100 826.050 137.550 ;
        RECT 829.950 137.100 832.050 137.550 ;
        RECT 838.950 136.950 841.050 139.050 ;
        RECT 844.950 138.600 849.000 139.050 ;
        RECT 844.950 136.950 849.600 138.600 ;
        RECT 839.400 133.050 840.600 136.950 ;
        RECT 808.950 132.600 811.050 132.900 ;
        RECT 791.400 131.400 811.050 132.600 ;
        RECT 754.950 130.800 757.050 131.400 ;
        RECT 808.950 130.800 811.050 131.400 ;
        RECT 814.950 130.800 817.050 132.900 ;
        RECT 838.950 130.950 841.050 133.050 ;
        RECT 848.400 132.900 849.600 136.950 ;
        RECT 847.950 130.800 850.050 132.900 ;
        RECT 574.950 129.600 577.050 130.050 ;
        RECT 553.950 128.400 564.600 129.600 ;
        RECT 569.400 128.400 577.050 129.600 ;
        RECT 553.950 127.950 556.050 128.400 ;
        RECT 100.950 126.600 103.050 127.050 ;
        RECT 136.950 126.600 139.050 127.050 ;
        RECT 100.950 125.400 139.050 126.600 ;
        RECT 100.950 124.950 103.050 125.400 ;
        RECT 136.950 124.950 139.050 125.400 ;
        RECT 214.950 126.600 217.050 127.050 ;
        RECT 229.950 126.600 232.050 127.050 ;
        RECT 214.950 125.400 232.050 126.600 ;
        RECT 214.950 124.950 217.050 125.400 ;
        RECT 229.950 124.950 232.050 125.400 ;
        RECT 235.950 126.600 238.050 127.050 ;
        RECT 265.950 126.600 268.050 127.050 ;
        RECT 235.950 125.400 268.050 126.600 ;
        RECT 235.950 124.950 238.050 125.400 ;
        RECT 265.950 124.950 268.050 125.400 ;
        RECT 337.950 126.600 340.050 127.050 ;
        RECT 349.950 126.600 352.050 127.050 ;
        RECT 337.950 125.400 352.050 126.600 ;
        RECT 337.950 124.950 340.050 125.400 ;
        RECT 349.950 124.950 352.050 125.400 ;
        RECT 463.950 126.600 466.050 127.050 ;
        RECT 469.950 126.600 472.050 127.050 ;
        RECT 463.950 125.400 472.050 126.600 ;
        RECT 463.950 124.950 466.050 125.400 ;
        RECT 469.950 124.950 472.050 125.400 ;
        RECT 475.950 126.600 478.050 127.050 ;
        RECT 511.950 126.600 514.050 127.050 ;
        RECT 475.950 125.400 514.050 126.600 ;
        RECT 475.950 124.950 478.050 125.400 ;
        RECT 511.950 124.950 514.050 125.400 ;
        RECT 526.950 126.600 529.050 127.050 ;
        RECT 538.950 126.600 541.050 127.050 ;
        RECT 526.950 125.400 541.050 126.600 ;
        RECT 526.950 124.950 529.050 125.400 ;
        RECT 538.950 124.950 541.050 125.400 ;
        RECT 547.950 126.600 550.050 127.050 ;
        RECT 569.400 126.600 570.600 128.400 ;
        RECT 574.950 127.950 577.050 128.400 ;
        RECT 664.950 129.600 667.050 130.050 ;
        RECT 673.950 129.600 676.050 130.050 ;
        RECT 664.950 128.400 676.050 129.600 ;
        RECT 664.950 127.950 667.050 128.400 ;
        RECT 673.950 127.950 676.050 128.400 ;
        RECT 733.950 129.600 736.050 130.050 ;
        RECT 745.950 129.600 748.050 130.050 ;
        RECT 733.950 128.400 748.050 129.600 ;
        RECT 733.950 127.950 736.050 128.400 ;
        RECT 745.950 127.950 748.050 128.400 ;
        RECT 751.950 129.600 754.050 130.050 ;
        RECT 772.950 129.600 775.050 130.050 ;
        RECT 751.950 128.400 775.050 129.600 ;
        RECT 751.950 127.950 754.050 128.400 ;
        RECT 772.950 127.950 775.050 128.400 ;
        RECT 547.950 125.400 570.600 126.600 ;
        RECT 724.950 126.600 727.050 127.050 ;
        RECT 808.950 126.600 811.050 127.050 ;
        RECT 724.950 125.400 811.050 126.600 ;
        RECT 547.950 124.950 550.050 125.400 ;
        RECT 724.950 124.950 727.050 125.400 ;
        RECT 808.950 124.950 811.050 125.400 ;
        RECT 838.950 126.600 841.050 127.050 ;
        RECT 850.950 126.600 853.050 127.050 ;
        RECT 838.950 125.400 853.050 126.600 ;
        RECT 838.950 124.950 841.050 125.400 ;
        RECT 850.950 124.950 853.050 125.400 ;
        RECT 22.950 123.600 25.050 124.050 ;
        RECT 49.950 123.600 52.050 124.050 ;
        RECT 88.950 123.600 91.050 124.050 ;
        RECT 22.950 122.400 91.050 123.600 ;
        RECT 22.950 121.950 25.050 122.400 ;
        RECT 49.950 121.950 52.050 122.400 ;
        RECT 88.950 121.950 91.050 122.400 ;
        RECT 103.950 123.600 106.050 124.050 ;
        RECT 127.950 123.600 130.050 124.050 ;
        RECT 103.950 122.400 130.050 123.600 ;
        RECT 103.950 121.950 106.050 122.400 ;
        RECT 127.950 121.950 130.050 122.400 ;
        RECT 199.950 123.600 202.050 124.050 ;
        RECT 328.950 123.600 331.050 124.050 ;
        RECT 343.950 123.600 346.050 124.050 ;
        RECT 421.800 123.600 423.900 124.050 ;
        RECT 199.950 122.400 210.600 123.600 ;
        RECT 199.950 121.950 202.050 122.400 ;
        RECT 25.950 120.600 28.050 121.050 ;
        RECT 34.950 120.600 37.050 121.050 ;
        RECT 40.950 120.600 43.050 121.050 ;
        RECT 73.950 120.600 76.050 121.050 ;
        RECT 25.950 119.400 76.050 120.600 ;
        RECT 25.950 118.950 28.050 119.400 ;
        RECT 34.950 118.950 37.050 119.400 ;
        RECT 40.950 118.950 43.050 119.400 ;
        RECT 73.950 118.950 76.050 119.400 ;
        RECT 109.950 120.600 112.050 121.050 ;
        RECT 121.950 120.600 124.050 121.050 ;
        RECT 109.950 119.400 124.050 120.600 ;
        RECT 109.950 118.950 112.050 119.400 ;
        RECT 121.950 118.950 124.050 119.400 ;
        RECT 133.950 120.600 136.050 121.050 ;
        RECT 209.400 120.600 210.600 122.400 ;
        RECT 328.950 122.400 346.050 123.600 ;
        RECT 328.950 121.950 331.050 122.400 ;
        RECT 343.950 121.950 346.050 122.400 ;
        RECT 362.400 122.400 423.900 123.600 ;
        RECT 235.950 120.600 238.050 121.050 ;
        RECT 133.950 119.400 177.600 120.600 ;
        RECT 209.400 119.400 238.050 120.600 ;
        RECT 133.950 118.950 136.050 119.400 ;
        RECT 176.400 118.050 177.600 119.400 ;
        RECT 235.950 118.950 238.050 119.400 ;
        RECT 253.950 120.600 256.050 121.050 ;
        RECT 274.950 120.600 277.050 121.050 ;
        RECT 253.950 119.400 277.050 120.600 ;
        RECT 253.950 118.950 256.050 119.400 ;
        RECT 274.950 118.950 277.050 119.400 ;
        RECT 304.950 120.600 307.050 121.050 ;
        RECT 319.950 120.600 322.050 121.050 ;
        RECT 304.950 119.400 322.050 120.600 ;
        RECT 304.950 118.950 307.050 119.400 ;
        RECT 319.950 118.950 322.050 119.400 ;
        RECT 331.950 120.600 334.050 121.050 ;
        RECT 362.400 120.600 363.600 122.400 ;
        RECT 421.800 121.950 423.900 122.400 ;
        RECT 424.950 123.600 427.050 124.050 ;
        RECT 448.950 123.600 451.050 124.050 ;
        RECT 424.950 122.400 451.050 123.600 ;
        RECT 424.950 121.950 427.050 122.400 ;
        RECT 448.950 121.950 451.050 122.400 ;
        RECT 514.950 123.600 517.050 124.050 ;
        RECT 544.950 123.600 547.050 124.050 ;
        RECT 562.950 123.600 565.050 124.050 ;
        RECT 571.950 123.600 574.050 124.050 ;
        RECT 514.950 122.400 574.050 123.600 ;
        RECT 514.950 121.950 517.050 122.400 ;
        RECT 544.950 121.950 547.050 122.400 ;
        RECT 562.950 121.950 565.050 122.400 ;
        RECT 571.950 121.950 574.050 122.400 ;
        RECT 643.950 123.600 646.050 124.050 ;
        RECT 772.950 123.600 775.050 124.050 ;
        RECT 784.950 123.600 787.050 124.050 ;
        RECT 643.950 122.400 660.600 123.600 ;
        RECT 643.950 121.950 646.050 122.400 ;
        RECT 331.950 119.400 363.600 120.600 ;
        RECT 376.950 120.600 379.050 121.050 ;
        RECT 439.950 120.600 442.050 121.050 ;
        RECT 469.950 120.600 472.050 121.050 ;
        RECT 376.950 119.400 472.050 120.600 ;
        RECT 331.950 118.950 334.050 119.400 ;
        RECT 376.950 118.950 379.050 119.400 ;
        RECT 439.950 118.950 442.050 119.400 ;
        RECT 469.950 118.950 472.050 119.400 ;
        RECT 580.950 120.600 583.050 121.050 ;
        RECT 622.950 120.600 625.050 121.050 ;
        RECT 580.950 119.400 625.050 120.600 ;
        RECT 659.400 120.600 660.600 122.400 ;
        RECT 772.950 122.400 787.050 123.600 ;
        RECT 772.950 121.950 775.050 122.400 ;
        RECT 784.950 121.950 787.050 122.400 ;
        RECT 685.950 120.600 688.050 121.050 ;
        RECT 659.400 119.400 688.050 120.600 ;
        RECT 580.950 118.950 583.050 119.400 ;
        RECT 622.950 118.950 625.050 119.400 ;
        RECT 685.950 118.950 688.050 119.400 ;
        RECT 694.950 120.600 697.050 121.050 ;
        RECT 721.950 120.600 724.050 121.050 ;
        RECT 694.950 119.400 724.050 120.600 ;
        RECT 694.950 118.950 697.050 119.400 ;
        RECT 721.950 118.950 724.050 119.400 ;
        RECT 793.950 120.600 796.050 121.050 ;
        RECT 805.950 120.600 808.050 121.050 ;
        RECT 832.950 120.600 835.050 121.050 ;
        RECT 793.950 119.400 835.050 120.600 ;
        RECT 793.950 118.950 796.050 119.400 ;
        RECT 805.950 118.950 808.050 119.400 ;
        RECT 832.950 118.950 835.050 119.400 ;
        RECT 844.950 120.600 847.050 121.050 ;
        RECT 853.950 120.600 856.050 121.050 ;
        RECT 844.950 119.400 856.050 120.600 ;
        RECT 844.950 118.950 847.050 119.400 ;
        RECT 853.950 118.950 856.050 119.400 ;
        RECT 16.950 117.600 19.050 118.050 ;
        RECT 28.950 117.600 31.050 118.050 ;
        RECT 16.950 116.400 31.050 117.600 ;
        RECT 16.950 115.950 19.050 116.400 ;
        RECT 28.950 115.950 31.050 116.400 ;
        RECT 145.950 117.600 148.050 118.050 ;
        RECT 175.950 117.600 178.050 118.050 ;
        RECT 193.950 117.600 196.050 118.050 ;
        RECT 205.950 117.600 208.050 118.050 ;
        RECT 145.950 116.400 165.600 117.600 ;
        RECT 145.950 115.950 148.050 116.400 ;
        RECT 164.400 115.050 165.600 116.400 ;
        RECT 175.950 116.400 208.050 117.600 ;
        RECT 175.950 115.950 178.050 116.400 ;
        RECT 193.950 115.950 196.050 116.400 ;
        RECT 205.950 115.950 208.050 116.400 ;
        RECT 268.950 117.600 271.050 118.050 ;
        RECT 280.950 117.600 283.050 118.050 ;
        RECT 292.950 117.600 295.050 118.050 ;
        RECT 268.950 116.400 295.050 117.600 ;
        RECT 268.950 115.950 271.050 116.400 ;
        RECT 280.950 115.950 283.050 116.400 ;
        RECT 292.950 115.950 295.050 116.400 ;
        RECT 478.950 117.600 481.050 118.050 ;
        RECT 520.950 117.600 523.050 118.050 ;
        RECT 478.950 116.400 523.050 117.600 ;
        RECT 478.950 115.950 481.050 116.400 ;
        RECT 520.950 115.950 523.050 116.400 ;
        RECT 535.950 117.600 538.050 118.050 ;
        RECT 553.950 117.600 556.050 118.050 ;
        RECT 535.950 116.400 556.050 117.600 ;
        RECT 535.950 115.950 538.050 116.400 ;
        RECT 553.950 115.950 556.050 116.400 ;
        RECT 808.950 117.600 811.050 118.050 ;
        RECT 823.950 117.600 826.050 118.050 ;
        RECT 808.950 116.400 826.050 117.600 ;
        RECT 808.950 115.950 811.050 116.400 ;
        RECT 823.950 115.950 826.050 116.400 ;
        RECT 835.950 117.600 838.050 118.050 ;
        RECT 841.950 117.600 844.050 118.050 ;
        RECT 835.950 116.400 844.050 117.600 ;
        RECT 835.950 115.950 838.050 116.400 ;
        RECT 841.950 115.950 844.050 116.400 ;
        RECT 52.950 114.600 55.050 115.050 ;
        RECT 58.950 114.600 61.050 115.050 ;
        RECT 94.950 114.600 97.050 115.050 ;
        RECT 52.950 113.400 97.050 114.600 ;
        RECT 52.950 112.950 55.050 113.400 ;
        RECT 58.950 112.950 61.050 113.400 ;
        RECT 94.950 112.950 97.050 113.400 ;
        RECT 124.950 114.600 127.050 115.050 ;
        RECT 130.950 114.600 133.050 115.050 ;
        RECT 160.800 114.600 162.900 115.050 ;
        RECT 124.950 113.400 133.050 114.600 ;
        RECT 124.950 112.950 127.050 113.400 ;
        RECT 130.950 112.950 133.050 113.400 ;
        RECT 134.400 113.400 162.900 114.600 ;
        RECT 10.950 111.600 13.050 112.050 ;
        RECT 31.950 111.600 34.050 112.050 ;
        RECT 10.950 110.400 34.050 111.600 ;
        RECT 10.950 109.950 13.050 110.400 ;
        RECT 31.950 109.950 34.050 110.400 ;
        RECT 112.950 111.600 115.050 112.050 ;
        RECT 121.950 111.600 124.050 112.050 ;
        RECT 112.950 110.400 124.050 111.600 ;
        RECT 112.950 109.950 115.050 110.400 ;
        RECT 121.950 109.950 124.050 110.400 ;
        RECT 127.950 111.600 130.050 112.050 ;
        RECT 134.400 111.600 135.600 113.400 ;
        RECT 160.800 112.950 162.900 113.400 ;
        RECT 163.950 114.600 166.050 115.050 ;
        RECT 172.950 114.600 175.050 115.050 ;
        RECT 163.950 113.400 175.050 114.600 ;
        RECT 163.950 112.950 166.050 113.400 ;
        RECT 172.950 112.950 175.050 113.400 ;
        RECT 211.950 114.600 214.050 115.050 ;
        RECT 220.950 114.600 223.050 115.050 ;
        RECT 211.950 113.400 223.050 114.600 ;
        RECT 211.950 112.950 214.050 113.400 ;
        RECT 220.950 112.950 223.050 113.400 ;
        RECT 250.950 114.600 253.050 115.050 ;
        RECT 256.950 114.600 259.050 115.050 ;
        RECT 250.950 113.400 259.050 114.600 ;
        RECT 250.950 112.950 253.050 113.400 ;
        RECT 256.950 112.950 259.050 113.400 ;
        RECT 265.950 114.600 268.050 115.050 ;
        RECT 280.950 114.600 283.050 114.900 ;
        RECT 265.950 113.400 283.050 114.600 ;
        RECT 265.950 112.950 268.050 113.400 ;
        RECT 280.950 112.800 283.050 113.400 ;
        RECT 295.950 114.600 298.050 115.050 ;
        RECT 322.950 114.600 325.050 115.050 ;
        RECT 355.950 114.600 358.050 115.050 ;
        RECT 295.950 113.400 358.050 114.600 ;
        RECT 295.950 112.950 298.050 113.400 ;
        RECT 322.950 112.950 325.050 113.400 ;
        RECT 355.950 112.950 358.050 113.400 ;
        RECT 361.950 114.600 364.050 115.050 ;
        RECT 373.950 114.600 376.050 115.050 ;
        RECT 361.950 113.400 376.050 114.600 ;
        RECT 361.950 112.950 364.050 113.400 ;
        RECT 373.950 112.950 376.050 113.400 ;
        RECT 385.950 114.600 388.050 115.050 ;
        RECT 403.950 114.600 406.050 115.050 ;
        RECT 385.950 113.400 406.050 114.600 ;
        RECT 385.950 112.950 388.050 113.400 ;
        RECT 403.950 112.950 406.050 113.400 ;
        RECT 409.950 114.600 412.050 115.050 ;
        RECT 418.950 114.600 421.050 115.050 ;
        RECT 436.950 114.600 439.050 115.050 ;
        RECT 448.950 114.600 451.050 115.050 ;
        RECT 409.950 113.400 429.600 114.600 ;
        RECT 409.950 112.950 412.050 113.400 ;
        RECT 418.950 112.950 421.050 113.400 ;
        RECT 127.950 110.400 135.600 111.600 ;
        RECT 157.950 111.600 160.050 112.050 ;
        RECT 169.950 111.600 172.050 112.050 ;
        RECT 157.950 110.400 172.050 111.600 ;
        RECT 127.950 109.950 130.050 110.400 ;
        RECT 157.950 109.950 160.050 110.400 ;
        RECT 169.950 109.950 172.050 110.400 ;
        RECT 184.950 111.600 187.050 112.050 ;
        RECT 196.950 111.600 199.050 112.050 ;
        RECT 184.950 110.400 199.050 111.600 ;
        RECT 184.950 109.950 187.050 110.400 ;
        RECT 196.950 109.950 199.050 110.400 ;
        RECT 208.950 111.600 211.050 112.050 ;
        RECT 235.950 111.600 238.050 112.050 ;
        RECT 208.950 110.400 238.050 111.600 ;
        RECT 208.950 109.950 211.050 110.400 ;
        RECT 235.950 109.950 238.050 110.400 ;
        RECT 241.950 111.600 244.050 112.050 ;
        RECT 262.950 111.600 265.050 112.050 ;
        RECT 289.950 111.600 292.050 112.050 ;
        RECT 424.950 111.600 427.050 112.050 ;
        RECT 241.950 110.400 292.050 111.600 ;
        RECT 241.950 109.950 244.050 110.400 ;
        RECT 262.950 109.950 265.050 110.400 ;
        RECT 289.950 109.950 292.050 110.400 ;
        RECT 392.400 110.400 427.050 111.600 ;
        RECT 428.400 111.600 429.600 113.400 ;
        RECT 436.950 113.400 451.050 114.600 ;
        RECT 436.950 112.950 439.050 113.400 ;
        RECT 448.950 112.950 451.050 113.400 ;
        RECT 496.950 114.600 499.050 115.050 ;
        RECT 505.800 114.600 507.900 115.050 ;
        RECT 496.950 113.400 507.900 114.600 ;
        RECT 496.950 112.950 499.050 113.400 ;
        RECT 505.800 112.950 507.900 113.400 ;
        RECT 508.950 114.600 511.050 115.050 ;
        RECT 532.950 114.600 535.050 115.050 ;
        RECT 508.950 113.400 535.050 114.600 ;
        RECT 508.950 112.950 511.050 113.400 ;
        RECT 532.950 112.950 535.050 113.400 ;
        RECT 538.950 114.600 541.050 115.050 ;
        RECT 544.950 114.600 547.050 115.050 ;
        RECT 538.950 113.400 547.050 114.600 ;
        RECT 538.950 112.950 541.050 113.400 ;
        RECT 544.950 112.950 547.050 113.400 ;
        RECT 556.950 114.600 559.050 115.050 ;
        RECT 601.950 114.600 604.050 115.050 ;
        RECT 640.950 114.600 643.050 115.050 ;
        RECT 556.950 113.400 643.050 114.600 ;
        RECT 556.950 112.950 559.050 113.400 ;
        RECT 601.950 112.950 604.050 113.400 ;
        RECT 640.950 112.950 643.050 113.400 ;
        RECT 679.950 114.600 682.050 115.050 ;
        RECT 727.950 114.600 730.050 115.050 ;
        RECT 679.950 113.400 730.050 114.600 ;
        RECT 679.950 112.950 682.050 113.400 ;
        RECT 727.950 112.950 730.050 113.400 ;
        RECT 736.950 114.600 739.050 115.050 ;
        RECT 765.000 114.600 768.900 115.050 ;
        RECT 736.950 113.400 768.900 114.600 ;
        RECT 736.950 112.950 739.050 113.400 ;
        RECT 764.400 112.950 768.900 113.400 ;
        RECT 769.950 114.600 772.050 115.050 ;
        RECT 778.950 114.600 781.050 115.050 ;
        RECT 769.950 113.400 781.050 114.600 ;
        RECT 769.950 112.950 772.050 113.400 ;
        RECT 778.950 112.950 781.050 113.400 ;
        RECT 802.950 114.600 805.050 115.050 ;
        RECT 826.950 114.600 829.050 115.050 ;
        RECT 802.950 113.400 829.050 114.600 ;
        RECT 802.950 112.950 805.050 113.400 ;
        RECT 826.950 112.950 829.050 113.400 ;
        RECT 445.950 111.600 448.050 112.050 ;
        RECT 428.400 110.400 448.050 111.600 ;
        RECT 46.950 108.600 49.050 109.050 ;
        RECT 32.400 107.400 49.050 108.600 ;
        RECT 22.950 105.600 27.000 106.050 ;
        RECT 22.950 103.950 27.600 105.600 ;
        RECT 13.950 99.600 16.050 99.900 ;
        RECT 19.950 99.600 22.050 100.050 ;
        RECT 26.400 99.900 27.600 103.950 ;
        RECT 32.400 99.900 33.600 107.400 ;
        RECT 46.950 106.950 49.050 107.400 ;
        RECT 52.950 108.600 55.050 109.050 ;
        RECT 67.950 108.600 70.050 109.050 ;
        RECT 52.950 107.400 70.050 108.600 ;
        RECT 52.950 106.950 55.050 107.400 ;
        RECT 67.950 106.950 70.050 107.400 ;
        RECT 73.950 108.600 76.050 109.050 ;
        RECT 103.950 108.600 106.050 109.050 ;
        RECT 73.950 107.400 106.050 108.600 ;
        RECT 73.950 106.950 76.050 107.400 ;
        RECT 103.950 106.950 106.050 107.400 ;
        RECT 151.950 108.600 154.050 109.050 ;
        RECT 199.950 108.600 202.050 109.050 ;
        RECT 265.950 108.600 268.050 109.050 ;
        RECT 151.950 107.400 159.600 108.600 ;
        RECT 151.950 106.950 154.050 107.400 ;
        RECT 34.950 105.600 37.050 106.200 ;
        RECT 49.950 105.600 52.050 106.200 ;
        RECT 94.950 105.750 97.050 106.200 ;
        RECT 100.950 105.750 103.050 106.200 ;
        RECT 34.950 104.400 39.600 105.600 ;
        RECT 34.950 104.100 37.050 104.400 ;
        RECT 38.400 100.050 39.600 104.400 ;
        RECT 49.950 104.400 60.600 105.600 ;
        RECT 49.950 104.100 52.050 104.400 ;
        RECT 13.950 98.400 22.050 99.600 ;
        RECT 13.950 97.800 16.050 98.400 ;
        RECT 19.950 97.950 22.050 98.400 ;
        RECT 25.950 97.800 28.050 99.900 ;
        RECT 31.950 97.800 34.050 99.900 ;
        RECT 37.950 97.950 40.050 100.050 ;
        RECT 59.400 99.600 60.600 104.400 ;
        RECT 94.950 104.550 103.050 105.750 ;
        RECT 94.950 104.100 97.050 104.550 ;
        RECT 100.950 104.100 103.050 104.550 ;
        RECT 106.950 105.600 109.050 106.050 ;
        RECT 112.950 105.600 115.050 106.200 ;
        RECT 106.950 104.400 115.050 105.600 ;
        RECT 106.950 103.950 109.050 104.400 ;
        RECT 112.950 104.100 115.050 104.400 ;
        RECT 118.950 104.100 121.050 106.200 ;
        RECT 154.950 105.600 157.050 106.050 ;
        RECT 143.400 104.400 157.050 105.600 ;
        RECT 119.400 102.600 120.600 104.100 ;
        RECT 139.950 102.600 142.050 103.050 ;
        RECT 119.400 101.400 142.050 102.600 ;
        RECT 139.950 100.950 142.050 101.400 ;
        RECT 143.400 100.050 144.600 104.400 ;
        RECT 154.950 103.950 157.050 104.400 ;
        RECT 79.950 99.600 82.050 100.050 ;
        RECT 59.400 98.400 82.050 99.600 ;
        RECT 79.950 97.950 82.050 98.400 ;
        RECT 97.950 99.450 100.050 99.900 ;
        RECT 103.950 99.450 106.050 99.900 ;
        RECT 97.950 98.250 106.050 99.450 ;
        RECT 97.950 97.800 100.050 98.250 ;
        RECT 103.950 97.800 106.050 98.250 ;
        RECT 142.950 97.950 145.050 100.050 ;
        RECT 158.400 99.600 159.600 107.400 ;
        RECT 194.400 107.400 202.050 108.600 ;
        RECT 181.950 105.600 184.050 106.050 ;
        RECT 190.950 105.600 193.050 106.200 ;
        RECT 181.950 104.400 193.050 105.600 ;
        RECT 181.950 103.950 184.050 104.400 ;
        RECT 190.950 104.100 193.050 104.400 ;
        RECT 194.400 99.900 195.600 107.400 ;
        RECT 199.950 106.950 202.050 107.400 ;
        RECT 224.400 107.400 268.050 108.600 ;
        RECT 196.950 105.750 199.050 106.200 ;
        RECT 202.800 105.750 204.900 106.200 ;
        RECT 196.950 104.550 204.900 105.750 ;
        RECT 196.950 104.100 199.050 104.550 ;
        RECT 202.800 104.100 204.900 104.550 ;
        RECT 205.950 105.750 208.050 106.200 ;
        RECT 214.950 105.750 217.050 106.200 ;
        RECT 205.950 104.550 217.050 105.750 ;
        RECT 205.950 104.100 208.050 104.550 ;
        RECT 214.950 104.100 217.050 104.550 ;
        RECT 203.400 102.600 204.600 104.100 ;
        RECT 203.400 101.400 216.600 102.600 ;
        RECT 166.950 99.600 169.050 99.900 ;
        RECT 158.400 98.400 169.050 99.600 ;
        RECT 166.950 97.800 169.050 98.400 ;
        RECT 172.950 99.450 175.050 99.900 ;
        RECT 184.950 99.450 187.050 99.900 ;
        RECT 172.950 98.250 187.050 99.450 ;
        RECT 172.950 97.800 175.050 98.250 ;
        RECT 184.950 97.800 187.050 98.250 ;
        RECT 193.950 97.800 196.050 99.900 ;
        RECT 215.400 99.600 216.600 101.400 ;
        RECT 224.400 99.900 225.600 107.400 ;
        RECT 265.950 106.950 268.050 107.400 ;
        RECT 307.950 108.600 310.050 109.050 ;
        RECT 325.950 108.600 328.050 109.050 ;
        RECT 334.950 108.600 337.050 109.050 ;
        RECT 307.950 107.400 328.050 108.600 ;
        RECT 307.950 106.950 310.050 107.400 ;
        RECT 325.950 106.950 328.050 107.400 ;
        RECT 329.400 107.400 337.050 108.600 ;
        RECT 267.000 105.600 271.050 106.050 ;
        RECT 286.950 105.600 289.050 106.200 ;
        RECT 239.400 104.400 271.050 105.600 ;
        RECT 239.400 99.900 240.600 104.400 ;
        RECT 266.400 103.950 271.050 104.400 ;
        RECT 278.400 104.400 289.050 105.600 ;
        RECT 266.400 99.900 267.600 103.950 ;
        RECT 278.400 100.050 279.600 104.400 ;
        RECT 286.950 104.100 289.050 104.400 ;
        RECT 292.950 103.950 295.050 106.050 ;
        RECT 313.950 105.600 316.050 106.050 ;
        RECT 329.400 105.600 330.600 107.400 ;
        RECT 334.950 106.950 337.050 107.400 ;
        RECT 313.950 104.400 330.600 105.600 ;
        RECT 313.950 103.950 316.050 104.400 ;
        RECT 337.950 103.950 340.050 106.050 ;
        RECT 346.950 103.950 349.050 106.050 ;
        RECT 367.950 105.600 370.050 106.200 ;
        RECT 385.950 105.600 388.050 106.200 ;
        RECT 367.950 104.400 388.050 105.600 ;
        RECT 367.950 104.100 370.050 104.400 ;
        RECT 385.950 104.100 388.050 104.400 ;
        RECT 217.950 99.600 220.050 99.900 ;
        RECT 215.400 98.400 220.050 99.600 ;
        RECT 217.950 97.800 220.050 98.400 ;
        RECT 223.950 97.800 226.050 99.900 ;
        RECT 238.950 97.800 241.050 99.900 ;
        RECT 244.950 99.600 247.050 99.900 ;
        RECT 259.950 99.600 262.050 99.900 ;
        RECT 244.950 98.400 262.050 99.600 ;
        RECT 244.950 97.800 247.050 98.400 ;
        RECT 259.950 97.800 262.050 98.400 ;
        RECT 265.950 97.800 268.050 99.900 ;
        RECT 277.950 97.950 280.050 100.050 ;
        RECT 289.950 99.600 292.050 99.900 ;
        RECT 293.400 99.600 294.600 103.950 ;
        RECT 289.950 98.400 294.600 99.600 ;
        RECT 295.950 99.450 298.050 99.900 ;
        RECT 304.950 99.450 307.050 99.900 ;
        RECT 289.950 97.800 292.050 98.400 ;
        RECT 295.950 98.250 307.050 99.450 ;
        RECT 295.950 97.800 298.050 98.250 ;
        RECT 304.950 97.800 307.050 98.250 ;
        RECT 334.950 99.600 337.050 99.900 ;
        RECT 338.400 99.600 339.600 103.950 ;
        RECT 334.950 98.400 339.600 99.600 ;
        RECT 347.400 99.600 348.600 103.950 ;
        RECT 373.950 99.600 376.050 100.050 ;
        RECT 347.400 98.400 376.050 99.600 ;
        RECT 334.950 97.800 337.050 98.400 ;
        RECT 373.950 97.950 376.050 98.400 ;
        RECT 388.950 99.600 391.050 99.900 ;
        RECT 392.400 99.600 393.600 110.400 ;
        RECT 424.950 109.950 427.050 110.400 ;
        RECT 445.950 109.950 448.050 110.400 ;
        RECT 451.950 111.600 454.050 112.050 ;
        RECT 490.950 111.600 493.050 111.900 ;
        RECT 553.950 111.600 556.050 112.050 ;
        RECT 451.950 110.400 493.050 111.600 ;
        RECT 451.950 109.950 454.050 110.400 ;
        RECT 427.950 105.750 430.050 106.200 ;
        RECT 439.950 105.750 442.050 106.200 ;
        RECT 427.950 104.550 442.050 105.750 ;
        RECT 427.950 104.100 430.050 104.550 ;
        RECT 439.950 104.100 442.050 104.550 ;
        RECT 448.950 104.100 451.050 106.200 ;
        RECT 418.950 102.600 423.000 103.050 ;
        RECT 418.950 100.950 423.600 102.600 ;
        RECT 388.950 98.400 393.600 99.600 ;
        RECT 422.400 99.600 423.600 100.950 ;
        RECT 424.950 99.600 427.050 99.900 ;
        RECT 422.400 98.400 427.050 99.600 ;
        RECT 388.950 97.800 391.050 98.400 ;
        RECT 424.950 97.800 427.050 98.400 ;
        RECT 430.950 99.450 433.050 99.900 ;
        RECT 436.950 99.600 439.050 99.900 ;
        RECT 449.400 99.600 450.600 104.100 ;
        RECT 452.400 99.900 453.600 109.950 ;
        RECT 490.950 109.800 493.050 110.400 ;
        RECT 509.400 110.400 556.050 111.600 ;
        RECT 502.950 108.600 505.050 109.050 ;
        RECT 509.400 108.600 510.600 110.400 ;
        RECT 553.950 109.950 556.050 110.400 ;
        RECT 568.950 111.600 571.050 112.050 ;
        RECT 598.950 111.600 601.050 112.050 ;
        RECT 568.950 110.400 601.050 111.600 ;
        RECT 568.950 109.950 571.050 110.400 ;
        RECT 598.950 109.950 601.050 110.400 ;
        RECT 607.950 111.600 610.050 112.050 ;
        RECT 622.950 111.600 625.050 112.050 ;
        RECT 760.950 111.600 763.050 112.050 ;
        RECT 607.950 110.400 763.050 111.600 ;
        RECT 764.400 111.600 765.600 112.950 ;
        RECT 793.950 111.600 796.050 112.050 ;
        RECT 764.400 110.400 796.050 111.600 ;
        RECT 607.950 109.950 610.050 110.400 ;
        RECT 622.950 109.950 625.050 110.400 ;
        RECT 760.950 109.950 763.050 110.400 ;
        RECT 793.950 109.950 796.050 110.400 ;
        RECT 494.400 107.400 510.600 108.600 ;
        RECT 511.950 108.600 514.050 109.050 ;
        RECT 517.950 108.600 520.050 109.050 ;
        RECT 511.950 107.400 520.050 108.600 ;
        RECT 454.950 105.600 457.050 106.200 ;
        RECT 475.950 105.600 478.050 106.200 ;
        RECT 454.950 104.400 474.600 105.600 ;
        RECT 454.950 104.100 457.050 104.400 ;
        RECT 473.400 102.600 474.600 104.400 ;
        RECT 475.950 104.400 489.600 105.600 ;
        RECT 475.950 104.100 478.050 104.400 ;
        RECT 473.400 101.400 480.600 102.600 ;
        RECT 479.400 99.900 480.600 101.400 ;
        RECT 488.400 100.050 489.600 104.400 ;
        RECT 436.950 99.450 450.600 99.600 ;
        RECT 430.950 98.400 450.600 99.450 ;
        RECT 430.950 98.250 439.050 98.400 ;
        RECT 430.950 97.800 433.050 98.250 ;
        RECT 436.950 97.800 439.050 98.250 ;
        RECT 451.950 97.800 454.050 99.900 ;
        RECT 478.950 97.800 481.050 99.900 ;
        RECT 487.950 97.950 490.050 100.050 ;
        RECT 494.400 99.900 495.600 107.400 ;
        RECT 502.950 106.950 505.050 107.400 ;
        RECT 511.950 106.950 514.050 107.400 ;
        RECT 517.950 106.950 520.050 107.400 ;
        RECT 496.950 105.600 499.050 106.200 ;
        RECT 529.950 105.600 532.050 106.200 ;
        RECT 496.950 104.400 532.050 105.600 ;
        RECT 496.950 104.100 499.050 104.400 ;
        RECT 512.400 99.900 513.600 104.400 ;
        RECT 529.950 104.100 532.050 104.400 ;
        RECT 535.950 104.100 538.050 106.200 ;
        RECT 589.950 104.100 592.050 106.200 ;
        RECT 610.950 104.100 613.050 106.200 ;
        RECT 616.950 105.600 619.050 106.200 ;
        RECT 628.950 105.600 631.050 106.200 ;
        RECT 616.950 104.400 631.050 105.600 ;
        RECT 616.950 104.100 619.050 104.400 ;
        RECT 628.950 104.100 631.050 104.400 ;
        RECT 634.950 104.100 637.050 106.200 ;
        RECT 640.950 105.600 643.050 106.050 ;
        RECT 655.950 105.600 658.050 106.200 ;
        RECT 667.950 105.600 670.050 109.050 ;
        RECT 700.950 108.600 703.050 109.200 ;
        RECT 706.950 108.600 709.050 109.050 ;
        RECT 700.950 107.400 709.050 108.600 ;
        RECT 700.950 107.100 703.050 107.400 ;
        RECT 706.950 106.950 709.050 107.400 ;
        RECT 763.950 108.600 766.050 109.050 ;
        RECT 775.950 108.600 778.050 109.050 ;
        RECT 790.950 108.600 793.050 109.050 ;
        RECT 763.950 107.400 793.050 108.600 ;
        RECT 763.950 106.950 766.050 107.400 ;
        RECT 775.950 106.950 778.050 107.400 ;
        RECT 790.950 106.950 793.050 107.400 ;
        RECT 799.950 108.600 802.050 109.050 ;
        RECT 811.800 108.600 813.900 109.050 ;
        RECT 799.950 107.400 813.900 108.600 ;
        RECT 799.950 106.950 802.050 107.400 ;
        RECT 811.800 106.950 813.900 107.400 ;
        RECT 673.950 105.600 676.050 106.200 ;
        RECT 640.950 104.400 654.600 105.600 ;
        RECT 536.400 102.600 537.600 104.100 ;
        RECT 590.400 102.600 591.600 104.100 ;
        RECT 611.400 102.600 612.600 104.100 ;
        RECT 635.400 102.600 636.600 104.100 ;
        RECT 640.950 103.950 643.050 104.400 ;
        RECT 536.400 101.400 558.600 102.600 ;
        RECT 590.400 102.000 597.600 102.600 ;
        RECT 590.400 101.400 598.050 102.000 ;
        RECT 611.400 101.400 618.600 102.600 ;
        RECT 635.400 102.000 648.600 102.600 ;
        RECT 635.400 101.400 649.050 102.000 ;
        RECT 557.400 99.900 558.600 101.400 ;
        RECT 493.950 97.800 496.050 99.900 ;
        RECT 511.950 97.800 514.050 99.900 ;
        RECT 538.950 99.600 541.050 99.900 ;
        RECT 550.950 99.600 553.050 99.900 ;
        RECT 538.950 98.400 553.050 99.600 ;
        RECT 538.950 97.800 541.050 98.400 ;
        RECT 550.950 97.800 553.050 98.400 ;
        RECT 556.950 97.800 559.050 99.900 ;
        RECT 580.950 99.450 583.050 99.900 ;
        RECT 586.950 99.450 589.050 99.900 ;
        RECT 580.950 98.250 589.050 99.450 ;
        RECT 580.950 97.800 583.050 98.250 ;
        RECT 586.950 97.800 589.050 98.250 ;
        RECT 595.950 97.950 598.050 101.400 ;
        RECT 617.400 100.050 618.600 101.400 ;
        RECT 601.950 99.450 604.050 99.900 ;
        RECT 607.950 99.450 610.050 99.900 ;
        RECT 601.950 98.250 610.050 99.450 ;
        RECT 617.400 98.400 622.050 100.050 ;
        RECT 601.950 97.800 604.050 98.250 ;
        RECT 607.950 97.800 610.050 98.250 ;
        RECT 618.000 97.950 622.050 98.400 ;
        RECT 646.950 97.950 649.050 101.400 ;
        RECT 653.400 99.900 654.600 104.400 ;
        RECT 655.950 104.400 676.050 105.600 ;
        RECT 655.950 104.100 658.050 104.400 ;
        RECT 673.950 104.100 676.050 104.400 ;
        RECT 700.950 105.600 703.050 106.050 ;
        RECT 712.950 105.600 715.050 106.200 ;
        RECT 700.950 104.400 715.050 105.600 ;
        RECT 700.950 103.950 703.050 104.400 ;
        RECT 712.950 104.100 715.050 104.400 ;
        RECT 718.950 105.600 721.050 106.200 ;
        RECT 736.950 105.600 739.050 106.200 ;
        RECT 718.950 104.400 739.050 105.600 ;
        RECT 718.950 104.100 721.050 104.400 ;
        RECT 736.950 104.100 739.050 104.400 ;
        RECT 742.950 105.600 745.050 106.200 ;
        RECT 748.950 105.600 751.050 106.050 ;
        RECT 757.950 105.600 760.050 106.200 ;
        RECT 742.950 104.400 751.050 105.600 ;
        RECT 742.950 104.100 745.050 104.400 ;
        RECT 748.950 103.950 751.050 104.400 ;
        RECT 752.400 104.400 760.050 105.600 ;
        RECT 752.400 102.600 753.600 104.400 ;
        RECT 757.950 104.100 760.050 104.400 ;
        RECT 781.950 105.600 784.050 106.200 ;
        RECT 793.950 105.600 796.050 106.050 ;
        RECT 808.950 105.600 811.050 106.050 ;
        RECT 781.950 104.400 792.600 105.600 ;
        RECT 781.950 104.100 784.050 104.400 ;
        RECT 740.400 101.400 753.600 102.600 ;
        RECT 791.400 102.600 792.600 104.400 ;
        RECT 793.950 104.400 811.050 105.600 ;
        RECT 814.950 105.600 817.050 109.050 ;
        RECT 823.950 108.600 826.050 109.050 ;
        RECT 838.950 108.600 841.050 109.050 ;
        RECT 823.950 107.400 841.050 108.600 ;
        RECT 823.950 106.950 826.050 107.400 ;
        RECT 838.950 106.950 841.050 107.400 ;
        RECT 820.950 105.600 823.050 106.200 ;
        RECT 814.950 105.000 823.050 105.600 ;
        RECT 815.400 104.400 823.050 105.000 ;
        RECT 793.950 103.950 796.050 104.400 ;
        RECT 808.950 102.600 811.050 104.400 ;
        RECT 820.950 104.100 823.050 104.400 ;
        RECT 826.950 105.600 829.050 106.200 ;
        RECT 844.950 105.600 847.050 106.200 ;
        RECT 826.950 104.400 831.600 105.600 ;
        RECT 826.950 104.100 829.050 104.400 ;
        RECT 791.400 101.400 807.600 102.600 ;
        RECT 808.950 102.000 822.600 102.600 ;
        RECT 809.400 101.400 822.600 102.000 ;
        RECT 740.400 99.900 741.600 101.400 ;
        RECT 652.950 97.800 655.050 99.900 ;
        RECT 658.950 99.450 661.050 99.900 ;
        RECT 664.950 99.600 667.050 99.900 ;
        RECT 676.950 99.600 679.050 99.900 ;
        RECT 664.950 99.450 679.050 99.600 ;
        RECT 658.950 98.400 679.050 99.450 ;
        RECT 658.950 98.250 667.050 98.400 ;
        RECT 658.950 97.800 661.050 98.250 ;
        RECT 664.950 97.800 667.050 98.250 ;
        RECT 676.950 97.800 679.050 98.400 ;
        RECT 721.950 99.600 724.050 99.900 ;
        RECT 739.950 99.600 742.050 99.900 ;
        RECT 721.950 98.400 742.050 99.600 ;
        RECT 721.950 97.800 724.050 98.400 ;
        RECT 739.950 97.800 742.050 98.400 ;
        RECT 760.950 99.600 763.050 99.900 ;
        RECT 769.950 99.600 772.050 99.900 ;
        RECT 760.950 99.450 772.050 99.600 ;
        RECT 778.950 99.450 781.050 99.900 ;
        RECT 760.950 98.400 781.050 99.450 ;
        RECT 806.400 99.600 807.600 101.400 ;
        RECT 814.950 99.600 817.050 100.050 ;
        RECT 806.400 98.400 817.050 99.600 ;
        RECT 760.950 97.800 763.050 98.400 ;
        RECT 769.950 98.250 781.050 98.400 ;
        RECT 769.950 97.800 772.050 98.250 ;
        RECT 778.950 97.800 781.050 98.250 ;
        RECT 814.950 97.950 817.050 98.400 ;
        RECT 82.950 96.600 85.050 97.050 ;
        RECT 91.950 96.600 94.050 97.050 ;
        RECT 82.950 95.400 94.050 96.600 ;
        RECT 82.950 94.950 85.050 95.400 ;
        RECT 91.950 94.950 94.050 95.400 ;
        RECT 109.950 96.600 112.050 97.050 ;
        RECT 124.950 96.600 127.050 97.050 ;
        RECT 130.950 96.600 133.050 97.050 ;
        RECT 109.950 95.400 133.050 96.600 ;
        RECT 109.950 94.950 112.050 95.400 ;
        RECT 124.950 94.950 127.050 95.400 ;
        RECT 130.950 94.950 133.050 95.400 ;
        RECT 157.950 96.600 160.050 97.050 ;
        RECT 163.950 96.600 166.050 97.050 ;
        RECT 296.400 96.600 297.600 97.800 ;
        RECT 821.400 97.050 822.600 101.400 ;
        RECT 830.400 99.600 831.600 104.400 ;
        RECT 844.950 104.400 852.600 105.600 ;
        RECT 844.950 104.100 847.050 104.400 ;
        RECT 851.400 100.050 852.600 104.400 ;
        RECT 830.400 98.400 846.600 99.600 ;
        RECT 845.400 97.050 846.600 98.400 ;
        RECT 850.950 97.950 853.050 100.050 ;
        RECT 859.950 99.600 862.050 99.900 ;
        RECT 868.950 99.600 871.050 100.050 ;
        RECT 859.950 98.400 871.050 99.600 ;
        RECT 859.950 97.800 862.050 98.400 ;
        RECT 868.950 97.950 871.050 98.400 ;
        RECT 157.950 95.400 166.050 96.600 ;
        RECT 157.950 94.950 160.050 95.400 ;
        RECT 163.950 94.950 166.050 95.400 ;
        RECT 263.400 95.400 297.600 96.600 ;
        RECT 322.950 96.600 325.050 97.050 ;
        RECT 442.950 96.600 445.050 97.050 ;
        RECT 457.950 96.600 460.050 97.050 ;
        RECT 322.950 96.000 333.600 96.600 ;
        RECT 322.950 95.400 334.050 96.000 ;
        RECT 263.400 94.050 264.600 95.400 ;
        RECT 322.950 94.950 325.050 95.400 ;
        RECT 76.950 93.600 79.050 94.050 ;
        RECT 100.950 93.600 103.050 94.050 ;
        RECT 76.950 92.400 103.050 93.600 ;
        RECT 76.950 91.950 79.050 92.400 ;
        RECT 100.950 91.950 103.050 92.400 ;
        RECT 139.950 93.600 142.050 94.050 ;
        RECT 172.950 93.600 175.050 94.050 ;
        RECT 139.950 92.400 175.050 93.600 ;
        RECT 139.950 91.950 142.050 92.400 ;
        RECT 172.950 91.950 175.050 92.400 ;
        RECT 223.950 93.600 226.050 94.050 ;
        RECT 223.950 92.400 258.600 93.600 ;
        RECT 223.950 91.950 226.050 92.400 ;
        RECT 115.950 90.600 118.050 91.050 ;
        RECT 121.950 90.600 124.050 91.050 ;
        RECT 148.950 90.600 151.050 91.050 ;
        RECT 115.950 89.400 151.050 90.600 ;
        RECT 115.950 88.950 118.050 89.400 ;
        RECT 121.950 88.950 124.050 89.400 ;
        RECT 148.950 88.950 151.050 89.400 ;
        RECT 178.950 90.600 181.050 91.050 ;
        RECT 250.950 90.600 253.050 91.050 ;
        RECT 178.950 89.400 253.050 90.600 ;
        RECT 257.400 90.600 258.600 92.400 ;
        RECT 259.950 92.400 264.600 94.050 ;
        RECT 283.950 93.600 286.050 94.050 ;
        RECT 325.950 93.600 328.050 94.050 ;
        RECT 283.950 92.400 328.050 93.600 ;
        RECT 259.950 91.950 264.000 92.400 ;
        RECT 283.950 91.950 286.050 92.400 ;
        RECT 325.950 91.950 328.050 92.400 ;
        RECT 331.950 91.950 334.050 95.400 ;
        RECT 442.950 95.400 460.050 96.600 ;
        RECT 442.950 94.950 445.050 95.400 ;
        RECT 457.950 94.950 460.050 95.400 ;
        RECT 499.950 96.600 502.050 97.050 ;
        RECT 505.950 96.600 508.050 97.050 ;
        RECT 526.950 96.600 529.050 97.050 ;
        RECT 499.950 95.400 529.050 96.600 ;
        RECT 499.950 94.950 502.050 95.400 ;
        RECT 505.950 94.950 508.050 95.400 ;
        RECT 526.950 94.950 529.050 95.400 ;
        RECT 790.950 96.600 793.050 97.050 ;
        RECT 805.950 96.600 808.050 97.050 ;
        RECT 790.950 95.400 808.050 96.600 ;
        RECT 790.950 94.950 793.050 95.400 ;
        RECT 805.950 94.950 808.050 95.400 ;
        RECT 820.950 94.950 823.050 97.050 ;
        RECT 845.400 95.400 850.050 97.050 ;
        RECT 846.000 94.950 850.050 95.400 ;
        RECT 412.950 93.600 415.050 94.050 ;
        RECT 439.950 93.600 442.050 94.050 ;
        RECT 445.950 93.600 448.050 94.050 ;
        RECT 502.950 93.600 505.050 94.050 ;
        RECT 412.950 92.400 505.050 93.600 ;
        RECT 412.950 91.950 415.050 92.400 ;
        RECT 439.950 91.950 442.050 92.400 ;
        RECT 445.950 91.950 448.050 92.400 ;
        RECT 502.950 91.950 505.050 92.400 ;
        RECT 508.950 93.600 511.050 94.050 ;
        RECT 517.950 93.600 520.050 94.050 ;
        RECT 508.950 92.400 520.050 93.600 ;
        RECT 508.950 91.950 511.050 92.400 ;
        RECT 517.950 91.950 520.050 92.400 ;
        RECT 697.950 93.600 700.050 94.050 ;
        RECT 736.950 93.600 739.050 94.050 ;
        RECT 697.950 92.400 739.050 93.600 ;
        RECT 697.950 91.950 700.050 92.400 ;
        RECT 736.950 91.950 739.050 92.400 ;
        RECT 817.950 93.600 820.050 94.050 ;
        RECT 829.950 93.600 832.050 94.050 ;
        RECT 817.950 92.400 832.050 93.600 ;
        RECT 817.950 91.950 820.050 92.400 ;
        RECT 829.950 91.950 832.050 92.400 ;
        RECT 835.950 93.600 838.050 94.050 ;
        RECT 853.950 93.600 856.050 94.050 ;
        RECT 835.950 92.400 856.050 93.600 ;
        RECT 835.950 91.950 838.050 92.400 ;
        RECT 853.950 91.950 856.050 92.400 ;
        RECT 271.950 90.600 274.050 91.050 ;
        RECT 257.400 89.400 274.050 90.600 ;
        RECT 178.950 88.950 181.050 89.400 ;
        RECT 250.950 88.950 253.050 89.400 ;
        RECT 271.950 88.950 274.050 89.400 ;
        RECT 364.950 90.600 367.050 91.050 ;
        RECT 376.950 90.600 379.050 91.050 ;
        RECT 382.950 90.600 385.050 91.050 ;
        RECT 364.950 89.400 385.050 90.600 ;
        RECT 364.950 88.950 367.050 89.400 ;
        RECT 376.950 88.950 379.050 89.400 ;
        RECT 382.950 88.950 385.050 89.400 ;
        RECT 451.950 90.600 454.050 91.050 ;
        RECT 472.950 90.600 475.050 91.050 ;
        RECT 451.950 89.400 475.050 90.600 ;
        RECT 451.950 88.950 454.050 89.400 ;
        RECT 472.950 88.950 475.050 89.400 ;
        RECT 520.950 90.600 523.050 91.050 ;
        RECT 538.950 90.600 541.050 91.050 ;
        RECT 520.950 89.400 541.050 90.600 ;
        RECT 520.950 88.950 523.050 89.400 ;
        RECT 538.950 88.950 541.050 89.400 ;
        RECT 598.950 90.600 601.050 91.050 ;
        RECT 712.950 90.600 715.050 91.050 ;
        RECT 598.950 89.400 715.050 90.600 ;
        RECT 598.950 88.950 601.050 89.400 ;
        RECT 712.950 88.950 715.050 89.400 ;
        RECT 727.950 90.600 730.050 91.050 ;
        RECT 787.950 90.600 790.050 91.050 ;
        RECT 727.950 89.400 790.050 90.600 ;
        RECT 727.950 88.950 730.050 89.400 ;
        RECT 787.950 88.950 790.050 89.400 ;
        RECT 805.950 90.600 808.050 91.050 ;
        RECT 823.950 90.600 826.050 91.050 ;
        RECT 805.950 89.400 826.050 90.600 ;
        RECT 805.950 88.950 808.050 89.400 ;
        RECT 823.950 88.950 826.050 89.400 ;
        RECT 190.950 87.600 193.050 88.050 ;
        RECT 247.950 87.600 250.050 88.050 ;
        RECT 190.950 86.400 250.050 87.600 ;
        RECT 190.950 85.950 193.050 86.400 ;
        RECT 247.950 85.950 250.050 86.400 ;
        RECT 256.950 87.600 259.050 88.050 ;
        RECT 268.950 87.600 271.050 88.050 ;
        RECT 256.950 86.400 271.050 87.600 ;
        RECT 256.950 85.950 259.050 86.400 ;
        RECT 268.950 85.950 271.050 86.400 ;
        RECT 277.950 87.600 280.050 88.050 ;
        RECT 358.950 87.600 361.050 88.050 ;
        RECT 277.950 86.400 361.050 87.600 ;
        RECT 277.950 85.950 280.050 86.400 ;
        RECT 358.950 85.950 361.050 86.400 ;
        RECT 529.950 87.600 532.050 88.050 ;
        RECT 544.950 87.600 547.050 88.050 ;
        RECT 529.950 86.400 547.050 87.600 ;
        RECT 529.950 85.950 532.050 86.400 ;
        RECT 544.950 85.950 547.050 86.400 ;
        RECT 595.950 87.600 598.050 88.050 ;
        RECT 715.950 87.600 718.050 88.050 ;
        RECT 733.950 87.600 736.050 88.050 ;
        RECT 856.950 87.600 859.050 88.050 ;
        RECT 595.950 86.400 859.050 87.600 ;
        RECT 595.950 85.950 598.050 86.400 ;
        RECT 715.950 85.950 718.050 86.400 ;
        RECT 733.950 85.950 736.050 86.400 ;
        RECT 856.950 85.950 859.050 86.400 ;
        RECT 61.950 84.600 64.050 85.050 ;
        RECT 157.950 84.600 160.050 85.050 ;
        RECT 223.800 84.600 225.900 85.050 ;
        RECT 61.950 83.400 225.900 84.600 ;
        RECT 61.950 82.950 64.050 83.400 ;
        RECT 157.950 82.950 160.050 83.400 ;
        RECT 223.800 82.950 225.900 83.400 ;
        RECT 319.950 84.600 322.050 85.050 ;
        RECT 355.950 84.600 358.050 85.050 ;
        RECT 319.950 83.400 358.050 84.600 ;
        RECT 319.950 82.950 322.050 83.400 ;
        RECT 355.950 82.950 358.050 83.400 ;
        RECT 364.950 84.600 367.050 85.050 ;
        RECT 454.950 84.600 457.050 85.050 ;
        RECT 364.950 83.400 457.050 84.600 ;
        RECT 364.950 82.950 367.050 83.400 ;
        RECT 454.950 82.950 457.050 83.400 ;
        RECT 532.950 84.600 535.050 85.050 ;
        RECT 637.950 84.600 640.050 85.050 ;
        RECT 655.950 84.600 658.050 85.050 ;
        RECT 532.950 83.400 658.050 84.600 ;
        RECT 532.950 82.950 535.050 83.400 ;
        RECT 637.950 82.950 640.050 83.400 ;
        RECT 655.950 82.950 658.050 83.400 ;
        RECT 673.950 84.600 676.050 85.050 ;
        RECT 685.950 84.600 688.050 85.050 ;
        RECT 673.950 83.400 688.050 84.600 ;
        RECT 673.950 82.950 676.050 83.400 ;
        RECT 685.950 82.950 688.050 83.400 ;
        RECT 736.950 84.600 739.050 85.050 ;
        RECT 793.950 84.600 796.050 85.050 ;
        RECT 736.950 83.400 796.050 84.600 ;
        RECT 736.950 82.950 739.050 83.400 ;
        RECT 793.950 82.950 796.050 83.400 ;
        RECT 166.950 81.600 169.050 82.050 ;
        RECT 259.950 81.600 262.050 82.050 ;
        RECT 166.950 80.400 262.050 81.600 ;
        RECT 166.950 79.950 169.050 80.400 ;
        RECT 259.950 79.950 262.050 80.400 ;
        RECT 373.950 81.600 376.050 82.050 ;
        RECT 382.950 81.600 385.050 82.050 ;
        RECT 373.950 80.400 385.050 81.600 ;
        RECT 373.950 79.950 376.050 80.400 ;
        RECT 382.950 79.950 385.050 80.400 ;
        RECT 691.950 81.600 694.050 82.050 ;
        RECT 742.950 81.600 745.050 82.050 ;
        RECT 691.950 80.400 745.050 81.600 ;
        RECT 691.950 79.950 694.050 80.400 ;
        RECT 742.950 79.950 745.050 80.400 ;
        RECT 199.950 78.600 202.050 79.050 ;
        RECT 292.950 78.600 295.050 79.050 ;
        RECT 199.950 77.400 295.050 78.600 ;
        RECT 199.950 76.950 202.050 77.400 ;
        RECT 292.950 76.950 295.050 77.400 ;
        RECT 358.950 78.600 361.050 79.050 ;
        RECT 436.950 78.600 439.050 79.050 ;
        RECT 358.950 77.400 439.050 78.600 ;
        RECT 358.950 76.950 361.050 77.400 ;
        RECT 436.950 76.950 439.050 77.400 ;
        RECT 484.950 78.600 487.050 79.050 ;
        RECT 514.950 78.600 517.050 79.050 ;
        RECT 484.950 77.400 517.050 78.600 ;
        RECT 484.950 76.950 487.050 77.400 ;
        RECT 514.950 76.950 517.050 77.400 ;
        RECT 643.950 78.600 646.050 79.050 ;
        RECT 781.950 78.600 784.050 79.050 ;
        RECT 643.950 77.400 784.050 78.600 ;
        RECT 643.950 76.950 646.050 77.400 ;
        RECT 781.950 76.950 784.050 77.400 ;
        RECT 37.950 75.600 40.050 76.050 ;
        RECT 61.950 75.600 64.050 76.050 ;
        RECT 76.950 75.600 79.050 76.050 ;
        RECT 37.950 74.400 79.050 75.600 ;
        RECT 37.950 73.950 40.050 74.400 ;
        RECT 61.950 73.950 64.050 74.400 ;
        RECT 76.950 73.950 79.050 74.400 ;
        RECT 151.950 75.600 154.050 76.050 ;
        RECT 238.950 75.600 241.050 76.050 ;
        RECT 151.950 74.400 241.050 75.600 ;
        RECT 151.950 73.950 154.050 74.400 ;
        RECT 238.950 73.950 241.050 74.400 ;
        RECT 250.950 75.600 253.050 76.050 ;
        RECT 283.950 75.600 286.050 76.050 ;
        RECT 250.950 74.400 286.050 75.600 ;
        RECT 250.950 73.950 253.050 74.400 ;
        RECT 283.950 73.950 286.050 74.400 ;
        RECT 322.950 75.600 325.050 76.050 ;
        RECT 352.950 75.600 355.050 76.050 ;
        RECT 322.950 74.400 355.050 75.600 ;
        RECT 322.950 73.950 325.050 74.400 ;
        RECT 352.950 73.950 355.050 74.400 ;
        RECT 367.950 75.600 370.050 76.050 ;
        RECT 406.950 75.600 409.050 76.050 ;
        RECT 442.950 75.600 445.050 76.050 ;
        RECT 367.950 74.400 445.050 75.600 ;
        RECT 367.950 73.950 370.050 74.400 ;
        RECT 406.950 73.950 409.050 74.400 ;
        RECT 442.950 73.950 445.050 74.400 ;
        RECT 481.950 75.600 484.050 76.050 ;
        RECT 568.950 75.600 571.050 76.050 ;
        RECT 481.950 74.400 571.050 75.600 ;
        RECT 481.950 73.950 484.050 74.400 ;
        RECT 568.950 73.950 571.050 74.400 ;
        RECT 22.950 72.600 25.050 73.050 ;
        RECT 28.950 72.600 31.050 73.050 ;
        RECT 115.950 72.600 118.050 73.050 ;
        RECT 22.950 71.400 118.050 72.600 ;
        RECT 22.950 70.950 25.050 71.400 ;
        RECT 28.950 70.950 31.050 71.400 ;
        RECT 115.950 70.950 118.050 71.400 ;
        RECT 127.950 72.600 130.050 73.050 ;
        RECT 241.950 72.600 244.050 73.050 ;
        RECT 316.950 72.600 319.050 73.050 ;
        RECT 127.950 71.400 147.600 72.600 ;
        RECT 127.950 70.950 130.050 71.400 ;
        RECT 146.400 70.050 147.600 71.400 ;
        RECT 241.950 71.400 319.050 72.600 ;
        RECT 241.950 70.950 244.050 71.400 ;
        RECT 316.950 70.950 319.050 71.400 ;
        RECT 328.950 72.600 331.050 73.050 ;
        RECT 346.950 72.600 349.050 73.050 ;
        RECT 328.950 71.400 349.050 72.600 ;
        RECT 328.950 70.950 331.050 71.400 ;
        RECT 346.950 70.950 349.050 71.400 ;
        RECT 355.950 72.600 358.050 73.050 ;
        RECT 373.950 72.600 376.050 73.050 ;
        RECT 379.950 72.600 382.050 73.050 ;
        RECT 355.950 71.400 382.050 72.600 ;
        RECT 355.950 70.950 358.050 71.400 ;
        RECT 373.950 70.950 376.050 71.400 ;
        RECT 379.950 70.950 382.050 71.400 ;
        RECT 487.950 72.600 490.050 73.050 ;
        RECT 613.950 72.600 616.050 73.050 ;
        RECT 487.950 71.400 616.050 72.600 ;
        RECT 487.950 70.950 490.050 71.400 ;
        RECT 613.950 70.950 616.050 71.400 ;
        RECT 619.950 72.600 622.050 73.050 ;
        RECT 682.950 72.600 685.050 73.050 ;
        RECT 619.950 71.400 685.050 72.600 ;
        RECT 619.950 70.950 622.050 71.400 ;
        RECT 682.950 70.950 685.050 71.400 ;
        RECT 145.950 69.600 148.050 70.050 ;
        RECT 178.950 69.600 181.050 70.050 ;
        RECT 145.950 68.400 181.050 69.600 ;
        RECT 145.950 67.950 148.050 68.400 ;
        RECT 178.950 67.950 181.050 68.400 ;
        RECT 271.950 69.600 274.050 70.050 ;
        RECT 301.950 69.600 304.050 70.050 ;
        RECT 271.950 68.400 304.050 69.600 ;
        RECT 271.950 67.950 274.050 68.400 ;
        RECT 301.950 67.950 304.050 68.400 ;
        RECT 334.950 69.600 337.050 70.050 ;
        RECT 349.950 69.600 352.050 70.050 ;
        RECT 445.950 69.600 448.050 70.050 ;
        RECT 334.950 68.400 448.050 69.600 ;
        RECT 334.950 67.950 337.050 68.400 ;
        RECT 349.950 67.950 352.050 68.400 ;
        RECT 445.950 67.950 448.050 68.400 ;
        RECT 784.950 69.600 787.050 70.050 ;
        RECT 841.950 69.600 844.050 70.050 ;
        RECT 844.950 69.600 847.050 70.050 ;
        RECT 784.950 68.400 847.050 69.600 ;
        RECT 784.950 67.950 787.050 68.400 ;
        RECT 841.950 67.950 844.050 68.400 ;
        RECT 844.950 67.950 847.050 68.400 ;
        RECT 31.950 66.600 34.050 67.050 ;
        RECT 49.950 66.600 52.050 67.050 ;
        RECT 31.950 65.400 52.050 66.600 ;
        RECT 31.950 64.950 34.050 65.400 ;
        RECT 49.950 64.950 52.050 65.400 ;
        RECT 115.950 66.600 118.050 67.050 ;
        RECT 142.950 66.600 145.050 67.050 ;
        RECT 115.950 65.400 145.050 66.600 ;
        RECT 115.950 64.950 118.050 65.400 ;
        RECT 142.950 64.950 145.050 65.400 ;
        RECT 169.950 66.600 172.050 67.050 ;
        RECT 190.950 66.600 193.050 67.050 ;
        RECT 169.950 65.400 193.050 66.600 ;
        RECT 169.950 64.950 172.050 65.400 ;
        RECT 190.950 64.950 193.050 65.400 ;
        RECT 238.950 66.600 241.050 67.050 ;
        RECT 277.950 66.600 280.050 67.050 ;
        RECT 238.950 65.400 280.050 66.600 ;
        RECT 238.950 64.950 241.050 65.400 ;
        RECT 277.950 64.950 280.050 65.400 ;
        RECT 358.950 66.600 361.050 67.050 ;
        RECT 367.950 66.600 370.050 67.050 ;
        RECT 358.950 65.400 370.050 66.600 ;
        RECT 358.950 64.950 361.050 65.400 ;
        RECT 367.950 64.950 370.050 65.400 ;
        RECT 379.950 66.600 382.050 67.050 ;
        RECT 385.950 66.600 388.050 67.050 ;
        RECT 394.950 66.600 397.050 67.050 ;
        RECT 379.950 65.400 397.050 66.600 ;
        RECT 379.950 64.950 382.050 65.400 ;
        RECT 385.950 64.950 388.050 65.400 ;
        RECT 394.950 64.950 397.050 65.400 ;
        RECT 457.950 66.600 460.050 67.050 ;
        RECT 481.950 66.600 484.050 67.050 ;
        RECT 457.950 65.400 484.050 66.600 ;
        RECT 457.950 64.950 460.050 65.400 ;
        RECT 481.950 64.950 484.050 65.400 ;
        RECT 595.950 66.600 598.050 67.050 ;
        RECT 607.950 66.600 610.050 67.050 ;
        RECT 595.950 65.400 610.050 66.600 ;
        RECT 595.950 64.950 598.050 65.400 ;
        RECT 607.950 64.950 610.050 65.400 ;
        RECT 616.950 66.600 619.050 67.050 ;
        RECT 643.950 66.600 646.050 67.050 ;
        RECT 652.950 66.600 655.050 67.050 ;
        RECT 616.950 65.400 655.050 66.600 ;
        RECT 616.950 64.950 619.050 65.400 ;
        RECT 643.950 64.950 646.050 65.400 ;
        RECT 652.950 64.950 655.050 65.400 ;
        RECT 694.950 66.600 697.050 67.050 ;
        RECT 706.950 66.600 709.050 67.050 ;
        RECT 721.950 66.600 724.050 67.050 ;
        RECT 694.950 65.400 724.050 66.600 ;
        RECT 694.950 64.950 697.050 65.400 ;
        RECT 706.950 64.950 709.050 65.400 ;
        RECT 721.950 64.950 724.050 65.400 ;
        RECT 796.950 66.600 799.050 67.050 ;
        RECT 832.950 66.600 835.050 67.050 ;
        RECT 796.950 65.400 835.050 66.600 ;
        RECT 796.950 64.950 799.050 65.400 ;
        RECT 832.950 64.950 835.050 65.400 ;
        RECT 79.950 63.600 82.050 64.050 ;
        RECT 94.950 63.600 97.050 64.050 ;
        RECT 100.950 63.600 103.050 64.050 ;
        RECT 79.950 62.400 103.050 63.600 ;
        RECT 79.950 61.950 82.050 62.400 ;
        RECT 94.950 61.950 97.050 62.400 ;
        RECT 100.950 61.950 103.050 62.400 ;
        RECT 127.950 61.950 130.050 64.050 ;
        RECT 163.950 63.600 166.050 64.050 ;
        RECT 199.950 63.600 202.050 64.050 ;
        RECT 205.950 63.600 208.050 64.050 ;
        RECT 232.950 63.600 235.050 64.050 ;
        RECT 163.950 62.400 235.050 63.600 ;
        RECT 163.950 61.950 166.050 62.400 ;
        RECT 199.950 61.950 202.050 62.400 ;
        RECT 205.950 61.950 208.050 62.400 ;
        RECT 232.950 61.950 235.050 62.400 ;
        RECT 352.950 61.950 355.050 64.050 ;
        RECT 415.950 63.600 418.050 64.050 ;
        RECT 442.950 63.600 445.050 64.050 ;
        RECT 415.950 62.400 445.050 63.600 ;
        RECT 415.950 61.950 418.050 62.400 ;
        RECT 442.950 61.950 445.050 62.400 ;
        RECT 454.950 61.950 457.050 64.050 ;
        RECT 472.950 63.600 475.050 64.050 ;
        RECT 478.950 63.600 481.050 64.050 ;
        RECT 487.950 63.600 490.050 64.050 ;
        RECT 472.950 62.400 490.050 63.600 ;
        RECT 472.950 61.950 475.050 62.400 ;
        RECT 478.950 61.950 481.050 62.400 ;
        RECT 487.950 61.950 490.050 62.400 ;
        RECT 493.950 63.600 496.050 64.050 ;
        RECT 535.950 63.600 538.050 64.050 ;
        RECT 493.950 62.400 538.050 63.600 ;
        RECT 493.950 61.950 496.050 62.400 ;
        RECT 535.950 61.950 538.050 62.400 ;
        RECT 784.950 61.950 787.050 64.050 ;
        RECT 847.950 61.950 850.050 64.050 ;
        RECT 862.950 63.600 865.050 64.050 ;
        RECT 871.950 63.600 874.050 64.050 ;
        RECT 862.950 62.400 874.050 63.600 ;
        RECT 862.950 61.950 865.050 62.400 ;
        RECT 871.950 61.950 874.050 62.400 ;
        RECT 16.950 59.100 19.050 61.200 ;
        RECT 4.950 54.600 7.050 55.050 ;
        RECT 13.950 54.600 16.050 54.900 ;
        RECT 4.950 53.400 16.050 54.600 ;
        RECT 4.950 52.950 7.050 53.400 ;
        RECT 13.950 52.800 16.050 53.400 ;
        RECT 17.400 52.050 18.600 59.100 ;
        RECT 25.950 58.950 28.050 61.050 ;
        RECT 43.950 59.100 46.050 61.200 ;
        RECT 67.950 60.750 70.050 61.200 ;
        RECT 73.950 60.750 76.050 61.200 ;
        RECT 67.950 59.550 76.050 60.750 ;
        RECT 67.950 59.100 70.050 59.550 ;
        RECT 73.950 59.100 76.050 59.550 ;
        RECT 85.950 59.100 88.050 61.200 ;
        RECT 106.950 59.100 109.050 61.200 ;
        RECT 26.400 54.600 27.600 58.950 ;
        RECT 34.950 54.600 37.050 54.900 ;
        RECT 44.400 54.600 45.600 59.100 ;
        RECT 86.400 57.600 87.600 59.100 ;
        RECT 107.400 57.600 108.600 59.100 ;
        RECT 86.400 56.400 108.600 57.600 ;
        RECT 26.400 53.400 37.050 54.600 ;
        RECT 38.400 54.000 45.600 54.600 ;
        RECT 34.950 52.800 37.050 53.400 ;
        RECT 37.950 53.400 45.600 54.000 ;
        RECT 49.950 54.600 52.050 55.050 ;
        RECT 58.950 54.600 61.050 54.900 ;
        RECT 49.950 53.400 61.050 54.600 ;
        RECT 107.400 54.600 108.600 56.400 ;
        RECT 112.950 54.600 115.050 55.050 ;
        RECT 128.400 54.900 129.600 61.950 ;
        RECT 130.800 59.100 132.900 61.200 ;
        RECT 133.950 60.600 136.050 61.050 ;
        RECT 151.950 60.600 154.050 61.200 ;
        RECT 174.000 60.600 178.050 61.050 ;
        RECT 133.950 59.400 154.050 60.600 ;
        RECT 107.400 53.400 115.050 54.600 ;
        RECT 16.950 49.950 19.050 52.050 ;
        RECT 37.950 49.950 40.050 53.400 ;
        RECT 49.950 52.950 52.050 53.400 ;
        RECT 58.950 52.800 61.050 53.400 ;
        RECT 112.950 52.950 115.050 53.400 ;
        RECT 127.950 52.800 130.050 54.900 ;
        RECT 131.400 54.600 132.600 59.100 ;
        RECT 133.950 58.950 136.050 59.400 ;
        RECT 151.950 59.100 154.050 59.400 ;
        RECT 148.950 54.600 151.050 54.900 ;
        RECT 131.400 53.400 151.050 54.600 ;
        RECT 148.950 52.800 151.050 53.400 ;
        RECT 46.950 51.600 49.050 52.050 ;
        RECT 82.950 51.600 85.050 52.050 ;
        RECT 46.950 50.400 85.050 51.600 ;
        RECT 46.950 49.950 49.050 50.400 ;
        RECT 82.950 49.950 85.050 50.400 ;
        RECT 88.950 51.600 91.050 52.050 ;
        RECT 152.400 51.600 153.600 59.100 ;
        RECT 173.400 58.950 178.050 60.600 ;
        RECT 202.950 58.950 205.050 61.050 ;
        RECT 211.950 60.600 214.050 61.200 ;
        RECT 220.950 60.600 223.050 61.050 ;
        RECT 226.950 60.600 229.050 61.200 ;
        RECT 211.950 59.400 229.050 60.600 ;
        RECT 211.950 59.100 214.050 59.400 ;
        RECT 220.950 58.950 223.050 59.400 ;
        RECT 226.950 59.100 229.050 59.400 ;
        RECT 256.950 60.600 259.050 61.200 ;
        RECT 271.950 60.600 274.050 61.200 ;
        RECT 289.950 60.600 292.050 61.200 ;
        RECT 256.950 59.400 270.600 60.600 ;
        RECT 256.950 59.100 259.050 59.400 ;
        RECT 173.400 54.900 174.600 58.950 ;
        RECT 172.950 54.600 175.050 54.900 ;
        RECT 193.950 54.600 196.050 54.900 ;
        RECT 172.950 53.400 196.050 54.600 ;
        RECT 203.400 54.600 204.600 58.950 ;
        RECT 269.400 57.600 270.600 59.400 ;
        RECT 271.950 59.400 292.050 60.600 ;
        RECT 271.950 59.100 274.050 59.400 ;
        RECT 289.950 59.100 292.050 59.400 ;
        RECT 310.950 60.600 313.050 61.200 ;
        RECT 328.950 60.600 331.050 61.200 ;
        RECT 310.950 59.400 331.050 60.600 ;
        RECT 310.950 59.100 313.050 59.400 ;
        RECT 328.950 59.100 331.050 59.400 ;
        RECT 343.950 60.750 346.050 61.200 ;
        RECT 349.950 60.750 352.050 61.200 ;
        RECT 343.950 59.550 352.050 60.750 ;
        RECT 343.950 59.100 346.050 59.550 ;
        RECT 349.950 59.100 352.050 59.550 ;
        RECT 215.400 56.400 270.600 57.600 ;
        RECT 215.400 54.900 216.600 56.400 ;
        RECT 269.400 54.900 270.600 56.400 ;
        RECT 353.400 54.900 354.600 61.950 ;
        RECT 382.950 58.950 385.050 61.050 ;
        RECT 400.950 60.600 403.050 61.200 ;
        RECT 421.950 60.600 424.050 61.200 ;
        RECT 400.950 59.400 424.050 60.600 ;
        RECT 400.950 59.100 403.050 59.400 ;
        RECT 208.950 54.600 211.050 54.900 ;
        RECT 203.400 53.400 211.050 54.600 ;
        RECT 172.950 52.800 175.050 53.400 ;
        RECT 193.950 52.800 196.050 53.400 ;
        RECT 208.950 52.800 211.050 53.400 ;
        RECT 214.950 52.800 217.050 54.900 ;
        RECT 268.950 52.800 271.050 54.900 ;
        RECT 277.950 54.450 280.050 54.900 ;
        RECT 286.950 54.450 289.050 54.900 ;
        RECT 277.950 53.250 289.050 54.450 ;
        RECT 277.950 52.800 280.050 53.250 ;
        RECT 286.950 52.800 289.050 53.250 ;
        RECT 313.950 54.450 316.050 54.900 ;
        RECT 322.800 54.450 324.900 54.900 ;
        RECT 313.950 53.250 324.900 54.450 ;
        RECT 313.950 52.800 316.050 53.250 ;
        RECT 322.800 52.800 324.900 53.250 ;
        RECT 352.950 52.800 355.050 54.900 ;
        RECT 383.400 54.600 384.600 58.950 ;
        RECT 410.400 55.050 411.600 59.400 ;
        RECT 421.950 59.100 424.050 59.400 ;
        RECT 427.950 60.750 430.050 61.200 ;
        RECT 436.950 60.750 439.050 61.200 ;
        RECT 427.950 59.550 439.050 60.750 ;
        RECT 427.950 59.100 430.050 59.550 ;
        RECT 436.950 59.100 439.050 59.550 ;
        RECT 442.950 59.100 445.050 61.200 ;
        RECT 388.950 54.600 391.050 55.050 ;
        RECT 383.400 53.400 391.050 54.600 ;
        RECT 388.950 52.950 391.050 53.400 ;
        RECT 409.950 52.950 412.050 55.050 ;
        RECT 443.400 54.600 444.600 59.100 ;
        RECT 451.800 54.600 453.900 55.050 ;
        RECT 455.400 54.900 456.600 61.950 ;
        RECT 463.950 60.600 466.050 61.200 ;
        RECT 469.950 60.600 472.050 61.050 ;
        RECT 463.950 59.400 472.050 60.600 ;
        RECT 463.950 59.100 466.050 59.400 ;
        RECT 469.950 58.950 472.050 59.400 ;
        RECT 502.950 60.600 505.050 61.200 ;
        RECT 520.950 60.600 523.050 61.200 ;
        RECT 502.950 59.400 523.050 60.600 ;
        RECT 502.950 59.100 505.050 59.400 ;
        RECT 520.950 59.100 523.050 59.400 ;
        RECT 541.950 59.100 544.050 61.200 ;
        RECT 547.950 60.750 550.050 61.200 ;
        RECT 556.950 60.750 559.050 61.200 ;
        RECT 547.950 59.550 559.050 60.750 ;
        RECT 547.950 59.100 550.050 59.550 ;
        RECT 556.950 59.100 559.050 59.550 ;
        RECT 562.950 60.600 565.050 61.200 ;
        RECT 568.950 60.600 571.050 61.050 ;
        RECT 562.950 59.400 571.050 60.600 ;
        RECT 562.950 59.100 565.050 59.400 ;
        RECT 542.400 55.050 543.600 59.100 ;
        RECT 568.950 58.950 571.050 59.400 ;
        RECT 577.950 60.600 580.050 61.200 ;
        RECT 586.950 60.600 589.050 61.050 ;
        RECT 577.950 59.400 589.050 60.600 ;
        RECT 577.950 59.100 580.050 59.400 ;
        RECT 586.950 58.950 589.050 59.400 ;
        RECT 601.950 59.100 604.050 61.200 ;
        RECT 622.950 59.100 625.050 61.200 ;
        RECT 637.950 59.100 640.050 61.200 ;
        RECT 655.950 60.600 658.050 61.050 ;
        RECT 688.950 60.600 691.050 61.200 ;
        RECT 706.950 60.600 709.050 61.200 ;
        RECT 655.950 59.400 663.600 60.600 ;
        RECT 443.400 53.400 453.900 54.600 ;
        RECT 451.800 52.950 453.900 53.400 ;
        RECT 454.950 52.800 457.050 54.900 ;
        RECT 460.950 54.450 463.050 54.900 ;
        RECT 472.950 54.450 475.050 54.900 ;
        RECT 460.950 53.250 475.050 54.450 ;
        RECT 460.950 52.800 463.050 53.250 ;
        RECT 472.950 52.800 475.050 53.250 ;
        RECT 484.950 54.600 487.050 54.900 ;
        RECT 517.950 54.600 520.050 54.900 ;
        RECT 484.950 53.400 520.050 54.600 ;
        RECT 484.950 52.800 487.050 53.400 ;
        RECT 517.950 52.800 520.050 53.400 ;
        RECT 529.950 54.600 532.050 55.050 ;
        RECT 538.950 54.600 541.050 54.900 ;
        RECT 529.950 53.400 541.050 54.600 ;
        RECT 542.400 53.400 547.050 55.050 ;
        RECT 529.950 52.950 532.050 53.400 ;
        RECT 538.950 52.800 541.050 53.400 ;
        RECT 543.000 52.950 547.050 53.400 ;
        RECT 568.950 54.450 571.050 54.900 ;
        RECT 574.950 54.450 577.050 54.900 ;
        RECT 568.950 53.250 577.050 54.450 ;
        RECT 568.950 52.800 571.050 53.250 ;
        RECT 574.950 52.800 577.050 53.250 ;
        RECT 586.950 54.450 589.050 54.900 ;
        RECT 592.950 54.450 595.050 54.900 ;
        RECT 586.950 53.250 595.050 54.450 ;
        RECT 602.400 54.600 603.600 59.100 ;
        RECT 623.400 57.600 624.600 59.100 ;
        RECT 638.400 57.600 639.600 59.100 ;
        RECT 655.950 58.950 658.050 59.400 ;
        RECT 623.400 56.400 639.600 57.600 ;
        RECT 634.950 54.600 637.050 54.900 ;
        RECT 602.400 53.400 637.050 54.600 ;
        RECT 638.400 54.600 639.600 56.400 ;
        RECT 646.950 54.600 649.050 55.050 ;
        RECT 662.400 54.900 663.600 59.400 ;
        RECT 688.950 59.400 709.050 60.600 ;
        RECT 688.950 59.100 691.050 59.400 ;
        RECT 706.950 59.100 709.050 59.400 ;
        RECT 712.950 60.750 715.050 61.200 ;
        RECT 727.950 60.750 730.050 61.200 ;
        RECT 712.950 59.550 730.050 60.750 ;
        RECT 712.950 59.100 715.050 59.550 ;
        RECT 727.950 59.100 730.050 59.550 ;
        RECT 733.950 60.750 736.050 61.200 ;
        RECT 757.950 60.750 760.050 61.200 ;
        RECT 733.950 59.550 760.050 60.750 ;
        RECT 733.950 59.100 736.050 59.550 ;
        RECT 757.950 59.100 760.050 59.550 ;
        RECT 763.950 60.750 766.050 61.200 ;
        RECT 769.950 60.750 772.050 61.200 ;
        RECT 763.950 59.550 772.050 60.750 ;
        RECT 763.950 59.100 766.050 59.550 ;
        RECT 769.950 59.100 772.050 59.550 ;
        RECT 707.400 57.600 708.600 59.100 ;
        RECT 707.400 56.400 780.600 57.600 ;
        RECT 638.400 53.400 649.050 54.600 ;
        RECT 586.950 52.800 589.050 53.250 ;
        RECT 592.950 52.800 595.050 53.250 ;
        RECT 634.950 52.800 637.050 53.400 ;
        RECT 646.950 52.950 649.050 53.400 ;
        RECT 661.950 52.800 664.050 54.900 ;
        RECT 676.950 54.450 679.050 54.900 ;
        RECT 685.950 54.600 688.050 54.900 ;
        RECT 703.950 54.600 706.050 54.900 ;
        RECT 685.950 54.450 706.050 54.600 ;
        RECT 676.950 53.400 706.050 54.450 ;
        RECT 707.400 54.600 708.600 56.400 ;
        RECT 724.950 54.600 727.050 54.900 ;
        RECT 707.400 53.400 727.050 54.600 ;
        RECT 676.950 53.250 688.050 53.400 ;
        RECT 676.950 52.800 679.050 53.250 ;
        RECT 685.950 52.800 688.050 53.250 ;
        RECT 703.950 52.800 706.050 53.400 ;
        RECT 724.950 52.800 727.050 53.400 ;
        RECT 733.950 54.600 736.050 55.050 ;
        RECT 779.400 54.900 780.600 56.400 ;
        RECT 785.400 54.900 786.600 61.950 ;
        RECT 787.950 60.600 790.050 61.200 ;
        RECT 787.950 59.400 792.600 60.600 ;
        RECT 787.950 59.100 790.050 59.400 ;
        RECT 791.400 55.050 792.600 59.400 ;
        RECT 796.950 58.950 799.050 61.050 ;
        RECT 802.950 59.100 805.050 61.200 ;
        RECT 808.950 59.100 811.050 61.200 ;
        RECT 826.950 59.100 829.050 61.200 ;
        RECT 797.400 55.050 798.600 58.950 ;
        RECT 739.950 54.600 742.050 54.900 ;
        RECT 733.950 53.400 742.050 54.600 ;
        RECT 733.950 52.950 736.050 53.400 ;
        RECT 739.950 52.800 742.050 53.400 ;
        RECT 748.950 54.450 751.050 54.900 ;
        RECT 760.950 54.450 763.050 54.900 ;
        RECT 748.950 53.250 763.050 54.450 ;
        RECT 748.950 52.800 751.050 53.250 ;
        RECT 760.950 52.800 763.050 53.250 ;
        RECT 778.950 52.800 781.050 54.900 ;
        RECT 784.950 52.800 787.050 54.900 ;
        RECT 790.950 52.950 793.050 55.050 ;
        RECT 796.950 52.950 799.050 55.050 ;
        RECT 803.400 54.600 804.600 59.100 ;
        RECT 809.400 57.600 810.600 59.100 ;
        RECT 809.400 56.400 816.600 57.600 ;
        RECT 815.400 55.050 816.600 56.400 ;
        RECT 811.950 54.600 814.050 55.050 ;
        RECT 803.400 53.400 814.050 54.600 ;
        RECT 815.400 53.400 820.050 55.050 ;
        RECT 827.400 54.600 828.600 59.100 ;
        RECT 848.400 54.900 849.600 61.950 ;
        RECT 850.950 59.100 853.050 61.200 ;
        RECT 841.950 54.600 844.050 54.900 ;
        RECT 827.400 53.400 844.050 54.600 ;
        RECT 811.950 52.950 814.050 53.400 ;
        RECT 816.000 52.950 820.050 53.400 ;
        RECT 841.950 52.800 844.050 53.400 ;
        RECT 847.950 52.800 850.050 54.900 ;
        RECT 187.950 51.600 190.050 52.050 ;
        RECT 88.950 50.400 111.600 51.600 ;
        RECT 152.400 50.400 190.050 51.600 ;
        RECT 88.950 49.950 91.050 50.400 ;
        RECT 110.400 49.050 111.600 50.400 ;
        RECT 187.950 49.950 190.050 50.400 ;
        RECT 295.950 51.600 298.050 52.050 ;
        RECT 307.950 51.600 310.050 52.050 ;
        RECT 295.950 50.400 310.050 51.600 ;
        RECT 323.400 51.600 324.600 52.800 ;
        RECT 331.950 51.600 334.050 52.050 ;
        RECT 370.950 51.600 373.050 52.050 ;
        RECT 391.950 51.600 394.050 52.050 ;
        RECT 323.400 50.400 334.050 51.600 ;
        RECT 295.950 49.950 298.050 50.400 ;
        RECT 307.950 49.950 310.050 50.400 ;
        RECT 331.950 49.950 334.050 50.400 ;
        RECT 344.400 50.400 369.600 51.600 ;
        RECT 344.400 49.050 345.600 50.400 ;
        RECT 31.950 48.600 34.050 49.050 ;
        RECT 40.950 48.600 43.050 49.050 ;
        RECT 31.950 47.400 43.050 48.600 ;
        RECT 31.950 46.950 34.050 47.400 ;
        RECT 40.950 46.950 43.050 47.400 ;
        RECT 52.950 48.600 55.050 49.050 ;
        RECT 61.950 48.600 64.050 49.050 ;
        RECT 52.950 47.400 64.050 48.600 ;
        RECT 52.950 46.950 55.050 47.400 ;
        RECT 61.950 46.950 64.050 47.400 ;
        RECT 91.950 48.600 94.050 49.050 ;
        RECT 103.950 48.600 106.050 49.050 ;
        RECT 91.950 47.400 106.050 48.600 ;
        RECT 91.950 46.950 94.050 47.400 ;
        RECT 103.950 46.950 106.050 47.400 ;
        RECT 109.950 48.600 112.050 49.050 ;
        RECT 142.950 48.600 145.050 49.050 ;
        RECT 109.950 47.400 145.050 48.600 ;
        RECT 109.950 46.950 112.050 47.400 ;
        RECT 142.950 46.950 145.050 47.400 ;
        RECT 175.950 48.600 178.050 49.050 ;
        RECT 211.950 48.600 214.050 49.050 ;
        RECT 175.950 47.400 214.050 48.600 ;
        RECT 175.950 46.950 178.050 47.400 ;
        RECT 211.950 46.950 214.050 47.400 ;
        RECT 223.950 48.600 226.050 49.050 ;
        RECT 241.950 48.600 244.050 49.050 ;
        RECT 247.950 48.600 250.050 49.050 ;
        RECT 223.950 47.400 250.050 48.600 ;
        RECT 223.950 46.950 226.050 47.400 ;
        RECT 241.950 46.950 244.050 47.400 ;
        RECT 247.950 46.950 250.050 47.400 ;
        RECT 253.950 48.600 256.050 49.050 ;
        RECT 343.950 48.600 346.050 49.050 ;
        RECT 253.950 47.400 346.050 48.600 ;
        RECT 253.950 46.950 256.050 47.400 ;
        RECT 343.950 46.950 346.050 47.400 ;
        RECT 358.950 48.600 361.050 49.050 ;
        RECT 364.950 48.600 367.050 49.050 ;
        RECT 358.950 47.400 367.050 48.600 ;
        RECT 368.400 48.600 369.600 50.400 ;
        RECT 370.950 50.400 394.050 51.600 ;
        RECT 473.400 51.600 474.600 52.800 ;
        RECT 851.400 52.050 852.600 59.100 ;
        RECT 499.950 51.600 502.050 52.050 ;
        RECT 473.400 50.400 502.050 51.600 ;
        RECT 370.950 49.950 373.050 50.400 ;
        RECT 391.950 49.950 394.050 50.400 ;
        RECT 499.950 49.950 502.050 50.400 ;
        RECT 673.950 51.600 676.050 52.050 ;
        RECT 766.950 51.600 769.050 52.050 ;
        RECT 673.950 50.400 769.050 51.600 ;
        RECT 673.950 49.950 676.050 50.400 ;
        RECT 766.950 49.950 769.050 50.400 ;
        RECT 793.950 51.600 796.050 52.050 ;
        RECT 799.950 51.600 802.050 52.050 ;
        RECT 793.950 50.400 802.050 51.600 ;
        RECT 793.950 49.950 796.050 50.400 ;
        RECT 799.950 49.950 802.050 50.400 ;
        RECT 850.950 49.950 853.050 52.050 ;
        RECT 418.950 48.600 421.050 49.050 ;
        RECT 427.950 48.600 430.050 49.050 ;
        RECT 368.400 47.400 430.050 48.600 ;
        RECT 358.950 46.950 361.050 47.400 ;
        RECT 364.950 46.950 367.050 47.400 ;
        RECT 418.950 46.950 421.050 47.400 ;
        RECT 427.950 46.950 430.050 47.400 ;
        RECT 475.950 48.600 478.050 49.050 ;
        RECT 484.950 48.600 487.050 49.050 ;
        RECT 475.950 47.400 487.050 48.600 ;
        RECT 475.950 46.950 478.050 47.400 ;
        RECT 484.950 46.950 487.050 47.400 ;
        RECT 619.950 48.600 622.050 49.050 ;
        RECT 640.950 48.600 643.050 49.050 ;
        RECT 652.950 48.600 655.050 49.050 ;
        RECT 679.950 48.600 682.050 49.050 ;
        RECT 619.950 47.400 682.050 48.600 ;
        RECT 619.950 46.950 622.050 47.400 ;
        RECT 640.950 46.950 643.050 47.400 ;
        RECT 652.950 46.950 655.050 47.400 ;
        RECT 679.950 46.950 682.050 47.400 ;
        RECT 751.950 48.600 754.050 49.050 ;
        RECT 775.950 48.600 778.050 49.050 ;
        RECT 751.950 47.400 778.050 48.600 ;
        RECT 751.950 46.950 754.050 47.400 ;
        RECT 775.950 46.950 778.050 47.400 ;
        RECT 823.950 48.600 826.050 49.050 ;
        RECT 835.950 48.600 838.050 49.050 ;
        RECT 823.950 47.400 838.050 48.600 ;
        RECT 823.950 46.950 826.050 47.400 ;
        RECT 835.950 46.950 838.050 47.400 ;
        RECT 865.950 48.600 868.050 49.050 ;
        RECT 874.950 48.600 877.050 49.050 ;
        RECT 865.950 47.400 877.050 48.600 ;
        RECT 865.950 46.950 868.050 47.400 ;
        RECT 874.950 46.950 877.050 47.400 ;
        RECT 16.950 45.600 19.050 46.050 ;
        RECT 46.950 45.600 49.050 46.050 ;
        RECT 16.950 44.400 49.050 45.600 ;
        RECT 16.950 43.950 19.050 44.400 ;
        RECT 46.950 43.950 49.050 44.400 ;
        RECT 64.950 45.600 67.050 46.050 ;
        RECT 70.950 45.600 73.050 46.050 ;
        RECT 88.950 45.600 91.050 46.050 ;
        RECT 121.950 45.600 124.050 46.050 ;
        RECT 64.950 44.400 124.050 45.600 ;
        RECT 64.950 43.950 67.050 44.400 ;
        RECT 70.950 43.950 73.050 44.400 ;
        RECT 88.950 43.950 91.050 44.400 ;
        RECT 121.950 43.950 124.050 44.400 ;
        RECT 148.950 45.600 151.050 46.050 ;
        RECT 214.950 45.600 217.050 46.050 ;
        RECT 148.950 44.400 217.050 45.600 ;
        RECT 148.950 43.950 151.050 44.400 ;
        RECT 214.950 43.950 217.050 44.400 ;
        RECT 268.950 45.600 271.050 46.050 ;
        RECT 274.950 45.600 277.050 46.050 ;
        RECT 268.950 44.400 277.050 45.600 ;
        RECT 268.950 43.950 271.050 44.400 ;
        RECT 274.950 43.950 277.050 44.400 ;
        RECT 301.950 45.600 304.050 46.050 ;
        RECT 319.950 45.600 322.050 46.050 ;
        RECT 301.950 44.400 322.050 45.600 ;
        RECT 301.950 43.950 304.050 44.400 ;
        RECT 319.950 43.950 322.050 44.400 ;
        RECT 346.950 45.600 349.050 46.050 ;
        RECT 370.950 45.600 373.050 46.050 ;
        RECT 346.950 44.400 373.050 45.600 ;
        RECT 346.950 43.950 349.050 44.400 ;
        RECT 370.950 43.950 373.050 44.400 ;
        RECT 379.950 45.600 382.050 46.050 ;
        RECT 385.950 45.600 388.050 46.050 ;
        RECT 379.950 44.400 388.050 45.600 ;
        RECT 379.950 43.950 382.050 44.400 ;
        RECT 385.950 43.950 388.050 44.400 ;
        RECT 409.950 45.600 412.050 46.050 ;
        RECT 439.950 45.600 442.050 46.050 ;
        RECT 409.950 44.400 442.050 45.600 ;
        RECT 409.950 43.950 412.050 44.400 ;
        RECT 439.950 43.950 442.050 44.400 ;
        RECT 667.950 45.600 670.050 46.050 ;
        RECT 676.950 45.600 679.050 46.050 ;
        RECT 667.950 44.400 679.050 45.600 ;
        RECT 667.950 43.950 670.050 44.400 ;
        RECT 676.950 43.950 679.050 44.400 ;
        RECT 703.950 45.600 706.050 46.050 ;
        RECT 718.950 45.600 721.050 46.050 ;
        RECT 703.950 44.400 721.050 45.600 ;
        RECT 776.400 45.600 777.600 46.950 ;
        RECT 838.950 45.600 841.050 46.050 ;
        RECT 776.400 44.400 841.050 45.600 ;
        RECT 703.950 43.950 706.050 44.400 ;
        RECT 718.950 43.950 721.050 44.400 ;
        RECT 838.950 43.950 841.050 44.400 ;
        RECT 67.950 42.600 70.050 43.050 ;
        RECT 85.950 42.600 88.050 43.050 ;
        RECT 67.950 41.400 88.050 42.600 ;
        RECT 67.950 40.950 70.050 41.400 ;
        RECT 85.950 40.950 88.050 41.400 ;
        RECT 157.950 42.600 160.050 43.050 ;
        RECT 196.950 42.600 199.050 43.050 ;
        RECT 157.950 41.400 199.050 42.600 ;
        RECT 157.950 40.950 160.050 41.400 ;
        RECT 196.950 40.950 199.050 41.400 ;
        RECT 211.950 42.600 214.050 43.050 ;
        RECT 223.950 42.600 226.050 43.050 ;
        RECT 211.950 41.400 226.050 42.600 ;
        RECT 320.400 42.600 321.600 43.950 ;
        RECT 343.950 42.600 346.050 43.050 ;
        RECT 320.400 41.400 346.050 42.600 ;
        RECT 211.950 40.950 214.050 41.400 ;
        RECT 223.950 40.950 226.050 41.400 ;
        RECT 343.950 40.950 346.050 41.400 ;
        RECT 376.950 42.600 379.050 43.050 ;
        RECT 391.950 42.600 394.050 43.050 ;
        RECT 400.950 42.600 403.050 43.050 ;
        RECT 376.950 41.400 403.050 42.600 ;
        RECT 376.950 40.950 379.050 41.400 ;
        RECT 391.950 40.950 394.050 41.400 ;
        RECT 400.950 40.950 403.050 41.400 ;
        RECT 478.950 42.600 481.050 43.050 ;
        RECT 493.950 42.600 496.050 43.050 ;
        RECT 478.950 41.400 496.050 42.600 ;
        RECT 478.950 40.950 481.050 41.400 ;
        RECT 493.950 40.950 496.050 41.400 ;
        RECT 646.950 42.600 649.050 43.050 ;
        RECT 745.950 42.600 748.050 43.050 ;
        RECT 646.950 41.400 748.050 42.600 ;
        RECT 646.950 40.950 649.050 41.400 ;
        RECT 745.950 40.950 748.050 41.400 ;
        RECT 817.950 42.600 820.050 43.050 ;
        RECT 835.950 42.600 838.050 43.050 ;
        RECT 817.950 41.400 838.050 42.600 ;
        RECT 817.950 40.950 820.050 41.400 ;
        RECT 835.950 40.950 838.050 41.400 ;
        RECT 13.950 39.600 16.050 40.050 ;
        RECT 19.950 39.600 22.050 40.050 ;
        RECT 64.950 39.600 67.050 40.050 ;
        RECT 13.950 38.400 67.050 39.600 ;
        RECT 13.950 37.950 16.050 38.400 ;
        RECT 19.950 37.950 22.050 38.400 ;
        RECT 64.950 37.950 67.050 38.400 ;
        RECT 133.950 39.600 136.050 40.050 ;
        RECT 154.950 39.600 157.050 40.050 ;
        RECT 133.950 38.400 157.050 39.600 ;
        RECT 133.950 37.950 136.050 38.400 ;
        RECT 154.950 37.950 157.050 38.400 ;
        RECT 172.950 39.600 175.050 40.050 ;
        RECT 199.800 39.600 201.900 40.050 ;
        RECT 172.950 38.400 201.900 39.600 ;
        RECT 172.950 37.950 175.050 38.400 ;
        RECT 199.800 37.950 201.900 38.400 ;
        RECT 202.950 39.600 205.050 40.050 ;
        RECT 208.950 39.600 211.050 40.050 ;
        RECT 229.950 39.600 232.050 40.050 ;
        RECT 202.950 38.400 232.050 39.600 ;
        RECT 202.950 37.950 205.050 38.400 ;
        RECT 208.950 37.950 211.050 38.400 ;
        RECT 229.950 37.950 232.050 38.400 ;
        RECT 292.950 39.600 295.050 40.050 ;
        RECT 373.950 39.600 376.050 40.050 ;
        RECT 292.950 38.400 376.050 39.600 ;
        RECT 292.950 37.950 295.050 38.400 ;
        RECT 373.950 37.950 376.050 38.400 ;
        RECT 394.950 39.600 397.050 40.050 ;
        RECT 451.950 39.600 454.050 40.050 ;
        RECT 475.950 39.600 478.050 40.050 ;
        RECT 394.950 38.400 478.050 39.600 ;
        RECT 394.950 37.950 397.050 38.400 ;
        RECT 451.950 37.950 454.050 38.400 ;
        RECT 475.950 37.950 478.050 38.400 ;
        RECT 496.950 39.600 499.050 40.050 ;
        RECT 508.950 39.600 511.050 40.050 ;
        RECT 532.950 39.600 535.050 40.050 ;
        RECT 496.950 38.400 535.050 39.600 ;
        RECT 496.950 37.950 499.050 38.400 ;
        RECT 508.950 37.950 511.050 38.400 ;
        RECT 532.950 37.950 535.050 38.400 ;
        RECT 559.950 39.600 562.050 40.050 ;
        RECT 583.950 39.600 586.050 40.050 ;
        RECT 634.950 39.600 637.050 40.050 ;
        RECT 559.950 38.400 637.050 39.600 ;
        RECT 559.950 37.950 562.050 38.400 ;
        RECT 583.950 37.950 586.050 38.400 ;
        RECT 634.950 37.950 637.050 38.400 ;
        RECT 655.950 39.600 658.050 40.050 ;
        RECT 664.950 39.600 667.050 40.050 ;
        RECT 655.950 38.400 667.050 39.600 ;
        RECT 655.950 37.950 658.050 38.400 ;
        RECT 664.950 37.950 667.050 38.400 ;
        RECT 700.950 39.600 703.050 40.050 ;
        RECT 709.950 39.600 712.050 40.050 ;
        RECT 700.950 38.400 712.050 39.600 ;
        RECT 700.950 37.950 703.050 38.400 ;
        RECT 709.950 37.950 712.050 38.400 ;
        RECT 715.950 39.600 718.050 40.050 ;
        RECT 730.950 39.600 733.050 40.050 ;
        RECT 715.950 38.400 733.050 39.600 ;
        RECT 715.950 37.950 718.050 38.400 ;
        RECT 730.950 37.950 733.050 38.400 ;
        RECT 805.950 39.600 808.050 40.050 ;
        RECT 826.950 39.600 829.050 40.050 ;
        RECT 805.950 38.400 829.050 39.600 ;
        RECT 805.950 37.950 808.050 38.400 ;
        RECT 826.950 37.950 829.050 38.400 ;
        RECT 112.950 36.600 115.050 37.050 ;
        RECT 127.950 36.600 130.050 37.050 ;
        RECT 217.950 36.600 220.050 37.050 ;
        RECT 244.950 36.600 247.050 37.050 ;
        RECT 112.950 35.400 130.050 36.600 ;
        RECT 112.950 34.950 115.050 35.400 ;
        RECT 127.950 34.950 130.050 35.400 ;
        RECT 131.400 35.400 220.050 36.600 ;
        RECT 64.950 33.600 67.050 34.050 ;
        RECT 103.950 33.600 106.050 34.050 ;
        RECT 64.950 32.400 106.050 33.600 ;
        RECT 64.950 31.950 67.050 32.400 ;
        RECT 103.950 31.950 106.050 32.400 ;
        RECT 109.950 33.600 112.050 34.050 ;
        RECT 131.400 33.600 132.600 35.400 ;
        RECT 217.950 34.950 220.050 35.400 ;
        RECT 239.400 35.400 247.050 36.600 ;
        RECT 109.950 32.400 132.600 33.600 ;
        RECT 154.950 33.600 157.050 34.050 ;
        RECT 184.950 33.600 187.050 34.050 ;
        RECT 154.950 32.400 187.050 33.600 ;
        RECT 109.950 31.950 112.050 32.400 ;
        RECT 154.950 31.950 157.050 32.400 ;
        RECT 184.950 31.950 187.050 32.400 ;
        RECT 199.950 33.600 202.050 34.050 ;
        RECT 214.950 33.600 217.050 34.050 ;
        RECT 228.000 33.600 232.050 34.050 ;
        RECT 239.400 33.600 240.600 35.400 ;
        RECT 244.950 34.950 247.050 35.400 ;
        RECT 307.950 36.600 310.050 37.050 ;
        RECT 355.950 36.600 358.050 37.050 ;
        RECT 370.950 36.600 373.050 37.050 ;
        RECT 307.950 35.400 336.600 36.600 ;
        RECT 307.950 34.950 310.050 35.400 ;
        RECT 199.950 32.400 217.050 33.600 ;
        RECT 199.950 31.950 202.050 32.400 ;
        RECT 214.950 31.950 217.050 32.400 ;
        RECT 227.400 32.400 240.600 33.600 ;
        RECT 301.950 33.600 304.050 34.050 ;
        RECT 328.950 33.600 331.050 34.050 ;
        RECT 301.950 32.400 331.050 33.600 ;
        RECT 335.400 33.600 336.600 35.400 ;
        RECT 355.950 35.400 373.050 36.600 ;
        RECT 355.950 34.950 358.050 35.400 ;
        RECT 370.950 34.950 373.050 35.400 ;
        RECT 382.950 36.600 385.050 37.050 ;
        RECT 412.950 36.600 415.050 37.050 ;
        RECT 382.950 35.400 415.050 36.600 ;
        RECT 382.950 34.950 385.050 35.400 ;
        RECT 412.950 34.950 415.050 35.400 ;
        RECT 439.950 36.600 442.050 37.050 ;
        RECT 487.950 36.600 490.050 37.050 ;
        RECT 439.950 35.400 490.050 36.600 ;
        RECT 439.950 34.950 442.050 35.400 ;
        RECT 487.950 34.950 490.050 35.400 ;
        RECT 523.950 36.600 526.050 37.050 ;
        RECT 643.950 36.600 646.050 37.050 ;
        RECT 676.950 36.600 679.050 37.050 ;
        RECT 523.950 35.400 679.050 36.600 ;
        RECT 523.950 34.950 526.050 35.400 ;
        RECT 643.950 34.950 646.050 35.400 ;
        RECT 676.950 34.950 679.050 35.400 ;
        RECT 718.950 36.600 721.050 37.050 ;
        RECT 757.950 36.600 760.050 37.050 ;
        RECT 718.950 35.400 760.050 36.600 ;
        RECT 718.950 34.950 721.050 35.400 ;
        RECT 757.950 34.950 760.050 35.400 ;
        RECT 769.950 36.600 772.050 37.050 ;
        RECT 811.950 36.600 814.050 37.050 ;
        RECT 829.950 36.600 832.050 37.050 ;
        RECT 853.950 36.600 856.050 37.050 ;
        RECT 769.950 35.400 801.600 36.600 ;
        RECT 769.950 34.950 772.050 35.400 ;
        RECT 376.950 33.600 379.050 34.050 ;
        RECT 335.400 32.400 379.050 33.600 ;
        RECT 227.400 31.950 232.050 32.400 ;
        RECT 301.950 31.950 304.050 32.400 ;
        RECT 328.950 31.950 331.050 32.400 ;
        RECT 376.950 31.950 379.050 32.400 ;
        RECT 433.950 33.600 436.050 34.050 ;
        RECT 445.950 33.600 448.050 34.050 ;
        RECT 433.950 32.400 448.050 33.600 ;
        RECT 433.950 31.950 436.050 32.400 ;
        RECT 445.950 31.950 448.050 32.400 ;
        RECT 538.950 33.600 541.050 34.050 ;
        RECT 553.950 33.600 556.050 34.050 ;
        RECT 538.950 32.400 556.050 33.600 ;
        RECT 538.950 31.950 541.050 32.400 ;
        RECT 553.950 31.950 556.050 32.400 ;
        RECT 649.950 33.600 652.050 34.050 ;
        RECT 703.950 33.600 706.050 34.050 ;
        RECT 649.950 32.400 706.050 33.600 ;
        RECT 649.950 31.950 652.050 32.400 ;
        RECT 703.950 31.950 706.050 32.400 ;
        RECT 709.950 33.600 712.050 34.050 ;
        RECT 760.950 33.600 763.050 34.050 ;
        RECT 709.950 32.400 763.050 33.600 ;
        RECT 800.400 33.600 801.600 35.400 ;
        RECT 811.950 35.400 856.050 36.600 ;
        RECT 811.950 34.950 814.050 35.400 ;
        RECT 829.950 34.950 832.050 35.400 ;
        RECT 853.950 34.950 856.050 35.400 ;
        RECT 820.950 33.600 823.050 34.050 ;
        RECT 800.400 32.400 823.050 33.600 ;
        RECT 709.950 31.950 712.050 32.400 ;
        RECT 760.950 31.950 763.050 32.400 ;
        RECT 820.950 31.950 823.050 32.400 ;
        RECT 73.950 30.600 76.050 31.050 ;
        RECT 93.000 30.600 97.050 31.050 ;
        RECT 73.950 29.400 84.600 30.600 ;
        RECT 73.950 28.950 76.050 29.400 ;
        RECT 52.950 27.600 55.050 28.200 ;
        RECT 79.950 27.600 82.050 28.050 ;
        RECT 52.950 26.400 82.050 27.600 ;
        RECT 52.950 26.100 55.050 26.400 ;
        RECT 79.950 25.950 82.050 26.400 ;
        RECT 31.950 21.600 34.050 21.900 ;
        RECT 37.950 21.600 40.050 22.050 ;
        RECT 43.950 21.600 46.050 21.900 ;
        RECT 31.950 20.400 46.050 21.600 ;
        RECT 83.400 21.600 84.600 29.400 ;
        RECT 92.400 28.950 97.050 30.600 ;
        RECT 121.950 30.600 124.050 31.050 ;
        RECT 148.950 30.600 151.050 31.050 ;
        RECT 121.950 29.400 151.050 30.600 ;
        RECT 121.950 28.950 124.050 29.400 ;
        RECT 148.950 28.950 151.050 29.400 ;
        RECT 190.950 30.600 193.050 31.050 ;
        RECT 220.950 30.600 223.050 31.050 ;
        RECT 190.950 29.400 223.050 30.600 ;
        RECT 190.950 28.950 193.050 29.400 ;
        RECT 220.950 28.950 223.050 29.400 ;
        RECT 92.400 21.900 93.600 28.950 ;
        RECT 103.950 27.600 108.000 28.050 ;
        RECT 163.950 27.600 166.050 28.050 ;
        RECT 175.950 27.600 178.050 28.050 ;
        RECT 202.950 27.600 205.050 28.050 ;
        RECT 103.950 25.950 108.600 27.600 ;
        RECT 163.950 26.400 178.050 27.600 ;
        RECT 163.950 25.950 166.050 26.400 ;
        RECT 175.950 25.950 178.050 26.400 ;
        RECT 194.400 26.400 205.050 27.600 ;
        RECT 107.400 21.900 108.600 25.950 ;
        RECT 85.950 21.600 88.050 21.900 ;
        RECT 83.400 20.400 88.050 21.600 ;
        RECT 31.950 19.800 34.050 20.400 ;
        RECT 37.950 19.950 40.050 20.400 ;
        RECT 43.950 19.800 46.050 20.400 ;
        RECT 85.950 19.800 88.050 20.400 ;
        RECT 91.950 19.800 94.050 21.900 ;
        RECT 106.950 19.800 109.050 21.900 ;
        RECT 130.950 21.600 133.050 21.900 ;
        RECT 157.950 21.600 160.050 21.900 ;
        RECT 130.950 21.450 160.050 21.600 ;
        RECT 163.950 21.450 166.050 21.900 ;
        RECT 130.950 20.400 166.050 21.450 ;
        RECT 130.950 19.800 133.050 20.400 ;
        RECT 157.950 20.250 166.050 20.400 ;
        RECT 157.950 19.800 160.050 20.250 ;
        RECT 163.950 19.800 166.050 20.250 ;
        RECT 172.950 21.600 175.050 21.900 ;
        RECT 178.950 21.600 181.050 22.050 ;
        RECT 194.400 21.900 195.600 26.400 ;
        RECT 202.950 25.950 205.050 26.400 ;
        RECT 211.950 27.600 214.050 28.200 ;
        RECT 227.400 27.600 228.600 31.950 ;
        RECT 241.950 30.600 244.050 31.050 ;
        RECT 277.950 30.600 280.050 31.050 ;
        RECT 241.950 29.400 280.050 30.600 ;
        RECT 241.950 28.950 244.050 29.400 ;
        RECT 277.950 28.950 280.050 29.400 ;
        RECT 331.950 30.600 334.050 31.050 ;
        RECT 337.800 30.600 339.900 31.050 ;
        RECT 331.950 29.400 339.900 30.600 ;
        RECT 331.950 28.950 334.050 29.400 ;
        RECT 337.800 28.950 339.900 29.400 ;
        RECT 340.950 28.950 343.050 31.050 ;
        RECT 421.950 30.600 424.050 31.050 ;
        RECT 592.950 30.600 595.050 31.050 ;
        RECT 421.950 29.400 444.600 30.600 ;
        RECT 421.950 28.950 424.050 29.400 ;
        RECT 211.950 26.400 228.600 27.600 ;
        RECT 247.950 27.750 250.050 28.200 ;
        RECT 253.950 27.750 256.050 28.200 ;
        RECT 247.950 26.550 256.050 27.750 ;
        RECT 211.950 26.100 214.050 26.400 ;
        RECT 247.950 26.100 250.050 26.550 ;
        RECT 253.950 26.100 256.050 26.550 ;
        RECT 286.950 27.600 289.050 28.050 ;
        RECT 295.950 27.600 298.050 28.200 ;
        RECT 313.950 27.600 316.050 28.200 ;
        RECT 286.950 26.400 298.050 27.600 ;
        RECT 286.950 25.950 289.050 26.400 ;
        RECT 295.950 26.100 298.050 26.400 ;
        RECT 311.400 26.400 316.050 27.600 ;
        RECT 268.950 24.600 271.050 25.050 ;
        RECT 311.400 24.600 312.600 26.400 ;
        RECT 313.950 26.100 316.050 26.400 ;
        RECT 263.400 23.400 312.600 24.600 ;
        RECT 187.950 21.600 190.050 21.900 ;
        RECT 172.950 20.400 190.050 21.600 ;
        RECT 172.950 19.800 175.050 20.400 ;
        RECT 178.950 19.950 181.050 20.400 ;
        RECT 187.950 19.800 190.050 20.400 ;
        RECT 193.950 19.800 196.050 21.900 ;
        RECT 199.950 21.600 202.050 22.050 ;
        RECT 263.400 21.900 264.600 23.400 ;
        RECT 268.950 22.950 271.050 23.400 ;
        RECT 341.400 21.900 342.600 28.950 ;
        RECT 343.950 27.600 346.050 28.200 ;
        RECT 355.950 27.600 358.050 28.200 ;
        RECT 343.950 26.400 358.050 27.600 ;
        RECT 343.950 26.100 346.050 26.400 ;
        RECT 355.950 26.100 358.050 26.400 ;
        RECT 361.950 27.600 364.050 28.200 ;
        RECT 382.950 27.600 385.050 28.200 ;
        RECT 361.950 26.400 385.050 27.600 ;
        RECT 361.950 26.100 364.050 26.400 ;
        RECT 382.950 26.100 385.050 26.400 ;
        RECT 388.950 25.950 391.050 28.050 ;
        RECT 412.950 27.750 415.050 28.050 ;
        RECT 421.950 27.750 424.050 28.200 ;
        RECT 412.950 26.550 424.050 27.750 ;
        RECT 412.950 25.950 415.050 26.550 ;
        RECT 421.950 26.100 424.050 26.550 ;
        RECT 430.950 27.600 433.050 28.050 ;
        RECT 430.950 26.400 438.600 27.600 ;
        RECT 430.950 25.950 433.050 26.400 ;
        RECT 208.950 21.600 211.050 21.900 ;
        RECT 199.950 20.400 211.050 21.600 ;
        RECT 199.950 19.950 202.050 20.400 ;
        RECT 208.950 19.800 211.050 20.400 ;
        RECT 241.950 21.450 244.050 21.900 ;
        RECT 256.950 21.450 259.050 21.900 ;
        RECT 241.950 20.250 259.050 21.450 ;
        RECT 241.950 19.800 244.050 20.250 ;
        RECT 256.950 19.800 259.050 20.250 ;
        RECT 262.950 19.800 265.050 21.900 ;
        RECT 280.950 21.450 283.050 21.900 ;
        RECT 286.950 21.450 289.050 21.900 ;
        RECT 280.950 20.250 289.050 21.450 ;
        RECT 280.950 19.800 283.050 20.250 ;
        RECT 286.950 19.800 289.050 20.250 ;
        RECT 292.950 21.450 295.050 21.900 ;
        RECT 307.950 21.450 310.050 21.900 ;
        RECT 292.950 20.250 310.050 21.450 ;
        RECT 292.950 19.800 295.050 20.250 ;
        RECT 307.950 19.800 310.050 20.250 ;
        RECT 322.950 21.450 325.050 21.900 ;
        RECT 328.950 21.450 331.050 21.900 ;
        RECT 322.950 20.250 331.050 21.450 ;
        RECT 322.950 19.800 325.050 20.250 ;
        RECT 328.950 19.800 331.050 20.250 ;
        RECT 340.950 19.800 343.050 21.900 ;
        RECT 364.950 21.600 367.050 21.900 ;
        RECT 379.950 21.600 382.050 21.900 ;
        RECT 364.950 20.400 382.050 21.600 ;
        RECT 364.950 19.800 367.050 20.400 ;
        RECT 379.950 19.800 382.050 20.400 ;
        RECT 385.950 21.600 388.050 21.900 ;
        RECT 389.400 21.600 390.600 25.950 ;
        RECT 437.400 21.900 438.600 26.400 ;
        RECT 443.400 21.900 444.600 29.400 ;
        RECT 592.950 29.400 630.600 30.600 ;
        RECT 592.950 28.950 595.050 29.400 ;
        RECT 457.950 27.750 460.050 28.200 ;
        RECT 487.950 27.750 490.050 28.200 ;
        RECT 457.950 26.550 490.050 27.750 ;
        RECT 457.950 26.100 460.050 26.550 ;
        RECT 487.950 26.100 490.050 26.550 ;
        RECT 526.950 27.600 529.050 28.050 ;
        RECT 544.950 27.600 547.050 28.050 ;
        RECT 559.950 27.600 562.050 28.200 ;
        RECT 526.950 26.400 562.050 27.600 ;
        RECT 526.950 25.950 529.050 26.400 ;
        RECT 544.950 25.950 547.050 26.400 ;
        RECT 559.950 26.100 562.050 26.400 ;
        RECT 565.950 27.600 568.050 28.200 ;
        RECT 577.950 27.600 580.050 28.200 ;
        RECT 598.950 27.600 601.050 28.200 ;
        RECT 565.950 26.400 580.050 27.600 ;
        RECT 565.950 26.100 568.050 26.400 ;
        RECT 577.950 26.100 580.050 26.400 ;
        RECT 581.400 26.400 601.050 27.600 ;
        RECT 581.400 24.600 582.600 26.400 ;
        RECT 598.950 26.100 601.050 26.400 ;
        RECT 482.400 23.400 510.600 24.600 ;
        RECT 482.400 21.900 483.600 23.400 ;
        RECT 397.950 21.600 400.050 21.900 ;
        RECT 385.950 20.400 400.050 21.600 ;
        RECT 385.950 19.800 388.050 20.400 ;
        RECT 397.950 19.800 400.050 20.400 ;
        RECT 436.950 19.800 439.050 21.900 ;
        RECT 442.950 19.800 445.050 21.900 ;
        RECT 481.950 19.800 484.050 21.900 ;
        RECT 487.950 21.600 490.050 22.050 ;
        RECT 509.400 21.900 510.600 23.400 ;
        RECT 563.400 23.400 582.600 24.600 ;
        RECT 563.400 21.900 564.600 23.400 ;
        RECT 602.400 21.900 603.600 29.400 ;
        RECT 604.950 27.750 607.050 28.200 ;
        RECT 613.950 27.750 616.050 28.200 ;
        RECT 604.950 27.600 616.050 27.750 ;
        RECT 625.950 27.600 628.050 28.200 ;
        RECT 604.950 26.550 628.050 27.600 ;
        RECT 604.950 26.100 607.050 26.550 ;
        RECT 613.950 26.400 628.050 26.550 ;
        RECT 613.950 26.100 616.050 26.400 ;
        RECT 625.950 26.100 628.050 26.400 ;
        RECT 629.400 21.900 630.600 29.400 ;
        RECT 643.950 28.950 646.050 31.050 ;
        RECT 670.950 30.600 673.050 31.050 ;
        RECT 691.950 30.600 694.050 31.050 ;
        RECT 670.950 29.400 694.050 30.600 ;
        RECT 670.950 28.950 673.050 29.400 ;
        RECT 691.950 28.950 694.050 29.400 ;
        RECT 772.950 30.600 775.050 31.050 ;
        RECT 796.950 30.600 799.050 30.900 ;
        RECT 772.950 29.400 799.050 30.600 ;
        RECT 772.950 28.950 775.050 29.400 ;
        RECT 634.950 27.600 637.050 28.050 ;
        RECT 640.950 27.600 643.050 28.200 ;
        RECT 634.950 26.400 643.050 27.600 ;
        RECT 634.950 25.950 637.050 26.400 ;
        RECT 640.950 26.100 643.050 26.400 ;
        RECT 644.400 21.900 645.600 28.950 ;
        RECT 796.950 28.800 799.050 29.400 ;
        RECT 838.950 28.950 841.050 31.050 ;
        RECT 850.950 28.950 853.050 31.050 ;
        RECT 856.950 30.600 859.050 31.050 ;
        RECT 865.950 30.600 868.050 31.050 ;
        RECT 856.950 29.400 868.050 30.600 ;
        RECT 856.950 28.950 859.050 29.400 ;
        RECT 865.950 28.950 868.050 29.400 ;
        RECT 651.000 27.600 655.050 28.050 ;
        RECT 650.400 25.950 655.050 27.600 ;
        RECT 650.400 21.900 651.600 25.950 ;
        RECT 658.950 24.600 661.050 28.050 ;
        RECT 685.950 27.600 688.050 28.200 ;
        RECT 674.250 26.400 688.050 27.600 ;
        RECT 658.950 24.000 663.600 24.600 ;
        RECT 659.400 23.400 663.600 24.000 ;
        RECT 662.400 21.900 663.600 23.400 ;
        RECT 674.250 22.050 675.450 26.400 ;
        RECT 685.950 26.100 688.050 26.400 ;
        RECT 691.950 27.600 694.050 28.200 ;
        RECT 703.950 27.600 706.050 28.200 ;
        RECT 691.950 26.400 706.050 27.600 ;
        RECT 691.950 26.100 694.050 26.400 ;
        RECT 703.950 26.100 706.050 26.400 ;
        RECT 751.950 26.100 754.050 28.200 ;
        RECT 756.000 27.600 760.050 28.050 ;
        RECT 739.950 24.600 742.050 25.050 ;
        RECT 752.400 24.600 753.600 26.100 ;
        RECT 739.950 23.400 753.600 24.600 ;
        RECT 755.400 25.950 760.050 27.600 ;
        RECT 781.950 27.600 784.050 28.050 ;
        RECT 790.950 27.600 793.050 28.200 ;
        RECT 781.950 26.400 793.050 27.600 ;
        RECT 781.950 25.950 784.050 26.400 ;
        RECT 790.950 26.100 793.050 26.400 ;
        RECT 808.950 27.750 811.050 28.200 ;
        RECT 814.950 27.750 817.050 28.200 ;
        RECT 808.950 26.550 817.050 27.750 ;
        RECT 831.000 27.600 835.050 28.050 ;
        RECT 808.950 26.100 811.050 26.550 ;
        RECT 814.950 26.100 817.050 26.550 ;
        RECT 830.400 25.950 835.050 27.600 ;
        RECT 739.950 22.950 742.050 23.400 ;
        RECT 493.950 21.600 496.050 21.900 ;
        RECT 487.950 20.400 496.050 21.600 ;
        RECT 487.950 19.950 490.050 20.400 ;
        RECT 493.950 19.800 496.050 20.400 ;
        RECT 508.950 21.450 511.050 21.900 ;
        RECT 514.950 21.450 517.050 21.900 ;
        RECT 508.950 20.250 517.050 21.450 ;
        RECT 508.950 19.800 511.050 20.250 ;
        RECT 514.950 19.800 517.050 20.250 ;
        RECT 562.950 19.800 565.050 21.900 ;
        RECT 574.950 21.450 577.050 21.900 ;
        RECT 580.950 21.450 583.050 21.900 ;
        RECT 574.950 20.250 583.050 21.450 ;
        RECT 574.950 19.800 577.050 20.250 ;
        RECT 580.950 19.800 583.050 20.250 ;
        RECT 586.950 21.450 589.050 21.900 ;
        RECT 595.950 21.450 598.050 21.900 ;
        RECT 586.950 20.250 598.050 21.450 ;
        RECT 586.950 19.800 589.050 20.250 ;
        RECT 595.950 19.800 598.050 20.250 ;
        RECT 601.950 19.800 604.050 21.900 ;
        RECT 607.950 21.600 610.050 21.900 ;
        RECT 622.950 21.600 625.050 21.900 ;
        RECT 607.950 20.400 625.050 21.600 ;
        RECT 607.950 19.800 610.050 20.400 ;
        RECT 622.950 19.800 625.050 20.400 ;
        RECT 628.950 19.800 631.050 21.900 ;
        RECT 643.950 19.800 646.050 21.900 ;
        RECT 649.950 19.800 652.050 21.900 ;
        RECT 661.950 19.800 664.050 21.900 ;
        RECT 673.800 19.950 675.900 22.050 ;
        RECT 676.950 21.450 679.050 21.900 ;
        RECT 682.950 21.450 685.050 21.900 ;
        RECT 676.950 20.250 685.050 21.450 ;
        RECT 676.950 19.800 679.050 20.250 ;
        RECT 682.950 19.800 685.050 20.250 ;
        RECT 712.950 21.450 715.050 21.900 ;
        RECT 718.950 21.450 721.050 21.900 ;
        RECT 712.950 20.250 721.050 21.450 ;
        RECT 712.950 19.800 715.050 20.250 ;
        RECT 718.950 19.800 721.050 20.250 ;
        RECT 748.950 21.600 751.050 21.900 ;
        RECT 755.400 21.600 756.600 25.950 ;
        RECT 748.950 20.400 756.600 21.600 ;
        RECT 772.950 21.600 775.050 21.900 ;
        RECT 787.950 21.600 790.050 21.900 ;
        RECT 772.950 20.400 790.050 21.600 ;
        RECT 748.950 19.800 751.050 20.400 ;
        RECT 772.950 19.800 775.050 20.400 ;
        RECT 787.950 19.800 790.050 20.400 ;
        RECT 796.950 21.600 799.050 22.050 ;
        RECT 830.400 21.900 831.600 25.950 ;
        RECT 839.400 24.600 840.600 28.950 ;
        RECT 839.400 23.400 846.600 24.600 ;
        RECT 845.400 21.900 846.600 23.400 ;
        RECT 851.400 21.900 852.600 28.950 ;
        RECT 805.950 21.600 808.050 21.900 ;
        RECT 796.950 20.400 808.050 21.600 ;
        RECT 796.950 19.950 799.050 20.400 ;
        RECT 805.950 19.800 808.050 20.400 ;
        RECT 829.950 19.800 832.050 21.900 ;
        RECT 844.950 19.800 847.050 21.900 ;
        RECT 850.950 19.800 853.050 21.900 ;
        RECT 856.950 21.600 859.050 22.050 ;
        RECT 862.950 21.600 865.050 21.900 ;
        RECT 856.950 20.400 865.050 21.600 ;
        RECT 856.950 19.950 859.050 20.400 ;
        RECT 862.950 19.800 865.050 20.400 ;
        RECT 136.950 18.600 139.050 19.050 ;
        RECT 151.950 18.600 154.050 19.050 ;
        RECT 136.950 17.400 154.050 18.600 ;
        RECT 136.950 16.950 139.050 17.400 ;
        RECT 151.950 16.950 154.050 17.400 ;
        RECT 214.950 18.600 217.050 19.050 ;
        RECT 247.950 18.600 250.050 19.050 ;
        RECT 214.950 17.400 250.050 18.600 ;
        RECT 214.950 16.950 217.050 17.400 ;
        RECT 247.950 16.950 250.050 17.400 ;
        RECT 370.950 18.600 373.050 19.050 ;
        RECT 376.950 18.600 379.050 19.050 ;
        RECT 370.950 17.400 379.050 18.600 ;
        RECT 370.950 16.950 373.050 17.400 ;
        RECT 376.950 16.950 379.050 17.400 ;
        RECT 403.950 18.600 406.050 19.050 ;
        RECT 418.950 18.600 421.050 19.050 ;
        RECT 403.950 17.400 421.050 18.600 ;
        RECT 403.950 16.950 406.050 17.400 ;
        RECT 418.950 16.950 421.050 17.400 ;
        RECT 457.950 18.600 460.050 19.050 ;
        RECT 475.950 18.600 478.050 19.050 ;
        RECT 457.950 17.400 478.050 18.600 ;
        RECT 457.950 16.950 460.050 17.400 ;
        RECT 475.950 16.950 478.050 17.400 ;
        RECT 706.950 18.600 709.050 19.050 ;
        RECT 733.950 18.600 736.050 19.050 ;
        RECT 739.950 18.600 742.050 19.050 ;
        RECT 745.950 18.600 748.050 18.750 ;
        RECT 706.950 17.400 748.050 18.600 ;
        RECT 706.950 16.950 709.050 17.400 ;
        RECT 733.950 16.950 736.050 17.400 ;
        RECT 739.950 16.950 742.050 17.400 ;
        RECT 745.950 16.650 748.050 17.400 ;
        RECT 16.950 15.600 19.050 16.050 ;
        RECT 49.950 15.600 52.050 16.050 ;
        RECT 16.950 14.400 52.050 15.600 ;
        RECT 16.950 13.950 19.050 14.400 ;
        RECT 49.950 13.950 52.050 14.400 ;
        RECT 73.950 15.600 76.050 16.050 ;
        RECT 85.950 15.600 88.050 16.050 ;
        RECT 121.950 15.600 124.050 16.050 ;
        RECT 73.950 14.400 124.050 15.600 ;
        RECT 73.950 13.950 76.050 14.400 ;
        RECT 85.950 13.950 88.050 14.400 ;
        RECT 121.950 13.950 124.050 14.400 ;
        RECT 274.950 15.600 277.050 16.050 ;
        RECT 292.950 15.600 295.050 16.050 ;
        RECT 274.950 14.400 295.050 15.600 ;
        RECT 274.950 13.950 277.050 14.400 ;
        RECT 292.950 13.950 295.050 14.400 ;
        RECT 319.950 15.600 322.050 16.050 ;
        RECT 334.950 15.600 337.050 16.050 ;
        RECT 319.950 14.400 337.050 15.600 ;
        RECT 319.950 13.950 322.050 14.400 ;
        RECT 334.950 13.950 337.050 14.400 ;
        RECT 358.950 15.600 361.050 16.050 ;
        RECT 385.950 15.600 388.050 16.050 ;
        RECT 358.950 14.400 388.050 15.600 ;
        RECT 358.950 13.950 361.050 14.400 ;
        RECT 385.950 13.950 388.050 14.400 ;
        RECT 394.950 15.600 397.050 16.050 ;
        RECT 400.950 15.600 403.050 16.050 ;
        RECT 394.950 14.400 403.050 15.600 ;
        RECT 394.950 13.950 397.050 14.400 ;
        RECT 400.950 13.950 403.050 14.400 ;
        RECT 412.950 15.600 415.050 16.050 ;
        RECT 454.950 15.600 457.050 16.050 ;
        RECT 412.950 14.400 457.050 15.600 ;
        RECT 412.950 13.950 415.050 14.400 ;
        RECT 454.950 13.950 457.050 14.400 ;
        RECT 490.950 15.600 493.050 16.050 ;
        RECT 541.950 15.600 544.050 16.050 ;
        RECT 490.950 14.400 544.050 15.600 ;
        RECT 490.950 13.950 493.050 14.400 ;
        RECT 541.950 13.950 544.050 14.400 ;
        RECT 547.950 15.600 550.050 16.050 ;
        RECT 586.950 15.600 589.050 16.050 ;
        RECT 547.950 14.400 589.050 15.600 ;
        RECT 547.950 13.950 550.050 14.400 ;
        RECT 586.950 13.950 589.050 14.400 ;
        RECT 613.950 15.600 616.050 16.050 ;
        RECT 655.950 15.600 658.050 16.050 ;
        RECT 613.950 14.400 658.050 15.600 ;
        RECT 613.950 13.950 616.050 14.400 ;
        RECT 655.950 13.950 658.050 14.400 ;
        RECT 667.950 15.600 670.050 16.050 ;
        RECT 688.950 15.600 691.050 16.050 ;
        RECT 667.950 14.400 691.050 15.600 ;
        RECT 667.950 13.950 670.050 14.400 ;
        RECT 688.950 13.950 691.050 14.400 ;
        RECT 754.950 15.600 757.050 16.050 ;
        RECT 760.950 15.600 763.050 16.050 ;
        RECT 781.950 15.600 784.050 16.050 ;
        RECT 754.950 14.400 784.050 15.600 ;
        RECT 754.950 13.950 757.050 14.400 ;
        RECT 760.950 13.950 763.050 14.400 ;
        RECT 781.950 13.950 784.050 14.400 ;
        RECT 244.950 12.600 247.050 13.050 ;
        RECT 460.950 12.600 463.050 13.050 ;
        RECT 244.950 11.400 463.050 12.600 ;
        RECT 244.950 10.950 247.050 11.400 ;
        RECT 460.950 10.950 463.050 11.400 ;
        RECT 502.950 12.600 505.050 13.050 ;
        RECT 520.950 12.600 523.050 13.050 ;
        RECT 502.950 11.400 523.050 12.600 ;
        RECT 502.950 10.950 505.050 11.400 ;
        RECT 520.950 10.950 523.050 11.400 ;
        RECT 535.950 12.600 538.050 13.050 ;
        RECT 610.950 12.600 613.050 13.050 ;
        RECT 535.950 11.400 613.050 12.600 ;
        RECT 535.950 10.950 538.050 11.400 ;
        RECT 610.950 10.950 613.050 11.400 ;
        RECT 697.950 12.600 700.050 13.050 ;
        RECT 724.950 12.600 727.050 13.050 ;
        RECT 697.950 11.400 727.050 12.600 ;
        RECT 697.950 10.950 700.050 11.400 ;
        RECT 724.950 10.950 727.050 11.400 ;
        RECT 247.950 9.600 250.050 10.050 ;
        RECT 319.950 9.600 322.050 10.050 ;
        RECT 247.950 8.400 322.050 9.600 ;
        RECT 247.950 7.950 250.050 8.400 ;
        RECT 319.950 7.950 322.050 8.400 ;
        RECT 328.950 9.600 331.050 10.050 ;
        RECT 457.950 9.600 460.050 10.050 ;
        RECT 328.950 8.400 460.050 9.600 ;
        RECT 328.950 7.950 331.050 8.400 ;
        RECT 457.950 7.950 460.050 8.400 ;
        RECT 79.950 6.600 82.050 7.050 ;
        RECT 214.950 6.600 217.050 7.050 ;
        RECT 79.950 5.400 217.050 6.600 ;
        RECT 79.950 4.950 82.050 5.400 ;
        RECT 214.950 4.950 217.050 5.400 ;
        RECT 220.950 6.600 223.050 7.050 ;
        RECT 298.950 6.600 301.050 7.050 ;
        RECT 220.950 5.400 301.050 6.600 ;
        RECT 220.950 4.950 223.050 5.400 ;
        RECT 298.950 4.950 301.050 5.400 ;
        RECT 412.950 6.600 415.050 7.050 ;
        RECT 451.950 6.600 454.050 7.050 ;
        RECT 412.950 5.400 454.050 6.600 ;
        RECT 412.950 4.950 415.050 5.400 ;
        RECT 451.950 4.950 454.050 5.400 ;
        RECT 460.950 6.600 463.050 7.050 ;
        RECT 556.950 6.600 559.050 7.050 ;
        RECT 460.950 5.400 559.050 6.600 ;
        RECT 460.950 4.950 463.050 5.400 ;
        RECT 556.950 4.950 559.050 5.400 ;
        RECT 592.950 6.600 595.050 7.050 ;
        RECT 736.950 6.600 739.050 7.050 ;
        RECT 592.950 5.400 739.050 6.600 ;
        RECT 592.950 4.950 595.050 5.400 ;
        RECT 736.950 4.950 739.050 5.400 ;
        RECT 595.950 3.600 598.050 4.050 ;
        RECT 673.950 3.600 676.050 4.050 ;
        RECT 595.950 2.400 676.050 3.600 ;
        RECT 595.950 1.950 598.050 2.400 ;
        RECT 673.950 1.950 676.050 2.400 ;
  END
END fir_pe
END LIBRARY

