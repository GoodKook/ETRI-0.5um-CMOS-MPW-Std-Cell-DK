magic
tech scmos
magscale 1 2
timestamp 1754220398
<< metal1 >>
rect -62 4338 -2 4578
rect 4750 4562 4842 4578
rect 3117 4517 3133 4523
rect 497 4447 503 4493
rect 3117 4447 3123 4517
rect -62 4322 30 4338
rect -62 3858 -2 4322
rect 4782 4098 4842 4562
rect 4750 4082 4842 4098
rect 4347 4017 4363 4023
rect 4357 3967 4363 4017
rect -62 3842 30 3858
rect -62 3378 -2 3842
rect 537 3757 553 3763
rect 537 3687 543 3757
rect 757 3703 763 3753
rect 747 3697 763 3703
rect 4782 3618 4842 4082
rect 4750 3602 4842 3618
rect 937 3557 953 3563
rect 937 3467 943 3557
rect 3397 3483 3403 3533
rect 3397 3477 3413 3483
rect -62 3362 30 3378
rect -62 2898 -2 3362
rect 1727 3297 1773 3303
rect 397 3283 403 3293
rect 377 3277 403 3283
rect 1577 3277 1593 3283
rect 377 3227 383 3277
rect 1577 3183 1583 3277
rect 1907 3277 1923 3283
rect 1917 3203 1923 3277
rect 1917 3197 1933 3203
rect 1567 3177 1583 3183
rect 4782 3138 4842 3602
rect 4750 3122 4842 3138
rect 557 3057 573 3063
rect 557 2963 563 3057
rect 1827 3037 1843 3043
rect 1837 2987 1843 3037
rect 4277 3007 4283 3073
rect 4737 3007 4743 3073
rect 547 2957 563 2963
rect -62 2882 30 2898
rect -62 2418 -2 2882
rect 1937 2727 1943 2773
rect 4782 2658 4842 3122
rect 4750 2642 4842 2658
rect 477 2597 493 2603
rect 477 2523 483 2597
rect 807 2577 823 2583
rect 547 2557 593 2563
rect 467 2517 483 2523
rect 817 2503 823 2577
rect 807 2497 823 2503
rect -62 2402 30 2418
rect -62 1938 -2 2402
rect 117 2337 133 2343
rect 117 2263 123 2337
rect 3737 2317 3773 2323
rect 3737 2287 3743 2317
rect 107 2257 123 2263
rect 3957 2243 3963 2293
rect 3947 2237 3963 2243
rect 4782 2178 4842 2642
rect 4750 2162 4842 2178
rect 1277 2097 1293 2103
rect 97 2077 113 2083
rect 97 2003 103 2077
rect 1087 2077 1113 2083
rect 1277 2047 1283 2097
rect 1447 2097 1463 2103
rect 1377 2023 1383 2053
rect 1367 2017 1383 2023
rect 1457 2023 1463 2097
rect 1457 2017 1473 2023
rect 97 1997 113 2003
rect -62 1922 30 1938
rect -62 1458 -2 1922
rect 1117 1857 1133 1863
rect 217 1783 223 1833
rect 207 1777 223 1783
rect 1117 1783 1123 1857
rect 3897 1857 3913 1863
rect 1117 1777 1153 1783
rect 3897 1783 3903 1857
rect 3897 1777 3913 1783
rect 4782 1698 4842 2162
rect 4750 1682 4842 1698
rect 1267 1637 1283 1643
rect 257 1617 273 1623
rect 257 1543 263 1617
rect 257 1537 273 1543
rect 1077 1543 1083 1613
rect 1277 1563 1283 1637
rect 1997 1597 2033 1603
rect 1277 1557 1293 1563
rect 1997 1547 2003 1597
rect 2117 1597 2133 1603
rect 1077 1537 1093 1543
rect 2117 1543 2123 1597
rect 3357 1597 3373 1603
rect 2107 1537 2123 1543
rect 3357 1523 3363 1597
rect 4217 1567 4223 1613
rect 3357 1517 3373 1523
rect 4677 1523 4683 1613
rect 4667 1517 4683 1523
rect -62 1442 30 1458
rect -62 978 -2 1442
rect 1417 1377 1433 1383
rect 197 1303 203 1353
rect 197 1297 213 1303
rect 297 1287 303 1353
rect 477 1307 483 1353
rect 1417 1303 1423 1377
rect 1417 1297 1433 1303
rect 4782 1218 4842 1682
rect 4750 1202 4842 1218
rect 487 1157 503 1163
rect 297 1087 303 1133
rect 497 1083 503 1157
rect 1587 1137 1603 1143
rect 867 1117 903 1123
rect 497 1077 513 1083
rect 897 1047 903 1117
rect 1597 1063 1603 1137
rect 2227 1117 2263 1123
rect 2257 1063 2263 1117
rect 1597 1057 1623 1063
rect 2257 1057 2273 1063
rect 1617 1047 1623 1057
rect -62 962 30 978
rect -62 498 -2 962
rect 1587 877 1603 883
rect 1597 867 1603 877
rect 1617 823 1623 933
rect 1617 817 1633 823
rect 4782 738 4842 1202
rect 4750 722 4842 738
rect 2137 677 2153 683
rect 2137 663 2143 677
rect 2117 657 2143 663
rect 1907 637 1923 643
rect 1917 563 1923 637
rect 2117 587 2123 657
rect 1907 557 1923 563
rect 2237 563 2243 633
rect 2227 557 2243 563
rect -62 482 30 498
rect -62 18 -2 482
rect 247 397 263 403
rect 257 347 263 397
rect 427 397 443 403
rect 437 307 443 397
rect 2187 397 2203 403
rect 1737 343 1743 353
rect 1737 337 1753 343
rect 2017 323 2023 373
rect 2097 327 2103 393
rect 2197 347 2203 397
rect 2017 317 2033 323
rect 4782 258 4842 722
rect 4750 242 4842 258
rect 597 107 603 173
rect 977 127 983 193
rect -62 2 30 18
rect 4782 2 4842 242
<< m2contact >>
rect 493 4493 507 4507
rect 3133 4513 3147 4527
rect 493 4433 507 4447
rect 3113 4433 3127 4447
rect 4333 4013 4347 4027
rect 4353 3953 4367 3967
rect 553 3753 567 3767
rect 753 3753 767 3767
rect 733 3693 747 3707
rect 533 3673 547 3687
rect 953 3553 967 3567
rect 3393 3533 3407 3547
rect 3413 3473 3427 3487
rect 933 3453 947 3467
rect 393 3293 407 3307
rect 1713 3293 1727 3307
rect 1773 3293 1787 3307
rect 373 3213 387 3227
rect 1553 3173 1567 3187
rect 1593 3273 1607 3287
rect 1893 3273 1907 3287
rect 1933 3193 1947 3207
rect 4273 3073 4287 3087
rect 4733 3073 4747 3087
rect 533 2953 547 2967
rect 573 3053 587 3067
rect 1813 3033 1827 3047
rect 4273 2993 4287 3007
rect 4733 2993 4747 3007
rect 1833 2973 1847 2987
rect 1933 2773 1947 2787
rect 1933 2713 1947 2727
rect 453 2513 467 2527
rect 493 2593 507 2607
rect 793 2573 807 2587
rect 533 2553 547 2567
rect 593 2553 607 2567
rect 793 2493 807 2507
rect 93 2253 107 2267
rect 133 2333 147 2347
rect 3773 2313 3787 2327
rect 3953 2293 3967 2307
rect 3733 2273 3747 2287
rect 3933 2233 3947 2247
rect 113 2073 127 2087
rect 1073 2073 1087 2087
rect 1113 2073 1127 2087
rect 1293 2093 1307 2107
rect 1433 2093 1447 2107
rect 1373 2053 1387 2067
rect 1273 2033 1287 2047
rect 1353 2013 1367 2027
rect 1473 2013 1487 2027
rect 113 1993 127 2007
rect 213 1833 227 1847
rect 193 1773 207 1787
rect 1133 1853 1147 1867
rect 1153 1773 1167 1787
rect 3913 1853 3927 1867
rect 3913 1773 3927 1787
rect 1253 1633 1267 1647
rect 273 1613 287 1627
rect 1073 1613 1087 1627
rect 273 1533 287 1547
rect 4213 1613 4227 1627
rect 4673 1613 4687 1627
rect 1293 1553 1307 1567
rect 2033 1593 2047 1607
rect 1093 1533 1107 1547
rect 1993 1533 2007 1547
rect 2093 1533 2107 1547
rect 2133 1593 2147 1607
rect 3373 1593 3387 1607
rect 4213 1553 4227 1567
rect 3373 1513 3387 1527
rect 4653 1513 4667 1527
rect 193 1353 207 1367
rect 293 1353 307 1367
rect 473 1353 487 1367
rect 213 1293 227 1307
rect 473 1293 487 1307
rect 1433 1373 1447 1387
rect 1433 1293 1447 1307
rect 293 1273 307 1287
rect 473 1153 487 1167
rect 293 1133 307 1147
rect 293 1073 307 1087
rect 1573 1133 1587 1147
rect 853 1113 867 1127
rect 513 1073 527 1087
rect 2213 1113 2227 1127
rect 2273 1053 2287 1067
rect 893 1033 907 1047
rect 1613 1033 1627 1047
rect 1613 933 1627 947
rect 1573 873 1587 887
rect 1593 853 1607 867
rect 1633 813 1647 827
rect 2153 673 2167 687
rect 1893 633 1907 647
rect 1893 553 1907 567
rect 2233 633 2247 647
rect 2113 573 2127 587
rect 2213 553 2227 567
rect 233 393 247 407
rect 413 393 427 407
rect 253 333 267 347
rect 2093 393 2107 407
rect 2173 393 2187 407
rect 2013 373 2027 387
rect 1733 353 1747 367
rect 1753 333 1767 347
rect 2193 333 2207 347
rect 2033 313 2047 327
rect 2093 313 2107 327
rect 433 293 447 307
rect 973 193 987 207
rect 593 173 607 187
rect 973 113 987 127
rect 593 93 607 107
<< metal2 >>
rect 3996 4616 4023 4623
rect 36 4476 43 4513
rect 56 4407 63 4463
rect 96 4427 103 4453
rect 116 4407 123 4533
rect 176 4487 183 4493
rect 176 4447 183 4473
rect 196 4456 203 4533
rect 496 4507 503 4513
rect 216 4456 223 4473
rect 136 4367 143 4443
rect 236 4436 243 4453
rect 36 4216 43 4233
rect 96 4207 103 4233
rect 156 4227 163 4413
rect 56 4147 63 4203
rect 56 3976 63 4033
rect 76 4027 83 4173
rect 116 3976 123 4153
rect 156 4107 163 4183
rect 176 4127 183 4393
rect 16 3956 33 3963
rect 16 3703 23 3956
rect 76 3956 103 3963
rect 56 3727 63 3893
rect 76 3747 83 3956
rect 136 3947 143 3963
rect 136 3747 143 3933
rect 156 3887 163 4073
rect 176 3943 183 4113
rect 196 4067 203 4413
rect 316 4227 323 4453
rect 376 4447 383 4493
rect 496 4476 523 4483
rect 556 4476 563 4493
rect 396 4456 403 4473
rect 496 4467 503 4476
rect 656 4476 663 4493
rect 336 4407 343 4443
rect 416 4287 423 4453
rect 456 4327 463 4453
rect 536 4447 543 4463
rect 576 4456 603 4463
rect 507 4436 513 4443
rect 596 4367 603 4456
rect 256 4216 283 4223
rect 216 3976 223 4013
rect 256 3987 263 4173
rect 276 4087 283 4216
rect 356 4187 363 4273
rect 296 4147 303 4173
rect 336 4087 343 4183
rect 376 4127 383 4203
rect 436 4176 463 4183
rect 436 4107 443 4176
rect 516 4127 523 4193
rect 556 4167 563 4353
rect 576 4196 583 4313
rect 616 4183 623 4433
rect 636 4427 643 4463
rect 656 4387 663 4433
rect 696 4407 703 4453
rect 716 4443 723 4513
rect 756 4496 863 4503
rect 756 4487 763 4496
rect 856 4487 863 4496
rect 716 4436 743 4443
rect 776 4436 783 4473
rect 836 4447 843 4473
rect 896 4423 903 4533
rect 1056 4516 1143 4523
rect 1056 4507 1063 4516
rect 1136 4507 1143 4516
rect 996 4456 1003 4473
rect 916 4427 923 4443
rect 876 4416 903 4423
rect 656 4196 663 4213
rect 616 4176 643 4183
rect 716 4167 723 4413
rect 736 4196 743 4373
rect 816 4367 823 4413
rect 856 4223 863 4413
rect 836 4216 863 4223
rect 596 4147 603 4163
rect 296 3996 303 4053
rect 376 4016 383 4033
rect 336 3996 343 4013
rect 416 3996 423 4033
rect 456 3996 483 4003
rect 176 3936 203 3943
rect 16 3696 43 3703
rect 36 3627 43 3696
rect 76 3667 83 3693
rect 96 3647 103 3703
rect 56 3496 63 3633
rect 116 3627 123 3673
rect 136 3667 143 3703
rect 16 3427 23 3473
rect 16 3207 23 3393
rect 36 3287 43 3483
rect 96 3463 103 3613
rect 116 3487 123 3593
rect 76 3456 103 3463
rect 36 3183 43 3273
rect 16 3176 43 3183
rect 16 2947 23 3176
rect 76 3036 83 3456
rect 96 3267 103 3433
rect 116 3267 123 3473
rect 96 3167 103 3193
rect 116 3123 123 3253
rect 136 3207 143 3223
rect 156 3187 163 3693
rect 176 3667 183 3873
rect 176 3516 183 3533
rect 196 3483 203 3936
rect 236 3903 243 3963
rect 256 3903 263 3913
rect 316 3907 323 3983
rect 356 3976 383 3983
rect 236 3896 263 3903
rect 256 3703 263 3896
rect 356 3727 363 3953
rect 376 3887 383 3976
rect 396 3907 403 3983
rect 436 3927 443 3993
rect 456 3947 463 3996
rect 536 3927 543 3963
rect 576 3947 583 3963
rect 596 3907 603 4113
rect 656 3996 663 4053
rect 256 3696 283 3703
rect 236 3647 243 3673
rect 216 3516 243 3523
rect 176 3476 203 3483
rect 176 3247 183 3476
rect 136 3147 143 3173
rect 176 3143 183 3213
rect 236 3207 243 3516
rect 256 3367 263 3673
rect 296 3447 303 3523
rect 296 3407 303 3433
rect 176 3136 203 3143
rect 116 3116 143 3123
rect 16 2707 23 2773
rect 36 2767 43 2993
rect 56 2987 63 3023
rect 136 3003 143 3116
rect 156 3036 163 3053
rect 136 2996 163 3003
rect 56 2767 63 2913
rect 76 2847 83 2993
rect 96 2823 103 2973
rect 76 2816 103 2823
rect 36 2587 43 2713
rect 56 2707 63 2723
rect 16 2536 23 2553
rect 36 2516 43 2573
rect 56 2547 63 2653
rect 76 2567 83 2816
rect 156 2787 163 2996
rect 176 2947 183 3003
rect 176 2843 183 2933
rect 196 2867 203 3136
rect 236 3043 243 3113
rect 256 3087 263 3333
rect 316 3327 323 3633
rect 356 3587 363 3693
rect 376 3667 383 3703
rect 416 3687 423 3753
rect 456 3736 483 3743
rect 436 3647 443 3703
rect 456 3647 463 3736
rect 536 3707 543 3893
rect 556 3736 563 3753
rect 596 3736 603 3753
rect 636 3716 643 3753
rect 516 3667 523 3693
rect 336 3503 343 3573
rect 376 3543 383 3613
rect 536 3587 543 3673
rect 376 3536 403 3543
rect 336 3496 363 3503
rect 376 3467 383 3493
rect 396 3343 403 3536
rect 516 3516 523 3533
rect 476 3483 483 3513
rect 416 3467 423 3483
rect 456 3476 483 3483
rect 376 3336 403 3343
rect 296 3236 303 3273
rect 336 3236 343 3273
rect 376 3247 383 3336
rect 456 3327 463 3476
rect 396 3307 403 3313
rect 396 3256 403 3273
rect 276 3127 283 3223
rect 316 3203 323 3223
rect 316 3196 343 3203
rect 336 3187 343 3196
rect 216 3036 243 3043
rect 176 2836 203 2843
rect 96 2667 103 2763
rect 136 2756 143 2773
rect 196 2767 203 2836
rect 216 2787 223 2993
rect 236 2827 243 3036
rect 256 2907 263 3043
rect 296 3027 303 3133
rect 276 2747 283 2813
rect 296 2787 303 2993
rect 316 2927 323 3173
rect 356 3043 363 3193
rect 376 3187 383 3213
rect 336 3036 363 3043
rect 356 2887 363 3036
rect 376 2967 383 2993
rect 396 2943 403 3153
rect 436 3127 443 3213
rect 456 3187 463 3293
rect 476 3227 483 3253
rect 436 2967 443 3113
rect 376 2936 403 2943
rect 336 2776 343 2793
rect 376 2787 383 2936
rect 396 2776 423 2783
rect 16 2327 23 2493
rect 36 2327 43 2393
rect 76 2343 83 2523
rect 96 2363 103 2613
rect 156 2607 163 2743
rect 176 2627 183 2733
rect 196 2683 203 2713
rect 216 2707 223 2743
rect 196 2676 223 2683
rect 176 2556 203 2563
rect 96 2356 123 2363
rect 76 2336 103 2343
rect 96 2327 103 2336
rect 16 2296 43 2303
rect 16 2187 23 2296
rect 76 2267 83 2303
rect 56 2256 73 2263
rect 16 2007 23 2173
rect 36 2076 43 2253
rect 56 2107 63 2256
rect 76 2076 83 2093
rect 16 1727 23 1873
rect 36 1823 43 1853
rect 56 1847 63 2073
rect 96 2063 103 2253
rect 116 2087 123 2356
rect 136 2347 143 2353
rect 196 2307 203 2556
rect 216 2407 223 2676
rect 256 2576 263 2593
rect 296 2563 303 2713
rect 316 2667 323 2763
rect 356 2727 363 2773
rect 396 2767 403 2776
rect 396 2723 403 2753
rect 376 2716 403 2723
rect 276 2556 303 2563
rect 256 2303 263 2533
rect 276 2367 283 2556
rect 336 2467 343 2693
rect 356 2556 363 2613
rect 376 2527 383 2716
rect 416 2667 423 2733
rect 436 2576 443 2613
rect 456 2587 463 3153
rect 476 3036 483 3093
rect 516 3087 523 3313
rect 536 3067 543 3353
rect 556 3307 563 3473
rect 556 3207 563 3223
rect 576 3167 583 3693
rect 656 3683 663 3933
rect 696 3927 703 4153
rect 776 4147 783 4193
rect 816 4187 823 4203
rect 856 4187 863 4216
rect 876 4167 883 4416
rect 956 4367 963 4433
rect 1056 4407 1063 4443
rect 1076 4367 1083 4493
rect 1096 4427 1103 4453
rect 1136 4447 1143 4463
rect 1176 4427 1183 4473
rect 1236 4456 1243 4553
rect 1276 4467 1283 4493
rect 1296 4476 1303 4533
rect 916 4227 923 4353
rect 996 4216 1023 4223
rect 916 4196 923 4213
rect 996 4183 1003 4216
rect 1156 4216 1163 4353
rect 1196 4223 1203 4453
rect 1216 4387 1223 4443
rect 1256 4407 1263 4433
rect 1356 4427 1363 4493
rect 1436 4476 1443 4513
rect 1456 4507 1463 4533
rect 1416 4407 1423 4463
rect 1456 4443 1463 4493
rect 1536 4476 1543 4553
rect 1496 4456 1503 4473
rect 1616 4456 1623 4513
rect 1456 4436 1483 4443
rect 1556 4407 1563 4453
rect 1596 4427 1603 4453
rect 1636 4436 1643 4533
rect 1696 4447 1703 4513
rect 1816 4496 1823 4513
rect 1956 4496 1963 4513
rect 1716 4476 1743 4483
rect 1676 4267 1683 4443
rect 1196 4216 1223 4223
rect 1256 4216 1283 4223
rect 936 4167 943 4183
rect 976 4176 1003 4183
rect 1036 4147 1043 4203
rect 716 3963 723 4013
rect 776 4007 783 4133
rect 796 3976 803 4053
rect 856 3976 863 4033
rect 716 3956 743 3963
rect 896 3963 903 4133
rect 936 3976 943 4033
rect 956 3996 963 4033
rect 1056 3996 1063 4213
rect 1076 4127 1083 4203
rect 1096 4196 1123 4203
rect 1076 3976 1083 4053
rect 876 3956 903 3963
rect 756 3767 763 3933
rect 836 3743 843 3773
rect 756 3736 783 3743
rect 816 3736 843 3743
rect 756 3707 763 3736
rect 716 3696 733 3703
rect 836 3687 843 3736
rect 596 3496 603 3573
rect 616 3516 623 3683
rect 656 3676 683 3683
rect 656 3527 663 3593
rect 676 3567 683 3676
rect 696 3627 703 3673
rect 596 3267 603 3293
rect 596 3107 603 3173
rect 616 3167 623 3393
rect 636 3347 643 3503
rect 676 3467 683 3483
rect 656 3187 663 3253
rect 316 2327 323 2353
rect 356 2327 363 2513
rect 416 2347 423 2413
rect 236 2296 263 2303
rect 236 2287 243 2296
rect 136 2267 143 2283
rect 156 2207 163 2263
rect 196 2247 203 2263
rect 216 2247 223 2263
rect 176 2087 183 2133
rect 216 2087 223 2213
rect 236 2087 243 2213
rect 256 2087 263 2263
rect 276 2227 283 2273
rect 296 2247 303 2293
rect 336 2267 343 2303
rect 376 2296 403 2303
rect 336 2247 343 2253
rect 256 2063 263 2073
rect 276 2067 283 2153
rect 316 2096 323 2173
rect 356 2107 363 2193
rect 96 2056 123 2063
rect 76 1827 83 2033
rect 96 1887 103 2033
rect 116 1847 123 1993
rect 36 1816 63 1823
rect 56 1796 63 1816
rect 96 1796 103 1813
rect 156 1807 163 2063
rect 236 2056 263 2063
rect 176 1987 183 2033
rect 216 1967 223 2043
rect 236 1947 243 2013
rect 216 1847 223 1853
rect 236 1847 243 1913
rect 296 1883 303 1933
rect 316 1907 323 2053
rect 336 2047 343 2063
rect 296 1876 323 1883
rect 236 1816 243 1833
rect 296 1823 303 1853
rect 276 1816 303 1823
rect 36 1747 43 1783
rect 96 1627 103 1753
rect 116 1707 123 1783
rect 136 1727 143 1783
rect 176 1747 183 1783
rect 136 1687 143 1713
rect 176 1627 183 1733
rect 56 1616 83 1623
rect 16 1147 23 1593
rect 76 1407 83 1616
rect 176 1576 183 1613
rect 116 1567 123 1573
rect 56 1347 63 1393
rect 136 1387 143 1573
rect 196 1567 203 1773
rect 216 1747 223 1813
rect 256 1767 263 1793
rect 276 1707 283 1773
rect 256 1563 263 1693
rect 276 1627 283 1633
rect 296 1627 303 1816
rect 316 1727 323 1876
rect 376 1867 383 2253
rect 396 2227 403 2296
rect 416 2276 423 2333
rect 436 2287 443 2533
rect 456 2527 463 2543
rect 476 2487 483 2973
rect 496 2947 503 3023
rect 536 2807 543 2953
rect 556 2927 563 3093
rect 576 3067 583 3093
rect 596 3047 603 3073
rect 616 2947 623 3003
rect 556 2827 563 2833
rect 556 2783 563 2813
rect 576 2787 583 2893
rect 636 2883 643 3133
rect 656 2907 663 3153
rect 676 3147 683 3353
rect 696 3243 703 3453
rect 716 3387 723 3483
rect 736 3367 743 3553
rect 756 3547 763 3613
rect 756 3516 763 3533
rect 796 3516 803 3633
rect 836 3527 843 3533
rect 696 3236 723 3243
rect 756 3236 763 3373
rect 776 3347 783 3503
rect 816 3447 823 3503
rect 776 3203 783 3223
rect 796 3207 803 3273
rect 816 3267 823 3433
rect 856 3407 863 3913
rect 876 3807 883 3933
rect 876 3736 883 3793
rect 896 3716 923 3723
rect 916 3687 923 3716
rect 936 3707 943 3723
rect 956 3716 963 3773
rect 976 3727 983 3953
rect 1036 3947 1043 3973
rect 1096 3967 1103 4173
rect 1116 3907 1123 4196
rect 1136 4147 1143 4203
rect 1196 4147 1203 4216
rect 1276 4187 1283 4216
rect 1336 4187 1343 4223
rect 1396 4216 1403 4233
rect 1516 4216 1543 4223
rect 1156 4016 1183 4023
rect 1176 3807 1183 4016
rect 1216 3976 1223 4033
rect 1236 4027 1243 4173
rect 1256 4016 1283 4023
rect 1236 3956 1243 4013
rect 1256 3983 1263 4016
rect 1336 3987 1343 4113
rect 1356 4107 1363 4203
rect 1256 3976 1283 3983
rect 1276 3907 1283 3976
rect 1356 3956 1363 4013
rect 1376 3976 1383 4033
rect 1396 4007 1403 4173
rect 1416 4127 1423 4203
rect 1416 3947 1423 4093
rect 1436 3976 1443 4013
rect 1456 3967 1463 4133
rect 1476 4027 1483 4213
rect 1496 4167 1503 4203
rect 1536 4087 1543 4216
rect 1556 4207 1563 4233
rect 1716 4223 1723 4476
rect 2016 4483 2023 4513
rect 2056 4496 2063 4513
rect 2096 4496 2123 4503
rect 2096 4483 2103 4496
rect 2016 4476 2043 4483
rect 2076 4476 2103 4483
rect 2176 4476 2183 4493
rect 2016 4467 2023 4476
rect 1756 4407 1763 4463
rect 1796 4327 1803 4463
rect 1836 4447 1843 4463
rect 1936 4327 1943 4463
rect 1976 4447 1983 4463
rect 1716 4216 1743 4223
rect 1736 4207 1743 4216
rect 1796 4203 1803 4233
rect 1896 4207 1903 4313
rect 1776 4196 1803 4203
rect 1556 4183 1563 4193
rect 1556 4176 1583 4183
rect 1496 4016 1563 4023
rect 1496 4003 1503 4016
rect 1476 3996 1503 4003
rect 1476 3976 1483 3996
rect 996 3716 1003 3753
rect 1036 3747 1043 3793
rect 1056 3707 1063 3713
rect 936 3687 943 3693
rect 1076 3687 1083 3733
rect 1136 3716 1163 3723
rect 836 3236 843 3293
rect 876 3267 883 3493
rect 916 3367 923 3673
rect 936 3483 943 3653
rect 976 3567 983 3673
rect 1076 3607 1083 3633
rect 1096 3607 1103 3713
rect 1136 3707 1143 3716
rect 1216 3687 1223 3703
rect 956 3523 963 3553
rect 996 3527 1003 3573
rect 956 3516 983 3523
rect 976 3496 983 3516
rect 1016 3507 1023 3533
rect 1096 3516 1103 3533
rect 1116 3507 1123 3573
rect 1136 3516 1143 3613
rect 1156 3536 1163 3573
rect 1236 3547 1243 3893
rect 1336 3736 1343 3853
rect 1396 3687 1403 3723
rect 1416 3687 1423 3753
rect 1476 3707 1483 3933
rect 1516 3867 1523 3993
rect 1556 3976 1563 4016
rect 1596 4007 1603 4163
rect 1616 4107 1623 4183
rect 1656 4107 1663 4183
rect 1696 4007 1703 4183
rect 1716 4127 1723 4183
rect 1716 3996 1723 4093
rect 1816 4067 1823 4193
rect 1856 4147 1863 4203
rect 1916 4196 1923 4213
rect 1936 4203 1943 4233
rect 1936 4196 1963 4203
rect 1536 3947 1543 3963
rect 1576 3867 1583 3963
rect 1716 3956 1743 3963
rect 1256 3667 1263 3673
rect 1176 3516 1203 3523
rect 1036 3487 1043 3493
rect 936 3476 963 3483
rect 936 3407 943 3453
rect 1076 3447 1083 3503
rect 916 3256 923 3273
rect 816 3207 823 3223
rect 756 3196 783 3203
rect 636 2876 663 2883
rect 536 2776 563 2783
rect 536 2756 543 2776
rect 616 2776 623 2833
rect 496 2747 503 2753
rect 516 2603 523 2743
rect 507 2596 523 2603
rect 516 2536 523 2573
rect 536 2567 543 2713
rect 536 2547 543 2553
rect 556 2536 563 2593
rect 496 2427 503 2523
rect 576 2507 583 2733
rect 596 2607 603 2763
rect 616 2707 623 2733
rect 656 2707 663 2876
rect 676 2827 683 2973
rect 696 2756 703 2953
rect 716 2807 723 2953
rect 736 2847 743 3193
rect 756 3167 763 3196
rect 776 3056 783 3173
rect 796 3036 803 3093
rect 836 3083 843 3193
rect 876 3167 883 3173
rect 836 3076 863 3083
rect 836 3047 843 3053
rect 856 3047 863 3076
rect 836 3016 843 3033
rect 736 2783 743 2833
rect 756 2807 763 2933
rect 776 2783 783 2973
rect 856 2847 863 3003
rect 876 2967 883 3153
rect 896 2987 903 3213
rect 976 3167 983 3353
rect 996 3247 1003 3273
rect 1016 3256 1023 3393
rect 1096 3387 1103 3473
rect 1096 3347 1103 3373
rect 1036 3236 1063 3243
rect 1056 3223 1063 3236
rect 1056 3216 1073 3223
rect 916 3016 923 3113
rect 936 3036 943 3153
rect 716 2776 743 2783
rect 756 2776 783 2783
rect 676 2683 683 2733
rect 656 2676 683 2683
rect 616 2587 623 2613
rect 616 2556 623 2573
rect 656 2556 663 2676
rect 716 2587 723 2776
rect 756 2756 763 2776
rect 836 2767 843 2813
rect 676 2556 703 2563
rect 596 2536 603 2553
rect 576 2427 583 2493
rect 456 2276 463 2353
rect 516 2303 523 2313
rect 496 2296 523 2303
rect 396 2103 403 2213
rect 396 2096 423 2103
rect 456 2076 463 2113
rect 476 2107 483 2233
rect 496 2083 503 2296
rect 516 2243 523 2263
rect 516 2236 543 2243
rect 476 2076 503 2083
rect 396 1887 403 2033
rect 416 1847 423 2053
rect 436 2047 443 2053
rect 456 1823 463 1853
rect 476 1847 483 2076
rect 516 2063 523 2213
rect 536 2167 543 2236
rect 576 2227 583 2283
rect 596 2267 603 2473
rect 616 2263 623 2513
rect 636 2327 643 2543
rect 676 2387 683 2556
rect 696 2363 703 2513
rect 716 2487 723 2543
rect 776 2536 783 2693
rect 796 2647 803 2763
rect 816 2667 823 2733
rect 796 2587 803 2613
rect 756 2407 763 2513
rect 796 2507 803 2523
rect 816 2487 823 2653
rect 836 2567 843 2653
rect 856 2536 863 2613
rect 876 2547 883 2893
rect 896 2776 903 2833
rect 896 2567 903 2733
rect 936 2647 943 2993
rect 956 2947 963 3023
rect 996 3007 1003 3093
rect 1016 3016 1023 3053
rect 1036 3036 1043 3073
rect 1076 3036 1083 3093
rect 1096 3043 1103 3333
rect 1136 3307 1143 3333
rect 1136 3256 1143 3293
rect 1116 3043 1123 3133
rect 1136 3056 1143 3153
rect 1156 3067 1163 3493
rect 1196 3487 1203 3516
rect 1216 3407 1223 3483
rect 1256 3427 1263 3473
rect 1216 3327 1223 3393
rect 1176 3267 1183 3293
rect 1276 3267 1283 3553
rect 1376 3516 1383 3633
rect 1396 3483 1403 3503
rect 1387 3476 1403 3483
rect 1376 3367 1383 3473
rect 1176 3207 1183 3223
rect 1176 3107 1183 3193
rect 1196 3087 1203 3243
rect 1216 3167 1223 3263
rect 1236 3167 1243 3243
rect 1176 3043 1183 3053
rect 1096 3036 1123 3043
rect 1156 3036 1183 3043
rect 1056 2967 1063 3023
rect 916 2543 923 2573
rect 896 2536 923 2543
rect 936 2536 943 2633
rect 956 2607 963 2773
rect 1016 2767 1023 2953
rect 1096 2947 1103 3036
rect 1176 3027 1183 3036
rect 1196 3016 1203 3073
rect 1216 3036 1223 3113
rect 1256 3036 1263 3073
rect 1276 3047 1283 3233
rect 1296 3087 1303 3223
rect 1336 3207 1343 3223
rect 1376 3123 1383 3353
rect 1436 3256 1443 3333
rect 1416 3167 1423 3243
rect 1356 3116 1383 3123
rect 1296 3016 1303 3073
rect 1176 2887 1183 3013
rect 1356 3003 1363 3116
rect 1396 3103 1403 3133
rect 1376 3096 1403 3103
rect 1376 3036 1383 3096
rect 1056 2776 1063 2813
rect 976 2747 983 2763
rect 1076 2747 1083 2763
rect 976 2587 983 2653
rect 996 2647 1003 2743
rect 956 2556 963 2573
rect 1016 2567 1023 2713
rect 1036 2707 1043 2743
rect 676 2356 703 2363
rect 656 2276 663 2293
rect 676 2287 683 2356
rect 736 2276 743 2293
rect 616 2256 643 2263
rect 656 2236 683 2243
rect 556 2083 563 2193
rect 576 2187 583 2213
rect 656 2207 663 2236
rect 616 2136 663 2143
rect 496 2056 523 2063
rect 536 2076 563 2083
rect 536 2056 543 2076
rect 456 1816 483 1823
rect 56 1316 63 1333
rect 96 1327 103 1373
rect 196 1367 203 1453
rect 236 1387 243 1563
rect 256 1556 283 1563
rect 256 1367 263 1556
rect 316 1547 323 1563
rect 276 1367 283 1533
rect 296 1367 303 1433
rect 336 1363 343 1773
rect 356 1767 363 1803
rect 396 1783 403 1803
rect 436 1796 443 1813
rect 476 1796 483 1816
rect 396 1776 423 1783
rect 356 1427 363 1653
rect 376 1607 383 1773
rect 416 1747 423 1776
rect 516 1747 523 1993
rect 556 1783 563 1913
rect 576 1867 583 2113
rect 616 2036 623 2136
rect 636 2067 643 2113
rect 656 2087 663 2136
rect 616 1787 623 1893
rect 547 1776 563 1783
rect 596 1767 603 1783
rect 636 1767 643 2013
rect 656 1987 663 2043
rect 676 1927 683 2213
rect 716 2187 723 2243
rect 756 2147 763 2353
rect 716 2096 723 2113
rect 776 2107 783 2453
rect 816 2296 823 2393
rect 796 2127 803 2253
rect 836 2247 843 2473
rect 876 2296 883 2393
rect 916 2307 923 2453
rect 756 2076 783 2083
rect 696 1967 703 2053
rect 716 1907 723 2033
rect 736 2007 743 2063
rect 676 1807 683 1813
rect 396 1596 403 1713
rect 416 1647 423 1733
rect 356 1367 363 1393
rect 316 1356 343 1363
rect 36 1127 43 1303
rect 136 1287 143 1343
rect 276 1336 303 1343
rect 156 1307 163 1323
rect 196 1316 223 1323
rect 56 1116 63 1253
rect 96 1116 103 1133
rect 116 1116 123 1133
rect 156 1116 163 1153
rect 176 1127 183 1293
rect 16 947 23 1113
rect 196 1103 203 1316
rect 216 1187 223 1293
rect 236 1147 243 1333
rect 176 1096 203 1103
rect 216 1096 223 1113
rect 16 856 43 863
rect 76 856 83 873
rect 16 807 23 856
rect 56 823 63 843
rect 36 816 63 823
rect 36 643 43 816
rect 96 803 103 1073
rect 196 1067 203 1096
rect 236 1076 243 1133
rect 256 1127 263 1313
rect 296 1303 303 1336
rect 276 1296 303 1303
rect 276 1227 283 1296
rect 316 1287 323 1356
rect 376 1336 383 1433
rect 396 1347 403 1373
rect 416 1347 423 1413
rect 436 1407 443 1553
rect 456 1467 463 1693
rect 476 1596 483 1613
rect 476 1367 483 1493
rect 496 1343 503 1633
rect 536 1627 543 1753
rect 656 1747 663 1783
rect 576 1616 583 1633
rect 516 1596 543 1603
rect 536 1563 543 1596
rect 476 1336 503 1343
rect 516 1556 543 1563
rect 476 1323 483 1336
rect 516 1327 523 1556
rect 536 1327 543 1533
rect 556 1527 563 1583
rect 596 1576 603 1633
rect 636 1627 643 1653
rect 636 1576 643 1613
rect 656 1607 663 1713
rect 696 1623 703 1773
rect 716 1647 723 1833
rect 736 1827 743 1993
rect 756 1747 763 2033
rect 776 2007 783 2076
rect 796 2027 803 2093
rect 816 2087 823 2193
rect 836 2076 843 2213
rect 896 2167 903 2283
rect 916 2207 923 2253
rect 936 2227 943 2493
rect 956 2487 963 2513
rect 976 2507 983 2543
rect 1036 2536 1043 2613
rect 1056 2567 1063 2733
rect 1116 2707 1123 2873
rect 1136 2687 1143 2813
rect 1196 2787 1203 2793
rect 1156 2747 1163 2763
rect 1196 2756 1203 2773
rect 1236 2743 1243 2973
rect 1256 2787 1263 2993
rect 1216 2707 1223 2743
rect 1236 2736 1263 2743
rect 1096 2607 1103 2653
rect 1236 2647 1243 2736
rect 1296 2727 1303 2953
rect 1316 2827 1323 3003
rect 1356 2996 1383 3003
rect 956 2307 963 2333
rect 976 2247 983 2433
rect 996 2387 1003 2513
rect 1016 2487 1023 2523
rect 1036 2287 1043 2393
rect 1056 2267 1063 2523
rect 1076 2447 1083 2513
rect 1096 2307 1103 2593
rect 1136 2536 1143 2633
rect 1156 2547 1163 2633
rect 1176 2536 1183 2593
rect 1236 2587 1243 2593
rect 1196 2543 1203 2573
rect 1196 2536 1223 2543
rect 1116 2467 1123 2523
rect 1136 2327 1143 2493
rect 1076 2267 1083 2283
rect 1116 2276 1123 2313
rect 1156 2263 1163 2373
rect 1196 2347 1203 2513
rect 1256 2407 1263 2693
rect 1316 2667 1323 2813
rect 1356 2767 1363 2873
rect 1376 2807 1383 2996
rect 1396 2987 1403 3023
rect 1436 3016 1443 3213
rect 1456 3207 1463 3673
rect 1556 3667 1563 3693
rect 1576 3687 1583 3733
rect 1636 3716 1643 3753
rect 1716 3707 1723 3956
rect 1756 3727 1763 3993
rect 1536 3463 1543 3593
rect 1536 3456 1563 3463
rect 1476 3167 1483 3393
rect 1496 3236 1503 3253
rect 1516 3187 1523 3253
rect 1556 3247 1563 3456
rect 1496 3107 1503 3173
rect 1476 3007 1483 3073
rect 1516 3027 1523 3073
rect 1556 3027 1563 3173
rect 1576 3123 1583 3613
rect 1596 3516 1603 3553
rect 1596 3287 1603 3473
rect 1636 3327 1643 3633
rect 1796 3547 1803 4033
rect 1816 3976 1823 4013
rect 1876 4003 1883 4073
rect 1936 4047 1943 4173
rect 1876 3996 1903 4003
rect 1936 3996 1943 4033
rect 1856 3967 1863 3983
rect 1816 3707 1823 3933
rect 1836 3743 1843 3953
rect 1836 3736 1863 3743
rect 1856 3716 1863 3736
rect 1896 3716 1903 3753
rect 1836 3667 1843 3703
rect 1916 3687 1923 3973
rect 1956 3767 1963 4013
rect 1976 3987 1983 4153
rect 1996 4107 2003 4203
rect 2036 4023 2043 4393
rect 2096 4327 2103 4476
rect 2236 4456 2263 4463
rect 2256 4447 2263 4456
rect 2056 4047 2063 4203
rect 2076 4147 2083 4223
rect 2116 4216 2123 4273
rect 2276 4223 2283 4533
rect 2296 4476 2303 4513
rect 2336 4476 2343 4533
rect 3147 4516 3163 4523
rect 2416 4476 2433 4483
rect 2356 4447 2363 4463
rect 2367 4436 2383 4443
rect 2256 4216 2283 4223
rect 2256 4183 2263 4216
rect 2236 4176 2263 4183
rect 2016 4016 2043 4023
rect 2036 3996 2043 4016
rect 2076 3996 2083 4093
rect 2136 4016 2143 4113
rect 1996 3967 2003 3983
rect 2056 3963 2063 3983
rect 2176 3963 2183 4113
rect 2276 4087 2283 4183
rect 2256 3963 2263 4053
rect 2276 4007 2283 4033
rect 2276 3976 2283 3993
rect 2316 3976 2323 4093
rect 2376 4047 2383 4436
rect 2436 4427 2443 4473
rect 2476 4463 2483 4493
rect 2556 4476 2583 4483
rect 2476 4456 2503 4463
rect 2536 4447 2543 4463
rect 2396 4027 2403 4183
rect 2376 3996 2403 4003
rect 2416 3996 2423 4393
rect 2456 4183 2463 4373
rect 2496 4207 2503 4433
rect 2576 4427 2583 4476
rect 2696 4476 2723 4483
rect 2716 4467 2723 4476
rect 2936 4483 2943 4493
rect 2816 4476 2843 4483
rect 2916 4476 2943 4483
rect 2636 4427 2643 4463
rect 2676 4447 2683 4463
rect 2676 4247 2683 4433
rect 2436 4176 2463 4183
rect 2556 4167 2563 4173
rect 2596 4167 2603 4173
rect 2576 4027 2583 4163
rect 2056 3956 2083 3963
rect 2176 3956 2203 3963
rect 2236 3956 2263 3963
rect 2296 3956 2303 3973
rect 1956 3707 1963 3723
rect 2016 3696 2043 3703
rect 1676 3487 1683 3513
rect 1676 3387 1683 3413
rect 1676 3236 1683 3373
rect 1696 3267 1703 3533
rect 1836 3516 1843 3533
rect 1716 3407 1723 3513
rect 1736 3467 1743 3483
rect 1716 3307 1723 3353
rect 1716 3227 1723 3243
rect 1636 3216 1663 3223
rect 1576 3116 1603 3123
rect 1416 2983 1423 2993
rect 1456 2987 1463 3003
rect 1416 2976 1443 2983
rect 1336 2667 1343 2743
rect 1296 2556 1303 2613
rect 1336 2556 1343 2593
rect 1356 2567 1363 2753
rect 1396 2663 1403 2973
rect 1396 2656 1423 2663
rect 1276 2536 1283 2553
rect 1096 2247 1103 2263
rect 1136 2256 1163 2263
rect 896 2083 903 2093
rect 936 2087 943 2113
rect 956 2087 963 2233
rect 1136 2227 1143 2256
rect 876 2076 903 2083
rect 856 2007 863 2063
rect 896 2056 903 2076
rect 936 2056 943 2073
rect 916 2047 923 2053
rect 776 1783 783 1913
rect 816 1827 823 1853
rect 836 1796 843 1873
rect 856 1847 863 1953
rect 876 1867 883 2033
rect 896 1987 903 2013
rect 896 1796 903 1873
rect 936 1863 943 2013
rect 956 1887 963 2043
rect 976 2007 983 2213
rect 996 2056 1003 2073
rect 1016 2067 1023 2093
rect 1036 2056 1043 2113
rect 1116 2087 1123 2093
rect 1156 2087 1163 2213
rect 1076 2043 1083 2073
rect 1056 2036 1083 2043
rect 1116 2036 1123 2073
rect 996 1987 1003 2013
rect 916 1856 943 1863
rect 916 1827 923 1856
rect 936 1787 943 1803
rect 776 1776 803 1783
rect 676 1616 703 1623
rect 456 1316 483 1323
rect 296 1207 303 1273
rect 336 1187 343 1293
rect 296 1147 303 1173
rect 356 1147 363 1273
rect 376 1187 383 1293
rect 396 1167 403 1303
rect 436 1247 443 1303
rect 456 1227 463 1316
rect 476 1167 483 1293
rect 556 1287 563 1303
rect 376 1143 383 1153
rect 376 1136 403 1143
rect 296 1103 303 1113
rect 296 1096 323 1103
rect 176 863 183 1053
rect 256 867 263 1053
rect 296 887 303 1073
rect 356 1067 363 1103
rect 396 1087 403 1136
rect 416 1127 423 1153
rect 416 1096 423 1113
rect 436 1107 443 1133
rect 436 1076 443 1093
rect 496 1067 503 1273
rect 516 1227 523 1283
rect 576 1247 583 1573
rect 616 1567 623 1573
rect 656 1547 663 1563
rect 596 1287 603 1303
rect 596 1267 603 1273
rect 556 1147 563 1193
rect 576 1116 583 1213
rect 616 1207 623 1273
rect 636 1247 643 1303
rect 656 1187 663 1313
rect 527 1076 533 1083
rect 136 856 163 863
rect 176 856 203 863
rect 96 796 123 803
rect 16 636 43 643
rect 76 636 103 643
rect 116 636 123 796
rect 136 667 143 813
rect 156 807 163 856
rect 196 827 203 856
rect 176 787 183 823
rect 216 707 223 843
rect 296 823 303 873
rect 376 836 383 853
rect 156 656 163 673
rect 16 376 23 636
rect 96 407 103 636
rect 56 376 83 383
rect 96 376 103 393
rect 156 387 163 613
rect 176 607 183 623
rect 196 403 203 613
rect 216 607 223 623
rect 236 427 243 633
rect 176 396 203 403
rect 136 376 153 383
rect 36 207 43 363
rect 76 327 83 376
rect 36 163 43 193
rect 36 156 63 163
rect 56 136 63 156
rect 76 147 83 173
rect 96 167 103 333
rect 116 187 123 363
rect 176 347 183 396
rect 236 376 243 393
rect 256 367 263 693
rect 276 667 283 823
rect 296 816 323 823
rect 296 787 303 816
rect 396 723 403 813
rect 376 716 403 723
rect 316 656 323 673
rect 356 647 363 673
rect 376 667 383 716
rect 416 707 423 873
rect 436 807 443 823
rect 296 607 303 623
rect 356 616 363 633
rect 396 627 403 693
rect 276 376 283 573
rect 316 527 323 613
rect 316 376 323 453
rect 296 347 303 363
rect 256 327 263 333
rect 136 176 143 193
rect 96 136 103 153
rect 236 136 243 193
rect 316 187 323 333
rect 336 187 343 413
rect 356 387 363 493
rect 396 367 403 433
rect 416 407 423 603
rect 436 507 443 673
rect 456 667 463 853
rect 496 847 503 893
rect 516 836 523 913
rect 476 747 483 823
rect 536 747 543 1053
rect 556 763 563 1033
rect 576 907 583 1073
rect 576 836 583 853
rect 596 847 603 1173
rect 616 823 623 1173
rect 656 1096 663 1153
rect 676 1123 683 1616
rect 756 1596 763 1693
rect 696 1507 703 1553
rect 716 1387 723 1573
rect 736 1527 743 1583
rect 736 1347 743 1453
rect 696 1267 703 1303
rect 756 1287 763 1323
rect 716 1227 723 1273
rect 676 1116 703 1123
rect 716 1116 723 1193
rect 736 1127 743 1173
rect 776 1143 783 1633
rect 796 1607 803 1776
rect 816 1727 823 1753
rect 856 1727 863 1753
rect 816 1587 823 1613
rect 876 1607 883 1753
rect 916 1747 923 1783
rect 936 1707 943 1773
rect 956 1747 963 1853
rect 1016 1847 1023 1893
rect 1036 1867 1043 2013
rect 1036 1847 1043 1853
rect 1056 1827 1063 2013
rect 1076 1803 1083 1993
rect 1096 1847 1103 2013
rect 1176 2007 1183 2253
rect 1196 2247 1203 2263
rect 1256 2227 1263 2293
rect 1276 2067 1283 2493
rect 1316 2347 1323 2543
rect 1376 2536 1383 2573
rect 1356 2487 1363 2523
rect 1396 2507 1403 2523
rect 1416 2507 1423 2656
rect 1436 2587 1443 2976
rect 1496 2927 1503 3003
rect 1536 2987 1543 3003
rect 1456 2767 1463 2913
rect 1556 2867 1563 2993
rect 1456 2587 1463 2753
rect 1556 2743 1563 2853
rect 1576 2847 1583 2973
rect 1596 2967 1603 3116
rect 1616 3047 1623 3153
rect 1456 2556 1463 2573
rect 1476 2567 1483 2673
rect 1496 2607 1503 2743
rect 1536 2736 1563 2743
rect 1496 2543 1503 2573
rect 1476 2536 1503 2543
rect 1316 2183 1323 2313
rect 1336 2247 1343 2263
rect 1296 2176 1323 2183
rect 1296 2107 1303 2176
rect 1316 2096 1323 2133
rect 1016 1787 1023 1803
rect 1056 1796 1083 1803
rect 1096 1796 1103 1813
rect 1036 1747 1043 1773
rect 916 1627 923 1633
rect 956 1596 963 1613
rect 876 1543 883 1573
rect 896 1567 903 1583
rect 856 1536 883 1543
rect 796 1347 803 1493
rect 796 1227 803 1293
rect 816 1287 823 1413
rect 836 1367 843 1473
rect 856 1467 863 1536
rect 896 1527 903 1553
rect 916 1507 923 1573
rect 756 1136 783 1143
rect 636 1027 643 1083
rect 696 887 703 1116
rect 756 927 763 1136
rect 776 1027 783 1073
rect 776 856 783 993
rect 656 836 663 853
rect 696 847 703 853
rect 716 836 743 843
rect 616 816 643 823
rect 596 767 603 803
rect 556 756 583 763
rect 436 407 443 473
rect 456 407 463 653
rect 536 636 543 713
rect 516 603 523 623
rect 516 596 543 603
rect 476 403 483 513
rect 496 487 503 593
rect 536 587 543 596
rect 516 507 523 573
rect 556 567 563 733
rect 576 663 583 756
rect 616 667 623 693
rect 576 656 603 663
rect 476 396 503 403
rect 356 327 363 343
rect 436 327 443 393
rect 456 387 463 393
rect 496 387 503 396
rect 476 327 483 363
rect 516 327 523 453
rect 596 427 603 656
rect 616 636 623 653
rect 636 647 643 793
rect 656 616 663 753
rect 676 687 683 793
rect 696 663 703 773
rect 676 656 703 663
rect 676 636 683 656
rect 716 647 723 793
rect 736 767 743 836
rect 756 827 763 843
rect 536 376 543 413
rect 356 287 363 313
rect 476 307 483 313
rect 256 156 263 173
rect 356 156 363 253
rect 376 136 383 153
rect 76 116 83 133
rect 416 123 423 233
rect 436 187 443 293
rect 556 267 563 363
rect 576 343 583 383
rect 576 336 603 343
rect 416 116 443 123
rect 476 116 483 173
rect 496 136 503 153
rect 536 116 543 173
rect 556 147 563 193
rect 596 187 603 336
rect 616 207 623 493
rect 636 447 643 613
rect 696 547 703 623
rect 656 356 663 393
rect 696 356 703 393
rect 636 327 643 343
rect 676 227 683 343
rect 696 203 703 313
rect 736 247 743 753
rect 776 663 783 733
rect 796 687 803 1193
rect 816 1127 823 1273
rect 836 1167 843 1293
rect 856 1287 863 1303
rect 876 1263 883 1453
rect 936 1427 943 1573
rect 856 1256 883 1263
rect 856 1247 863 1256
rect 836 1096 843 1133
rect 856 1127 863 1213
rect 876 1096 883 1233
rect 896 1227 903 1353
rect 956 1336 963 1373
rect 976 1367 983 1673
rect 996 1576 1003 1633
rect 1016 1607 1023 1733
rect 1056 1603 1063 1796
rect 1116 1763 1123 1993
rect 1147 1856 1153 1863
rect 1196 1816 1203 2053
rect 1136 1796 1163 1803
rect 1156 1787 1163 1796
rect 1096 1756 1123 1763
rect 1076 1627 1083 1753
rect 1056 1596 1083 1603
rect 1027 1576 1043 1583
rect 1076 1543 1083 1596
rect 1096 1567 1103 1756
rect 1136 1667 1143 1773
rect 1176 1747 1183 1803
rect 1116 1587 1123 1633
rect 1136 1596 1143 1653
rect 1196 1576 1203 1593
rect 1216 1587 1223 2053
rect 1236 1847 1243 2063
rect 1276 1847 1283 2033
rect 1296 1847 1303 2013
rect 1236 1767 1243 1803
rect 1256 1727 1263 1813
rect 1276 1747 1283 1803
rect 1256 1647 1263 1673
rect 1276 1567 1283 1693
rect 1296 1687 1303 1773
rect 1316 1707 1323 2053
rect 1356 2043 1363 2333
rect 1416 2267 1423 2473
rect 1436 2427 1443 2533
rect 1476 2367 1483 2536
rect 1376 2207 1383 2263
rect 1416 2107 1423 2253
rect 1476 2223 1483 2333
rect 1496 2283 1503 2373
rect 1576 2347 1583 2833
rect 1616 2827 1623 2953
rect 1636 2787 1643 3216
rect 1716 3207 1723 3213
rect 1656 3036 1663 3093
rect 1696 3036 1703 3153
rect 1736 3147 1743 3353
rect 1636 2707 1643 2743
rect 1656 2667 1663 2973
rect 1676 2887 1683 3023
rect 1716 3016 1723 3073
rect 1696 2927 1703 2993
rect 1736 2983 1743 3113
rect 1756 3107 1763 3453
rect 1776 3407 1783 3483
rect 1816 3467 1823 3503
rect 1796 3303 1803 3373
rect 1787 3296 1803 3303
rect 1776 3167 1783 3243
rect 1816 3236 1823 3273
rect 1836 3267 1843 3293
rect 1856 3256 1863 3433
rect 1876 3423 1883 3673
rect 1916 3516 1923 3633
rect 1896 3487 1903 3503
rect 1896 3447 1903 3473
rect 1876 3416 1903 3423
rect 1896 3287 1903 3416
rect 1876 3227 1883 3243
rect 1876 3207 1883 3213
rect 1796 3036 1803 3153
rect 1816 3047 1823 3133
rect 1836 3007 1843 3193
rect 1896 3123 1903 3213
rect 1916 3147 1923 3473
rect 1936 3367 1943 3613
rect 1956 3487 1963 3673
rect 1996 3507 2003 3593
rect 2036 3523 2043 3696
rect 2076 3683 2083 3956
rect 2336 3763 2343 3963
rect 2316 3756 2343 3763
rect 2096 3696 2123 3703
rect 2076 3676 2103 3683
rect 2036 3516 2063 3523
rect 2036 3483 2043 3516
rect 2016 3476 2043 3483
rect 1956 3236 1963 3273
rect 1976 3267 1983 3373
rect 1896 3116 1923 3123
rect 1856 3036 1863 3093
rect 1876 3056 1883 3093
rect 1716 2976 1743 2983
rect 1696 2827 1703 2893
rect 1696 2743 1703 2813
rect 1676 2736 1703 2743
rect 1696 2687 1703 2736
rect 1596 2527 1603 2593
rect 1656 2556 1663 2613
rect 1496 2276 1523 2283
rect 1536 2227 1543 2263
rect 1576 2247 1583 2253
rect 1456 2216 1483 2223
rect 1436 2083 1443 2093
rect 1416 2076 1443 2083
rect 1376 2067 1383 2073
rect 1416 2056 1423 2076
rect 1356 2036 1383 2043
rect 1356 1987 1363 2013
rect 1376 1803 1383 2036
rect 1396 2027 1403 2043
rect 1456 1927 1463 2216
rect 1556 2056 1563 2073
rect 1476 2027 1483 2043
rect 1516 2007 1523 2043
rect 1576 2007 1583 2043
rect 1336 1796 1383 1803
rect 1336 1627 1343 1796
rect 1376 1727 1383 1763
rect 1356 1596 1363 1653
rect 1296 1576 1323 1583
rect 1056 1536 1083 1543
rect 996 1507 1003 1533
rect 1036 1447 1043 1533
rect 916 1287 923 1293
rect 996 1287 1003 1323
rect 816 1027 823 1083
rect 856 1076 863 1093
rect 896 1067 903 1153
rect 916 1096 923 1273
rect 996 1207 1003 1253
rect 976 1116 983 1153
rect 996 1116 1003 1193
rect 1036 1187 1043 1333
rect 1056 1267 1063 1536
rect 1096 1367 1103 1533
rect 1036 1116 1043 1133
rect 1056 1123 1063 1193
rect 1096 1167 1103 1293
rect 1056 1116 1083 1123
rect 956 1087 963 1103
rect 816 707 823 913
rect 836 867 843 973
rect 856 856 863 893
rect 776 656 803 663
rect 756 636 783 643
rect 796 636 803 656
rect 776 607 783 636
rect 776 367 783 533
rect 836 403 843 653
rect 856 647 863 813
rect 876 787 883 1053
rect 896 987 903 1033
rect 896 867 903 933
rect 916 856 923 893
rect 936 807 943 843
rect 976 827 983 853
rect 996 727 1003 953
rect 1016 927 1023 1103
rect 1076 967 1083 1116
rect 1076 887 1083 933
rect 1096 867 1103 1153
rect 1116 1147 1123 1313
rect 1136 1207 1143 1323
rect 1156 1307 1163 1553
rect 1176 1447 1183 1553
rect 1256 1547 1263 1563
rect 1196 1487 1203 1533
rect 1236 1507 1243 1533
rect 1296 1527 1303 1553
rect 1316 1507 1323 1576
rect 1176 1316 1183 1333
rect 1196 1327 1203 1373
rect 1196 1247 1203 1283
rect 1196 1227 1203 1233
rect 1216 1187 1223 1353
rect 1256 1336 1263 1393
rect 1136 1116 1143 1153
rect 1176 1116 1183 1173
rect 1116 1096 1123 1113
rect 1156 1087 1163 1103
rect 1156 987 1163 1073
rect 1116 867 1123 913
rect 1036 767 1043 843
rect 876 636 883 653
rect 896 627 903 693
rect 916 636 923 673
rect 956 636 963 693
rect 856 407 863 593
rect 876 467 883 593
rect 896 587 903 613
rect 876 443 883 453
rect 876 436 903 443
rect 816 396 843 403
rect 816 347 823 396
rect 876 376 883 413
rect 896 387 903 436
rect 936 376 943 393
rect 756 307 763 343
rect 796 327 803 343
rect 776 203 783 323
rect 816 227 823 293
rect 856 227 863 363
rect 916 327 923 363
rect 916 267 923 313
rect 956 287 963 353
rect 896 227 903 233
rect 676 196 703 203
rect 756 196 803 203
rect 676 156 683 196
rect 756 187 763 196
rect 796 187 803 196
rect 816 176 823 213
rect 596 127 603 153
rect 576 103 583 123
rect 616 107 623 143
rect 656 127 663 143
rect 836 107 843 133
rect 576 96 593 103
rect 856 47 863 193
rect 876 127 883 153
rect 896 136 903 213
rect 976 207 983 433
rect 996 427 1003 653
rect 1016 647 1023 673
rect 1056 667 1063 833
rect 1076 787 1083 843
rect 1116 836 1123 853
rect 1176 843 1183 953
rect 1196 947 1203 1153
rect 1236 1147 1243 1303
rect 1256 1267 1263 1293
rect 1256 967 1263 1083
rect 1196 847 1203 913
rect 1216 887 1223 893
rect 1276 887 1283 1333
rect 1336 1327 1343 1553
rect 1376 1367 1383 1613
rect 1396 1407 1403 1913
rect 1436 1827 1443 1873
rect 1576 1816 1583 1993
rect 1436 1796 1443 1813
rect 1516 1787 1523 1803
rect 1456 1747 1463 1783
rect 1496 1767 1503 1783
rect 1536 1647 1543 1793
rect 1436 1616 1463 1623
rect 1456 1583 1463 1616
rect 1436 1576 1463 1583
rect 1416 1487 1423 1553
rect 1436 1507 1443 1576
rect 1476 1556 1483 1633
rect 1576 1616 1583 1633
rect 1596 1627 1603 2493
rect 1636 2387 1643 2533
rect 1616 1827 1623 2273
rect 1656 2267 1663 2513
rect 1676 2487 1683 2633
rect 1696 2567 1703 2673
rect 1716 2483 1723 2976
rect 1796 2947 1803 2993
rect 1756 2807 1763 2873
rect 1776 2687 1783 2793
rect 1836 2787 1843 2973
rect 1796 2607 1803 2743
rect 1856 2707 1863 2733
rect 1696 2476 1723 2483
rect 1676 2227 1683 2263
rect 1696 2187 1703 2476
rect 1736 2263 1743 2553
rect 1776 2427 1783 2563
rect 1836 2536 1843 2653
rect 1816 2507 1823 2513
rect 1856 2487 1863 2523
rect 1876 2483 1883 3013
rect 1916 2847 1923 3116
rect 1936 3067 1943 3193
rect 1976 3147 1983 3223
rect 1996 3187 2003 3243
rect 2016 3163 2023 3453
rect 2036 3243 2043 3273
rect 2076 3267 2083 3483
rect 2096 3467 2103 3676
rect 2116 3547 2123 3696
rect 2156 3607 2163 3733
rect 2316 3727 2323 3756
rect 2176 3716 2203 3723
rect 2176 3587 2183 3716
rect 2336 3716 2343 3733
rect 2176 3567 2183 3573
rect 2156 3496 2163 3513
rect 2196 3496 2223 3503
rect 2196 3483 2203 3496
rect 2036 3236 2063 3243
rect 2096 3236 2103 3413
rect 2116 3267 2123 3473
rect 2136 3463 2143 3483
rect 2176 3476 2203 3483
rect 2236 3476 2243 3513
rect 2136 3456 2163 3463
rect 2156 3347 2163 3456
rect 2136 3247 2143 3313
rect 2156 3247 2163 3333
rect 1996 3156 2023 3163
rect 1956 3056 1963 3113
rect 1996 3036 2003 3156
rect 2036 3143 2043 3213
rect 2016 3136 2043 3143
rect 1896 2767 1903 2793
rect 1936 2787 1943 3023
rect 1976 3007 1983 3023
rect 2016 2967 2023 3136
rect 2036 3056 2043 3093
rect 2076 3027 2083 3193
rect 2096 3036 2103 3073
rect 2116 3067 2123 3213
rect 2136 3087 2143 3203
rect 2156 3027 2163 3113
rect 2176 3107 2183 3476
rect 2276 3307 2283 3483
rect 2276 3227 2283 3273
rect 2296 3267 2303 3553
rect 2316 3536 2323 3593
rect 2356 3367 2363 3993
rect 2376 3707 2383 3913
rect 2396 3683 2403 3996
rect 2376 3676 2403 3683
rect 2376 3627 2383 3676
rect 2396 3543 2403 3653
rect 2436 3567 2443 4013
rect 2476 3907 2483 3983
rect 2476 3747 2483 3893
rect 2616 3707 2623 3973
rect 2676 3967 2683 4233
rect 2716 4087 2723 4183
rect 2756 4127 2763 4183
rect 2816 4087 2823 4476
rect 3016 4427 3023 4513
rect 3056 4476 3063 4513
rect 3096 4476 3103 4513
rect 3156 4496 3163 4516
rect 3176 4507 3183 4513
rect 3116 4467 3123 4493
rect 3136 4476 3143 4493
rect 3176 4476 3183 4493
rect 3236 4476 3243 4513
rect 3336 4496 3343 4533
rect 3296 4476 3323 4483
rect 3296 4467 3303 4476
rect 3196 4456 3223 4463
rect 2916 4147 2923 4213
rect 2996 4147 3003 4183
rect 2736 3996 2743 4033
rect 2876 4016 2903 4023
rect 2876 4003 2883 4016
rect 2956 4003 2963 4133
rect 3036 4127 3043 4183
rect 3076 4167 3083 4433
rect 3116 4267 3123 4433
rect 3196 4427 3203 4456
rect 3376 4463 3383 4473
rect 3376 4456 3393 4463
rect 3136 4216 3163 4223
rect 3196 4216 3203 4273
rect 2856 3996 2883 4003
rect 2936 3996 2963 4003
rect 2996 3996 3003 4033
rect 3056 3996 3063 4013
rect 3096 4007 3103 4153
rect 3156 4127 3163 4216
rect 3216 4187 3223 4203
rect 3256 4167 3263 4253
rect 3276 4216 3283 4233
rect 3336 4167 3343 4183
rect 3376 4167 3383 4183
rect 3356 4067 3363 4163
rect 2716 3716 2743 3723
rect 2716 3707 2723 3716
rect 2456 3687 2463 3703
rect 2576 3696 2603 3703
rect 2396 3536 2423 3543
rect 2336 3247 2343 3293
rect 2356 3256 2363 3273
rect 2396 3256 2403 3293
rect 2296 3236 2323 3243
rect 2216 3056 2263 3063
rect 1916 2756 1933 2763
rect 1976 2756 1983 2773
rect 2016 2756 2023 2793
rect 1936 2743 1943 2753
rect 1936 2736 1963 2743
rect 1916 2536 1923 2673
rect 1936 2567 1943 2713
rect 1896 2507 1903 2523
rect 1876 2476 1903 2483
rect 1796 2267 1803 2473
rect 1716 2256 1743 2263
rect 1716 2207 1723 2256
rect 1816 2207 1823 2453
rect 1836 2276 1863 2283
rect 1836 2247 1843 2276
rect 1876 2227 1883 2243
rect 1636 2067 1643 2173
rect 1656 2076 1663 2113
rect 1696 2087 1703 2153
rect 1756 2107 1763 2133
rect 1776 2076 1783 2173
rect 1816 2076 1823 2153
rect 1836 2096 1843 2153
rect 1856 2076 1863 2093
rect 1616 1687 1623 1763
rect 1296 1147 1303 1293
rect 1316 1287 1323 1303
rect 1316 1067 1323 1083
rect 1216 856 1223 873
rect 1256 847 1263 863
rect 1296 847 1303 1013
rect 1156 836 1183 843
rect 1096 807 1103 813
rect 1036 616 1043 653
rect 1096 647 1103 793
rect 1136 767 1143 823
rect 1236 747 1243 843
rect 1276 767 1283 843
rect 1316 836 1323 913
rect 1336 867 1343 1253
rect 1356 1207 1363 1303
rect 1376 1267 1383 1323
rect 1396 1243 1403 1353
rect 1376 1236 1403 1243
rect 1356 1116 1363 1133
rect 1376 1127 1383 1236
rect 1396 1096 1403 1213
rect 1416 1127 1423 1393
rect 1436 1387 1443 1413
rect 1456 1347 1463 1493
rect 1476 1316 1483 1373
rect 1496 1367 1503 1473
rect 1516 1347 1523 1433
rect 1536 1427 1543 1613
rect 1636 1583 1643 1753
rect 1656 1747 1663 1973
rect 1716 1907 1723 2053
rect 1736 2027 1743 2053
rect 1876 2007 1883 2153
rect 1896 2127 1903 2476
rect 1936 2427 1943 2523
rect 1956 2487 1963 2693
rect 2036 2687 2043 2743
rect 2056 2707 2063 2793
rect 2076 2647 2083 2993
rect 2216 2787 2223 3013
rect 2256 2847 2263 3056
rect 2096 2727 2103 2743
rect 2156 2743 2163 2753
rect 2236 2743 2243 2793
rect 2276 2767 2283 3073
rect 2296 3047 2303 3236
rect 2376 3147 2383 3243
rect 2356 3047 2363 3093
rect 2396 3036 2403 3213
rect 2416 3043 2423 3536
rect 2436 3523 2443 3533
rect 2436 3516 2463 3523
rect 2436 3067 2443 3516
rect 2456 3087 2463 3173
rect 2456 3056 2463 3073
rect 2416 3036 2443 3043
rect 2396 2983 2403 2993
rect 2396 2976 2423 2983
rect 2156 2736 2183 2743
rect 2216 2736 2243 2743
rect 2256 2727 2263 2743
rect 2116 2687 2123 2723
rect 2276 2707 2283 2723
rect 2296 2687 2303 2743
rect 2096 2576 2103 2673
rect 2196 2576 2203 2633
rect 1976 2536 1983 2573
rect 2076 2556 2083 2573
rect 2036 2507 2043 2523
rect 1976 2287 1983 2293
rect 2036 2263 2043 2473
rect 1956 2243 1963 2263
rect 1996 2256 2043 2263
rect 1916 2127 1923 2233
rect 1936 2207 1943 2243
rect 1956 2236 1983 2243
rect 1936 2167 1943 2193
rect 1916 2087 1923 2113
rect 1956 2107 1963 2213
rect 1976 2127 1983 2236
rect 1936 2076 1943 2093
rect 1976 2076 1983 2113
rect 1996 2076 2003 2173
rect 2056 2147 2063 2513
rect 2096 2467 2103 2533
rect 2136 2523 2143 2573
rect 2216 2556 2243 2563
rect 2276 2556 2283 2653
rect 2216 2547 2223 2556
rect 2116 2516 2143 2523
rect 1896 2056 1923 2063
rect 1896 2027 1903 2056
rect 2056 2063 2063 2113
rect 2076 2083 2083 2293
rect 2116 2227 2123 2516
rect 2076 2076 2103 2083
rect 2096 2067 2103 2076
rect 2136 2076 2143 2263
rect 2156 2147 2163 2413
rect 2176 2203 2183 2263
rect 2196 2227 2203 2533
rect 2256 2287 2263 2353
rect 2176 2196 2203 2203
rect 2176 2076 2183 2173
rect 1896 1983 1903 2013
rect 1876 1976 1903 1983
rect 1676 1627 1683 1813
rect 1716 1807 1723 1833
rect 1756 1816 1763 1893
rect 1876 1823 1883 1976
rect 1856 1816 1883 1823
rect 1696 1707 1703 1783
rect 1556 1467 1563 1573
rect 1556 1336 1563 1393
rect 1436 1223 1443 1293
rect 1496 1287 1503 1303
rect 1536 1267 1543 1313
rect 1436 1216 1463 1223
rect 1356 927 1363 1073
rect 1376 887 1383 1073
rect 1396 907 1403 1053
rect 1436 987 1443 1113
rect 1456 1087 1463 1216
rect 1376 836 1383 853
rect 1296 787 1303 803
rect 1336 723 1343 833
rect 1356 807 1363 823
rect 1396 767 1403 823
rect 1336 716 1363 723
rect 1116 627 1123 673
rect 1196 656 1203 693
rect 1236 636 1243 713
rect 1016 583 1023 613
rect 1076 607 1083 613
rect 1016 576 1043 583
rect 996 376 1003 413
rect 1036 383 1043 576
rect 1156 547 1163 623
rect 1036 376 1063 383
rect 1076 376 1083 493
rect 1116 387 1123 533
rect 1056 327 1063 376
rect 1136 367 1143 413
rect 956 156 963 193
rect 996 187 1003 313
rect 1016 176 1023 213
rect 1036 207 1043 293
rect 1096 227 1103 363
rect 1176 356 1183 393
rect 1216 356 1223 493
rect 1256 387 1263 613
rect 1276 447 1283 673
rect 1316 656 1323 693
rect 1336 636 1343 693
rect 1356 687 1363 716
rect 1416 647 1423 753
rect 1436 747 1443 913
rect 1436 636 1443 673
rect 1456 667 1463 893
rect 1476 867 1483 1073
rect 1496 987 1503 1093
rect 1516 1083 1523 1153
rect 1556 1127 1563 1253
rect 1576 1247 1583 1573
rect 1596 1507 1603 1583
rect 1636 1576 1663 1583
rect 1636 1567 1643 1576
rect 1676 1556 1683 1573
rect 1736 1563 1743 1773
rect 1776 1767 1783 1803
rect 1796 1763 1803 1793
rect 1816 1787 1823 1803
rect 1856 1787 1863 1816
rect 1836 1767 1843 1783
rect 1916 1783 1923 1973
rect 1936 1827 1943 2033
rect 1896 1776 1923 1783
rect 1796 1756 1823 1763
rect 1776 1743 1783 1753
rect 1776 1736 1803 1743
rect 1796 1596 1803 1736
rect 1816 1607 1823 1756
rect 1836 1627 1843 1713
rect 1836 1583 1843 1593
rect 1716 1556 1743 1563
rect 1616 1327 1623 1513
rect 1576 1147 1583 1173
rect 1516 1076 1543 1083
rect 1536 1007 1543 1076
rect 1576 1047 1583 1083
rect 1536 883 1543 933
rect 1596 887 1603 1293
rect 1616 1147 1623 1193
rect 1636 1187 1643 1303
rect 1656 1287 1663 1323
rect 1676 1147 1683 1353
rect 1696 1336 1703 1473
rect 1736 1336 1743 1393
rect 1756 1347 1763 1553
rect 1776 1547 1783 1583
rect 1816 1576 1843 1583
rect 1796 1487 1803 1553
rect 1836 1407 1843 1553
rect 1856 1547 1863 1653
rect 1936 1627 1943 1813
rect 1956 1616 1963 1633
rect 1896 1567 1903 1583
rect 1696 1267 1703 1293
rect 1716 1287 1723 1323
rect 1696 1147 1703 1153
rect 1636 1096 1643 1133
rect 1676 1096 1683 1113
rect 1696 1076 1703 1133
rect 1616 1067 1623 1073
rect 1616 947 1623 1033
rect 1516 876 1543 883
rect 1516 856 1523 876
rect 1567 876 1573 883
rect 1496 787 1503 843
rect 1596 827 1603 853
rect 1476 636 1483 733
rect 1356 527 1363 623
rect 1396 616 1423 623
rect 1356 427 1363 433
rect 1376 427 1383 593
rect 1416 587 1423 616
rect 1456 607 1463 623
rect 1496 616 1503 693
rect 1516 547 1523 653
rect 1496 523 1503 533
rect 1536 527 1543 673
rect 1556 636 1563 813
rect 1616 767 1623 913
rect 1636 907 1643 1013
rect 1656 1007 1663 1073
rect 1756 1047 1763 1113
rect 1656 907 1663 933
rect 1636 827 1643 843
rect 1656 707 1663 823
rect 1696 727 1703 823
rect 1716 807 1723 813
rect 1716 703 1723 773
rect 1736 767 1743 873
rect 1756 867 1763 973
rect 1776 947 1783 1193
rect 1796 1147 1803 1273
rect 1836 1267 1843 1303
rect 1856 1227 1863 1393
rect 1916 1367 1923 1573
rect 1936 1387 1943 1583
rect 1876 1307 1883 1323
rect 1856 1096 1863 1133
rect 1876 1127 1883 1293
rect 1896 1287 1903 1343
rect 1916 1123 1923 1313
rect 1936 1267 1943 1293
rect 1956 1267 1963 1573
rect 1976 1567 1983 1583
rect 1996 1567 2003 2013
rect 2016 2007 2023 2063
rect 2056 2056 2083 2063
rect 2076 1947 2083 2056
rect 2116 2056 2123 2073
rect 2196 2063 2203 2196
rect 2216 2127 2223 2273
rect 2276 2247 2283 2313
rect 2296 2267 2303 2633
rect 2336 2276 2343 2513
rect 2356 2307 2363 2773
rect 2416 2767 2423 2976
rect 2436 2787 2443 3036
rect 2456 2987 2463 3013
rect 2476 2807 2483 3013
rect 2496 2827 2503 3573
rect 2536 3547 2543 3693
rect 2596 3667 2603 3696
rect 2656 3687 2663 3703
rect 2696 3696 2713 3703
rect 2536 3523 2543 3533
rect 2536 3516 2563 3523
rect 2576 3516 2583 3553
rect 2676 3527 2683 3673
rect 2756 3667 2763 3673
rect 2776 3627 2783 3953
rect 2856 3703 2863 3996
rect 2936 3967 2943 3996
rect 2796 3687 2803 3703
rect 2836 3696 2863 3703
rect 2816 3647 2823 3683
rect 2516 3127 2523 3353
rect 2556 3223 2563 3516
rect 2716 3516 2723 3553
rect 2756 3516 2783 3523
rect 2536 3216 2563 3223
rect 2556 3207 2563 3216
rect 2516 3047 2523 3113
rect 2576 3043 2583 3223
rect 2676 3167 2683 3223
rect 2556 3036 2583 3043
rect 2616 3036 2623 3053
rect 2576 3016 2603 3023
rect 2476 2756 2483 2773
rect 2376 2607 2383 2753
rect 2396 2647 2403 2743
rect 2416 2583 2423 2723
rect 2456 2707 2463 2723
rect 2416 2576 2443 2583
rect 2436 2563 2443 2576
rect 2496 2583 2503 2793
rect 2536 2723 2543 2993
rect 2596 2987 2603 3016
rect 2636 2807 2643 3133
rect 2696 3047 2703 3493
rect 2756 3427 2763 3516
rect 2836 3483 2843 3513
rect 2836 3476 2863 3483
rect 2716 3187 2723 3223
rect 2716 3107 2723 3173
rect 2756 3067 2763 3413
rect 2676 3003 2683 3033
rect 2676 2996 2703 3003
rect 2596 2743 2603 2773
rect 2696 2763 2703 2996
rect 2776 2867 2783 3153
rect 2676 2756 2703 2763
rect 2596 2736 2623 2743
rect 2516 2716 2543 2723
rect 2516 2667 2523 2716
rect 2496 2576 2523 2583
rect 2436 2556 2463 2563
rect 2516 2347 2523 2576
rect 2536 2556 2543 2693
rect 2556 2507 2563 2733
rect 2656 2727 2663 2743
rect 2716 2727 2723 2743
rect 2796 2707 2803 3053
rect 2836 3007 2843 3213
rect 2856 3207 2863 3223
rect 2856 3107 2863 3193
rect 2896 3167 2903 3223
rect 2856 3036 2863 3073
rect 2816 2776 2823 2793
rect 2876 2727 2883 3093
rect 2896 3036 2903 3093
rect 2916 2787 2923 3613
rect 2936 3527 2943 3953
rect 2976 3727 2983 3973
rect 3176 3947 3183 3963
rect 3156 3727 3163 3753
rect 3216 3743 3223 4013
rect 3236 3996 3243 4033
rect 3316 3996 3323 4013
rect 3216 3736 3243 3743
rect 3036 3716 3063 3723
rect 2956 3687 2963 3703
rect 2956 3667 2963 3673
rect 2976 3623 2983 3683
rect 2996 3647 3003 3703
rect 3016 3623 3023 3683
rect 2976 3616 3023 3623
rect 3056 3607 3063 3716
rect 3076 3716 3103 3723
rect 3076 3687 3083 3716
rect 3116 3667 3123 3683
rect 3136 3647 3143 3703
rect 3176 3587 3183 3703
rect 3196 3687 3203 3723
rect 3216 3567 3223 3713
rect 3236 3547 3243 3736
rect 3276 3727 3283 3733
rect 3296 3727 3303 3983
rect 3336 3727 3343 4013
rect 3356 4007 3363 4053
rect 3376 3716 3383 3953
rect 3396 3747 3403 4233
rect 3436 4167 3443 4533
rect 3496 4247 3503 4513
rect 3516 4476 3543 4483
rect 3516 4183 3523 4476
rect 3616 4187 3623 4213
rect 3516 4176 3543 4183
rect 3536 4087 3543 4176
rect 3556 4023 3563 4093
rect 3536 4016 3563 4023
rect 3476 3996 3483 4013
rect 3296 3627 3303 3683
rect 3356 3667 3363 3683
rect 2956 3487 2963 3523
rect 3036 3516 3043 3533
rect 2956 3247 2963 3473
rect 2976 3127 2983 3213
rect 2976 2987 2983 3043
rect 2996 3007 3003 3453
rect 3096 3247 3103 3273
rect 3136 3267 3143 3513
rect 3156 3327 3163 3533
rect 3216 3516 3223 3533
rect 3176 3487 3183 3513
rect 3236 3467 3243 3493
rect 3276 3307 3283 3553
rect 3356 3536 3363 3553
rect 3336 3516 3343 3533
rect 3376 3523 3383 3673
rect 3396 3647 3403 3703
rect 3416 3627 3423 3993
rect 3576 3947 3583 4003
rect 3636 3927 3643 4493
rect 3656 4476 3683 4483
rect 3656 4447 3663 4476
rect 3656 4167 3663 4233
rect 3716 4216 3723 4233
rect 3696 4107 3703 4203
rect 3736 4167 3743 4183
rect 3656 3996 3663 4073
rect 3676 3967 3683 4033
rect 3756 4027 3763 4163
rect 3776 3907 3783 4153
rect 3456 3716 3483 3723
rect 3396 3547 3403 3553
rect 3436 3547 3443 3613
rect 3376 3516 3403 3523
rect 3396 3507 3403 3516
rect 3296 3487 3303 3503
rect 3296 3283 3303 3393
rect 3276 3276 3303 3283
rect 3036 3047 3043 3193
rect 3076 3187 3083 3223
rect 3096 3207 3103 3233
rect 3116 3227 3123 3243
rect 3216 3236 3223 3273
rect 3176 3207 3183 3223
rect 3076 3047 3083 3173
rect 2596 2556 2623 2563
rect 2636 2556 2643 2673
rect 2156 1947 2163 2063
rect 2196 2056 2223 2063
rect 2076 1783 2083 1813
rect 2016 1627 2023 1783
rect 2056 1776 2083 1783
rect 2036 1607 2043 1633
rect 2096 1607 2103 1933
rect 2196 1867 2203 2056
rect 2236 1987 2243 2153
rect 2156 1647 2163 1833
rect 2196 1827 2203 1853
rect 2256 1807 2263 2213
rect 2276 1847 2283 2093
rect 2176 1627 2183 1793
rect 2196 1623 2203 1773
rect 2236 1763 2243 1783
rect 2236 1756 2283 1763
rect 2196 1616 2223 1623
rect 2156 1596 2163 1613
rect 2276 1603 2283 1756
rect 2296 1727 2303 2133
rect 2336 1827 2343 2053
rect 2356 1847 2363 2063
rect 2376 1987 2383 2233
rect 2396 2107 2403 2293
rect 2496 2243 2503 2283
rect 2536 2247 2543 2273
rect 2576 2267 2583 2493
rect 2616 2327 2623 2556
rect 2696 2547 2703 2593
rect 2656 2507 2663 2543
rect 2716 2507 2723 2693
rect 2796 2576 2823 2583
rect 2796 2567 2803 2576
rect 2836 2556 2843 2573
rect 2736 2523 2743 2553
rect 2856 2527 2863 2573
rect 2736 2516 2763 2523
rect 2876 2507 2883 2543
rect 2636 2296 2643 2353
rect 2616 2263 2623 2293
rect 2596 2256 2623 2263
rect 2456 2236 2503 2243
rect 2456 2043 2463 2193
rect 2496 2076 2503 2236
rect 2396 1947 2403 2043
rect 2436 2036 2463 2043
rect 2516 1967 2523 2043
rect 2316 1763 2323 1783
rect 2316 1756 2343 1763
rect 2276 1596 2303 1603
rect 2016 1576 2023 1593
rect 2096 1567 2103 1593
rect 2136 1576 2143 1593
rect 2076 1543 2083 1563
rect 2116 1547 2123 1573
rect 2176 1567 2183 1583
rect 2336 1567 2343 1756
rect 2356 1747 2363 1783
rect 2076 1536 2093 1543
rect 1996 1347 2003 1533
rect 1976 1287 1983 1303
rect 1916 1116 1943 1123
rect 1796 1067 1803 1083
rect 1836 1067 1843 1083
rect 1936 1067 1943 1116
rect 1976 1096 1983 1273
rect 2016 1247 2023 1303
rect 1756 747 1763 813
rect 1796 807 1803 973
rect 1816 967 1823 1033
rect 1816 827 1823 953
rect 1836 927 1843 1053
rect 1956 1047 1963 1083
rect 1996 1063 2003 1083
rect 1976 1056 2003 1063
rect 1836 836 1843 873
rect 1896 856 1903 1013
rect 1936 887 1943 893
rect 1936 856 1943 873
rect 1976 867 1983 1056
rect 2016 1027 2023 1213
rect 2056 1147 2063 1373
rect 2096 1316 2103 1373
rect 2356 1347 2363 1633
rect 2396 1603 2403 1853
rect 2416 1767 2423 1783
rect 2376 1596 2403 1603
rect 2416 1596 2423 1733
rect 2436 1647 2443 1763
rect 2456 1747 2463 1783
rect 2476 1743 2483 1833
rect 2536 1823 2543 2153
rect 2596 2076 2603 2153
rect 2616 2007 2623 2233
rect 2656 2227 2663 2263
rect 2676 2167 2683 2333
rect 2696 2256 2723 2263
rect 2696 2207 2703 2256
rect 2656 2063 2663 2133
rect 2636 2056 2663 2063
rect 2676 2047 2683 2073
rect 2696 2007 2703 2043
rect 2536 1816 2563 1823
rect 2496 1767 2503 1773
rect 2516 1747 2523 1763
rect 2476 1736 2503 1743
rect 2156 1327 2163 1343
rect 2216 1336 2243 1343
rect 2136 1287 2143 1323
rect 2036 1116 2063 1123
rect 2096 1116 2103 1253
rect 2136 1127 2143 1233
rect 2036 1067 2043 1116
rect 2156 1107 2163 1293
rect 2216 1247 2223 1336
rect 2256 1307 2263 1323
rect 2376 1316 2383 1533
rect 2436 1363 2443 1613
rect 2416 1356 2443 1363
rect 2296 1276 2323 1283
rect 2216 1127 2223 1133
rect 2076 1087 2083 1103
rect 2216 1076 2223 1113
rect 2236 1096 2263 1103
rect 2296 1096 2303 1276
rect 2256 1067 2263 1096
rect 2336 1083 2343 1103
rect 2316 1076 2343 1083
rect 2316 1067 2323 1076
rect 1856 787 1863 803
rect 1696 696 1723 703
rect 1596 667 1603 673
rect 1696 636 1703 696
rect 1576 607 1583 623
rect 1616 616 1643 623
rect 1496 516 1523 523
rect 1276 356 1283 373
rect 1116 227 1123 313
rect 976 147 983 173
rect 1036 156 1043 193
rect 1076 156 1083 193
rect 1096 167 1103 213
rect 1136 156 1143 293
rect 1176 156 1183 313
rect 1196 287 1203 343
rect 1256 307 1263 333
rect 996 127 1003 143
rect 1096 136 1103 153
rect 1116 123 1123 133
rect 1156 123 1163 143
rect 1116 116 1163 123
rect 976 87 983 113
rect 1216 67 1223 193
rect 1276 136 1283 233
rect 1296 207 1303 343
rect 1336 287 1343 373
rect 1356 367 1363 413
rect 1396 367 1403 453
rect 1456 356 1463 393
rect 1376 267 1383 343
rect 1396 267 1403 323
rect 1416 247 1423 313
rect 1436 287 1443 343
rect 1316 27 1323 173
rect 1336 136 1343 153
rect 1376 136 1383 233
rect 1436 167 1443 173
rect 1456 156 1463 313
rect 1476 267 1483 313
rect 1496 307 1503 363
rect 1516 187 1523 516
rect 1536 367 1543 513
rect 1556 387 1563 513
rect 1576 387 1583 593
rect 1596 527 1603 613
rect 1636 527 1643 616
rect 1676 603 1683 623
rect 1716 607 1723 653
rect 1736 623 1743 673
rect 1736 616 1753 623
rect 1776 616 1783 653
rect 1676 596 1703 603
rect 1556 356 1583 363
rect 1536 287 1543 323
rect 1576 267 1583 356
rect 1596 287 1603 433
rect 1656 407 1663 533
rect 1636 367 1643 393
rect 1676 387 1683 573
rect 1696 527 1703 596
rect 1716 463 1723 473
rect 1696 456 1723 463
rect 1696 427 1703 456
rect 1716 367 1723 413
rect 1736 367 1743 493
rect 1776 487 1783 573
rect 1796 487 1803 603
rect 1816 547 1823 653
rect 1836 636 1843 753
rect 1876 687 1883 853
rect 1916 807 1923 843
rect 1976 836 1983 853
rect 1876 636 1893 643
rect 1836 527 1843 593
rect 1856 587 1863 623
rect 1896 616 1923 623
rect 1896 567 1903 573
rect 1616 207 1623 343
rect 1656 267 1663 323
rect 1676 243 1683 313
rect 1696 307 1703 313
rect 1736 283 1743 333
rect 1756 307 1763 333
rect 1736 276 1763 283
rect 1656 236 1683 243
rect 1436 147 1443 153
rect 1536 147 1543 193
rect 1516 127 1523 143
rect 1396 107 1403 123
rect 1556 116 1563 153
rect 1616 147 1623 193
rect 1636 127 1643 233
rect 1656 156 1663 236
rect 1696 203 1703 233
rect 1676 196 1703 203
rect 1676 187 1683 196
rect 1736 147 1743 173
rect 1756 167 1763 276
rect 1776 267 1783 383
rect 1816 376 1823 393
rect 1796 287 1803 363
rect 1836 347 1843 493
rect 1916 467 1923 616
rect 1856 356 1863 433
rect 1876 367 1883 453
rect 1896 356 1903 413
rect 1916 407 1923 433
rect 1936 403 1943 773
rect 1956 727 1963 793
rect 1996 787 2003 873
rect 2036 856 2043 1053
rect 1976 703 1983 733
rect 1956 696 1983 703
rect 1956 636 1963 696
rect 1996 656 2003 753
rect 2016 667 2023 793
rect 2036 636 2043 713
rect 2056 707 2063 773
rect 2076 636 2083 863
rect 2096 803 2103 843
rect 2096 796 2123 803
rect 2096 627 2103 693
rect 2116 667 2123 796
rect 1976 607 1983 623
rect 1996 487 2003 613
rect 2016 563 2023 623
rect 2016 556 2043 563
rect 2036 547 2043 556
rect 1936 396 1953 403
rect 1956 376 1963 393
rect 2016 387 2023 533
rect 2056 527 2063 623
rect 2116 607 2123 633
rect 2036 376 2043 413
rect 2096 407 2103 553
rect 2116 427 2123 573
rect 2136 527 2143 733
rect 2156 687 2163 933
rect 2236 807 2243 843
rect 2276 827 2283 1053
rect 2416 887 2423 1356
rect 2476 1347 2483 1673
rect 2496 1507 2503 1736
rect 2536 1607 2543 1773
rect 2556 1687 2563 1816
rect 2656 1783 2663 1973
rect 2576 1767 2583 1783
rect 2616 1776 2663 1783
rect 2676 1823 2683 1953
rect 2736 1847 2743 2033
rect 2676 1816 2703 1823
rect 2556 1596 2563 1653
rect 2676 1647 2683 1816
rect 2716 1783 2723 1803
rect 2707 1776 2723 1783
rect 2756 1647 2763 1993
rect 2816 1947 2823 2493
rect 2856 2263 2863 2273
rect 2836 2256 2863 2263
rect 2896 2187 2903 2573
rect 2916 2567 2923 2773
rect 2956 2563 2963 2833
rect 2996 2647 3003 2853
rect 3016 2727 3023 2743
rect 3036 2687 3043 2993
rect 2956 2556 2983 2563
rect 2996 2556 3003 2633
rect 3036 2556 3043 2573
rect 2956 2507 2963 2523
rect 2976 2427 2983 2556
rect 2916 2167 2923 2413
rect 3056 2323 3063 2973
rect 3096 2947 3103 3053
rect 3116 3036 3123 3073
rect 3156 3056 3163 3073
rect 3196 3047 3203 3223
rect 3256 3127 3263 3243
rect 3276 3207 3283 3276
rect 3236 3036 3263 3043
rect 3136 3007 3143 3023
rect 3096 2887 3103 2933
rect 3096 2736 3103 2793
rect 3116 2556 3123 2693
rect 3156 2667 3163 3013
rect 3256 2987 3263 3036
rect 3216 2707 3223 2743
rect 3256 2727 3263 2743
rect 3276 2703 3283 3193
rect 3296 3007 3303 3233
rect 3316 3227 3323 3243
rect 3416 3236 3423 3473
rect 3456 3283 3463 3653
rect 3476 3567 3483 3716
rect 3516 3703 3523 3753
rect 3496 3696 3523 3703
rect 3576 3703 3583 3733
rect 3616 3716 3623 3753
rect 3676 3723 3683 3833
rect 3656 3716 3683 3723
rect 3576 3696 3603 3703
rect 3636 3696 3703 3703
rect 3596 3607 3603 3696
rect 3476 3347 3483 3533
rect 3496 3516 3503 3593
rect 3536 3516 3543 3553
rect 3576 3536 3583 3553
rect 3436 3276 3463 3283
rect 3436 3267 3443 3276
rect 3456 3227 3463 3243
rect 3336 3167 3343 3223
rect 3376 3087 3383 3213
rect 3396 3207 3403 3223
rect 3396 3036 3403 3093
rect 3436 3047 3443 3223
rect 3476 3207 3483 3313
rect 3496 3256 3503 3473
rect 3536 3267 3543 3333
rect 3496 3043 3503 3073
rect 3476 3036 3503 3043
rect 3256 2696 3283 2703
rect 3036 2316 3063 2323
rect 2936 2247 2943 2253
rect 2936 2083 2943 2233
rect 2956 2207 2963 2283
rect 2996 2276 3003 2293
rect 3016 2187 3023 2263
rect 2936 2076 2963 2083
rect 2916 1787 2923 2033
rect 2936 1867 2943 2076
rect 2776 1687 2783 1773
rect 2816 1767 2823 1783
rect 2836 1767 2843 1783
rect 2596 1596 2603 1613
rect 2616 1567 2623 1633
rect 2716 1596 2723 1633
rect 2796 1623 2803 1753
rect 2836 1627 2843 1673
rect 2936 1647 2943 1763
rect 2796 1616 2823 1623
rect 2767 1596 2783 1603
rect 2776 1567 2783 1596
rect 2456 1287 2463 1323
rect 2556 1303 2563 1553
rect 2796 1547 2803 1573
rect 2596 1307 2603 1333
rect 2656 1316 2663 1353
rect 2716 1323 2723 1333
rect 2816 1327 2823 1333
rect 2696 1316 2723 1323
rect 2556 1296 2583 1303
rect 2616 1147 2623 1303
rect 2796 1247 2803 1303
rect 2476 1136 2503 1143
rect 2496 967 2503 1136
rect 2636 1116 2643 1173
rect 2676 1116 2683 1153
rect 2696 1147 2703 1193
rect 2696 1116 2703 1133
rect 2856 1116 2863 1173
rect 2876 1167 2883 1573
rect 2896 1567 2903 1593
rect 2896 1116 2903 1153
rect 2656 1087 2663 1093
rect 2356 836 2363 853
rect 2296 807 2303 823
rect 2176 627 2183 793
rect 2196 607 2203 753
rect 2236 647 2243 673
rect 2256 647 2263 773
rect 2276 636 2283 733
rect 2336 687 2343 803
rect 2376 707 2383 803
rect 2316 636 2323 653
rect 2336 636 2343 653
rect 2376 636 2383 673
rect 2216 623 2223 633
rect 2216 616 2263 623
rect 2176 547 2183 573
rect 2136 403 2143 473
rect 2176 407 2183 473
rect 2116 396 2143 403
rect 2116 376 2123 396
rect 2156 376 2183 383
rect 1476 -24 1483 73
rect 1516 67 1523 113
rect 1696 107 1703 133
rect 1716 127 1723 143
rect 1776 136 1783 193
rect 1816 127 1823 333
rect 1856 136 1863 313
rect 1876 267 1883 323
rect 1796 107 1803 123
rect 1836 87 1843 123
rect 1756 -24 1763 53
rect 1876 47 1883 123
rect 1896 -24 1903 113
rect 1916 87 1923 113
rect 1936 47 1943 373
rect 1956 187 1963 293
rect 1976 267 1983 363
rect 2016 327 2023 353
rect 2096 343 2103 373
rect 2096 336 2123 343
rect 2036 307 2043 313
rect 1956 156 1963 173
rect 1936 -24 1943 33
rect 1976 27 1983 153
rect 1996 107 2003 293
rect 2016 167 2023 213
rect 2056 187 2063 333
rect 2076 187 2083 233
rect 2096 207 2103 313
rect 2056 123 2063 173
rect 2076 156 2083 173
rect 2096 156 2103 193
rect 2036 116 2063 123
rect 2056 87 2063 116
rect 2116 67 2123 336
rect 2136 307 2143 353
rect 2176 227 2183 376
rect 2196 367 2203 453
rect 2216 387 2223 553
rect 2236 367 2243 616
rect 2396 616 2403 633
rect 2276 447 2283 593
rect 2296 487 2303 593
rect 2416 507 2423 653
rect 2436 616 2443 753
rect 2456 707 2463 863
rect 2476 687 2483 843
rect 2516 667 2523 973
rect 2556 867 2563 953
rect 2796 867 2803 1113
rect 2916 1067 2923 1533
rect 2976 1367 2983 2173
rect 3036 2127 3043 2316
rect 3056 2267 3063 2283
rect 3096 2276 3103 2353
rect 3156 2307 3163 2653
rect 3156 2276 3163 2293
rect 3196 2267 3203 2283
rect 3116 2207 3123 2263
rect 2996 1627 3003 2113
rect 3116 2103 3123 2193
rect 3136 2187 3143 2263
rect 3216 2227 3223 2673
rect 3236 2556 3243 2593
rect 3256 2467 3263 2696
rect 3296 2627 3303 2993
rect 3336 2736 3363 2743
rect 3356 2587 3363 2736
rect 3336 2556 3343 2573
rect 3376 2556 3383 2953
rect 3396 2756 3403 2993
rect 3436 2727 3443 2933
rect 3496 2783 3503 3013
rect 3516 2803 3523 3243
rect 3556 3223 3563 3473
rect 3596 3327 3603 3503
rect 3636 3323 3643 3633
rect 3656 3547 3663 3573
rect 3676 3516 3683 3553
rect 3696 3487 3703 3673
rect 3756 3547 3763 3723
rect 3776 3687 3783 3893
rect 3796 3687 3803 4413
rect 3816 4207 3823 4443
rect 3836 4176 3843 4193
rect 3876 4187 3883 4463
rect 3956 4387 3963 4533
rect 3936 4183 3943 4213
rect 3936 4176 3963 4183
rect 3876 4087 3883 4173
rect 3916 4147 3923 4173
rect 3856 4016 3863 4033
rect 3936 3996 3943 4033
rect 3976 4023 3983 4513
rect 3996 4463 4003 4616
rect 3996 4456 4023 4463
rect 4016 4167 4023 4456
rect 4036 4407 4043 4553
rect 4056 4427 4063 4573
rect 4076 4476 4083 4623
rect 4116 4587 4123 4623
rect 4136 4507 4143 4573
rect 4156 4567 4163 4623
rect 4196 4547 4203 4623
rect 4236 4587 4243 4623
rect 4256 4616 4283 4623
rect 4196 4496 4223 4503
rect 4096 4476 4113 4483
rect 4096 4447 4103 4476
rect 4156 4456 4163 4493
rect 4096 4307 4103 4433
rect 4136 4307 4143 4443
rect 4196 4407 4203 4496
rect 4036 4107 4043 4293
rect 4196 4247 4203 4393
rect 4136 4183 4143 4213
rect 4216 4196 4223 4233
rect 4096 4067 4103 4183
rect 4136 4176 4163 4183
rect 4196 4067 4203 4153
rect 4236 4123 4243 4183
rect 4256 4163 4263 4616
rect 4316 4587 4323 4623
rect 4556 4616 4583 4623
rect 4636 4616 4663 4623
rect 4336 4456 4343 4493
rect 4256 4156 4283 4163
rect 4236 4116 4263 4123
rect 3956 4016 3983 4023
rect 3856 3947 3863 3973
rect 3876 3927 3883 3983
rect 3816 3667 3823 3913
rect 3896 3683 3903 3713
rect 3876 3676 3903 3683
rect 3756 3516 3783 3523
rect 3816 3516 3823 3593
rect 3756 3507 3763 3516
rect 3836 3467 3843 3503
rect 3776 3327 3783 3453
rect 3636 3316 3663 3323
rect 3596 3307 3603 3313
rect 3576 3256 3583 3293
rect 3536 3216 3563 3223
rect 3536 3027 3543 3216
rect 3636 3147 3643 3293
rect 3656 3256 3663 3316
rect 3716 3256 3743 3263
rect 3776 3256 3783 3313
rect 3516 2796 3543 2803
rect 3536 2787 3543 2796
rect 3496 2776 3523 2783
rect 3416 2556 3423 2713
rect 3456 2687 3463 2743
rect 3476 2647 3483 2723
rect 3456 2556 3463 2633
rect 3476 2567 3483 2593
rect 3496 2556 3503 2693
rect 3276 2507 3283 2523
rect 3116 2096 3143 2103
rect 3056 2083 3063 2093
rect 3176 2087 3183 2173
rect 3196 2096 3203 2113
rect 3036 2076 3063 2083
rect 3056 1827 3063 2076
rect 3216 2076 3223 2093
rect 3116 2047 3123 2063
rect 3136 2007 3143 2053
rect 3016 1623 3023 1783
rect 3016 1616 3043 1623
rect 3076 1616 3083 1773
rect 3136 1707 3143 1813
rect 3156 1783 3163 1853
rect 3156 1776 3183 1783
rect 3216 1647 3223 1783
rect 3036 1423 3043 1616
rect 3136 1596 3143 1633
rect 3236 1607 3243 2253
rect 3296 2207 3303 2313
rect 3336 2247 3343 2263
rect 3356 2227 3363 2543
rect 3396 2527 3403 2533
rect 3256 2067 3263 2153
rect 3276 2076 3283 2133
rect 3356 2076 3383 2083
rect 3176 1547 3183 1593
rect 3196 1547 3203 1563
rect 3016 1416 3043 1423
rect 2936 1267 2943 1303
rect 2976 1287 2983 1303
rect 2976 1167 2983 1273
rect 2996 1147 3003 1313
rect 2996 1083 3003 1133
rect 3016 1127 3023 1416
rect 3256 1387 3263 1693
rect 3076 1083 3083 1293
rect 3096 1283 3103 1333
rect 3176 1303 3183 1353
rect 3216 1316 3223 1333
rect 3256 1316 3263 1353
rect 3156 1296 3183 1303
rect 3096 1276 3143 1283
rect 3196 1267 3203 1303
rect 3236 1267 3243 1283
rect 3276 1207 3283 1933
rect 3336 1847 3343 2053
rect 3376 2047 3383 2076
rect 3436 2027 3443 2513
rect 3296 1783 3303 1833
rect 3456 1816 3463 1833
rect 3296 1776 3323 1783
rect 3356 1747 3363 1783
rect 3316 1576 3323 1633
rect 3336 1607 3343 1653
rect 3296 1527 3303 1563
rect 3336 1547 3343 1553
rect 3136 1116 3143 1153
rect 3176 1116 3183 1133
rect 3216 1116 3223 1133
rect 2996 1076 3023 1083
rect 3056 1076 3083 1083
rect 3156 1083 3163 1103
rect 3156 1076 3183 1083
rect 2596 847 2603 863
rect 2576 807 2583 833
rect 2596 763 2603 833
rect 2616 827 2623 843
rect 2896 836 2903 853
rect 2616 783 2623 813
rect 2616 776 2643 783
rect 2596 756 2623 763
rect 2456 627 2463 653
rect 2476 627 2483 633
rect 2536 616 2543 713
rect 2576 616 2583 733
rect 2336 387 2343 393
rect 2276 376 2303 383
rect 2276 347 2283 376
rect 2316 347 2323 363
rect 2196 287 2203 333
rect 2216 327 2223 343
rect 2136 156 2143 213
rect 2156 27 2163 193
rect 2176 147 2183 193
rect 2196 147 2203 213
rect 2236 163 2243 323
rect 2256 307 2263 343
rect 2396 307 2403 343
rect 2256 207 2263 273
rect 2256 183 2263 193
rect 2356 187 2363 193
rect 2256 176 2283 183
rect 2236 156 2263 163
rect 2276 156 2283 176
rect 2216 136 2223 153
rect 2196 116 2203 133
rect 2256 127 2263 156
rect 2356 156 2363 173
rect 2396 156 2403 253
rect 2416 207 2423 413
rect 2436 156 2443 333
rect 2456 227 2463 383
rect 2476 347 2483 363
rect 2516 156 2523 613
rect 2616 603 2623 756
rect 2596 596 2623 603
rect 2636 427 2643 776
rect 2876 636 2883 823
rect 2916 636 2923 713
rect 2936 647 2943 853
rect 2996 767 3003 1053
rect 3176 843 3183 1076
rect 3176 836 3203 843
rect 3016 807 3023 823
rect 2656 607 2663 623
rect 2696 616 2703 633
rect 2676 547 2683 613
rect 2536 307 2543 373
rect 2556 356 2563 413
rect 2576 367 2583 393
rect 2596 376 2623 383
rect 2596 323 2603 376
rect 2576 316 2603 323
rect 2556 176 2563 193
rect 2596 167 2603 173
rect 2636 156 2643 353
rect 2656 327 2663 383
rect 2696 356 2703 393
rect 2736 387 2743 533
rect 2756 407 2763 603
rect 2736 356 2743 373
rect 2776 367 2783 633
rect 2856 327 2863 373
rect 2876 347 2883 413
rect 2936 387 2943 633
rect 2236 107 2243 123
rect 2296 87 2303 143
rect 2456 136 2483 143
rect 2476 107 2483 136
rect 2536 127 2543 143
rect 2616 127 2623 143
rect 2656 136 2663 253
rect 2696 176 2703 253
rect 2716 243 2723 313
rect 2956 247 2963 713
rect 3016 643 3023 793
rect 3036 667 3043 803
rect 3076 787 3083 833
rect 3096 807 3103 823
rect 3116 787 3123 803
rect 3136 787 3143 823
rect 3196 787 3203 836
rect 2996 636 3023 643
rect 3036 636 3043 653
rect 3076 636 3083 753
rect 3116 663 3123 773
rect 3216 667 3223 823
rect 3276 667 3283 843
rect 3116 656 3143 663
rect 3056 607 3063 623
rect 2976 307 2983 363
rect 3016 356 3023 373
rect 2716 236 2743 243
rect 2736 87 2743 236
rect 2776 167 2783 193
rect 2996 156 3003 343
rect 3016 183 3023 233
rect 3036 207 3043 343
rect 3056 327 3063 593
rect 3176 587 3183 633
rect 3216 587 3223 623
rect 3236 607 3243 653
rect 3296 647 3303 1373
rect 3336 1147 3343 1533
rect 3356 1527 3363 1613
rect 3376 1607 3383 1773
rect 3396 1596 3403 1613
rect 3416 1567 3423 1583
rect 3356 1247 3363 1303
rect 3376 1223 3383 1513
rect 3456 1507 3463 1753
rect 3476 1727 3483 2553
rect 3516 2527 3523 2776
rect 3556 2756 3563 2773
rect 3536 2667 3543 2743
rect 3536 2367 3543 2613
rect 3576 2563 3583 3133
rect 3636 3047 3643 3093
rect 3676 3067 3683 3243
rect 3716 3107 3723 3256
rect 3756 3227 3763 3243
rect 3836 3223 3843 3433
rect 3876 3407 3883 3676
rect 3916 3587 3923 3703
rect 3956 3547 3963 4016
rect 3976 3996 3993 4003
rect 3976 3967 3983 3996
rect 4036 3996 4043 4053
rect 4076 3963 4083 4053
rect 4096 4047 4103 4053
rect 4136 3963 4143 4053
rect 4156 3996 4163 4013
rect 4216 3987 4223 4093
rect 4076 3956 4103 3963
rect 4116 3956 4143 3963
rect 4056 3703 4063 3833
rect 4116 3703 4123 3956
rect 4236 3867 4243 4093
rect 4256 3747 4263 4116
rect 4276 4087 4283 4156
rect 4296 4107 4303 4433
rect 4356 4227 4363 4573
rect 4396 4407 4403 4483
rect 4476 4476 4503 4483
rect 4316 4143 4323 4193
rect 4336 4167 4343 4183
rect 4356 4143 4363 4163
rect 4316 4136 4363 4143
rect 4376 4127 4383 4173
rect 4416 4127 4423 4183
rect 4496 4147 4503 4476
rect 4336 4027 4343 4073
rect 4396 4016 4423 4023
rect 4416 4003 4423 4016
rect 4336 3996 4363 4003
rect 4416 3996 4443 4003
rect 4516 3996 4523 4133
rect 4556 4103 4563 4233
rect 4536 4096 4563 4103
rect 4276 3976 4283 3993
rect 4356 3983 4363 3996
rect 4356 3976 4383 3983
rect 3996 3696 4023 3703
rect 3916 3496 3923 3533
rect 3896 3467 3903 3483
rect 3936 3467 3943 3483
rect 3956 3287 3963 3513
rect 3976 3287 3983 3523
rect 4016 3467 4023 3696
rect 4036 3567 4043 3703
rect 4056 3696 4083 3703
rect 4116 3696 4143 3703
rect 3816 3167 3823 3223
rect 3836 3216 3863 3223
rect 3716 3087 3723 3093
rect 3776 3056 3783 3073
rect 3596 3036 3623 3043
rect 3616 3027 3623 3036
rect 3596 2747 3603 2773
rect 3556 2556 3583 2563
rect 3576 2507 3583 2556
rect 3536 2276 3543 2353
rect 3556 2307 3563 2493
rect 3576 2263 3583 2353
rect 3616 2287 3623 2633
rect 3636 2327 3643 2873
rect 3656 2787 3663 2993
rect 3676 2867 3683 3033
rect 3716 3007 3723 3033
rect 3676 2743 3683 2853
rect 3676 2736 3703 2743
rect 3676 2367 3683 2593
rect 3656 2287 3663 2313
rect 3556 2256 3583 2263
rect 3496 2076 3503 2233
rect 3496 1767 3503 2013
rect 3516 1827 3523 2213
rect 3576 2187 3583 2256
rect 3596 2247 3603 2253
rect 3536 2087 3543 2113
rect 3516 1776 3523 1813
rect 3476 1547 3483 1593
rect 3396 1287 3403 1303
rect 3396 1247 3403 1273
rect 3356 1216 3383 1223
rect 3336 1116 3343 1133
rect 3356 1083 3363 1216
rect 3376 1187 3383 1193
rect 3376 1123 3383 1173
rect 3376 1116 3403 1123
rect 3416 1107 3423 1493
rect 3456 1123 3463 1213
rect 3436 1116 3463 1123
rect 3356 1076 3383 1083
rect 3376 847 3383 1076
rect 3396 767 3403 853
rect 3256 616 3263 633
rect 3276 596 3283 613
rect 3336 603 3343 753
rect 3316 596 3343 603
rect 3356 387 3363 673
rect 3456 667 3463 1116
rect 3476 827 3483 1153
rect 3496 807 3503 823
rect 3496 727 3503 793
rect 3516 687 3523 1633
rect 3536 1596 3543 1613
rect 3556 1603 3563 1853
rect 3596 1823 3603 2193
rect 3616 2107 3623 2243
rect 3636 2007 3643 2063
rect 3676 2056 3683 2133
rect 3576 1816 3603 1823
rect 3576 1783 3583 1816
rect 3576 1776 3603 1783
rect 3616 1763 3623 1933
rect 3596 1756 3623 1763
rect 3576 1727 3583 1753
rect 3576 1627 3583 1713
rect 3556 1596 3583 1603
rect 3576 1127 3583 1553
rect 3596 1467 3603 1756
rect 3636 1747 3643 1783
rect 3616 1507 3623 1673
rect 3656 1647 3663 1853
rect 3696 1623 3703 2353
rect 3716 2327 3723 2973
rect 3776 2927 3783 3013
rect 3816 2967 3823 3013
rect 3736 2707 3743 2913
rect 3836 2887 3843 3153
rect 3856 3047 3863 3113
rect 3876 3036 3883 3253
rect 3896 3067 3903 3273
rect 3916 3256 3923 3273
rect 3956 3256 3983 3263
rect 3916 3036 3923 3133
rect 3936 3023 3943 3243
rect 3956 3047 3963 3213
rect 3976 3187 3983 3256
rect 4016 3247 4023 3273
rect 4036 3267 4043 3533
rect 4056 3527 4063 3573
rect 4076 3447 4083 3673
rect 4116 3667 4123 3696
rect 4096 3516 4103 3593
rect 3976 3087 3983 3173
rect 3996 3147 4003 3213
rect 4016 3127 4023 3153
rect 3996 3063 4003 3113
rect 4036 3087 4043 3223
rect 4056 3167 4063 3223
rect 4076 3127 4083 3313
rect 4116 3207 4123 3653
rect 4156 3627 4163 3683
rect 4176 3647 4183 3703
rect 4156 3427 4163 3553
rect 4176 3247 4183 3593
rect 4136 3236 4163 3243
rect 3976 3056 4003 3063
rect 3976 3036 3983 3056
rect 4016 3036 4023 3073
rect 4036 3036 4043 3073
rect 3936 3016 3963 3023
rect 4096 3016 4103 3053
rect 4116 3027 4123 3093
rect 4136 3087 4143 3236
rect 4196 3227 4203 3673
rect 4216 3667 4223 3683
rect 4276 3627 4283 3713
rect 4296 3703 4303 3853
rect 4316 3847 4323 3973
rect 4296 3696 4323 3703
rect 4296 3647 4303 3696
rect 4216 3427 4223 3523
rect 4316 3267 4323 3613
rect 4356 3607 4363 3953
rect 4376 3607 4383 3976
rect 4396 3527 4403 3703
rect 4416 3627 4423 3973
rect 4536 3767 4543 4096
rect 4576 3963 4583 4616
rect 4616 4476 4623 4513
rect 4656 4476 4663 4616
rect 4596 4147 4603 4183
rect 4556 3956 4583 3963
rect 4336 3516 4363 3523
rect 4356 3467 4363 3516
rect 4396 3507 4403 3513
rect 4336 3267 4343 3453
rect 4416 3287 4423 3593
rect 4456 3307 4463 3493
rect 4476 3283 4483 3513
rect 4496 3327 4503 3753
rect 4556 3703 4563 3956
rect 4456 3276 4483 3283
rect 4216 3203 4223 3243
rect 4296 3236 4323 3243
rect 4176 3187 4183 3203
rect 4216 3196 4243 3203
rect 4136 3036 4143 3073
rect 3776 2736 3783 2813
rect 3796 2667 3803 2773
rect 3736 2556 3763 2563
rect 3716 1947 3723 2233
rect 3736 1823 3743 2273
rect 3756 2207 3763 2556
rect 3776 2547 3783 2613
rect 3816 2607 3823 2833
rect 3856 2756 3863 2793
rect 3896 2756 3903 2773
rect 3836 2727 3843 2743
rect 3916 2723 3923 2743
rect 3896 2716 3923 2723
rect 3816 2507 3823 2563
rect 3776 2327 3783 2393
rect 3816 2307 3823 2373
rect 3776 1823 3783 2253
rect 3796 2147 3803 2283
rect 3836 2263 3843 2713
rect 3896 2707 3903 2716
rect 3936 2707 3943 2813
rect 3976 2767 3983 2993
rect 4036 2756 4043 2813
rect 3856 2487 3863 2693
rect 3916 2576 3923 2593
rect 3956 2587 3963 2743
rect 3996 2707 4003 2743
rect 4016 2727 4023 2743
rect 3996 2647 4003 2693
rect 4056 2627 4063 2713
rect 4076 2707 4083 2763
rect 3976 2576 3983 2613
rect 4096 2607 4103 2973
rect 4116 2727 4123 2993
rect 4136 2827 4143 2993
rect 4156 2967 4163 3023
rect 4196 3016 4203 3053
rect 4176 2756 4183 2993
rect 4216 2787 4223 3153
rect 4236 3127 4243 3196
rect 4256 3167 4263 3193
rect 4256 3063 4263 3133
rect 4276 3087 4283 3193
rect 4296 3147 4303 3236
rect 4256 3056 4283 3063
rect 4276 3023 4283 3056
rect 4296 3047 4303 3113
rect 4336 3083 4343 3193
rect 4356 3187 4363 3223
rect 4356 3127 4363 3173
rect 4396 3167 4403 3223
rect 4336 3076 4363 3083
rect 4256 3016 4283 3023
rect 4236 2947 4243 3013
rect 4256 2996 4273 3003
rect 4256 2847 4263 2996
rect 4316 2996 4323 3073
rect 4336 3016 4343 3053
rect 4356 3047 4363 3076
rect 4276 2927 4283 2973
rect 3936 2487 3943 2533
rect 3876 2276 3883 2353
rect 3936 2307 3943 2473
rect 3956 2307 3963 2473
rect 3976 2327 3983 2533
rect 4016 2407 4023 2593
rect 4036 2507 4043 2553
rect 4056 2527 4063 2543
rect 4076 2467 4083 2573
rect 3996 2276 4003 2373
rect 4056 2307 4063 2433
rect 3836 2256 3863 2263
rect 3816 2147 3823 2253
rect 3856 2247 3863 2256
rect 3896 2243 3903 2263
rect 3896 2236 3933 2243
rect 3836 2107 3843 2193
rect 3816 2027 3823 2093
rect 3836 2076 3843 2093
rect 3936 2083 3943 2133
rect 3916 2076 3943 2083
rect 3676 1616 3703 1623
rect 3716 1816 3743 1823
rect 3756 1816 3783 1823
rect 3716 1623 3723 1816
rect 3736 1767 3743 1783
rect 3756 1767 3763 1816
rect 3796 1743 3803 2013
rect 3816 1823 3823 1833
rect 3816 1816 3843 1823
rect 3876 1816 3883 2073
rect 3816 1787 3823 1816
rect 3776 1736 3803 1743
rect 3776 1647 3783 1736
rect 3796 1687 3803 1713
rect 3716 1616 3743 1623
rect 3676 1603 3683 1616
rect 3656 1596 3683 1603
rect 3716 1547 3723 1583
rect 3616 1327 3623 1493
rect 3596 1263 3603 1273
rect 3636 1263 3643 1273
rect 3596 1256 3643 1263
rect 3596 827 3603 1113
rect 3616 1103 3623 1233
rect 3616 1096 3643 1103
rect 3636 867 3643 1096
rect 3656 987 3663 1453
rect 3736 1347 3743 1616
rect 3796 1616 3803 1673
rect 3756 1583 3763 1613
rect 3756 1576 3783 1583
rect 3676 1287 3683 1303
rect 3716 1283 3723 1293
rect 3716 1276 3743 1283
rect 3676 687 3683 823
rect 3716 807 3723 853
rect 3416 603 3423 633
rect 3496 603 3503 653
rect 3576 636 3583 653
rect 3716 636 3723 793
rect 3776 727 3783 1553
rect 3796 1287 3803 1573
rect 3816 1567 3823 1753
rect 3876 1747 3883 1773
rect 3836 1607 3843 1653
rect 3856 1596 3863 1693
rect 3896 1687 3903 1933
rect 3916 1867 3923 2053
rect 3956 1827 3963 2273
rect 3976 2247 3983 2263
rect 4056 2243 4063 2263
rect 4007 2236 4063 2243
rect 3927 1776 3943 1783
rect 3996 1763 4003 1953
rect 4016 1947 4023 2213
rect 4036 2087 4043 2213
rect 4056 2076 4063 2093
rect 3976 1756 4003 1763
rect 3896 1603 3903 1653
rect 3896 1596 3923 1603
rect 3956 1596 3963 1713
rect 3976 1563 3983 1756
rect 3996 1703 4003 1733
rect 4016 1727 4023 1803
rect 4056 1796 4063 2013
rect 4076 1967 4083 2453
rect 4096 2103 4103 2493
rect 4116 2447 4123 2693
rect 4156 2687 4163 2743
rect 4196 2727 4203 2743
rect 4136 2347 4143 2653
rect 4156 2303 4163 2613
rect 4136 2296 4163 2303
rect 4136 2163 4143 2296
rect 4156 2247 4163 2263
rect 4136 2156 4163 2163
rect 4096 2096 4123 2103
rect 4116 1867 4123 2096
rect 4156 1963 4163 2156
rect 4136 1956 4163 1963
rect 3996 1696 4023 1703
rect 4016 1616 4023 1696
rect 4036 1596 4043 1753
rect 4056 1667 4063 1753
rect 4076 1747 4083 1783
rect 4096 1707 4103 1763
rect 4076 1643 4083 1693
rect 4116 1667 4123 1773
rect 4056 1636 4083 1643
rect 3956 1556 3983 1563
rect 3956 1347 3963 1556
rect 3856 1147 3863 1333
rect 3876 1267 3883 1333
rect 3896 1147 3903 1303
rect 4016 1207 4023 1573
rect 4056 1547 4063 1636
rect 4096 1627 4103 1653
rect 4136 1623 4143 1956
rect 4156 1796 4163 1933
rect 4116 1616 4143 1623
rect 4156 1616 4163 1653
rect 4176 1627 4183 2713
rect 4216 2647 4223 2743
rect 4216 2267 4223 2533
rect 4236 2487 4243 2693
rect 4256 2527 4263 2743
rect 4276 2727 4283 2853
rect 4196 2256 4213 2263
rect 4196 2107 4203 2256
rect 4296 2263 4303 2973
rect 4316 2707 4323 2933
rect 4376 2783 4383 3133
rect 4396 3067 4403 3113
rect 4416 3087 4423 3213
rect 4436 3187 4443 3273
rect 4356 2776 4383 2783
rect 4356 2583 4363 2776
rect 4396 2647 4403 3053
rect 4416 2967 4423 3013
rect 4416 2727 4423 2743
rect 4436 2727 4443 2873
rect 4356 2576 4383 2583
rect 4336 2556 4363 2563
rect 4336 2547 4343 2556
rect 4276 2256 4303 2263
rect 4236 2183 4243 2233
rect 4316 2223 4323 2513
rect 4336 2256 4343 2293
rect 4316 2216 4343 2223
rect 4236 2176 4263 2183
rect 4196 2076 4223 2083
rect 4256 2076 4263 2176
rect 4296 2076 4303 2133
rect 4316 2096 4323 2113
rect 4336 2107 4343 2216
rect 4376 2147 4383 2576
rect 4436 2547 4443 2563
rect 4416 2147 4423 2253
rect 4196 1947 4203 2076
rect 4236 1927 4243 2063
rect 4036 1247 4043 1303
rect 3816 667 3823 1133
rect 3896 1107 3903 1133
rect 3856 823 3863 1093
rect 3836 816 3863 823
rect 3916 816 3923 973
rect 3936 963 3943 1193
rect 4016 1083 4023 1113
rect 3956 987 3963 1083
rect 3996 1076 4023 1083
rect 3936 956 3963 963
rect 3856 807 3863 816
rect 3936 787 3943 853
rect 3416 596 3443 603
rect 3476 596 3503 603
rect 3476 427 3483 596
rect 3796 547 3803 643
rect 3836 636 3843 673
rect 3476 387 3483 413
rect 3116 356 3123 373
rect 3236 356 3263 363
rect 3236 347 3243 356
rect 3096 307 3103 343
rect 3216 336 3233 343
rect 3396 343 3403 373
rect 3476 356 3503 363
rect 3016 176 3033 183
rect 3036 156 3043 173
rect 3076 167 3083 213
rect 2776 116 2783 153
rect 3136 147 3143 333
rect 3196 287 3203 323
rect 3276 267 3283 323
rect 3336 247 3343 343
rect 3376 336 3403 343
rect 3416 327 3423 343
rect 3496 307 3503 356
rect 3616 347 3623 393
rect 3636 356 3643 393
rect 3656 376 3683 383
rect 3716 376 3743 383
rect 3156 176 3163 213
rect 3196 143 3203 193
rect 3256 176 3283 183
rect 3276 167 3283 176
rect 3356 156 3363 293
rect 3516 287 3523 333
rect 3556 176 3563 343
rect 3596 327 3603 343
rect 3656 327 3663 376
rect 3576 307 3583 323
rect 3736 307 3743 376
rect 3796 376 3803 393
rect 3396 156 3403 173
rect 3576 167 3583 253
rect 3696 156 3703 173
rect 3736 156 3743 233
rect 3796 147 3803 173
rect 3816 167 3823 613
rect 3856 603 3863 623
rect 3836 596 3863 603
rect 3836 367 3843 596
rect 3916 587 3923 633
rect 3936 603 3943 673
rect 3956 647 3963 956
rect 4036 867 4043 1093
rect 4056 1087 4063 1123
rect 4016 836 4023 853
rect 4036 687 4043 823
rect 4116 823 4123 1616
rect 4196 1596 4203 1913
rect 4276 1847 4283 2063
rect 4316 2023 4323 2053
rect 4336 2047 4343 2053
rect 4316 2016 4343 2023
rect 4336 1787 4343 2016
rect 4356 1807 4363 2093
rect 4436 2083 4443 2513
rect 4456 2507 4463 3276
rect 4516 3256 4523 3273
rect 4476 2867 4483 3073
rect 4496 3036 4503 3073
rect 4536 3063 4543 3703
rect 4556 3696 4583 3703
rect 4516 3056 4543 3063
rect 4496 2736 4503 2773
rect 4516 2687 4523 3056
rect 4556 2987 4563 3493
rect 4596 3487 4603 3503
rect 4616 3463 4623 4433
rect 4676 4307 4683 4453
rect 4636 4127 4643 4183
rect 4636 4016 4663 4023
rect 4636 3967 4643 4016
rect 4636 3727 4643 3913
rect 4696 3783 4703 4443
rect 4716 3987 4723 4193
rect 4696 3776 4723 3783
rect 4696 3716 4703 3753
rect 4656 3667 4663 3683
rect 4596 3456 4623 3463
rect 4596 3007 4603 3456
rect 4636 3223 4643 3293
rect 4656 3267 4663 3453
rect 4676 3287 4683 3473
rect 4716 3343 4723 3776
rect 4696 3336 4723 3343
rect 4616 3047 4623 3223
rect 4636 3216 4663 3223
rect 4636 3087 4643 3216
rect 4656 3107 4663 3193
rect 4656 3063 4663 3073
rect 4676 3067 4683 3233
rect 4696 3227 4703 3336
rect 4736 3247 4743 4293
rect 4636 3056 4663 3063
rect 4636 3036 4643 3056
rect 4696 3043 4703 3213
rect 4736 3087 4743 3173
rect 4696 3036 4723 3043
rect 4616 2927 4623 3013
rect 4656 3007 4663 3023
rect 4676 2807 4683 2993
rect 4556 2756 4563 2793
rect 4536 2727 4543 2743
rect 4596 2727 4603 2763
rect 4476 2556 4483 2573
rect 4496 2487 4503 2543
rect 4536 2536 4543 2553
rect 4556 2527 4563 2693
rect 4616 2567 4623 2793
rect 4676 2776 4683 2793
rect 4596 2536 4603 2553
rect 4636 2527 4643 2733
rect 4656 2727 4663 2763
rect 4676 2536 4683 2733
rect 4696 2707 4703 2973
rect 4576 2347 4583 2513
rect 4616 2487 4623 2513
rect 4656 2507 4663 2523
rect 4656 2343 4663 2493
rect 4636 2336 4663 2343
rect 4536 2167 4543 2293
rect 4576 2276 4583 2313
rect 4556 2187 4563 2263
rect 4636 2183 4643 2336
rect 4696 2327 4703 2473
rect 4696 2296 4703 2313
rect 4636 2176 4663 2183
rect 4376 2076 4403 2083
rect 4436 2076 4463 2083
rect 4476 2076 4483 2113
rect 4376 2067 4383 2076
rect 4456 1823 4463 2076
rect 4436 1816 4463 1823
rect 4216 1627 4223 1693
rect 4236 1603 4243 1733
rect 4276 1707 4283 1763
rect 4216 1596 4243 1603
rect 4276 1596 4283 1653
rect 4216 1587 4223 1596
rect 4136 1547 4143 1583
rect 4176 1407 4183 1583
rect 4136 1336 4143 1353
rect 4176 1336 4183 1373
rect 4136 1116 4143 1133
rect 4176 1116 4183 1133
rect 4196 1087 4203 1533
rect 4216 1507 4223 1553
rect 4256 1547 4263 1573
rect 4296 1427 4303 1673
rect 4316 1667 4323 1783
rect 4356 1783 4363 1793
rect 4356 1776 4383 1783
rect 4336 1763 4343 1773
rect 4336 1756 4363 1763
rect 4336 1627 4343 1693
rect 4356 1627 4363 1756
rect 4316 1567 4323 1583
rect 4216 1303 4223 1353
rect 4216 1296 4243 1303
rect 4256 827 4263 1413
rect 4296 1343 4303 1393
rect 4296 1336 4323 1343
rect 4356 1336 4363 1553
rect 4276 1187 4283 1303
rect 4296 1127 4303 1336
rect 4376 1307 4383 1513
rect 4396 1387 4403 1733
rect 4416 1667 4423 1673
rect 4436 1667 4443 1816
rect 4456 1776 4463 1793
rect 4496 1787 4503 2053
rect 4416 1616 4423 1653
rect 4456 1567 4463 1713
rect 4476 1616 4483 1693
rect 4516 1627 4523 1833
rect 4536 1823 4543 2133
rect 4556 1847 4563 2073
rect 4536 1816 4563 1823
rect 4556 1783 4563 1816
rect 4536 1776 4563 1783
rect 4596 1747 4603 2153
rect 4636 2076 4643 2133
rect 4656 1827 4663 2176
rect 4676 2076 4683 2253
rect 4716 2163 4723 3036
rect 4736 3027 4743 3053
rect 4736 2267 4743 2993
rect 4756 2747 4763 3493
rect 4776 3087 4783 3713
rect 4776 2927 4783 3053
rect 4696 2156 4723 2163
rect 4696 1816 4703 2156
rect 4656 1727 4663 1813
rect 4476 1367 4483 1553
rect 4476 1323 4483 1353
rect 4516 1343 4523 1593
rect 4536 1583 4543 1653
rect 4536 1576 4563 1583
rect 4656 1576 4663 1673
rect 4676 1627 4683 1773
rect 4716 1607 4723 1803
rect 4776 1607 4783 2333
rect 4647 1516 4653 1523
rect 4676 1367 4683 1593
rect 4516 1336 4543 1343
rect 4536 1327 4543 1336
rect 4476 1316 4503 1323
rect 4456 1267 4463 1303
rect 4396 1116 4403 1133
rect 4336 1083 4343 1113
rect 4436 1087 4443 1153
rect 4476 1123 4483 1316
rect 4496 1127 4503 1293
rect 4516 1287 4523 1303
rect 4636 1303 4643 1353
rect 4556 1147 4563 1293
rect 4576 1287 4583 1303
rect 4616 1296 4643 1303
rect 4596 1267 4603 1283
rect 4536 1136 4553 1143
rect 4456 1116 4483 1123
rect 4316 1076 4343 1083
rect 4456 827 4463 1116
rect 4536 1116 4543 1136
rect 4576 1116 4583 1153
rect 4636 1127 4643 1296
rect 4656 1103 4663 1273
rect 4696 1127 4703 1353
rect 4736 1316 4743 1333
rect 4756 1327 4763 1593
rect 4776 1367 4783 1573
rect 4616 1096 4663 1103
rect 4676 1096 4683 1113
rect 4516 1047 4523 1083
rect 4116 816 4143 823
rect 3936 596 3963 603
rect 3856 347 3863 363
rect 3896 356 3903 413
rect 3936 356 3963 363
rect 3936 343 3943 356
rect 3876 287 3883 343
rect 3916 336 3943 343
rect 3916 267 3923 336
rect 3976 307 3983 323
rect 3936 156 3943 293
rect 3176 136 3203 143
rect 3876 143 3883 153
rect 3856 136 3883 143
rect 3916 127 3923 143
rect 3956 136 3963 213
rect 3976 127 3983 253
rect 3996 187 4003 533
rect 4016 356 4023 653
rect 4036 607 4043 633
rect 4076 367 4083 773
rect 4116 636 4123 793
rect 4096 587 4103 633
rect 4116 307 4123 333
rect 4136 327 4143 816
rect 4156 807 4163 823
rect 4176 343 4183 793
rect 4196 767 4203 823
rect 4216 607 4223 713
rect 4236 463 4243 613
rect 4316 603 4323 813
rect 4376 787 4383 823
rect 4416 807 4423 823
rect 4496 816 4503 913
rect 4556 907 4563 1073
rect 4616 927 4623 1096
rect 4556 836 4563 893
rect 4616 843 4623 873
rect 4596 836 4623 843
rect 4656 836 4663 913
rect 4676 867 4683 1053
rect 4696 1047 4703 1083
rect 4716 843 4723 1313
rect 4776 1283 4783 1313
rect 4756 1276 4783 1283
rect 4736 887 4743 1113
rect 4756 927 4763 1133
rect 4696 836 4723 843
rect 4396 603 4403 673
rect 4456 636 4463 753
rect 4496 636 4503 673
rect 4236 456 4263 463
rect 4256 347 4263 456
rect 4296 427 4303 603
rect 4316 596 4343 603
rect 4376 596 4403 603
rect 4476 527 4483 623
rect 4536 427 4543 823
rect 4576 816 4603 823
rect 4596 636 4603 816
rect 4676 816 4703 823
rect 4636 643 4643 793
rect 4676 647 4683 793
rect 4696 787 4703 816
rect 4616 636 4643 643
rect 4156 336 4183 343
rect 4036 156 4043 253
rect 4056 176 4103 183
rect 4056 147 4063 176
rect 4116 156 4123 293
rect 4196 287 4203 343
rect 4176 196 4223 203
rect 4176 187 4183 196
rect 4216 183 4223 196
rect 4216 176 4243 183
rect 4176 156 4183 173
rect 4236 156 4243 176
rect 4276 156 4283 393
rect 4356 376 4363 393
rect 4376 227 4383 373
rect 4396 347 4403 363
rect 4476 343 4483 413
rect 4616 343 4623 636
rect 4416 307 4423 343
rect 4456 336 4483 343
rect 4536 336 4563 343
rect 4616 336 4643 343
rect 4536 323 4543 336
rect 4516 316 4543 323
rect 2816 87 2823 123
rect 4336 123 4343 173
rect 4376 136 4383 213
rect 4416 123 4423 173
rect 4476 167 4483 313
rect 4516 187 4523 193
rect 4656 183 4663 633
rect 4676 307 4683 343
rect 4696 263 4703 513
rect 4696 256 4723 263
rect 4656 176 4683 183
rect 4516 156 4523 173
rect 4336 116 4363 123
rect 4396 116 4423 123
rect 4436 107 4443 133
rect 4536 123 4543 153
rect 4616 123 4623 173
rect 4716 136 4723 256
rect 4756 147 4763 893
rect 4536 116 4563 123
rect 4596 116 4623 123
rect 4736 107 4743 123
rect 1976 -24 1983 13
rect 2116 -24 2123 13
<< m3contact >>
rect 1233 4553 1247 4567
rect 1533 4553 1547 4567
rect 113 4533 127 4547
rect 193 4533 207 4547
rect 893 4533 907 4547
rect 33 4513 47 4527
rect 73 4493 87 4507
rect 93 4453 107 4467
rect 93 4413 107 4427
rect 173 4493 187 4507
rect 173 4473 187 4487
rect 153 4453 167 4467
rect 493 4513 507 4527
rect 713 4513 727 4527
rect 373 4493 387 4507
rect 433 4493 447 4507
rect 553 4493 567 4507
rect 653 4493 667 4507
rect 213 4473 227 4487
rect 233 4453 247 4467
rect 253 4453 267 4467
rect 313 4453 327 4467
rect 353 4453 367 4467
rect 53 4393 67 4407
rect 113 4393 127 4407
rect 173 4433 187 4447
rect 273 4433 287 4447
rect 153 4413 167 4427
rect 193 4413 207 4427
rect 133 4353 147 4367
rect 33 4233 47 4247
rect 93 4233 107 4247
rect 73 4213 87 4227
rect 173 4393 187 4407
rect 153 4213 167 4227
rect 93 4193 107 4207
rect 133 4193 147 4207
rect 73 4173 87 4187
rect 53 4133 67 4147
rect 53 4033 67 4047
rect 113 4153 127 4167
rect 73 4013 87 4027
rect 173 4113 187 4127
rect 153 4093 167 4107
rect 153 4073 167 4087
rect 33 3953 47 3967
rect 53 3893 67 3907
rect 133 3933 147 3947
rect 393 4473 407 4487
rect 473 4473 487 4487
rect 613 4473 627 4487
rect 413 4453 427 4467
rect 453 4453 467 4467
rect 493 4453 507 4467
rect 373 4433 387 4447
rect 333 4393 347 4407
rect 513 4433 527 4447
rect 533 4433 547 4447
rect 613 4433 627 4447
rect 553 4353 567 4367
rect 593 4353 607 4367
rect 453 4313 467 4327
rect 353 4273 367 4287
rect 413 4273 427 4287
rect 213 4213 227 4227
rect 233 4193 247 4207
rect 253 4173 267 4187
rect 193 4053 207 4067
rect 213 4013 227 4027
rect 313 4213 327 4227
rect 293 4173 307 4187
rect 313 4153 327 4167
rect 293 4133 307 4147
rect 353 4173 367 4187
rect 413 4193 427 4207
rect 473 4193 487 4207
rect 513 4193 527 4207
rect 393 4173 407 4187
rect 373 4113 387 4127
rect 493 4173 507 4187
rect 573 4313 587 4327
rect 673 4453 687 4467
rect 693 4453 707 4467
rect 653 4433 667 4447
rect 633 4413 647 4427
rect 753 4473 767 4487
rect 773 4473 787 4487
rect 833 4473 847 4487
rect 853 4473 867 4487
rect 753 4453 767 4467
rect 793 4453 807 4467
rect 813 4453 827 4467
rect 853 4453 867 4467
rect 833 4433 847 4447
rect 873 4433 887 4447
rect 713 4413 727 4427
rect 813 4413 827 4427
rect 853 4413 867 4427
rect 1053 4493 1067 4507
rect 1073 4493 1087 4507
rect 1113 4493 1127 4507
rect 1133 4493 1147 4507
rect 993 4473 1007 4487
rect 933 4453 947 4467
rect 1033 4453 1047 4467
rect 953 4433 967 4447
rect 1013 4433 1027 4447
rect 693 4393 707 4407
rect 653 4373 667 4387
rect 653 4213 667 4227
rect 693 4193 707 4207
rect 733 4373 747 4387
rect 813 4353 827 4367
rect 793 4213 807 4227
rect 773 4193 787 4207
rect 553 4153 567 4167
rect 673 4153 687 4167
rect 693 4153 707 4167
rect 713 4153 727 4167
rect 753 4153 767 4167
rect 593 4133 607 4147
rect 513 4113 527 4127
rect 593 4113 607 4127
rect 433 4093 447 4107
rect 273 4073 287 4087
rect 333 4073 347 4087
rect 293 4053 307 4067
rect 373 4033 387 4047
rect 413 4033 427 4047
rect 333 4013 347 4027
rect 493 4013 507 4027
rect 433 3993 447 4007
rect 253 3973 267 3987
rect 273 3973 287 3987
rect 193 3953 207 3967
rect 153 3873 167 3887
rect 173 3873 187 3887
rect 73 3733 87 3747
rect 133 3733 147 3747
rect 53 3713 67 3727
rect 113 3713 127 3727
rect 153 3713 167 3727
rect 73 3693 87 3707
rect 53 3673 67 3687
rect 73 3653 87 3667
rect 113 3673 127 3687
rect 53 3633 67 3647
rect 93 3633 107 3647
rect 33 3613 47 3627
rect 153 3693 167 3707
rect 133 3653 147 3667
rect 93 3613 107 3627
rect 113 3613 127 3627
rect 13 3473 27 3487
rect 13 3413 27 3427
rect 13 3393 27 3407
rect 73 3473 87 3487
rect 113 3593 127 3607
rect 113 3473 127 3487
rect 33 3273 47 3287
rect 13 3193 27 3207
rect 33 3033 47 3047
rect 93 3433 107 3447
rect 93 3253 107 3267
rect 113 3253 127 3267
rect 93 3213 107 3227
rect 93 3193 107 3207
rect 93 3153 107 3167
rect 133 3193 147 3207
rect 173 3653 187 3667
rect 173 3533 187 3547
rect 253 3913 267 3927
rect 353 3953 367 3967
rect 213 3713 227 3727
rect 313 3893 327 3907
rect 513 3993 527 4007
rect 553 3973 567 3987
rect 453 3933 467 3947
rect 573 3933 587 3947
rect 433 3913 447 3927
rect 533 3913 547 3927
rect 653 4053 667 4067
rect 613 3993 627 4007
rect 633 3973 647 3987
rect 673 3973 687 3987
rect 653 3933 667 3947
rect 393 3893 407 3907
rect 533 3893 547 3907
rect 593 3893 607 3907
rect 373 3873 387 3887
rect 413 3753 427 3767
rect 393 3733 407 3747
rect 293 3713 307 3727
rect 333 3713 347 3727
rect 353 3713 367 3727
rect 353 3693 367 3707
rect 233 3673 247 3687
rect 253 3673 267 3687
rect 313 3673 327 3687
rect 233 3633 247 3647
rect 173 3233 187 3247
rect 173 3213 187 3227
rect 213 3213 227 3227
rect 133 3173 147 3187
rect 153 3173 167 3187
rect 133 3133 147 3147
rect 313 3633 327 3647
rect 293 3433 307 3447
rect 293 3393 307 3407
rect 253 3353 267 3367
rect 253 3333 267 3347
rect 233 3193 247 3207
rect 113 3033 127 3047
rect 33 2993 47 3007
rect 13 2933 27 2947
rect 13 2773 27 2787
rect 93 3013 107 3027
rect 73 2993 87 3007
rect 153 3053 167 3067
rect 53 2973 67 2987
rect 53 2913 67 2927
rect 93 2973 107 2987
rect 73 2833 87 2847
rect 33 2753 47 2767
rect 53 2753 67 2767
rect 33 2713 47 2727
rect 13 2693 27 2707
rect 53 2693 67 2707
rect 53 2653 67 2667
rect 33 2573 47 2587
rect 13 2553 27 2567
rect 173 2933 187 2947
rect 233 3113 247 3127
rect 413 3673 427 3687
rect 373 3653 387 3667
rect 513 3733 527 3747
rect 493 3713 507 3727
rect 593 3753 607 3767
rect 633 3753 647 3767
rect 573 3713 587 3727
rect 513 3693 527 3707
rect 533 3693 547 3707
rect 573 3693 587 3707
rect 513 3653 527 3667
rect 433 3633 447 3647
rect 453 3633 467 3647
rect 373 3613 387 3627
rect 333 3573 347 3587
rect 353 3573 367 3587
rect 533 3573 547 3587
rect 373 3493 387 3507
rect 373 3453 387 3467
rect 513 3533 527 3547
rect 473 3513 487 3527
rect 553 3513 567 3527
rect 433 3493 447 3507
rect 493 3493 507 3507
rect 533 3493 547 3507
rect 413 3453 427 3467
rect 313 3313 327 3327
rect 293 3273 307 3287
rect 333 3273 347 3287
rect 553 3473 567 3487
rect 533 3353 547 3367
rect 393 3313 407 3327
rect 453 3313 467 3327
rect 513 3313 527 3327
rect 453 3293 467 3307
rect 393 3273 407 3287
rect 433 3253 447 3267
rect 373 3233 387 3247
rect 413 3233 427 3247
rect 353 3213 367 3227
rect 433 3213 447 3227
rect 353 3193 367 3207
rect 313 3173 327 3187
rect 333 3173 347 3187
rect 293 3133 307 3147
rect 273 3113 287 3127
rect 253 3073 267 3087
rect 213 2993 227 3007
rect 193 2853 207 2867
rect 133 2773 147 2787
rect 153 2773 167 2787
rect 293 3013 307 3027
rect 293 2993 307 3007
rect 253 2893 267 2907
rect 233 2813 247 2827
rect 273 2813 287 2827
rect 213 2773 227 2787
rect 193 2753 207 2767
rect 233 2753 247 2767
rect 373 3173 387 3187
rect 393 3153 407 3167
rect 313 2913 327 2927
rect 373 3033 387 3047
rect 373 2993 387 3007
rect 373 2953 387 2967
rect 473 3253 487 3267
rect 473 3213 487 3227
rect 453 3173 467 3187
rect 453 3153 467 3167
rect 433 3113 447 3127
rect 433 2953 447 2967
rect 353 2873 367 2887
rect 333 2793 347 2807
rect 293 2773 307 2787
rect 353 2773 367 2787
rect 373 2773 387 2787
rect 113 2733 127 2747
rect 93 2653 107 2667
rect 93 2613 107 2627
rect 73 2553 87 2567
rect 53 2533 67 2547
rect 13 2493 27 2507
rect 33 2393 47 2407
rect 173 2733 187 2747
rect 193 2713 207 2727
rect 253 2733 267 2747
rect 273 2733 287 2747
rect 293 2713 307 2727
rect 213 2693 227 2707
rect 173 2613 187 2627
rect 153 2593 167 2607
rect 133 2573 147 2587
rect 113 2533 127 2547
rect 153 2533 167 2547
rect 13 2313 27 2327
rect 33 2313 47 2327
rect 93 2313 107 2327
rect 53 2273 67 2287
rect 93 2273 107 2287
rect 33 2253 47 2267
rect 13 2173 27 2187
rect 73 2253 87 2267
rect 53 2093 67 2107
rect 73 2093 87 2107
rect 53 2073 67 2087
rect 13 1993 27 2007
rect 13 1873 27 1887
rect 33 1853 47 1867
rect 133 2353 147 2367
rect 253 2593 267 2607
rect 393 2753 407 2767
rect 373 2733 387 2747
rect 353 2713 367 2727
rect 413 2733 427 2747
rect 433 2733 447 2747
rect 333 2693 347 2707
rect 313 2653 327 2667
rect 233 2533 247 2547
rect 253 2533 267 2547
rect 213 2393 227 2407
rect 193 2293 207 2307
rect 313 2513 327 2527
rect 353 2613 367 2627
rect 413 2653 427 2667
rect 433 2613 447 2627
rect 473 3093 487 3107
rect 513 3073 527 3087
rect 553 3293 567 3307
rect 553 3193 567 3207
rect 813 4173 827 4187
rect 853 4173 867 4187
rect 913 4413 927 4427
rect 1053 4393 1067 4407
rect 1153 4473 1167 4487
rect 1173 4473 1187 4487
rect 1093 4453 1107 4467
rect 1133 4433 1147 4447
rect 1193 4453 1207 4467
rect 1293 4533 1307 4547
rect 1453 4533 1467 4547
rect 1273 4493 1287 4507
rect 1433 4513 1447 4527
rect 1313 4493 1327 4507
rect 1353 4493 1367 4507
rect 1333 4473 1347 4487
rect 1273 4453 1287 4467
rect 1093 4413 1107 4427
rect 1173 4413 1187 4427
rect 913 4353 927 4367
rect 953 4353 967 4367
rect 1073 4353 1087 4367
rect 1153 4353 1167 4367
rect 913 4213 927 4227
rect 953 4193 967 4207
rect 893 4173 907 4187
rect 1053 4213 1067 4227
rect 1113 4213 1127 4227
rect 1253 4433 1267 4447
rect 1393 4473 1407 4487
rect 1453 4493 1467 4507
rect 1373 4453 1387 4467
rect 1353 4413 1367 4427
rect 1493 4473 1507 4487
rect 1633 4533 1647 4547
rect 2273 4533 2287 4547
rect 2333 4533 2347 4547
rect 3333 4533 3347 4547
rect 3433 4533 3447 4547
rect 3953 4533 3967 4547
rect 1613 4513 1627 4527
rect 1553 4493 1567 4507
rect 1573 4473 1587 4487
rect 1553 4453 1567 4467
rect 1593 4453 1607 4467
rect 1513 4433 1527 4447
rect 1693 4513 1707 4527
rect 1813 4513 1827 4527
rect 1953 4513 1967 4527
rect 2013 4513 2027 4527
rect 2053 4513 2067 4527
rect 1653 4453 1667 4467
rect 1773 4493 1787 4507
rect 1913 4493 1927 4507
rect 1593 4413 1607 4427
rect 1253 4393 1267 4407
rect 1413 4393 1427 4407
rect 1553 4393 1567 4407
rect 1213 4373 1227 4387
rect 1693 4433 1707 4447
rect 1673 4253 1687 4267
rect 1393 4233 1407 4247
rect 1553 4233 1567 4247
rect 873 4153 887 4167
rect 933 4153 947 4167
rect 773 4133 787 4147
rect 893 4133 907 4147
rect 1033 4133 1047 4147
rect 713 4013 727 4027
rect 793 4053 807 4067
rect 773 3993 787 4007
rect 753 3973 767 3987
rect 853 4033 867 4047
rect 813 3973 827 3987
rect 773 3953 787 3967
rect 833 3953 847 3967
rect 933 4033 947 4047
rect 953 4033 967 4047
rect 993 3993 1007 4007
rect 1013 3993 1027 4007
rect 1093 4173 1107 4187
rect 1073 4113 1087 4127
rect 1073 4053 1087 4067
rect 973 3973 987 3987
rect 1033 3973 1047 3987
rect 973 3953 987 3967
rect 753 3933 767 3947
rect 873 3933 887 3947
rect 693 3913 707 3927
rect 853 3913 867 3927
rect 833 3773 847 3787
rect 693 3713 707 3727
rect 733 3713 747 3727
rect 793 3713 807 3727
rect 673 3693 687 3707
rect 753 3693 767 3707
rect 593 3573 607 3587
rect 653 3593 667 3607
rect 693 3673 707 3687
rect 833 3673 847 3687
rect 793 3633 807 3647
rect 693 3613 707 3627
rect 753 3613 767 3627
rect 673 3553 687 3567
rect 733 3553 747 3567
rect 653 3513 667 3527
rect 613 3393 627 3407
rect 593 3293 607 3307
rect 593 3253 607 3267
rect 593 3213 607 3227
rect 593 3173 607 3187
rect 573 3153 587 3167
rect 693 3493 707 3507
rect 673 3453 687 3467
rect 693 3453 707 3467
rect 673 3353 687 3367
rect 633 3333 647 3347
rect 653 3253 667 3267
rect 653 3173 667 3187
rect 613 3153 627 3167
rect 653 3153 667 3167
rect 633 3133 647 3147
rect 553 3093 567 3107
rect 573 3093 587 3107
rect 593 3093 607 3107
rect 533 3053 547 3067
rect 513 3033 527 3047
rect 473 2973 487 2987
rect 453 2573 467 2587
rect 393 2553 407 2567
rect 413 2533 427 2547
rect 433 2533 447 2547
rect 353 2513 367 2527
rect 373 2513 387 2527
rect 333 2453 347 2467
rect 273 2353 287 2367
rect 313 2353 327 2367
rect 413 2413 427 2427
rect 413 2333 427 2347
rect 313 2313 327 2327
rect 353 2313 367 2327
rect 293 2293 307 2307
rect 173 2273 187 2287
rect 233 2273 247 2287
rect 273 2273 287 2287
rect 133 2253 147 2267
rect 193 2233 207 2247
rect 213 2233 227 2247
rect 213 2213 227 2227
rect 233 2213 247 2227
rect 153 2193 167 2207
rect 173 2133 187 2147
rect 313 2273 327 2287
rect 353 2273 367 2287
rect 333 2253 347 2267
rect 373 2253 387 2267
rect 293 2233 307 2247
rect 333 2233 347 2247
rect 273 2213 287 2227
rect 353 2193 367 2207
rect 313 2173 327 2187
rect 273 2153 287 2167
rect 133 2073 147 2087
rect 173 2073 187 2087
rect 213 2073 227 2087
rect 233 2073 247 2087
rect 253 2073 267 2087
rect 353 2093 367 2107
rect 353 2073 367 2087
rect 73 2033 87 2047
rect 93 2033 107 2047
rect 53 1833 67 1847
rect 93 1873 107 1887
rect 113 1833 127 1847
rect 73 1813 87 1827
rect 93 1813 107 1827
rect 273 2053 287 2067
rect 293 2053 307 2067
rect 313 2053 327 2067
rect 173 2033 187 2047
rect 173 1973 187 1987
rect 253 2033 267 2047
rect 233 2013 247 2027
rect 213 1953 227 1967
rect 233 1933 247 1947
rect 293 1933 307 1947
rect 233 1913 247 1927
rect 213 1853 227 1867
rect 333 2033 347 2047
rect 313 1893 327 1907
rect 293 1853 307 1867
rect 233 1833 247 1847
rect 213 1813 227 1827
rect 153 1793 167 1807
rect 193 1793 207 1807
rect 73 1773 87 1787
rect 93 1753 107 1767
rect 33 1733 47 1747
rect 13 1713 27 1727
rect 173 1733 187 1747
rect 133 1713 147 1727
rect 113 1693 127 1707
rect 133 1673 147 1687
rect 13 1593 27 1607
rect 33 1573 47 1587
rect 93 1613 107 1627
rect 133 1613 147 1627
rect 173 1613 187 1627
rect 93 1593 107 1607
rect 113 1573 127 1587
rect 133 1573 147 1587
rect 153 1573 167 1587
rect 113 1553 127 1567
rect 53 1393 67 1407
rect 73 1393 87 1407
rect 253 1793 267 1807
rect 273 1773 287 1787
rect 253 1753 267 1767
rect 213 1733 227 1747
rect 253 1693 267 1707
rect 273 1693 287 1707
rect 213 1573 227 1587
rect 193 1553 207 1567
rect 273 1633 287 1647
rect 453 2513 467 2527
rect 533 3013 547 3027
rect 493 2933 507 2947
rect 593 3073 607 3087
rect 593 3033 607 3047
rect 593 3013 607 3027
rect 573 2993 587 3007
rect 613 2933 627 2947
rect 553 2913 567 2927
rect 573 2893 587 2907
rect 553 2833 567 2847
rect 553 2813 567 2827
rect 533 2793 547 2807
rect 713 3373 727 3387
rect 753 3533 767 3547
rect 833 3533 847 3547
rect 833 3513 847 3527
rect 753 3373 767 3387
rect 733 3353 747 3367
rect 813 3433 827 3447
rect 773 3333 787 3347
rect 793 3273 807 3287
rect 733 3213 747 3227
rect 733 3193 747 3207
rect 873 3793 887 3807
rect 953 3773 967 3787
rect 913 3733 927 3747
rect 1093 3953 1107 3967
rect 1033 3933 1047 3947
rect 1233 4193 1247 4207
rect 1293 4213 1307 4227
rect 1313 4193 1327 4207
rect 1433 4213 1447 4227
rect 1473 4213 1487 4227
rect 1233 4173 1247 4187
rect 1273 4173 1287 4187
rect 1333 4173 1347 4187
rect 1133 4133 1147 4147
rect 1193 4133 1207 4147
rect 1213 4033 1227 4047
rect 1133 3973 1147 3987
rect 1113 3893 1127 3907
rect 1333 4113 1347 4127
rect 1233 4013 1247 4027
rect 1193 3953 1207 3967
rect 1393 4173 1407 4187
rect 1353 4093 1367 4107
rect 1373 4033 1387 4047
rect 1353 4013 1367 4027
rect 1293 3973 1307 3987
rect 1333 3973 1347 3987
rect 1453 4193 1467 4207
rect 1453 4133 1467 4147
rect 1413 4113 1427 4127
rect 1413 4093 1427 4107
rect 1393 3993 1407 4007
rect 1393 3953 1407 3967
rect 1433 4013 1447 4027
rect 1493 4153 1507 4167
rect 1993 4473 2007 4487
rect 2173 4493 2187 4507
rect 1753 4393 1767 4407
rect 1893 4453 1907 4467
rect 1833 4433 1847 4447
rect 2013 4453 2027 4467
rect 1973 4433 1987 4447
rect 2033 4393 2047 4407
rect 1793 4313 1807 4327
rect 1893 4313 1907 4327
rect 1933 4313 1947 4327
rect 1793 4233 1807 4247
rect 1553 4193 1567 4207
rect 1733 4193 1747 4207
rect 1833 4213 1847 4227
rect 1873 4213 1887 4227
rect 1933 4233 1947 4247
rect 1913 4213 1927 4227
rect 1813 4193 1827 4207
rect 1533 4073 1547 4087
rect 1473 4013 1487 4027
rect 1513 3993 1527 4007
rect 1453 3953 1467 3967
rect 1493 3953 1507 3967
rect 1413 3933 1427 3947
rect 1473 3933 1487 3947
rect 1233 3893 1247 3907
rect 1273 3893 1287 3907
rect 1033 3793 1047 3807
rect 1173 3793 1187 3807
rect 993 3753 1007 3767
rect 973 3713 987 3727
rect 1033 3733 1047 3747
rect 1073 3733 1087 3747
rect 1113 3733 1127 3747
rect 1053 3713 1067 3727
rect 933 3693 947 3707
rect 1013 3693 1027 3707
rect 1053 3693 1067 3707
rect 1093 3713 1107 3727
rect 913 3673 927 3687
rect 933 3673 947 3687
rect 973 3673 987 3687
rect 1073 3673 1087 3687
rect 873 3533 887 3547
rect 873 3493 887 3507
rect 893 3493 907 3507
rect 853 3393 867 3407
rect 833 3293 847 3307
rect 813 3253 827 3267
rect 933 3653 947 3667
rect 1073 3633 1087 3647
rect 1193 3713 1207 3727
rect 1133 3693 1147 3707
rect 1173 3673 1187 3687
rect 1213 3673 1227 3687
rect 1133 3613 1147 3627
rect 1073 3593 1087 3607
rect 1093 3593 1107 3607
rect 993 3573 1007 3587
rect 1113 3573 1127 3587
rect 973 3553 987 3567
rect 1013 3533 1027 3547
rect 1053 3533 1067 3547
rect 1093 3533 1107 3547
rect 993 3513 1007 3527
rect 1153 3573 1167 3587
rect 1333 3853 1347 3867
rect 1413 3753 1427 3767
rect 1373 3733 1387 3747
rect 1273 3713 1287 3727
rect 1353 3713 1367 3727
rect 1433 3713 1447 3727
rect 1673 4153 1687 4167
rect 1613 4093 1627 4107
rect 1653 4093 1667 4107
rect 1653 4013 1667 4027
rect 1753 4173 1767 4187
rect 1713 4113 1727 4127
rect 1713 4093 1727 4107
rect 1593 3993 1607 4007
rect 1633 3993 1647 4007
rect 1673 3993 1687 4007
rect 1693 3993 1707 4007
rect 1893 4193 1907 4207
rect 1973 4213 1987 4227
rect 2013 4213 2027 4227
rect 1933 4173 1947 4187
rect 1893 4153 1907 4167
rect 1853 4133 1867 4147
rect 1873 4073 1887 4087
rect 1813 4053 1827 4067
rect 1793 4033 1807 4047
rect 1753 3993 1767 4007
rect 1773 3993 1787 4007
rect 1533 3933 1547 3947
rect 1513 3853 1527 3867
rect 1573 3853 1587 3867
rect 1633 3753 1647 3767
rect 1573 3733 1587 3747
rect 1493 3713 1507 3727
rect 1533 3713 1547 3727
rect 1473 3693 1487 3707
rect 1513 3693 1527 3707
rect 1553 3693 1567 3707
rect 1253 3673 1267 3687
rect 1393 3673 1407 3687
rect 1413 3673 1427 3687
rect 1453 3673 1467 3687
rect 1253 3653 1267 3667
rect 1373 3633 1387 3647
rect 1273 3553 1287 3567
rect 1233 3533 1247 3547
rect 1013 3493 1027 3507
rect 1033 3493 1047 3507
rect 993 3473 1007 3487
rect 1033 3473 1047 3487
rect 1113 3493 1127 3507
rect 1153 3493 1167 3507
rect 1093 3473 1107 3487
rect 1073 3433 1087 3447
rect 933 3393 947 3407
rect 1013 3393 1027 3407
rect 913 3353 927 3367
rect 973 3353 987 3367
rect 913 3273 927 3287
rect 873 3253 887 3267
rect 953 3253 967 3267
rect 873 3233 887 3247
rect 933 3233 947 3247
rect 853 3213 867 3227
rect 893 3213 907 3227
rect 673 3133 687 3147
rect 693 3013 707 3027
rect 673 2993 687 3007
rect 713 2993 727 3007
rect 673 2973 687 2987
rect 653 2893 667 2907
rect 613 2833 627 2847
rect 493 2753 507 2767
rect 573 2773 587 2787
rect 493 2733 507 2747
rect 553 2733 567 2747
rect 573 2733 587 2747
rect 533 2713 547 2727
rect 513 2573 527 2587
rect 553 2593 567 2607
rect 533 2533 547 2547
rect 473 2473 487 2487
rect 533 2513 547 2527
rect 613 2733 627 2747
rect 693 2953 707 2967
rect 713 2953 727 2967
rect 673 2813 687 2827
rect 793 3193 807 3207
rect 813 3193 827 3207
rect 833 3193 847 3207
rect 773 3173 787 3187
rect 753 3153 767 3167
rect 793 3093 807 3107
rect 753 3033 767 3047
rect 873 3173 887 3187
rect 873 3153 887 3167
rect 833 3053 847 3067
rect 833 3033 847 3047
rect 853 3033 867 3047
rect 813 2993 827 3007
rect 773 2973 787 2987
rect 753 2933 767 2947
rect 733 2833 747 2847
rect 713 2793 727 2807
rect 753 2793 767 2807
rect 993 3273 1007 3287
rect 1093 3373 1107 3387
rect 1093 3333 1107 3347
rect 1133 3333 1147 3347
rect 1053 3253 1067 3267
rect 993 3233 1007 3247
rect 1073 3233 1087 3247
rect 1073 3213 1087 3227
rect 933 3153 947 3167
rect 973 3153 987 3167
rect 913 3113 927 3127
rect 993 3093 1007 3107
rect 1073 3093 1087 3107
rect 973 3033 987 3047
rect 933 2993 947 3007
rect 893 2973 907 2987
rect 873 2953 887 2967
rect 873 2893 887 2907
rect 853 2833 867 2847
rect 833 2813 847 2827
rect 673 2733 687 2747
rect 613 2693 627 2707
rect 653 2693 667 2707
rect 613 2613 627 2627
rect 593 2593 607 2607
rect 613 2573 627 2587
rect 813 2773 827 2787
rect 733 2733 747 2747
rect 773 2693 787 2707
rect 713 2573 727 2587
rect 613 2513 627 2527
rect 573 2493 587 2507
rect 593 2473 607 2487
rect 493 2413 507 2427
rect 573 2413 587 2427
rect 453 2353 467 2367
rect 433 2273 447 2287
rect 513 2313 527 2327
rect 473 2253 487 2267
rect 433 2233 447 2247
rect 473 2233 487 2247
rect 393 2213 407 2227
rect 453 2113 467 2127
rect 473 2093 487 2107
rect 533 2273 547 2287
rect 553 2253 567 2267
rect 513 2213 527 2227
rect 393 2053 407 2067
rect 413 2053 427 2067
rect 433 2053 447 2067
rect 393 2033 407 2047
rect 393 1873 407 1887
rect 373 1853 387 1867
rect 433 2033 447 2047
rect 453 1853 467 1867
rect 413 1833 427 1847
rect 333 1813 347 1827
rect 373 1813 387 1827
rect 433 1813 447 1827
rect 593 2253 607 2267
rect 693 2513 707 2527
rect 673 2373 687 2387
rect 833 2753 847 2767
rect 813 2733 827 2747
rect 853 2733 867 2747
rect 813 2653 827 2667
rect 833 2653 847 2667
rect 793 2633 807 2647
rect 793 2613 807 2627
rect 753 2513 767 2527
rect 713 2473 727 2487
rect 853 2613 867 2627
rect 833 2553 847 2567
rect 893 2833 907 2847
rect 893 2733 907 2747
rect 913 2733 927 2747
rect 1033 3073 1047 3087
rect 1013 3053 1027 3067
rect 1133 3293 1147 3307
rect 1113 3213 1127 3227
rect 1133 3153 1147 3167
rect 1113 3133 1127 3147
rect 1233 3493 1247 3507
rect 1193 3473 1207 3487
rect 1253 3473 1267 3487
rect 1253 3413 1267 3427
rect 1213 3393 1227 3407
rect 1213 3313 1227 3327
rect 1173 3293 1187 3307
rect 1413 3513 1427 3527
rect 1313 3493 1327 3507
rect 1293 3473 1307 3487
rect 1333 3473 1347 3487
rect 1373 3473 1387 3487
rect 1433 3493 1447 3507
rect 1373 3353 1387 3367
rect 1173 3253 1187 3267
rect 1173 3193 1187 3207
rect 1173 3093 1187 3107
rect 1253 3253 1267 3267
rect 1273 3253 1287 3267
rect 1273 3233 1287 3247
rect 1313 3233 1327 3247
rect 1353 3233 1367 3247
rect 1213 3153 1227 3167
rect 1233 3153 1247 3167
rect 1213 3113 1227 3127
rect 1193 3073 1207 3087
rect 1153 3053 1167 3067
rect 1173 3053 1187 3067
rect 993 2993 1007 3007
rect 1013 2953 1027 2967
rect 1053 2953 1067 2967
rect 953 2933 967 2947
rect 953 2773 967 2787
rect 933 2633 947 2647
rect 913 2573 927 2587
rect 893 2553 907 2567
rect 873 2533 887 2547
rect 1173 3013 1187 3027
rect 1253 3073 1267 3087
rect 1333 3193 1347 3207
rect 1433 3333 1447 3347
rect 1393 3253 1407 3267
rect 1433 3213 1447 3227
rect 1413 3153 1427 3167
rect 1393 3133 1407 3147
rect 1293 3073 1307 3087
rect 1273 3033 1287 3047
rect 1233 3013 1247 3027
rect 1093 2933 1107 2947
rect 1253 2993 1267 3007
rect 1273 2993 1287 3007
rect 1233 2973 1247 2987
rect 1113 2873 1127 2887
rect 1173 2873 1187 2887
rect 1053 2813 1067 2827
rect 1093 2773 1107 2787
rect 1013 2753 1027 2767
rect 973 2733 987 2747
rect 973 2653 987 2667
rect 953 2593 967 2607
rect 1013 2713 1027 2727
rect 993 2633 1007 2647
rect 953 2573 967 2587
rect 973 2573 987 2587
rect 1053 2733 1067 2747
rect 1073 2733 1087 2747
rect 1033 2693 1047 2707
rect 1033 2613 1047 2627
rect 993 2553 1007 2567
rect 1013 2553 1027 2567
rect 833 2513 847 2527
rect 873 2513 887 2527
rect 953 2513 967 2527
rect 933 2493 947 2507
rect 813 2473 827 2487
rect 833 2473 847 2487
rect 773 2453 787 2467
rect 753 2393 767 2407
rect 633 2313 647 2327
rect 653 2293 667 2307
rect 753 2353 767 2367
rect 733 2293 747 2307
rect 673 2273 687 2287
rect 693 2273 707 2287
rect 573 2213 587 2227
rect 553 2193 567 2207
rect 533 2153 547 2167
rect 673 2213 687 2227
rect 653 2193 667 2207
rect 573 2173 587 2187
rect 573 2113 587 2127
rect 513 2033 527 2047
rect 553 2033 567 2047
rect 513 1993 527 2007
rect 473 1833 487 1847
rect 333 1773 347 1787
rect 313 1713 327 1727
rect 293 1613 307 1627
rect 293 1573 307 1587
rect 193 1453 207 1467
rect 93 1373 107 1387
rect 133 1373 147 1387
rect 53 1333 67 1347
rect 233 1373 247 1387
rect 313 1533 327 1547
rect 293 1433 307 1447
rect 253 1353 267 1367
rect 273 1353 287 1367
rect 373 1773 387 1787
rect 353 1753 367 1767
rect 353 1653 367 1667
rect 453 1773 467 1787
rect 493 1773 507 1787
rect 553 1913 567 1927
rect 533 1773 547 1787
rect 593 2053 607 2067
rect 633 2113 647 2127
rect 653 2073 667 2087
rect 633 2053 647 2067
rect 633 2013 647 2027
rect 613 1893 627 1907
rect 573 1853 587 1867
rect 573 1813 587 1827
rect 613 1773 627 1787
rect 653 1973 667 1987
rect 713 2173 727 2187
rect 753 2133 767 2147
rect 713 2113 727 2127
rect 813 2393 827 2407
rect 793 2253 807 2267
rect 913 2453 927 2467
rect 873 2393 887 2407
rect 913 2293 927 2307
rect 853 2253 867 2267
rect 833 2233 847 2247
rect 833 2213 847 2227
rect 813 2193 827 2207
rect 793 2113 807 2127
rect 773 2093 787 2107
rect 793 2093 807 2107
rect 693 2053 707 2067
rect 713 2033 727 2047
rect 693 1953 707 1967
rect 673 1913 687 1927
rect 753 2033 767 2047
rect 733 1993 747 2007
rect 713 1893 727 1907
rect 713 1833 727 1847
rect 673 1813 687 1827
rect 673 1793 687 1807
rect 533 1753 547 1767
rect 593 1753 607 1767
rect 633 1753 647 1767
rect 413 1733 427 1747
rect 513 1733 527 1747
rect 393 1713 407 1727
rect 373 1593 387 1607
rect 453 1693 467 1707
rect 413 1633 427 1647
rect 433 1593 447 1607
rect 373 1573 387 1587
rect 413 1573 427 1587
rect 433 1553 447 1567
rect 373 1433 387 1447
rect 353 1413 367 1427
rect 353 1393 367 1407
rect 93 1313 107 1327
rect 113 1313 127 1327
rect 13 1133 27 1147
rect 173 1333 187 1347
rect 233 1333 247 1347
rect 153 1293 167 1307
rect 173 1293 187 1307
rect 73 1273 87 1287
rect 133 1273 147 1287
rect 53 1253 67 1267
rect 13 1113 27 1127
rect 33 1113 47 1127
rect 153 1153 167 1167
rect 93 1133 107 1147
rect 113 1133 127 1147
rect 173 1113 187 1127
rect 33 1093 47 1107
rect 73 1093 87 1107
rect 133 1093 147 1107
rect 213 1173 227 1187
rect 253 1313 267 1327
rect 233 1133 247 1147
rect 213 1113 227 1127
rect 93 1073 107 1087
rect 13 933 27 947
rect 73 873 87 887
rect 13 793 27 807
rect 353 1353 367 1367
rect 333 1333 347 1347
rect 413 1413 427 1427
rect 393 1373 407 1387
rect 493 1633 507 1647
rect 473 1613 487 1627
rect 473 1493 487 1507
rect 453 1453 467 1467
rect 433 1393 447 1407
rect 393 1333 407 1347
rect 413 1333 427 1347
rect 693 1773 707 1787
rect 653 1733 667 1747
rect 653 1713 667 1727
rect 633 1653 647 1667
rect 573 1633 587 1647
rect 593 1633 607 1647
rect 533 1613 547 1627
rect 353 1313 367 1327
rect 413 1313 427 1327
rect 533 1533 547 1547
rect 573 1573 587 1587
rect 633 1613 647 1627
rect 613 1573 627 1587
rect 733 1813 747 1827
rect 733 1773 747 1787
rect 813 2073 827 2087
rect 913 2253 927 2267
rect 1133 2813 1147 2827
rect 1113 2693 1127 2707
rect 1193 2793 1207 2807
rect 1193 2773 1207 2787
rect 1153 2733 1167 2747
rect 1173 2733 1187 2747
rect 1293 2953 1307 2967
rect 1253 2773 1267 2787
rect 1213 2693 1227 2707
rect 1133 2673 1147 2687
rect 1093 2653 1107 2667
rect 1353 2873 1367 2887
rect 1313 2813 1327 2827
rect 1293 2713 1307 2727
rect 1253 2693 1267 2707
rect 1133 2633 1147 2647
rect 1153 2633 1167 2647
rect 1233 2633 1247 2647
rect 1093 2593 1107 2607
rect 1053 2553 1067 2567
rect 993 2513 1007 2527
rect 973 2493 987 2507
rect 953 2473 967 2487
rect 973 2433 987 2447
rect 953 2333 967 2347
rect 953 2293 967 2307
rect 953 2253 967 2267
rect 1013 2473 1027 2487
rect 1033 2393 1047 2407
rect 993 2373 1007 2387
rect 993 2293 1007 2307
rect 1033 2273 1047 2287
rect 1073 2513 1087 2527
rect 1073 2433 1087 2447
rect 1173 2593 1187 2607
rect 1233 2593 1247 2607
rect 1153 2533 1167 2547
rect 1193 2573 1207 2587
rect 1233 2573 1247 2587
rect 1153 2513 1167 2527
rect 1193 2513 1207 2527
rect 1133 2493 1147 2507
rect 1113 2453 1127 2467
rect 1153 2373 1167 2387
rect 1113 2313 1127 2327
rect 1133 2313 1147 2327
rect 1093 2293 1107 2307
rect 1013 2253 1027 2267
rect 1053 2253 1067 2267
rect 1073 2253 1087 2267
rect 1593 3713 1607 3727
rect 1673 3713 1687 3727
rect 1753 3713 1767 3727
rect 1693 3693 1707 3707
rect 1713 3693 1727 3707
rect 1733 3693 1747 3707
rect 1773 3693 1787 3707
rect 1573 3673 1587 3687
rect 1613 3673 1627 3687
rect 1653 3673 1667 3687
rect 1753 3673 1767 3687
rect 1553 3653 1567 3667
rect 1633 3633 1647 3647
rect 1573 3613 1587 3627
rect 1533 3593 1547 3607
rect 1553 3513 1567 3527
rect 1473 3393 1487 3407
rect 1453 3193 1467 3207
rect 1493 3253 1507 3267
rect 1513 3253 1527 3267
rect 1553 3233 1567 3247
rect 1533 3213 1547 3227
rect 1553 3193 1567 3207
rect 1493 3173 1507 3187
rect 1513 3173 1527 3187
rect 1473 3153 1487 3167
rect 1493 3093 1507 3107
rect 1473 3073 1487 3087
rect 1513 3073 1527 3087
rect 1593 3553 1607 3567
rect 1593 3473 1607 3487
rect 1813 4013 1827 4027
rect 1833 3993 1847 4007
rect 1973 4153 1987 4167
rect 1933 4033 1947 4047
rect 1913 4013 1927 4027
rect 1953 4013 1967 4027
rect 1913 3973 1927 3987
rect 1833 3953 1847 3967
rect 1853 3953 1867 3967
rect 1813 3933 1827 3947
rect 1893 3753 1907 3767
rect 1813 3693 1827 3707
rect 1993 4093 2007 4107
rect 2213 4473 2227 4487
rect 2133 4453 2147 4467
rect 2193 4453 2207 4467
rect 2253 4433 2267 4447
rect 2093 4313 2107 4327
rect 2113 4273 2127 4287
rect 2293 4513 2307 4527
rect 3013 4513 3027 4527
rect 3053 4513 3067 4527
rect 3093 4513 3107 4527
rect 2393 4493 2407 4507
rect 2473 4493 2487 4507
rect 2513 4493 2527 4507
rect 2933 4493 2947 4507
rect 2993 4493 3007 4507
rect 2373 4473 2387 4487
rect 2433 4473 2447 4487
rect 2313 4453 2327 4467
rect 2353 4433 2367 4447
rect 2093 4193 2107 4207
rect 2073 4133 2087 4147
rect 2133 4113 2147 4127
rect 2173 4113 2187 4127
rect 2073 4093 2087 4107
rect 2053 4033 2067 4047
rect 1973 3973 1987 3987
rect 1993 3953 2007 3967
rect 2093 3973 2107 3987
rect 2153 3973 2167 3987
rect 2353 4173 2367 4187
rect 2313 4093 2327 4107
rect 2273 4073 2287 4087
rect 2253 4053 2267 4067
rect 2213 3973 2227 3987
rect 2273 4033 2287 4047
rect 2273 3993 2287 4007
rect 2293 3973 2307 3987
rect 2453 4453 2467 4467
rect 2493 4433 2507 4447
rect 2533 4433 2547 4447
rect 2433 4413 2447 4427
rect 2413 4393 2427 4407
rect 2373 4033 2387 4047
rect 2393 4013 2407 4027
rect 2353 3993 2367 4007
rect 2453 4373 2467 4387
rect 2613 4473 2627 4487
rect 2653 4473 2667 4487
rect 2793 4473 2807 4487
rect 2713 4453 2727 4467
rect 2673 4433 2687 4447
rect 2573 4413 2587 4427
rect 2633 4413 2647 4427
rect 2673 4233 2687 4247
rect 2493 4193 2507 4207
rect 2553 4173 2567 4187
rect 2593 4173 2607 4187
rect 2633 4173 2647 4187
rect 2513 4153 2527 4167
rect 2553 4153 2567 4167
rect 2593 4153 2607 4167
rect 2433 4013 2447 4027
rect 2573 4013 2587 4027
rect 1953 3753 1967 3767
rect 1933 3733 1947 3747
rect 1973 3733 1987 3747
rect 2053 3713 2067 3727
rect 1953 3693 1967 3707
rect 1873 3673 1887 3687
rect 1913 3673 1927 3687
rect 1953 3673 1967 3687
rect 1993 3673 2007 3687
rect 1833 3653 1847 3667
rect 1693 3533 1707 3547
rect 1793 3533 1807 3547
rect 1833 3533 1847 3547
rect 1673 3513 1687 3527
rect 1673 3473 1687 3487
rect 1673 3413 1687 3427
rect 1673 3373 1687 3387
rect 1633 3313 1647 3327
rect 1593 3253 1607 3267
rect 1633 3253 1647 3267
rect 1613 3233 1627 3247
rect 1713 3513 1727 3527
rect 1793 3513 1807 3527
rect 1753 3493 1767 3507
rect 1733 3453 1747 3467
rect 1753 3453 1767 3467
rect 1713 3393 1727 3407
rect 1713 3353 1727 3367
rect 1733 3353 1747 3367
rect 1693 3253 1707 3267
rect 1613 3153 1627 3167
rect 1573 3033 1587 3047
rect 1513 3013 1527 3027
rect 1553 3013 1567 3027
rect 1413 2993 1427 3007
rect 1393 2973 1407 2987
rect 1473 2993 1487 3007
rect 1373 2793 1387 2807
rect 1353 2753 1367 2767
rect 1313 2653 1327 2667
rect 1333 2653 1347 2667
rect 1293 2613 1307 2627
rect 1273 2553 1287 2567
rect 1333 2593 1347 2607
rect 1373 2733 1387 2747
rect 1373 2573 1387 2587
rect 1353 2553 1367 2567
rect 1273 2493 1287 2507
rect 1253 2393 1267 2407
rect 1193 2333 1207 2347
rect 1253 2293 1267 2307
rect 1173 2273 1187 2287
rect 1213 2273 1227 2287
rect 953 2233 967 2247
rect 973 2233 987 2247
rect 1093 2233 1107 2247
rect 933 2213 947 2227
rect 913 2193 927 2207
rect 893 2153 907 2167
rect 933 2113 947 2127
rect 893 2093 907 2107
rect 1173 2253 1187 2267
rect 973 2213 987 2227
rect 1133 2213 1147 2227
rect 1153 2213 1167 2227
rect 813 2053 827 2067
rect 793 2013 807 2027
rect 933 2073 947 2087
rect 953 2073 967 2087
rect 913 2053 927 2067
rect 873 2033 887 2047
rect 913 2033 927 2047
rect 773 1993 787 2007
rect 853 1993 867 2007
rect 853 1953 867 1967
rect 773 1913 787 1927
rect 833 1873 847 1887
rect 813 1853 827 1867
rect 813 1813 827 1827
rect 793 1793 807 1807
rect 893 2013 907 2027
rect 933 2013 947 2027
rect 893 1973 907 1987
rect 893 1873 907 1887
rect 873 1853 887 1867
rect 853 1833 867 1847
rect 1033 2113 1047 2127
rect 1013 2093 1027 2107
rect 993 2073 1007 2087
rect 1013 2053 1027 2067
rect 1113 2093 1127 2107
rect 1153 2073 1167 2087
rect 1013 2033 1027 2047
rect 1093 2053 1107 2067
rect 1133 2053 1147 2067
rect 1153 2033 1167 2047
rect 993 2013 1007 2027
rect 1033 2013 1047 2027
rect 1053 2013 1067 2027
rect 1093 2013 1107 2027
rect 973 1993 987 2007
rect 993 1973 1007 1987
rect 1013 1893 1027 1907
rect 953 1873 967 1887
rect 953 1853 967 1867
rect 913 1813 927 1827
rect 753 1733 767 1747
rect 753 1693 767 1707
rect 713 1633 727 1647
rect 653 1593 667 1607
rect 553 1513 567 1527
rect 333 1293 347 1307
rect 373 1293 387 1307
rect 313 1273 327 1287
rect 273 1213 287 1227
rect 293 1193 307 1207
rect 353 1273 367 1287
rect 293 1173 307 1187
rect 333 1173 347 1187
rect 373 1173 387 1187
rect 433 1233 447 1247
rect 493 1313 507 1327
rect 513 1313 527 1327
rect 533 1313 547 1327
rect 453 1213 467 1227
rect 493 1273 507 1287
rect 373 1153 387 1167
rect 393 1153 407 1167
rect 413 1153 427 1167
rect 333 1133 347 1147
rect 353 1133 367 1147
rect 253 1113 267 1127
rect 293 1113 307 1127
rect 373 1113 387 1127
rect 253 1093 267 1107
rect 273 1073 287 1087
rect 173 1053 187 1067
rect 193 1053 207 1067
rect 253 1053 267 1067
rect 433 1133 447 1147
rect 413 1113 427 1127
rect 433 1093 447 1107
rect 453 1093 467 1107
rect 393 1073 407 1087
rect 473 1073 487 1087
rect 553 1273 567 1287
rect 613 1553 627 1567
rect 653 1533 667 1547
rect 613 1313 627 1327
rect 653 1313 667 1327
rect 593 1273 607 1287
rect 613 1273 627 1287
rect 593 1253 607 1267
rect 573 1233 587 1247
rect 513 1213 527 1227
rect 573 1213 587 1227
rect 553 1193 567 1207
rect 533 1133 547 1147
rect 553 1133 567 1147
rect 633 1233 647 1247
rect 613 1193 627 1207
rect 593 1173 607 1187
rect 613 1173 627 1187
rect 653 1173 667 1187
rect 513 1093 527 1107
rect 553 1093 567 1107
rect 533 1073 547 1087
rect 573 1073 587 1087
rect 353 1053 367 1067
rect 493 1053 507 1067
rect 533 1053 547 1067
rect 513 913 527 927
rect 493 893 507 907
rect 293 873 307 887
rect 413 873 427 887
rect 113 813 127 827
rect 133 813 147 827
rect 53 653 67 667
rect 253 853 267 867
rect 153 793 167 807
rect 193 813 207 827
rect 173 773 187 787
rect 253 833 267 847
rect 233 813 247 827
rect 373 853 387 867
rect 333 833 347 847
rect 213 693 227 707
rect 253 693 267 707
rect 153 673 167 687
rect 133 653 147 667
rect 193 653 207 667
rect 233 633 247 647
rect 133 613 147 627
rect 153 613 167 627
rect 93 393 107 407
rect 193 613 207 627
rect 173 593 187 607
rect 213 593 227 607
rect 233 413 247 427
rect 153 373 167 387
rect 93 333 107 347
rect 73 313 87 327
rect 33 193 47 207
rect 73 173 87 187
rect 193 373 207 387
rect 353 813 367 827
rect 393 813 407 827
rect 293 773 307 787
rect 313 673 327 687
rect 353 673 367 687
rect 273 653 287 667
rect 453 853 467 867
rect 433 793 447 807
rect 393 693 407 707
rect 413 693 427 707
rect 373 653 387 667
rect 273 633 287 647
rect 353 633 367 647
rect 313 613 327 627
rect 333 613 347 627
rect 433 673 447 687
rect 393 613 407 627
rect 293 593 307 607
rect 273 573 287 587
rect 373 593 387 607
rect 313 513 327 527
rect 353 493 367 507
rect 313 453 327 467
rect 333 413 347 427
rect 213 353 227 367
rect 253 353 267 367
rect 173 333 187 347
rect 293 333 307 347
rect 313 333 327 347
rect 253 313 267 327
rect 133 193 147 207
rect 233 193 247 207
rect 113 173 127 187
rect 93 153 107 167
rect 173 153 187 167
rect 73 133 87 147
rect 113 133 127 147
rect 153 133 167 147
rect 393 433 407 447
rect 353 373 367 387
rect 373 373 387 387
rect 493 833 507 847
rect 493 793 507 807
rect 553 1033 567 1047
rect 573 893 587 907
rect 573 853 587 867
rect 593 833 607 847
rect 653 1153 667 1167
rect 713 1613 727 1627
rect 773 1633 787 1647
rect 693 1573 707 1587
rect 713 1573 727 1587
rect 693 1553 707 1567
rect 693 1493 707 1507
rect 733 1513 747 1527
rect 733 1453 747 1467
rect 713 1373 727 1387
rect 733 1333 747 1347
rect 713 1313 727 1327
rect 733 1293 747 1307
rect 713 1273 727 1287
rect 753 1273 767 1287
rect 693 1253 707 1267
rect 713 1213 727 1227
rect 713 1193 727 1207
rect 733 1173 747 1187
rect 813 1773 827 1787
rect 853 1773 867 1787
rect 873 1773 887 1787
rect 813 1753 827 1767
rect 853 1753 867 1767
rect 873 1753 887 1767
rect 813 1713 827 1727
rect 853 1713 867 1727
rect 813 1613 827 1627
rect 793 1593 807 1607
rect 933 1773 947 1787
rect 913 1733 927 1747
rect 1033 1853 1047 1867
rect 1013 1833 1027 1847
rect 1033 1833 1047 1847
rect 1073 1993 1087 2007
rect 993 1813 1007 1827
rect 1033 1813 1047 1827
rect 1053 1813 1067 1827
rect 973 1793 987 1807
rect 1233 2253 1247 2267
rect 1193 2233 1207 2247
rect 1253 2213 1267 2227
rect 1213 2093 1227 2107
rect 1253 2073 1267 2087
rect 1453 2973 1467 2987
rect 1553 2993 1567 3007
rect 1533 2973 1547 2987
rect 1453 2913 1467 2927
rect 1493 2913 1507 2927
rect 1573 2973 1587 2987
rect 1553 2853 1567 2867
rect 1453 2753 1467 2767
rect 1613 3033 1627 3047
rect 1593 2953 1607 2967
rect 1613 2953 1627 2967
rect 1573 2833 1587 2847
rect 1473 2673 1487 2687
rect 1433 2573 1447 2587
rect 1453 2573 1467 2587
rect 1493 2593 1507 2607
rect 1493 2573 1507 2587
rect 1473 2553 1487 2567
rect 1433 2533 1447 2547
rect 1393 2493 1407 2507
rect 1413 2493 1427 2507
rect 1353 2473 1367 2487
rect 1413 2473 1427 2487
rect 1313 2333 1327 2347
rect 1353 2333 1367 2347
rect 1313 2313 1327 2327
rect 1333 2233 1347 2247
rect 1313 2133 1327 2147
rect 1293 2073 1307 2087
rect 1333 2073 1347 2087
rect 1193 2053 1207 2067
rect 1213 2053 1227 2067
rect 1113 1993 1127 2007
rect 1173 1993 1187 2007
rect 1093 1833 1107 1847
rect 1093 1813 1107 1827
rect 1013 1773 1027 1787
rect 1033 1773 1047 1787
rect 953 1733 967 1747
rect 1013 1733 1027 1747
rect 1033 1733 1047 1747
rect 933 1693 947 1707
rect 973 1673 987 1687
rect 913 1633 927 1647
rect 913 1613 927 1627
rect 953 1613 967 1627
rect 873 1593 887 1607
rect 793 1573 807 1587
rect 813 1573 827 1587
rect 833 1573 847 1587
rect 873 1573 887 1587
rect 813 1553 827 1567
rect 853 1553 867 1567
rect 913 1573 927 1587
rect 933 1573 947 1587
rect 893 1553 907 1567
rect 793 1493 807 1507
rect 833 1473 847 1487
rect 813 1413 827 1427
rect 793 1333 807 1347
rect 793 1293 807 1307
rect 893 1513 907 1527
rect 913 1493 927 1507
rect 853 1453 867 1467
rect 873 1453 887 1467
rect 833 1353 847 1367
rect 833 1333 847 1347
rect 833 1293 847 1307
rect 813 1273 827 1287
rect 793 1213 807 1227
rect 793 1193 807 1207
rect 673 1073 687 1087
rect 633 1013 647 1027
rect 733 1113 747 1127
rect 733 1073 747 1087
rect 773 1113 787 1127
rect 773 1073 787 1087
rect 773 1013 787 1027
rect 773 993 787 1007
rect 753 913 767 927
rect 693 873 707 887
rect 653 853 667 867
rect 693 853 707 867
rect 733 853 747 867
rect 693 833 707 847
rect 633 793 647 807
rect 673 793 687 807
rect 713 793 727 807
rect 473 733 487 747
rect 533 733 547 747
rect 553 733 567 747
rect 533 713 547 727
rect 453 653 467 667
rect 433 493 447 507
rect 433 473 447 487
rect 493 633 507 647
rect 473 613 487 627
rect 493 593 507 607
rect 473 513 487 527
rect 433 393 447 407
rect 453 393 467 407
rect 513 573 527 587
rect 533 573 547 587
rect 593 753 607 767
rect 613 693 627 707
rect 573 633 587 647
rect 553 553 567 567
rect 513 493 527 507
rect 493 473 507 487
rect 513 453 527 467
rect 393 353 407 367
rect 413 333 427 347
rect 453 373 467 387
rect 493 373 507 387
rect 613 653 627 667
rect 653 753 667 767
rect 633 633 647 647
rect 633 613 647 627
rect 693 773 707 787
rect 673 673 687 687
rect 753 813 767 827
rect 733 753 747 767
rect 713 633 727 647
rect 613 493 627 507
rect 533 413 547 427
rect 593 413 607 427
rect 353 313 367 327
rect 433 313 447 327
rect 473 313 487 327
rect 513 313 527 327
rect 473 293 487 307
rect 353 273 367 287
rect 353 253 367 267
rect 253 173 267 187
rect 313 173 327 187
rect 333 173 347 187
rect 293 153 307 167
rect 313 153 327 167
rect 413 233 427 247
rect 373 153 387 167
rect 273 133 287 147
rect 333 133 347 147
rect 33 113 47 127
rect 593 353 607 367
rect 553 253 567 267
rect 553 193 567 207
rect 433 173 447 187
rect 473 173 487 187
rect 533 173 547 187
rect 453 133 467 147
rect 493 153 507 167
rect 513 133 527 147
rect 693 533 707 547
rect 633 433 647 447
rect 653 393 667 407
rect 693 393 707 407
rect 633 313 647 327
rect 713 333 727 347
rect 693 313 707 327
rect 673 213 687 227
rect 613 193 627 207
rect 773 733 787 747
rect 853 1273 867 1287
rect 933 1413 947 1427
rect 953 1373 967 1387
rect 893 1353 907 1367
rect 853 1233 867 1247
rect 873 1233 887 1247
rect 853 1213 867 1227
rect 833 1153 847 1167
rect 833 1133 847 1147
rect 813 1113 827 1127
rect 853 1093 867 1107
rect 913 1333 927 1347
rect 993 1633 1007 1647
rect 1013 1593 1027 1607
rect 1073 1753 1087 1767
rect 1153 1853 1167 1867
rect 1153 1813 1167 1827
rect 1133 1773 1147 1787
rect 1013 1573 1027 1587
rect 1013 1553 1027 1567
rect 1053 1553 1067 1567
rect 993 1533 1007 1547
rect 1033 1533 1047 1547
rect 1173 1733 1187 1747
rect 1133 1653 1147 1667
rect 1113 1633 1127 1647
rect 1173 1593 1187 1607
rect 1193 1593 1207 1607
rect 1113 1573 1127 1587
rect 1153 1573 1167 1587
rect 1273 2053 1287 2067
rect 1313 2053 1327 2067
rect 1293 2013 1307 2027
rect 1233 1833 1247 1847
rect 1273 1833 1287 1847
rect 1293 1833 1307 1847
rect 1253 1813 1267 1827
rect 1293 1813 1307 1827
rect 1233 1753 1247 1767
rect 1293 1773 1307 1787
rect 1273 1733 1287 1747
rect 1253 1713 1267 1727
rect 1273 1693 1287 1707
rect 1253 1673 1267 1687
rect 1213 1573 1227 1587
rect 1233 1573 1247 1587
rect 1433 2413 1447 2427
rect 1533 2533 1547 2547
rect 1513 2513 1527 2527
rect 1553 2513 1567 2527
rect 1493 2373 1507 2387
rect 1473 2353 1487 2367
rect 1473 2333 1487 2347
rect 1413 2253 1427 2267
rect 1453 2253 1467 2267
rect 1373 2193 1387 2207
rect 1613 2813 1627 2827
rect 1693 3213 1707 3227
rect 1713 3213 1727 3227
rect 1713 3193 1727 3207
rect 1693 3153 1707 3167
rect 1653 3093 1667 3107
rect 1733 3133 1747 3147
rect 1733 3113 1747 3127
rect 1713 3073 1727 3087
rect 1653 2973 1667 2987
rect 1633 2773 1647 2787
rect 1633 2693 1647 2707
rect 1693 2993 1707 3007
rect 1853 3493 1867 3507
rect 1813 3453 1827 3467
rect 1853 3433 1867 3447
rect 1773 3393 1787 3407
rect 1793 3373 1807 3387
rect 1833 3293 1847 3307
rect 1813 3273 1827 3287
rect 1833 3253 1847 3267
rect 1913 3633 1927 3647
rect 1933 3613 1947 3627
rect 1893 3473 1907 3487
rect 1913 3473 1927 3487
rect 1893 3433 1907 3447
rect 1893 3253 1907 3267
rect 1793 3213 1807 3227
rect 1833 3213 1847 3227
rect 1873 3213 1887 3227
rect 1893 3213 1907 3227
rect 1833 3193 1847 3207
rect 1873 3193 1887 3207
rect 1773 3153 1787 3167
rect 1793 3153 1807 3167
rect 1753 3093 1767 3107
rect 1753 3033 1767 3047
rect 1813 3133 1827 3147
rect 1773 3013 1787 3027
rect 1813 3013 1827 3027
rect 1993 3593 2007 3607
rect 2153 3733 2167 3747
rect 1993 3493 2007 3507
rect 1953 3473 1967 3487
rect 1973 3473 1987 3487
rect 2013 3453 2027 3467
rect 1973 3373 1987 3387
rect 1933 3353 1947 3367
rect 1953 3273 1967 3287
rect 1973 3253 1987 3267
rect 1933 3213 1947 3227
rect 1913 3133 1927 3147
rect 1853 3093 1867 3107
rect 1873 3093 1887 3107
rect 1893 3033 1907 3047
rect 1873 3013 1887 3027
rect 1793 2993 1807 3007
rect 1833 2993 1847 3007
rect 1693 2913 1707 2927
rect 1693 2893 1707 2907
rect 1673 2873 1687 2887
rect 1693 2813 1707 2827
rect 1693 2673 1707 2687
rect 1653 2653 1667 2667
rect 1673 2633 1687 2647
rect 1653 2613 1667 2627
rect 1593 2593 1607 2607
rect 1633 2533 1647 2547
rect 1593 2513 1607 2527
rect 1593 2493 1607 2507
rect 1573 2333 1587 2347
rect 1553 2273 1567 2287
rect 1573 2253 1587 2267
rect 1573 2233 1587 2247
rect 1413 2093 1427 2107
rect 1373 2073 1387 2087
rect 1353 1973 1367 1987
rect 1433 2033 1447 2047
rect 1393 2013 1407 2027
rect 1533 2213 1547 2227
rect 1553 2073 1567 2087
rect 1493 2053 1507 2067
rect 1533 2033 1547 2047
rect 1513 1993 1527 2007
rect 1573 1993 1587 2007
rect 1393 1913 1407 1927
rect 1453 1913 1467 1927
rect 1313 1693 1327 1707
rect 1293 1673 1307 1687
rect 1373 1713 1387 1727
rect 1353 1653 1367 1667
rect 1313 1613 1327 1627
rect 1333 1613 1347 1627
rect 1373 1613 1387 1627
rect 1093 1553 1107 1567
rect 1153 1553 1167 1567
rect 1173 1553 1187 1567
rect 1213 1553 1227 1567
rect 993 1493 1007 1507
rect 1033 1433 1047 1447
rect 973 1353 987 1367
rect 973 1333 987 1347
rect 1013 1333 1027 1347
rect 1033 1333 1047 1347
rect 933 1313 947 1327
rect 913 1293 927 1307
rect 913 1273 927 1287
rect 993 1273 1007 1287
rect 893 1213 907 1227
rect 893 1153 907 1167
rect 993 1253 1007 1267
rect 993 1193 1007 1207
rect 973 1153 987 1167
rect 933 1113 947 1127
rect 1093 1353 1107 1367
rect 1073 1333 1087 1347
rect 1113 1333 1127 1347
rect 1093 1313 1107 1327
rect 1113 1313 1127 1327
rect 1093 1293 1107 1307
rect 1053 1253 1067 1267
rect 1053 1193 1067 1207
rect 1033 1173 1047 1187
rect 1033 1133 1047 1147
rect 1093 1153 1107 1167
rect 953 1073 967 1087
rect 873 1053 887 1067
rect 893 1053 907 1067
rect 813 1013 827 1027
rect 833 973 847 987
rect 813 913 827 927
rect 853 893 867 907
rect 833 853 847 867
rect 833 813 847 827
rect 853 813 867 827
rect 813 693 827 707
rect 793 673 807 687
rect 833 653 847 667
rect 813 633 827 647
rect 773 593 787 607
rect 773 533 787 547
rect 893 973 907 987
rect 993 953 1007 967
rect 893 933 907 947
rect 913 893 927 907
rect 893 853 907 867
rect 953 853 967 867
rect 973 853 987 867
rect 893 813 907 827
rect 973 813 987 827
rect 933 793 947 807
rect 873 773 887 787
rect 1053 1093 1067 1107
rect 1073 953 1087 967
rect 1073 933 1087 947
rect 1013 913 1027 927
rect 1073 873 1087 887
rect 1273 1553 1287 1567
rect 1193 1533 1207 1547
rect 1233 1533 1247 1547
rect 1253 1533 1267 1547
rect 1293 1513 1307 1527
rect 1333 1573 1347 1587
rect 1333 1553 1347 1567
rect 1233 1493 1247 1507
rect 1313 1493 1327 1507
rect 1193 1473 1207 1487
rect 1173 1433 1187 1447
rect 1253 1393 1267 1407
rect 1193 1373 1207 1387
rect 1173 1333 1187 1347
rect 1213 1353 1227 1367
rect 1193 1313 1207 1327
rect 1153 1293 1167 1307
rect 1193 1233 1207 1247
rect 1193 1213 1207 1227
rect 1133 1193 1147 1207
rect 1273 1333 1287 1347
rect 1173 1173 1187 1187
rect 1213 1173 1227 1187
rect 1133 1153 1147 1167
rect 1113 1133 1127 1147
rect 1113 1113 1127 1127
rect 1193 1153 1207 1167
rect 1153 1073 1167 1087
rect 1153 973 1167 987
rect 1173 953 1187 967
rect 1113 913 1127 927
rect 1013 853 1027 867
rect 1053 853 1067 867
rect 1093 853 1107 867
rect 1113 853 1127 867
rect 1053 833 1067 847
rect 1033 753 1047 767
rect 993 713 1007 727
rect 893 693 907 707
rect 953 693 967 707
rect 873 653 887 667
rect 853 633 867 647
rect 913 673 927 687
rect 1013 673 1027 687
rect 993 653 1007 667
rect 893 613 907 627
rect 933 613 947 627
rect 973 613 987 627
rect 853 593 867 607
rect 873 593 887 607
rect 893 573 907 587
rect 873 453 887 467
rect 873 413 887 427
rect 773 353 787 367
rect 853 393 867 407
rect 833 373 847 387
rect 973 433 987 447
rect 933 393 947 407
rect 893 373 907 387
rect 813 333 827 347
rect 753 293 767 307
rect 733 233 747 247
rect 793 313 807 327
rect 813 293 827 307
rect 953 353 967 367
rect 913 313 927 327
rect 953 273 967 287
rect 913 253 927 267
rect 893 233 907 247
rect 813 213 827 227
rect 853 213 867 227
rect 893 213 907 227
rect 633 173 647 187
rect 593 153 607 167
rect 753 173 767 187
rect 773 173 787 187
rect 793 173 807 187
rect 853 193 867 207
rect 733 153 747 167
rect 553 133 567 147
rect 593 113 607 127
rect 753 133 767 147
rect 793 133 807 147
rect 833 133 847 147
rect 653 113 667 127
rect 613 93 627 107
rect 833 93 847 107
rect 873 153 887 167
rect 1253 1293 1267 1307
rect 1253 1253 1267 1267
rect 1233 1133 1247 1147
rect 1233 1093 1247 1107
rect 1213 1073 1227 1087
rect 1253 953 1267 967
rect 1193 933 1207 947
rect 1193 913 1207 927
rect 1213 893 1227 907
rect 1433 1873 1447 1887
rect 1433 1813 1447 1827
rect 1533 1813 1547 1827
rect 1473 1793 1487 1807
rect 1533 1793 1547 1807
rect 1553 1793 1567 1807
rect 1413 1773 1427 1787
rect 1513 1773 1527 1787
rect 1493 1753 1507 1767
rect 1453 1733 1467 1747
rect 1473 1633 1487 1647
rect 1533 1633 1547 1647
rect 1573 1633 1587 1647
rect 1413 1573 1427 1587
rect 1413 1553 1427 1567
rect 1533 1613 1547 1627
rect 1653 2513 1667 2527
rect 1633 2373 1647 2387
rect 1613 2273 1627 2287
rect 1693 2553 1707 2567
rect 1673 2473 1687 2487
rect 1793 2933 1807 2947
rect 1753 2873 1767 2887
rect 1753 2793 1767 2807
rect 1773 2793 1787 2807
rect 1753 2733 1767 2747
rect 1833 2773 1847 2787
rect 1813 2753 1827 2767
rect 1853 2753 1867 2767
rect 1773 2673 1787 2687
rect 1833 2733 1847 2747
rect 1853 2733 1867 2747
rect 1853 2693 1867 2707
rect 1833 2653 1847 2667
rect 1793 2593 1807 2607
rect 1733 2553 1747 2567
rect 1653 2253 1667 2267
rect 1673 2213 1687 2227
rect 1813 2513 1827 2527
rect 1813 2493 1827 2507
rect 1793 2473 1807 2487
rect 1853 2473 1867 2487
rect 1993 3173 2007 3187
rect 2033 3273 2047 3287
rect 2133 3693 2147 3707
rect 2333 3733 2347 3747
rect 2153 3593 2167 3607
rect 2313 3713 2327 3727
rect 2313 3593 2327 3607
rect 2173 3573 2187 3587
rect 2173 3553 2187 3567
rect 2293 3553 2307 3567
rect 2113 3533 2127 3547
rect 2113 3513 2127 3527
rect 2153 3513 2167 3527
rect 2233 3513 2247 3527
rect 2113 3473 2127 3487
rect 2093 3453 2107 3467
rect 2093 3413 2107 3427
rect 2073 3253 2087 3267
rect 2253 3493 2267 3507
rect 2153 3333 2167 3347
rect 2133 3313 2147 3327
rect 2113 3253 2127 3267
rect 2133 3233 2147 3247
rect 2153 3233 2167 3247
rect 2033 3213 2047 3227
rect 2073 3213 2087 3227
rect 2113 3213 2127 3227
rect 1973 3133 1987 3147
rect 1953 3113 1967 3127
rect 1933 3053 1947 3067
rect 2073 3193 2087 3207
rect 1913 2833 1927 2847
rect 1893 2793 1907 2807
rect 1973 2993 1987 3007
rect 2033 3093 2047 3107
rect 2093 3073 2107 3087
rect 2153 3113 2167 3127
rect 2133 3073 2147 3087
rect 2113 3053 2127 3067
rect 2133 3033 2147 3047
rect 2273 3293 2287 3307
rect 2273 3273 2287 3287
rect 2213 3233 2227 3247
rect 2253 3233 2267 3247
rect 2333 3493 2347 3507
rect 2373 3913 2387 3927
rect 2373 3693 2387 3707
rect 2393 3653 2407 3667
rect 2373 3613 2387 3627
rect 2373 3533 2387 3547
rect 2613 3973 2627 3987
rect 2473 3893 2487 3907
rect 2473 3733 2487 3747
rect 2753 4113 2767 4127
rect 2973 4453 2987 4467
rect 3113 4493 3127 4507
rect 3133 4493 3147 4507
rect 3173 4513 3187 4527
rect 3233 4513 3247 4527
rect 3173 4493 3187 4507
rect 3413 4493 3427 4507
rect 3273 4473 3287 4487
rect 3353 4473 3367 4487
rect 3373 4473 3387 4487
rect 3033 4453 3047 4467
rect 3073 4453 3087 4467
rect 3113 4453 3127 4467
rect 3073 4433 3087 4447
rect 3013 4413 3027 4427
rect 2913 4213 2927 4227
rect 2873 4193 2887 4207
rect 2853 4153 2867 4167
rect 3013 4193 3027 4207
rect 3053 4193 3067 4207
rect 2933 4173 2947 4187
rect 2973 4173 2987 4187
rect 2953 4153 2967 4167
rect 2913 4133 2927 4147
rect 2953 4133 2967 4147
rect 2993 4133 3007 4147
rect 2713 4073 2727 4087
rect 2813 4073 2827 4087
rect 2733 4033 2747 4047
rect 2773 3993 2787 4007
rect 3253 4453 3267 4467
rect 3293 4453 3307 4467
rect 3393 4453 3407 4467
rect 3193 4413 3207 4427
rect 3193 4273 3207 4287
rect 3113 4253 3127 4267
rect 3093 4213 3107 4227
rect 3253 4253 3267 4267
rect 3113 4193 3127 4207
rect 3073 4153 3087 4167
rect 3093 4153 3107 4167
rect 3033 4113 3047 4127
rect 2993 4033 3007 4047
rect 3053 4013 3067 4027
rect 3073 4013 3087 4027
rect 3233 4213 3247 4227
rect 3213 4173 3227 4187
rect 3273 4233 3287 4247
rect 3393 4233 3407 4247
rect 3313 4213 3327 4227
rect 3293 4193 3307 4207
rect 3253 4153 3267 4167
rect 3333 4153 3347 4167
rect 3153 4113 3167 4127
rect 3373 4153 3387 4167
rect 3353 4053 3367 4067
rect 3233 4033 3247 4047
rect 3213 4013 3227 4027
rect 2673 3953 2687 3967
rect 2773 3953 2787 3967
rect 2633 3713 2647 3727
rect 2673 3713 2687 3727
rect 2493 3693 2507 3707
rect 2533 3693 2547 3707
rect 2453 3673 2467 3687
rect 2493 3573 2507 3587
rect 2433 3553 2447 3567
rect 2393 3493 2407 3507
rect 2353 3353 2367 3367
rect 2333 3293 2347 3307
rect 2393 3293 2407 3307
rect 2293 3253 2307 3267
rect 2353 3273 2367 3287
rect 2193 3213 2207 3227
rect 2233 3213 2247 3227
rect 2273 3213 2287 3227
rect 2173 3093 2187 3107
rect 2273 3073 2287 3087
rect 2193 3033 2207 3047
rect 2233 3033 2247 3047
rect 2053 3013 2067 3027
rect 2073 3013 2087 3027
rect 2113 3013 2127 3027
rect 2153 3013 2167 3027
rect 2213 3013 2227 3027
rect 2073 2993 2087 3007
rect 2013 2953 2027 2967
rect 2013 2793 2027 2807
rect 2053 2793 2067 2807
rect 1973 2773 1987 2787
rect 1893 2753 1907 2767
rect 1933 2753 1947 2767
rect 1993 2733 2007 2747
rect 1893 2713 1907 2727
rect 1913 2673 1927 2687
rect 1953 2693 1967 2707
rect 1933 2553 1947 2567
rect 1893 2493 1907 2507
rect 1773 2413 1787 2427
rect 1813 2453 1827 2467
rect 1793 2253 1807 2267
rect 1833 2233 1847 2247
rect 1873 2213 1887 2227
rect 1713 2193 1727 2207
rect 1813 2193 1827 2207
rect 1633 2173 1647 2187
rect 1693 2173 1707 2187
rect 1773 2173 1787 2187
rect 1693 2153 1707 2167
rect 1653 2113 1667 2127
rect 1753 2133 1767 2147
rect 1733 2093 1747 2107
rect 1753 2093 1767 2107
rect 1693 2073 1707 2087
rect 1813 2153 1827 2167
rect 1833 2153 1847 2167
rect 1873 2153 1887 2167
rect 1853 2093 1867 2107
rect 1633 2053 1647 2067
rect 1673 2053 1687 2067
rect 1713 2053 1727 2067
rect 1733 2053 1747 2067
rect 1753 2053 1767 2067
rect 1653 1973 1667 1987
rect 1613 1813 1627 1827
rect 1633 1793 1647 1807
rect 1633 1753 1647 1767
rect 1613 1673 1627 1687
rect 1593 1613 1607 1627
rect 1493 1573 1507 1587
rect 1513 1553 1527 1567
rect 1433 1493 1447 1507
rect 1453 1493 1467 1507
rect 1413 1473 1427 1487
rect 1433 1413 1447 1427
rect 1393 1393 1407 1407
rect 1413 1393 1427 1407
rect 1373 1353 1387 1367
rect 1393 1353 1407 1367
rect 1333 1313 1347 1327
rect 1293 1293 1307 1307
rect 1313 1273 1327 1287
rect 1333 1253 1347 1267
rect 1293 1133 1307 1147
rect 1293 1113 1307 1127
rect 1313 1053 1327 1067
rect 1293 1013 1307 1027
rect 1213 873 1227 887
rect 1273 873 1287 887
rect 1313 913 1327 927
rect 1193 833 1207 847
rect 1093 813 1107 827
rect 1093 793 1107 807
rect 1073 773 1087 787
rect 1033 653 1047 667
rect 1053 653 1067 667
rect 1013 633 1027 647
rect 1013 613 1027 627
rect 1133 753 1147 767
rect 1253 833 1267 847
rect 1293 833 1307 847
rect 1373 1253 1387 1267
rect 1353 1193 1367 1207
rect 1353 1133 1367 1147
rect 1393 1213 1407 1227
rect 1373 1113 1387 1127
rect 1493 1473 1507 1487
rect 1473 1373 1487 1387
rect 1453 1333 1467 1347
rect 1433 1313 1447 1327
rect 1513 1433 1527 1447
rect 1493 1353 1507 1367
rect 1613 1593 1627 1607
rect 1553 1573 1567 1587
rect 1573 1573 1587 1587
rect 1733 2013 1747 2027
rect 2053 2693 2067 2707
rect 2033 2673 2047 2687
rect 2253 2833 2267 2847
rect 2233 2793 2247 2807
rect 2213 2773 2227 2787
rect 2153 2753 2167 2767
rect 2133 2733 2147 2747
rect 2333 3233 2347 3247
rect 2333 3193 2347 3207
rect 2393 3213 2407 3227
rect 2373 3133 2387 3147
rect 2353 3093 2367 3107
rect 2293 3033 2307 3047
rect 2353 3033 2367 3047
rect 2433 3533 2447 3547
rect 2453 3213 2467 3227
rect 2453 3173 2467 3187
rect 2453 3073 2467 3087
rect 2433 3053 2447 3067
rect 2313 3013 2327 3027
rect 2373 3013 2387 3027
rect 2413 3013 2427 3027
rect 2293 2993 2307 3007
rect 2333 2993 2347 3007
rect 2393 2993 2407 3007
rect 2353 2773 2367 2787
rect 2273 2753 2287 2767
rect 2333 2753 2347 2767
rect 2093 2713 2107 2727
rect 2193 2713 2207 2727
rect 2253 2713 2267 2727
rect 2273 2693 2287 2707
rect 2313 2713 2327 2727
rect 2093 2673 2107 2687
rect 2113 2673 2127 2687
rect 2293 2673 2307 2687
rect 2073 2633 2087 2647
rect 1973 2573 1987 2587
rect 2073 2573 2087 2587
rect 2273 2653 2287 2667
rect 2193 2633 2207 2647
rect 2133 2573 2147 2587
rect 2253 2573 2267 2587
rect 2113 2553 2127 2567
rect 2013 2533 2027 2547
rect 2093 2533 2107 2547
rect 1993 2513 2007 2527
rect 2053 2513 2067 2527
rect 2033 2493 2047 2507
rect 1953 2473 1967 2487
rect 2033 2473 2047 2487
rect 1933 2413 1947 2427
rect 1973 2293 1987 2307
rect 1913 2273 1927 2287
rect 1973 2273 1987 2287
rect 2013 2273 2027 2287
rect 1913 2233 1927 2247
rect 1953 2213 1967 2227
rect 1933 2193 1947 2207
rect 1933 2153 1947 2167
rect 1893 2113 1907 2127
rect 1913 2113 1927 2127
rect 1993 2173 2007 2187
rect 1973 2113 1987 2127
rect 1933 2093 1947 2107
rect 1953 2093 1967 2107
rect 1913 2073 1927 2087
rect 2293 2633 2307 2647
rect 2173 2533 2187 2547
rect 2193 2533 2207 2547
rect 2213 2533 2227 2547
rect 2093 2453 2107 2467
rect 2073 2293 2087 2307
rect 2053 2133 2067 2147
rect 2053 2113 2067 2127
rect 2033 2073 2047 2087
rect 1953 2053 1967 2067
rect 2153 2413 2167 2427
rect 2113 2213 2127 2227
rect 2113 2073 2127 2087
rect 2253 2353 2267 2367
rect 2273 2313 2287 2327
rect 2213 2273 2227 2287
rect 2253 2273 2267 2287
rect 2193 2213 2207 2227
rect 2173 2173 2187 2187
rect 2153 2133 2167 2147
rect 1933 2033 1947 2047
rect 1893 2013 1907 2027
rect 1873 1993 1887 2007
rect 1713 1893 1727 1907
rect 1753 1893 1767 1907
rect 1713 1833 1727 1847
rect 1673 1813 1687 1827
rect 1653 1733 1667 1747
rect 1793 1813 1807 1827
rect 1913 1973 1927 1987
rect 1713 1793 1727 1807
rect 1733 1773 1747 1787
rect 1693 1693 1707 1707
rect 1673 1613 1687 1627
rect 1553 1453 1567 1467
rect 1533 1413 1547 1427
rect 1553 1393 1567 1407
rect 1513 1333 1527 1347
rect 1533 1313 1547 1327
rect 1453 1293 1467 1307
rect 1493 1273 1507 1287
rect 1533 1253 1547 1267
rect 1553 1253 1567 1267
rect 1413 1113 1427 1127
rect 1433 1113 1447 1127
rect 1353 1073 1367 1087
rect 1373 1073 1387 1087
rect 1413 1073 1427 1087
rect 1353 913 1367 927
rect 1393 1053 1407 1067
rect 1513 1153 1527 1167
rect 1473 1113 1487 1127
rect 1493 1093 1507 1107
rect 1453 1073 1467 1087
rect 1473 1073 1487 1087
rect 1433 973 1447 987
rect 1433 913 1447 927
rect 1393 893 1407 907
rect 1373 873 1387 887
rect 1333 853 1347 867
rect 1373 853 1387 867
rect 1333 833 1347 847
rect 1413 833 1427 847
rect 1293 773 1307 787
rect 1273 753 1287 767
rect 1233 733 1247 747
rect 1233 713 1247 727
rect 1353 793 1367 807
rect 1393 753 1407 767
rect 1413 753 1427 767
rect 1193 693 1207 707
rect 1113 673 1127 687
rect 1053 633 1067 647
rect 1093 633 1107 647
rect 1133 633 1147 647
rect 1313 693 1327 707
rect 1333 693 1347 707
rect 1273 673 1287 687
rect 1073 613 1087 627
rect 1113 613 1127 627
rect 1073 593 1087 607
rect 993 413 1007 427
rect 1173 613 1187 627
rect 1213 613 1227 627
rect 1253 613 1267 627
rect 1113 533 1127 547
rect 1153 533 1167 547
rect 1073 493 1087 507
rect 1213 493 1227 507
rect 1133 413 1147 427
rect 1013 353 1027 367
rect 1113 373 1127 387
rect 1173 393 1187 407
rect 993 313 1007 327
rect 1053 313 1067 327
rect 953 193 967 207
rect 913 153 927 167
rect 1033 293 1047 307
rect 1013 213 1027 227
rect 973 173 987 187
rect 993 173 1007 187
rect 1133 353 1147 367
rect 1353 673 1367 687
rect 1453 893 1467 907
rect 1433 733 1447 747
rect 1433 673 1447 687
rect 1373 633 1387 647
rect 1413 633 1427 647
rect 1673 1573 1687 1587
rect 1693 1573 1707 1587
rect 1633 1553 1647 1567
rect 1793 1793 1807 1807
rect 1773 1753 1787 1767
rect 1813 1773 1827 1787
rect 1853 1773 1867 1787
rect 1993 2013 2007 2027
rect 1933 1813 1947 1827
rect 1753 1593 1767 1607
rect 1833 1753 1847 1767
rect 1833 1713 1847 1727
rect 1853 1653 1867 1667
rect 1833 1613 1847 1627
rect 1813 1593 1827 1607
rect 1833 1593 1847 1607
rect 1753 1553 1767 1567
rect 1613 1513 1627 1527
rect 1593 1493 1607 1507
rect 1693 1473 1707 1487
rect 1673 1353 1687 1367
rect 1613 1313 1627 1327
rect 1593 1293 1607 1307
rect 1573 1233 1587 1247
rect 1573 1173 1587 1187
rect 1553 1113 1567 1127
rect 1553 1093 1567 1107
rect 1573 1033 1587 1047
rect 1533 993 1547 1007
rect 1493 973 1507 987
rect 1533 933 1547 947
rect 1613 1193 1627 1207
rect 1653 1273 1667 1287
rect 1633 1173 1647 1187
rect 1733 1393 1747 1407
rect 1793 1553 1807 1567
rect 1833 1553 1847 1567
rect 1773 1533 1787 1547
rect 1793 1473 1807 1487
rect 1953 1633 1967 1647
rect 1913 1613 1927 1627
rect 1933 1613 1947 1627
rect 1873 1593 1887 1607
rect 1913 1573 1927 1587
rect 1893 1553 1907 1567
rect 1853 1533 1867 1547
rect 1833 1393 1847 1407
rect 1853 1393 1867 1407
rect 1753 1333 1767 1347
rect 1693 1293 1707 1307
rect 1773 1313 1787 1327
rect 1813 1313 1827 1327
rect 1713 1273 1727 1287
rect 1793 1273 1807 1287
rect 1693 1253 1707 1267
rect 1773 1193 1787 1207
rect 1693 1153 1707 1167
rect 1613 1133 1627 1147
rect 1633 1133 1647 1147
rect 1673 1133 1687 1147
rect 1693 1133 1707 1147
rect 1673 1113 1687 1127
rect 1613 1073 1627 1087
rect 1653 1073 1667 1087
rect 1753 1113 1767 1127
rect 1713 1093 1727 1107
rect 1733 1073 1747 1087
rect 1613 1053 1627 1067
rect 1633 1013 1647 1027
rect 1613 913 1627 927
rect 1473 853 1487 867
rect 1553 873 1567 887
rect 1593 873 1607 887
rect 1533 853 1547 867
rect 1573 853 1587 867
rect 1553 833 1567 847
rect 1553 813 1567 827
rect 1593 813 1607 827
rect 1493 773 1507 787
rect 1473 733 1487 747
rect 1453 653 1467 667
rect 1493 693 1507 707
rect 1293 613 1307 627
rect 1373 593 1387 607
rect 1353 513 1367 527
rect 1273 433 1287 447
rect 1353 433 1367 447
rect 1533 673 1547 687
rect 1513 653 1527 667
rect 1453 593 1467 607
rect 1413 573 1427 587
rect 1493 533 1507 547
rect 1513 533 1527 547
rect 1753 1033 1767 1047
rect 1653 993 1667 1007
rect 1753 973 1767 987
rect 1653 933 1667 947
rect 1633 893 1647 907
rect 1653 893 1667 907
rect 1733 873 1747 887
rect 1673 833 1687 847
rect 1613 753 1627 767
rect 1713 813 1727 827
rect 1713 793 1727 807
rect 1713 773 1727 787
rect 1693 713 1707 727
rect 1653 693 1667 707
rect 1833 1253 1847 1267
rect 1953 1573 1967 1587
rect 1933 1373 1947 1387
rect 1913 1353 1927 1367
rect 1873 1293 1887 1307
rect 1853 1213 1867 1227
rect 1793 1133 1807 1147
rect 1853 1133 1867 1147
rect 1813 1093 1827 1107
rect 1933 1333 1947 1347
rect 1913 1313 1927 1327
rect 1893 1273 1907 1287
rect 1873 1113 1887 1127
rect 1933 1293 1947 1307
rect 2013 1993 2027 2007
rect 2093 2053 2107 2067
rect 2253 2253 2267 2267
rect 2333 2573 2347 2587
rect 2313 2533 2327 2547
rect 2333 2513 2347 2527
rect 2453 3013 2467 3027
rect 2473 3013 2487 3027
rect 2453 2973 2467 2987
rect 2613 3693 2627 3707
rect 2713 3693 2727 3707
rect 2653 3673 2667 3687
rect 2673 3673 2687 3687
rect 2753 3673 2767 3687
rect 2593 3653 2607 3667
rect 2573 3553 2587 3567
rect 2533 3533 2547 3547
rect 2753 3653 2767 3667
rect 2913 3973 2927 3987
rect 3093 3993 3107 4007
rect 2973 3973 2987 3987
rect 3013 3973 3027 3987
rect 3153 3973 3167 3987
rect 2933 3953 2947 3967
rect 2873 3693 2887 3707
rect 2913 3693 2927 3707
rect 2793 3673 2807 3687
rect 2893 3673 2907 3687
rect 2813 3633 2827 3647
rect 2773 3613 2787 3627
rect 2913 3613 2927 3627
rect 2713 3553 2727 3567
rect 2513 3353 2527 3367
rect 2673 3513 2687 3527
rect 2693 3493 2707 3507
rect 2733 3493 2747 3507
rect 2553 3193 2567 3207
rect 2513 3113 2527 3127
rect 2513 3033 2527 3047
rect 2673 3153 2687 3167
rect 2633 3133 2647 3147
rect 2613 3053 2627 3067
rect 2533 3013 2547 3027
rect 2533 2993 2547 3007
rect 2493 2813 2507 2827
rect 2473 2793 2487 2807
rect 2493 2793 2507 2807
rect 2433 2773 2447 2787
rect 2473 2773 2487 2787
rect 2373 2753 2387 2767
rect 2413 2753 2427 2767
rect 2433 2733 2447 2747
rect 2393 2633 2407 2647
rect 2373 2593 2387 2607
rect 2453 2693 2467 2707
rect 2393 2553 2407 2567
rect 2473 2573 2487 2587
rect 2513 2733 2527 2747
rect 2593 2973 2607 2987
rect 2813 3513 2827 3527
rect 2833 3513 2847 3527
rect 2873 3493 2887 3507
rect 2893 3473 2907 3487
rect 2753 3413 2767 3427
rect 2713 3173 2727 3187
rect 2713 3093 2727 3107
rect 2773 3213 2787 3227
rect 2833 3213 2847 3227
rect 2773 3153 2787 3167
rect 2753 3053 2767 3067
rect 2653 3033 2667 3047
rect 2673 3033 2687 3047
rect 2693 3033 2707 3047
rect 2713 3013 2727 3027
rect 2633 2793 2647 2807
rect 2553 2773 2567 2787
rect 2593 2773 2607 2787
rect 2553 2733 2567 2747
rect 2573 2733 2587 2747
rect 2633 2753 2647 2767
rect 2733 2993 2747 3007
rect 2793 3053 2807 3067
rect 2773 2853 2787 2867
rect 2733 2753 2747 2767
rect 2773 2753 2787 2767
rect 2533 2693 2547 2707
rect 2513 2653 2527 2667
rect 2493 2553 2507 2567
rect 2373 2533 2387 2547
rect 2413 2533 2427 2547
rect 2753 2733 2767 2747
rect 2653 2713 2667 2727
rect 2713 2713 2727 2727
rect 2853 3193 2867 3207
rect 2893 3153 2907 3167
rect 2853 3093 2867 3107
rect 2873 3093 2887 3107
rect 2893 3093 2907 3107
rect 2853 3073 2867 3087
rect 2833 2993 2847 3007
rect 2813 2793 2827 2807
rect 2853 2773 2867 2787
rect 2833 2753 2847 2767
rect 3133 3953 3147 3967
rect 3173 3933 3187 3947
rect 3153 3753 3167 3767
rect 3273 4013 3287 4027
rect 3313 4013 3327 4027
rect 3333 4013 3347 4027
rect 3253 3973 3267 3987
rect 2973 3713 2987 3727
rect 2953 3673 2967 3687
rect 2953 3653 2967 3667
rect 2993 3633 3007 3647
rect 3153 3713 3167 3727
rect 3073 3673 3087 3687
rect 3113 3653 3127 3667
rect 3133 3633 3147 3647
rect 3053 3593 3067 3607
rect 3213 3713 3227 3727
rect 3193 3673 3207 3687
rect 3173 3573 3187 3587
rect 3213 3553 3227 3567
rect 3273 3733 3287 3747
rect 3353 3993 3367 4007
rect 3373 3993 3387 4007
rect 3353 3953 3367 3967
rect 3373 3953 3387 3967
rect 3273 3713 3287 3727
rect 3293 3713 3307 3727
rect 3313 3713 3327 3727
rect 3333 3713 3347 3727
rect 3493 4513 3507 4527
rect 3453 4473 3467 4487
rect 3633 4493 3647 4507
rect 3493 4233 3507 4247
rect 3493 4173 3507 4187
rect 3573 4473 3587 4487
rect 3613 4213 3627 4227
rect 3433 4153 3447 4167
rect 3613 4173 3627 4187
rect 3553 4093 3567 4107
rect 3533 4073 3547 4087
rect 3453 4013 3467 4027
rect 3473 4013 3487 4027
rect 3413 3993 3427 4007
rect 3433 3993 3447 4007
rect 3393 3733 3407 3747
rect 3253 3693 3267 3707
rect 3373 3673 3387 3687
rect 3353 3653 3367 3667
rect 3293 3613 3307 3627
rect 3273 3553 3287 3567
rect 3353 3553 3367 3567
rect 3033 3533 3047 3547
rect 3153 3533 3167 3547
rect 3213 3533 3227 3547
rect 3233 3533 3247 3547
rect 2933 3513 2947 3527
rect 3073 3513 3087 3527
rect 3133 3513 3147 3527
rect 2953 3473 2967 3487
rect 2993 3453 3007 3467
rect 2953 3233 2967 3247
rect 2973 3213 2987 3227
rect 2973 3113 2987 3127
rect 3093 3273 3107 3287
rect 3173 3513 3187 3527
rect 3253 3513 3267 3527
rect 3193 3493 3207 3507
rect 3233 3493 3247 3507
rect 3173 3473 3187 3487
rect 3233 3453 3247 3467
rect 3153 3313 3167 3327
rect 3313 3533 3327 3547
rect 3333 3533 3347 3547
rect 3393 3633 3407 3647
rect 3513 3973 3527 3987
rect 3573 3933 3587 3947
rect 3713 4473 3727 4487
rect 3693 4453 3707 4467
rect 3733 4453 3747 4467
rect 3793 4453 3807 4467
rect 3653 4433 3667 4447
rect 3773 4433 3787 4447
rect 3793 4413 3807 4427
rect 3653 4233 3667 4247
rect 3713 4233 3727 4247
rect 3673 4213 3687 4227
rect 3653 4153 3667 4167
rect 3773 4173 3787 4187
rect 3733 4153 3747 4167
rect 3693 4093 3707 4107
rect 3653 4073 3667 4087
rect 3673 4033 3687 4047
rect 3773 4153 3787 4167
rect 3753 4013 3767 4027
rect 3693 3993 3707 4007
rect 3673 3953 3687 3967
rect 3633 3913 3647 3927
rect 3773 3893 3787 3907
rect 3673 3833 3687 3847
rect 3513 3753 3527 3767
rect 3613 3753 3627 3767
rect 3433 3673 3447 3687
rect 3453 3653 3467 3667
rect 3413 3613 3427 3627
rect 3433 3613 3447 3627
rect 3393 3553 3407 3567
rect 3413 3533 3427 3547
rect 3433 3533 3447 3547
rect 3393 3493 3407 3507
rect 3433 3493 3447 3507
rect 3293 3473 3307 3487
rect 3293 3393 3307 3407
rect 3273 3293 3287 3307
rect 3213 3273 3227 3287
rect 3133 3253 3147 3267
rect 3013 3233 3027 3247
rect 3053 3233 3067 3247
rect 3093 3233 3107 3247
rect 3033 3213 3047 3227
rect 3033 3193 3047 3207
rect 3153 3233 3167 3247
rect 3113 3213 3127 3227
rect 3133 3213 3147 3227
rect 3093 3193 3107 3207
rect 3173 3193 3187 3207
rect 3073 3173 3087 3187
rect 3053 3053 3067 3067
rect 3113 3073 3127 3087
rect 3153 3073 3167 3087
rect 3093 3053 3107 3067
rect 3033 3033 3047 3047
rect 3073 3033 3087 3047
rect 2993 2993 3007 3007
rect 3033 2993 3047 3007
rect 2973 2973 2987 2987
rect 2993 2853 3007 2867
rect 2953 2833 2967 2847
rect 2913 2773 2927 2787
rect 2873 2713 2887 2727
rect 2713 2693 2727 2707
rect 2793 2693 2807 2707
rect 2633 2673 2647 2687
rect 2693 2593 2707 2607
rect 2573 2513 2587 2527
rect 2553 2493 2567 2507
rect 2573 2493 2587 2507
rect 2513 2333 2527 2347
rect 2353 2293 2367 2307
rect 2393 2293 2407 2307
rect 2513 2293 2527 2307
rect 2553 2293 2567 2307
rect 2373 2273 2387 2287
rect 2293 2253 2307 2267
rect 2313 2253 2327 2267
rect 2273 2233 2287 2247
rect 2353 2233 2367 2247
rect 2373 2233 2387 2247
rect 2253 2213 2267 2227
rect 2233 2153 2247 2167
rect 2213 2113 2227 2127
rect 2073 1933 2087 1947
rect 2093 1933 2107 1947
rect 2153 1933 2167 1947
rect 2073 1813 2087 1827
rect 2033 1633 2047 1647
rect 2013 1613 2027 1627
rect 2233 1973 2247 1987
rect 2193 1853 2207 1867
rect 2153 1833 2167 1847
rect 2133 1773 2147 1787
rect 2193 1813 2207 1827
rect 2293 2133 2307 2147
rect 2273 2093 2287 2107
rect 2273 1833 2287 1847
rect 2173 1793 2187 1807
rect 2253 1793 2267 1807
rect 2273 1793 2287 1807
rect 2153 1633 2167 1647
rect 2193 1773 2207 1787
rect 2153 1613 2167 1627
rect 2173 1613 2187 1627
rect 2213 1753 2227 1767
rect 2013 1593 2027 1607
rect 2093 1593 2107 1607
rect 2193 1593 2207 1607
rect 2333 2053 2347 2067
rect 2433 2273 2447 2287
rect 2473 2273 2487 2287
rect 2413 2253 2427 2267
rect 2533 2273 2547 2287
rect 2673 2553 2687 2567
rect 2693 2533 2707 2547
rect 2833 2573 2847 2587
rect 2853 2573 2867 2587
rect 2893 2573 2907 2587
rect 2733 2553 2747 2567
rect 2793 2553 2807 2567
rect 2773 2533 2787 2547
rect 2793 2513 2807 2527
rect 2853 2513 2867 2527
rect 2653 2493 2667 2507
rect 2713 2493 2727 2507
rect 2813 2493 2827 2507
rect 2873 2493 2887 2507
rect 2633 2353 2647 2367
rect 2613 2313 2627 2327
rect 2613 2293 2627 2307
rect 2673 2333 2687 2347
rect 2573 2253 2587 2267
rect 2453 2193 2467 2207
rect 2393 2093 2407 2107
rect 2413 2053 2427 2067
rect 2533 2233 2547 2247
rect 2613 2233 2627 2247
rect 2533 2153 2547 2167
rect 2593 2153 2607 2167
rect 2373 1973 2387 1987
rect 2513 1953 2527 1967
rect 2393 1933 2407 1947
rect 2393 1853 2407 1867
rect 2353 1833 2367 1847
rect 2333 1813 2347 1827
rect 2333 1793 2347 1807
rect 2373 1793 2387 1807
rect 2293 1713 2307 1727
rect 2053 1573 2067 1587
rect 2113 1573 2127 1587
rect 1973 1553 1987 1567
rect 1993 1553 2007 1567
rect 2033 1553 2047 1567
rect 2093 1553 2107 1567
rect 2233 1573 2247 1587
rect 2353 1733 2367 1747
rect 2353 1633 2367 1647
rect 2173 1553 2187 1567
rect 2333 1553 2347 1567
rect 2113 1533 2127 1547
rect 2053 1373 2067 1387
rect 2093 1373 2107 1387
rect 1993 1333 2007 1347
rect 1993 1313 2007 1327
rect 2033 1313 2047 1327
rect 1973 1273 1987 1287
rect 1933 1253 1947 1267
rect 1953 1253 1967 1267
rect 1893 1093 1907 1107
rect 1873 1073 1887 1087
rect 1913 1073 1927 1087
rect 2013 1233 2027 1247
rect 2013 1213 2027 1227
rect 1793 1053 1807 1067
rect 1833 1053 1847 1067
rect 1933 1053 1947 1067
rect 1813 1033 1827 1047
rect 1793 973 1807 987
rect 1773 933 1787 947
rect 1753 853 1767 867
rect 1753 813 1767 827
rect 1773 813 1787 827
rect 1733 753 1747 767
rect 1813 953 1827 967
rect 1953 1033 1967 1047
rect 1893 1013 1907 1027
rect 1833 913 1847 927
rect 1833 873 1847 887
rect 1873 853 1887 867
rect 1933 893 1947 907
rect 1933 873 1947 887
rect 2473 1833 2487 1847
rect 2413 1753 2427 1767
rect 2413 1733 2427 1747
rect 2453 1733 2467 1747
rect 2573 2093 2587 2107
rect 2553 2073 2567 2087
rect 2653 2213 2667 2227
rect 2793 2253 2807 2267
rect 2693 2193 2707 2207
rect 2673 2153 2687 2167
rect 2653 2133 2667 2147
rect 2673 2073 2687 2087
rect 2713 2053 2727 2067
rect 2773 2053 2787 2067
rect 2673 2033 2687 2047
rect 2733 2033 2747 2047
rect 2753 2033 2767 2047
rect 2793 2033 2807 2047
rect 2613 1993 2627 2007
rect 2693 1993 2707 2007
rect 2653 1973 2667 1987
rect 2493 1773 2507 1787
rect 2533 1773 2547 1787
rect 2493 1753 2507 1767
rect 2473 1673 2487 1687
rect 2433 1633 2447 1647
rect 2433 1613 2447 1627
rect 2373 1533 2387 1547
rect 2193 1333 2207 1347
rect 2153 1313 2167 1327
rect 2173 1313 2187 1327
rect 2153 1293 2167 1307
rect 2073 1273 2087 1287
rect 2133 1273 2147 1287
rect 2093 1253 2107 1267
rect 2053 1133 2067 1147
rect 2133 1233 2147 1247
rect 2133 1113 2147 1127
rect 2273 1333 2287 1347
rect 2353 1333 2367 1347
rect 2253 1293 2267 1307
rect 2333 1293 2347 1307
rect 2213 1233 2227 1247
rect 2213 1133 2227 1147
rect 2113 1093 2127 1107
rect 2153 1093 2167 1107
rect 2193 1093 2207 1107
rect 2073 1073 2087 1087
rect 2173 1073 2187 1087
rect 2353 1133 2367 1147
rect 2393 1113 2407 1127
rect 2273 1073 2287 1087
rect 2373 1093 2387 1107
rect 2033 1053 2047 1067
rect 2253 1053 2267 1067
rect 2313 1053 2327 1067
rect 2013 1013 2027 1027
rect 1993 873 2007 887
rect 1973 853 1987 867
rect 1813 813 1827 827
rect 1793 793 1807 807
rect 1853 773 1867 787
rect 1833 753 1847 767
rect 1753 733 1767 747
rect 1593 673 1607 687
rect 1593 653 1607 667
rect 1653 653 1667 667
rect 1733 673 1747 687
rect 1713 653 1727 667
rect 1593 613 1607 627
rect 1573 593 1587 607
rect 1393 453 1407 467
rect 1353 413 1367 427
rect 1373 413 1387 427
rect 1253 373 1267 387
rect 1273 373 1287 387
rect 1333 373 1347 387
rect 1313 353 1327 367
rect 1153 333 1167 347
rect 1113 313 1127 327
rect 1173 313 1187 327
rect 1133 293 1147 307
rect 1093 213 1107 227
rect 1113 213 1127 227
rect 1033 193 1047 207
rect 1073 193 1087 207
rect 1093 153 1107 167
rect 1233 333 1247 347
rect 1253 333 1267 347
rect 1253 293 1267 307
rect 1193 273 1207 287
rect 1273 233 1287 247
rect 1213 193 1227 207
rect 933 133 947 147
rect 973 133 987 147
rect 1053 133 1067 147
rect 1113 133 1127 147
rect 873 113 887 127
rect 993 113 1007 127
rect 1193 133 1207 147
rect 973 73 987 87
rect 1233 133 1247 147
rect 1453 393 1467 407
rect 1353 353 1367 367
rect 1393 353 1407 367
rect 1333 273 1347 287
rect 1413 333 1427 347
rect 1413 313 1427 327
rect 1373 253 1387 267
rect 1393 253 1407 267
rect 1473 333 1487 347
rect 1453 313 1467 327
rect 1473 313 1487 327
rect 1433 273 1447 287
rect 1373 233 1387 247
rect 1413 233 1427 247
rect 1293 193 1307 207
rect 1313 173 1327 187
rect 1253 113 1267 127
rect 1293 113 1307 127
rect 1213 53 1227 67
rect 853 33 867 47
rect 1333 153 1347 167
rect 1433 173 1447 187
rect 1433 153 1447 167
rect 1493 293 1507 307
rect 1473 253 1487 267
rect 1533 513 1547 527
rect 1553 513 1567 527
rect 1773 653 1787 667
rect 1813 653 1827 667
rect 1753 613 1767 627
rect 1673 573 1687 587
rect 1653 533 1667 547
rect 1593 513 1607 527
rect 1633 513 1647 527
rect 1593 433 1607 447
rect 1553 373 1567 387
rect 1573 373 1587 387
rect 1533 353 1547 367
rect 1533 273 1547 287
rect 1633 393 1647 407
rect 1653 393 1667 407
rect 1713 593 1727 607
rect 1753 593 1767 607
rect 1773 573 1787 587
rect 1693 513 1707 527
rect 1733 493 1747 507
rect 1713 473 1727 487
rect 1693 413 1707 427
rect 1713 413 1727 427
rect 1673 373 1687 387
rect 1913 793 1927 807
rect 1953 793 1967 807
rect 1933 773 1947 787
rect 1873 673 1887 687
rect 1833 593 1847 607
rect 1813 533 1827 547
rect 1853 573 1867 587
rect 1893 573 1907 587
rect 1833 513 1847 527
rect 1833 493 1847 507
rect 1773 473 1787 487
rect 1793 473 1807 487
rect 1813 393 1827 407
rect 1633 353 1647 367
rect 1673 353 1687 367
rect 1713 353 1727 367
rect 1753 353 1767 367
rect 1593 273 1607 287
rect 1573 253 1587 267
rect 1733 333 1747 347
rect 1673 313 1687 327
rect 1693 313 1707 327
rect 1653 253 1667 267
rect 1633 233 1647 247
rect 1693 293 1707 307
rect 1753 293 1767 307
rect 1533 193 1547 207
rect 1613 193 1627 207
rect 1493 173 1507 187
rect 1513 173 1527 187
rect 1553 153 1567 167
rect 1433 133 1447 147
rect 1473 133 1487 147
rect 1533 133 1547 147
rect 1353 113 1367 127
rect 1513 113 1527 127
rect 1573 133 1587 147
rect 1613 133 1627 147
rect 1693 233 1707 247
rect 1673 173 1687 187
rect 1693 173 1707 187
rect 1733 173 1747 187
rect 1873 453 1887 467
rect 1913 453 1927 467
rect 1853 433 1867 447
rect 1913 433 1927 447
rect 1893 413 1907 427
rect 1873 353 1887 367
rect 1913 393 1927 407
rect 2153 933 2167 947
rect 2053 833 2067 847
rect 2013 793 2027 807
rect 1993 773 2007 787
rect 1993 753 2007 767
rect 1973 733 1987 747
rect 1953 713 1967 727
rect 2053 773 2067 787
rect 2033 713 2047 727
rect 2013 653 2027 667
rect 2053 693 2067 707
rect 2133 833 2147 847
rect 2093 693 2107 707
rect 2133 733 2147 747
rect 2113 653 2127 667
rect 2113 633 2127 647
rect 1993 613 2007 627
rect 1973 593 1987 607
rect 2013 533 2027 547
rect 2033 533 2047 547
rect 1993 473 2007 487
rect 1953 393 1967 407
rect 1933 373 1947 387
rect 2093 613 2107 627
rect 2113 593 2127 607
rect 2093 553 2107 567
rect 2053 513 2067 527
rect 2033 413 2047 427
rect 1993 373 2007 387
rect 2193 833 2207 847
rect 2173 813 2187 827
rect 2213 813 2227 827
rect 2513 1733 2527 1747
rect 2593 1793 2607 1807
rect 2633 1793 2647 1807
rect 2673 1953 2687 1967
rect 2753 1993 2767 2007
rect 2733 1833 2747 1847
rect 2573 1753 2587 1767
rect 2553 1673 2567 1687
rect 2553 1653 2567 1667
rect 2533 1593 2547 1607
rect 2733 1813 2747 1827
rect 2693 1773 2707 1787
rect 2853 2273 2867 2287
rect 2913 2553 2927 2567
rect 2973 2733 2987 2747
rect 3013 2713 3027 2727
rect 3053 2973 3067 2987
rect 3033 2673 3047 2687
rect 2993 2633 3007 2647
rect 3033 2573 3047 2587
rect 2933 2533 2947 2547
rect 2913 2513 2927 2527
rect 2953 2493 2967 2507
rect 2913 2413 2927 2427
rect 2973 2413 2987 2427
rect 2893 2173 2907 2187
rect 3233 3213 3247 3227
rect 3293 3233 3307 3247
rect 3273 3193 3287 3207
rect 3253 3113 3267 3127
rect 3213 3053 3227 3067
rect 3193 3033 3207 3047
rect 3153 3013 3167 3027
rect 3173 3013 3187 3027
rect 3133 2993 3147 3007
rect 3093 2933 3107 2947
rect 3093 2873 3107 2887
rect 3093 2793 3107 2807
rect 3113 2693 3127 2707
rect 3073 2553 3087 2567
rect 3253 2973 3267 2987
rect 3253 2713 3267 2727
rect 3213 2693 3227 2707
rect 3353 3233 3367 3247
rect 3533 3733 3547 3747
rect 3573 3733 3587 3747
rect 3553 3693 3567 3707
rect 3713 3713 3727 3727
rect 3733 3693 3747 3707
rect 3693 3673 3707 3687
rect 3633 3633 3647 3647
rect 3493 3593 3507 3607
rect 3593 3593 3607 3607
rect 3473 3553 3487 3567
rect 3473 3533 3487 3547
rect 3533 3553 3547 3567
rect 3573 3553 3587 3567
rect 3513 3533 3527 3547
rect 3613 3513 3627 3527
rect 3553 3493 3567 3507
rect 3493 3473 3507 3487
rect 3553 3473 3567 3487
rect 3473 3333 3487 3347
rect 3473 3313 3487 3327
rect 3433 3253 3447 3267
rect 3313 3213 3327 3227
rect 3373 3213 3387 3227
rect 3333 3153 3347 3167
rect 3393 3193 3407 3207
rect 3393 3093 3407 3107
rect 3373 3073 3387 3087
rect 3353 3033 3367 3047
rect 3453 3213 3467 3227
rect 3533 3333 3547 3347
rect 3533 3253 3547 3267
rect 3473 3193 3487 3207
rect 3493 3073 3507 3087
rect 3433 3033 3447 3047
rect 3493 3013 3507 3027
rect 3293 2993 3307 3007
rect 3393 2993 3407 3007
rect 3213 2673 3227 2687
rect 3153 2653 3167 2667
rect 3093 2533 3107 2547
rect 3133 2533 3147 2547
rect 3093 2353 3107 2367
rect 2993 2293 3007 2307
rect 2933 2253 2947 2267
rect 2933 2233 2947 2247
rect 2913 2153 2927 2167
rect 2913 2073 2927 2087
rect 2973 2253 2987 2267
rect 2953 2193 2967 2207
rect 2973 2173 2987 2187
rect 3013 2173 3027 2187
rect 2913 2033 2927 2047
rect 2813 1933 2827 1947
rect 2853 1793 2867 1807
rect 2893 1793 2907 1807
rect 2933 1853 2947 1867
rect 2953 1793 2967 1807
rect 2773 1773 2787 1787
rect 2873 1773 2887 1787
rect 2913 1773 2927 1787
rect 2793 1753 2807 1767
rect 2813 1753 2827 1767
rect 2833 1753 2847 1767
rect 2773 1673 2787 1687
rect 2613 1633 2627 1647
rect 2673 1633 2687 1647
rect 2713 1633 2727 1647
rect 2753 1633 2767 1647
rect 2593 1613 2607 1627
rect 2533 1573 2547 1587
rect 2573 1573 2587 1587
rect 2633 1593 2647 1607
rect 2693 1593 2707 1607
rect 2733 1613 2747 1627
rect 2833 1673 2847 1687
rect 2933 1633 2947 1647
rect 2833 1613 2847 1627
rect 2933 1613 2947 1627
rect 2753 1593 2767 1607
rect 2853 1593 2867 1607
rect 2893 1593 2907 1607
rect 2913 1593 2927 1607
rect 2953 1593 2967 1607
rect 2793 1573 2807 1587
rect 2833 1573 2847 1587
rect 2873 1573 2887 1587
rect 2553 1553 2567 1567
rect 2613 1553 2627 1567
rect 2653 1553 2667 1567
rect 2773 1553 2787 1567
rect 2493 1493 2507 1507
rect 2433 1333 2447 1347
rect 2473 1333 2487 1347
rect 2513 1313 2527 1327
rect 2793 1533 2807 1547
rect 2653 1353 2667 1367
rect 2593 1333 2607 1347
rect 2713 1333 2727 1347
rect 2813 1333 2827 1347
rect 2773 1313 2787 1327
rect 2813 1313 2827 1327
rect 2593 1293 2607 1307
rect 2453 1273 2467 1287
rect 2493 1273 2507 1287
rect 2633 1293 2647 1307
rect 2673 1293 2687 1307
rect 2753 1293 2767 1307
rect 2833 1293 2847 1307
rect 2793 1233 2807 1247
rect 2693 1193 2707 1207
rect 2633 1173 2647 1187
rect 2453 1093 2467 1107
rect 2613 1133 2627 1147
rect 2593 1113 2607 1127
rect 2673 1153 2687 1167
rect 2853 1173 2867 1187
rect 2693 1133 2707 1147
rect 2733 1113 2747 1127
rect 2793 1113 2807 1127
rect 2893 1553 2907 1567
rect 2913 1533 2927 1547
rect 2873 1153 2887 1167
rect 2893 1153 2907 1167
rect 2533 1093 2547 1107
rect 2613 1093 2627 1107
rect 2653 1093 2667 1107
rect 2513 1073 2527 1087
rect 2553 1073 2567 1087
rect 2653 1073 2667 1087
rect 2513 973 2527 987
rect 2493 953 2507 967
rect 2413 873 2427 887
rect 2353 853 2367 867
rect 2313 833 2327 847
rect 2393 833 2407 847
rect 2433 833 2447 847
rect 2273 813 2287 827
rect 2173 793 2187 807
rect 2233 793 2247 807
rect 2293 793 2307 807
rect 2253 773 2267 787
rect 2193 753 2207 767
rect 2173 613 2187 627
rect 2233 673 2247 687
rect 2273 733 2287 747
rect 2213 633 2227 647
rect 2253 633 2267 647
rect 2433 753 2447 767
rect 2373 693 2387 707
rect 2333 673 2347 687
rect 2373 673 2387 687
rect 2313 653 2327 667
rect 2333 653 2347 667
rect 2413 653 2427 667
rect 2393 633 2407 647
rect 2153 593 2167 607
rect 2193 593 2207 607
rect 2173 573 2187 587
rect 2173 533 2187 547
rect 2133 513 2147 527
rect 2133 473 2147 487
rect 2173 473 2187 487
rect 2113 413 2127 427
rect 2193 453 2207 467
rect 2073 373 2087 387
rect 2093 373 2107 387
rect 1813 333 1827 347
rect 1833 333 1847 347
rect 1913 333 1927 347
rect 1793 273 1807 287
rect 1773 253 1787 267
rect 1773 193 1787 207
rect 1753 153 1767 167
rect 1673 133 1687 147
rect 1693 133 1707 147
rect 1593 113 1607 127
rect 1633 113 1647 127
rect 1393 93 1407 107
rect 1473 73 1487 87
rect 1313 13 1327 27
rect 1733 133 1747 147
rect 1853 313 1867 327
rect 1873 253 1887 267
rect 1913 153 1927 167
rect 1713 113 1727 127
rect 1753 113 1767 127
rect 1813 113 1827 127
rect 1693 93 1707 107
rect 1793 93 1807 107
rect 1833 73 1847 87
rect 1513 53 1527 67
rect 1753 53 1767 67
rect 1893 113 1907 127
rect 1913 113 1927 127
rect 1873 33 1887 47
rect 1913 73 1927 87
rect 1953 293 1967 307
rect 2013 353 2027 367
rect 2053 353 2067 367
rect 2053 333 2067 347
rect 2133 353 2147 367
rect 2013 313 2027 327
rect 1993 293 2007 307
rect 2033 293 2047 307
rect 1973 253 1987 267
rect 1953 173 1967 187
rect 1973 153 1987 167
rect 1933 33 1947 47
rect 2013 213 2027 227
rect 2073 233 2087 247
rect 2093 193 2107 207
rect 2053 173 2067 187
rect 2073 173 2087 187
rect 2013 153 2027 167
rect 1993 93 2007 107
rect 2053 73 2067 87
rect 2133 293 2147 307
rect 2213 373 2227 387
rect 2293 613 2307 627
rect 2353 613 2367 627
rect 2273 593 2287 607
rect 2293 593 2307 607
rect 2493 853 2507 867
rect 2453 693 2467 707
rect 2473 673 2487 687
rect 2553 953 2567 967
rect 3193 2553 3207 2567
rect 3153 2293 3167 2307
rect 3053 2253 3067 2267
rect 3073 2253 3087 2267
rect 3113 2193 3127 2207
rect 2993 2113 3007 2127
rect 3033 2113 3047 2127
rect 3053 2093 3067 2107
rect 3173 2253 3187 2267
rect 3193 2253 3207 2267
rect 3233 2593 3247 2607
rect 3373 2953 3387 2967
rect 3293 2613 3307 2627
rect 3333 2573 3347 2587
rect 3353 2573 3367 2587
rect 3433 2933 3447 2947
rect 3593 3313 3607 3327
rect 3653 3573 3667 3587
rect 3673 3553 3687 3567
rect 3653 3533 3667 3547
rect 3813 4193 3827 4207
rect 3833 4193 3847 4207
rect 3973 4513 3987 4527
rect 3953 4373 3967 4387
rect 3933 4213 3947 4227
rect 3873 4173 3887 4187
rect 3913 4173 3927 4187
rect 3913 4133 3927 4147
rect 3873 4073 3887 4087
rect 3853 4033 3867 4047
rect 3933 4033 3947 4047
rect 3913 4013 3927 4027
rect 3813 3993 3827 4007
rect 3893 3993 3907 4007
rect 4053 4573 4067 4587
rect 4033 4553 4047 4567
rect 4113 4573 4127 4587
rect 4133 4573 4147 4587
rect 4153 4553 4167 4567
rect 4233 4573 4247 4587
rect 4193 4533 4207 4547
rect 4133 4493 4147 4507
rect 4153 4493 4167 4507
rect 4113 4473 4127 4487
rect 4093 4433 4107 4447
rect 4053 4413 4067 4427
rect 4033 4393 4047 4407
rect 4173 4433 4187 4447
rect 4233 4453 4247 4467
rect 4193 4393 4207 4407
rect 4033 4293 4047 4307
rect 4093 4293 4107 4307
rect 4133 4293 4147 4307
rect 4013 4153 4027 4167
rect 4193 4233 4207 4247
rect 4213 4233 4227 4247
rect 4133 4213 4147 4227
rect 4053 4173 4067 4187
rect 4173 4193 4187 4207
rect 4073 4153 4087 4167
rect 4033 4093 4047 4107
rect 4193 4153 4207 4167
rect 4313 4573 4327 4587
rect 4353 4573 4367 4587
rect 4333 4493 4347 4507
rect 4273 4473 4287 4487
rect 4313 4473 4327 4487
rect 4293 4453 4307 4467
rect 4293 4433 4307 4447
rect 4273 4173 4287 4187
rect 4213 4093 4227 4107
rect 4233 4093 4247 4107
rect 4033 4053 4047 4067
rect 4073 4053 4087 4067
rect 4093 4053 4107 4067
rect 4133 4053 4147 4067
rect 4193 4053 4207 4067
rect 3833 3973 3847 3987
rect 3853 3973 3867 3987
rect 3853 3933 3867 3947
rect 3813 3913 3827 3927
rect 3873 3913 3887 3927
rect 3773 3673 3787 3687
rect 3793 3673 3807 3687
rect 3893 3713 3907 3727
rect 3873 3693 3887 3707
rect 3813 3653 3827 3667
rect 3813 3593 3827 3607
rect 3753 3533 3767 3547
rect 3853 3513 3867 3527
rect 3713 3493 3727 3507
rect 3753 3493 3767 3507
rect 3793 3493 3807 3507
rect 3693 3473 3707 3487
rect 3773 3453 3787 3467
rect 3833 3453 3847 3467
rect 3833 3433 3847 3447
rect 3573 3293 3587 3307
rect 3593 3293 3607 3307
rect 3633 3293 3647 3307
rect 3613 3253 3627 3267
rect 3593 3233 3607 3247
rect 3773 3313 3787 3327
rect 3693 3253 3707 3267
rect 3573 3133 3587 3147
rect 3633 3133 3647 3147
rect 3533 3013 3547 3027
rect 3413 2713 3427 2727
rect 3433 2713 3447 2727
rect 3493 2733 3507 2747
rect 3453 2673 3467 2687
rect 3493 2693 3507 2707
rect 3453 2633 3467 2647
rect 3473 2633 3487 2647
rect 3473 2593 3487 2607
rect 3473 2553 3487 2567
rect 3293 2533 3307 2547
rect 3313 2513 3327 2527
rect 3273 2493 3287 2507
rect 3253 2453 3267 2467
rect 3293 2313 3307 2327
rect 3233 2253 3247 2267
rect 3253 2253 3267 2267
rect 3213 2213 3227 2227
rect 3133 2173 3147 2187
rect 3173 2173 3187 2187
rect 3193 2113 3207 2127
rect 3213 2093 3227 2107
rect 3093 2073 3107 2087
rect 3173 2073 3187 2087
rect 3133 2053 3147 2067
rect 3153 2053 3167 2067
rect 3113 2033 3127 2047
rect 3133 1993 3147 2007
rect 3153 1853 3167 1867
rect 3053 1813 3067 1827
rect 3133 1813 3147 1827
rect 2993 1613 3007 1627
rect 3053 1773 3067 1787
rect 3073 1773 3087 1787
rect 3093 1773 3107 1787
rect 3033 1753 3047 1767
rect 3133 1693 3147 1707
rect 3133 1633 3147 1647
rect 3213 1633 3227 1647
rect 2993 1573 3007 1587
rect 3093 1593 3107 1607
rect 3333 2233 3347 2247
rect 3393 2533 3407 2547
rect 3393 2513 3407 2527
rect 3433 2513 3447 2527
rect 3373 2253 3387 2267
rect 3353 2213 3367 2227
rect 3293 2193 3307 2207
rect 3253 2153 3267 2167
rect 3273 2133 3287 2147
rect 3313 2073 3327 2087
rect 3253 2053 3267 2067
rect 3293 2053 3307 2067
rect 3333 2053 3347 2067
rect 3273 1933 3287 1947
rect 3253 1693 3267 1707
rect 3173 1593 3187 1607
rect 3233 1593 3247 1607
rect 3053 1573 3067 1587
rect 3113 1573 3127 1587
rect 3153 1573 3167 1587
rect 3213 1573 3227 1587
rect 3233 1553 3247 1567
rect 3173 1533 3187 1547
rect 3193 1533 3207 1547
rect 2973 1353 2987 1367
rect 2993 1313 3007 1327
rect 2973 1273 2987 1287
rect 2933 1253 2947 1267
rect 2973 1153 2987 1167
rect 2993 1133 3007 1147
rect 2973 1113 2987 1127
rect 3253 1373 3267 1387
rect 3173 1353 3187 1367
rect 3253 1353 3267 1367
rect 3093 1333 3107 1347
rect 3053 1293 3067 1307
rect 3073 1293 3087 1307
rect 3013 1113 3027 1127
rect 3033 1093 3047 1107
rect 3113 1293 3127 1307
rect 3213 1333 3227 1347
rect 3193 1253 3207 1267
rect 3233 1253 3247 1267
rect 3373 2033 3387 2047
rect 3453 2073 3467 2087
rect 3433 2013 3447 2027
rect 3293 1833 3307 1847
rect 3333 1833 3347 1847
rect 3453 1833 3467 1847
rect 3413 1813 3427 1827
rect 3333 1793 3347 1807
rect 3373 1793 3387 1807
rect 3433 1793 3447 1807
rect 3373 1773 3387 1787
rect 3353 1733 3367 1747
rect 3333 1653 3347 1667
rect 3313 1633 3327 1647
rect 3353 1613 3367 1627
rect 3333 1593 3347 1607
rect 3333 1553 3347 1567
rect 3333 1533 3347 1547
rect 3293 1513 3307 1527
rect 3293 1373 3307 1387
rect 3273 1193 3287 1207
rect 3133 1153 3147 1167
rect 3173 1133 3187 1147
rect 3213 1133 3227 1147
rect 3253 1113 3267 1127
rect 3113 1093 3127 1107
rect 2913 1053 2927 1067
rect 2993 1053 3007 1067
rect 2553 853 2567 867
rect 2753 853 2767 867
rect 2793 853 2807 867
rect 2893 853 2907 867
rect 2933 853 2947 867
rect 2573 833 2587 847
rect 2593 833 2607 847
rect 2573 793 2587 807
rect 2633 833 2647 847
rect 2673 833 2687 847
rect 2773 833 2787 847
rect 2853 833 2867 847
rect 2613 813 2627 827
rect 2693 813 2707 827
rect 2833 813 2847 827
rect 2653 793 2667 807
rect 2573 733 2587 747
rect 2533 713 2547 727
rect 2453 653 2467 667
rect 2513 653 2527 667
rect 2473 633 2487 647
rect 2453 613 2467 627
rect 2473 613 2487 627
rect 2513 613 2527 627
rect 2453 593 2467 607
rect 2493 593 2507 607
rect 2413 493 2427 507
rect 2293 473 2307 487
rect 2273 433 2287 447
rect 2413 413 2427 427
rect 2333 393 2347 407
rect 2193 353 2207 367
rect 2233 353 2247 367
rect 2333 373 2347 387
rect 2213 313 2227 327
rect 2193 273 2207 287
rect 2133 213 2147 227
rect 2173 213 2187 227
rect 2193 213 2207 227
rect 2153 193 2167 207
rect 2173 193 2187 207
rect 2113 53 2127 67
rect 2213 153 2227 167
rect 2273 333 2287 347
rect 2313 333 2327 347
rect 2353 333 2367 347
rect 2373 313 2387 327
rect 2253 293 2267 307
rect 2393 293 2407 307
rect 2253 273 2267 287
rect 2393 253 2407 267
rect 2253 193 2267 207
rect 2353 193 2367 207
rect 2353 173 2367 187
rect 2173 133 2187 147
rect 2193 133 2207 147
rect 2313 153 2327 167
rect 2433 353 2447 367
rect 2433 333 2447 347
rect 2413 193 2427 207
rect 2493 373 2507 387
rect 2473 333 2487 347
rect 2453 213 2467 227
rect 2553 593 2567 607
rect 2673 653 2687 667
rect 2693 633 2707 647
rect 2773 633 2787 647
rect 2913 813 2927 827
rect 2913 713 2927 727
rect 2953 833 2967 847
rect 2973 793 2987 807
rect 3073 833 3087 847
rect 3053 813 3067 827
rect 3013 793 3027 807
rect 2993 753 3007 767
rect 2953 713 2967 727
rect 2933 633 2947 647
rect 2673 613 2687 627
rect 2733 613 2747 627
rect 2653 593 2667 607
rect 2713 593 2727 607
rect 2673 533 2687 547
rect 2733 533 2747 547
rect 2553 413 2567 427
rect 2633 413 2647 427
rect 2533 373 2547 387
rect 2573 393 2587 407
rect 2693 393 2707 407
rect 2573 353 2587 367
rect 2633 353 2647 367
rect 2533 293 2547 307
rect 2553 193 2567 207
rect 2593 173 2607 187
rect 2593 153 2607 167
rect 2673 353 2687 367
rect 2753 393 2767 407
rect 2733 373 2747 387
rect 2873 413 2887 427
rect 2853 373 2867 387
rect 2773 353 2787 367
rect 2753 333 2767 347
rect 2793 333 2807 347
rect 2833 333 2847 347
rect 2893 373 2907 387
rect 2933 373 2947 387
rect 2913 353 2927 367
rect 2873 333 2887 347
rect 2653 313 2667 327
rect 2713 313 2727 327
rect 2813 313 2827 327
rect 2853 313 2867 327
rect 2653 253 2667 267
rect 2693 253 2707 267
rect 2253 113 2267 127
rect 2233 93 2247 107
rect 2333 133 2347 147
rect 2413 133 2427 147
rect 2573 133 2587 147
rect 3093 793 3107 807
rect 3153 793 3167 807
rect 3233 833 3247 847
rect 3073 773 3087 787
rect 3113 773 3127 787
rect 3133 773 3147 787
rect 3193 773 3207 787
rect 3073 753 3087 767
rect 3033 653 3047 667
rect 3253 813 3267 827
rect 3193 653 3207 667
rect 3213 653 3227 667
rect 3233 653 3247 667
rect 3273 653 3287 667
rect 3173 633 3187 647
rect 3093 613 3107 627
rect 3153 613 3167 627
rect 3053 593 3067 607
rect 3013 373 3027 387
rect 2973 293 2987 307
rect 2713 133 2727 147
rect 2533 113 2547 127
rect 2613 113 2627 127
rect 2473 93 2487 107
rect 2953 233 2967 247
rect 2773 193 2787 207
rect 2853 173 2867 187
rect 2773 153 2787 167
rect 3013 233 3027 247
rect 3453 1753 3467 1767
rect 3393 1613 3407 1627
rect 3433 1593 3447 1607
rect 3373 1573 3387 1587
rect 3413 1553 3427 1567
rect 3353 1513 3367 1527
rect 3353 1233 3367 1247
rect 3533 2773 3547 2787
rect 3553 2773 3567 2787
rect 3533 2653 3547 2667
rect 3533 2613 3547 2627
rect 3513 2513 3527 2527
rect 3633 3093 3647 3107
rect 3753 3213 3767 3227
rect 3913 3573 3927 3587
rect 4013 4013 4027 4027
rect 3993 3993 4007 4007
rect 4053 3993 4067 4007
rect 3973 3953 3987 3967
rect 4093 4033 4107 4047
rect 4113 3993 4127 4007
rect 4153 4013 4167 4027
rect 4193 3993 4207 4007
rect 4173 3973 4187 3987
rect 4213 3973 4227 3987
rect 4053 3833 4067 3847
rect 4233 3853 4247 3867
rect 4393 4393 4407 4407
rect 4353 4213 4367 4227
rect 4313 4193 4327 4207
rect 4433 4193 4447 4207
rect 4473 4193 4487 4207
rect 4373 4173 4387 4187
rect 4333 4153 4347 4167
rect 4453 4153 4467 4167
rect 4513 4473 4527 4487
rect 4553 4233 4567 4247
rect 4513 4173 4527 4187
rect 4493 4133 4507 4147
rect 4513 4133 4527 4147
rect 4373 4113 4387 4127
rect 4413 4113 4427 4127
rect 4293 4093 4307 4107
rect 4273 4073 4287 4087
rect 4333 4073 4347 4087
rect 4273 3993 4287 4007
rect 4293 3993 4307 4007
rect 4313 3973 4327 3987
rect 4293 3853 4307 3867
rect 4253 3733 4267 3747
rect 4193 3713 4207 3727
rect 4233 3713 4247 3727
rect 4273 3713 4287 3727
rect 3913 3533 3927 3547
rect 3953 3533 3967 3547
rect 3953 3513 3967 3527
rect 3893 3453 3907 3467
rect 3933 3453 3947 3467
rect 3873 3393 3887 3407
rect 4073 3673 4087 3687
rect 4053 3573 4067 3587
rect 4033 3553 4047 3567
rect 4033 3533 4047 3547
rect 4013 3453 4027 3467
rect 3893 3273 3907 3287
rect 3913 3273 3927 3287
rect 3953 3273 3967 3287
rect 3973 3273 3987 3287
rect 4013 3273 4027 3287
rect 3873 3253 3887 3267
rect 3813 3153 3827 3167
rect 3833 3153 3847 3167
rect 3713 3093 3727 3107
rect 3713 3073 3727 3087
rect 3773 3073 3787 3087
rect 3673 3053 3687 3067
rect 3633 3033 3647 3047
rect 3673 3033 3687 3047
rect 3713 3033 3727 3047
rect 3753 3033 3767 3047
rect 3793 3033 3807 3047
rect 3613 3013 3627 3027
rect 3653 2993 3667 3007
rect 3633 2873 3647 2887
rect 3593 2773 3607 2787
rect 3593 2733 3607 2747
rect 3613 2633 3627 2647
rect 3593 2553 3607 2567
rect 3553 2493 3567 2507
rect 3573 2493 3587 2507
rect 3533 2353 3547 2367
rect 3493 2273 3507 2287
rect 3573 2353 3587 2367
rect 3553 2293 3567 2307
rect 3513 2253 3527 2267
rect 3773 3013 3787 3027
rect 3813 3013 3827 3027
rect 3713 2993 3727 3007
rect 3713 2973 3727 2987
rect 3673 2853 3687 2867
rect 3653 2773 3667 2787
rect 3653 2733 3667 2747
rect 3673 2593 3687 2607
rect 3693 2553 3707 2567
rect 3673 2353 3687 2367
rect 3693 2353 3707 2367
rect 3633 2313 3647 2327
rect 3653 2313 3667 2327
rect 3613 2273 3627 2287
rect 3653 2273 3667 2287
rect 3493 2233 3507 2247
rect 3513 2213 3527 2227
rect 3493 2013 3507 2027
rect 3593 2253 3607 2267
rect 3633 2253 3647 2267
rect 3673 2253 3687 2267
rect 3593 2233 3607 2247
rect 3593 2193 3607 2207
rect 3573 2173 3587 2187
rect 3533 2113 3547 2127
rect 3533 2073 3547 2087
rect 3573 2073 3587 2087
rect 3553 1853 3567 1867
rect 3513 1813 3527 1827
rect 3493 1753 3507 1767
rect 3473 1713 3487 1727
rect 3513 1633 3527 1647
rect 3473 1593 3487 1607
rect 3473 1533 3487 1547
rect 3413 1493 3427 1507
rect 3453 1493 3467 1507
rect 3393 1273 3407 1287
rect 3393 1233 3407 1247
rect 3333 1133 3347 1147
rect 3373 1193 3387 1207
rect 3373 1173 3387 1187
rect 3473 1293 3487 1307
rect 3453 1213 3467 1227
rect 3473 1153 3487 1167
rect 3413 1093 3427 1107
rect 3313 853 3327 867
rect 3353 853 3367 867
rect 3393 853 3407 867
rect 3333 833 3347 847
rect 3373 833 3387 847
rect 3413 813 3427 827
rect 3333 753 3347 767
rect 3393 753 3407 767
rect 3253 633 3267 647
rect 3293 633 3307 647
rect 3273 613 3287 627
rect 3293 613 3307 627
rect 3233 593 3247 607
rect 3353 673 3367 687
rect 3173 573 3187 587
rect 3213 573 3227 587
rect 3493 1093 3507 1107
rect 3473 813 3487 827
rect 3493 793 3507 807
rect 3493 713 3507 727
rect 3533 1613 3547 1627
rect 3653 2233 3667 2247
rect 3673 2133 3687 2147
rect 3613 2093 3627 2107
rect 3613 2073 3627 2087
rect 3653 2073 3667 2087
rect 3633 1993 3647 2007
rect 3613 1933 3627 1947
rect 3573 1753 3587 1767
rect 3653 1853 3667 1867
rect 3573 1713 3587 1727
rect 3573 1613 3587 1627
rect 3573 1553 3587 1567
rect 3533 1313 3547 1327
rect 3553 1273 3567 1287
rect 3633 1733 3647 1747
rect 3613 1673 3627 1687
rect 3653 1633 3667 1647
rect 3813 2953 3827 2967
rect 3733 2913 3747 2927
rect 3773 2913 3787 2927
rect 3853 3113 3867 3127
rect 3853 3033 3867 3047
rect 3913 3133 3927 3147
rect 3893 3053 3907 3067
rect 3853 3013 3867 3027
rect 3893 3013 3907 3027
rect 3953 3213 3967 3227
rect 4053 3513 4067 3527
rect 4113 3653 4127 3667
rect 4093 3593 4107 3607
rect 4073 3433 4087 3447
rect 4073 3313 4087 3327
rect 4033 3253 4047 3267
rect 4013 3233 4027 3247
rect 3993 3213 4007 3227
rect 3973 3173 3987 3187
rect 4013 3193 4027 3207
rect 4013 3153 4027 3167
rect 3993 3133 4007 3147
rect 3993 3113 4007 3127
rect 4013 3113 4027 3127
rect 3973 3073 3987 3087
rect 4053 3153 4067 3167
rect 4093 3213 4107 3227
rect 4253 3693 4267 3707
rect 4193 3673 4207 3687
rect 4173 3633 4187 3647
rect 4153 3613 4167 3627
rect 4173 3593 4187 3607
rect 4153 3553 4167 3567
rect 4153 3413 4167 3427
rect 4113 3193 4127 3207
rect 4073 3113 4087 3127
rect 4113 3093 4127 3107
rect 4013 3073 4027 3087
rect 4033 3073 4047 3087
rect 3953 3033 3967 3047
rect 4093 3053 4107 3067
rect 4073 3033 4087 3047
rect 3993 3013 4007 3027
rect 4053 3013 4067 3027
rect 4173 3233 4187 3247
rect 4213 3653 4227 3667
rect 4313 3833 4327 3847
rect 4293 3633 4307 3647
rect 4273 3613 4287 3627
rect 4313 3613 4327 3627
rect 4293 3513 4307 3527
rect 4213 3413 4227 3427
rect 4413 3973 4427 3987
rect 4353 3593 4367 3607
rect 4373 3593 4387 3607
rect 4553 3993 4567 4007
rect 4613 4513 4627 4527
rect 4673 4453 4687 4467
rect 4713 4453 4727 4467
rect 4613 4433 4627 4447
rect 4593 4133 4607 4147
rect 4493 3753 4507 3767
rect 4533 3753 4547 3767
rect 4433 3693 4447 3707
rect 4413 3613 4427 3627
rect 4413 3593 4427 3607
rect 4393 3513 4407 3527
rect 4393 3493 4407 3507
rect 4333 3453 4347 3467
rect 4353 3453 4367 3467
rect 4473 3513 4487 3527
rect 4453 3493 4467 3507
rect 4453 3293 4467 3307
rect 4413 3273 4427 3287
rect 4433 3273 4447 3287
rect 4493 3313 4507 3327
rect 4313 3253 4327 3267
rect 4333 3253 4347 3267
rect 4193 3213 4207 3227
rect 4253 3233 4267 3247
rect 4233 3213 4247 3227
rect 4273 3213 4287 3227
rect 4173 3173 4187 3187
rect 4213 3153 4227 3167
rect 4133 3073 4147 3087
rect 4193 3053 4207 3067
rect 4173 3033 4187 3047
rect 4113 3013 4127 3027
rect 3973 2993 3987 3007
rect 4113 2993 4127 3007
rect 4133 2993 4147 3007
rect 3833 2873 3847 2887
rect 3813 2833 3827 2847
rect 3773 2813 3787 2827
rect 3793 2773 3807 2787
rect 3733 2693 3747 2707
rect 3793 2653 3807 2667
rect 3773 2613 3787 2627
rect 3713 2313 3727 2327
rect 3713 2273 3727 2287
rect 3713 2233 3727 2247
rect 3713 1933 3727 1947
rect 3933 2813 3947 2827
rect 3853 2793 3867 2807
rect 3893 2773 3907 2787
rect 3873 2733 3887 2747
rect 3833 2713 3847 2727
rect 3813 2593 3827 2607
rect 3773 2533 3787 2547
rect 3813 2493 3827 2507
rect 3773 2393 3787 2407
rect 3813 2373 3827 2387
rect 3773 2293 3787 2307
rect 3813 2293 3827 2307
rect 3773 2253 3787 2267
rect 3753 2193 3767 2207
rect 3813 2253 3827 2267
rect 4093 2973 4107 2987
rect 4033 2813 4047 2827
rect 3973 2753 3987 2767
rect 3853 2693 3867 2707
rect 3893 2693 3907 2707
rect 3933 2693 3947 2707
rect 3913 2593 3927 2607
rect 3973 2713 3987 2727
rect 4053 2733 4067 2747
rect 4013 2713 4027 2727
rect 4053 2713 4067 2727
rect 3993 2693 4007 2707
rect 3993 2633 4007 2647
rect 4073 2693 4087 2707
rect 3973 2613 3987 2627
rect 4053 2613 4067 2627
rect 3953 2573 3967 2587
rect 4173 2993 4187 3007
rect 4153 2953 4167 2967
rect 4133 2813 4147 2827
rect 4133 2753 4147 2767
rect 4253 3193 4267 3207
rect 4273 3193 4287 3207
rect 4253 3153 4267 3167
rect 4253 3133 4267 3147
rect 4233 3113 4247 3127
rect 4233 3053 4247 3067
rect 4373 3233 4387 3247
rect 4413 3233 4427 3247
rect 4333 3193 4347 3207
rect 4293 3133 4307 3147
rect 4293 3113 4307 3127
rect 4233 3013 4247 3027
rect 4313 3073 4327 3087
rect 4353 3173 4367 3187
rect 4413 3213 4427 3227
rect 4393 3153 4407 3167
rect 4373 3133 4387 3147
rect 4353 3113 4367 3127
rect 4293 3033 4307 3047
rect 4293 3013 4307 3027
rect 4233 2933 4247 2947
rect 4333 3053 4347 3067
rect 4353 3033 4367 3047
rect 4353 2993 4367 3007
rect 4273 2973 4287 2987
rect 4293 2973 4307 2987
rect 4273 2913 4287 2927
rect 4273 2853 4287 2867
rect 4253 2833 4267 2847
rect 4213 2773 4227 2787
rect 4113 2713 4127 2727
rect 4113 2693 4127 2707
rect 4013 2593 4027 2607
rect 4093 2593 4107 2607
rect 3873 2553 3887 2567
rect 3953 2553 3967 2567
rect 3993 2553 4007 2567
rect 3893 2533 3907 2547
rect 3933 2533 3947 2547
rect 3973 2533 3987 2547
rect 3853 2473 3867 2487
rect 3933 2473 3947 2487
rect 3953 2473 3967 2487
rect 3873 2353 3887 2367
rect 4073 2573 4087 2587
rect 4033 2553 4047 2567
rect 4053 2513 4067 2527
rect 4033 2493 4047 2507
rect 4093 2493 4107 2507
rect 4073 2453 4087 2467
rect 4053 2433 4067 2447
rect 4013 2393 4027 2407
rect 3993 2373 4007 2387
rect 3973 2313 3987 2327
rect 3933 2293 3947 2307
rect 3913 2273 3927 2287
rect 3953 2273 3967 2287
rect 4053 2293 4067 2307
rect 4033 2273 4047 2287
rect 3853 2233 3867 2247
rect 3933 2253 3947 2267
rect 3833 2193 3847 2207
rect 3793 2133 3807 2147
rect 3813 2133 3827 2147
rect 3933 2133 3947 2147
rect 3813 2093 3827 2107
rect 3833 2093 3847 2107
rect 3793 2073 3807 2087
rect 3873 2073 3887 2087
rect 3793 2013 3807 2027
rect 3813 2013 3827 2027
rect 3773 1773 3787 1787
rect 3733 1753 3747 1767
rect 3753 1753 3767 1767
rect 3813 1833 3827 1847
rect 3913 2053 3927 2067
rect 3893 1933 3907 1947
rect 3853 1793 3867 1807
rect 3813 1773 3827 1787
rect 3873 1773 3887 1787
rect 3813 1753 3827 1767
rect 3793 1713 3807 1727
rect 3793 1673 3807 1687
rect 3773 1633 3787 1647
rect 3713 1533 3727 1547
rect 3613 1493 3627 1507
rect 3593 1453 3607 1467
rect 3653 1453 3667 1467
rect 3613 1313 3627 1327
rect 3593 1293 3607 1307
rect 3633 1293 3647 1307
rect 3593 1273 3607 1287
rect 3613 1273 3627 1287
rect 3633 1273 3647 1287
rect 3613 1233 3627 1247
rect 3573 1113 3587 1127
rect 3593 1113 3607 1127
rect 3753 1613 3767 1627
rect 3793 1573 3807 1587
rect 3773 1553 3787 1567
rect 3733 1333 3747 1347
rect 3753 1313 3767 1327
rect 3713 1293 3727 1307
rect 3673 1273 3687 1287
rect 3693 1273 3707 1287
rect 3693 1093 3707 1107
rect 3653 973 3667 987
rect 3633 853 3647 867
rect 3713 853 3727 867
rect 3533 813 3547 827
rect 3593 813 3607 827
rect 3633 813 3647 827
rect 3713 793 3727 807
rect 3513 673 3527 687
rect 3673 673 3687 687
rect 3393 653 3407 667
rect 3453 653 3467 667
rect 3493 653 3507 667
rect 3573 653 3587 667
rect 3413 633 3427 647
rect 3373 613 3387 627
rect 3453 613 3467 627
rect 3533 633 3547 647
rect 3673 633 3687 647
rect 3873 1733 3887 1747
rect 3853 1693 3867 1707
rect 3833 1653 3847 1667
rect 3833 1593 3847 1607
rect 4013 2253 4027 2267
rect 3973 2233 3987 2247
rect 3993 2233 4007 2247
rect 4013 2213 4027 2227
rect 4033 2213 4047 2227
rect 3973 2073 3987 2087
rect 3993 1953 4007 1967
rect 3953 1813 3967 1827
rect 3913 1793 3927 1807
rect 3953 1793 3967 1807
rect 3973 1773 3987 1787
rect 4053 2093 4067 2107
rect 4033 2073 4047 2087
rect 4053 2013 4067 2027
rect 4013 1933 4027 1947
rect 3953 1713 3967 1727
rect 3893 1673 3907 1687
rect 3893 1653 3907 1667
rect 3933 1613 3947 1627
rect 3833 1573 3847 1587
rect 3873 1573 3887 1587
rect 3813 1553 3827 1567
rect 3993 1733 4007 1747
rect 4173 2713 4187 2727
rect 4193 2713 4207 2727
rect 4153 2673 4167 2687
rect 4133 2653 4147 2667
rect 4113 2433 4127 2447
rect 4153 2613 4167 2627
rect 4133 2333 4147 2347
rect 4153 2233 4167 2247
rect 4093 2073 4107 2087
rect 4073 1953 4087 1967
rect 4113 1853 4127 1867
rect 4033 1773 4047 1787
rect 4033 1753 4047 1767
rect 4053 1753 4067 1767
rect 4013 1713 4027 1727
rect 3993 1593 4007 1607
rect 4113 1773 4127 1787
rect 4073 1733 4087 1747
rect 4073 1693 4087 1707
rect 4093 1693 4107 1707
rect 4053 1653 4067 1667
rect 4093 1653 4107 1667
rect 4113 1653 4127 1667
rect 4013 1573 4027 1587
rect 3853 1333 3867 1347
rect 3873 1333 3887 1347
rect 3953 1333 3967 1347
rect 3813 1293 3827 1307
rect 3793 1273 3807 1287
rect 3873 1253 3887 1267
rect 3933 1293 3947 1307
rect 4073 1613 4087 1627
rect 4093 1613 4107 1627
rect 4153 1933 4167 1947
rect 4153 1653 4167 1667
rect 4233 2713 4247 2727
rect 4233 2693 4247 2707
rect 4213 2633 4227 2647
rect 4193 2533 4207 2547
rect 4213 2533 4227 2547
rect 4273 2713 4287 2727
rect 4253 2513 4267 2527
rect 4233 2473 4247 2487
rect 4213 2253 4227 2267
rect 4313 2933 4327 2947
rect 4393 3113 4407 3127
rect 4433 3173 4447 3187
rect 4413 3073 4427 3087
rect 4393 3053 4407 3067
rect 4313 2693 4327 2707
rect 4373 2733 4387 2747
rect 4413 3033 4427 3047
rect 4413 3013 4427 3027
rect 4413 2953 4427 2967
rect 4433 2873 4447 2887
rect 4413 2713 4427 2727
rect 4433 2713 4447 2727
rect 4393 2633 4407 2647
rect 4313 2553 4327 2567
rect 4333 2533 4347 2547
rect 4313 2513 4327 2527
rect 4233 2233 4247 2247
rect 4333 2293 4347 2307
rect 4193 2093 4207 2107
rect 4293 2133 4307 2147
rect 4313 2113 4327 2127
rect 4433 2533 4447 2547
rect 4433 2513 4447 2527
rect 4413 2253 4427 2267
rect 4373 2133 4387 2147
rect 4413 2133 4427 2147
rect 4333 2093 4347 2107
rect 4353 2093 4367 2107
rect 4413 2093 4427 2107
rect 4193 1933 4207 1947
rect 4193 1913 4207 1927
rect 4233 1913 4247 1927
rect 4093 1573 4107 1587
rect 4053 1533 4067 1547
rect 4053 1313 4067 1327
rect 4093 1313 4107 1327
rect 4073 1293 4087 1307
rect 4033 1233 4047 1247
rect 3933 1193 3947 1207
rect 4013 1193 4027 1207
rect 3813 1133 3827 1147
rect 3853 1133 3867 1147
rect 3893 1133 3907 1147
rect 3793 813 3807 827
rect 3773 713 3787 727
rect 3873 1113 3887 1127
rect 3913 1113 3927 1127
rect 3833 1093 3847 1107
rect 3853 1093 3867 1107
rect 3893 1093 3907 1107
rect 3913 973 3927 987
rect 4013 1113 4027 1127
rect 3973 1093 3987 1107
rect 4033 1093 4047 1107
rect 3953 973 3967 987
rect 3933 853 3947 867
rect 3853 793 3867 807
rect 3933 773 3947 787
rect 3833 673 3847 687
rect 3933 673 3947 687
rect 3813 653 3827 667
rect 3513 613 3527 627
rect 3553 613 3567 627
rect 3873 633 3887 647
rect 3913 633 3927 647
rect 3813 613 3827 627
rect 3793 533 3807 547
rect 3473 413 3487 427
rect 3613 393 3627 407
rect 3633 393 3647 407
rect 3793 393 3807 407
rect 3113 373 3127 387
rect 3353 373 3367 387
rect 3393 373 3407 387
rect 3473 373 3487 387
rect 3073 353 3087 367
rect 3313 353 3327 367
rect 3353 353 3367 367
rect 3053 313 3067 327
rect 3133 333 3147 347
rect 3173 333 3187 347
rect 3233 333 3247 347
rect 3433 353 3447 367
rect 3093 293 3107 307
rect 3073 213 3087 227
rect 3033 193 3047 207
rect 3033 173 3047 187
rect 3073 153 3087 167
rect 3113 153 3127 167
rect 2753 133 2767 147
rect 3193 273 3207 287
rect 3273 253 3287 267
rect 3413 313 3427 327
rect 3453 313 3467 327
rect 3513 333 3527 347
rect 3353 293 3367 307
rect 3493 293 3507 307
rect 3333 233 3347 247
rect 3153 213 3167 227
rect 3193 193 3207 207
rect 2793 133 2807 147
rect 2873 133 2887 147
rect 3133 133 3147 147
rect 3273 153 3287 167
rect 3533 313 3547 327
rect 3513 273 3527 287
rect 3393 173 3407 187
rect 3613 333 3627 347
rect 3693 353 3707 367
rect 3593 313 3607 327
rect 3653 313 3667 327
rect 3753 373 3767 387
rect 3773 353 3787 367
rect 3573 293 3587 307
rect 3733 293 3747 307
rect 3573 253 3587 267
rect 3733 233 3747 247
rect 3693 173 3707 187
rect 3473 153 3487 167
rect 3533 153 3547 167
rect 3573 153 3587 167
rect 3613 153 3627 167
rect 3793 173 3807 187
rect 3893 613 3907 627
rect 4053 1073 4067 1087
rect 4013 853 4027 867
rect 4033 853 4047 867
rect 3973 833 3987 847
rect 3993 813 4007 827
rect 4073 813 4087 827
rect 4173 1613 4187 1627
rect 4313 2053 4327 2067
rect 4333 2053 4347 2067
rect 4333 2033 4347 2047
rect 4273 1833 4287 1847
rect 4213 1793 4227 1807
rect 4253 1793 4267 1807
rect 4293 1793 4307 1807
rect 4513 3273 4527 3287
rect 4473 3253 4487 3267
rect 4493 3233 4507 3247
rect 4473 3073 4487 3087
rect 4493 3073 4507 3087
rect 4553 3493 4567 3507
rect 4473 2853 4487 2867
rect 4493 2773 4507 2787
rect 4533 3033 4547 3047
rect 4593 3473 4607 3487
rect 4673 4293 4687 4307
rect 4633 4113 4647 4127
rect 4673 3973 4687 3987
rect 4633 3953 4647 3967
rect 4633 3913 4647 3927
rect 4733 4433 4747 4447
rect 4733 4293 4747 4307
rect 4713 4193 4727 4207
rect 4713 3973 4727 3987
rect 4693 3753 4707 3767
rect 4633 3713 4647 3727
rect 4673 3673 4687 3687
rect 4653 3653 4667 3667
rect 4633 3513 4647 3527
rect 4673 3513 4687 3527
rect 4653 3493 4667 3507
rect 4693 3493 4707 3507
rect 4673 3473 4687 3487
rect 4653 3453 4667 3467
rect 4633 3293 4647 3307
rect 4673 3273 4687 3287
rect 4653 3253 4667 3267
rect 4673 3233 4687 3247
rect 4653 3193 4667 3207
rect 4653 3093 4667 3107
rect 4633 3073 4647 3087
rect 4653 3073 4667 3087
rect 4773 3713 4787 3727
rect 4753 3493 4767 3507
rect 4733 3233 4747 3247
rect 4693 3213 4707 3227
rect 4733 3213 4747 3227
rect 4613 3033 4627 3047
rect 4673 3053 4687 3067
rect 4673 3033 4687 3047
rect 4733 3173 4747 3187
rect 4733 3053 4747 3067
rect 4613 3013 4627 3027
rect 4593 2993 4607 3007
rect 4553 2973 4567 2987
rect 4693 3013 4707 3027
rect 4653 2993 4667 3007
rect 4673 2993 4687 3007
rect 4613 2913 4627 2927
rect 4693 2973 4707 2987
rect 4553 2793 4567 2807
rect 4613 2793 4627 2807
rect 4673 2793 4687 2807
rect 4573 2733 4587 2747
rect 4533 2713 4547 2727
rect 4593 2713 4607 2727
rect 4553 2693 4567 2707
rect 4513 2673 4527 2687
rect 4473 2573 4487 2587
rect 4513 2553 4527 2567
rect 4533 2553 4547 2567
rect 4453 2493 4467 2507
rect 4633 2773 4647 2787
rect 4633 2733 4647 2747
rect 4593 2553 4607 2567
rect 4613 2553 4627 2567
rect 4673 2733 4687 2747
rect 4653 2713 4667 2727
rect 4693 2693 4707 2707
rect 4553 2513 4567 2527
rect 4573 2513 4587 2527
rect 4613 2513 4627 2527
rect 4633 2513 4647 2527
rect 4493 2473 4507 2487
rect 4693 2513 4707 2527
rect 4653 2493 4667 2507
rect 4613 2473 4627 2487
rect 4573 2333 4587 2347
rect 4693 2473 4707 2487
rect 4573 2313 4587 2327
rect 4533 2293 4547 2307
rect 4453 2253 4467 2267
rect 4613 2273 4627 2287
rect 4593 2253 4607 2267
rect 4553 2173 4567 2187
rect 4693 2313 4707 2327
rect 4653 2293 4667 2307
rect 4673 2273 4687 2287
rect 4673 2253 4687 2267
rect 4533 2153 4547 2167
rect 4593 2153 4607 2167
rect 4533 2133 4547 2147
rect 4473 2113 4487 2127
rect 4493 2093 4507 2107
rect 4373 2053 4387 2067
rect 4513 2073 4527 2087
rect 4493 2053 4507 2067
rect 4353 1793 4367 1807
rect 4233 1753 4247 1767
rect 4233 1733 4247 1747
rect 4213 1693 4227 1707
rect 4273 1693 4287 1707
rect 4293 1673 4307 1687
rect 4273 1653 4287 1667
rect 4253 1613 4267 1627
rect 4133 1533 4147 1547
rect 4213 1573 4227 1587
rect 4253 1573 4267 1587
rect 4193 1533 4207 1547
rect 4173 1393 4187 1407
rect 4173 1373 4187 1387
rect 4133 1353 4147 1367
rect 4153 1313 4167 1327
rect 4133 1133 4147 1147
rect 4173 1133 4187 1147
rect 4253 1533 4267 1547
rect 4213 1493 4227 1507
rect 4333 1773 4347 1787
rect 4413 1773 4427 1787
rect 4333 1693 4347 1707
rect 4313 1653 4327 1667
rect 4393 1753 4407 1767
rect 4393 1733 4407 1747
rect 4333 1613 4347 1627
rect 4353 1613 4367 1627
rect 4373 1593 4387 1607
rect 4353 1573 4367 1587
rect 4313 1553 4327 1567
rect 4353 1553 4367 1567
rect 4253 1413 4267 1427
rect 4293 1413 4307 1427
rect 4213 1353 4227 1367
rect 4193 1073 4207 1087
rect 4293 1393 4307 1407
rect 4373 1513 4387 1527
rect 4273 1173 4287 1187
rect 4333 1313 4347 1327
rect 4413 1673 4427 1687
rect 4453 1793 4467 1807
rect 4513 1833 4527 1847
rect 4493 1773 4507 1787
rect 4453 1713 4467 1727
rect 4413 1653 4427 1667
rect 4433 1653 4447 1667
rect 4433 1573 4447 1587
rect 4473 1693 4487 1707
rect 4553 2073 4567 2087
rect 4553 1833 4567 1847
rect 4573 1773 4587 1787
rect 4633 2133 4647 2147
rect 4733 3013 4747 3027
rect 4773 3073 4787 3087
rect 4773 3053 4787 3067
rect 4773 2913 4787 2927
rect 4753 2733 4767 2747
rect 4773 2333 4787 2347
rect 4733 2253 4747 2267
rect 4653 1813 4667 1827
rect 4733 1813 4747 1827
rect 4593 1733 4607 1747
rect 4673 1773 4687 1787
rect 4653 1713 4667 1727
rect 4653 1673 4667 1687
rect 4533 1653 4547 1667
rect 4513 1613 4527 1627
rect 4513 1593 4527 1607
rect 4493 1573 4507 1587
rect 4453 1553 4467 1567
rect 4473 1553 4487 1567
rect 4393 1373 4407 1387
rect 4473 1353 4487 1367
rect 4393 1313 4407 1327
rect 4433 1313 4447 1327
rect 4573 1613 4587 1627
rect 4593 1593 4607 1607
rect 4633 1593 4647 1607
rect 4613 1573 4627 1587
rect 4673 1593 4687 1607
rect 4713 1593 4727 1607
rect 4753 1593 4767 1607
rect 4773 1593 4787 1607
rect 4633 1513 4647 1527
rect 4713 1573 4727 1587
rect 4693 1553 4707 1567
rect 4733 1553 4747 1567
rect 4633 1353 4647 1367
rect 4673 1353 4687 1367
rect 4693 1353 4707 1367
rect 4373 1293 4387 1307
rect 4413 1293 4427 1307
rect 4453 1253 4467 1267
rect 4433 1153 4447 1167
rect 4393 1133 4407 1147
rect 4293 1113 4307 1127
rect 4333 1113 4347 1127
rect 4353 1113 4367 1127
rect 4293 1093 4307 1107
rect 4273 1073 4287 1087
rect 4373 1093 4387 1107
rect 4413 1093 4427 1107
rect 4533 1313 4547 1327
rect 4493 1293 4507 1307
rect 4553 1293 4567 1307
rect 4673 1313 4687 1327
rect 4513 1273 4527 1287
rect 4573 1273 4587 1287
rect 4593 1253 4607 1267
rect 4573 1153 4587 1167
rect 4433 1073 4447 1087
rect 4493 1113 4507 1127
rect 4553 1133 4567 1147
rect 4653 1273 4667 1287
rect 4633 1113 4647 1127
rect 4493 1093 4507 1107
rect 4553 1093 4567 1107
rect 4593 1093 4607 1107
rect 4733 1333 4747 1347
rect 4713 1313 4727 1327
rect 4773 1573 4787 1587
rect 4773 1353 4787 1367
rect 4753 1313 4767 1327
rect 4773 1313 4787 1327
rect 4673 1113 4687 1127
rect 4693 1113 4707 1127
rect 4473 1073 4487 1087
rect 4553 1073 4567 1087
rect 4513 1033 4527 1047
rect 4493 913 4507 927
rect 4113 793 4127 807
rect 4073 773 4087 787
rect 4033 673 4047 687
rect 4013 653 4027 667
rect 3953 633 3967 647
rect 3973 613 3987 627
rect 3993 593 4007 607
rect 3913 573 3927 587
rect 3993 533 4007 547
rect 3893 413 3907 427
rect 3833 353 3847 367
rect 3853 333 3867 347
rect 3873 273 3887 287
rect 3933 293 3947 307
rect 3973 293 3987 307
rect 3913 253 3927 267
rect 3833 173 3847 187
rect 3813 153 3827 167
rect 3873 153 3887 167
rect 3893 153 3907 167
rect 3973 253 3987 267
rect 3953 213 3967 227
rect 3233 133 3247 147
rect 3793 133 3807 147
rect 4033 633 4047 647
rect 4033 593 4047 607
rect 4093 633 4107 647
rect 4093 573 4107 587
rect 4073 353 4087 367
rect 4073 333 4087 347
rect 4113 333 4127 347
rect 4033 313 4047 327
rect 4153 793 4167 807
rect 4173 793 4187 807
rect 4153 633 4167 647
rect 4253 813 4267 827
rect 4313 813 4327 827
rect 4193 753 4207 767
rect 4213 713 4227 727
rect 4233 613 4247 627
rect 4273 613 4287 627
rect 4213 593 4227 607
rect 4253 593 4267 607
rect 4453 813 4467 827
rect 4653 1073 4667 1087
rect 4673 1053 4687 1067
rect 4613 913 4627 927
rect 4653 913 4667 927
rect 4553 893 4567 907
rect 4613 873 4627 887
rect 4693 1033 4707 1047
rect 4673 853 4687 867
rect 4753 1133 4767 1147
rect 4733 1113 4747 1127
rect 4753 913 4767 927
rect 4753 893 4767 907
rect 4733 873 4747 887
rect 4413 793 4427 807
rect 4373 773 4387 787
rect 4453 753 4467 767
rect 4393 673 4407 687
rect 4353 613 4367 627
rect 4493 673 4507 687
rect 4433 613 4447 627
rect 4473 513 4487 527
rect 4633 813 4647 827
rect 4633 793 4647 807
rect 4673 793 4687 807
rect 4693 773 4707 787
rect 4293 413 4307 427
rect 4473 413 4487 427
rect 4533 413 4547 427
rect 4273 393 4287 407
rect 4353 393 4367 407
rect 4133 313 4147 327
rect 4113 293 4127 307
rect 4033 253 4047 267
rect 3993 173 4007 187
rect 4013 173 4027 187
rect 3993 153 4007 167
rect 4073 153 4087 167
rect 4253 333 4267 347
rect 4193 273 4207 287
rect 4173 173 4187 187
rect 4193 173 4207 187
rect 4213 153 4227 167
rect 4313 373 4327 387
rect 4373 373 4387 387
rect 4333 353 4347 367
rect 4433 353 4447 367
rect 4393 333 4407 347
rect 4493 353 4507 367
rect 4653 633 4667 647
rect 4673 633 4687 647
rect 4713 633 4727 647
rect 4473 313 4487 327
rect 4413 293 4427 307
rect 4373 213 4387 227
rect 4333 173 4347 187
rect 4053 133 4067 147
rect 4253 133 4267 147
rect 4293 133 4307 147
rect 3913 113 3927 127
rect 3973 113 3987 127
rect 4413 173 4427 187
rect 4453 173 4467 187
rect 4513 193 4527 207
rect 4493 173 4507 187
rect 4513 173 4527 187
rect 4613 173 4627 187
rect 4693 513 4707 527
rect 4673 293 4687 307
rect 4473 153 4487 167
rect 4533 153 4547 167
rect 4433 133 4447 147
rect 4573 133 4587 147
rect 4653 133 4667 147
rect 4753 133 4767 147
rect 4693 113 4707 127
rect 4433 93 4447 107
rect 4733 93 4747 107
rect 2293 73 2307 87
rect 2733 73 2747 87
rect 2813 73 2827 87
rect 1973 13 1987 27
rect 2113 13 2127 27
rect 2153 13 2167 27
<< metal3 >>
rect 4067 4576 4113 4584
rect 4147 4576 4233 4584
rect 4327 4576 4353 4584
rect 1247 4556 1533 4564
rect 4047 4556 4153 4564
rect 127 4536 193 4544
rect 907 4536 1293 4544
rect 1467 4536 1633 4544
rect 2287 4536 2333 4544
rect 3347 4536 3433 4544
rect 3967 4536 4193 4544
rect 47 4516 493 4524
rect 727 4516 1433 4524
rect 1447 4516 1613 4524
rect 1627 4516 1693 4524
rect 1707 4516 1813 4524
rect 1967 4516 2013 4524
rect 2067 4516 2293 4524
rect 3027 4516 3053 4524
rect 3107 4516 3173 4524
rect 3247 4516 3493 4524
rect 3987 4516 4613 4524
rect 87 4496 173 4504
rect 387 4496 433 4504
rect 567 4496 644 4504
rect 187 4476 213 4484
rect 407 4476 444 4484
rect 107 4456 153 4464
rect 167 4456 233 4464
rect 267 4456 313 4464
rect 367 4456 413 4464
rect 436 4464 444 4476
rect 487 4476 604 4484
rect 436 4456 453 4464
rect 467 4456 493 4464
rect 287 4436 373 4444
rect 496 4436 513 4444
rect 527 4436 533 4444
rect 107 4416 153 4424
rect 176 4424 184 4433
rect 176 4416 193 4424
rect 596 4424 604 4476
rect 636 4484 644 4496
rect 667 4496 1053 4504
rect 1087 4496 1113 4504
rect 1147 4496 1273 4504
rect 1327 4496 1353 4504
rect 1376 4496 1453 4504
rect 636 4476 753 4484
rect 787 4476 833 4484
rect 867 4476 984 4484
rect 616 4447 624 4473
rect 707 4456 753 4464
rect 867 4456 933 4464
rect 976 4464 984 4476
rect 1007 4476 1104 4484
rect 1096 4467 1104 4476
rect 1167 4476 1173 4484
rect 1187 4476 1333 4484
rect 1376 4484 1384 4496
rect 1567 4496 1773 4504
rect 1896 4496 1913 4504
rect 1356 4476 1384 4484
rect 976 4456 1033 4464
rect 1047 4456 1084 4464
rect 676 4444 684 4453
rect 667 4436 684 4444
rect 596 4416 633 4424
rect 796 4424 804 4453
rect 816 4427 824 4453
rect 847 4436 864 4444
rect 856 4427 864 4436
rect 887 4436 904 4444
rect 727 4416 804 4424
rect 67 4396 113 4404
rect 127 4396 173 4404
rect 347 4396 693 4404
rect 896 4404 904 4436
rect 967 4436 1013 4444
rect 1076 4444 1084 4456
rect 1107 4456 1193 4464
rect 1356 4464 1364 4476
rect 1407 4476 1484 4484
rect 1287 4456 1364 4464
rect 1476 4464 1484 4476
rect 1507 4476 1573 4484
rect 1896 4484 1904 4496
rect 1927 4496 2173 4504
rect 2196 4496 2393 4504
rect 1587 4476 1904 4484
rect 2196 4484 2204 4496
rect 2407 4496 2473 4504
rect 2947 4496 2993 4504
rect 3007 4496 3113 4504
rect 3127 4496 3133 4504
rect 3187 4496 3413 4504
rect 3427 4496 3464 4504
rect 2007 4476 2204 4484
rect 2227 4476 2324 4484
rect 2316 4467 2324 4476
rect 2516 4484 2524 4493
rect 3456 4487 3464 4496
rect 3647 4496 4133 4504
rect 4167 4496 4333 4504
rect 2447 4476 2524 4484
rect 2667 4476 2793 4484
rect 3016 4476 3144 4484
rect 1476 4456 1553 4464
rect 1607 4456 1653 4464
rect 1907 4456 2013 4464
rect 2147 4456 2193 4464
rect 1076 4436 1133 4444
rect 1376 4444 1384 4453
rect 1267 4436 1384 4444
rect 1527 4436 1693 4444
rect 1847 4436 1973 4444
rect 2267 4436 2353 4444
rect 2376 4444 2384 4473
rect 2616 4464 2624 4473
rect 2467 4456 2624 4464
rect 2727 4456 2973 4464
rect 3016 4464 3024 4476
rect 2987 4456 3024 4464
rect 3087 4456 3113 4464
rect 3136 4464 3144 4476
rect 3287 4476 3353 4484
rect 3367 4476 3373 4484
rect 3587 4476 3713 4484
rect 4127 4476 4273 4484
rect 4327 4476 4513 4484
rect 3136 4456 3253 4464
rect 3267 4456 3293 4464
rect 3407 4456 3693 4464
rect 3747 4456 3793 4464
rect 4247 4456 4293 4464
rect 4687 4456 4713 4464
rect 2376 4436 2493 4444
rect 2547 4436 2673 4444
rect 3036 4444 3044 4453
rect 3036 4436 3073 4444
rect 3667 4436 3773 4444
rect 3787 4436 4093 4444
rect 4187 4436 4293 4444
rect 4627 4436 4733 4444
rect 927 4416 1093 4424
rect 1187 4416 1284 4424
rect 896 4396 1044 4404
rect 667 4376 733 4384
rect 1036 4384 1044 4396
rect 1067 4396 1253 4404
rect 1276 4404 1284 4416
rect 1367 4416 1593 4424
rect 1607 4416 2433 4424
rect 2587 4416 2633 4424
rect 3027 4416 3193 4424
rect 3807 4416 4053 4424
rect 1276 4396 1413 4404
rect 1567 4396 1753 4404
rect 1767 4396 2033 4404
rect 2427 4396 4033 4404
rect 4207 4396 4393 4404
rect 1036 4376 1213 4384
rect 2467 4376 3953 4384
rect 147 4356 553 4364
rect 567 4356 593 4364
rect 607 4356 813 4364
rect 827 4356 913 4364
rect 967 4356 1073 4364
rect 1087 4356 1153 4364
rect 467 4316 573 4324
rect 1807 4316 1893 4324
rect 1907 4316 1933 4324
rect 1947 4316 2093 4324
rect 4047 4296 4093 4304
rect 4107 4296 4133 4304
rect 4687 4296 4733 4304
rect 367 4276 413 4284
rect 2127 4276 3193 4284
rect 1687 4256 2004 4264
rect 47 4236 93 4244
rect 1407 4236 1484 4244
rect 1476 4227 1484 4236
rect 1567 4236 1793 4244
rect 1807 4236 1933 4244
rect 87 4216 124 4224
rect 96 4184 104 4193
rect 87 4176 104 4184
rect 116 4167 124 4216
rect 167 4216 184 4224
rect 176 4204 184 4216
rect 227 4216 264 4224
rect 147 4196 164 4204
rect 176 4196 233 4204
rect 156 4184 164 4196
rect 256 4204 264 4216
rect 327 4216 504 4224
rect 256 4196 284 4204
rect 156 4176 253 4184
rect 276 4184 284 4196
rect 316 4196 413 4204
rect 276 4176 293 4184
rect 316 4167 324 4196
rect 427 4196 473 4204
rect 496 4204 504 4216
rect 667 4216 724 4224
rect 496 4196 513 4204
rect 716 4204 724 4216
rect 807 4216 913 4224
rect 1067 4216 1113 4224
rect 1307 4216 1433 4224
rect 1447 4216 1464 4224
rect 1456 4207 1464 4216
rect 1927 4216 1973 4224
rect 716 4196 773 4204
rect 1247 4196 1313 4204
rect 1467 4196 1553 4204
rect 1747 4196 1813 4204
rect 367 4176 393 4184
rect 696 4184 704 4193
rect 507 4176 813 4184
rect 867 4176 893 4184
rect 956 4184 964 4193
rect 956 4176 1093 4184
rect 1247 4176 1273 4184
rect 1347 4176 1393 4184
rect 1836 4184 1844 4213
rect 1767 4176 1844 4184
rect 567 4156 673 4164
rect 707 4156 713 4164
rect 727 4156 753 4164
rect 887 4156 933 4164
rect 1507 4156 1673 4164
rect 1876 4164 1884 4213
rect 1996 4204 2004 4256
rect 3127 4256 3253 4264
rect 2687 4236 3273 4244
rect 3407 4236 3493 4244
rect 3667 4236 3713 4244
rect 3727 4236 4193 4244
rect 4227 4236 4553 4244
rect 2027 4216 2104 4224
rect 2096 4207 2104 4216
rect 2927 4216 3093 4224
rect 3327 4216 3613 4224
rect 3627 4216 3673 4224
rect 3947 4216 4133 4224
rect 4296 4216 4353 4224
rect 1936 4196 2004 4204
rect 1896 4184 1904 4193
rect 1936 4187 1944 4196
rect 2507 4196 2864 4204
rect 1896 4176 1924 4184
rect 1687 4156 1893 4164
rect 1916 4164 1924 4176
rect 2367 4176 2553 4184
rect 2607 4176 2633 4184
rect 2856 4184 2864 4196
rect 2887 4196 3013 4204
rect 3067 4196 3113 4204
rect 3236 4204 3244 4213
rect 3236 4196 3293 4204
rect 3827 4196 3833 4204
rect 3847 4196 3944 4204
rect 2856 4176 2933 4184
rect 3016 4184 3024 4193
rect 2987 4176 3024 4184
rect 3227 4176 3493 4184
rect 3627 4176 3773 4184
rect 3887 4176 3913 4184
rect 3936 4184 3944 4196
rect 3936 4176 4053 4184
rect 1916 4156 1973 4164
rect 2527 4156 2553 4164
rect 2607 4156 2853 4164
rect 2967 4156 3073 4164
rect 3087 4156 3093 4164
rect 3267 4156 3333 4164
rect 3387 4156 3433 4164
rect 3667 4156 3733 4164
rect 3787 4156 4013 4164
rect 4176 4164 4184 4193
rect 4296 4184 4304 4216
rect 4327 4196 4433 4204
rect 4487 4196 4713 4204
rect 4287 4176 4304 4184
rect 4387 4176 4513 4184
rect 4087 4156 4184 4164
rect 4207 4156 4333 4164
rect 4347 4156 4453 4164
rect 67 4136 293 4144
rect 607 4136 773 4144
rect 907 4136 1033 4144
rect 1047 4136 1133 4144
rect 1207 4136 1453 4144
rect 1867 4136 2073 4144
rect 2927 4136 2953 4144
rect 2967 4136 2993 4144
rect 3927 4136 4493 4144
rect 4507 4136 4513 4144
rect 4527 4136 4593 4144
rect 187 4116 373 4124
rect 527 4116 593 4124
rect 1087 4116 1333 4124
rect 1427 4116 1713 4124
rect 1727 4116 2133 4124
rect 2147 4116 2173 4124
rect 2767 4116 3033 4124
rect 3167 4116 4373 4124
rect 4427 4116 4633 4124
rect 167 4096 433 4104
rect 1367 4096 1413 4104
rect 1627 4096 1653 4104
rect 1667 4096 1713 4104
rect 2007 4096 2073 4104
rect 2087 4096 2313 4104
rect 3567 4096 3693 4104
rect 4047 4096 4213 4104
rect 4247 4096 4293 4104
rect 167 4076 273 4084
rect 287 4076 333 4084
rect 1547 4076 1873 4084
rect 2287 4076 2713 4084
rect 2727 4076 2813 4084
rect 2827 4076 3533 4084
rect 3547 4076 3653 4084
rect 3667 4076 3873 4084
rect 4287 4076 4333 4084
rect 207 4056 293 4064
rect 667 4056 793 4064
rect 807 4056 1073 4064
rect 1827 4056 2253 4064
rect 3367 4056 4033 4064
rect 4047 4056 4073 4064
rect 4107 4056 4133 4064
rect 4147 4056 4193 4064
rect 67 4036 373 4044
rect 427 4036 853 4044
rect 867 4036 933 4044
rect 967 4036 1213 4044
rect 1227 4036 1373 4044
rect 1807 4036 1933 4044
rect 2067 4036 2273 4044
rect 2287 4036 2373 4044
rect 2747 4036 2993 4044
rect 3247 4036 3673 4044
rect 3867 4036 3933 4044
rect 3947 4036 4093 4044
rect 87 4016 213 4024
rect 347 4016 493 4024
rect 507 4016 644 4024
rect 447 3996 513 4004
rect 536 3996 613 4004
rect 267 3976 273 3984
rect 536 3984 544 3996
rect 636 3987 644 4016
rect 727 4016 1233 4024
rect 1247 4016 1353 4024
rect 1367 4016 1433 4024
rect 1487 4016 1544 4024
rect 736 3996 773 4004
rect 287 3976 544 3984
rect 567 3976 624 3984
rect 47 3956 193 3964
rect 276 3964 284 3973
rect 276 3956 353 3964
rect 616 3964 624 3976
rect 676 3964 684 3973
rect 616 3956 684 3964
rect 147 3936 453 3944
rect 467 3936 573 3944
rect 736 3944 744 3996
rect 1007 3996 1013 4004
rect 1407 3996 1513 4004
rect 767 3976 813 3984
rect 956 3976 973 3984
rect 756 3947 764 3973
rect 787 3956 833 3964
rect 667 3936 744 3944
rect 836 3944 844 3953
rect 836 3936 873 3944
rect 956 3944 964 3976
rect 996 3964 1004 3993
rect 1047 3976 1133 3984
rect 1307 3976 1333 3984
rect 987 3956 1004 3964
rect 1107 3956 1193 3964
rect 1407 3956 1453 3964
rect 1536 3964 1544 4016
rect 1667 4016 1813 4024
rect 1927 4016 1953 4024
rect 2407 4016 2433 4024
rect 2587 4016 3053 4024
rect 3087 4016 3213 4024
rect 3227 4016 3273 4024
rect 3287 4016 3313 4024
rect 3347 4016 3453 4024
rect 3487 4016 3753 4024
rect 3836 4016 3913 4024
rect 1607 3996 1633 4004
rect 1687 3996 1693 4004
rect 1707 3996 1753 4004
rect 2287 3996 2353 4004
rect 3107 3996 3244 4004
rect 1507 3956 1544 3964
rect 956 3936 1033 3944
rect 1427 3936 1473 3944
rect 1487 3936 1533 3944
rect 1776 3944 1784 3993
rect 1836 3967 1844 3993
rect 1927 3976 1973 3984
rect 2107 3976 2153 3984
rect 2227 3976 2293 3984
rect 2776 3984 2784 3993
rect 2627 3976 2784 3984
rect 2927 3976 2973 3984
rect 3027 3976 3153 3984
rect 3236 3984 3244 3996
rect 3387 3996 3413 4004
rect 3707 3996 3813 4004
rect 3236 3976 3253 3984
rect 3356 3967 3364 3993
rect 3436 3984 3444 3993
rect 3836 3987 3844 4016
rect 4027 4016 4153 4024
rect 3856 3996 3893 4004
rect 3856 3987 3864 3996
rect 4007 3996 4053 4004
rect 4127 3996 4184 4004
rect 4176 3987 4184 3996
rect 4207 3996 4273 4004
rect 4307 3996 4553 4004
rect 3376 3976 3513 3984
rect 3376 3967 3384 3976
rect 4227 3976 4313 3984
rect 4427 3976 4673 3984
rect 4687 3976 4713 3984
rect 1867 3956 1993 3964
rect 2687 3956 2773 3964
rect 2947 3956 3133 3964
rect 3687 3956 3973 3964
rect 4647 3956 4824 3964
rect 1776 3936 1813 3944
rect 3187 3936 3573 3944
rect 3587 3936 3853 3944
rect 267 3916 433 3924
rect 447 3916 533 3924
rect 707 3916 853 3924
rect 2387 3916 3633 3924
rect 3827 3916 3873 3924
rect 3887 3916 4633 3924
rect 67 3896 313 3904
rect 327 3896 393 3904
rect 547 3896 593 3904
rect 1127 3896 1233 3904
rect 1247 3896 1273 3904
rect 2487 3896 3773 3904
rect 167 3876 173 3884
rect 187 3876 373 3884
rect 1347 3856 1513 3864
rect 1527 3856 1573 3864
rect 4247 3856 4293 3864
rect 3687 3836 4053 3844
rect 4067 3836 4313 3844
rect 887 3796 1033 3804
rect 1047 3796 1173 3804
rect 847 3776 953 3784
rect 427 3756 593 3764
rect 647 3756 993 3764
rect 916 3747 924 3756
rect 1427 3756 1633 3764
rect 1907 3756 1953 3764
rect 3167 3756 3513 3764
rect 3527 3756 3613 3764
rect 4507 3756 4533 3764
rect 4547 3756 4693 3764
rect 407 3736 513 3744
rect 676 3736 844 3744
rect 56 3687 64 3713
rect 76 3707 84 3733
rect 116 3687 124 3713
rect 136 3704 144 3733
rect 167 3716 213 3724
rect 367 3716 493 3724
rect 136 3696 153 3704
rect 296 3704 304 3713
rect 236 3696 304 3704
rect 336 3704 344 3713
rect 516 3707 524 3733
rect 676 3724 684 3736
rect 587 3716 684 3724
rect 747 3716 793 3724
rect 836 3724 844 3736
rect 956 3736 1024 3744
rect 956 3724 964 3736
rect 836 3716 964 3724
rect 1016 3724 1024 3736
rect 1047 3736 1073 3744
rect 1127 3736 1373 3744
rect 1387 3736 1573 3744
rect 1987 3736 2153 3744
rect 2347 3736 2473 3744
rect 3287 3736 3393 3744
rect 3547 3736 3573 3744
rect 4216 3736 4253 3744
rect 1016 3716 1053 3724
rect 1107 3716 1193 3724
rect 1287 3716 1353 3724
rect 1447 3716 1493 3724
rect 1547 3716 1593 3724
rect 1936 3724 1944 3733
rect 1936 3716 2053 3724
rect 2327 3716 2633 3724
rect 3227 3716 3273 3724
rect 3307 3716 3313 3724
rect 3347 3716 3444 3724
rect 336 3696 353 3704
rect 236 3687 244 3696
rect 547 3696 573 3704
rect 267 3676 313 3684
rect 327 3676 413 3684
rect 676 3684 684 3693
rect 696 3687 704 3713
rect 767 3696 933 3704
rect 976 3704 984 3713
rect 976 3696 1013 3704
rect 1067 3696 1133 3704
rect 1487 3696 1513 3704
rect 1676 3704 1684 3713
rect 1567 3696 1684 3704
rect 1707 3696 1713 3704
rect 1727 3696 1733 3704
rect 1756 3687 1764 3713
rect 1787 3696 1813 3704
rect 1827 3696 1953 3704
rect 2147 3696 2373 3704
rect 2507 3696 2533 3704
rect 2547 3696 2613 3704
rect 2676 3687 2684 3713
rect 2727 3696 2873 3704
rect 2976 3704 2984 3713
rect 2927 3696 2984 3704
rect 3156 3704 3164 3713
rect 3156 3696 3253 3704
rect 3316 3704 3324 3713
rect 3316 3696 3344 3704
rect 427 3676 684 3684
rect 847 3676 913 3684
rect 947 3676 973 3684
rect 1087 3676 1173 3684
rect 1227 3676 1253 3684
rect 1407 3676 1413 3684
rect 1427 3676 1453 3684
rect 1587 3676 1613 3684
rect 1627 3676 1653 3684
rect 1887 3676 1913 3684
rect 1967 3676 1993 3684
rect 2467 3676 2653 3684
rect 2767 3676 2793 3684
rect 2907 3676 2953 3684
rect 3087 3676 3193 3684
rect 3336 3684 3344 3696
rect 3436 3687 3444 3716
rect 3907 3716 4193 3724
rect 3716 3704 3724 3713
rect 3567 3696 3724 3704
rect 3747 3696 3873 3704
rect 4216 3704 4224 3736
rect 4247 3716 4273 3724
rect 4647 3716 4773 3724
rect 4196 3696 4224 3704
rect 4196 3687 4204 3696
rect 4267 3696 4433 3704
rect 4816 3704 4824 3724
rect 4796 3696 4824 3704
rect 3336 3676 3373 3684
rect 3707 3676 3773 3684
rect 3807 3676 4073 3684
rect 4796 3684 4804 3696
rect 4687 3676 4804 3684
rect 87 3656 133 3664
rect 187 3656 373 3664
rect 527 3656 933 3664
rect 1267 3656 1553 3664
rect 1847 3656 2393 3664
rect 2607 3656 2753 3664
rect 2967 3656 3113 3664
rect 3127 3656 3353 3664
rect 3467 3656 3813 3664
rect 4127 3656 4213 3664
rect 4816 3664 4824 3684
rect 4667 3656 4824 3664
rect 67 3636 93 3644
rect 247 3636 313 3644
rect 447 3636 453 3644
rect 467 3636 793 3644
rect 1087 3636 1373 3644
rect 1387 3636 1633 3644
rect 1647 3636 1913 3644
rect 2827 3636 2993 3644
rect 3007 3636 3133 3644
rect 3407 3636 3633 3644
rect 4187 3636 4293 3644
rect 47 3616 93 3624
rect 127 3616 373 3624
rect 387 3616 693 3624
rect 767 3616 1133 3624
rect 1147 3616 1573 3624
rect 1947 3616 2373 3624
rect 2787 3616 2913 3624
rect 3307 3616 3413 3624
rect 3427 3616 3433 3624
rect 4167 3616 4273 3624
rect 4327 3616 4413 3624
rect 127 3596 644 3604
rect 347 3576 353 3584
rect 367 3576 533 3584
rect 547 3576 593 3584
rect 636 3584 644 3596
rect 667 3596 1073 3604
rect 1107 3596 1533 3604
rect 2007 3596 2153 3604
rect 2167 3596 2313 3604
rect 3067 3596 3493 3604
rect 3507 3596 3593 3604
rect 3827 3596 4093 3604
rect 4187 3596 4353 3604
rect 4387 3596 4413 3604
rect 636 3576 993 3584
rect 1127 3576 1153 3584
rect 2187 3576 2493 3584
rect 3187 3576 3653 3584
rect 3927 3576 4053 3584
rect -24 3544 -16 3564
rect 687 3556 733 3564
rect 987 3556 1273 3564
rect 1607 3556 2173 3564
rect 2307 3556 2433 3564
rect 2587 3556 2713 3564
rect 3227 3556 3273 3564
rect 3367 3556 3393 3564
rect 3487 3556 3533 3564
rect 3547 3556 3573 3564
rect 3587 3556 3673 3564
rect 4047 3556 4153 3564
rect -44 3536 -16 3544
rect -44 3444 -36 3536
rect 187 3536 513 3544
rect 576 3536 753 3544
rect -24 3504 -16 3524
rect 487 3516 553 3524
rect -24 3496 373 3504
rect 447 3496 493 3504
rect 576 3504 584 3536
rect 847 3536 873 3544
rect 1027 3536 1053 3544
rect 1107 3536 1233 3544
rect 1396 3536 1684 3544
rect 1396 3524 1404 3536
rect 1676 3527 1684 3536
rect 1707 3536 1793 3544
rect 1847 3536 2113 3544
rect 2387 3536 2433 3544
rect 2547 3536 3033 3544
rect 3167 3536 3213 3544
rect 3247 3536 3313 3544
rect 3327 3536 3333 3544
rect 3356 3536 3413 3544
rect 1007 3516 1404 3524
rect 1427 3516 1553 3524
rect 1727 3516 1793 3524
rect 2127 3516 2153 3524
rect 2167 3516 2233 3524
rect 2687 3516 2813 3524
rect 2827 3516 2833 3524
rect 2847 3516 2933 3524
rect 2947 3516 3064 3524
rect 547 3496 584 3504
rect -24 3476 13 3484
rect 87 3476 113 3484
rect 656 3484 664 3513
rect 836 3504 844 3513
rect 836 3496 873 3504
rect 907 3496 1013 3504
rect 1047 3496 1113 3504
rect 1167 3496 1233 3504
rect 1327 3496 1433 3504
rect 1767 3496 1853 3504
rect 2007 3496 2124 3504
rect 567 3476 664 3484
rect 696 3467 704 3493
rect 2116 3487 2124 3496
rect 2267 3496 2333 3504
rect 2407 3496 2693 3504
rect 2747 3496 2873 3504
rect 3056 3504 3064 3516
rect 3087 3516 3133 3524
rect 3187 3516 3253 3524
rect 3356 3524 3364 3536
rect 3447 3536 3464 3544
rect 3336 3516 3364 3524
rect 3456 3524 3464 3536
rect 3487 3536 3513 3544
rect 3556 3536 3653 3544
rect 3456 3516 3504 3524
rect 3056 3496 3193 3504
rect 3336 3504 3344 3516
rect 3247 3496 3344 3504
rect 3407 3496 3433 3504
rect 3496 3487 3504 3516
rect 3556 3507 3564 3536
rect 3767 3536 3913 3544
rect 3967 3536 4033 3544
rect 3627 3516 3804 3524
rect 3796 3507 3804 3516
rect 3867 3516 3953 3524
rect 4067 3516 4293 3524
rect 4307 3516 4393 3524
rect 4487 3516 4633 3524
rect 3727 3496 3753 3504
rect 4407 3496 4453 3504
rect 4567 3496 4653 3504
rect 4676 3487 4684 3513
rect 4707 3496 4753 3504
rect 1007 3476 1033 3484
rect 1107 3476 1193 3484
rect 1267 3476 1293 3484
rect 1347 3476 1373 3484
rect 1607 3476 1673 3484
rect 1687 3476 1893 3484
rect 1927 3476 1953 3484
rect 1967 3476 1973 3484
rect 2907 3476 2953 3484
rect 3187 3476 3293 3484
rect 3567 3476 3693 3484
rect 3707 3476 4593 3484
rect 387 3456 413 3464
rect 427 3456 673 3464
rect 796 3456 1733 3464
rect -44 3436 93 3444
rect 796 3444 804 3456
rect 1767 3456 1813 3464
rect 2027 3456 2093 3464
rect 3007 3456 3233 3464
rect 3787 3456 3833 3464
rect 3847 3456 3893 3464
rect 3947 3456 4013 3464
rect 4027 3456 4333 3464
rect 4367 3456 4653 3464
rect 307 3436 804 3444
rect 827 3436 1073 3444
rect 1867 3436 1893 3444
rect 3847 3436 4073 3444
rect 27 3416 1253 3424
rect 1687 3416 2093 3424
rect 2767 3416 4153 3424
rect 4167 3416 4213 3424
rect 27 3396 293 3404
rect 627 3396 853 3404
rect 947 3396 1013 3404
rect 1227 3396 1473 3404
rect 1487 3396 1713 3404
rect 1727 3396 1773 3404
rect 3307 3396 3873 3404
rect 727 3376 753 3384
rect 767 3376 1004 3384
rect 267 3356 533 3364
rect 687 3356 733 3364
rect 927 3356 973 3364
rect 996 3364 1004 3376
rect 1107 3376 1673 3384
rect 1807 3376 1973 3384
rect 996 3356 1373 3364
rect 1396 3356 1713 3364
rect 267 3336 633 3344
rect 787 3336 1093 3344
rect 1396 3344 1404 3356
rect 1747 3356 1933 3364
rect 2367 3356 2513 3364
rect 1147 3336 1404 3344
rect 1447 3336 2153 3344
rect 3487 3336 3533 3344
rect 327 3316 393 3324
rect 467 3316 513 3324
rect 527 3316 1213 3324
rect 1647 3316 2133 3324
rect 3167 3316 3473 3324
rect 3607 3316 3773 3324
rect 4087 3316 4493 3324
rect 467 3296 553 3304
rect 607 3296 824 3304
rect 47 3276 293 3284
rect 347 3276 393 3284
rect 407 3276 793 3284
rect 816 3284 824 3296
rect 847 3296 1133 3304
rect 1187 3296 1833 3304
rect 2287 3296 2333 3304
rect 2347 3296 2393 3304
rect 3287 3296 3573 3304
rect 3607 3296 3633 3304
rect 4467 3296 4633 3304
rect 816 3276 913 3284
rect 1007 3276 1813 3284
rect 1827 3276 1953 3284
rect 1967 3276 2033 3284
rect 2287 3276 2353 3284
rect 3107 3276 3213 3284
rect 3907 3276 3913 3284
rect 3927 3276 3953 3284
rect 3987 3276 4013 3284
rect 4447 3276 4513 3284
rect 4636 3276 4673 3284
rect 127 3256 364 3264
rect 96 3227 104 3253
rect 156 3236 173 3244
rect 156 3224 164 3236
rect 356 3227 364 3256
rect 447 3256 473 3264
rect 487 3256 593 3264
rect 667 3256 813 3264
rect 856 3256 873 3264
rect 387 3236 413 3244
rect 856 3227 864 3256
rect 896 3256 953 3264
rect 896 3244 904 3256
rect 967 3256 1053 3264
rect 1067 3256 1173 3264
rect 1267 3256 1273 3264
rect 1287 3256 1364 3264
rect 1356 3247 1364 3256
rect 1507 3256 1513 3264
rect 1527 3256 1593 3264
rect 1707 3256 1824 3264
rect 887 3236 904 3244
rect 947 3236 993 3244
rect 1056 3236 1073 3244
rect 116 3216 164 3224
rect 27 3196 93 3204
rect 116 3184 124 3216
rect 187 3216 213 3224
rect 447 3216 473 3224
rect 607 3216 733 3224
rect 1056 3224 1064 3236
rect 1287 3236 1313 3244
rect 907 3216 1064 3224
rect 1087 3216 1113 3224
rect 1396 3224 1404 3253
rect 1567 3236 1613 3244
rect 1127 3216 1404 3224
rect 1447 3216 1533 3224
rect 1636 3224 1644 3253
rect 1636 3216 1693 3224
rect 1727 3216 1793 3224
rect 147 3196 233 3204
rect 247 3196 353 3204
rect 367 3196 553 3204
rect 747 3196 793 3204
rect 827 3196 833 3204
rect 847 3196 1173 3204
rect 1347 3196 1453 3204
rect 1567 3196 1713 3204
rect 1816 3204 1824 3256
rect 1907 3256 1973 3264
rect 1836 3244 1844 3253
rect 1916 3244 1924 3256
rect 2127 3256 2264 3264
rect 1836 3236 1904 3244
rect 1916 3236 2044 3244
rect 1896 3227 1904 3236
rect 2036 3227 2044 3236
rect 2076 3227 2084 3253
rect 2256 3247 2264 3256
rect 2307 3256 2404 3264
rect 2116 3236 2133 3244
rect 2116 3227 2124 3236
rect 2167 3236 2204 3244
rect 2196 3227 2204 3236
rect 1847 3216 1873 3224
rect 1816 3196 1833 3204
rect 1936 3204 1944 3213
rect 1887 3196 1944 3204
rect 2216 3204 2224 3233
rect 2247 3216 2273 3224
rect 2336 3207 2344 3233
rect 2396 3227 2404 3256
rect 3376 3256 3433 3264
rect 2967 3236 3013 3244
rect 3067 3236 3093 3244
rect 3136 3227 3144 3253
rect 3167 3236 3293 3244
rect 3307 3236 3353 3244
rect 3376 3227 3384 3256
rect 3547 3256 3613 3264
rect 3887 3256 4033 3264
rect 4156 3256 4284 3264
rect 3696 3244 3704 3253
rect 3607 3236 3704 3244
rect 3956 3236 4013 3244
rect 3956 3227 3964 3236
rect 4156 3244 4164 3256
rect 4076 3236 4164 3244
rect 2787 3216 2833 3224
rect 2847 3216 2973 3224
rect 3047 3216 3113 3224
rect 3247 3216 3313 3224
rect 3467 3216 3753 3224
rect 4076 3224 4084 3236
rect 4007 3216 4084 3224
rect 4176 3224 4184 3233
rect 4107 3216 4184 3224
rect 4207 3216 4233 3224
rect 2087 3196 2224 3204
rect 2456 3187 2464 3213
rect 4256 3207 4264 3233
rect 4276 3227 4284 3256
rect 4296 3256 4313 3264
rect 2567 3196 2853 3204
rect 3047 3196 3093 3204
rect 3187 3196 3273 3204
rect 3407 3196 3473 3204
rect 4027 3196 4113 3204
rect 4296 3204 4304 3256
rect 4416 3264 4424 3273
rect 4347 3256 4404 3264
rect 4416 3256 4473 3264
rect 4287 3196 4304 3204
rect 4376 3204 4384 3233
rect 4396 3224 4404 3256
rect 4427 3236 4493 3244
rect 4396 3216 4413 3224
rect 4347 3196 4384 3204
rect 116 3176 133 3184
rect 167 3176 313 3184
rect 347 3176 373 3184
rect 467 3176 593 3184
rect 667 3176 773 3184
rect 887 3176 1493 3184
rect 1527 3176 1993 3184
rect 2727 3176 3073 3184
rect 3987 3176 4173 3184
rect 4187 3176 4353 3184
rect 4367 3176 4433 3184
rect 4636 3184 4644 3276
rect 4656 3207 4664 3253
rect 4687 3236 4733 3244
rect 4707 3216 4733 3224
rect 4636 3176 4733 3184
rect 107 3156 393 3164
rect 467 3156 573 3164
rect 627 3156 653 3164
rect 767 3156 873 3164
rect 947 3156 973 3164
rect 1147 3156 1213 3164
rect 1247 3156 1413 3164
rect 1487 3156 1613 3164
rect 1707 3156 1773 3164
rect 1807 3156 2664 3164
rect 147 3136 293 3144
rect 647 3136 673 3144
rect 1127 3136 1393 3144
rect 1747 3136 1813 3144
rect 1927 3136 1973 3144
rect 2387 3136 2633 3144
rect 2656 3144 2664 3156
rect 2687 3156 2773 3164
rect 2907 3156 3333 3164
rect 3356 3156 3813 3164
rect 3356 3144 3364 3156
rect 3847 3156 4013 3164
rect 4067 3156 4213 3164
rect 4267 3156 4393 3164
rect 2656 3136 3364 3144
rect 3587 3136 3633 3144
rect 3927 3136 3993 3144
rect 4007 3136 4253 3144
rect 4307 3136 4373 3144
rect 247 3116 273 3124
rect 287 3116 433 3124
rect 927 3116 1213 3124
rect 1747 3116 1953 3124
rect 2167 3116 2513 3124
rect 2987 3116 3253 3124
rect 3867 3116 3993 3124
rect 4027 3116 4073 3124
rect 4247 3116 4293 3124
rect 4367 3116 4393 3124
rect 487 3096 553 3104
rect 587 3096 593 3104
rect 607 3096 784 3104
rect 76 3076 253 3084
rect 36 3007 44 3033
rect 76 3007 84 3076
rect 527 3076 593 3084
rect 776 3084 784 3096
rect 807 3096 993 3104
rect 1016 3096 1073 3104
rect 1016 3084 1024 3096
rect 1187 3096 1324 3104
rect 776 3076 1024 3084
rect 1047 3076 1193 3084
rect 1267 3076 1293 3084
rect 1316 3084 1324 3096
rect 1507 3096 1653 3104
rect 1667 3096 1753 3104
rect 1767 3096 1853 3104
rect 1887 3096 2033 3104
rect 2047 3096 2173 3104
rect 2367 3096 2713 3104
rect 2867 3096 2873 3104
rect 2887 3096 2893 3104
rect 3407 3096 3633 3104
rect 3727 3096 4113 3104
rect 4667 3096 4804 3104
rect 1316 3076 1473 3084
rect 1527 3076 1713 3084
rect 1727 3076 2093 3084
rect 2107 3076 2133 3084
rect 2287 3076 2453 3084
rect 2867 3076 3113 3084
rect 3167 3076 3373 3084
rect 3507 3076 3713 3084
rect 3787 3076 3924 3084
rect 96 3056 153 3064
rect 96 3027 104 3056
rect 356 3056 533 3064
rect -24 2964 -16 3004
rect 116 3004 124 3033
rect 276 3016 293 3024
rect 116 2996 213 3004
rect 67 2976 93 2984
rect 276 2984 284 3016
rect 356 3004 364 3056
rect 847 3056 1013 3064
rect 1187 3056 1784 3064
rect 387 3036 513 3044
rect 607 3036 724 3044
rect 547 3016 593 3024
rect 307 2996 364 3004
rect 387 2996 573 3004
rect 587 2996 673 3004
rect 276 2976 473 2984
rect 696 2984 704 3013
rect 716 3007 724 3036
rect 767 3036 833 3044
rect 1156 3044 1164 3053
rect 1156 3036 1224 3044
rect 856 3024 864 3033
rect 816 3016 864 3024
rect 976 3024 984 3033
rect 976 3016 1173 3024
rect 816 3007 824 3016
rect 947 2996 993 3004
rect 1216 3004 1224 3036
rect 1536 3036 1573 3044
rect 1276 3024 1284 3033
rect 1247 3016 1513 3024
rect 1216 2996 1253 3004
rect 1287 2996 1413 3004
rect 1427 2996 1473 3004
rect 1536 3004 1544 3036
rect 1627 3036 1753 3044
rect 1776 3027 1784 3056
rect 2127 3056 2384 3064
rect 1796 3036 1893 3044
rect 1567 3016 1704 3024
rect 1696 3007 1704 3016
rect 1796 3007 1804 3036
rect 1936 3024 1944 3053
rect 2147 3036 2193 3044
rect 2247 3036 2293 3044
rect 2336 3036 2353 3044
rect 1887 3016 1944 3024
rect 2067 3016 2073 3024
rect 2087 3016 2113 3024
rect 2167 3016 2213 3024
rect 1536 2996 1553 3004
rect 687 2976 704 2984
rect 787 2976 893 2984
rect 907 2976 1233 2984
rect 1407 2976 1453 2984
rect 1547 2976 1573 2984
rect 1816 2984 1824 3013
rect 1847 2996 1973 3004
rect 2087 2996 2293 3004
rect 1667 2976 1824 2984
rect 2316 2984 2324 3013
rect 2336 3007 2344 3036
rect 2376 3027 2384 3056
rect 2627 3056 2753 3064
rect 2767 3056 2793 3064
rect 3067 3056 3093 3064
rect 3596 3056 3673 3064
rect 2436 3044 2444 3053
rect 2396 3036 2444 3044
rect 2396 3007 2404 3036
rect 2527 3036 2653 3044
rect 2667 3036 2673 3044
rect 3087 3036 3193 3044
rect 2427 3016 2453 3024
rect 2487 3016 2533 3024
rect 2696 3004 2704 3033
rect 3036 3024 3044 3033
rect 3176 3027 3184 3036
rect 3036 3016 3153 3024
rect 3216 3024 3224 3053
rect 3367 3036 3433 3044
rect 3196 3016 3224 3024
rect 2547 2996 2704 3004
rect 2316 2976 2453 2984
rect 2716 2984 2724 3013
rect 2747 2996 2833 3004
rect 3007 2996 3033 3004
rect 3196 3004 3204 3016
rect 3507 3016 3533 3024
rect 3147 2996 3204 3004
rect 3307 2996 3393 3004
rect 2607 2976 2724 2984
rect 2987 2976 3053 2984
rect 3067 2976 3253 2984
rect 3596 2984 3604 3056
rect 3916 3064 3924 3076
rect 3987 3076 4013 3084
rect 4047 3076 4133 3084
rect 4147 3076 4313 3084
rect 4376 3076 4413 3084
rect 3916 3056 4093 3064
rect 4107 3056 4193 3064
rect 4207 3056 4233 3064
rect 4247 3056 4333 3064
rect 3647 3036 3673 3044
rect 3727 3036 3753 3044
rect 3896 3044 3904 3053
rect 3867 3036 3884 3044
rect 3896 3036 3944 3044
rect 3627 3016 3773 3024
rect 3796 3024 3804 3033
rect 3787 3016 3804 3024
rect 3827 3016 3853 3024
rect 3876 3024 3884 3036
rect 3876 3016 3893 3024
rect 3936 3024 3944 3036
rect 3967 3036 3984 3044
rect 3936 3016 3964 3024
rect 3667 2996 3713 3004
rect 3596 2976 3713 2984
rect 3956 2984 3964 3016
rect 3976 3007 3984 3036
rect 4087 3036 4144 3044
rect 4007 3016 4024 3024
rect 4016 3004 4024 3016
rect 4067 3016 4113 3024
rect 4136 3007 4144 3036
rect 4256 3036 4293 3044
rect 4176 3007 4184 3033
rect 4256 3024 4264 3036
rect 4316 3036 4353 3044
rect 4247 3016 4264 3024
rect 4276 3016 4293 3024
rect 4016 2996 4113 3004
rect 4276 2987 4284 3016
rect 4316 3004 4324 3036
rect 4376 3044 4384 3076
rect 4487 3076 4493 3084
rect 4507 3076 4633 3084
rect 4667 3076 4773 3084
rect 4407 3056 4544 3064
rect 4536 3047 4544 3056
rect 4687 3056 4733 3064
rect 4796 3064 4804 3096
rect 4787 3056 4804 3064
rect 4376 3036 4404 3044
rect 4396 3024 4404 3036
rect 4427 3036 4444 3044
rect 4396 3016 4413 3024
rect 4436 3024 4444 3036
rect 4627 3036 4673 3044
rect 4436 3016 4613 3024
rect 4707 3016 4733 3024
rect 4296 2996 4324 3004
rect 4296 2987 4304 2996
rect 4367 2996 4593 3004
rect 4607 2996 4653 3004
rect 4667 2996 4673 3004
rect 3956 2976 4093 2984
rect 4567 2976 4693 2984
rect -24 2956 373 2964
rect 447 2956 693 2964
rect 727 2956 873 2964
rect 1027 2956 1053 2964
rect 1307 2956 1593 2964
rect 1627 2956 2013 2964
rect 3387 2956 3813 2964
rect 4167 2956 4413 2964
rect 27 2936 173 2944
rect 507 2936 613 2944
rect 627 2936 753 2944
rect 967 2936 1093 2944
rect 1107 2936 1793 2944
rect 3107 2936 3433 2944
rect 4247 2936 4313 2944
rect 67 2916 313 2924
rect 567 2916 1453 2924
rect 1507 2916 1693 2924
rect 3747 2916 3773 2924
rect 4287 2916 4613 2924
rect 4627 2916 4773 2924
rect 267 2896 573 2904
rect 667 2896 873 2904
rect 896 2896 1693 2904
rect 896 2884 904 2896
rect 367 2876 904 2884
rect 1127 2876 1173 2884
rect 1367 2876 1673 2884
rect 1767 2876 3093 2884
rect 3647 2876 3833 2884
rect 3847 2876 4433 2884
rect 207 2856 1553 2864
rect 1567 2856 2773 2864
rect 2787 2856 2993 2864
rect 3687 2856 4273 2864
rect 4287 2856 4473 2864
rect 87 2836 553 2844
rect 627 2836 733 2844
rect 867 2836 893 2844
rect 907 2836 1573 2844
rect 1587 2836 1913 2844
rect 2267 2836 2953 2844
rect 3827 2836 4253 2844
rect 247 2816 273 2824
rect 567 2816 624 2824
rect 347 2796 444 2804
rect 27 2776 133 2784
rect 307 2776 353 2784
rect 387 2776 424 2784
rect -24 2684 -16 2764
rect 36 2727 44 2753
rect 56 2744 64 2753
rect 56 2736 113 2744
rect 156 2744 164 2773
rect 156 2736 173 2744
rect 196 2727 204 2753
rect 216 2724 224 2773
rect 247 2756 393 2764
rect 416 2747 424 2776
rect 436 2764 444 2796
rect 616 2804 624 2816
rect 687 2816 833 2824
rect 1067 2816 1133 2824
rect 1327 2816 1613 2824
rect 1707 2816 2493 2824
rect 3787 2816 3933 2824
rect 4047 2816 4133 2824
rect 616 2796 664 2804
rect 436 2756 493 2764
rect 267 2736 273 2744
rect 287 2736 373 2744
rect 447 2736 493 2744
rect 536 2744 544 2793
rect 576 2747 584 2773
rect 656 2764 664 2796
rect 767 2796 1193 2804
rect 1207 2796 1373 2804
rect 1387 2796 1753 2804
rect 1787 2796 1893 2804
rect 2027 2796 2053 2804
rect 2247 2796 2473 2804
rect 2507 2796 2633 2804
rect 2827 2796 3093 2804
rect 3107 2796 3853 2804
rect 4567 2796 4613 2804
rect 4627 2796 4673 2804
rect 636 2756 664 2764
rect 536 2736 553 2744
rect 636 2744 644 2756
rect 627 2736 644 2744
rect 716 2744 724 2793
rect 827 2776 953 2784
rect 1107 2776 1193 2784
rect 1267 2776 1404 2784
rect 847 2756 1004 2764
rect 687 2736 724 2744
rect 747 2736 764 2744
rect 216 2716 293 2724
rect 367 2716 533 2724
rect 756 2724 764 2736
rect 827 2736 853 2744
rect 907 2736 913 2744
rect 927 2736 973 2744
rect 996 2744 1004 2756
rect 1027 2756 1353 2764
rect 996 2736 1053 2744
rect 1087 2736 1153 2744
rect 1187 2736 1373 2744
rect 756 2716 804 2724
rect 27 2696 53 2704
rect 67 2696 213 2704
rect 347 2696 613 2704
rect 667 2696 773 2704
rect 796 2704 804 2716
rect 1027 2716 1293 2724
rect 1396 2724 1404 2776
rect 1987 2776 2213 2784
rect 2367 2776 2433 2784
rect 2487 2776 2553 2784
rect 2567 2776 2593 2784
rect 2867 2776 2913 2784
rect 3496 2776 3533 2784
rect 1636 2764 1644 2773
rect 1467 2756 1813 2764
rect 1836 2747 1844 2773
rect 1867 2756 1893 2764
rect 1947 2756 2153 2764
rect 2216 2756 2273 2764
rect 1867 2736 1993 2744
rect 2216 2744 2224 2756
rect 2347 2756 2373 2764
rect 2556 2756 2633 2764
rect 2147 2736 2224 2744
rect 2416 2744 2424 2753
rect 2556 2747 2564 2756
rect 2787 2756 2833 2764
rect 2416 2736 2433 2744
rect 2527 2736 2553 2744
rect 2736 2744 2744 2753
rect 3496 2747 3504 2776
rect 3567 2776 3593 2784
rect 3607 2776 3653 2784
rect 3807 2776 3893 2784
rect 3956 2776 4144 2784
rect 2587 2736 2744 2744
rect 2767 2736 2973 2744
rect 3607 2736 3653 2744
rect 3956 2744 3964 2776
rect 4136 2767 4144 2776
rect 4196 2776 4213 2784
rect 3987 2756 4024 2764
rect 3887 2736 3964 2744
rect 4016 2744 4024 2756
rect 4196 2764 4204 2776
rect 4507 2776 4633 2784
rect 4176 2756 4204 2764
rect 4016 2736 4044 2744
rect 1316 2716 1404 2724
rect 1756 2724 1764 2733
rect 1756 2716 1893 2724
rect 796 2696 1033 2704
rect 1047 2696 1113 2704
rect 1127 2696 1213 2704
rect 1316 2704 1324 2716
rect 1907 2716 2093 2724
rect 2207 2716 2253 2724
rect 2267 2716 2313 2724
rect 2667 2716 2713 2724
rect 2887 2716 3013 2724
rect 3027 2716 3253 2724
rect 3427 2716 3433 2724
rect 3447 2716 3833 2724
rect 3987 2716 4013 2724
rect 4036 2724 4044 2736
rect 4176 2744 4184 2756
rect 4636 2747 4644 2773
rect 4067 2736 4184 2744
rect 4387 2736 4573 2744
rect 4687 2736 4753 2744
rect 4036 2716 4053 2724
rect 4127 2716 4173 2724
rect 4207 2716 4233 2724
rect 4287 2716 4413 2724
rect 4447 2716 4533 2724
rect 4607 2716 4653 2724
rect 1267 2696 1324 2704
rect 1647 2696 1853 2704
rect 1967 2696 2053 2704
rect 2287 2696 2453 2704
rect 2467 2696 2533 2704
rect 2727 2696 2793 2704
rect 3127 2696 3213 2704
rect 3507 2696 3733 2704
rect 3747 2696 3853 2704
rect 3867 2696 3893 2704
rect 3947 2696 3993 2704
rect 4087 2696 4113 2704
rect 4247 2696 4313 2704
rect 4567 2696 4693 2704
rect -24 2676 1133 2684
rect 1147 2676 1473 2684
rect 1496 2676 1693 2684
rect 67 2656 93 2664
rect 107 2656 313 2664
rect 427 2656 813 2664
rect 847 2656 973 2664
rect 1107 2656 1313 2664
rect 1496 2664 1504 2676
rect 1787 2676 1913 2684
rect 2047 2676 2093 2684
rect 2127 2676 2293 2684
rect 2307 2676 2633 2684
rect 3047 2676 3213 2684
rect 3227 2676 3453 2684
rect 4167 2676 4513 2684
rect 1347 2656 1504 2664
rect 1667 2656 1833 2664
rect 2287 2656 2513 2664
rect 3167 2656 3533 2664
rect 3807 2656 4133 2664
rect 807 2636 933 2644
rect 1007 2636 1133 2644
rect 1167 2636 1233 2644
rect 1687 2636 2073 2644
rect 2207 2636 2293 2644
rect 2307 2636 2393 2644
rect 3007 2636 3453 2644
rect 3487 2636 3613 2644
rect 4007 2636 4213 2644
rect 4227 2636 4393 2644
rect 107 2616 173 2624
rect 187 2616 353 2624
rect 447 2616 613 2624
rect 807 2616 853 2624
rect 867 2616 1033 2624
rect 1307 2616 1653 2624
rect 3307 2616 3533 2624
rect 3787 2616 3973 2624
rect 4067 2616 4153 2624
rect 167 2596 253 2604
rect 267 2596 553 2604
rect 47 2576 133 2584
rect 27 2556 73 2564
rect 87 2556 144 2564
rect 67 2536 113 2544
rect 136 2544 144 2556
rect 256 2556 393 2564
rect 256 2547 264 2556
rect 416 2547 424 2596
rect 567 2596 593 2604
rect 967 2596 1093 2604
rect 1187 2596 1233 2604
rect 1347 2596 1493 2604
rect 1507 2596 1593 2604
rect 1607 2596 1793 2604
rect 2387 2596 2693 2604
rect 3247 2596 3473 2604
rect 3687 2596 3813 2604
rect 3827 2596 3913 2604
rect 4027 2596 4093 2604
rect 527 2576 613 2584
rect 927 2576 953 2584
rect 987 2576 1193 2584
rect 1247 2576 1373 2584
rect 1467 2576 1493 2584
rect 1987 2576 2073 2584
rect 2087 2576 2133 2584
rect 2267 2576 2333 2584
rect 2347 2576 2464 2584
rect 456 2564 464 2573
rect 456 2556 564 2564
rect 136 2536 153 2544
rect 167 2536 233 2544
rect 447 2536 533 2544
rect 327 2516 353 2524
rect 367 2516 373 2524
rect 467 2516 533 2524
rect 556 2524 564 2556
rect 556 2516 613 2524
rect 716 2524 724 2573
rect 847 2556 864 2564
rect 707 2516 724 2524
rect 767 2516 833 2524
rect 856 2524 864 2556
rect 907 2556 964 2564
rect 887 2536 904 2544
rect 856 2516 873 2524
rect 27 2496 573 2504
rect 896 2504 904 2536
rect 956 2527 964 2556
rect 1007 2556 1013 2564
rect 1067 2556 1273 2564
rect 996 2527 1004 2553
rect 1167 2536 1184 2544
rect 1087 2516 1153 2524
rect 1176 2524 1184 2536
rect 1176 2516 1193 2524
rect 896 2496 933 2504
rect 987 2496 1133 2504
rect 1356 2504 1364 2553
rect 1436 2547 1444 2573
rect 1707 2556 1733 2564
rect 2456 2564 2464 2576
rect 2487 2576 2833 2584
rect 2847 2576 2853 2584
rect 2907 2576 3033 2584
rect 3047 2576 3333 2584
rect 3967 2576 3984 2584
rect 2456 2556 2493 2564
rect 2687 2556 2733 2564
rect 2747 2556 2793 2564
rect 2927 2556 3073 2564
rect 3087 2556 3193 2564
rect 1476 2524 1484 2553
rect 1547 2536 1633 2544
rect 1476 2516 1513 2524
rect 1567 2516 1593 2524
rect 1607 2516 1653 2524
rect 1667 2516 1813 2524
rect 1287 2496 1364 2504
rect 1407 2496 1413 2504
rect 1427 2496 1593 2504
rect 1827 2496 1893 2504
rect 1936 2504 1944 2553
rect 2027 2536 2093 2544
rect 2116 2544 2124 2553
rect 2107 2536 2124 2544
rect 2187 2536 2193 2544
rect 2207 2536 2213 2544
rect 2327 2536 2373 2544
rect 2007 2516 2053 2524
rect 2396 2524 2404 2553
rect 2427 2536 2693 2544
rect 2787 2536 2924 2544
rect 2916 2527 2924 2536
rect 2947 2536 3093 2544
rect 3147 2536 3293 2544
rect 3356 2544 3364 2573
rect 3487 2556 3593 2564
rect 3707 2556 3873 2564
rect 3356 2536 3393 2544
rect 3787 2536 3893 2544
rect 3956 2544 3964 2553
rect 3976 2547 3984 2576
rect 4087 2576 4473 2584
rect 4007 2556 4033 2564
rect 4327 2556 4513 2564
rect 4547 2556 4593 2564
rect 3947 2536 3964 2544
rect 4207 2536 4213 2544
rect 4227 2536 4333 2544
rect 4447 2536 4584 2544
rect 4576 2527 4584 2536
rect 4616 2527 4624 2553
rect 2347 2516 2404 2524
rect 2587 2516 2793 2524
rect 2807 2516 2853 2524
rect 3327 2516 3393 2524
rect 3447 2516 3513 2524
rect 3527 2516 4053 2524
rect 4267 2516 4313 2524
rect 4447 2516 4553 2524
rect 4647 2516 4693 2524
rect 1936 2496 2033 2504
rect 2567 2496 2573 2504
rect 2587 2496 2653 2504
rect 2727 2496 2813 2504
rect 2887 2496 2953 2504
rect 3287 2496 3553 2504
rect 3567 2496 3573 2504
rect 3827 2496 4033 2504
rect 4047 2496 4093 2504
rect 4467 2496 4653 2504
rect 487 2476 593 2484
rect 727 2476 813 2484
rect 827 2476 833 2484
rect 967 2476 1013 2484
rect 1367 2476 1413 2484
rect 1427 2476 1673 2484
rect 1807 2476 1853 2484
rect 1967 2476 2033 2484
rect 3867 2476 3933 2484
rect 3967 2476 4233 2484
rect 4507 2476 4613 2484
rect 4627 2476 4693 2484
rect 347 2456 773 2464
rect 927 2456 1113 2464
rect 1827 2456 2093 2464
rect 3267 2456 4073 2464
rect 987 2436 1073 2444
rect 4067 2436 4113 2444
rect 427 2416 493 2424
rect 587 2416 1433 2424
rect 1787 2416 1933 2424
rect 1947 2416 2153 2424
rect 2927 2416 2973 2424
rect 47 2396 213 2404
rect 767 2396 813 2404
rect 827 2396 873 2404
rect 1047 2396 1253 2404
rect 3787 2396 4013 2404
rect 687 2376 993 2384
rect 1007 2376 1153 2384
rect 1507 2376 1633 2384
rect 3827 2376 3993 2384
rect 147 2356 273 2364
rect 327 2356 453 2364
rect 767 2356 1473 2364
rect 2267 2356 2633 2364
rect 3107 2356 3533 2364
rect 3587 2356 3673 2364
rect 3707 2356 3873 2364
rect 76 2336 413 2344
rect 16 2224 24 2313
rect 36 2267 44 2313
rect 76 2284 84 2336
rect 96 2287 104 2313
rect 207 2296 293 2304
rect 316 2287 324 2313
rect 67 2276 84 2284
rect 107 2276 164 2284
rect 87 2256 133 2264
rect 156 2264 164 2276
rect 187 2276 233 2284
rect 287 2276 313 2284
rect 336 2284 344 2336
rect 967 2336 1193 2344
rect 1327 2336 1353 2344
rect 1487 2336 1573 2344
rect 2527 2336 2673 2344
rect 3956 2336 4133 2344
rect 527 2316 633 2324
rect 1127 2316 1133 2324
rect 1147 2316 1313 2324
rect 2287 2316 2613 2324
rect 356 2304 364 2313
rect 356 2296 384 2304
rect 336 2276 353 2284
rect 376 2267 384 2296
rect 667 2296 733 2304
rect 856 2296 913 2304
rect 156 2256 333 2264
rect 436 2264 444 2273
rect 436 2256 464 2264
rect 207 2236 213 2244
rect 227 2236 293 2244
rect 347 2236 433 2244
rect 456 2244 464 2256
rect 536 2264 544 2273
rect 487 2256 544 2264
rect 567 2256 593 2264
rect 456 2236 473 2244
rect 676 2227 684 2273
rect 696 2264 704 2273
rect 856 2267 864 2296
rect 1007 2296 1093 2304
rect 1107 2296 1253 2304
rect 1987 2296 2073 2304
rect 2367 2296 2393 2304
rect 2536 2304 2544 2316
rect 3307 2316 3633 2324
rect 3667 2316 3713 2324
rect 2527 2296 2544 2304
rect 2567 2296 2613 2304
rect 3007 2296 3153 2304
rect 3567 2296 3773 2304
rect 956 2267 964 2293
rect 1047 2276 1173 2284
rect 1567 2276 1613 2284
rect 1927 2276 1973 2284
rect 2027 2276 2213 2284
rect 2267 2276 2324 2284
rect 696 2256 793 2264
rect 927 2256 953 2264
rect 1027 2256 1053 2264
rect 1067 2256 1073 2264
rect 1216 2264 1224 2273
rect 2316 2267 2324 2276
rect 2387 2276 2433 2284
rect 2487 2276 2533 2284
rect 2867 2276 3084 2284
rect 1187 2256 1224 2264
rect 1247 2256 1384 2264
rect 847 2236 953 2244
rect 987 2236 1093 2244
rect 1207 2236 1333 2244
rect 1376 2244 1384 2256
rect 1427 2256 1453 2264
rect 1587 2256 1653 2264
rect 1807 2256 2244 2264
rect 1376 2236 1573 2244
rect 1847 2236 1913 2244
rect 2236 2244 2244 2256
rect 2267 2256 2293 2264
rect 2376 2247 2384 2273
rect 3076 2267 3084 2276
rect 3176 2276 3493 2284
rect 3176 2267 3184 2276
rect 3596 2276 3613 2284
rect 3596 2267 3604 2276
rect 3667 2276 3684 2284
rect 3676 2267 3684 2276
rect 3727 2276 3784 2284
rect 3776 2267 3784 2276
rect 3816 2267 3824 2293
rect 2427 2256 2573 2264
rect 2807 2256 2933 2264
rect 2987 2256 3053 2264
rect 3207 2256 3233 2264
rect 3247 2256 3253 2264
rect 3387 2256 3513 2264
rect 3647 2256 3673 2264
rect 3916 2264 3924 2273
rect 3936 2267 3944 2293
rect 3956 2287 3964 2336
rect 4587 2336 4773 2344
rect 3987 2316 4084 2324
rect 4016 2296 4053 2304
rect 4016 2267 4024 2296
rect 3836 2256 3924 2264
rect 2236 2236 2264 2244
rect 2256 2227 2264 2236
rect 2287 2236 2353 2244
rect 2547 2236 2613 2244
rect 2947 2236 3333 2244
rect 3347 2236 3493 2244
rect 3607 2236 3653 2244
rect 3836 2244 3844 2256
rect 3947 2256 4004 2264
rect 3996 2247 4004 2256
rect 3727 2236 3844 2244
rect 3867 2236 3973 2244
rect 4036 2244 4044 2273
rect 4016 2236 4044 2244
rect 4016 2227 4024 2236
rect 16 2216 213 2224
rect 247 2216 273 2224
rect 407 2216 513 2224
rect 527 2216 573 2224
rect 847 2216 933 2224
rect 987 2216 1133 2224
rect 1167 2216 1253 2224
rect 1547 2216 1673 2224
rect 1887 2216 1953 2224
rect 1967 2216 2113 2224
rect 2176 2216 2193 2224
rect 167 2196 353 2204
rect 367 2196 553 2204
rect 567 2196 653 2204
rect 827 2196 913 2204
rect 1387 2196 1713 2204
rect 1827 2196 1933 2204
rect 2176 2187 2184 2216
rect 2667 2216 3213 2224
rect 3367 2216 3513 2224
rect 4076 2224 4084 2316
rect 4587 2316 4693 2324
rect 4347 2296 4533 2304
rect 4547 2296 4653 2304
rect 4627 2276 4673 2284
rect 4227 2256 4413 2264
rect 4467 2256 4593 2264
rect 4687 2256 4733 2264
rect 4167 2236 4233 2244
rect 4047 2216 4084 2224
rect 2467 2196 2693 2204
rect 2707 2196 2953 2204
rect 3127 2196 3293 2204
rect 3607 2196 3753 2204
rect 3767 2196 3833 2204
rect 27 2176 313 2184
rect 587 2176 713 2184
rect 1647 2176 1693 2184
rect 1787 2176 1993 2184
rect 2907 2176 2973 2184
rect 2987 2176 3013 2184
rect 3027 2176 3133 2184
rect 3147 2176 3173 2184
rect 3587 2176 4553 2184
rect 287 2156 533 2164
rect 547 2156 893 2164
rect 1707 2156 1813 2164
rect 1847 2156 1873 2164
rect 1947 2156 2233 2164
rect 2547 2156 2593 2164
rect 2607 2156 2673 2164
rect 2927 2156 3253 2164
rect 4547 2156 4593 2164
rect 187 2136 753 2144
rect 1327 2136 1753 2144
rect 1767 2136 2053 2144
rect 2167 2136 2293 2144
rect 2667 2136 3273 2144
rect 3687 2136 3793 2144
rect 3827 2136 3933 2144
rect 4307 2136 4373 2144
rect 4427 2136 4533 2144
rect 4547 2136 4633 2144
rect 467 2116 573 2124
rect 647 2116 713 2124
rect 736 2116 793 2124
rect 36 2096 53 2104
rect 36 2044 44 2096
rect 87 2096 324 2104
rect 67 2076 133 2084
rect 156 2076 173 2084
rect 156 2064 164 2076
rect 267 2076 304 2084
rect 96 2056 164 2064
rect 96 2047 104 2056
rect 36 2036 73 2044
rect 216 2044 224 2073
rect 187 2036 224 2044
rect 236 2027 244 2073
rect 296 2067 304 2076
rect 316 2067 324 2096
rect 367 2096 404 2104
rect 367 2076 384 2084
rect 276 2044 284 2053
rect 276 2036 333 2044
rect 376 2044 384 2076
rect 396 2067 404 2096
rect 416 2096 473 2104
rect 416 2067 424 2096
rect 736 2104 744 2116
rect 947 2116 1033 2124
rect 1667 2116 1893 2124
rect 1927 2116 1973 2124
rect 2067 2116 2213 2124
rect 3007 2116 3033 2124
rect 3207 2116 3244 2124
rect 496 2096 744 2104
rect 496 2084 504 2096
rect 807 2096 884 2104
rect 436 2076 504 2084
rect 436 2067 444 2076
rect 776 2084 784 2093
rect 756 2076 784 2084
rect 796 2076 813 2084
rect 536 2056 593 2064
rect 376 2036 393 2044
rect 447 2036 513 2044
rect 256 2004 264 2033
rect 536 2024 544 2056
rect 656 2064 664 2073
rect 656 2056 693 2064
rect 636 2044 644 2053
rect 756 2047 764 2076
rect 567 2036 713 2044
rect 796 2044 804 2076
rect 876 2084 884 2096
rect 907 2096 1013 2104
rect 1127 2096 1213 2104
rect 1236 2096 1413 2104
rect 876 2076 933 2084
rect 1007 2076 1064 2084
rect 827 2056 913 2064
rect 796 2036 873 2044
rect 956 2044 964 2073
rect 1027 2056 1044 2064
rect 936 2036 964 2044
rect 536 2016 564 2024
rect 27 1996 264 2004
rect 276 1996 513 2004
rect 276 1984 284 1996
rect 556 2004 564 2016
rect 647 2016 793 2024
rect 916 2024 924 2033
rect 936 2027 944 2036
rect 907 2016 924 2024
rect 1016 2024 1024 2033
rect 1036 2027 1044 2056
rect 1056 2027 1064 2076
rect 1116 2076 1153 2084
rect 1096 2027 1104 2053
rect 1007 2016 1024 2024
rect 1116 2024 1124 2076
rect 1147 2056 1193 2064
rect 1236 2064 1244 2096
rect 1867 2096 1933 2104
rect 2287 2096 2393 2104
rect 2407 2096 2573 2104
rect 3067 2096 3213 2104
rect 1267 2076 1293 2084
rect 1347 2076 1373 2084
rect 1567 2076 1693 2084
rect 1736 2067 1744 2093
rect 1756 2067 1764 2093
rect 1956 2084 1964 2093
rect 1936 2076 1964 2084
rect 1227 2056 1244 2064
rect 1287 2056 1313 2064
rect 1507 2056 1633 2064
rect 1687 2056 1713 2064
rect 1167 2036 1433 2044
rect 1447 2036 1533 2044
rect 1116 2016 1293 2024
rect 1407 2016 1733 2024
rect 1747 2016 1893 2024
rect 1916 2024 1924 2073
rect 1936 2047 1944 2076
rect 2047 2076 2113 2084
rect 2567 2076 2673 2084
rect 2927 2076 3093 2084
rect 3156 2076 3173 2084
rect 3156 2067 3164 2076
rect 3236 2084 3244 2116
rect 3547 2116 4313 2124
rect 4327 2116 4473 2124
rect 3627 2096 3813 2104
rect 3847 2096 4053 2104
rect 4067 2096 4193 2104
rect 4367 2096 4413 2104
rect 3196 2076 3244 2084
rect 1967 2056 2093 2064
rect 2347 2056 2413 2064
rect 2727 2056 2764 2064
rect 2756 2047 2764 2056
rect 2787 2056 3133 2064
rect 3196 2064 3204 2076
rect 3327 2076 3453 2084
rect 3547 2076 3573 2084
rect 3667 2076 3793 2084
rect 3887 2076 3973 2084
rect 3987 2076 4033 2084
rect 4336 2084 4344 2093
rect 4316 2076 4344 2084
rect 3176 2056 3204 2064
rect 2687 2036 2733 2044
rect 2807 2036 2913 2044
rect 3176 2044 3184 2056
rect 3267 2056 3293 2064
rect 3616 2064 3624 2073
rect 3347 2056 3624 2064
rect 4096 2064 4104 2073
rect 4316 2067 4324 2076
rect 4496 2067 4504 2093
rect 4527 2076 4553 2084
rect 3927 2056 4104 2064
rect 4347 2056 4373 2064
rect 3127 2036 3184 2044
rect 3387 2036 4333 2044
rect 1916 2016 1993 2024
rect 3447 2016 3493 2024
rect 3807 2016 3813 2024
rect 3827 2016 4053 2024
rect 556 1996 733 2004
rect 787 1996 853 2004
rect 987 1996 1073 2004
rect 1127 1996 1173 2004
rect 1527 1996 1573 2004
rect 1887 1996 2013 2004
rect 2627 1996 2693 2004
rect 2707 1996 2753 2004
rect 3147 1996 3633 2004
rect 187 1976 284 1984
rect 667 1976 893 1984
rect 907 1976 993 1984
rect 1367 1976 1653 1984
rect 1927 1976 2233 1984
rect 2387 1976 2653 1984
rect 227 1956 693 1964
rect 707 1956 853 1964
rect 2527 1956 2673 1964
rect 4007 1956 4073 1964
rect 247 1936 293 1944
rect 2087 1936 2093 1944
rect 2107 1936 2153 1944
rect 2167 1936 2393 1944
rect 2827 1936 3273 1944
rect 3627 1936 3713 1944
rect 3907 1936 4013 1944
rect 4167 1936 4193 1944
rect 247 1916 553 1924
rect 687 1916 773 1924
rect 1407 1916 1453 1924
rect 4207 1916 4233 1924
rect 327 1896 613 1904
rect 727 1896 1013 1904
rect 1727 1896 1753 1904
rect 27 1876 93 1884
rect 407 1876 833 1884
rect 847 1876 893 1884
rect 967 1876 1433 1884
rect 47 1856 213 1864
rect 307 1856 373 1864
rect 387 1856 453 1864
rect 587 1856 813 1864
rect 887 1856 953 1864
rect 1047 1856 1153 1864
rect 2207 1856 2393 1864
rect 2407 1856 2933 1864
rect 2947 1856 3153 1864
rect 3167 1856 3553 1864
rect 3667 1856 4113 1864
rect 127 1836 233 1844
rect 316 1836 413 1844
rect 56 1764 64 1833
rect 107 1816 213 1824
rect 316 1824 324 1836
rect 487 1836 713 1844
rect 867 1836 984 1844
rect 227 1816 324 1824
rect 387 1816 433 1824
rect 447 1816 573 1824
rect 587 1816 673 1824
rect 747 1816 804 1824
rect 76 1787 84 1813
rect 167 1796 184 1804
rect 176 1784 184 1796
rect 207 1796 253 1804
rect 336 1787 344 1813
rect 796 1807 804 1816
rect 827 1816 864 1824
rect 687 1796 724 1804
rect 176 1776 273 1784
rect 387 1776 453 1784
rect 507 1776 533 1784
rect 627 1776 693 1784
rect 716 1784 724 1796
rect 716 1776 733 1784
rect 56 1756 93 1764
rect 267 1756 353 1764
rect 376 1756 533 1764
rect 47 1736 173 1744
rect 376 1744 384 1756
rect 547 1756 593 1764
rect 796 1764 804 1793
rect 856 1787 864 1816
rect 827 1776 844 1784
rect 647 1756 784 1764
rect 796 1756 813 1764
rect 227 1736 384 1744
rect 427 1736 513 1744
rect 596 1736 653 1744
rect 27 1716 133 1724
rect 327 1716 393 1724
rect 596 1724 604 1736
rect 667 1736 753 1744
rect 776 1744 784 1756
rect 836 1764 844 1776
rect 867 1776 873 1784
rect 836 1756 853 1764
rect 916 1764 924 1813
rect 976 1807 984 1836
rect 996 1836 1013 1844
rect 996 1827 1004 1836
rect 1047 1836 1084 1844
rect 1076 1824 1084 1836
rect 1107 1836 1233 1844
rect 1076 1816 1093 1824
rect 1036 1787 1044 1813
rect 947 1776 1013 1784
rect 887 1756 924 1764
rect 1056 1764 1064 1813
rect 1136 1787 1144 1836
rect 1307 1836 1713 1844
rect 2167 1836 2273 1844
rect 2367 1836 2473 1844
rect 2716 1836 2733 1844
rect 1167 1816 1253 1824
rect 1276 1784 1284 1833
rect 1307 1816 1404 1824
rect 1396 1804 1404 1816
rect 1447 1816 1533 1824
rect 1627 1816 1673 1824
rect 1807 1816 1933 1824
rect 2087 1816 2193 1824
rect 2347 1816 2384 1824
rect 2376 1807 2384 1816
rect 1396 1796 1424 1804
rect 1416 1787 1424 1796
rect 1487 1796 1533 1804
rect 1567 1796 1633 1804
rect 1727 1796 1793 1804
rect 2187 1796 2253 1804
rect 2287 1796 2333 1804
rect 1276 1776 1293 1784
rect 1427 1776 1513 1784
rect 1747 1776 1813 1784
rect 1827 1776 1853 1784
rect 2147 1776 2193 1784
rect 2336 1784 2344 1793
rect 2336 1776 2493 1784
rect 2596 1784 2604 1793
rect 2547 1776 2604 1784
rect 2636 1784 2644 1793
rect 2636 1776 2693 1784
rect 1056 1756 1073 1764
rect 1087 1756 1233 1764
rect 1507 1756 1633 1764
rect 1787 1756 1833 1764
rect 2227 1756 2413 1764
rect 2507 1756 2573 1764
rect 2716 1764 2724 1836
rect 3307 1836 3333 1844
rect 3347 1836 3453 1844
rect 3467 1836 3813 1844
rect 3827 1836 4273 1844
rect 4527 1836 4553 1844
rect 2747 1816 2804 1824
rect 2796 1804 2804 1816
rect 3067 1816 3133 1824
rect 3427 1816 3513 1824
rect 3967 1816 3984 1824
rect 2796 1796 2853 1804
rect 2796 1784 2804 1796
rect 2907 1796 2953 1804
rect 3387 1796 3433 1804
rect 3867 1796 3913 1804
rect 3976 1804 3984 1816
rect 4667 1816 4733 1824
rect 3976 1796 4064 1804
rect 2787 1776 2804 1784
rect 2887 1776 2913 1784
rect 3067 1776 3073 1784
rect 3087 1776 3093 1784
rect 3336 1784 3344 1793
rect 3336 1776 3373 1784
rect 3787 1776 3813 1784
rect 3956 1784 3964 1793
rect 3887 1776 3964 1784
rect 3987 1776 4033 1784
rect 4056 1767 4064 1796
rect 4116 1796 4213 1804
rect 4116 1787 4124 1796
rect 4307 1796 4353 1804
rect 4396 1796 4453 1804
rect 2716 1756 2793 1764
rect 2827 1756 2833 1764
rect 2847 1756 3033 1764
rect 3467 1756 3493 1764
rect 3587 1756 3733 1764
rect 3767 1756 3813 1764
rect 3827 1756 4033 1764
rect 4256 1764 4264 1793
rect 4396 1784 4404 1796
rect 4347 1776 4404 1784
rect 4427 1776 4493 1784
rect 4587 1776 4673 1784
rect 4247 1756 4393 1764
rect 776 1736 913 1744
rect 967 1736 1013 1744
rect 1047 1736 1173 1744
rect 1187 1736 1273 1744
rect 1467 1736 1653 1744
rect 2367 1736 2413 1744
rect 2467 1736 2513 1744
rect 3367 1736 3633 1744
rect 3887 1736 3993 1744
rect 4087 1736 4233 1744
rect 4407 1736 4593 1744
rect 476 1716 604 1724
rect 127 1696 253 1704
rect 287 1696 453 1704
rect 476 1704 484 1716
rect 667 1716 813 1724
rect 867 1716 1253 1724
rect 1387 1716 1833 1724
rect 1847 1716 2293 1724
rect 3487 1716 3573 1724
rect 3807 1716 3953 1724
rect 4027 1716 4453 1724
rect 4467 1716 4653 1724
rect 467 1696 484 1704
rect 767 1696 933 1704
rect 1287 1696 1313 1704
rect 1327 1696 1693 1704
rect 3147 1696 3253 1704
rect 3867 1696 4073 1704
rect 4087 1696 4093 1704
rect 4227 1696 4273 1704
rect 4347 1696 4473 1704
rect 147 1676 973 1684
rect 1267 1676 1293 1684
rect 1336 1676 1613 1684
rect 367 1656 633 1664
rect 1336 1664 1344 1676
rect 2487 1676 2553 1684
rect 2787 1676 2833 1684
rect 3627 1676 3793 1684
rect 3907 1676 4293 1684
rect 4427 1676 4653 1684
rect 1147 1656 1344 1664
rect 1367 1656 1853 1664
rect 2567 1656 3333 1664
rect 3847 1656 3893 1664
rect 4067 1656 4093 1664
rect 4127 1656 4153 1664
rect 4167 1656 4273 1664
rect 4327 1656 4413 1664
rect 4447 1656 4533 1664
rect 287 1636 413 1644
rect 507 1636 573 1644
rect 587 1636 593 1644
rect 727 1636 773 1644
rect 927 1636 993 1644
rect 1127 1636 1473 1644
rect 1487 1636 1533 1644
rect 1547 1636 1573 1644
rect 1967 1636 2033 1644
rect 2167 1636 2353 1644
rect 2447 1636 2613 1644
rect 2627 1636 2673 1644
rect 2687 1636 2713 1644
rect 2767 1636 2933 1644
rect 107 1616 124 1624
rect 27 1596 93 1604
rect 116 1604 124 1616
rect 147 1616 173 1624
rect 307 1616 473 1624
rect 496 1616 533 1624
rect 116 1596 144 1604
rect 136 1587 144 1596
rect 387 1596 424 1604
rect 416 1587 424 1596
rect 496 1604 504 1616
rect 647 1616 713 1624
rect 827 1616 913 1624
rect 967 1616 1164 1624
rect 476 1596 504 1604
rect 596 1596 653 1604
rect 47 1576 113 1584
rect 167 1576 213 1584
rect 227 1576 293 1584
rect 307 1576 373 1584
rect 436 1567 444 1593
rect 476 1584 484 1596
rect 456 1576 484 1584
rect 127 1556 193 1564
rect 456 1544 464 1576
rect 596 1584 604 1596
rect 776 1596 793 1604
rect 587 1576 604 1584
rect 627 1576 693 1584
rect 776 1584 784 1596
rect 887 1596 904 1604
rect 727 1576 784 1584
rect 807 1576 813 1584
rect 847 1576 873 1584
rect 896 1584 904 1596
rect 1027 1596 1044 1604
rect 896 1576 913 1584
rect 947 1576 1013 1584
rect 796 1564 804 1573
rect 707 1556 804 1564
rect 867 1556 884 1564
rect 327 1536 464 1544
rect 616 1544 624 1553
rect 547 1536 624 1544
rect 816 1544 824 1553
rect 876 1544 884 1556
rect 907 1556 1013 1564
rect 1036 1547 1044 1596
rect 1156 1587 1164 1616
rect 1347 1616 1373 1624
rect 1547 1616 1593 1624
rect 1687 1616 1784 1624
rect 1187 1596 1193 1604
rect 1316 1604 1324 1613
rect 1207 1596 1264 1604
rect 1316 1596 1444 1604
rect 1076 1576 1113 1584
rect 1076 1564 1084 1576
rect 1196 1576 1213 1584
rect 1067 1556 1084 1564
rect 1107 1556 1153 1564
rect 1196 1564 1204 1576
rect 1256 1584 1264 1596
rect 1256 1576 1333 1584
rect 1347 1576 1413 1584
rect 1187 1556 1204 1564
rect 667 1536 864 1544
rect 876 1536 993 1544
rect 567 1516 733 1524
rect 856 1524 864 1536
rect 1216 1544 1224 1553
rect 1236 1547 1244 1573
rect 1287 1556 1333 1564
rect 1436 1564 1444 1596
rect 1627 1596 1753 1604
rect 1507 1576 1553 1584
rect 1587 1576 1673 1584
rect 1776 1584 1784 1616
rect 1756 1576 1784 1584
rect 1796 1616 1833 1624
rect 1427 1556 1444 1564
rect 1527 1556 1633 1564
rect 1207 1536 1224 1544
rect 1696 1544 1704 1573
rect 1756 1567 1764 1576
rect 1796 1567 1804 1616
rect 2027 1616 2153 1624
rect 2187 1616 2433 1624
rect 2607 1616 2733 1624
rect 1847 1596 1873 1604
rect 1816 1564 1824 1593
rect 1916 1587 1924 1613
rect 1936 1584 1944 1613
rect 2027 1596 2093 1604
rect 2207 1596 2533 1604
rect 2236 1587 2244 1596
rect 2576 1596 2633 1604
rect 2576 1587 2584 1596
rect 2707 1596 2753 1604
rect 1936 1576 1953 1584
rect 2067 1576 2113 1584
rect 2816 1584 2824 1636
rect 3147 1636 3213 1644
rect 3327 1636 3513 1644
rect 3667 1636 3744 1644
rect 2847 1616 2933 1624
rect 3007 1616 3353 1624
rect 3407 1616 3533 1624
rect 2836 1587 2844 1613
rect 2867 1596 2893 1604
rect 2927 1596 2944 1604
rect 2807 1576 2824 1584
rect 2936 1584 2944 1596
rect 2967 1596 3064 1604
rect 3056 1587 3064 1596
rect 3107 1596 3173 1604
rect 3347 1596 3384 1604
rect 2887 1576 2993 1584
rect 3067 1576 3113 1584
rect 3167 1576 3213 1584
rect 1816 1556 1833 1564
rect 1907 1556 1973 1564
rect 2007 1556 2033 1564
rect 2107 1556 2173 1564
rect 2187 1556 2333 1564
rect 2536 1564 2544 1573
rect 3236 1567 3244 1593
rect 3376 1587 3384 1596
rect 3447 1596 3473 1604
rect 3576 1567 3584 1613
rect 3736 1604 3744 1636
rect 3787 1636 4624 1644
rect 3767 1616 3864 1624
rect 3736 1596 3784 1604
rect 3776 1567 3784 1596
rect 3816 1596 3833 1604
rect 3816 1584 3824 1596
rect 3807 1576 3824 1584
rect 3856 1584 3864 1616
rect 3876 1587 3884 1636
rect 3947 1616 4073 1624
rect 3996 1607 4004 1616
rect 4267 1616 4333 1624
rect 4527 1616 4573 1624
rect 4096 1604 4104 1613
rect 4076 1596 4104 1604
rect 4176 1604 4184 1613
rect 4356 1604 4364 1613
rect 4176 1596 4244 1604
rect 3847 1576 3864 1584
rect 4076 1584 4084 1596
rect 4027 1576 4084 1584
rect 4107 1576 4213 1584
rect 4236 1584 4244 1596
rect 4336 1596 4364 1604
rect 4236 1576 4253 1584
rect 2347 1556 2553 1564
rect 2627 1556 2653 1564
rect 2787 1556 2893 1564
rect 3347 1556 3413 1564
rect 3827 1556 4313 1564
rect 4336 1564 4344 1596
rect 4387 1596 4513 1604
rect 4367 1576 4433 1584
rect 4596 1584 4604 1593
rect 4616 1587 4624 1636
rect 4647 1596 4673 1604
rect 4727 1596 4753 1604
rect 4787 1596 4804 1604
rect 4507 1576 4604 1584
rect 4727 1576 4773 1584
rect 4336 1556 4353 1564
rect 4467 1556 4473 1564
rect 4487 1556 4693 1564
rect 4796 1564 4804 1596
rect 4747 1556 4804 1564
rect 1267 1536 1704 1544
rect 1787 1536 1853 1544
rect 2127 1536 2373 1544
rect 2807 1536 2913 1544
rect 3187 1536 3193 1544
rect 3207 1536 3333 1544
rect 3487 1536 3713 1544
rect 4067 1536 4133 1544
rect 4207 1536 4253 1544
rect 856 1516 893 1524
rect 1307 1516 1613 1524
rect 3307 1516 3353 1524
rect 4387 1516 4633 1524
rect 487 1496 693 1504
rect 807 1496 913 1504
rect 1007 1496 1233 1504
rect 1247 1496 1313 1504
rect 1447 1496 1453 1504
rect 1467 1496 1593 1504
rect 2507 1496 3413 1504
rect 3427 1496 3453 1504
rect 3627 1496 4213 1504
rect 847 1476 1193 1484
rect 1207 1476 1413 1484
rect 1507 1476 1693 1484
rect 1707 1476 1793 1484
rect 207 1456 453 1464
rect 747 1456 853 1464
rect 887 1456 1553 1464
rect 3607 1456 3653 1464
rect 307 1436 373 1444
rect 387 1436 1033 1444
rect 1187 1436 1513 1444
rect 367 1416 413 1424
rect 827 1416 933 1424
rect 1447 1416 1533 1424
rect 4267 1416 4293 1424
rect 67 1396 73 1404
rect 87 1396 353 1404
rect 367 1396 433 1404
rect 1267 1396 1393 1404
rect 1407 1396 1413 1404
rect 1427 1396 1553 1404
rect 1747 1396 1833 1404
rect 1847 1396 1853 1404
rect 4187 1396 4293 1404
rect 107 1376 133 1384
rect 336 1376 393 1384
rect 236 1347 244 1373
rect 287 1356 324 1364
rect 67 1336 124 1344
rect 116 1327 124 1336
rect 187 1336 224 1344
rect 216 1324 224 1336
rect 256 1344 264 1353
rect 256 1336 284 1344
rect 216 1316 253 1324
rect 96 1304 104 1313
rect 96 1296 153 1304
rect 276 1304 284 1336
rect 316 1324 324 1356
rect 336 1347 344 1376
rect 407 1376 713 1384
rect 967 1376 1193 1384
rect 1487 1376 1524 1384
rect 776 1356 833 1364
rect 356 1327 364 1353
rect 376 1336 393 1344
rect 316 1316 344 1324
rect 336 1307 344 1316
rect 376 1307 384 1336
rect 427 1336 504 1344
rect 496 1327 504 1336
rect 696 1336 733 1344
rect 627 1316 644 1324
rect 187 1296 284 1304
rect 87 1276 133 1284
rect 147 1276 313 1284
rect 416 1284 424 1313
rect 496 1304 504 1313
rect 367 1276 424 1284
rect 476 1296 504 1304
rect 476 1264 484 1296
rect 516 1284 524 1313
rect 536 1304 544 1313
rect 636 1304 644 1316
rect 696 1324 704 1336
rect 667 1316 704 1324
rect 716 1304 724 1313
rect 536 1296 624 1304
rect 636 1296 724 1304
rect 616 1287 624 1296
rect 716 1287 724 1296
rect 776 1304 784 1356
rect 907 1356 973 1364
rect 1107 1356 1204 1364
rect 1027 1336 1033 1344
rect 1047 1336 1073 1344
rect 1127 1336 1173 1344
rect 1196 1344 1204 1356
rect 1227 1356 1373 1364
rect 1407 1356 1493 1364
rect 1516 1364 1524 1376
rect 1947 1376 2053 1384
rect 2067 1376 2093 1384
rect 3267 1376 3293 1384
rect 4187 1376 4393 1384
rect 1516 1356 1544 1364
rect 1196 1336 1224 1344
rect 796 1307 804 1333
rect 836 1307 844 1333
rect 916 1307 924 1333
rect 976 1324 984 1333
rect 947 1316 1093 1324
rect 1127 1316 1193 1324
rect 747 1296 784 1304
rect 1107 1296 1153 1304
rect 507 1276 524 1284
rect 567 1276 593 1284
rect 767 1276 813 1284
rect 867 1276 913 1284
rect 1216 1284 1224 1336
rect 1287 1336 1364 1344
rect 1276 1316 1333 1324
rect 1276 1304 1284 1316
rect 1356 1324 1364 1336
rect 1476 1336 1513 1344
rect 1356 1316 1433 1324
rect 1456 1307 1464 1333
rect 1267 1296 1284 1304
rect 1307 1296 1344 1304
rect 1007 1276 1224 1284
rect 1236 1276 1313 1284
rect 67 1256 484 1264
rect 607 1256 693 1264
rect 1007 1256 1053 1264
rect 1236 1264 1244 1276
rect 1336 1284 1344 1296
rect 1476 1284 1484 1336
rect 1536 1327 1544 1356
rect 1687 1356 1913 1364
rect 1927 1356 2184 1364
rect 1596 1336 1753 1344
rect 1596 1307 1604 1336
rect 1947 1336 1993 1344
rect 2007 1336 2024 1344
rect 1787 1316 1804 1324
rect 1616 1304 1624 1313
rect 1616 1296 1693 1304
rect 1796 1304 1804 1316
rect 1827 1316 1913 1324
rect 2016 1324 2024 1336
rect 2176 1327 2184 1356
rect 2456 1356 2653 1364
rect 2207 1336 2273 1344
rect 2367 1336 2433 1344
rect 2456 1344 2464 1356
rect 2987 1356 3173 1364
rect 3187 1356 3253 1364
rect 4147 1356 4213 1364
rect 4227 1356 4473 1364
rect 4647 1356 4673 1364
rect 4707 1356 4773 1364
rect 2447 1336 2464 1344
rect 2487 1336 2593 1344
rect 2727 1336 2813 1344
rect 3107 1336 3213 1344
rect 3747 1336 3853 1344
rect 3887 1336 3953 1344
rect 3967 1336 4733 1344
rect 2016 1316 2033 1324
rect 2047 1316 2153 1324
rect 1796 1296 1873 1304
rect 1996 1304 2004 1313
rect 1947 1296 2004 1304
rect 2196 1304 2204 1333
rect 2527 1316 2773 1324
rect 2827 1316 2993 1324
rect 3016 1316 3533 1324
rect 2167 1296 2204 1304
rect 2267 1296 2333 1304
rect 2607 1296 2633 1304
rect 2687 1296 2753 1304
rect 3016 1304 3024 1316
rect 3547 1316 3604 1324
rect 3596 1307 3604 1316
rect 3696 1316 3753 1324
rect 2847 1296 3024 1304
rect 3067 1296 3073 1304
rect 3087 1296 3113 1304
rect 1336 1276 1484 1284
rect 1507 1276 1653 1284
rect 1667 1276 1713 1284
rect 1807 1276 1893 1284
rect 1987 1276 2073 1284
rect 2087 1276 2133 1284
rect 2467 1276 2493 1284
rect 2987 1276 3393 1284
rect 3476 1284 3484 1293
rect 3616 1287 3624 1313
rect 3696 1304 3704 1316
rect 3767 1316 4053 1324
rect 4107 1316 4153 1324
rect 4347 1316 4393 1324
rect 4496 1316 4533 1324
rect 3647 1296 3704 1304
rect 3727 1296 3813 1304
rect 3947 1296 4073 1304
rect 4387 1296 4413 1304
rect 3476 1276 3553 1284
rect 3567 1276 3593 1284
rect 3647 1276 3673 1284
rect 3707 1276 3793 1284
rect 4436 1284 4444 1313
rect 4496 1307 4504 1316
rect 4727 1316 4753 1324
rect 4787 1316 4824 1324
rect 4676 1304 4684 1313
rect 4567 1296 4684 1304
rect 4436 1276 4513 1284
rect 4587 1276 4653 1284
rect 1067 1256 1244 1264
rect 1267 1256 1333 1264
rect 1387 1256 1533 1264
rect 1567 1256 1693 1264
rect 1847 1256 1933 1264
rect 1967 1256 2093 1264
rect 2947 1256 3193 1264
rect 3247 1256 3873 1264
rect 4467 1256 4593 1264
rect 447 1236 573 1244
rect 647 1236 853 1244
rect 887 1236 1193 1244
rect 1587 1236 2013 1244
rect 2147 1236 2213 1244
rect 2807 1236 3353 1244
rect 3407 1236 3613 1244
rect 3956 1236 4033 1244
rect 287 1216 453 1224
rect 467 1216 513 1224
rect 587 1216 713 1224
rect 807 1216 853 1224
rect 907 1216 1024 1224
rect 307 1196 553 1204
rect 627 1196 713 1204
rect 807 1196 993 1204
rect 1016 1204 1024 1216
rect 1207 1216 1393 1224
rect 1867 1216 2013 1224
rect 3956 1224 3964 1236
rect 3467 1216 3964 1224
rect 1016 1196 1053 1204
rect 1147 1196 1353 1204
rect 1627 1196 1773 1204
rect 2707 1196 3273 1204
rect 3287 1196 3373 1204
rect 3947 1196 4013 1204
rect -4 1176 213 1184
rect -4 1124 4 1176
rect 307 1176 333 1184
rect 387 1176 593 1184
rect 627 1176 653 1184
rect 747 1176 1033 1184
rect 1187 1176 1213 1184
rect 1587 1176 1633 1184
rect 2647 1176 2853 1184
rect 3387 1176 4273 1184
rect 167 1156 373 1164
rect 407 1156 413 1164
rect 427 1156 653 1164
rect 847 1156 893 1164
rect 987 1156 1093 1164
rect 1147 1156 1193 1164
rect 1527 1156 1693 1164
rect 2687 1156 2873 1164
rect 2907 1156 2973 1164
rect 3147 1156 3473 1164
rect 4447 1156 4573 1164
rect 27 1136 93 1144
rect 107 1136 113 1144
rect 156 1136 204 1144
rect -4 1116 13 1124
rect 47 1116 84 1124
rect 76 1107 84 1116
rect 87 1096 133 1104
rect 36 1084 44 1093
rect 36 1076 93 1084
rect 156 1084 164 1136
rect 107 1076 164 1084
rect 176 1067 184 1113
rect 196 1104 204 1136
rect 247 1136 333 1144
rect 447 1136 533 1144
rect 567 1136 584 1144
rect 227 1116 253 1124
rect 267 1116 293 1124
rect 356 1124 364 1133
rect 356 1116 373 1124
rect 427 1116 564 1124
rect 556 1107 564 1116
rect 196 1096 253 1104
rect 376 1096 433 1104
rect 376 1084 384 1096
rect 467 1096 513 1104
rect 287 1076 384 1084
rect 456 1084 464 1093
rect 576 1087 584 1136
rect 847 1136 1033 1144
rect 1056 1136 1113 1144
rect 856 1116 933 1124
rect 736 1087 744 1113
rect 776 1087 784 1113
rect 407 1076 464 1084
rect 487 1076 533 1084
rect 687 1076 733 1084
rect 207 1056 253 1064
rect 267 1056 353 1064
rect 507 1056 533 1064
rect 816 1064 824 1113
rect 856 1107 864 1116
rect 1056 1107 1064 1136
rect 1127 1136 1233 1144
rect 1307 1136 1353 1144
rect 1367 1136 1613 1144
rect 1647 1136 1673 1144
rect 1707 1136 1793 1144
rect 1867 1136 2053 1144
rect 2227 1136 2353 1144
rect 2627 1136 2693 1144
rect 3007 1136 3173 1144
rect 3187 1136 3213 1144
rect 3227 1136 3333 1144
rect 3827 1136 3853 1144
rect 3907 1136 4133 1144
rect 4187 1136 4393 1144
rect 4567 1136 4753 1144
rect 1127 1116 1293 1124
rect 1216 1087 1224 1116
rect 1447 1116 1473 1124
rect 1487 1116 1553 1124
rect 1687 1116 1753 1124
rect 1767 1116 1873 1124
rect 1936 1116 2133 1124
rect 1247 1096 1364 1104
rect 1356 1087 1364 1096
rect 1376 1087 1384 1113
rect 1416 1104 1424 1113
rect 1416 1096 1493 1104
rect 1567 1096 1624 1104
rect 1616 1087 1624 1096
rect 1827 1096 1893 1104
rect 1936 1104 1944 1116
rect 2407 1116 2593 1124
rect 2656 1116 2733 1124
rect 2656 1107 2664 1116
rect 2747 1116 2793 1124
rect 2987 1116 3013 1124
rect 3267 1116 3573 1124
rect 3587 1116 3593 1124
rect 3607 1116 3873 1124
rect 3927 1116 4013 1124
rect 4027 1116 4293 1124
rect 4307 1116 4333 1124
rect 4347 1116 4353 1124
rect 4376 1116 4444 1124
rect 4376 1107 4384 1116
rect 1916 1096 1944 1104
rect 967 1076 1153 1084
rect 1427 1076 1453 1084
rect 1467 1076 1473 1084
rect 1716 1084 1724 1093
rect 1916 1087 1924 1096
rect 2127 1096 2153 1104
rect 2207 1096 2373 1104
rect 2387 1096 2453 1104
rect 2547 1096 2613 1104
rect 3047 1096 3113 1104
rect 3427 1096 3493 1104
rect 3507 1096 3693 1104
rect 3847 1096 3853 1104
rect 3867 1096 3893 1104
rect 3987 1096 4033 1104
rect 4307 1096 4364 1104
rect 1667 1076 1724 1084
rect 1747 1076 1873 1084
rect 2087 1076 2173 1084
rect 2187 1076 2273 1084
rect 2287 1076 2513 1084
rect 2567 1076 2653 1084
rect 4067 1076 4193 1084
rect 4207 1076 4273 1084
rect 4356 1084 4364 1096
rect 4436 1104 4444 1116
rect 4507 1116 4564 1124
rect 4556 1107 4564 1116
rect 4647 1116 4673 1124
rect 4707 1116 4733 1124
rect 4436 1096 4493 1104
rect 4576 1096 4593 1104
rect 4416 1084 4424 1093
rect 4356 1076 4424 1084
rect 4447 1076 4473 1084
rect 4576 1084 4584 1096
rect 4567 1076 4584 1084
rect 4667 1076 4684 1084
rect 4676 1067 4684 1076
rect 816 1056 873 1064
rect 907 1056 1313 1064
rect 1327 1056 1393 1064
rect 1627 1056 1793 1064
rect 1847 1056 1933 1064
rect 2047 1056 2253 1064
rect 2267 1056 2313 1064
rect 2927 1056 2993 1064
rect 567 1036 1573 1044
rect 1587 1036 1753 1044
rect 1827 1036 1953 1044
rect 4527 1036 4693 1044
rect 647 1016 773 1024
rect 787 1016 813 1024
rect 1307 1016 1624 1024
rect 787 996 1533 1004
rect 1616 1004 1624 1016
rect 1647 1016 1893 1024
rect 1907 1016 2013 1024
rect 1616 996 1653 1004
rect 847 976 893 984
rect 1167 976 1433 984
rect 1507 976 1753 984
rect 1807 976 2513 984
rect 3667 976 3913 984
rect 3927 976 3953 984
rect 1007 956 1073 964
rect 1187 956 1253 964
rect 1267 956 1813 964
rect 2507 956 2553 964
rect 27 936 893 944
rect 1087 936 1193 944
rect 1547 936 1653 944
rect 1787 936 2153 944
rect 527 916 753 924
rect 767 916 813 924
rect 1027 916 1113 924
rect 1207 916 1313 924
rect 1367 916 1433 924
rect 1496 916 1604 924
rect 507 896 573 904
rect 867 896 913 904
rect 927 896 1213 904
rect 1407 896 1453 904
rect 1496 904 1504 916
rect 1467 896 1504 904
rect 1596 904 1604 916
rect 1627 916 1833 924
rect 4507 916 4613 924
rect 4667 916 4753 924
rect 1596 896 1633 904
rect 1667 896 1933 904
rect 4567 896 4753 904
rect 87 876 293 884
rect 427 876 693 884
rect 1056 876 1073 884
rect 1056 867 1064 876
rect 1227 876 1273 884
rect 1387 876 1553 884
rect 1536 867 1544 876
rect 1607 876 1733 884
rect 1747 876 1833 884
rect 1947 876 1993 884
rect 2007 876 2413 884
rect 4627 876 4733 884
rect 236 856 253 864
rect 236 827 244 856
rect 276 856 364 864
rect 276 844 284 856
rect 267 836 284 844
rect 127 816 133 824
rect 147 816 193 824
rect 27 796 153 804
rect 336 804 344 833
rect 356 827 364 856
rect 387 856 453 864
rect 587 856 653 864
rect 707 856 733 864
rect 847 856 864 864
rect 396 836 493 844
rect 396 827 404 836
rect 607 836 644 844
rect 636 807 644 836
rect 707 836 844 844
rect 836 827 844 836
rect 856 827 864 856
rect 907 856 944 864
rect 936 844 944 856
rect 967 856 973 864
rect 987 856 1013 864
rect 1127 856 1333 864
rect 1347 856 1373 864
rect 1396 856 1473 864
rect 936 836 1053 844
rect 1096 827 1104 853
rect 1207 836 1253 844
rect 1396 844 1404 856
rect 1587 856 1753 864
rect 1767 856 1873 864
rect 1987 856 2353 864
rect 2367 856 2444 864
rect 2436 847 2444 856
rect 2507 856 2544 864
rect 1347 836 1404 844
rect 1427 836 1553 844
rect 1567 836 1673 844
rect 1756 836 2053 844
rect 696 816 753 824
rect 167 796 433 804
rect 447 796 493 804
rect 696 804 704 816
rect 907 816 973 824
rect 1296 824 1304 833
rect 1756 827 1764 836
rect 2147 836 2193 844
rect 2327 836 2393 844
rect 2536 844 2544 856
rect 2567 856 2753 864
rect 2807 856 2893 864
rect 2907 856 2933 864
rect 3367 856 3393 864
rect 3647 856 3713 864
rect 3947 856 4013 864
rect 2536 836 2573 844
rect 2607 836 2633 844
rect 2787 836 2853 844
rect 3087 836 3233 844
rect 1296 816 1553 824
rect 1607 816 1713 824
rect 1787 816 1813 824
rect 1896 816 2173 824
rect 687 796 704 804
rect 727 796 933 804
rect 1107 796 1353 804
rect 1727 796 1793 804
rect 1896 804 1904 816
rect 2227 816 2273 824
rect 2676 824 2684 833
rect 2627 816 2684 824
rect 2707 816 2833 824
rect 2956 824 2964 833
rect 2927 816 3044 824
rect 1836 796 1904 804
rect 187 776 293 784
rect 707 776 873 784
rect 1087 776 1293 784
rect 1307 776 1493 784
rect 1836 784 1844 796
rect 1927 796 1953 804
rect 2027 796 2173 804
rect 2247 796 2293 804
rect 2587 796 2653 804
rect 2987 796 3013 804
rect 3036 804 3044 816
rect 3067 816 3164 824
rect 3156 807 3164 816
rect 3316 824 3324 853
rect 3347 836 3373 844
rect 4036 844 4044 853
rect 3987 836 4044 844
rect 3267 816 3324 824
rect 3487 816 3533 824
rect 3607 816 3633 824
rect 3807 816 3993 824
rect 4087 816 4253 824
rect 4267 816 4313 824
rect 4467 816 4633 824
rect 3036 796 3093 804
rect 3416 804 3424 813
rect 4676 807 4684 853
rect 3167 796 3424 804
rect 3507 796 3713 804
rect 3867 796 4113 804
rect 4127 796 4153 804
rect 4167 796 4173 804
rect 4187 796 4413 804
rect 4427 796 4633 804
rect 1727 776 1844 784
rect 1867 776 1933 784
rect 1947 776 1993 784
rect 2067 776 2253 784
rect 3087 776 3113 784
rect 3147 776 3193 784
rect 3947 776 4073 784
rect 4387 776 4693 784
rect 607 756 653 764
rect 667 756 733 764
rect 1047 756 1133 764
rect 1287 756 1393 764
rect 1427 756 1613 764
rect 1747 756 1833 764
rect 2007 756 2193 764
rect 2207 756 2433 764
rect 3007 756 3073 764
rect 3347 756 3393 764
rect 4207 756 4453 764
rect 487 736 533 744
rect 547 736 553 744
rect 567 736 773 744
rect 1247 736 1433 744
rect 1487 736 1753 744
rect 1987 736 2133 744
rect 2287 736 2573 744
rect 547 716 993 724
rect 1247 716 1684 724
rect 227 696 253 704
rect 267 696 393 704
rect 427 696 613 704
rect 827 696 893 704
rect 967 696 1193 704
rect 1327 696 1333 704
rect 1347 696 1493 704
rect 1507 696 1653 704
rect 1676 704 1684 716
rect 1707 716 1953 724
rect 1967 716 2033 724
rect 2047 716 2533 724
rect 2927 716 2953 724
rect 2967 716 3493 724
rect 3787 716 4213 724
rect 1676 696 2053 704
rect 2107 696 2373 704
rect 2387 696 2453 704
rect 167 676 313 684
rect 327 676 353 684
rect 447 676 673 684
rect 807 676 913 684
rect 1027 676 1113 684
rect 1287 676 1353 684
rect 1447 676 1533 684
rect 1607 676 1733 684
rect 1887 676 2233 684
rect 2347 676 2373 684
rect 2387 676 2473 684
rect 3367 676 3513 684
rect 3687 676 3833 684
rect 3847 676 3933 684
rect 3947 676 4033 684
rect 4047 676 4393 684
rect 4407 676 4493 684
rect 67 656 104 664
rect 96 624 104 656
rect 147 656 164 664
rect 156 627 164 656
rect 207 656 273 664
rect 316 656 373 664
rect 196 627 204 653
rect 247 636 273 644
rect 316 627 324 656
rect 467 656 524 664
rect 367 636 493 644
rect 516 644 524 656
rect 627 656 833 664
rect 887 656 993 664
rect 1007 656 1033 664
rect 1067 656 1084 664
rect 516 636 573 644
rect 596 636 633 644
rect 96 616 133 624
rect 347 616 393 624
rect 596 624 604 636
rect 656 636 713 644
rect 487 616 504 624
rect 496 607 504 616
rect 516 616 604 624
rect 187 596 213 604
rect 227 596 293 604
rect 307 596 373 604
rect 516 587 524 616
rect 656 624 664 636
rect 827 636 853 644
rect 867 636 884 644
rect 647 616 664 624
rect 876 607 884 636
rect 1027 636 1053 644
rect 1076 627 1084 656
rect 1467 656 1513 664
rect 1576 656 1593 664
rect 1107 636 1133 644
rect 1387 636 1413 644
rect 1576 644 1584 656
rect 1667 656 1713 664
rect 1787 656 1813 664
rect 2096 656 2113 664
rect 2016 644 2024 653
rect 2096 644 2104 656
rect 2327 656 2333 664
rect 2347 656 2413 664
rect 2467 656 2513 664
rect 3047 656 3193 664
rect 3207 656 3213 664
rect 3247 656 3273 664
rect 3287 656 3393 664
rect 3467 656 3493 664
rect 3507 656 3573 664
rect 3827 656 4013 664
rect 1476 636 1584 644
rect 1736 636 2024 644
rect 2076 636 2104 644
rect 907 616 933 624
rect 987 616 1013 624
rect 1127 616 1173 624
rect 1227 616 1253 624
rect 1476 624 1484 636
rect 1307 616 1484 624
rect 1736 624 1744 636
rect 1607 616 1744 624
rect 1767 616 1844 624
rect 1836 607 1844 616
rect 2076 624 2084 636
rect 2127 636 2213 644
rect 2267 636 2304 644
rect 2296 627 2304 636
rect 2407 636 2473 644
rect 2676 627 2684 653
rect 2707 636 2773 644
rect 2787 636 2933 644
rect 3187 636 3253 644
rect 3307 636 3413 644
rect 3547 636 3673 644
rect 3887 636 3913 644
rect 3967 636 4033 644
rect 4107 636 4153 644
rect 4667 636 4673 644
rect 4687 636 4713 644
rect 2007 616 2084 624
rect 2107 616 2144 624
rect 787 596 853 604
rect 1087 596 1373 604
rect 1467 596 1573 604
rect 1727 596 1753 604
rect 1987 596 2113 604
rect 2136 604 2144 616
rect 2307 616 2353 624
rect 2376 616 2453 624
rect 2136 596 2153 604
rect 287 576 513 584
rect 547 576 893 584
rect 1427 576 1673 584
rect 1756 584 1764 593
rect 2176 587 2184 613
rect 2207 596 2273 604
rect 2376 604 2384 616
rect 2487 616 2513 624
rect 2696 616 2733 624
rect 2307 596 2384 604
rect 2507 596 2553 604
rect 2696 604 2704 616
rect 3107 616 3153 624
rect 3167 616 3273 624
rect 3307 616 3373 624
rect 3467 616 3513 624
rect 3567 616 3813 624
rect 3907 616 3973 624
rect 4247 616 4273 624
rect 4367 616 4433 624
rect 2667 596 2704 604
rect 3067 596 3233 604
rect 4007 596 4033 604
rect 4227 596 4253 604
rect 1687 576 1764 584
rect 1787 576 1853 584
rect 1907 576 2164 584
rect 567 556 2093 564
rect 2156 564 2164 576
rect 2456 584 2464 593
rect 2187 576 2464 584
rect 2716 564 2724 593
rect 3187 576 3213 584
rect 3927 576 4093 584
rect 2156 556 2724 564
rect 707 536 773 544
rect 1127 536 1153 544
rect 1167 536 1493 544
rect 1527 536 1653 544
rect 1676 536 1813 544
rect 327 516 473 524
rect 1367 516 1533 524
rect 1567 516 1593 524
rect 1676 524 1684 536
rect 1827 536 2013 544
rect 2047 536 2173 544
rect 2687 536 2733 544
rect 3807 536 3993 544
rect 1647 516 1684 524
rect 1707 516 1833 524
rect 2067 516 2133 524
rect 4487 516 4693 524
rect 367 496 433 504
rect 527 496 613 504
rect 627 496 1073 504
rect 1227 496 1733 504
rect 1847 496 2413 504
rect 447 476 493 484
rect 1727 476 1773 484
rect 1807 476 1993 484
rect 2147 476 2173 484
rect 2187 476 2293 484
rect 327 456 513 464
rect 527 456 873 464
rect 1407 456 1873 464
rect 1927 456 2193 464
rect 407 436 633 444
rect 987 436 1273 444
rect 1367 436 1593 444
rect 1607 436 1853 444
rect 1927 436 2273 444
rect 247 416 333 424
rect 547 416 593 424
rect 887 416 993 424
rect 1147 416 1353 424
rect 1387 416 1693 424
rect 1727 416 1893 424
rect 2047 416 2113 424
rect 2127 416 2413 424
rect 2567 416 2633 424
rect 2647 416 2873 424
rect 3487 416 3893 424
rect 3907 416 4293 424
rect 4307 416 4473 424
rect 4487 416 4533 424
rect 107 396 433 404
rect 467 396 653 404
rect 707 396 853 404
rect 867 396 933 404
rect 947 396 1173 404
rect 1467 396 1633 404
rect 1667 396 1804 404
rect 167 376 193 384
rect 316 376 353 384
rect 227 356 253 364
rect 316 347 324 376
rect 387 376 453 384
rect 507 376 724 384
rect 407 356 593 364
rect 716 347 724 376
rect 907 376 1004 384
rect 836 364 844 373
rect 836 356 953 364
rect 107 336 173 344
rect 187 336 293 344
rect 427 336 713 344
rect 87 316 253 324
rect 267 316 353 324
rect 447 316 473 324
rect 527 316 633 324
rect 776 324 784 353
rect 996 344 1004 376
rect 1127 376 1244 384
rect 1027 356 1133 364
rect 1236 347 1244 376
rect 1287 376 1333 384
rect 1587 376 1664 384
rect 1256 347 1264 373
rect 1327 356 1353 364
rect 1407 356 1424 364
rect 1416 347 1424 356
rect 1456 356 1533 364
rect 827 336 964 344
rect 996 336 1153 344
rect 707 316 784 324
rect 807 316 913 324
rect 956 324 964 336
rect 1456 327 1464 356
rect 1556 344 1564 373
rect 1487 336 1564 344
rect 956 316 993 324
rect 1067 316 1113 324
rect 1187 316 1413 324
rect 1636 324 1644 353
rect 1487 316 1644 324
rect 1656 324 1664 376
rect 1796 384 1804 396
rect 1827 396 1913 404
rect 1967 396 2333 404
rect 2587 396 2693 404
rect 2767 396 3613 404
rect 3647 396 3793 404
rect 4287 396 4353 404
rect 1687 376 1784 384
rect 1796 376 1824 384
rect 1687 356 1713 364
rect 1727 356 1753 364
rect 1776 344 1784 376
rect 1816 347 1824 376
rect 1947 376 1993 384
rect 2107 376 2213 384
rect 2347 376 2444 384
rect 1887 356 2013 364
rect 2027 356 2053 364
rect 1747 336 1784 344
rect 1847 336 1913 344
rect 2076 344 2084 373
rect 2436 367 2444 376
rect 2507 376 2533 384
rect 2556 376 2733 384
rect 2147 356 2193 364
rect 2247 356 2384 364
rect 2067 336 2273 344
rect 2327 336 2353 344
rect 2376 344 2384 356
rect 2556 364 2564 376
rect 2676 367 2684 376
rect 2867 376 2893 384
rect 2947 376 3013 384
rect 3027 376 3113 384
rect 3316 376 3353 384
rect 3316 367 3324 376
rect 3407 376 3473 384
rect 4327 376 4373 384
rect 2456 356 2564 364
rect 2376 336 2433 344
rect 1656 316 1673 324
rect 1707 316 1853 324
rect 2027 316 2213 324
rect 2456 324 2464 356
rect 2587 356 2633 364
rect 2696 356 2773 364
rect 2696 344 2704 356
rect 2927 356 3073 364
rect 3756 364 3764 373
rect 3707 356 3764 364
rect 3787 356 3833 364
rect 4087 356 4333 364
rect 4447 356 4493 364
rect 2487 336 2704 344
rect 2767 336 2793 344
rect 2847 336 2873 344
rect 3147 336 3173 344
rect 3356 344 3364 353
rect 3247 336 3364 344
rect 3436 344 3444 353
rect 3436 336 3513 344
rect 3627 336 3853 344
rect 4087 336 4113 344
rect 4267 336 4393 344
rect 2387 316 2464 324
rect 2667 316 2713 324
rect 2827 316 2853 324
rect 3067 316 3413 324
rect 3467 316 3533 324
rect 3547 316 3593 324
rect 3607 316 3653 324
rect 4047 316 4133 324
rect 4496 324 4504 353
rect 4487 316 4504 324
rect 487 296 753 304
rect 827 296 1033 304
rect 1047 296 1133 304
rect 1267 296 1493 304
rect 1507 296 1693 304
rect 1767 296 1953 304
rect 2007 296 2033 304
rect 2147 296 2253 304
rect 2267 296 2393 304
rect 2547 296 2973 304
rect 3107 296 3353 304
rect 3507 296 3573 304
rect 3587 296 3733 304
rect 3747 296 3933 304
rect 3987 296 4113 304
rect 4427 296 4673 304
rect 367 276 953 284
rect 1207 276 1333 284
rect 1347 276 1433 284
rect 1447 276 1533 284
rect 1607 276 1793 284
rect 2207 276 2253 284
rect 3207 276 3513 284
rect 3887 276 4193 284
rect 367 256 553 264
rect 927 256 1373 264
rect 1407 256 1473 264
rect 1587 256 1653 264
rect 1667 256 1773 264
rect 1787 256 1873 264
rect 1987 256 2393 264
rect 2407 256 2653 264
rect 2667 256 2693 264
rect 3287 256 3573 264
rect 3927 256 3973 264
rect 3987 256 4033 264
rect 427 236 733 244
rect 907 236 1273 244
rect 1287 236 1373 244
rect 1427 236 1633 244
rect 1707 236 2073 244
rect 2967 236 3013 244
rect 3347 236 3733 244
rect 687 216 813 224
rect 867 216 893 224
rect 1027 216 1093 224
rect 1127 216 2013 224
rect 2147 216 2173 224
rect 2187 216 2193 224
rect 2207 216 2453 224
rect 3087 216 3153 224
rect 3967 216 4373 224
rect 47 196 133 204
rect 247 196 553 204
rect 627 196 853 204
rect 967 196 1033 204
rect 1087 196 1213 204
rect 1307 196 1533 204
rect 1627 196 1773 204
rect 2107 196 2153 204
rect 2187 196 2253 204
rect 2367 196 2413 204
rect 2567 196 2773 204
rect 3047 196 3193 204
rect 3207 196 4513 204
rect 87 176 113 184
rect 267 176 313 184
rect 447 176 473 184
rect 487 176 533 184
rect 547 176 633 184
rect 807 176 973 184
rect 1007 176 1313 184
rect 1447 176 1493 184
rect 1527 176 1673 184
rect 1707 176 1733 184
rect 1967 176 2053 184
rect 2087 176 2353 184
rect 2607 176 2853 184
rect 3047 176 3393 184
rect 3407 176 3693 184
rect 3807 176 3833 184
rect 3847 176 3993 184
rect 4027 176 4173 184
rect 4207 176 4333 184
rect 4427 176 4453 184
rect 4467 176 4493 184
rect 4527 176 4613 184
rect 107 156 164 164
rect 156 147 164 156
rect 187 156 293 164
rect 307 156 313 164
rect 336 147 344 173
rect 387 156 493 164
rect 507 156 593 164
rect 616 156 733 164
rect 87 136 113 144
rect 287 136 333 144
rect 467 136 513 144
rect 616 144 624 156
rect 756 147 764 173
rect 776 164 784 173
rect 776 156 864 164
rect 567 136 624 144
rect 807 136 833 144
rect 856 144 864 156
rect 887 156 913 164
rect 936 156 1093 164
rect 936 147 944 156
rect 1107 156 1333 164
rect 1447 156 1553 164
rect 1596 156 1753 164
rect 856 136 904 144
rect 516 124 524 133
rect 47 116 524 124
rect 516 104 524 116
rect 607 116 653 124
rect 667 116 873 124
rect 896 124 904 136
rect 987 136 1053 144
rect 1067 136 1113 144
rect 1156 136 1193 144
rect 896 116 993 124
rect 1156 124 1164 136
rect 1207 136 1233 144
rect 1336 136 1433 144
rect 1007 116 1164 124
rect 1236 116 1253 124
rect 516 96 613 104
rect 1236 104 1244 116
rect 1336 124 1344 136
rect 1487 136 1533 144
rect 1307 116 1344 124
rect 1576 124 1584 133
rect 1596 127 1604 156
rect 1927 156 1973 164
rect 2027 156 2213 164
rect 2327 156 2593 164
rect 2416 147 2424 156
rect 2787 156 2824 164
rect 1627 136 1673 144
rect 1707 136 1733 144
rect 1936 136 2173 144
rect 1527 116 1584 124
rect 1647 116 1713 124
rect 1727 116 1753 124
rect 1827 116 1893 124
rect 1936 124 1944 136
rect 2207 136 2333 144
rect 2587 136 2713 144
rect 2727 136 2753 144
rect 2816 144 2824 156
rect 3087 156 3113 164
rect 3287 156 3473 164
rect 3487 156 3533 164
rect 3587 156 3613 164
rect 3827 156 3873 164
rect 3887 156 3893 164
rect 3907 156 3993 164
rect 4016 156 4073 164
rect 2816 136 2873 144
rect 3147 136 3233 144
rect 4016 144 4024 156
rect 4487 156 4533 164
rect 3807 136 4024 144
rect 4216 144 4224 153
rect 4067 136 4253 144
rect 4307 136 4433 144
rect 4587 136 4644 144
rect 1927 116 1944 124
rect 2267 116 2533 124
rect 2547 116 2613 124
rect 1356 104 1364 113
rect 847 96 1364 104
rect 1407 96 1693 104
rect 1807 96 1993 104
rect 2247 96 2473 104
rect 2796 104 2804 133
rect 3927 116 3973 124
rect 4636 124 4644 136
rect 4667 136 4753 144
rect 4636 116 4693 124
rect 2487 96 2804 104
rect 4447 96 4733 104
rect 987 76 1473 84
rect 1847 76 1913 84
rect 2067 76 2293 84
rect 2747 76 2813 84
rect 1227 56 1513 64
rect 1767 56 2113 64
rect 867 36 1873 44
rect 1887 36 1933 44
rect 1327 16 1973 24
rect 2127 16 2153 24
use NOR2X1  _760_
timestamp 0
transform -1 0 4010 0 1 2650
box -6 -8 86 248
use INVX1  _761_
timestamp 0
transform -1 0 4190 0 1 3130
box -6 -8 66 248
use NOR2X1  _762_
timestamp 0
transform 1 0 3750 0 -1 3130
box -6 -8 86 248
use OAI21X1  _763_
timestamp 0
transform 1 0 4030 0 -1 3130
box -6 -8 106 248
use INVX2  _764_
timestamp 0
transform -1 0 3570 0 1 2650
box -6 -8 66 248
use NOR2X1  _765_
timestamp 0
transform -1 0 3090 0 -1 3130
box -6 -8 86 248
use AOI22X1  _766_
timestamp 0
transform -1 0 4070 0 1 2170
box -6 -8 126 248
use OAI21X1  _767_
timestamp 0
transform 1 0 4010 0 1 2650
box -6 -8 106 248
use INVX1  _768_
timestamp 0
transform 1 0 4230 0 -1 3130
box -6 -8 66 248
use INVX1  _769_
timestamp 0
transform -1 0 4410 0 -1 4090
box -6 -8 66 248
use NAND2X1  _770_
timestamp 0
transform -1 0 4530 0 1 3130
box -6 -8 86 248
use OAI21X1  _771_
timestamp 0
transform 1 0 4350 0 1 3130
box -6 -8 106 248
use AOI22X1  _772_
timestamp 0
transform -1 0 3950 0 1 2170
box -6 -8 126 248
use OAI21X1  _773_
timestamp 0
transform -1 0 4290 0 1 3130
box -6 -8 106 248
use NOR2X1  _774_
timestamp 0
transform 1 0 4210 0 1 2650
box -6 -8 86 248
use OAI21X1  _775_
timestamp 0
transform 1 0 4130 0 -1 3130
box -6 -8 106 248
use AOI22X1  _776_
timestamp 0
transform -1 0 3930 0 1 2650
box -6 -8 126 248
use OAI21X1  _777_
timestamp 0
transform -1 0 4210 0 1 2650
box -6 -8 106 248
use INVX1  _778_
timestamp 0
transform -1 0 4050 0 1 250
box -6 -8 66 248
use NAND2X1  _779_
timestamp 0
transform -1 0 3970 0 1 3130
box -6 -8 86 248
use OAI21X1  _780_
timestamp 0
transform -1 0 4030 0 -1 3130
box -6 -8 106 248
use AOI22X1  _781_
timestamp 0
transform 1 0 3330 0 -1 2650
box -6 -8 126 248
use OAI21X1  _782_
timestamp 0
transform -1 0 3930 0 -1 3130
box -6 -8 106 248
use INVX2  _783_
timestamp 0
transform -1 0 770 0 1 2650
box -6 -8 66 248
use NAND2X1  _784_
timestamp 0
transform 1 0 1810 0 -1 2650
box -6 -8 86 248
use OAI21X1  _785_
timestamp 0
transform 1 0 1750 0 -1 3130
box -6 -8 106 248
use INVX2  _786_
timestamp 0
transform 1 0 1430 0 -1 2650
box -6 -8 66 248
use NAND2X1  _787_
timestamp 0
transform 1 0 1890 0 -1 2650
box -6 -8 86 248
use OAI21X1  _788_
timestamp 0
transform 1 0 1790 0 1 2650
box -6 -8 106 248
use INVX2  _789_
timestamp 0
transform 1 0 1890 0 -1 3610
box -6 -8 66 248
use NAND2X1  _790_
timestamp 0
transform -1 0 2350 0 -1 3130
box -6 -8 86 248
use OAI21X1  _791_
timestamp 0
transform 1 0 2350 0 -1 3130
box -6 -8 106 248
use INVX2  _792_
timestamp 0
transform -1 0 710 0 1 2650
box -6 -8 66 248
use NAND2X1  _793_
timestamp 0
transform -1 0 1790 0 -1 3610
box -6 -8 86 248
use OAI21X1  _794_
timestamp 0
transform 1 0 1790 0 -1 3610
box -6 -8 106 248
use NAND2X1  _795_
timestamp 0
transform 1 0 1050 0 1 2650
box -6 -8 86 248
use OAI21X1  _796_
timestamp 0
transform -1 0 1230 0 1 2650
box -6 -8 106 248
use NAND2X1  _797_
timestamp 0
transform 1 0 570 0 -1 3130
box -6 -8 86 248
use OAI21X1  _798_
timestamp 0
transform 1 0 470 0 -1 3130
box -6 -8 106 248
use NAND2X1  _799_
timestamp 0
transform 1 0 1290 0 -1 3610
box -6 -8 86 248
use OAI21X1  _800_
timestamp 0
transform 1 0 1370 0 -1 3610
box -6 -8 106 248
use NAND2X1  _801_
timestamp 0
transform 1 0 670 0 -1 3610
box -6 -8 86 248
use OAI21X1  _802_
timestamp 0
transform -1 0 790 0 1 3130
box -6 -8 106 248
use INVX1  _803_
timestamp 0
transform -1 0 4530 0 1 250
box -6 -8 66 248
use NAND2X1  _804_
timestamp 0
transform 1 0 4250 0 -1 730
box -6 -8 86 248
use OAI21X1  _805_
timestamp 0
transform -1 0 4470 0 1 250
box -6 -8 106 248
use INVX1  _806_
timestamp 0
transform 1 0 3830 0 -1 250
box -6 -8 66 248
use NAND2X1  _807_
timestamp 0
transform -1 0 3490 0 -1 730
box -6 -8 86 248
use OAI21X1  _808_
timestamp 0
transform -1 0 3590 0 -1 730
box -6 -8 106 248
use INVX1  _809_
timestamp 0
transform -1 0 3290 0 1 250
box -6 -8 66 248
use NAND2X1  _810_
timestamp 0
transform -1 0 3350 0 -1 1690
box -6 -8 86 248
use OAI21X1  _811_
timestamp 0
transform -1 0 3390 0 1 250
box -6 -8 106 248
use INVX1  _812_
timestamp 0
transform 1 0 3150 0 1 730
box -6 -8 66 248
use NAND2X1  _813_
timestamp 0
transform 1 0 3010 0 -1 1210
box -6 -8 86 248
use OAI21X1  _814_
timestamp 0
transform -1 0 3190 0 -1 1210
box -6 -8 106 248
use INVX1  _815_
timestamp 0
transform -1 0 3090 0 -1 1690
box -6 -8 66 248
use NAND2X1  _816_
timestamp 0
transform 1 0 3190 0 -1 1690
box -6 -8 86 248
use OAI21X1  _817_
timestamp 0
transform 1 0 3090 0 -1 1690
box -6 -8 106 248
use INVX1  _818_
timestamp 0
transform 1 0 2250 0 1 1690
box -6 -8 66 248
use NAND2X1  _819_
timestamp 0
transform 1 0 2390 0 -1 2170
box -6 -8 86 248
use OAI21X1  _820_
timestamp 0
transform 1 0 2310 0 1 1690
box -6 -8 106 248
use INVX1  _821_
timestamp 0
transform 1 0 2450 0 -1 3130
box -6 -8 66 248
use NAND2X1  _822_
timestamp 0
transform 1 0 2690 0 -1 3130
box -6 -8 86 248
use OAI21X1  _823_
timestamp 0
transform 1 0 2510 0 -1 3130
box -6 -8 106 248
use INVX1  _824_
timestamp 0
transform 1 0 2370 0 -1 3610
box -6 -8 66 248
use NAND2X1  _825_
timestamp 0
transform 1 0 2850 0 -1 3610
box -6 -8 86 248
use OAI21X1  _826_
timestamp 0
transform 1 0 2670 0 -1 3610
box -6 -8 106 248
use INVX1  _827_
timestamp 0
transform 1 0 2850 0 1 4090
box -6 -8 66 248
use NAND2X1  _828_
timestamp 0
transform 1 0 3090 0 1 4090
box -6 -8 86 248
use OAI21X1  _829_
timestamp 0
transform 1 0 2990 0 1 4090
box -6 -8 106 248
use INVX1  _830_
timestamp 0
transform -1 0 3430 0 -1 4570
box -6 -8 66 248
use NAND2X1  _831_
timestamp 0
transform 1 0 3770 0 -1 4570
box -6 -8 86 248
use OAI21X1  _832_
timestamp 0
transform 1 0 3670 0 -1 4570
box -6 -8 106 248
use INVX1  _833_
timestamp 0
transform 1 0 2890 0 -1 4090
box -6 -8 66 248
use NAND2X1  _834_
timestamp 0
transform 1 0 3130 0 -1 4090
box -6 -8 86 248
use OAI21X1  _835_
timestamp 0
transform 1 0 2950 0 -1 4090
box -6 -8 106 248
use INVX1  _836_
timestamp 0
transform 1 0 4210 0 -1 4570
box -6 -8 66 248
use NAND2X1  _837_
timestamp 0
transform 1 0 4130 0 -1 4570
box -6 -8 86 248
use OAI21X1  _838_
timestamp 0
transform 1 0 4270 0 -1 4570
box -6 -8 106 248
use INVX1  _839_
timestamp 0
transform 1 0 3730 0 1 1210
box -6 -8 66 248
use NAND2X1  _840_
timestamp 0
transform 1 0 4130 0 1 1210
box -6 -8 86 248
use OAI21X1  _841_
timestamp 0
transform 1 0 4030 0 1 1210
box -6 -8 106 248
use INVX1  _842_
timestamp 0
transform -1 0 4590 0 -1 1690
box -6 -8 66 248
use NAND2X1  _843_
timestamp 0
transform 1 0 4650 0 -1 2650
box -6 -8 86 248
use OAI21X1  _844_
timestamp 0
transform 1 0 4630 0 -1 3610
box -6 -8 106 248
use INVX1  _845_
timestamp 0
transform 1 0 4650 0 1 1210
box -6 -8 66 248
use NAND2X1  _846_
timestamp 0
transform -1 0 4750 0 1 1690
box -6 -8 86 248
use OAI21X1  _847_
timestamp 0
transform 1 0 4630 0 1 730
box -6 -8 106 248
use INVX1  _848_
timestamp 0
transform -1 0 4690 0 -1 250
box -6 -8 66 248
use NAND2X1  _849_
timestamp 0
transform 1 0 4690 0 -1 1690
box -6 -8 86 248
use OAI21X1  _850_
timestamp 0
transform 1 0 4530 0 1 730
box -6 -8 106 248
use INVX1  _851_
timestamp 0
transform 1 0 3150 0 -1 250
box -6 -8 66 248
use NAND3X1  _852_
timestamp 0
transform 1 0 2430 0 1 250
box -6 -8 106 248
use OAI21X1  _853_
timestamp 0
transform -1 0 3050 0 1 250
box -6 -8 106 248
use INVX1  _854_
timestamp 0
transform -1 0 3990 0 1 250
box -6 -8 66 248
use NAND2X1  _855_
timestamp 0
transform -1 0 2350 0 1 250
box -6 -8 86 248
use NAND2X1  _856_
timestamp 0
transform 1 0 2110 0 1 250
box -6 -8 86 248
use NOR2X1  _857_
timestamp 0
transform 1 0 2350 0 1 250
box -6 -8 86 248
use INVX1  _858_
timestamp 0
transform -1 0 2690 0 -1 730
box -6 -8 66 248
use INVX1  _859_
timestamp 0
transform -1 0 1870 0 1 730
box -6 -8 66 248
use INVX2  _860_
timestamp 0
transform -1 0 690 0 1 1690
box -6 -8 66 248
use OAI21X1  _861_
timestamp 0
transform 1 0 1830 0 -1 730
box -6 -8 106 248
use NAND3X1  _862_
timestamp 0
transform 1 0 2690 0 -1 730
box -6 -8 106 248
use OAI21X1  _863_
timestamp 0
transform -1 0 3930 0 1 250
box -6 -8 106 248
use INVX1  _864_
timestamp 0
transform -1 0 3270 0 -1 250
box -6 -8 66 248
use NAND2X1  _865_
timestamp 0
transform 1 0 1950 0 1 250
box -6 -8 86 248
use NAND2X1  _866_
timestamp 0
transform 1 0 2030 0 1 250
box -6 -8 86 248
use NOR2X1  _867_
timestamp 0
transform -1 0 2270 0 1 250
box -6 -8 86 248
use AOI22X1  _868_
timestamp 0
transform 1 0 2270 0 -1 250
box -6 -8 126 248
use OAI21X1  _869_
timestamp 0
transform 1 0 2590 0 -1 250
box -6 -8 106 248
use INVX1  _870_
timestamp 0
transform 1 0 2690 0 -1 250
box -6 -8 66 248
use AND2X2  _871_
timestamp 0
transform -1 0 2090 0 -1 250
box -6 -8 106 248
use NAND3X1  _872_
timestamp 0
transform 1 0 2170 0 -1 250
box -6 -8 106 248
use INVX1  _873_
timestamp 0
transform 1 0 2850 0 -1 250
box -6 -8 66 248
use NAND3X1  _874_
timestamp 0
transform 1 0 2750 0 -1 250
box -6 -8 106 248
use NAND3X1  _875_
timestamp 0
transform -1 0 2690 0 1 250
box -6 -8 106 248
use INVX1  _876_
timestamp 0
transform -1 0 2590 0 1 250
box -6 -8 66 248
use AOI21X1  _877_
timestamp 0
transform 1 0 2690 0 1 250
box -6 -8 106 248
use NOR2X1  _878_
timestamp 0
transform 1 0 2790 0 1 250
box -6 -8 86 248
use NAND2X1  _879_
timestamp 0
transform -1 0 2950 0 1 250
box -6 -8 86 248
use OAI21X1  _880_
timestamp 0
transform -1 0 3150 0 1 250
box -6 -8 106 248
use INVX1  _881_
timestamp 0
transform -1 0 2990 0 1 730
box -6 -8 66 248
use NAND2X1  _882_
timestamp 0
transform -1 0 1950 0 1 730
box -6 -8 86 248
use AOI21X1  _883_
timestamp 0
transform -1 0 2590 0 -1 250
box -6 -8 106 248
use NAND2X1  _884_
timestamp 0
transform 1 0 1830 0 -1 250
box -6 -8 86 248
use NAND2X1  _885_
timestamp 0
transform 1 0 890 0 1 250
box -6 -8 86 248
use NOR2X1  _886_
timestamp 0
transform -1 0 1430 0 1 250
box -6 -8 86 248
use AOI22X1  _887_
timestamp 0
transform -1 0 1250 0 1 250
box -6 -8 126 248
use OAI21X1  _888_
timestamp 0
transform 1 0 1430 0 1 250
box -6 -8 106 248
use INVX1  _889_
timestamp 0
transform 1 0 1690 0 1 250
box -6 -8 66 248
use AND2X2  _890_
timestamp 0
transform 1 0 810 0 -1 730
box -6 -8 106 248
use NAND2X1  _891_
timestamp 0
transform -1 0 1050 0 1 250
box -6 -8 86 248
use INVX1  _892_
timestamp 0
transform 1 0 1530 0 1 250
box -6 -8 66 248
use NAND3X1  _893_
timestamp 0
transform 1 0 1750 0 1 250
box -6 -8 106 248
use NAND3X1  _894_
timestamp 0
transform 1 0 2430 0 -1 730
box -6 -8 106 248
use OAI21X1  _895_
timestamp 0
transform 1 0 2390 0 -1 250
box -6 -8 106 248
use AOI21X1  _896_
timestamp 0
transform 1 0 1850 0 1 250
box -6 -8 106 248
use INVX2  _897_
timestamp 0
transform -1 0 1170 0 -1 730
box -6 -8 66 248
use OAI21X1  _898_
timestamp 0
transform -1 0 1110 0 -1 730
box -6 -8 106 248
use INVX2  _899_
timestamp 0
transform -1 0 730 0 -1 2650
box -6 -8 66 248
use INVX1  _900_
timestamp 0
transform 1 0 490 0 1 730
box -6 -8 66 248
use OAI21X1  _901_
timestamp 0
transform 1 0 910 0 -1 730
box -6 -8 106 248
use AOI21X1  _902_
timestamp 0
transform 1 0 1170 0 -1 730
box -6 -8 106 248
use OAI21X1  _903_
timestamp 0
transform -1 0 2330 0 -1 730
box -6 -8 106 248
use NAND3X1  _904_
timestamp 0
transform 1 0 2530 0 -1 730
box -6 -8 106 248
use INVX1  _905_
timestamp 0
transform 1 0 1950 0 1 730
box -6 -8 66 248
use NAND3X1  _906_
timestamp 0
transform -1 0 2230 0 -1 730
box -6 -8 106 248
use OAI21X1  _907_
timestamp 0
transform 1 0 2330 0 -1 730
box -6 -8 106 248
use NAND3X1  _908_
timestamp 0
transform 1 0 2430 0 1 730
box -6 -8 106 248
use AOI21X1  _909_
timestamp 0
transform 1 0 2630 0 1 730
box -6 -8 106 248
use NAND3X1  _910_
timestamp 0
transform -1 0 2630 0 1 730
box -6 -8 106 248
use NAND2X1  _911_
timestamp 0
transform -1 0 2810 0 1 730
box -6 -8 86 248
use OAI22X1  _912_
timestamp 0
transform -1 0 2930 0 1 730
box -6 -8 126 248
use INVX1  _913_
timestamp 0
transform -1 0 3030 0 -1 1690
box -6 -8 66 248
use INVX1  _914_
timestamp 0
transform -1 0 2490 0 -1 1210
box -6 -8 66 248
use AOI21X1  _915_
timestamp 0
transform -1 0 2030 0 -1 730
box -6 -8 106 248
use OAI21X1  _916_
timestamp 0
transform 1 0 2030 0 -1 730
box -6 -8 106 248
use OAI21X1  _917_
timestamp 0
transform 1 0 1250 0 1 250
box -6 -8 106 248
use AND2X2  _918_
timestamp 0
transform -1 0 430 0 1 250
box -6 -8 106 248
use NAND2X1  _919_
timestamp 0
transform -1 0 890 0 1 250
box -6 -8 86 248
use AOI22X1  _920_
timestamp 0
transform -1 0 730 0 1 250
box -6 -8 126 248
use INVX1  _921_
timestamp 0
transform 1 0 810 0 -1 250
box -6 -8 66 248
use NAND2X1  _922_
timestamp 0
transform -1 0 1130 0 1 250
box -6 -8 86 248
use INVX1  _923_
timestamp 0
transform -1 0 1030 0 -1 250
box -6 -8 66 248
use NAND3X1  _924_
timestamp 0
transform 1 0 1230 0 -1 250
box -6 -8 106 248
use NAND2X1  _925_
timestamp 0
transform -1 0 510 0 1 250
box -6 -8 86 248
use NOR2X1  _926_
timestamp 0
transform -1 0 810 0 1 250
box -6 -8 86 248
use OAI21X1  _927_
timestamp 0
transform 1 0 1030 0 -1 250
box -6 -8 106 248
use AOI21X1  _928_
timestamp 0
transform -1 0 1530 0 -1 250
box -6 -8 106 248
use AOI21X1  _929_
timestamp 0
transform -1 0 1690 0 1 250
box -6 -8 106 248
use NAND3X1  _930_
timestamp 0
transform 1 0 1330 0 -1 250
box -6 -8 106 248
use OAI21X1  _931_
timestamp 0
transform 1 0 1130 0 -1 250
box -6 -8 106 248
use AOI21X1  _932_
timestamp 0
transform -1 0 1730 0 -1 250
box -6 -8 106 248
use NAND2X1  _933_
timestamp 0
transform 1 0 1530 0 1 730
box -6 -8 86 248
use INVX2  _934_
timestamp 0
transform -1 0 1510 0 -1 1210
box -6 -8 66 248
use NAND2X1  _935_
timestamp 0
transform 1 0 1690 0 1 1210
box -6 -8 86 248
use OAI21X1  _936_
timestamp 0
transform 1 0 1590 0 1 1210
box -6 -8 106 248
use OAI21X1  _937_
timestamp 0
transform -1 0 1710 0 1 730
box -6 -8 106 248
use OAI21X1  _938_
timestamp 0
transform 1 0 1430 0 -1 730
box -6 -8 106 248
use NAND3X1  _939_
timestamp 0
transform 1 0 1730 0 -1 250
box -6 -8 106 248
use NAND3X1  _940_
timestamp 0
transform 1 0 1530 0 -1 250
box -6 -8 106 248
use INVX1  _941_
timestamp 0
transform -1 0 1330 0 -1 730
box -6 -8 66 248
use NAND3X1  _942_
timestamp 0
transform 1 0 1730 0 -1 730
box -6 -8 106 248
use NAND3X1  _943_
timestamp 0
transform -1 0 2110 0 1 730
box -6 -8 106 248
use INVX1  _944_
timestamp 0
transform 1 0 2370 0 1 730
box -6 -8 66 248
use AOI21X1  _945_
timestamp 0
transform -1 0 2370 0 1 730
box -6 -8 106 248
use AOI21X1  _946_
timestamp 0
transform 1 0 1630 0 -1 730
box -6 -8 106 248
use INVX1  _947_
timestamp 0
transform 1 0 2110 0 1 730
box -6 -8 66 248
use OAI21X1  _948_
timestamp 0
transform 1 0 2170 0 1 730
box -6 -8 106 248
use AOI21X1  _949_
timestamp 0
transform 1 0 2330 0 -1 1210
box -6 -8 106 248
use NAND3X1  _950_
timestamp 0
transform -1 0 2250 0 -1 1210
box -6 -8 106 248
use NAND2X1  _951_
timestamp 0
transform -1 0 2570 0 -1 1210
box -6 -8 86 248
use OAI22X1  _952_
timestamp 0
transform -1 0 2690 0 -1 1210
box -6 -8 126 248
use INVX1  _953_
timestamp 0
transform 1 0 2210 0 -1 1690
box -6 -8 66 248
use AND2X2  _954_
timestamp 0
transform 1 0 1710 0 1 730
box -6 -8 106 248
use NAND2X1  _955_
timestamp 0
transform 1 0 1950 0 -1 1210
box -6 -8 86 248
use INVX1  _956_
timestamp 0
transform 1 0 2070 0 1 1210
box -6 -8 66 248
use AOI21X1  _957_
timestamp 0
transform -1 0 1630 0 -1 730
box -6 -8 106 248
use NAND2X1  _958_
timestamp 0
transform -1 0 1530 0 1 730
box -6 -8 86 248
use INVX1  _959_
timestamp 0
transform -1 0 1390 0 1 1690
box -6 -8 66 248
use AND2X2  _960_
timestamp 0
transform -1 0 1370 0 -1 1210
box -6 -8 106 248
use OAI21X1  _961_
timestamp 0
transform -1 0 1190 0 -1 1210
box -6 -8 106 248
use INVX2  _962_
timestamp 0
transform -1 0 1730 0 1 1690
box -6 -8 66 248
use OAI21X1  _963_
timestamp 0
transform 1 0 1090 0 1 730
box -6 -8 106 248
use NAND3X1  _964_
timestamp 0
transform -1 0 1090 0 1 730
box -6 -8 106 248
use INVX1  _965_
timestamp 0
transform 1 0 1290 0 1 730
box -6 -8 66 248
use NAND2X1  _966_
timestamp 0
transform -1 0 1270 0 -1 1210
box -6 -8 86 248
use OAI21X1  _967_
timestamp 0
transform 1 0 1350 0 1 730
box -6 -8 106 248
use NAND3X1  _968_
timestamp 0
transform -1 0 1290 0 1 730
box -6 -8 106 248
use NAND2X1  _969_
timestamp 0
transform 1 0 910 0 1 730
box -6 -8 86 248
use AOI21X1  _970_
timestamp 0
transform -1 0 810 0 -1 250
box -6 -8 106 248
use NAND2X1  _971_
timestamp 0
transform -1 0 330 0 1 250
box -6 -8 86 248
use AND2X2  _972_
timestamp 0
transform -1 0 190 0 1 730
box -6 -8 106 248
use NAND2X1  _973_
timestamp 0
transform 1 0 90 0 1 250
box -6 -8 86 248
use NAND2X1  _974_
timestamp 0
transform -1 0 90 0 1 730
box -6 -8 86 248
use NAND2X1  _975_
timestamp 0
transform 1 0 10 0 1 250
box -6 -8 86 248
use NAND3X1  _976_
timestamp 0
transform -1 0 110 0 -1 250
box -6 -8 106 248
use INVX1  _977_
timestamp 0
transform 1 0 190 0 -1 730
box -6 -8 66 248
use NAND2X1  _978_
timestamp 0
transform -1 0 250 0 1 250
box -6 -8 86 248
use OAI21X1  _979_
timestamp 0
transform -1 0 550 0 -1 730
box -6 -8 106 248
use NAND3X1  _980_
timestamp 0
transform 1 0 350 0 -1 730
box -6 -8 106 248
use NAND3X1  _981_
timestamp 0
transform 1 0 510 0 -1 250
box -6 -8 106 248
use OAI21X1  _982_
timestamp 0
transform -1 0 970 0 -1 250
box -6 -8 106 248
use AOI21X1  _983_
timestamp 0
transform -1 0 350 0 -1 730
box -6 -8 106 248
use AOI21X1  _984_
timestamp 0
transform 1 0 110 0 -1 250
box -6 -8 106 248
use OAI21X1  _985_
timestamp 0
transform 1 0 310 0 -1 250
box -6 -8 106 248
use NAND3X1  _986_
timestamp 0
transform -1 0 610 0 1 250
box -6 -8 106 248
use AND2X2  _987_
timestamp 0
transform -1 0 910 0 1 730
box -6 -8 106 248
use NAND3X1  _988_
timestamp 0
transform -1 0 510 0 -1 250
box -6 -8 106 248
use OAI21X1  _989_
timestamp 0
transform -1 0 310 0 -1 250
box -6 -8 106 248
use NAND3X1  _990_
timestamp 0
transform 1 0 710 0 1 730
box -6 -8 106 248
use NAND3X1  _991_
timestamp 0
transform 1 0 1670 0 -1 1210
box -6 -8 106 248
use OAI21X1  _992_
timestamp 0
transform 1 0 1330 0 -1 730
box -6 -8 106 248
use NAND2X1  _993_
timestamp 0
transform -1 0 1590 0 -1 1210
box -6 -8 86 248
use NAND2X1  _994_
timestamp 0
transform -1 0 1850 0 -1 1210
box -6 -8 86 248
use NAND3X1  _995_
timestamp 0
transform 1 0 1850 0 -1 1210
box -6 -8 106 248
use NAND3X1  _996_
timestamp 0
transform 1 0 1870 0 1 1210
box -6 -8 106 248
use NAND2X1  _997_
timestamp 0
transform -1 0 1670 0 -1 1210
box -6 -8 86 248
use NAND3X1  _998_
timestamp 0
transform 1 0 2130 0 1 1210
box -6 -8 106 248
use NAND2X1  _999_
timestamp 0
transform 1 0 2230 0 1 1210
box -6 -8 86 248
use NAND2X1  _1000_
timestamp 0
transform -1 0 2330 0 -1 1210
box -6 -8 86 248
use OR2X2  _1001_
timestamp 0
transform 1 0 2310 0 1 1210
box -6 -8 106 248
use AOI22X1  _1002_
timestamp 0
transform -1 0 2150 0 -1 1210
box -6 -8 126 248
use INVX1  _1003_
timestamp 0
transform -1 0 1890 0 1 2170
box -6 -8 66 248
use NAND3X1  _1004_
timestamp 0
transform 1 0 2010 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1005_
timestamp 0
transform -1 0 2210 0 -1 1690
box -6 -8 106 248
use INVX1  _1006_
timestamp 0
transform 1 0 1890 0 1 2650
box -6 -8 66 248
use AOI21X1  _1007_
timestamp 0
transform 1 0 1770 0 1 1210
box -6 -8 106 248
use OAI21X1  _1008_
timestamp 0
transform 1 0 1970 0 1 1210
box -6 -8 106 248
use NAND2X1  _1009_
timestamp 0
transform 1 0 1510 0 1 1210
box -6 -8 86 248
use OAI21X1  _1010_
timestamp 0
transform -1 0 1510 0 1 1210
box -6 -8 106 248
use INVX1  _1011_
timestamp 0
transform -1 0 1450 0 -1 1690
box -6 -8 66 248
use INVX1  _1012_
timestamp 0
transform -1 0 610 0 1 730
box -6 -8 66 248
use AOI21X1  _1013_
timestamp 0
transform -1 0 710 0 1 730
box -6 -8 106 248
use NAND2X1  _1014_
timestamp 0
transform 1 0 1370 0 -1 1210
box -6 -8 86 248
use AND2X2  _1015_
timestamp 0
transform 1 0 790 0 1 1210
box -6 -8 106 248
use OAI21X1  _1016_
timestamp 0
transform -1 0 990 0 -1 1210
box -6 -8 106 248
use AND2X2  _1017_
timestamp 0
transform -1 0 1310 0 1 1210
box -6 -8 106 248
use OAI21X1  _1018_
timestamp 0
transform 1 0 990 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1019_
timestamp 0
transform -1 0 890 0 -1 1210
box -6 -8 106 248
use INVX1  _1020_
timestamp 0
transform -1 0 1210 0 1 1210
box -6 -8 66 248
use NAND2X1  _1021_
timestamp 0
transform -1 0 970 0 1 1210
box -6 -8 86 248
use OAI21X1  _1022_
timestamp 0
transform 1 0 1310 0 1 1210
box -6 -8 106 248
use NAND3X1  _1023_
timestamp 0
transform -1 0 1150 0 1 1210
box -6 -8 106 248
use NAND2X1  _1024_
timestamp 0
transform -1 0 690 0 -1 1210
box -6 -8 86 248
use NOR2X1  _1025_
timestamp 0
transform -1 0 90 0 -1 730
box -6 -8 86 248
use AOI21X1  _1026_
timestamp 0
transform -1 0 190 0 -1 730
box -6 -8 106 248
use NAND2X1  _1027_
timestamp 0
transform -1 0 390 0 1 1210
box -6 -8 86 248
use AND2X2  _1028_
timestamp 0
transform -1 0 370 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1029_
timestamp 0
transform -1 0 190 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1030_
timestamp 0
transform 1 0 230 0 1 1690
box -6 -8 86 248
use NAND3X1  _1031_
timestamp 0
transform -1 0 410 0 1 1690
box -6 -8 106 248
use NAND3X1  _1032_
timestamp 0
transform 1 0 110 0 1 1210
box -6 -8 106 248
use INVX1  _1033_
timestamp 0
transform -1 0 70 0 -1 1690
box -6 -8 66 248
use AND2X2  _1034_
timestamp 0
transform 1 0 530 0 1 1690
box -6 -8 106 248
use NAND2X1  _1035_
timestamp 0
transform 1 0 270 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1036_
timestamp 0
transform 1 0 130 0 1 1690
box -6 -8 106 248
use NAND3X1  _1037_
timestamp 0
transform 1 0 170 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1038_
timestamp 0
transform 1 0 210 0 -1 1210
box -6 -8 106 248
use AOI22X1  _1039_
timestamp 0
transform -1 0 410 0 1 730
box -6 -8 126 248
use OAI21X1  _1040_
timestamp 0
transform -1 0 290 0 1 730
box -6 -8 106 248
use AOI21X1  _1041_
timestamp 0
transform -1 0 170 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1042_
timestamp 0
transform -1 0 110 0 1 1210
box -6 -8 106 248
use OAI21X1  _1043_
timestamp 0
transform 1 0 110 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1044_
timestamp 0
transform 1 0 410 0 -1 1210
box -6 -8 106 248
use AND2X2  _1045_
timestamp 0
transform -1 0 790 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1046_
timestamp 0
transform 1 0 210 0 1 1210
box -6 -8 106 248
use OAI21X1  _1047_
timestamp 0
transform -1 0 110 0 -1 1210
box -6 -8 106 248
use NAND3X1  _1048_
timestamp 0
transform 1 0 590 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1049_
timestamp 0
transform 1 0 790 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1050_
timestamp 0
transform 1 0 610 0 -1 250
box -6 -8 106 248
use OAI21X1  _1051_
timestamp 0
transform -1 0 730 0 -1 730
box -6 -8 106 248
use AOI21X1  _1052_
timestamp 0
transform 1 0 490 0 1 1210
box -6 -8 106 248
use AOI21X1  _1053_
timestamp 0
transform 1 0 510 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1054_
timestamp 0
transform 1 0 690 0 1 1210
box -6 -8 106 248
use NAND3X1  _1055_
timestamp 0
transform 1 0 1190 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1056_
timestamp 0
transform 1 0 990 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1057_
timestamp 0
transform 1 0 590 0 1 1210
box -6 -8 106 248
use NAND3X1  _1058_
timestamp 0
transform 1 0 1450 0 -1 1690
box -6 -8 106 248
use NAND3X1  _1059_
timestamp 0
transform 1 0 1650 0 -1 1690
box -6 -8 106 248
use INVX1  _1060_
timestamp 0
transform 1 0 1950 0 -1 1690
box -6 -8 66 248
use AOI21X1  _1061_
timestamp 0
transform -1 0 1950 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1062_
timestamp 0
transform 1 0 1550 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1063_
timestamp 0
transform 1 0 1290 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1064_
timestamp 0
transform 1 0 1750 0 -1 1690
box -6 -8 106 248
use AND2X2  _1065_
timestamp 0
transform 1 0 1830 0 1 1690
box -6 -8 106 248
use NOR2X1  _1066_
timestamp 0
transform 1 0 2070 0 -1 2650
box -6 -8 86 248
use INVX1  _1067_
timestamp 0
transform -1 0 1950 0 1 2170
box -6 -8 66 248
use OAI21X1  _1068_
timestamp 0
transform 1 0 1950 0 1 2170
box -6 -8 106 248
use OAI22X1  _1069_
timestamp 0
transform 1 0 1950 0 1 2650
box -6 -8 126 248
use INVX1  _1070_
timestamp 0
transform -1 0 2210 0 -1 2650
box -6 -8 66 248
use NAND3X1  _1071_
timestamp 0
transform -1 0 1830 0 1 1690
box -6 -8 106 248
use AOI21X1  _1072_
timestamp 0
transform 1 0 890 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1073_
timestamp 0
transform -1 0 1190 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1074_
timestamp 0
transform 1 0 970 0 1 1210
box -6 -8 86 248
use AOI21X1  _1075_
timestamp 0
transform 1 0 310 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1076_
timestamp 0
transform 1 0 390 0 1 1210
box -6 -8 106 248
use NAND2X1  _1077_
timestamp 0
transform 1 0 1350 0 -1 2650
box -6 -8 86 248
use AND2X2  _1078_
timestamp 0
transform 1 0 950 0 1 2170
box -6 -8 106 248
use OAI21X1  _1079_
timestamp 0
transform -1 0 1150 0 1 2170
box -6 -8 106 248
use AND2X2  _1080_
timestamp 0
transform 1 0 850 0 1 2650
box -6 -8 106 248
use OAI21X1  _1081_
timestamp 0
transform -1 0 1050 0 1 2650
box -6 -8 106 248
use NAND3X1  _1082_
timestamp 0
transform -1 0 1190 0 -1 2650
box -6 -8 106 248
use INVX1  _1083_
timestamp 0
transform -1 0 1250 0 -1 2650
box -6 -8 66 248
use NAND2X1  _1084_
timestamp 0
transform 1 0 1010 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1085_
timestamp 0
transform 1 0 770 0 1 2650
box -6 -8 86 248
use OAI21X1  _1086_
timestamp 0
transform -1 0 1010 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1087_
timestamp 0
transform -1 0 910 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1088_
timestamp 0
transform 1 0 870 0 1 2170
box -6 -8 86 248
use AOI22X1  _1089_
timestamp 0
transform -1 0 130 0 1 1690
box -6 -8 126 248
use NAND2X1  _1090_
timestamp 0
transform 1 0 570 0 1 2650
box -6 -8 86 248
use AND2X2  _1091_
timestamp 0
transform 1 0 370 0 1 2650
box -6 -8 106 248
use OAI21X1  _1092_
timestamp 0
transform -1 0 570 0 1 2650
box -6 -8 106 248
use OAI21X1  _1093_
timestamp 0
transform -1 0 670 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1094_
timestamp 0
transform -1 0 570 0 -1 2650
box -6 -8 106 248
use INVX1  _1095_
timestamp 0
transform -1 0 270 0 -1 2650
box -6 -8 66 248
use NAND2X1  _1096_
timestamp 0
transform 1 0 290 0 1 2650
box -6 -8 86 248
use AOI22X1  _1097_
timestamp 0
transform 1 0 170 0 1 2650
box -6 -8 126 248
use INVX1  _1098_
timestamp 0
transform -1 0 70 0 1 2650
box -6 -8 66 248
use NAND3X1  _1099_
timestamp 0
transform 1 0 10 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1100_
timestamp 0
transform -1 0 110 0 1 2170
box -6 -8 106 248
use AOI22X1  _1101_
timestamp 0
transform 1 0 410 0 1 1690
box -6 -8 126 248
use OAI21X1  _1102_
timestamp 0
transform -1 0 450 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1103_
timestamp 0
transform 1 0 110 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1104_
timestamp 0
transform -1 0 470 0 -1 2650
box -6 -8 106 248
use OAI21X1  _1105_
timestamp 0
transform 1 0 210 0 1 2170
box -6 -8 106 248
use NAND3X1  _1106_
timestamp 0
transform -1 0 290 0 -1 2170
box -6 -8 106 248
use AND2X2  _1107_
timestamp 0
transform -1 0 870 0 1 2170
box -6 -8 106 248
use NAND3X1  _1108_
timestamp 0
transform 1 0 310 0 1 2170
box -6 -8 106 248
use OAI21X1  _1109_
timestamp 0
transform -1 0 210 0 1 2170
box -6 -8 106 248
use NAND3X1  _1110_
timestamp 0
transform 1 0 490 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1111_
timestamp 0
transform 1 0 590 0 -1 2170
box -6 -8 106 248
use INVX1  _1112_
timestamp 0
transform -1 0 590 0 -1 1690
box -6 -8 66 248
use AOI21X1  _1113_
timestamp 0
transform 1 0 690 0 -1 1690
box -6 -8 106 248
use AOI21X1  _1114_
timestamp 0
transform 1 0 390 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1115_
timestamp 0
transform 1 0 290 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1116_
timestamp 0
transform 1 0 870 0 1 1690
box -6 -8 106 248
use NAND3X1  _1117_
timestamp 0
transform 1 0 990 0 -1 2170
box -6 -8 106 248
use INVX1  _1118_
timestamp 0
transform 1 0 1070 0 1 1690
box -6 -8 66 248
use NAND3X1  _1119_
timestamp 0
transform 1 0 970 0 1 1690
box -6 -8 106 248
use OAI21X1  _1120_
timestamp 0
transform -1 0 870 0 1 1690
box -6 -8 106 248
use NAND3X1  _1121_
timestamp 0
transform 1 0 1130 0 1 1690
box -6 -8 106 248
use AOI21X1  _1122_
timestamp 0
transform 1 0 1190 0 -1 2170
box -6 -8 106 248
use NAND3X1  _1123_
timestamp 0
transform 1 0 1230 0 1 1690
box -6 -8 106 248
use NAND3X1  _1124_
timestamp 0
transform 1 0 890 0 -1 2170
box -6 -8 106 248
use AOI22X1  _1125_
timestamp 0
transform -1 0 1510 0 1 1690
box -6 -8 126 248
use NOR2X1  _1126_
timestamp 0
transform 1 0 1290 0 -1 2170
box -6 -8 86 248
use AOI21X1  _1127_
timestamp 0
transform 1 0 1710 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1128_
timestamp 0
transform -1 0 1990 0 -1 2170
box -6 -8 106 248
use INVX1  _1129_
timestamp 0
transform 1 0 1610 0 1 1690
box -6 -8 66 248
use NAND3X1  _1130_
timestamp 0
transform 1 0 1510 0 1 1690
box -6 -8 106 248
use NAND3X1  _1131_
timestamp 0
transform 1 0 1090 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1132_
timestamp 0
transform 1 0 1530 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1133_
timestamp 0
transform 1 0 1810 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1134_
timestamp 0
transform 1 0 1990 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1135_
timestamp 0
transform -1 0 2190 0 -1 2170
box -6 -8 106 248
use INVX1  _1136_
timestamp 0
transform -1 0 2530 0 1 4090
box -6 -8 66 248
use NAND2X1  _1137_
timestamp 0
transform -1 0 1450 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1138_
timestamp 0
transform -1 0 1530 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1139_
timestamp 0
transform -1 0 1710 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1140_
timestamp 0
transform 1 0 690 0 -1 2170
box -6 -8 106 248
use OAI21X1  _1141_
timestamp 0
transform -1 0 890 0 -1 2170
box -6 -8 106 248
use NAND2X1  _1142_
timestamp 0
transform -1 0 810 0 -1 2650
box -6 -8 86 248
use INVX1  _1143_
timestamp 0
transform -1 0 610 0 1 4090
box -6 -8 66 248
use INVX1  _1144_
timestamp 0
transform 1 0 710 0 1 2170
box -6 -8 66 248
use AOI21X1  _1145_
timestamp 0
transform -1 0 710 0 1 2170
box -6 -8 106 248
use INVX2  _1146_
timestamp 0
transform -1 0 1410 0 -1 3130
box -6 -8 66 248
use NOR2X1  _1147_
timestamp 0
transform 1 0 1130 0 -1 3610
box -6 -8 86 248
use AND2X2  _1148_
timestamp 0
transform -1 0 1190 0 1 3130
box -6 -8 106 248
use NAND3X1  _1149_
timestamp 0
transform -1 0 1090 0 1 3130
box -6 -8 106 248
use AOI22X1  _1150_
timestamp 0
transform -1 0 910 0 1 3130
box -6 -8 126 248
use INVX1  _1151_
timestamp 0
transform 1 0 870 0 -1 3610
box -6 -8 66 248
use NAND3X1  _1152_
timestamp 0
transform -1 0 1030 0 -1 3610
box -6 -8 106 248
use NAND2X1  _1153_
timestamp 0
transform 1 0 810 0 -1 3130
box -6 -8 86 248
use NOR2X1  _1154_
timestamp 0
transform -1 0 810 0 -1 3130
box -6 -8 86 248
use OAI22X1  _1155_
timestamp 0
transform 1 0 750 0 -1 3610
box -6 -8 126 248
use NAND2X1  _1156_
timestamp 0
transform -1 0 530 0 1 3610
box -6 -8 86 248
use AND2X2  _1157_
timestamp 0
transform -1 0 230 0 -1 3130
box -6 -8 106 248
use AOI22X1  _1158_
timestamp 0
transform -1 0 130 0 -1 3130
box -6 -8 126 248
use NAND2X1  _1159_
timestamp 0
transform -1 0 90 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1160_
timestamp 0
transform -1 0 450 0 1 3130
box -6 -8 86 248
use AOI22X1  _1161_
timestamp 0
transform -1 0 370 0 1 3130
box -6 -8 126 248
use INVX1  _1162_
timestamp 0
transform -1 0 250 0 1 3610
box -6 -8 66 248
use OAI21X1  _1163_
timestamp 0
transform 1 0 90 0 1 3610
box -6 -8 106 248
use NOR2X1  _1164_
timestamp 0
transform -1 0 90 0 1 3610
box -6 -8 86 248
use OAI21X1  _1165_
timestamp 0
transform -1 0 170 0 1 2650
box -6 -8 106 248
use INVX1  _1166_
timestamp 0
transform -1 0 390 0 -1 3610
box -6 -8 66 248
use AOI21X1  _1167_
timestamp 0
transform -1 0 350 0 1 3610
box -6 -8 106 248
use NOR2X1  _1168_
timestamp 0
transform -1 0 530 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1169_
timestamp 0
transform -1 0 350 0 -1 4090
box -6 -8 106 248
use AND2X2  _1170_
timestamp 0
transform -1 0 450 0 1 3610
box -6 -8 106 248
use NAND2X1  _1171_
timestamp 0
transform -1 0 250 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1172_
timestamp 0
transform 1 0 90 0 -1 4090
box -6 -8 86 248
use NAND2X1  _1173_
timestamp 0
transform -1 0 90 0 1 4090
box -6 -8 86 248
use NAND2X1  _1174_
timestamp 0
transform -1 0 270 0 1 4090
box -6 -8 86 248
use NAND3X1  _1175_
timestamp 0
transform 1 0 210 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1176_
timestamp 0
transform 1 0 410 0 1 2170
box -6 -8 106 248
use OAI21X1  _1177_
timestamp 0
transform 1 0 510 0 1 2170
box -6 -8 106 248
use NOR2X1  _1178_
timestamp 0
transform -1 0 350 0 1 4090
box -6 -8 86 248
use AOI21X1  _1179_
timestamp 0
transform 1 0 90 0 1 4090
box -6 -8 106 248
use OAI21X1  _1180_
timestamp 0
transform -1 0 450 0 1 4090
box -6 -8 106 248
use NAND3X1  _1181_
timestamp 0
transform -1 0 410 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1182_
timestamp 0
transform -1 0 210 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1183_
timestamp 0
transform 1 0 450 0 1 4090
box -6 -8 106 248
use NAND3X1  _1184_
timestamp 0
transform 1 0 770 0 1 4090
box -6 -8 106 248
use NAND3X1  _1185_
timestamp 0
transform -1 0 810 0 -1 4570
box -6 -8 106 248
use INVX1  _1186_
timestamp 0
transform -1 0 770 0 1 4090
box -6 -8 66 248
use AOI21X1  _1187_
timestamp 0
transform -1 0 710 0 1 4090
box -6 -8 106 248
use AOI21X1  _1188_
timestamp 0
transform 1 0 410 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1189_
timestamp 0
transform 1 0 610 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1190_
timestamp 0
transform -1 0 1530 0 -1 4570
box -6 -8 86 248
use INVX1  _1191_
timestamp 0
transform -1 0 1930 0 -1 4570
box -6 -8 66 248
use NOR2X1  _1192_
timestamp 0
transform 1 0 2030 0 -1 4570
box -6 -8 86 248
use INVX1  _1193_
timestamp 0
transform 1 0 2110 0 -1 4570
box -6 -8 66 248
use OAI21X1  _1194_
timestamp 0
transform 1 0 2170 0 -1 4570
box -6 -8 106 248
use OAI22X1  _1195_
timestamp 0
transform -1 0 2390 0 -1 4570
box -6 -8 126 248
use INVX1  _1196_
timestamp 0
transform -1 0 3010 0 -1 4570
box -6 -8 66 248
use INVX8  _1197_
timestamp 0
transform 1 0 3190 0 -1 1210
box -6 -8 126 248
use INVX1  _1198_
timestamp 0
transform 1 0 1810 0 -1 4570
box -6 -8 66 248
use AOI21X1  _1199_
timestamp 0
transform 1 0 1930 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1200_
timestamp 0
transform -1 0 110 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1201_
timestamp 0
transform 1 0 510 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1202_
timestamp 0
transform 1 0 1030 0 -1 3610
box -6 -8 106 248
use INVX1  _1203_
timestamp 0
transform 1 0 1270 0 -1 4090
box -6 -8 66 248
use NAND2X1  _1204_
timestamp 0
transform 1 0 530 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1205_
timestamp 0
transform 1 0 610 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1206_
timestamp 0
transform -1 0 1170 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1207_
timestamp 0
transform 1 0 1490 0 -1 3130
box -6 -8 86 248
use INVX1  _1208_
timestamp 0
transform 1 0 2130 0 1 3130
box -6 -8 66 248
use NAND2X1  _1209_
timestamp 0
transform 1 0 1390 0 1 3130
box -6 -8 86 248
use OAI21X1  _1210_
timestamp 0
transform -1 0 1090 0 -1 3130
box -6 -8 106 248
use NAND3X1  _1211_
timestamp 0
transform 1 0 1190 0 1 3130
box -6 -8 106 248
use NAND2X1  _1212_
timestamp 0
transform 1 0 1270 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1213_
timestamp 0
transform -1 0 1270 0 -1 3130
box -6 -8 106 248
use OAI21X1  _1214_
timestamp 0
transform -1 0 990 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1215_
timestamp 0
transform 1 0 770 0 1 3610
box -6 -8 86 248
use OAI21X1  _1216_
timestamp 0
transform 1 0 670 0 1 3610
box -6 -8 106 248
use OAI21X1  _1217_
timestamp 0
transform -1 0 670 0 -1 3610
box -6 -8 106 248
use INVX1  _1218_
timestamp 0
transform 1 0 610 0 1 3610
box -6 -8 66 248
use NAND3X1  _1219_
timestamp 0
transform -1 0 950 0 1 3610
box -6 -8 106 248
use NAND3X1  _1220_
timestamp 0
transform -1 0 810 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1221_
timestamp 0
transform -1 0 90 0 -1 4090
box -6 -8 86 248
use AOI21X1  _1222_
timestamp 0
transform 1 0 350 0 -1 4090
box -6 -8 106 248
use AOI21X1  _1223_
timestamp 0
transform 1 0 950 0 1 3610
box -6 -8 106 248
use INVX1  _1224_
timestamp 0
transform -1 0 1170 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1225_
timestamp 0
transform -1 0 1010 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1226_
timestamp 0
transform 1 0 1330 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1227_
timestamp 0
transform 1 0 810 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1228_
timestamp 0
transform 1 0 1010 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1229_
timestamp 0
transform 1 0 1090 0 1 4090
box -6 -8 106 248
use AOI21X1  _1230_
timestamp 0
transform 1 0 1090 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1231_
timestamp 0
transform -1 0 1090 0 1 4090
box -6 -8 106 248
use NAND3X1  _1232_
timestamp 0
transform -1 0 1270 0 -1 4090
box -6 -8 106 248
use AOI22X1  _1233_
timestamp 0
transform -1 0 990 0 1 4090
box -6 -8 126 248
use NOR2X1  _1234_
timestamp 0
transform -1 0 1350 0 -1 4570
box -6 -8 86 248
use OR2X2  _1235_
timestamp 0
transform 1 0 2390 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1236_
timestamp 0
transform 1 0 2490 0 -1 4570
box -6 -8 106 248
use AOI22X1  _1237_
timestamp 0
transform -1 0 2710 0 -1 4570
box -6 -8 126 248
use INVX1  _1238_
timestamp 0
transform -1 0 2770 0 1 3610
box -6 -8 66 248
use NAND2X1  _1239_
timestamp 0
transform 1 0 910 0 -1 4570
box -6 -8 86 248
use NAND3X1  _1240_
timestamp 0
transform 1 0 810 0 -1 4570
box -6 -8 106 248
use NAND3X1  _1241_
timestamp 0
transform 1 0 990 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1242_
timestamp 0
transform -1 0 1270 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1243_
timestamp 0
transform 1 0 1530 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1244_
timestamp 0
transform -1 0 1450 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1245_
timestamp 0
transform -1 0 1810 0 -1 4570
box -6 -8 106 248
use NAND2X1  _1246_
timestamp 0
transform -1 0 1270 0 1 4090
box -6 -8 86 248
use OAI21X1  _1247_
timestamp 0
transform 1 0 1290 0 1 3130
box -6 -8 106 248
use INVX1  _1248_
timestamp 0
transform -1 0 1470 0 1 3610
box -6 -8 66 248
use NAND2X1  _1249_
timestamp 0
transform -1 0 610 0 1 3610
box -6 -8 86 248
use NAND2X1  _1250_
timestamp 0
transform 1 0 1410 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1251_
timestamp 0
transform 1 0 1850 0 1 3130
box -6 -8 86 248
use OAI21X1  _1252_
timestamp 0
transform 1 0 1650 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1253_
timestamp 0
transform 1 0 910 0 1 3130
box -6 -8 86 248
use OAI21X1  _1254_
timestamp 0
transform -1 0 1850 0 1 3130
box -6 -8 106 248
use OR2X2  _1255_
timestamp 0
transform -1 0 1570 0 1 3130
box -6 -8 106 248
use OAI21X1  _1256_
timestamp 0
transform 1 0 1650 0 1 3130
box -6 -8 106 248
use NAND2X1  _1257_
timestamp 0
transform -1 0 1650 0 1 3130
box -6 -8 86 248
use AOI21X1  _1258_
timestamp 0
transform 1 0 1150 0 1 3610
box -6 -8 106 248
use NAND3X1  _1259_
timestamp 0
transform 1 0 1050 0 1 3610
box -6 -8 106 248
use INVX1  _1260_
timestamp 0
transform -1 0 1630 0 1 3610
box -6 -8 66 248
use OAI21X1  _1261_
timestamp 0
transform -1 0 1570 0 1 3610
box -6 -8 106 248
use INVX1  _1262_
timestamp 0
transform 1 0 1250 0 1 3610
box -6 -8 66 248
use NAND3X1  _1263_
timestamp 0
transform -1 0 1410 0 1 3610
box -6 -8 106 248
use NAND3X1  _1264_
timestamp 0
transform -1 0 1370 0 1 4090
box -6 -8 106 248
use NAND2X1  _1265_
timestamp 0
transform 1 0 1530 0 -1 4090
box -6 -8 86 248
use NAND3X1  _1266_
timestamp 0
transform 1 0 1430 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1267_
timestamp 0
transform -1 0 1450 0 1 4090
box -6 -8 86 248
use NAND2X1  _1268_
timestamp 0
transform 1 0 2190 0 -1 4090
box -6 -8 86 248
use NAND3X1  _1269_
timestamp 0
transform 1 0 1970 0 -1 2650
box -6 -8 106 248
use NAND3X1  _1270_
timestamp 0
transform 1 0 1610 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1271_
timestamp 0
transform 1 0 1930 0 -1 3130
box -6 -8 106 248
use INVX1  _1272_
timestamp 0
transform 1 0 2130 0 -1 4090
box -6 -8 66 248
use OAI21X1  _1273_
timestamp 0
transform 1 0 2030 0 -1 4090
box -6 -8 106 248
use NAND3X1  _1274_
timestamp 0
transform 1 0 2270 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1275_
timestamp 0
transform -1 0 2710 0 1 3610
box -6 -8 106 248
use NAND2X1  _1276_
timestamp 0
transform -1 0 3330 0 1 4090
box -6 -8 86 248
use AOI21X1  _1277_
timestamp 0
transform 1 0 1630 0 1 3610
box -6 -8 106 248
use OAI21X1  _1278_
timestamp 0
transform 1 0 1930 0 1 3130
box -6 -8 106 248
use OAI21X1  _1279_
timestamp 0
transform -1 0 2130 0 1 3130
box -6 -8 106 248
use NOR2X1  _1280_
timestamp 0
transform 1 0 1850 0 -1 3130
box -6 -8 86 248
use NAND2X1  _1281_
timestamp 0
transform 1 0 2130 0 -1 3610
box -6 -8 86 248
use AND2X2  _1282_
timestamp 0
transform -1 0 2130 0 -1 3610
box -6 -8 106 248
use OR2X2  _1283_
timestamp 0
transform 1 0 1990 0 1 3610
box -6 -8 106 248
use NAND2X1  _1284_
timestamp 0
transform -1 0 2030 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1285_
timestamp 0
transform -1 0 1990 0 1 3610
box -6 -8 86 248
use NOR2X1  _1286_
timestamp 0
transform 1 0 1730 0 1 3610
box -6 -8 86 248
use AND2X2  _1287_
timestamp 0
transform -1 0 1790 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1288_
timestamp 0
transform -1 0 1710 0 1 4090
box -6 -8 86 248
use INVX1  _1289_
timestamp 0
transform 1 0 1890 0 1 4090
box -6 -8 66 248
use NAND3X1  _1290_
timestamp 0
transform 1 0 1950 0 1 4090
box -6 -8 106 248
use OAI21X1  _1291_
timestamp 0
transform 1 0 1710 0 1 4090
box -6 -8 106 248
use NAND2X1  _1292_
timestamp 0
transform -1 0 1890 0 1 4090
box -6 -8 86 248
use NAND3X1  _1293_
timestamp 0
transform 1 0 2050 0 1 4090
box -6 -8 106 248
use NAND2X1  _1294_
timestamp 0
transform -1 0 3250 0 1 4090
box -6 -8 86 248
use INVX1  _1295_
timestamp 0
transform -1 0 3570 0 1 1210
box -6 -8 66 248
use NAND3X1  _1296_
timestamp 0
transform 1 0 1450 0 1 4090
box -6 -8 106 248
use NOR2X1  _1297_
timestamp 0
transform 1 0 1890 0 -1 4090
box -6 -8 86 248
use INVX1  _1298_
timestamp 0
transform -1 0 2030 0 -1 4090
box -6 -8 66 248
use NOR2X1  _1299_
timestamp 0
transform -1 0 1630 0 1 4090
box -6 -8 86 248
use NOR2X1  _1300_
timestamp 0
transform -1 0 1690 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1301_
timestamp 0
transform -1 0 1890 0 -1 4090
box -6 -8 106 248
use AOI21X1  _1302_
timestamp 0
transform -1 0 1910 0 1 3610
box -6 -8 106 248
use INVX1  _1303_
timestamp 0
transform 1 0 2310 0 -1 3610
box -6 -8 66 248
use NAND3X1  _1304_
timestamp 0
transform 1 0 2210 0 -1 3610
box -6 -8 106 248
use INVX1  _1305_
timestamp 0
transform 1 0 2030 0 -1 3130
box -6 -8 66 248
use OAI21X1  _1306_
timestamp 0
transform 1 0 2190 0 1 3130
box -6 -8 106 248
use NAND2X1  _1307_
timestamp 0
transform 1 0 2350 0 1 3130
box -6 -8 86 248
use NAND2X1  _1308_
timestamp 0
transform -1 0 2490 0 1 1210
box -6 -8 86 248
use INVX1  _1309_
timestamp 0
transform 1 0 2490 0 1 1210
box -6 -8 66 248
use OAI21X1  _1310_
timestamp 0
transform 1 0 2630 0 1 1210
box -6 -8 106 248
use OAI22X1  _1311_
timestamp 0
transform -1 0 2850 0 1 1210
box -6 -8 126 248
use INVX1  _1312_
timestamp 0
transform 1 0 4310 0 -1 2170
box -6 -8 66 248
use OR2X2  _1313_
timestamp 0
transform 1 0 2570 0 -1 2170
box -6 -8 106 248
use INVX1  _1314_
timestamp 0
transform -1 0 2350 0 1 3130
box -6 -8 66 248
use OAI21X1  _1315_
timestamp 0
transform 1 0 2090 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1316_
timestamp 0
transform 1 0 2190 0 -1 3130
box -6 -8 86 248
use AOI22X1  _1317_
timestamp 0
transform -1 0 3370 0 -1 2170
box -6 -8 126 248
use NOR2X1  _1318_
timestamp 0
transform 1 0 4470 0 -1 250
box -6 -8 86 248
use INVX1  _1319_
timestamp 0
transform -1 0 4470 0 -1 250
box -6 -8 66 248
use NAND2X1  _1320_
timestamp 0
transform 1 0 4550 0 -1 250
box -6 -8 86 248
use NAND2X1  _1321_
timestamp 0
transform 1 0 4690 0 -1 250
box -6 -8 86 248
use NAND2X1  _1322_
timestamp 0
transform 1 0 4330 0 -1 730
box -6 -8 86 248
use OAI21X1  _1323_
timestamp 0
transform -1 0 4510 0 -1 730
box -6 -8 106 248
use NOR2X1  _1324_
timestamp 0
transform 1 0 3990 0 -1 250
box -6 -8 86 248
use NOR2X1  _1325_
timestamp 0
transform 1 0 4070 0 -1 250
box -6 -8 86 248
use NOR2X1  _1326_
timestamp 0
transform -1 0 4230 0 -1 250
box -6 -8 86 248
use NAND2X1  _1327_
timestamp 0
transform -1 0 4410 0 -1 250
box -6 -8 86 248
use OAI21X1  _1328_
timestamp 0
transform 1 0 4230 0 -1 250
box -6 -8 106 248
use NAND2X1  _1329_
timestamp 0
transform -1 0 4370 0 1 250
box -6 -8 86 248
use NAND2X1  _1330_
timestamp 0
transform 1 0 3950 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1331_
timestamp 0
transform -1 0 4050 0 1 730
box -6 -8 106 248
use OAI21X1  _1332_
timestamp 0
transform 1 0 3890 0 -1 250
box -6 -8 106 248
use NOR2X1  _1333_
timestamp 0
transform -1 0 3590 0 -1 250
box -6 -8 86 248
use NOR2X1  _1334_
timestamp 0
transform -1 0 3230 0 1 250
box -6 -8 86 248
use NOR2X1  _1335_
timestamp 0
transform -1 0 3570 0 1 250
box -6 -8 86 248
use NAND2X1  _1336_
timestamp 0
transform 1 0 3670 0 1 250
box -6 -8 86 248
use OR2X2  _1337_
timestamp 0
transform 1 0 3570 0 1 250
box -6 -8 106 248
use NAND2X1  _1338_
timestamp 0
transform 1 0 3750 0 1 250
box -6 -8 86 248
use NAND2X1  _1339_
timestamp 0
transform -1 0 4010 0 -1 730
box -6 -8 86 248
use OAI21X1  _1340_
timestamp 0
transform 1 0 3830 0 -1 730
box -6 -8 106 248
use AOI21X1  _1341_
timestamp 0
transform -1 0 3490 0 1 250
box -6 -8 106 248
use NOR2X1  _1342_
timestamp 0
transform -1 0 3070 0 1 730
box -6 -8 86 248
use NOR2X1  _1343_
timestamp 0
transform -1 0 3150 0 1 730
box -6 -8 86 248
use OAI21X1  _1344_
timestamp 0
transform 1 0 3210 0 1 730
box -6 -8 106 248
use INVX1  _1345_
timestamp 0
transform -1 0 3410 0 -1 730
box -6 -8 66 248
use INVX1  _1346_
timestamp 0
transform 1 0 3190 0 -1 730
box -6 -8 66 248
use INVX1  _1347_
timestamp 0
transform 1 0 3130 0 -1 730
box -6 -8 66 248
use NAND3X1  _1348_
timestamp 0
transform 1 0 3250 0 -1 730
box -6 -8 106 248
use NAND2X1  _1349_
timestamp 0
transform 1 0 3310 0 1 730
box -6 -8 86 248
use NAND2X1  _1350_
timestamp 0
transform 1 0 3410 0 1 1690
box -6 -8 86 248
use OAI21X1  _1351_
timestamp 0
transform 1 0 3310 0 1 1690
box -6 -8 106 248
use NAND2X1  _1352_
timestamp 0
transform -1 0 3830 0 1 2170
box -6 -8 86 248
use NOR2X1  _1353_
timestamp 0
transform -1 0 3070 0 1 1690
box -6 -8 86 248
use NOR2X1  _1354_
timestamp 0
transform -1 0 2970 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1355_
timestamp 0
transform 1 0 3030 0 -1 730
box -6 -8 106 248
use INVX1  _1356_
timestamp 0
transform 1 0 2930 0 1 1690
box -6 -8 66 248
use OAI21X1  _1357_
timestamp 0
transform 1 0 2830 0 1 1690
box -6 -8 106 248
use NOR2X1  _1358_
timestamp 0
transform -1 0 2830 0 1 1690
box -6 -8 86 248
use NAND2X1  _1359_
timestamp 0
transform -1 0 2750 0 -1 2170
box -6 -8 86 248
use NAND2X1  _1360_
timestamp 0
transform 1 0 2750 0 -1 2170
box -6 -8 86 248
use OAI21X1  _1361_
timestamp 0
transform 1 0 3610 0 -1 2170
box -6 -8 106 248
use INVX1  _1362_
timestamp 0
transform 1 0 3690 0 -1 1690
box -6 -8 66 248
use AOI21X1  _1363_
timestamp 0
transform 1 0 2790 0 -1 1690
box -6 -8 106 248
use NOR2X1  _1364_
timestamp 0
transform -1 0 2250 0 1 1690
box -6 -8 86 248
use NOR2X1  _1365_
timestamp 0
transform 1 0 2490 0 1 1690
box -6 -8 86 248
use NOR2X1  _1366_
timestamp 0
transform 1 0 2410 0 1 1690
box -6 -8 86 248
use AND2X2  _1367_
timestamp 0
transform -1 0 2710 0 -1 1690
box -6 -8 106 248
use NOR2X1  _1368_
timestamp 0
transform 1 0 2710 0 -1 1690
box -6 -8 86 248
use OAI21X1  _1369_
timestamp 0
transform -1 0 2610 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1370_
timestamp 0
transform -1 0 3450 0 -1 1690
box -6 -8 106 248
use NAND2X1  _1371_
timestamp 0
transform 1 0 2810 0 1 2650
box -6 -8 86 248
use NAND2X1  _1372_
timestamp 0
transform -1 0 2750 0 1 1690
box -6 -8 86 248
use OAI21X1  _1373_
timestamp 0
transform 1 0 2570 0 1 1690
box -6 -8 106 248
use AND2X2  _1374_
timestamp 0
transform -1 0 2570 0 -1 2170
box -6 -8 106 248
use AOI21X1  _1375_
timestamp 0
transform -1 0 2490 0 1 2170
box -6 -8 106 248
use NOR2X1  _1376_
timestamp 0
transform -1 0 2150 0 1 2650
box -6 -8 86 248
use NOR2X1  _1377_
timestamp 0
transform -1 0 2230 0 1 2650
box -6 -8 86 248
use NOR2X1  _1378_
timestamp 0
transform -1 0 2310 0 1 2650
box -6 -8 86 248
use INVX1  _1379_
timestamp 0
transform 1 0 2450 0 1 2650
box -6 -8 66 248
use AND2X2  _1380_
timestamp 0
transform 1 0 2510 0 1 2650
box -6 -8 106 248
use OAI21X1  _1381_
timestamp 0
transform 1 0 2610 0 1 2650
box -6 -8 106 248
use OAI21X1  _1382_
timestamp 0
transform 1 0 2710 0 1 2650
box -6 -8 106 248
use INVX1  _1383_
timestamp 0
transform 1 0 2310 0 1 2650
box -6 -8 66 248
use OAI21X1  _1384_
timestamp 0
transform 1 0 2630 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1385_
timestamp 0
transform -1 0 2450 0 1 2650
box -6 -8 86 248
use NOR2X1  _1386_
timestamp 0
transform -1 0 2290 0 -1 2650
box -6 -8 86 248
use NOR2X1  _1387_
timestamp 0
transform 1 0 2450 0 -1 2650
box -6 -8 86 248
use OR2X2  _1388_
timestamp 0
transform 1 0 2810 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1389_
timestamp 0
transform -1 0 2810 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1390_
timestamp 0
transform 1 0 2910 0 -1 2650
box -6 -8 86 248
use NAND2X1  _1391_
timestamp 0
transform -1 0 3330 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1392_
timestamp 0
transform 1 0 3070 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1393_
timestamp 0
transform 1 0 3730 0 1 3130
box -6 -8 86 248
use INVX1  _1394_
timestamp 0
transform -1 0 2350 0 -1 2650
box -6 -8 66 248
use OAI21X1  _1395_
timestamp 0
transform -1 0 2450 0 -1 2650
box -6 -8 106 248
use AND2X2  _1396_
timestamp 0
transform 1 0 2530 0 -1 2650
box -6 -8 106 248
use AOI21X1  _1397_
timestamp 0
transform -1 0 2390 0 1 2170
box -6 -8 106 248
use NAND3X1  _1398_
timestamp 0
transform 1 0 2490 0 1 2170
box -6 -8 106 248
use AND2X2  _1399_
timestamp 0
transform 1 0 2590 0 1 2170
box -6 -8 106 248
use INVX1  _1400_
timestamp 0
transform 1 0 3410 0 -1 3610
box -6 -8 66 248
use NOR2X1  _1401_
timestamp 0
transform -1 0 2610 0 1 4090
box -6 -8 86 248
use NOR2X1  _1402_
timestamp 0
transform -1 0 2990 0 1 4090
box -6 -8 86 248
use NOR2X1  _1403_
timestamp 0
transform 1 0 3050 0 -1 4090
box -6 -8 86 248
use NOR2X1  _1404_
timestamp 0
transform 1 0 3330 0 -1 3610
box -6 -8 86 248
use INVX1  _1405_
timestamp 0
transform -1 0 3330 0 -1 3610
box -6 -8 66 248
use OAI21X1  _1406_
timestamp 0
transform -1 0 3270 0 -1 3610
box -6 -8 106 248
use OAI21X1  _1407_
timestamp 0
transform 1 0 3390 0 1 3130
box -6 -8 106 248
use AOI21X1  _1408_
timestamp 0
transform -1 0 3310 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1409_
timestamp 0
transform -1 0 3190 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1410_
timestamp 0
transform -1 0 3370 0 -1 4570
box -6 -8 86 248
use NOR2X1  _1411_
timestamp 0
transform 1 0 3330 0 1 4090
box -6 -8 86 248
use AND2X2  _1412_
timestamp 0
transform 1 0 4050 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1413_
timestamp 0
transform -1 0 4050 0 -1 4090
box -6 -8 86 248
use OAI21X1  _1414_
timestamp 0
transform 1 0 4150 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1415_
timestamp 0
transform -1 0 4350 0 -1 4090
box -6 -8 106 248
use NAND2X1  _1416_
timestamp 0
transform -1 0 3950 0 -1 3610
box -6 -8 86 248
use AND2X2  _1417_
timestamp 0
transform 1 0 3310 0 -1 4090
box -6 -8 106 248
use OAI21X1  _1418_
timestamp 0
transform -1 0 3110 0 -1 4570
box -6 -8 106 248
use OAI21X1  _1419_
timestamp 0
transform -1 0 3290 0 -1 4570
box -6 -8 106 248
use AOI21X1  _1420_
timestamp 0
transform -1 0 3330 0 1 3610
box -6 -8 106 248
use NOR2X1  _1421_
timestamp 0
transform -1 0 2850 0 1 3610
box -6 -8 86 248
use NOR2X1  _1422_
timestamp 0
transform -1 0 2930 0 1 3610
box -6 -8 86 248
use NOR2X1  _1423_
timestamp 0
transform -1 0 3010 0 1 3610
box -6 -8 86 248
use INVX1  _1424_
timestamp 0
transform 1 0 3010 0 1 3610
box -6 -8 66 248
use AND2X2  _1425_
timestamp 0
transform 1 0 3490 0 1 3610
box -6 -8 106 248
use OAI21X1  _1426_
timestamp 0
transform 1 0 3590 0 1 3610
box -6 -8 106 248
use OAI21X1  _1427_
timestamp 0
transform 1 0 3690 0 1 3610
box -6 -8 106 248
use INVX1  _1428_
timestamp 0
transform -1 0 3130 0 1 3610
box -6 -8 66 248
use OAI21X1  _1429_
timestamp 0
transform 1 0 3130 0 1 3610
box -6 -8 106 248
use NOR2X1  _1430_
timestamp 0
transform 1 0 3730 0 1 4090
box -6 -8 86 248
use NAND2X1  _1431_
timestamp 0
transform -1 0 3730 0 1 4090
box -6 -8 86 248
use INVX1  _1432_
timestamp 0
transform -1 0 3550 0 -1 4090
box -6 -8 66 248
use NOR2X1  _1433_
timestamp 0
transform -1 0 3490 0 -1 4090
box -6 -8 86 248
use INVX1  _1434_
timestamp 0
transform 1 0 3430 0 1 3610
box -6 -8 66 248
use OR2X2  _1435_
timestamp 0
transform 1 0 3650 0 -1 3610
box -6 -8 106 248
use AOI21X1  _1436_
timestamp 0
transform 1 0 3550 0 -1 3610
box -6 -8 106 248
use AOI22X1  _1437_
timestamp 0
transform -1 0 3870 0 -1 3610
box -6 -8 126 248
use NAND2X1  _1438_
timestamp 0
transform -1 0 3890 0 1 1690
box -6 -8 86 248
use AOI21X1  _1439_
timestamp 0
transform 1 0 3330 0 1 3610
box -6 -8 106 248
use NOR2X1  _1440_
timestamp 0
transform -1 0 3550 0 -1 3610
box -6 -8 86 248
use NAND2X1  _1441_
timestamp 0
transform 1 0 3570 0 1 3130
box -6 -8 86 248
use NAND2X1  _1442_
timestamp 0
transform 1 0 3650 0 1 3130
box -6 -8 86 248
use NAND2X1  _1443_
timestamp 0
transform 1 0 3490 0 1 3130
box -6 -8 86 248
use NOR2X1  _1444_
timestamp 0
transform -1 0 3510 0 1 2650
box -6 -8 86 248
use OR2X2  _1445_
timestamp 0
transform 1 0 3650 0 1 2170
box -6 -8 106 248
use NOR2X1  _1446_
timestamp 0
transform -1 0 3730 0 1 1210
box -6 -8 86 248
use NOR2X1  _1447_
timestamp 0
transform -1 0 3650 0 1 1210
box -6 -8 86 248
use NOR2X1  _1448_
timestamp 0
transform 1 0 3910 0 -1 1690
box -6 -8 86 248
use NOR2X1  _1449_
timestamp 0
transform 1 0 3990 0 -1 1690
box -6 -8 86 248
use NOR2X1  _1450_
timestamp 0
transform -1 0 3650 0 1 2170
box -6 -8 86 248
use INVX1  _1451_
timestamp 0
transform 1 0 4070 0 -1 1690
box -6 -8 66 248
use OAI21X1  _1452_
timestamp 0
transform -1 0 4090 0 1 1690
box -6 -8 106 248
use OAI21X1  _1453_
timestamp 0
transform -1 0 3990 0 1 1690
box -6 -8 106 248
use INVX1  _1454_
timestamp 0
transform -1 0 4350 0 1 3130
box -6 -8 66 248
use INVX1  _1455_
timestamp 0
transform -1 0 3810 0 -1 1690
box -6 -8 66 248
use OAI21X1  _1456_
timestamp 0
transform -1 0 3910 0 -1 1690
box -6 -8 106 248
use NOR2X1  _1457_
timestamp 0
transform -1 0 4530 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1458_
timestamp 0
transform -1 0 4450 0 -1 2170
box -6 -8 86 248
use NOR2X1  _1459_
timestamp 0
transform -1 0 4430 0 1 1690
box -6 -8 86 248
use INVX1  _1460_
timestamp 0
transform -1 0 4250 0 1 1690
box -6 -8 66 248
use OR2X2  _1461_
timestamp 0
transform 1 0 4090 0 1 1690
box -6 -8 106 248
use AOI21X1  _1462_
timestamp 0
transform 1 0 4130 0 -1 1690
box -6 -8 106 248
use AOI22X1  _1463_
timestamp 0
transform -1 0 4310 0 -1 2170
box -6 -8 126 248
use NAND2X1  _1464_
timestamp 0
transform -1 0 4370 0 1 1210
box -6 -8 86 248
use AOI21X1  _1465_
timestamp 0
transform 1 0 4250 0 1 1690
box -6 -8 106 248
use NOR2X1  _1466_
timestamp 0
transform 1 0 4230 0 -1 1690
box -6 -8 86 248
use INVX1  _1467_
timestamp 0
transform 1 0 4470 0 -1 1690
box -6 -8 66 248
use OAI21X1  _1468_
timestamp 0
transform 1 0 4590 0 -1 1690
box -6 -8 106 248
use NOR2X1  _1469_
timestamp 0
transform 1 0 4570 0 1 1210
box -6 -8 86 248
use INVX1  _1470_
timestamp 0
transform 1 0 4410 0 -1 1690
box -6 -8 66 248
use AOI21X1  _1471_
timestamp 0
transform 1 0 4310 0 -1 1690
box -6 -8 106 248
use OAI21X1  _1472_
timestamp 0
transform -1 0 4570 0 1 1210
box -6 -8 106 248
use OAI21X1  _1473_
timestamp 0
transform -1 0 4470 0 1 1210
box -6 -8 106 248
use NAND2X1  _1474_
timestamp 0
transform 1 0 4270 0 -1 1210
box -6 -8 86 248
use NAND3X1  _1475_
timestamp 0
transform 1 0 4630 0 -1 1210
box -6 -8 106 248
use OAI21X1  _1476_
timestamp 0
transform 1 0 4530 0 -1 1210
box -6 -8 106 248
use NAND2X1  _1477_
timestamp 0
transform -1 0 4530 0 -1 1210
box -6 -8 86 248
use OAI21X1  _1478_
timestamp 0
transform 1 0 4350 0 -1 1210
box -6 -8 106 248
use INVX1  _1479_
timestamp 0
transform 1 0 4650 0 -1 4090
box -6 -8 66 248
use NAND3X1  _1480_
timestamp 0
transform 1 0 4290 0 -1 3130
box -6 -8 106 248
use NAND2X1  _1481_
timestamp 0
transform 1 0 4650 0 1 2170
box -6 -8 86 248
use OAI21X1  _1482_
timestamp 0
transform 1 0 4550 0 1 2170
box -6 -8 106 248
use INVX1  _1483_
timestamp 0
transform 1 0 4670 0 1 3610
box -6 -8 66 248
use NAND2X1  _1484_
timestamp 0
transform 1 0 4630 0 1 2650
box -6 -8 86 248
use OAI21X1  _1485_
timestamp 0
transform 1 0 4530 0 1 2650
box -6 -8 106 248
use INVX1  _1486_
timestamp 0
transform -1 0 4670 0 1 3610
box -6 -8 66 248
use NAND2X1  _1487_
timestamp 0
transform 1 0 4690 0 -1 4570
box -6 -8 86 248
use OAI21X1  _1488_
timestamp 0
transform 1 0 4630 0 -1 3130
box -6 -8 106 248
use INVX1  _1489_
timestamp 0
transform -1 0 4770 0 1 1210
box -6 -8 66 248
use NAND2X1  _1490_
timestamp 0
transform 1 0 4570 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1491_
timestamp 0
transform 1 0 4470 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1492_
timestamp 0
transform -1 0 4050 0 1 3130
box -6 -8 86 248
use NOR2X1  _1493_
timestamp 0
transform -1 0 4390 0 1 4090
box -6 -8 86 248
use AOI21X1  _1494_
timestamp 0
transform -1 0 4490 0 1 4090
box -6 -8 106 248
use NOR2X1  _1495_
timestamp 0
transform 1 0 4050 0 1 4090
box -6 -8 86 248
use AOI21X1  _1496_
timestamp 0
transform -1 0 4230 0 1 4090
box -6 -8 106 248
use NOR2X1  _1497_
timestamp 0
transform 1 0 3890 0 -1 4090
box -6 -8 86 248
use AOI21X1  _1498_
timestamp 0
transform -1 0 3890 0 -1 4090
box -6 -8 106 248
use NOR2X1  _1499_
timestamp 0
transform -1 0 4190 0 1 3610
box -6 -8 86 248
use AOI21X1  _1500_
timestamp 0
transform 1 0 4190 0 1 3610
box -6 -8 106 248
use INVX1  _1501_
timestamp 0
transform -1 0 3430 0 1 2650
box -6 -8 66 248
use OAI21X1  _1502_
timestamp 0
transform 1 0 3130 0 1 2170
box -6 -8 106 248
use OAI21X1  _1503_
timestamp 0
transform -1 0 3570 0 1 2170
box -6 -8 106 248
use OAI21X1  _1504_
timestamp 0
transform -1 0 3030 0 1 2170
box -6 -8 106 248
use OAI21X1  _1505_
timestamp 0
transform -1 0 3130 0 1 2170
box -6 -8 106 248
use OAI21X1  _1506_
timestamp 0
transform 1 0 3190 0 1 3130
box -6 -8 106 248
use OAI21X1  _1507_
timestamp 0
transform -1 0 3390 0 1 3130
box -6 -8 106 248
use OAI21X1  _1508_
timestamp 0
transform -1 0 3090 0 1 3130
box -6 -8 106 248
use OAI21X1  _1509_
timestamp 0
transform -1 0 3190 0 1 3130
box -6 -8 106 248
use NOR2X1  _1510_
timestamp 0
transform 1 0 3950 0 -1 2650
box -6 -8 86 248
use AOI21X1  _1511_
timestamp 0
transform -1 0 3950 0 -1 2650
box -6 -8 106 248
use NOR2X1  _1512_
timestamp 0
transform 1 0 3170 0 -1 2170
box -6 -8 86 248
use AOI21X1  _1513_
timestamp 0
transform -1 0 3170 0 -1 2170
box -6 -8 106 248
use NOR2X1  _1514_
timestamp 0
transform 1 0 3190 0 -1 3130
box -6 -8 86 248
use AOI21X1  _1515_
timestamp 0
transform -1 0 3190 0 -1 3130
box -6 -8 106 248
use NOR2X1  _1516_
timestamp 0
transform -1 0 3170 0 1 1210
box -6 -8 86 248
use AOI21X1  _1517_
timestamp 0
transform -1 0 3270 0 1 1210
box -6 -8 106 248
use NAND2X1  _1518_
timestamp 0
transform -1 0 1570 0 -1 2650
box -6 -8 86 248
use OAI21X1  _1519_
timestamp 0
transform -1 0 1590 0 1 2170
box -6 -8 106 248
use NAND2X1  _1520_
timestamp 0
transform -1 0 730 0 -1 3130
box -6 -8 86 248
use OAI21X1  _1521_
timestamp 0
transform -1 0 1350 0 -1 2650
box -6 -8 106 248
use NAND2X1  _1522_
timestamp 0
transform 1 0 1210 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1523_
timestamp 0
transform -1 0 1250 0 1 2170
box -6 -8 106 248
use NAND2X1  _1524_
timestamp 0
transform -1 0 470 0 -1 3610
box -6 -8 86 248
use OAI21X1  _1525_
timestamp 0
transform -1 0 570 0 -1 3610
box -6 -8 106 248
use DFFPOSX1  _1526_
timestamp 0
transform -1 0 1470 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1527_
timestamp 0
transform -1 0 470 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1528_
timestamp 0
transform 1 0 1470 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1529_
timestamp 0
transform -1 0 690 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1530_
timestamp 0
transform -1 0 4770 0 1 250
box -6 -8 246 248
use DFFPOSX1  _1531_
timestamp 0
transform 1 0 3590 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1532_
timestamp 0
transform -1 0 3830 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _1533_
timestamp 0
transform -1 0 3630 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1534_
timestamp 0
transform -1 0 3310 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1535_
timestamp 0
transform -1 0 2510 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _1536_
timestamp 0
transform -1 0 2670 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1537_
timestamp 0
transform -1 0 2670 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1538_
timestamp 0
transform -1 0 2850 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1539_
timestamp 0
transform -1 0 3670 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1540_
timestamp 0
transform 1 0 2650 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1541_
timestamp 0
transform -1 0 4610 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1542_
timestamp 0
transform -1 0 4030 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1543_
timestamp 0
transform -1 0 4770 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _1544_
timestamp 0
transform 1 0 4290 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1545_
timestamp 0
transform 1 0 4510 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1546_
timestamp 0
transform 1 0 2910 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _1547_
timestamp 0
transform -1 0 4290 0 1 250
box -6 -8 246 248
use DFFPOSX1  _1548_
timestamp 0
transform 1 0 3270 0 -1 250
box -6 -8 246 248
use DFFPOSX1  _1549_
timestamp 0
transform 1 0 2790 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1550_
timestamp 0
transform 1 0 2770 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1551_
timestamp 0
transform 1 0 1930 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1552_
timestamp 0
transform 1 0 1550 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1553_
timestamp 0
transform 1 0 2050 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1554_
timestamp 0
transform 1 0 2150 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1555_
timestamp 0
transform 1 0 2710 0 -1 4570
box -6 -8 246 248
use DFFPOSX1  _1556_
timestamp 0
transform 1 0 2370 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1557_
timestamp 0
transform 1 0 3410 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1558_
timestamp 0
transform 1 0 3270 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1559_
timestamp 0
transform 1 0 3370 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _1560_
timestamp 0
transform -1 0 4290 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1561_
timestamp 0
transform 1 0 3710 0 1 730
box -6 -8 246 248
use DFFPOSX1  _1562_
timestamp 0
transform -1 0 4250 0 -1 730
box -6 -8 246 248
use DFFPOSX1  _1563_
timestamp 0
transform -1 0 3730 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1564_
timestamp 0
transform 1 0 3710 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _1565_
timestamp 0
transform 1 0 3450 0 -1 1690
box -6 -8 246 248
use DFFPOSX1  _1566_
timestamp 0
transform 1 0 2890 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1567_
timestamp 0
transform 1 0 3130 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1568_
timestamp 0
transform 1 0 3270 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1569_
timestamp 0
transform -1 0 4650 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1570_
timestamp 0
transform 1 0 3790 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1571_
timestamp 0
transform -1 0 4190 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1572_
timestamp 0
transform -1 0 4190 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _1573_
timestamp 0
transform 1 0 4070 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1574_
timestamp 0
transform -1 0 4670 0 1 1690
box -6 -8 246 248
use DFFPOSX1  _1575_
timestamp 0
transform -1 0 4270 0 -1 1210
box -6 -8 246 248
use DFFPOSX1  _1576_
timestamp 0
transform -1 0 4550 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1577_
timestamp 0
transform 1 0 4290 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1578_
timestamp 0
transform 1 0 4530 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1579_
timestamp 0
transform 1 0 4230 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1580_
timestamp 0
transform -1 0 4730 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1581_
timestamp 0
transform -1 0 4050 0 1 4090
box -6 -8 246 248
use DFFPOSX1  _1582_
timestamp 0
transform -1 0 3790 0 -1 4090
box -6 -8 246 248
use DFFPOSX1  _1583_
timestamp 0
transform -1 0 4530 0 1 3610
box -6 -8 246 248
use DFFPOSX1  _1584_
timestamp 0
transform -1 0 3470 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1585_
timestamp 0
transform -1 0 2930 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1586_
timestamp 0
transform -1 0 2990 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1587_
timestamp 0
transform -1 0 3170 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1588_
timestamp 0
transform 1 0 3610 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1589_
timestamp 0
transform 1 0 2830 0 -1 2170
box -6 -8 246 248
use DFFPOSX1  _1590_
timestamp 0
transform 1 0 2770 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1591_
timestamp 0
transform 1 0 2850 0 1 1210
box -6 -8 246 248
use DFFPOSX1  _1592_
timestamp 0
transform 1 0 1590 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1593_
timestamp 0
transform 1 0 1570 0 -1 2650
box -6 -8 246 248
use DFFPOSX1  _1594_
timestamp 0
transform 1 0 1250 0 1 2170
box -6 -8 246 248
use DFFPOSX1  _1595_
timestamp 0
transform 1 0 90 0 -1 3610
box -6 -8 246 248
use DFFPOSX1  _1596_
timestamp 0
transform 1 0 10 0 1 3130
box -6 -8 246 248
use DFFPOSX1  _1597_
timestamp 0
transform 1 0 3510 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1598_
timestamp 0
transform 1 0 3570 0 1 2650
box -6 -8 246 248
use DFFPOSX1  _1599_
timestamp 0
transform -1 0 4630 0 -1 3130
box -6 -8 246 248
use DFFPOSX1  _1600_
timestamp 0
transform -1 0 4430 0 -1 3610
box -6 -8 246 248
use BUFX2  _1601_
timestamp 0
transform -1 0 4130 0 -1 4570
box -6 -8 86 248
use BUFX2  _1602_
timestamp 0
transform 1 0 3810 0 1 3130
box -6 -8 86 248
use BUFX2  _1603_
timestamp 0
transform 1 0 2370 0 -1 4090
box -6 -8 86 248
use BUFX2  _1604_
timestamp 0
transform 1 0 2390 0 1 4090
box -6 -8 86 248
use BUFX2  _1605_
timestamp 0
transform 1 0 2090 0 1 3610
box -6 -8 86 248
use BUFX2  _1606_
timestamp 0
transform 1 0 4050 0 1 3130
box -6 -8 86 248
use BUFX2  _1607_
timestamp 0
transform 1 0 4230 0 1 4090
box -6 -8 86 248
use BUFX2  _1608_
timestamp 0
transform 1 0 4530 0 1 3610
box -6 -8 86 248
use BUFX2  _1609_
timestamp 0
transform 1 0 4610 0 -1 4570
box -6 -8 86 248
use BUFX2  BUFX2_insert0
timestamp 0
transform 1 0 2690 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert1
timestamp 0
transform 1 0 2610 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert2
timestamp 0
transform -1 0 3390 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert3
timestamp 0
transform 1 0 2770 0 -1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert4
timestamp 0
transform 1 0 3390 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert5
timestamp 0
transform 1 0 4030 0 1 3610
box -6 -8 86 248
use BUFX2  BUFX2_insert6
timestamp 0
transform -1 0 4290 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert7
timestamp 0
transform -1 0 2630 0 1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert16
timestamp 0
transform 1 0 3730 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert17
timestamp 0
transform -1 0 3610 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert18
timestamp 0
transform 1 0 3630 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert19
timestamp 0
transform -1 0 3250 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert20
timestamp 0
transform 1 0 3870 0 -1 1210
box -6 -8 86 248
use BUFX2  BUFX2_insert21
timestamp 0
transform -1 0 530 0 -1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert22
timestamp 0
transform -1 0 490 0 1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert23
timestamp 0
transform 1 0 2090 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert24
timestamp 0
transform -1 0 810 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert25
timestamp 0
transform 1 0 1570 0 -1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert26
timestamp 0
transform 1 0 2670 0 1 3130
box -6 -8 86 248
use BUFX2  BUFX2_insert27
timestamp 0
transform 1 0 2990 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert28
timestamp 0
transform 1 0 3450 0 -1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert29
timestamp 0
transform -1 0 1550 0 1 2650
box -6 -8 86 248
use BUFX2  BUFX2_insert30
timestamp 0
transform 1 0 1910 0 -1 250
box -6 -8 86 248
use BUFX2  BUFX2_insert31
timestamp 0
transform 1 0 690 0 1 1690
box -6 -8 86 248
use BUFX2  BUFX2_insert32
timestamp 0
transform -1 0 630 0 -1 730
box -6 -8 86 248
use BUFX2  BUFX2_insert33
timestamp 0
transform -1 0 90 0 -1 2170
box -6 -8 86 248
use CLKBUF1  CLKBUF1_insert8
timestamp 0
transform -1 0 2370 0 1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert9
timestamp 0
transform -1 0 4630 0 -1 3610
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert10
timestamp 0
transform -1 0 4050 0 -1 4570
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert11
timestamp 0
transform -1 0 2390 0 -1 2170
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert12
timestamp 0
transform 1 0 2450 0 -1 4090
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert13
timestamp 0
transform 1 0 3670 0 -1 1210
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert14
timestamp 0
transform 1 0 4030 0 -1 2650
box -6 -8 206 248
use CLKBUF1  CLKBUF1_insert15
timestamp 0
transform 1 0 3470 0 -1 1210
box -6 -8 206 248
use FILL  FILL70650x39750
timestamp 0
transform 1 0 4710 0 1 2650
box -6 -8 26 248
use FILL  FILL70650x57750
timestamp 0
transform -1 0 4730 0 -1 4090
box -6 -8 26 248
use FILL  FILL70950x10950
timestamp 0
transform 1 0 4730 0 1 730
box -6 -8 26 248
use FILL  FILL70950x14550
timestamp 0
transform -1 0 4750 0 -1 1210
box -6 -8 26 248
use FILL  FILL70950x32550
timestamp 0
transform 1 0 4730 0 1 2170
box -6 -8 26 248
use FILL  FILL70950x36150
timestamp 0
transform -1 0 4750 0 -1 2650
box -6 -8 26 248
use FILL  FILL70950x39750
timestamp 0
transform 1 0 4730 0 1 2650
box -6 -8 26 248
use FILL  FILL70950x43350
timestamp 0
transform -1 0 4750 0 -1 3130
box -6 -8 26 248
use FILL  FILL70950x50550
timestamp 0
transform -1 0 4750 0 -1 3610
box -6 -8 26 248
use FILL  FILL70950x54150
timestamp 0
transform 1 0 4730 0 1 3610
box -6 -8 26 248
use FILL  FILL70950x57750
timestamp 0
transform -1 0 4750 0 -1 4090
box -6 -8 26 248
use FILL  FILL70950x61350
timestamp 0
transform 1 0 4730 0 1 4090
box -6 -8 26 248
use FILL  FILL71250x7350
timestamp 0
transform -1 0 4770 0 -1 730
box -6 -8 26 248
use FILL  FILL71250x10950
timestamp 0
transform 1 0 4750 0 1 730
box -6 -8 26 248
use FILL  FILL71250x14550
timestamp 0
transform -1 0 4770 0 -1 1210
box -6 -8 26 248
use FILL  FILL71250x25350
timestamp 0
transform 1 0 4750 0 1 1690
box -6 -8 26 248
use FILL  FILL71250x32550
timestamp 0
transform 1 0 4750 0 1 2170
box -6 -8 26 248
use FILL  FILL71250x36150
timestamp 0
transform -1 0 4770 0 -1 2650
box -6 -8 26 248
use FILL  FILL71250x39750
timestamp 0
transform 1 0 4750 0 1 2650
box -6 -8 26 248
use FILL  FILL71250x43350
timestamp 0
transform -1 0 4770 0 -1 3130
box -6 -8 26 248
use FILL  FILL71250x50550
timestamp 0
transform -1 0 4770 0 -1 3610
box -6 -8 26 248
use FILL  FILL71250x54150
timestamp 0
transform 1 0 4750 0 1 3610
box -6 -8 26 248
use FILL  FILL71250x57750
timestamp 0
transform -1 0 4770 0 -1 4090
box -6 -8 26 248
use FILL  FILL71250x61350
timestamp 0
transform 1 0 4750 0 1 4090
box -6 -8 26 248
<< labels >>
flabel metal1 s 4782 2 4842 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -62 2 -2 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 1477 -23 1483 -17 7 FreeSans 16 270 0 0 Cin[5]
port 2 nsew
flabel metal2 s 1757 -23 1763 -17 7 FreeSans 16 270 0 0 Cin[4]
port 3 nsew
flabel metal2 s 1897 -23 1903 -17 7 FreeSans 16 270 0 0 Cin[3]
port 4 nsew
flabel metal2 s 1937 -23 1943 -17 7 FreeSans 16 270 0 0 Cin[2]
port 5 nsew
flabel metal2 s 1977 -23 1983 -17 7 FreeSans 16 270 0 0 Cin[1]
port 6 nsew
flabel metal2 s 2117 -23 2123 -17 7 FreeSans 16 270 0 0 Cin[0]
port 7 nsew
flabel metal3 s -24 3556 -16 3564 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal2 s 4077 4617 4083 4623 3 FreeSans 16 90 0 0 Vld
port 9 nsew
flabel metal3 s -24 3516 -16 3524 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -24 3476 -16 3484 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -24 2996 -16 3004 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -24 2756 -16 2764 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal2 s 4237 4617 4243 4623 3 FreeSans 16 90 0 0 Xout[3]
port 14 nsew
flabel metal2 s 4197 4617 4203 4623 3 FreeSans 16 90 0 0 Xout[2]
port 15 nsew
flabel metal2 s 4157 4617 4163 4623 3 FreeSans 16 90 0 0 Xout[1]
port 16 nsew
flabel metal2 s 4117 4617 4123 4623 3 FreeSans 16 90 0 0 Xout[0]
port 17 nsew
flabel metal3 s 4816 1316 4824 1324 3 FreeSans 16 0 0 0 Yin[3]
port 18 nsew
flabel metal3 s 4816 3676 4824 3684 3 FreeSans 16 0 0 0 Yin[2]
port 19 nsew
flabel metal3 s 4816 3716 4824 3724 3 FreeSans 16 0 0 0 Yin[1]
port 20 nsew
flabel metal3 s 4816 3956 4824 3964 3 FreeSans 16 0 0 0 Yin[0]
port 21 nsew
flabel metal2 s 4637 4617 4643 4623 3 FreeSans 16 90 0 0 Yout[3]
port 22 nsew
flabel metal2 s 4557 4617 4563 4623 3 FreeSans 16 90 0 0 Yout[2]
port 23 nsew
flabel metal2 s 4317 4617 4323 4623 3 FreeSans 16 90 0 0 Yout[1]
port 24 nsew
flabel metal2 s 4277 4617 4283 4623 3 FreeSans 16 90 0 0 Yout[0]
port 25 nsew
flabel metal2 s 4017 4617 4023 4623 3 FreeSans 16 90 0 0 clk
port 26 nsew
<< properties >>
string FIXED_BBOX -40 -40 4820 4620
<< end >>
