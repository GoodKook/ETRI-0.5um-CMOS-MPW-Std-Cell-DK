magic
tech scmos
magscale 1 2
timestamp 1727271071
<< nwell >>
rect -12 154 131 272
rect 14 146 80 154
<< ntransistor >>
rect 20 22 24 42
rect 40 22 44 62
rect 50 22 54 62
rect 70 22 74 62
rect 80 22 84 62
<< ptransistor >>
rect 20 198 24 238
rect 40 158 44 238
rect 50 158 54 238
rect 70 166 74 246
rect 80 166 84 246
<< ndiffusion >>
rect 28 42 40 62
rect 18 22 20 42
rect 24 22 26 42
rect 38 22 40 42
rect 44 22 50 62
rect 54 54 70 62
rect 54 22 56 54
rect 68 22 70 54
rect 74 22 80 62
rect 84 22 86 62
<< pdiffusion >>
rect 61 238 70 246
rect 18 198 20 238
rect 24 198 26 238
rect 38 198 40 238
rect 30 158 40 198
rect 44 158 50 238
rect 54 174 56 238
rect 68 174 70 238
rect 54 166 70 174
rect 74 166 80 246
rect 84 166 86 246
rect 54 158 62 166
<< ndcontact >>
rect 6 22 18 42
rect 26 22 38 42
rect 56 22 68 54
rect 86 22 98 62
<< pdcontact >>
rect 6 198 18 238
rect 26 198 38 238
rect 56 174 68 238
rect 86 166 98 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 125 266
<< polysilicon >>
rect 20 246 54 250
rect 70 246 74 250
rect 80 246 84 250
rect 20 238 24 246
rect 40 238 44 242
rect 50 238 54 246
rect 20 194 24 198
rect 10 190 24 194
rect 10 103 14 190
rect 40 144 44 158
rect 50 154 54 158
rect 70 144 74 166
rect 28 140 44 144
rect 53 140 74 144
rect 28 109 32 140
rect 53 129 57 140
rect 10 51 14 91
rect 28 70 32 97
rect 28 66 44 70
rect 40 62 44 66
rect 50 62 54 117
rect 70 62 74 66
rect 80 62 84 166
rect 10 46 24 51
rect 20 42 24 46
rect 20 14 24 22
rect 40 18 44 22
rect 50 18 54 22
rect 70 14 74 22
rect 80 18 84 22
rect 20 10 74 14
<< polycontact >>
rect 45 117 57 129
rect 4 91 16 103
rect 24 97 36 109
rect 84 97 96 109
<< metal1 >>
rect -6 266 125 268
rect -6 252 125 254
rect 26 238 38 252
rect 86 246 98 252
rect 6 164 12 198
rect 68 174 70 176
rect 56 170 70 174
rect 6 158 55 164
rect 47 129 55 158
rect 64 117 70 170
rect 46 70 54 117
rect 6 64 54 70
rect 6 42 12 64
rect 64 58 70 103
rect 56 54 70 58
rect 68 52 70 54
rect 26 8 38 22
rect 86 8 98 22
rect -6 6 126 8
rect -6 -8 126 -6
<< m2contact >>
rect 3 103 17 117
rect 23 83 37 97
rect 63 103 77 117
rect 83 83 97 97
<< metal2 >>
rect 6 117 14 134
rect 66 117 74 134
rect 26 66 34 83
rect 86 66 94 83
<< m1p >>
rect -6 252 125 268
rect -6 -8 126 8
<< m2p >>
rect 6 117 14 134
rect 66 117 74 134
rect 26 66 34 83
rect 86 66 94 83
<< labels >>
rlabel metal1 -6 252 106 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 106 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal2 10 131 10 131 1 S
port 3 n signal input
rlabel metal2 70 133 70 133 5 Y
port 4 n signal output
rlabel metal2 30 71 30 71 1 B
port 2 n signal input
rlabel metal2 90 71 90 71 1 A
port 1 n signal input
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
