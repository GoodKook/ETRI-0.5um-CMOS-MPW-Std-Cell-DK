magic
tech scmos
magscale 1 2
timestamp 1727401709
<< nwell >>
rect -14 154 132 272
<< ntransistor >>
rect 24 14 28 54
rect 32 14 36 54
rect 52 14 56 54
rect 60 14 64 54
<< ptransistor >>
rect 20 166 24 246
rect 40 166 44 246
rect 60 166 64 246
rect 80 166 84 246
<< ndiffusion >>
rect 22 14 24 54
rect 28 14 32 54
rect 36 14 38 54
rect 50 14 52 54
rect 56 14 60 54
rect 64 14 66 54
<< pdiffusion >>
rect 18 168 20 246
rect 6 166 20 168
rect 24 180 26 246
rect 38 180 40 246
rect 24 166 40 180
rect 44 168 46 246
rect 58 168 60 246
rect 44 166 60 168
rect 64 234 80 246
rect 64 166 66 234
rect 78 166 80 234
rect 84 166 86 246
<< ndcontact >>
rect 10 14 22 54
rect 38 14 50 54
rect 66 14 78 54
<< pdcontact >>
rect 6 168 18 246
rect 26 180 38 246
rect 46 168 58 246
rect 66 166 78 234
rect 86 166 98 246
<< psubstratepcontact >>
rect -6 -6 126 6
<< nsubstratencontact >>
rect -6 254 126 266
<< polysilicon >>
rect 20 246 24 250
rect 40 246 44 250
rect 60 246 64 250
rect 80 246 84 250
rect 20 144 24 166
rect 40 144 44 166
rect 11 138 24 144
rect 32 138 44 144
rect 11 109 17 138
rect 32 123 36 138
rect 60 123 64 166
rect 80 144 84 166
rect 80 138 90 144
rect 60 111 63 123
rect 11 83 17 97
rect 11 71 28 83
rect 24 54 28 71
rect 32 54 36 111
rect 60 82 64 111
rect 52 71 64 82
rect 84 109 90 138
rect 52 54 56 71
rect 84 63 90 97
rect 60 59 90 63
rect 60 54 64 59
rect 24 10 28 14
rect 32 10 36 14
rect 52 10 56 14
rect 60 10 64 14
<< polycontact >>
rect 25 111 37 123
rect 63 111 75 123
rect 5 97 17 109
rect 84 97 96 109
<< metal1 >>
rect -6 266 126 268
rect -6 252 126 254
rect 26 246 38 252
rect 18 168 46 174
rect 58 240 86 246
rect 66 160 78 166
rect 51 154 78 160
rect 23 123 37 137
rect 51 97 57 154
rect 63 123 77 137
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
rect 43 54 50 83
rect 10 8 22 14
rect 66 8 78 14
rect -6 6 126 8
rect -6 -8 126 -6
<< m1p >>
rect 23 123 37 137
rect 63 123 77 137
rect 3 83 17 97
rect 43 83 57 97
rect 83 83 97 97
<< labels >>
rlabel metal1 -6 252 126 268 0 vdd
port 5 nsew power bidirectional abutment
rlabel metal1 -6 -8 126 8 0 gnd
port 6 nsew ground bidirectional abutment
rlabel metal1 23 123 37 137 0 B
port 1 nsew signal input
rlabel metal1 3 83 17 97 0 A
port 0 nsew signal input
rlabel metal1 43 83 57 97 0 Y
port 4 nsew signal output
rlabel metal1 63 123 77 137 0 D
port 3 nsew signal input
rlabel metal1 83 83 97 97 0 C
port 2 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 120 260
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
