magic
tech scmos
magscale 1 30
timestamp 1754274956
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
rect 147800 8500 172930 8670
rect 150400 8300 172930 8500
<< metal1 >>
rect 131200 103900 143000 113100
rect 45650 64600 58100 71400
<< m2contact >>
rect 143000 103900 144500 113100
rect 44300 64600 45650 71400
<< metal2 >>
rect 49000 133700 49300 145900
rect 62500 134300 62800 145900
rect 76000 134900 76300 145900
rect 89500 144600 89800 145900
rect 89502 135500 89798 144600
rect 103000 136100 103350 145900
rect 116500 136700 116800 145900
rect 47500 130200 47800 132800
rect 44100 129900 47800 130200
rect 118650 129700 119050 132500
rect 119600 129700 119950 133100
rect 120250 129700 120550 133700
rect 120850 129700 121150 134300
rect 121450 129945 121750 134900
rect 122050 129945 122350 135500
rect 121450 129840 121755 129945
rect 122050 129840 122355 129945
rect 122550 129850 122950 136400
rect 130000 133800 130300 145900
rect 123400 129900 123700 133500
rect 127000 132300 139800 132600
rect 121450 129700 121750 129840
rect 122050 129700 122350 129840
rect 127000 129800 127500 132300
rect 128200 131700 139100 132000
rect 128200 129800 128700 131700
rect 140700 130000 145900 130300
rect 44100 116400 49400 116700
rect 140000 116500 145900 116800
rect 144500 103900 145900 113100
rect 44100 102900 48800 103200
rect 138000 100300 145900 100600
rect 44100 89400 50300 89700
rect 137400 86800 145900 87100
rect 44100 75900 50900 76200
rect 136800 73300 145900 73600
rect 44150 64600 44300 71400
rect 80800 59500 81100 60300
rect 44100 48900 49700 49200
rect 73300 44100 73600 59200
rect 84900 56900 85200 60300
rect 87000 57700 87300 60300
rect 87600 58300 87900 60300
rect 88300 58900 88600 60300
rect 90400 59500 90700 60300
rect 136200 59800 145900 60100
rect 86800 44100 87100 56600
rect 100300 44100 100600 57400
rect 113800 44100 114100 58000
rect 127300 44100 127600 58600
rect 134300 45800 134600 59200
rect 140800 44100 141100 45500
<< m3contact >>
rect 116500 136400 117100 136700
rect 122250 136400 122950 136700
rect 103000 135800 103650 136100
rect 122050 135500 122350 136100
rect 89500 135200 90100 135500
rect 121450 134900 121750 135500
rect 76000 134600 76600 134900
rect 120850 134300 121150 134900
rect 62500 134000 63100 134300
rect 120250 133700 120550 134300
rect 49000 133400 49600 133700
rect 119600 133100 119950 133700
rect 47500 132800 48100 133100
rect 118650 132500 119050 133100
rect 123400 133500 124000 133800
rect 129700 133500 130300 133800
rect 139800 132300 140400 132600
rect 139100 131700 139700 132000
rect 140100 130000 140700 130300
rect 49400 116400 50000 116700
rect 139400 116500 140000 116800
rect 48800 102900 49400 103200
rect 137400 100300 138000 100600
rect 50300 89400 50600 90000
rect 136800 86800 137400 87100
rect 50900 75900 51200 76500
rect 136200 73300 136800 73600
rect 73300 59200 73900 59500
rect 80500 59200 81100 59500
rect 49700 48900 50000 49500
rect 135600 59800 136200 60100
rect 90400 59200 91000 59500
rect 134000 59200 134600 59500
rect 88300 58600 88900 58900
rect 127000 58600 127600 58900
rect 87600 58000 88200 58300
rect 113500 58000 114100 58300
rect 87000 57400 87600 57700
rect 100000 57400 100600 57700
rect 84900 56600 85500 56900
rect 86500 56600 87100 56900
rect 134300 45500 134600 45800
rect 140800 45500 141100 45800
<< metal3 >>
rect 117100 136400 122250 136700
rect 103650 135800 122050 136100
rect 90100 135200 121450 135500
rect 76600 134600 120850 134900
rect 63100 134000 120250 134300
rect 49600 133400 119600 133700
rect 124000 133500 129700 133800
rect 48100 132800 118650 133100
rect 131000 119800 137700 120100
rect 49700 113500 50000 116400
rect 131000 116100 137100 116400
rect 131000 115500 136500 115800
rect 49700 113200 58500 113500
rect 49100 112600 58400 112900
rect 49100 103200 49400 112600
rect 49700 112000 58400 112300
rect 49700 49500 50000 112000
rect 50300 105300 58400 105700
rect 50300 90000 50600 105300
rect 50900 101700 58400 102000
rect 50900 76500 51200 101700
rect 131000 80300 135900 80600
rect 135600 60100 135900 80300
rect 136200 73600 136500 115500
rect 136800 87100 137100 116100
rect 137400 100600 137700 119800
rect 139400 116800 139700 131700
rect 140100 130300 140400 132300
rect 73900 59200 80500 59500
rect 91000 59200 134000 59500
rect 88900 58600 127000 58900
rect 88200 58000 113500 58300
rect 87600 57400 100000 57700
rect 85500 56600 86500 56900
rect 134600 45500 140800 45800
use PIC  CIN_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 129500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_1
timestamp 1569139307
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_2
timestamp 1569139307
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_3
timestamp 1569139307
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_4
timestamp 1569139307
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use PIC  CIN_5
timestamp 1569139307
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use PIC  CLK
timestamp 1569139307
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use fir_pe_Core  fir_pe_Core_0
timestamp 1754220398
transform 1 0 58710 0 1 60600
box -930 -360 72630 69345
use PVSS  GND ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 -1 171100 1 0 102500
box 0 -9150 12000 25300
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1569139307
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1569139307
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1569139307
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use MY_LOGO  MY_LOGO_0
timestamp 1724157349
transform 1 0 156620 0 1 9565
box 180 225 21510 9045
use PIC  PAD_0
timestamp 1569139307
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1569139307
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1569139307
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use PIC  RDY
timestamp 1569139307
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use PVDD  VDD ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 74000
box 0 -9150 12000 25300
use POB8  VLD ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  XIN_0
timestamp 1569139307
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use PIC  XIN_1
timestamp 1569139307
transform 0 1 18900 -1 0 101000
box -100 -9150 12100 25300
use PIC  XIN_2
timestamp 1569139307
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PIC  XIN_3
timestamp 1569139307
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use POB8  XOUT_0
timestamp 1569139307
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT_1
timestamp 1569139307
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT_2
timestamp 1569139307
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB8  XOUT_3
timestamp 1569139307
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  YIN_0
timestamp 1569139307
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC  YIN_1
timestamp 1569139307
transform 0 -1 171100 1 0 75500
box -100 -9150 12100 25300
use PIC  YIN_2
timestamp 1569139307
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PIC  YIN_3
timestamp 1569139307
transform 0 -1 171100 1 0 48500
box -100 -9150 12100 25300
use POB8  YOUT_0
timestamp 1569139307
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT_1
timestamp 1569139307
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use POB8  YOUT_2
timestamp 1569139307
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use POB8  YOUT_3
timestamp 1569139307
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
<< end >>
