magic
tech scmos
magscale 1 30
timestamp 1740713424
<< checkpaint >>
rect 18300 186927 44800 197000
rect 13915 181835 44800 186927
rect 46919 186419 142100 190000
rect 46919 181835 143266 186419
rect 6771 176042 185015 181835
rect 6771 175958 328570 176042
rect 205 167042 328570 175958
rect 205 160774 185015 167042
rect 6771 143081 185015 160774
rect 0 142100 185015 143081
rect 0 102896 190000 142100
rect -13866 102380 190000 102896
rect -25613 89180 190000 102380
rect -24170 89077 190000 89180
rect -17472 83925 190000 89077
rect 0 47900 190000 83925
rect 6771 46919 190000 47900
rect 6771 32547 185015 46919
rect 6771 31724 186496 32547
rect -4457 10781 186496 31724
rect -4457 8670 185015 10781
rect -4457 7765 35955 8670
rect 205 1458 35955 7765
rect -600 -600 630 630
rect 46919 0 142100 8670
<< metal1 >>
rect 44700 91600 50500 98400
rect 139500 76800 145200 86100
rect 145800 76800 145900 86100
rect 142400 54200 145500 58400
rect 145800 54200 145900 58400
rect 142400 49100 143000 54200
rect 142400 47600 143000 47700
<< m2contact >>
rect 44100 91600 44700 98400
rect 145200 76800 145800 86100
rect 145500 54200 145800 58400
rect 142400 47300 143000 47600
<< metal2 >>
rect 59800 141900 60200 145900
rect 60200 140100 72400 140500
rect 44800 130200 45200 140100
rect 73300 139800 73700 145900
rect 74400 141500 86100 141900
rect 86800 141200 87200 145900
rect 87200 140100 99600 140500
rect 87200 139400 99600 139800
rect 100300 138400 100700 145900
rect 101400 141500 113100 141900
rect 101400 140800 113100 141200
rect 113800 139100 114200 145900
rect 114900 140100 121300 140500
rect 114900 139400 121300 139800
rect 114200 138000 121300 138400
rect 122000 137600 122400 141500
rect 127300 139800 127700 145900
rect 140800 143400 141200 145900
rect 132200 143000 141200 143400
rect 125600 138800 126000 139400
rect 125600 138400 127700 138800
rect 127300 137600 127700 138400
rect 128500 137600 128900 141500
rect 129500 137600 129900 140800
rect 132200 137600 132600 143000
rect 144100 140800 145900 141200
rect 134000 137600 134400 140100
rect 135700 137600 136100 139400
rect 136600 137600 137000 138700
rect 137300 137600 137700 138000
rect 44100 129800 45200 130200
rect 141900 127300 145900 127700
rect 44100 116300 47500 116700
rect 44100 102800 46800 103200
rect 47100 97600 47500 116300
rect 141200 113800 145900 114200
rect 141500 101500 141900 113100
rect 140500 100300 145900 100700
rect 44100 86600 48200 87000
rect 47800 74900 48200 86600
rect 48500 73500 48900 84100
rect 44100 73100 48900 73500
rect 49200 60000 49600 81400
rect 145800 77700 145900 86100
rect 140500 73300 145900 73700
rect 44100 59600 49600 60000
rect 145800 54200 145900 58400
rect 85300 49600 85700 50100
rect 62900 49200 76000 49600
rect 49000 44100 49400 49200
rect 83100 48500 93000 48900
rect 62500 44100 62900 48500
rect 76000 47800 85300 48200
rect 76000 44100 76400 47800
rect 89500 44100 89900 47100
rect 95600 46100 96000 50100
rect 103300 48900 103700 50100
rect 107800 48200 108200 50100
rect 101700 47800 108200 48200
rect 109300 47500 109700 50100
rect 110000 46800 110400 50100
rect 103000 44100 103400 46400
rect 110900 45700 121400 46100
rect 127300 44100 127700 45700
rect 142400 45300 143000 47300
rect 134900 45000 143000 45300
rect 134900 44000 139500 45000
<< m3contact >>
rect 59800 141500 60200 141900
rect 44800 140100 45200 140500
rect 59800 140100 60200 140500
rect 72400 140100 72800 140500
rect 74000 141500 74400 141900
rect 86100 141500 86500 141900
rect 86800 140800 87200 141200
rect 86800 140100 87200 140500
rect 99600 140100 100000 140500
rect 73300 139400 73700 139800
rect 86800 139400 87200 139800
rect 99600 139400 100000 139800
rect 101000 141500 101400 141900
rect 113100 141500 113500 141900
rect 101000 140800 101400 141200
rect 113100 140800 113500 141200
rect 122000 141500 122400 141900
rect 114500 140100 114900 140500
rect 121300 140100 121700 140500
rect 114500 139400 114900 139800
rect 121300 139400 121700 139800
rect 113800 138700 114200 139100
rect 100300 138000 100700 138400
rect 113800 138000 114200 138400
rect 121300 138000 121700 138400
rect 125600 139400 126000 139800
rect 127300 139400 127700 139800
rect 128500 141500 128900 141900
rect 129500 140800 129900 141200
rect 143700 140800 144100 141200
rect 134000 140100 134400 140500
rect 135700 139400 136100 139800
rect 136600 138700 137000 139100
rect 137300 138000 137700 138400
rect 141500 127300 141900 127700
rect 46400 102400 46800 102800
rect 140800 113800 141200 114200
rect 141500 113100 141900 113500
rect 141500 101100 141900 101500
rect 140100 100300 140500 100700
rect 47100 97200 47500 97600
rect 47800 74500 48200 74900
rect 48500 84100 48900 84500
rect 49200 81400 49600 81800
rect 140100 73300 140500 73700
rect 49000 49200 49400 49600
rect 62500 49200 62900 49600
rect 76000 49200 76400 49600
rect 85300 49200 85700 49600
rect 62500 48500 62900 48900
rect 82700 48500 83100 48900
rect 93000 48500 93400 48900
rect 85300 47800 85700 48200
rect 89500 47100 89900 47500
rect 103300 48500 103700 48900
rect 101300 47800 101700 48200
rect 109300 47100 109700 47500
rect 95600 45700 96000 46100
rect 103000 46400 103400 46800
rect 110000 46400 110400 46800
rect 110500 45700 110900 46100
rect 121400 45700 121800 46100
rect 127300 45700 127700 46100
<< metal3 >>
rect 60200 141500 74000 141900
rect 86500 141500 101000 141900
rect 113500 141500 122000 141900
rect 128900 141500 144100 141900
rect 143700 141200 144100 141500
rect 87200 140800 101000 141200
rect 113500 140800 129500 141200
rect 45200 140100 59800 140500
rect 72800 140100 86800 140500
rect 100000 140100 114500 140500
rect 121700 140100 134000 140500
rect 73700 139400 86800 139800
rect 100000 139400 114500 139800
rect 121700 139400 125600 139800
rect 127700 139400 135700 139800
rect 114200 138700 136600 139100
rect 100700 138000 113800 138400
rect 121700 138000 137300 138400
rect 139600 135100 141200 135500
rect 140800 114200 141200 135100
rect 141500 113500 141900 127300
rect 139600 109300 140500 109700
rect 46800 102400 50300 102800
rect 140100 100700 140500 109300
rect 47500 97200 50300 97600
rect 141500 92300 141900 101100
rect 139600 91900 141900 92300
rect 48900 84100 50300 84500
rect 49600 81400 50300 81800
rect 139600 77200 140500 77600
rect 48200 74500 50400 74900
rect 49900 72990 50400 74500
rect 140100 73700 140500 77200
rect 49890 72690 50400 72990
rect 49400 49200 62500 49600
rect 76400 49200 85300 49600
rect 62900 48500 82700 48900
rect 93400 48500 103300 48900
rect 85700 47800 101300 48200
rect 89900 47100 109300 47500
rect 103400 46400 110000 46800
rect 96000 45700 110500 46100
rect 121800 45700 127300 46100
use PIC  ABCMD_I_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 -1 171100 1 0 89000
box -100 -9150 12100 25300
use PIC  ABCMD_I_1
timestamp 1569139307
transform 0 -1 171100 1 0 102500
box -100 -9150 12100 25300
use PIC  ABCMD_I_2
timestamp 1569139307
transform 0 -1 171100 1 0 116000
box -100 -9150 12100 25300
use PIC  ABCMD_I_3
timestamp 1569139307
transform 0 -1 171100 1 0 129500
box -100 -9150 12100 25300
use PIC  ABCMD_I_4
timestamp 1569139307
transform 1 0 129500 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_5
timestamp 1569139307
transform 1 0 116000 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_6
timestamp 1569139307
transform 1 0 102500 0 -1 171100
box -100 -9150 12100 25300
use PIC  ABCMD_I_7
timestamp 1569139307
transform 1 0 89000 0 -1 171100
box -100 -9150 12100 25300
use POB4  ACC_O_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 87500
box -100 -9150 12100 25300
use POB4  ACC_O_1
timestamp 1569139307
transform 0 1 18900 -1 0 74000
box -100 -9150 12100 25300
use POB4  ACC_O_2
timestamp 1569139307
transform 0 1 18900 -1 0 60500
box -100 -9150 12100 25300
use POB4  ACC_O_3
timestamp 1569139307
transform 1 0 48500 0 1 18900
box -100 -9150 12100 25300
use POB4  ACC_O_4
timestamp 1569139307
transform 1 0 62000 0 1 18900
box -100 -9150 12100 25300
use POB4  ACC_O_5
timestamp 1569139307
transform 1 0 75500 0 1 18900
box -100 -9150 12100 25300
use POB4  ACC_O_6
timestamp 1569139307
transform 1 0 89000 0 1 18900
box -100 -9150 12100 25300
use POB4  ACC_O_7
timestamp 1569139307
transform 1 0 102500 0 1 18900
box -100 -9150 12100 25300
use ALU8_Mult_Core  ALU8_Mult_Core_0
timestamp 1740459297
transform 1 0 51330 0 1 50340
box -1050 -360 88350 87345
use PANA  ANA_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 129500 0 1 18900
box -100 -9150 12095 25300
use PANA  ANA_1
timestamp 1569139307
transform 0 -1 171100 1 0 48500
box -100 -9150 12095 25300
use PIC  CLK
timestamp 1569139307
transform 1 0 48500 0 -1 171100
box -100 -9150 12100 25300
use PIC  FLAG_I
timestamp 1569139307
transform 1 0 116000 0 1 18900
box -100 -9150 12100 25300
use IOFILLER18  IOFILLER18_0 ~/ETRI050_DesignKit/pads_ETRI
timestamp 1725930584
transform 0 -1 171100 -1 0 75646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_1
timestamp 1725930584
transform 0 -1 171098 -1 0 62146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_2
timestamp 1725930584
transform 0 -1 171100 -1 0 102646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_3
timestamp 1725930584
transform 0 -1 171100 -1 0 89146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_4
timestamp 1725930584
transform 0 -1 171102 -1 0 129646
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_5
timestamp 1725930584
transform 0 -1 171100 -1 0 116146
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_6
timestamp 1725930584
transform 1 0 73845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_7
timestamp 1725930584
transform 1 0 60345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_8
timestamp 1725930584
transform 1 0 100845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_9
timestamp 1725930584
transform 1 0 87345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_10
timestamp 1725930584
transform 1 0 127845 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_11
timestamp 1725930584
transform 1 0 114345 0 1 18900
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_12
timestamp 1725930584
transform 0 1 18899 -1 0 75655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_13
timestamp 1725930584
transform 0 1 18899 -1 0 62155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_14
timestamp 1725930584
transform 0 1 18900 -1 0 102655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_15
timestamp 1725930584
transform 0 1 18900 -1 0 89155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_16
timestamp 1725930584
transform 1 0 73845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_17
timestamp 1725930584
transform 0 1 18897 -1 0 116155
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_18
timestamp 1725930584
transform 0 1 18900 -1 0 129655
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_19
timestamp 1725930584
transform 1 0 60345 0 -1 171101
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_20
timestamp 1725930584
transform 1 0 100845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_21
timestamp 1725930584
transform 1 0 87344 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_22
timestamp 1725930584
transform 1 0 127845 0 -1 171100
box -60 0 1860 25060
use IOFILLER18  IOFILLER18_23
timestamp 1725930584
transform 1 0 114345 0 -1 171100
box -60 0 1860 25060
use IOFILLER50  IOFILLER50_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 43621 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_1
timestamp 1569139307
transform 1 0 141360 0 1 18900
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_2
timestamp 1569139307
transform 1 0 141345 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_3
timestamp 1569139307
transform 1 0 43638 0 -1 171100
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_4
timestamp 1569139307
transform 0 1 18900 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_5
timestamp 1569139307
transform 0 1 18900 -1 0 146379
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_6
timestamp 1569139307
transform 0 -1 171100 -1 0 48655
box -35 0 5035 25060
use IOFILLER50  IOFILLER50_7
timestamp 1569139307
transform 0 -1 171100 -1 0 146346
box -35 0 5035 25060
use PIC  LOADA_I
timestamp 1569139307
transform 1 0 75500 0 -1 171100
box -100 -9150 12100 25300
use PIC  LOADB_I
timestamp 1569139307
transform 1 0 62000 0 -1 171100
box -100 -9150 12100 25300
use PIC  LOADCMD_I
timestamp 1569139307
transform 0 1 18900 -1 0 141500
box -100 -9150 12100 25300
use PIC  MULH_I
timestamp 1569139307
transform 0 1 18900 -1 0 128000
box -100 -9150 12100 25300
use PIC  MULL_I
timestamp 1569139307
transform 0 1 18900 -1 0 114500
box -100 -9150 12100 25300
use PCORNER  PCORNER_0 ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 1 0 18900 0 1 18900
box 0 0 25300 25300
use PCORNER  PCORNER_1
timestamp 1569139307
transform 1 0 18900 0 -1 171100
box 0 0 25300 25300
use PCORNER  PCORNER_2
timestamp 1569139307
transform 0 -1 171100 1 0 18900
box 0 0 25300 25300
use PCORNER  PCORNER_3
timestamp 1569139307
transform -1 0 171100 0 -1 171100
box 0 0 25300 25300
use pdiode  pdiode_0 ~/ETRI050_DesignKit/analog_ETRI/GDS_Magic
timestamp 1569140870
transform 1 0 141330 0 1 46770
box 0 0 2700 2700
use PIC  RESET
timestamp 1569139307
transform 0 -1 171100 1 0 62000
box -100 -9150 12100 25300
use PVDD  VDD ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 1 18900 -1 0 101000
box 0 -9150 12000 25300
use PVSS  VSS ~/ETRI050_DesignKit/pads_ETRI/GDS_Magic
timestamp 1569139307
transform 0 -1 171100 1 0 75500
box 0 -9150 12000 25300
<< end >>
