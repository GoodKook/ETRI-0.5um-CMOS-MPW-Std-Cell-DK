magic
tech scmos
magscale 1 2
timestamp 1727833531
<< nwell >>
rect -12 134 92 252
<< ntransistor >>
rect 20 14 24 54
rect 40 14 44 54
<< ptransistor >>
rect 20 146 24 226
rect 40 146 44 226
<< ndiffusion >>
rect 18 14 20 54
rect 24 14 26 54
rect 38 14 40 54
rect 44 14 46 54
<< pdiffusion >>
rect 6 224 20 226
rect 18 146 20 224
rect 24 146 26 226
rect 38 146 40 226
rect 44 146 46 226
<< ndcontact >>
rect 6 14 18 54
rect 26 14 38 54
rect 46 14 58 54
<< pdcontact >>
rect 6 146 18 224
rect 26 146 38 226
rect 46 146 58 226
<< psubstratepcontact >>
rect -6 -6 86 6
<< nsubstratencontact >>
rect -6 234 86 246
<< polysilicon >>
rect 20 226 24 230
rect 40 226 44 230
rect 20 142 24 146
rect 40 142 44 146
rect 20 138 44 142
rect 20 89 24 138
rect 16 77 24 89
rect 20 62 24 77
rect 20 58 44 62
rect 20 54 24 58
rect 40 54 44 58
rect 20 10 24 14
rect 40 10 44 14
<< polycontact >>
rect 4 77 16 89
<< metal1 >>
rect -6 246 86 248
rect -6 232 86 234
rect 6 224 18 232
rect 46 226 58 232
rect 28 103 37 146
rect 28 89 43 103
rect 28 54 37 89
rect 6 8 18 14
rect 46 8 58 14
rect -6 6 86 8
rect -6 -8 86 -6
<< m2contact >>
rect 3 89 17 103
rect 43 89 57 103
<< metal2 >>
rect 3 103 17 117
rect 43 103 57 117
<< m2p >>
rect 3 103 17 117
rect 43 103 57 117
<< labels >>
rlabel metal1 -6 -8 86 8 0 gnd
port 3 nsew ground bidirectional abutment
rlabel metal1 -6 232 86 248 0 vdd
port 2 nsew power bidirectional abutment
rlabel metal2 3 103 17 117 0 A
port 0 nsew signal input
rlabel metal2 43 103 57 117 0 Y
port 1 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 80 240
string LEFclass CORE
string LEFsite core
string LEFsymmetry X Y
<< end >>
