** sch_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1_TB.sch
**.subckt inverter_x1_TB
Vdd VDD GND 5
R1 VDD Vout 1mega m=1
Vin Vin GND pulse(0 5 0 1n 1n 5n 12n)
x1 Vin Vout VDD GND inverter_x1
**** begin user architecture code



* ngspice commands
.include ~/ETRI050_DesignKit/devel/tech/05cmos_model_240201.lib
.dc vin 0 5 0.01
.tran 0.01 70n
.save all



**** end user architecture code
**.ends

* expanding   symbol:  /home/goodkook/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1.sym # of pins=4
** sym_path: /home/goodkook/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1.sym
.include ~/ETRI050_DesignKit/Tutorials/1-2_Inverter_Magic/inverter_x1.spice
.GLOBAL VDD
.GLOBAL GND
.end
