magic
tech scmos
magscale 1 2
timestamp 1725247039
<< checkpaint >>
rect -114 -64 5934 5563
<< metal1 >>
rect -63 5218 -3 5478
rect 5790 5462 5883 5478
rect 3107 5437 3133 5443
rect 3687 5437 3713 5443
rect 1507 5397 1533 5403
rect 2967 5397 3003 5403
rect 1773 5383 1787 5393
rect 1747 5380 1787 5383
rect 1747 5377 1783 5380
rect 2587 5383 2600 5387
rect 2740 5383 2753 5387
rect 2587 5373 2603 5383
rect 2597 5347 2603 5373
rect 2737 5373 2753 5383
rect 2997 5383 3003 5397
rect 3417 5397 3473 5403
rect 3120 5383 3133 5387
rect 2997 5377 3023 5383
rect 2737 5347 2743 5373
rect 2597 5337 2613 5347
rect 2600 5333 2613 5337
rect 2727 5337 2743 5347
rect 3017 5347 3023 5377
rect 3117 5373 3133 5383
rect 3417 5383 3423 5397
rect 3647 5397 3773 5403
rect 3397 5377 3423 5383
rect 3017 5337 3033 5347
rect 2727 5333 2740 5337
rect 3020 5333 3033 5337
rect 3117 5343 3123 5373
rect 3397 5347 3403 5377
rect 4067 5383 4080 5387
rect 4067 5373 4083 5383
rect 5727 5383 5740 5387
rect 5727 5373 5743 5383
rect 3097 5340 3123 5343
rect 3093 5337 3123 5340
rect 3093 5327 3107 5337
rect 3387 5337 3403 5347
rect 4077 5346 4083 5373
rect 5737 5347 5743 5373
rect 3387 5333 3400 5337
rect 5737 5337 5753 5347
rect 5740 5333 5753 5337
rect 2747 5317 2773 5323
rect 2827 5317 2913 5323
rect 3247 5317 3313 5323
rect 4727 5317 4773 5323
rect 5427 5317 5519 5323
rect 3087 5297 3113 5303
rect 2747 5277 2773 5283
rect -63 5202 30 5218
rect -63 4698 -3 5202
rect 2867 5177 2893 5183
rect 3307 5177 3353 5183
rect 2647 5117 2673 5123
rect 3567 5117 3633 5123
rect 527 5097 633 5103
rect 2007 5097 2053 5103
rect 2567 5097 2673 5103
rect 3267 5097 3373 5103
rect 4141 5097 4273 5103
rect 4427 5097 4493 5103
rect 4887 5097 4933 5103
rect 5067 5097 5113 5103
rect 867 5083 880 5087
rect 1940 5083 1953 5087
rect 867 5073 883 5083
rect 877 5047 883 5073
rect 1937 5073 1953 5083
rect 2167 5083 2180 5087
rect 2600 5083 2613 5087
rect 2167 5073 2183 5083
rect 877 5037 893 5047
rect 880 5033 893 5037
rect 547 5017 653 5023
rect 1937 5026 1943 5073
rect 2177 5023 2183 5073
rect 2597 5073 2613 5083
rect 2740 5086 2760 5087
rect 2740 5083 2753 5086
rect 2737 5073 2753 5083
rect 2597 5047 2603 5073
rect 2737 5047 2743 5073
rect 3620 5083 3633 5087
rect 3617 5073 3633 5083
rect 3887 5083 3900 5087
rect 3887 5073 3903 5083
rect 4327 5083 4340 5087
rect 4327 5073 4343 5083
rect 4467 5083 4480 5087
rect 4467 5073 4483 5083
rect 2587 5037 2603 5047
rect 2587 5033 2600 5037
rect 2727 5037 2743 5047
rect 3617 5047 3623 5073
rect 3897 5047 3903 5073
rect 4337 5047 4343 5073
rect 3617 5037 3633 5047
rect 2727 5033 2740 5037
rect 3620 5033 3633 5037
rect 3897 5037 3913 5047
rect 3900 5033 3913 5037
rect 4327 5037 4343 5047
rect 4477 5043 4483 5073
rect 4457 5037 4483 5043
rect 5177 5047 5183 5093
rect 5300 5083 5313 5087
rect 5297 5073 5313 5083
rect 5620 5083 5633 5087
rect 5617 5073 5633 5083
rect 5297 5047 5303 5073
rect 5177 5037 5193 5047
rect 4327 5033 4340 5037
rect 2177 5017 2213 5023
rect 2547 5017 2613 5023
rect 3267 5017 3313 5023
rect 4457 5023 4463 5037
rect 5180 5033 5193 5037
rect 5287 5037 5303 5047
rect 5287 5033 5300 5037
rect 4427 5017 4463 5023
rect 5597 5023 5603 5053
rect 5617 5047 5623 5073
rect 5597 5017 5633 5023
rect 5607 4977 5633 4983
rect 5823 4958 5883 5462
rect 5790 4942 5883 4958
rect 2440 4863 2453 4867
rect 2437 4853 2453 4863
rect 2680 4863 2693 4867
rect 2677 4860 2693 4863
rect 2673 4853 2693 4860
rect 2960 4863 2973 4867
rect 2957 4853 2973 4863
rect 3920 4863 3933 4867
rect 3917 4853 3933 4863
rect 4060 4863 4073 4867
rect 4057 4853 4073 4863
rect 4187 4863 4200 4867
rect 4580 4863 4593 4867
rect 4187 4853 4203 4863
rect 737 4827 743 4853
rect 727 4817 743 4827
rect 2437 4823 2443 4853
rect 2673 4847 2687 4853
rect 2957 4827 2963 4853
rect 3917 4827 3923 4853
rect 4057 4827 4063 4853
rect 4197 4827 4203 4853
rect 2417 4820 2443 4823
rect 2413 4817 2443 4820
rect 727 4813 740 4817
rect 2413 4807 2427 4817
rect 2947 4817 2963 4827
rect 2947 4813 2960 4817
rect 3907 4817 3923 4827
rect 3907 4813 3920 4817
rect 4047 4817 4063 4827
rect 4047 4813 4060 4817
rect 4187 4817 4203 4827
rect 4577 4853 4593 4863
rect 5220 4863 5233 4867
rect 5217 4853 5233 4863
rect 5307 4863 5320 4867
rect 5460 4863 5473 4867
rect 5307 4853 5323 4863
rect 4577 4823 4583 4853
rect 5217 4827 5223 4853
rect 4577 4817 4603 4823
rect 4187 4813 4200 4817
rect 667 4797 773 4803
rect 827 4797 893 4803
rect 3047 4797 3173 4803
rect 4001 4797 4073 4803
rect 4597 4803 4603 4817
rect 5207 4817 5223 4827
rect 5317 4827 5323 4853
rect 5457 4853 5473 4863
rect 5600 4863 5613 4867
rect 5597 4853 5613 4863
rect 5457 4827 5463 4853
rect 5317 4817 5333 4827
rect 5207 4813 5220 4817
rect 5320 4813 5333 4817
rect 5447 4817 5463 4827
rect 5447 4813 5460 4817
rect 4597 4797 4633 4803
rect 5047 4797 5073 4803
rect 5307 4797 5393 4803
rect 5597 4803 5603 4853
rect 5567 4797 5603 4803
rect -63 4682 30 4698
rect -63 4178 -3 4682
rect 2847 4637 2893 4643
rect 2827 4617 2853 4623
rect 427 4577 453 4583
rect 1067 4577 1113 4583
rect 1767 4583 1780 4587
rect 1767 4573 1783 4583
rect 1887 4577 1913 4583
rect 2687 4583 2700 4587
rect 2687 4573 2703 4583
rect 2907 4577 2933 4583
rect 1777 4567 1783 4573
rect 1367 4563 1380 4567
rect 1777 4566 1800 4567
rect 1367 4553 1383 4563
rect 1777 4557 1793 4566
rect 1780 4553 1793 4557
rect 1377 4527 1383 4553
rect 1920 4563 1933 4567
rect 1917 4553 1933 4563
rect 1917 4527 1923 4553
rect 1377 4517 1393 4527
rect 1380 4513 1393 4517
rect 1907 4517 1923 4527
rect 1907 4513 1920 4517
rect 1347 4497 1413 4503
rect 1787 4497 1833 4503
rect 2697 4503 2703 4573
rect 3667 4577 3753 4583
rect 4517 4577 4553 4583
rect 3120 4563 3133 4567
rect 3117 4553 3133 4563
rect 3600 4563 3613 4567
rect 3597 4553 3613 4563
rect 2853 4527 2867 4533
rect 3117 4527 3123 4553
rect 2847 4520 2867 4527
rect 2847 4517 2863 4520
rect 2847 4513 2860 4517
rect 3107 4517 3123 4527
rect 3597 4527 3603 4553
rect 4380 4543 4393 4547
rect 4377 4533 4393 4543
rect 3597 4517 3613 4527
rect 3107 4513 3120 4517
rect 3600 4513 3613 4517
rect 4377 4523 4383 4533
rect 4517 4527 4523 4577
rect 4607 4577 4653 4583
rect 4727 4560 4763 4563
rect 4727 4557 4767 4560
rect 4753 4546 4767 4557
rect 4400 4523 4413 4527
rect 4357 4517 4383 4523
rect 2697 4497 2773 4503
rect 3247 4497 3293 4503
rect 4047 4497 4073 4503
rect 4357 4483 4363 4517
rect 4397 4513 4413 4523
rect 4517 4517 4533 4527
rect 4520 4513 4533 4517
rect 4397 4507 4403 4513
rect 4380 4506 4403 4507
rect 4387 4497 4403 4506
rect 4387 4493 4400 4497
rect 4357 4477 4413 4483
rect 4627 4457 4653 4463
rect 5823 4438 5883 4942
rect 5790 4422 5883 4438
rect 967 4357 1013 4363
rect 1367 4357 1453 4363
rect 4467 4357 4523 4363
rect 687 4343 700 4347
rect 687 4333 703 4343
rect 1527 4343 1540 4347
rect 1680 4343 1693 4347
rect 1527 4333 1543 4343
rect 697 4307 703 4333
rect 1537 4307 1543 4333
rect 1677 4333 1693 4343
rect 1787 4343 1800 4347
rect 1787 4333 1803 4343
rect 2307 4343 2320 4347
rect 2307 4340 2323 4343
rect 2307 4333 2327 4340
rect 3267 4343 3280 4347
rect 3267 4333 3283 4343
rect 3387 4343 3400 4347
rect 3513 4343 3527 4353
rect 3387 4333 3403 4343
rect 3513 4340 3543 4343
rect 3517 4337 3543 4340
rect 1677 4307 1683 4333
rect 687 4297 703 4307
rect 687 4293 700 4297
rect 1527 4297 1543 4307
rect 1527 4293 1540 4297
rect 1667 4297 1683 4307
rect 1797 4307 1803 4333
rect 2313 4326 2327 4333
rect 1797 4297 1813 4307
rect 1667 4293 1680 4297
rect 1800 4293 1813 4297
rect 2337 4303 2343 4333
rect 2307 4297 2343 4303
rect 3157 4307 3163 4333
rect 3277 4307 3283 4333
rect 3157 4297 3173 4307
rect 3160 4293 3173 4297
rect 3267 4297 3283 4307
rect 3267 4293 3280 4297
rect 3397 4287 3403 4333
rect 3537 4307 3543 4337
rect 3667 4343 3680 4347
rect 3667 4333 3683 4343
rect 3537 4297 3553 4307
rect 3540 4293 3553 4297
rect 3677 4303 3683 4333
rect 4517 4307 4523 4357
rect 5027 4357 5053 4363
rect 4780 4343 4793 4347
rect 4777 4333 4793 4343
rect 5427 4337 5453 4343
rect 4777 4307 4783 4333
rect 3677 4297 3703 4303
rect 4517 4297 4533 4307
rect 27 4277 113 4283
rect 1087 4277 1133 4283
rect 1280 4283 1293 4287
rect 1277 4273 1293 4283
rect 3247 4277 3273 4283
rect 3607 4277 3659 4283
rect 3697 4283 3703 4297
rect 4520 4293 4533 4297
rect 4777 4297 4793 4307
rect 4780 4293 4793 4297
rect 3697 4277 3733 4283
rect 1277 4263 1283 4273
rect 1247 4257 1283 4263
rect 3697 4263 3703 4277
rect 3627 4257 3703 4263
rect 4087 4237 4113 4243
rect -63 4162 30 4178
rect -63 3658 -3 4162
rect 4407 4117 4433 4123
rect 3187 4097 3273 4103
rect 3587 4097 3613 4103
rect 567 4077 593 4083
rect 2807 4077 2873 4083
rect 3077 4077 3133 4083
rect 67 4057 133 4063
rect 967 4057 1013 4063
rect 1127 4057 1153 4063
rect 1240 4043 1253 4047
rect 1237 4033 1253 4043
rect 1640 4043 1653 4047
rect 1637 4033 1653 4043
rect 2367 4037 2403 4043
rect 1237 3987 1243 4033
rect 1637 4007 1643 4033
rect 1627 3997 1643 4007
rect 2397 4007 2403 4037
rect 2487 4043 2500 4047
rect 2820 4043 2833 4047
rect 2487 4033 2503 4043
rect 2497 4007 2503 4033
rect 2817 4033 2833 4043
rect 2947 4043 2960 4047
rect 3077 4043 3083 4077
rect 3267 4077 3293 4083
rect 5007 4077 5073 4083
rect 3107 4057 3133 4063
rect 3207 4057 3313 4063
rect 3547 4057 3603 4063
rect 3240 4043 3253 4047
rect 2947 4033 2963 4043
rect 3077 4037 3103 4043
rect 2817 4007 2823 4033
rect 2957 4007 2963 4033
rect 2397 3997 2413 4007
rect 1627 3993 1640 3997
rect 2400 3993 2413 3997
rect 2497 3997 2513 4007
rect 2500 3993 2513 3997
rect 2807 3997 2823 4007
rect 2807 3993 2820 3997
rect 2947 3997 2963 4007
rect 3097 4007 3103 4037
rect 3237 4033 3253 4043
rect 3380 4043 3393 4047
rect 3377 4033 3393 4043
rect 3597 4043 3603 4057
rect 4727 4057 4833 4063
rect 5041 4057 5093 4063
rect 3760 4043 3773 4047
rect 3597 4037 3623 4043
rect 3097 3997 3113 4007
rect 2947 3993 2960 3997
rect 3100 3993 3113 3997
rect 3237 4003 3243 4033
rect 3377 4007 3383 4033
rect 3207 3997 3243 4003
rect 3367 3997 3383 4007
rect 3617 4007 3623 4037
rect 3757 4033 3773 4043
rect 3880 4043 3893 4047
rect 3877 4033 3893 4043
rect 4007 4043 4020 4047
rect 4160 4043 4173 4047
rect 4007 4033 4023 4043
rect 3757 4007 3763 4033
rect 3877 4007 3883 4033
rect 4017 4007 4023 4033
rect 4157 4033 4173 4043
rect 4420 4043 4433 4047
rect 4417 4033 4433 4043
rect 4627 4043 4640 4047
rect 4627 4033 4643 4043
rect 5607 4043 5620 4047
rect 5607 4033 5623 4043
rect 4157 4007 4163 4033
rect 3617 3997 3633 4007
rect 3367 3993 3380 3997
rect 3620 3993 3633 3997
rect 3747 3997 3763 4007
rect 3747 3993 3760 3997
rect 3867 3997 3883 4007
rect 3867 3993 3880 3997
rect 4007 3997 4023 4007
rect 4007 3993 4020 3997
rect 4147 3997 4163 4007
rect 4417 4007 4423 4033
rect 4637 4007 4643 4033
rect 5617 4007 5623 4033
rect 4417 3997 4433 4007
rect 4147 3993 4160 3997
rect 4420 3993 4433 3997
rect 4637 3997 4653 4007
rect 4640 3993 4653 3997
rect 5617 3997 5633 4007
rect 5620 3993 5633 3997
rect 4593 3969 4607 3973
rect 4593 3963 4633 3969
rect 5823 3918 5883 4422
rect 5790 3902 5883 3918
rect 3187 3876 3223 3882
rect 287 3853 293 3867
rect 1767 3837 1813 3843
rect 407 3823 420 3827
rect 1080 3823 1093 3827
rect 407 3813 423 3823
rect 417 3787 423 3813
rect 1077 3813 1093 3823
rect 1607 3817 1633 3823
rect 2920 3823 2933 3827
rect 2917 3813 2933 3823
rect 1077 3787 1083 3813
rect 2917 3787 2923 3813
rect 417 3777 433 3787
rect 420 3773 433 3777
rect 1077 3777 1093 3787
rect 1080 3773 1093 3777
rect 2917 3777 2933 3787
rect 2920 3773 2933 3777
rect 647 3757 713 3763
rect 3217 3763 3223 3876
rect 4487 3837 4533 3843
rect 3340 3823 3353 3827
rect 3337 3813 3353 3823
rect 4187 3823 4200 3827
rect 4640 3823 4653 3827
rect 4187 3813 4203 3823
rect 3337 3787 3343 3813
rect 3337 3777 3353 3787
rect 3340 3773 3353 3777
rect 4197 3783 4203 3813
rect 4637 3813 4653 3823
rect 5027 3823 5040 3827
rect 5180 3823 5193 3827
rect 5027 3813 5043 3823
rect 4637 3787 4643 3813
rect 4177 3777 4203 3783
rect 4177 3767 4183 3777
rect 4627 3777 4643 3787
rect 5037 3787 5043 3813
rect 5177 3813 5193 3823
rect 5720 3823 5733 3827
rect 5717 3813 5733 3823
rect 5177 3787 5183 3813
rect 5037 3777 5053 3787
rect 4627 3773 4640 3777
rect 5040 3773 5053 3777
rect 5167 3777 5183 3787
rect 5717 3787 5723 3813
rect 5717 3777 5733 3787
rect 5167 3773 5180 3777
rect 5720 3773 5733 3777
rect 4160 3765 4183 3767
rect 3217 3757 3253 3763
rect 4167 3757 4183 3765
rect 4167 3753 4180 3757
rect 4907 3757 4973 3763
rect 5567 3757 5653 3763
rect 5587 3737 5633 3743
rect -63 3642 30 3658
rect -63 3138 -3 3642
rect 247 3537 313 3543
rect 1427 3537 1473 3543
rect 3587 3537 3623 3543
rect 1547 3523 1560 3527
rect 1547 3513 1563 3523
rect 1557 3487 1563 3513
rect 1547 3477 1563 3487
rect 2337 3483 2343 3533
rect 2447 3523 2460 3527
rect 3617 3523 3623 3537
rect 4207 3537 4233 3543
rect 5097 3537 5153 3543
rect 2447 3513 2463 3523
rect 3617 3517 3643 3523
rect 2457 3487 2463 3513
rect 3637 3487 3643 3517
rect 4567 3523 4580 3527
rect 4960 3523 4973 3527
rect 4567 3513 4583 3523
rect 3813 3503 3827 3513
rect 3787 3500 3827 3503
rect 3787 3497 3823 3500
rect 4577 3487 4583 3513
rect 2317 3480 2343 3483
rect 2313 3477 2343 3480
rect 1547 3473 1560 3477
rect 2313 3467 2327 3477
rect 2447 3477 2463 3487
rect 2447 3473 2460 3477
rect 3627 3477 3643 3487
rect 3627 3473 3640 3477
rect 4567 3477 4583 3487
rect 4957 3513 4973 3523
rect 4957 3483 4963 3513
rect 5097 3487 5103 3537
rect 5447 3537 5513 3543
rect 5240 3523 5253 3527
rect 5237 3513 5253 3523
rect 5380 3523 5393 3527
rect 5377 3513 5393 3523
rect 5520 3523 5533 3527
rect 5517 3513 5533 3523
rect 5660 3523 5673 3527
rect 5657 3513 5673 3523
rect 5237 3487 5243 3513
rect 4957 3480 4983 3483
rect 4957 3477 4987 3480
rect 5097 3477 5113 3487
rect 4567 3473 4580 3477
rect 4973 3467 4987 3477
rect 5100 3473 5113 3477
rect 5227 3477 5243 3487
rect 5377 3487 5383 3513
rect 5517 3487 5523 3513
rect 5377 3477 5393 3487
rect 5227 3473 5240 3477
rect 5380 3473 5393 3477
rect 5507 3477 5523 3487
rect 5657 3487 5663 3513
rect 5657 3477 5673 3487
rect 5507 3473 5520 3477
rect 5660 3473 5673 3477
rect 3107 3457 3133 3463
rect 5823 3398 5883 3902
rect 5790 3382 5883 3398
rect 1087 3337 1113 3343
rect 1307 3337 1353 3343
rect 1487 3323 1500 3327
rect 1487 3313 1503 3323
rect 1100 3303 1113 3307
rect 1097 3293 1113 3303
rect 1497 3303 1503 3313
rect 4527 3317 4603 3323
rect 2860 3303 2873 3307
rect 1497 3297 1523 3303
rect 1097 3267 1103 3293
rect 1097 3257 1113 3267
rect 1100 3253 1113 3257
rect 1087 3237 1153 3243
rect 1517 3243 1523 3297
rect 2857 3293 2873 3303
rect 2980 3303 2993 3307
rect 2977 3293 2993 3303
rect 3353 3303 3367 3313
rect 3520 3303 3533 3307
rect 3353 3300 3383 3303
rect 3357 3297 3383 3300
rect 2857 3267 2863 3293
rect 2847 3257 2863 3267
rect 2977 3263 2983 3293
rect 2957 3257 2983 3263
rect 3377 3263 3383 3297
rect 3517 3293 3533 3303
rect 3767 3303 3780 3307
rect 3767 3293 3783 3303
rect 4447 3303 4460 3307
rect 4447 3293 4463 3303
rect 3517 3267 3523 3293
rect 3377 3257 3403 3263
rect 2847 3253 2860 3257
rect 1517 3237 1553 3243
rect 2957 3227 2963 3257
rect 2987 3237 3013 3243
rect 3397 3243 3403 3257
rect 3507 3257 3523 3267
rect 3777 3267 3783 3293
rect 4457 3267 4463 3293
rect 4597 3267 4603 3317
rect 5287 3317 5333 3323
rect 4740 3303 4753 3307
rect 3777 3257 3793 3267
rect 3507 3253 3520 3257
rect 3780 3253 3793 3257
rect 4457 3257 4473 3267
rect 4460 3253 4473 3257
rect 4587 3257 4603 3267
rect 4737 3293 4753 3303
rect 4893 3303 4907 3313
rect 4877 3300 4907 3303
rect 4877 3297 4903 3300
rect 4737 3263 4743 3293
rect 4877 3267 4883 3297
rect 5147 3303 5160 3307
rect 5700 3303 5713 3307
rect 5147 3293 5163 3303
rect 5157 3267 5163 3293
rect 4737 3257 4763 3263
rect 4877 3257 4893 3267
rect 4587 3253 4600 3257
rect 4757 3247 4763 3257
rect 4880 3253 4893 3257
rect 5147 3257 5163 3267
rect 5697 3293 5713 3303
rect 5697 3267 5703 3293
rect 5697 3257 5713 3267
rect 5147 3253 5160 3257
rect 5700 3253 5713 3257
rect 3397 3237 3433 3243
rect 3627 3237 3693 3243
rect 4567 3237 4673 3243
rect 4767 3237 4813 3243
rect 5647 3237 5673 3243
rect 2957 3226 2980 3227
rect 2957 3217 2973 3226
rect 2960 3213 2973 3217
rect -63 3122 30 3138
rect -63 2618 -3 3122
rect 1287 3017 1333 3023
rect 3367 3017 3393 3023
rect 3417 3017 3453 3023
rect 1507 3003 1520 3007
rect 2760 3003 2773 3007
rect 1507 2993 1523 3003
rect 1517 2967 1523 2993
rect 1507 2957 1523 2967
rect 2757 2993 2773 3003
rect 3417 3003 3423 3017
rect 4007 3017 4053 3023
rect 4147 3017 4213 3023
rect 3397 2997 3423 3003
rect 2757 2967 2763 2993
rect 3397 2967 3403 2997
rect 3527 3003 3540 3007
rect 4160 3003 4173 3007
rect 3527 2993 3543 3003
rect 3537 2967 3543 2993
rect 2757 2957 2773 2967
rect 1507 2953 1520 2957
rect 2760 2953 2773 2957
rect 3387 2957 3403 2967
rect 3387 2953 3400 2957
rect 3527 2957 3543 2967
rect 4157 2993 4173 3003
rect 4867 3003 4880 3007
rect 4867 3000 4883 3003
rect 4867 2993 4887 3000
rect 5507 3003 5520 3007
rect 5507 2993 5523 3003
rect 4157 2963 4163 2993
rect 4873 2986 4887 2993
rect 5517 2967 5523 2993
rect 4137 2960 4163 2963
rect 4133 2957 4163 2960
rect 3527 2953 3540 2957
rect 4133 2947 4147 2957
rect 307 2937 353 2943
rect 673 2903 687 2913
rect 673 2900 713 2903
rect 677 2897 713 2900
rect 5823 2878 5883 3382
rect 5790 2862 5883 2878
rect 407 2797 433 2803
rect 1227 2797 1253 2803
rect 4407 2797 4433 2803
rect 5047 2797 5113 2803
rect 647 2773 663 2787
rect 4807 2777 4833 2783
rect 4960 2783 4973 2787
rect 4957 2773 4973 2783
rect 5060 2783 5073 2787
rect 5057 2773 5073 2783
rect 5460 2783 5473 2787
rect 5457 2773 5473 2783
rect 5587 2783 5600 2787
rect 5587 2773 5603 2783
rect 657 2747 663 2773
rect 4957 2747 4963 2773
rect 5057 2747 5063 2773
rect 647 2737 663 2747
rect 647 2733 660 2737
rect 4947 2737 4963 2747
rect 4947 2733 4960 2737
rect 5047 2737 5063 2747
rect 5457 2747 5463 2773
rect 5597 2747 5603 2773
rect 5457 2737 5473 2747
rect 5047 2733 5060 2737
rect 5460 2733 5473 2737
rect 5587 2737 5603 2747
rect 5587 2733 5600 2737
rect 907 2717 1013 2723
rect 3667 2717 3693 2723
rect 5447 2717 5533 2723
rect 5627 2717 5673 2723
rect -63 2602 30 2618
rect -63 2098 -3 2602
rect 347 2497 373 2503
rect 1567 2497 1593 2503
rect 5700 2483 5713 2487
rect 5697 2473 5713 2483
rect 5787 2483 5800 2487
rect 5787 2473 5803 2483
rect 5697 2447 5703 2473
rect 5797 2447 5803 2473
rect 5697 2437 5713 2447
rect 5700 2433 5713 2437
rect 5787 2437 5803 2447
rect 5787 2433 5800 2437
rect 2080 2386 2093 2387
rect 2087 2373 2093 2386
rect 5823 2358 5883 2862
rect 5790 2342 5883 2358
rect 787 2197 813 2203
rect 1387 2197 1433 2203
rect 1737 2206 1743 2273
rect 3367 2263 3380 2267
rect 3367 2253 3383 2263
rect 4247 2263 4260 2267
rect 4247 2253 4263 2263
rect 3377 2227 3383 2253
rect 3377 2217 3393 2227
rect 3380 2213 3393 2217
rect 4257 2206 4263 2253
rect -63 2082 30 2098
rect -63 1578 -3 2082
rect 847 1963 860 1967
rect 847 1953 863 1963
rect 967 1963 980 1967
rect 967 1953 983 1963
rect 2887 1963 2900 1967
rect 2887 1953 2903 1963
rect 3127 1963 3140 1967
rect 3127 1953 3143 1963
rect 5447 1963 5460 1967
rect 5447 1953 5463 1963
rect 857 1927 863 1953
rect 977 1927 983 1953
rect 857 1917 873 1927
rect 860 1913 873 1917
rect 967 1917 983 1927
rect 2897 1923 2903 1953
rect 3137 1927 3143 1953
rect 2897 1917 2933 1923
rect 967 1913 980 1917
rect 3137 1917 3153 1927
rect 3140 1913 3153 1917
rect 5457 1923 5463 1953
rect 5457 1920 5483 1923
rect 5457 1917 5487 1920
rect 5473 1907 5487 1917
rect 4527 1897 4573 1903
rect 5823 1838 5883 2342
rect 5790 1822 5883 1838
rect 887 1757 913 1763
rect 1467 1757 1493 1763
rect 400 1743 413 1747
rect 397 1733 413 1743
rect 4187 1743 4200 1747
rect 4187 1733 4203 1743
rect 4327 1743 4340 1747
rect 4920 1743 4933 1747
rect 4327 1733 4343 1743
rect 397 1723 403 1733
rect 387 1717 403 1723
rect 4197 1707 4203 1733
rect 4197 1697 4213 1707
rect 4200 1693 4213 1697
rect 4337 1703 4343 1733
rect 4917 1733 4933 1743
rect 4917 1707 4923 1733
rect 4317 1697 4343 1703
rect 1087 1677 1153 1683
rect 2227 1677 2293 1683
rect 4317 1683 4323 1697
rect 4907 1697 4923 1707
rect 4907 1693 4920 1697
rect 4287 1677 4323 1683
rect -63 1562 30 1578
rect -63 1058 -3 1562
rect 2967 1457 3003 1463
rect 1260 1443 1273 1447
rect 1257 1433 1273 1443
rect 2997 1443 3003 1457
rect 5127 1457 5173 1463
rect 2997 1437 3023 1443
rect 1257 1407 1263 1433
rect 3017 1407 3023 1437
rect 5247 1443 5260 1447
rect 5247 1433 5263 1443
rect 5257 1407 5263 1433
rect 1247 1397 1263 1407
rect 1247 1393 1260 1397
rect 3007 1397 3023 1407
rect 3007 1393 3020 1397
rect 5247 1397 5263 1407
rect 5247 1393 5260 1397
rect 1507 1377 1553 1383
rect 5823 1318 5883 1822
rect 5790 1302 5883 1318
rect 367 1257 393 1263
rect 3307 1237 3333 1243
rect 267 1223 280 1227
rect 1540 1223 1553 1227
rect 267 1213 283 1223
rect 277 1187 283 1213
rect 1537 1213 1553 1223
rect 2787 1223 2800 1227
rect 2787 1213 2803 1223
rect 3647 1223 3660 1227
rect 4280 1223 4293 1227
rect 3647 1213 3663 1223
rect 1537 1187 1543 1213
rect 277 1177 293 1187
rect 280 1173 293 1177
rect 1527 1177 1543 1187
rect 1527 1173 1540 1177
rect 2797 1167 2803 1213
rect 3657 1187 3663 1213
rect 4277 1213 4293 1223
rect 5127 1223 5140 1227
rect 5127 1213 5143 1223
rect 4277 1187 4283 1213
rect 5137 1187 5143 1213
rect 3657 1177 3673 1187
rect 3660 1173 3673 1177
rect 4277 1177 4293 1187
rect 4280 1173 4293 1177
rect 5127 1177 5143 1187
rect 5127 1173 5140 1177
rect -63 1042 30 1058
rect -63 538 -3 1042
rect 3487 937 3553 943
rect 287 917 313 923
rect 3517 887 3523 937
rect 4227 937 4333 943
rect 3900 923 3913 927
rect 3897 913 3913 923
rect 4140 923 4153 927
rect 4137 913 4153 923
rect 3897 887 3903 913
rect 4137 887 4143 913
rect 3507 877 3523 887
rect 3507 873 3520 877
rect 3887 877 3903 887
rect 3887 873 3900 877
rect 4127 877 4143 887
rect 4127 873 4140 877
rect 5823 798 5883 1302
rect 5790 782 5883 798
rect 1927 703 1940 707
rect 1927 693 1943 703
rect 2047 703 2060 707
rect 2047 693 2063 703
rect 5407 697 5433 703
rect 1937 663 1943 693
rect 2057 663 2063 693
rect 1937 660 1963 663
rect 1937 657 1967 660
rect 1953 647 1967 657
rect 627 637 673 643
rect 2037 657 2063 663
rect 2037 627 2043 657
rect 2067 637 2113 643
rect 3667 637 3713 643
rect 4307 637 4373 643
rect 4587 637 4633 643
rect 2037 626 2060 627
rect 2037 617 2053 626
rect 2040 613 2053 617
rect -63 522 30 538
rect -63 18 -3 522
rect 1247 417 1273 423
rect 3307 417 3333 423
rect 4067 417 4133 423
rect 2040 403 2053 407
rect 2037 393 2053 403
rect 2287 403 2300 407
rect 2287 393 2303 403
rect 2787 403 2800 407
rect 2787 400 2803 403
rect 2787 393 2807 400
rect 3207 403 3220 407
rect 3207 393 3223 403
rect 2037 367 2043 393
rect 2297 367 2303 393
rect 2793 386 2807 393
rect 3217 367 3223 393
rect 2037 357 2053 367
rect 2040 353 2053 357
rect 2297 357 2313 367
rect 2300 353 2313 357
rect 3207 357 3223 367
rect 3207 353 3220 357
rect 867 337 933 343
rect 2187 337 2213 343
rect 5823 278 5883 782
rect 5790 262 5883 278
rect 4447 197 4493 203
rect 3207 183 3220 187
rect 3207 180 3223 183
rect 3207 173 3227 180
rect 3213 166 3227 173
rect 4747 77 4773 83
rect -63 2 30 18
rect 5823 2 5883 262
<< m2contact >>
rect 3093 5433 3107 5447
rect 3133 5433 3147 5447
rect 3673 5433 3687 5447
rect 3713 5433 3727 5447
rect 1493 5393 1507 5407
rect 1533 5393 1547 5407
rect 1773 5393 1787 5407
rect 2953 5393 2967 5407
rect 1733 5373 1747 5387
rect 2573 5373 2587 5387
rect 2753 5373 2767 5387
rect 2613 5333 2627 5347
rect 2713 5333 2727 5347
rect 3133 5373 3147 5387
rect 3473 5393 3487 5407
rect 3633 5393 3647 5407
rect 3773 5393 3787 5407
rect 3033 5333 3047 5347
rect 4053 5373 4067 5387
rect 5713 5373 5727 5387
rect 3373 5333 3387 5347
rect 4073 5332 4087 5346
rect 5753 5333 5767 5347
rect 2733 5313 2747 5327
rect 2773 5313 2787 5327
rect 2813 5311 2827 5325
rect 2913 5313 2927 5327
rect 3093 5313 3107 5327
rect 3233 5313 3247 5327
rect 3313 5313 3327 5327
rect 4713 5313 4727 5327
rect 4773 5313 4787 5327
rect 5413 5313 5427 5327
rect 5519 5313 5533 5327
rect 3073 5293 3087 5307
rect 3113 5293 3127 5307
rect 2733 5273 2747 5287
rect 2773 5273 2787 5287
rect 2853 5173 2867 5187
rect 2893 5173 2907 5187
rect 3293 5173 3307 5187
rect 3353 5173 3367 5187
rect 2633 5113 2647 5127
rect 2673 5113 2687 5127
rect 3553 5113 3567 5127
rect 3633 5113 3647 5127
rect 513 5093 527 5107
rect 633 5093 647 5107
rect 1993 5093 2007 5107
rect 2053 5093 2067 5107
rect 2553 5093 2567 5107
rect 2673 5092 2687 5106
rect 3253 5093 3267 5107
rect 3373 5093 3387 5107
rect 4127 5093 4141 5107
rect 4273 5093 4287 5107
rect 4413 5093 4427 5107
rect 4493 5093 4507 5107
rect 4873 5093 4887 5107
rect 4933 5093 4947 5107
rect 5053 5093 5067 5107
rect 5113 5093 5127 5107
rect 5173 5093 5187 5107
rect 853 5073 867 5087
rect 1953 5073 1967 5087
rect 2153 5073 2167 5087
rect 893 5033 907 5047
rect 533 5013 547 5027
rect 653 5013 667 5027
rect 1933 5012 1947 5026
rect 2613 5073 2627 5087
rect 2753 5072 2767 5086
rect 3633 5073 3647 5087
rect 3873 5073 3887 5087
rect 4313 5073 4327 5087
rect 4453 5073 4467 5087
rect 2573 5033 2587 5047
rect 2713 5033 2727 5047
rect 3633 5033 3647 5047
rect 3913 5033 3927 5047
rect 4313 5033 4327 5047
rect 5313 5073 5327 5087
rect 5633 5073 5647 5087
rect 5593 5053 5607 5067
rect 2213 5013 2227 5027
rect 2533 5013 2547 5027
rect 2613 5013 2627 5027
rect 3253 5013 3267 5027
rect 3313 5013 3327 5027
rect 4413 5013 4427 5027
rect 5193 5033 5207 5047
rect 5273 5033 5287 5047
rect 5613 5033 5627 5047
rect 5633 5013 5647 5027
rect 5593 4973 5607 4987
rect 5633 4973 5647 4987
rect 733 4853 747 4867
rect 2453 4853 2467 4867
rect 2693 4853 2707 4867
rect 2973 4853 2987 4867
rect 3933 4853 3947 4867
rect 4073 4853 4087 4867
rect 4173 4853 4187 4867
rect 713 4813 727 4827
rect 2673 4833 2687 4847
rect 2933 4813 2947 4827
rect 3893 4813 3907 4827
rect 4033 4813 4047 4827
rect 4173 4813 4187 4827
rect 4593 4853 4607 4867
rect 5233 4853 5247 4867
rect 5293 4853 5307 4867
rect 653 4793 667 4807
rect 773 4793 787 4807
rect 813 4793 827 4807
rect 893 4793 907 4807
rect 2413 4793 2427 4807
rect 3033 4793 3047 4807
rect 3173 4793 3187 4807
rect 3987 4793 4001 4807
rect 4073 4793 4087 4807
rect 5193 4813 5207 4827
rect 5473 4853 5487 4867
rect 5613 4853 5627 4867
rect 5333 4813 5347 4827
rect 5433 4813 5447 4827
rect 4633 4793 4647 4807
rect 5033 4793 5047 4807
rect 5073 4793 5087 4807
rect 5293 4793 5307 4807
rect 5393 4793 5407 4807
rect 5553 4793 5567 4807
rect 2833 4633 2847 4647
rect 2893 4633 2907 4647
rect 2813 4613 2827 4627
rect 2853 4613 2867 4627
rect 413 4573 427 4587
rect 453 4573 467 4587
rect 1053 4573 1067 4587
rect 1113 4573 1127 4587
rect 1753 4573 1767 4587
rect 1873 4573 1887 4587
rect 1913 4573 1927 4587
rect 2673 4573 2687 4587
rect 2893 4573 2907 4587
rect 1353 4553 1367 4567
rect 1793 4552 1807 4566
rect 1933 4553 1947 4567
rect 1393 4513 1407 4527
rect 1893 4513 1907 4527
rect 1333 4493 1347 4507
rect 1413 4493 1427 4507
rect 1773 4493 1787 4507
rect 1833 4493 1847 4507
rect 2933 4572 2947 4586
rect 3653 4573 3667 4587
rect 3753 4573 3767 4587
rect 3133 4553 3147 4567
rect 3613 4553 3627 4567
rect 2853 4533 2867 4547
rect 2833 4513 2847 4527
rect 3093 4513 3107 4527
rect 4393 4533 4407 4547
rect 3613 4513 3627 4527
rect 4553 4574 4567 4588
rect 4593 4573 4607 4587
rect 4653 4573 4667 4587
rect 4713 4553 4727 4567
rect 4753 4532 4767 4546
rect 2773 4493 2787 4507
rect 3233 4493 3247 4507
rect 3293 4493 3307 4507
rect 4033 4493 4047 4507
rect 4073 4493 4087 4507
rect 4413 4513 4427 4527
rect 4533 4513 4547 4527
rect 4373 4492 4387 4506
rect 4413 4473 4427 4487
rect 4613 4453 4627 4467
rect 4653 4453 4667 4467
rect 953 4353 967 4367
rect 1013 4353 1027 4367
rect 1353 4353 1367 4367
rect 1453 4353 1467 4367
rect 3513 4353 3527 4367
rect 4453 4354 4467 4368
rect 673 4333 687 4347
rect 1513 4333 1527 4347
rect 1693 4333 1707 4347
rect 1773 4333 1787 4347
rect 2293 4333 2307 4347
rect 2333 4333 2347 4347
rect 3153 4333 3167 4347
rect 3253 4333 3267 4347
rect 3373 4333 3387 4347
rect 673 4293 687 4307
rect 1513 4293 1527 4307
rect 1653 4293 1667 4307
rect 2313 4312 2327 4326
rect 1813 4293 1827 4307
rect 2293 4293 2307 4307
rect 3173 4293 3187 4307
rect 3253 4293 3267 4307
rect 3653 4333 3667 4347
rect 3553 4293 3567 4307
rect 5013 4352 5027 4366
rect 5053 4353 5067 4367
rect 4793 4333 4807 4347
rect 5413 4333 5427 4347
rect 5453 4332 5467 4346
rect 13 4273 27 4287
rect 113 4273 127 4287
rect 1073 4273 1087 4287
rect 1133 4273 1147 4287
rect 1293 4273 1307 4287
rect 3233 4273 3247 4287
rect 3273 4273 3287 4287
rect 3393 4273 3407 4287
rect 3593 4273 3607 4287
rect 3659 4273 3673 4287
rect 4533 4293 4547 4307
rect 4793 4293 4807 4307
rect 1233 4253 1247 4267
rect 3613 4253 3627 4267
rect 3733 4273 3747 4287
rect 4073 4232 4087 4246
rect 4113 4233 4127 4247
rect 4393 4113 4407 4127
rect 4433 4112 4447 4126
rect 3173 4093 3187 4107
rect 3273 4093 3287 4107
rect 3573 4093 3587 4107
rect 3613 4093 3627 4107
rect 553 4073 567 4087
rect 593 4073 607 4087
rect 2793 4073 2807 4087
rect 2873 4073 2887 4087
rect 53 4053 67 4067
rect 133 4053 147 4067
rect 953 4053 967 4067
rect 1013 4053 1027 4067
rect 1113 4053 1127 4067
rect 1153 4053 1167 4067
rect 1253 4033 1267 4047
rect 1653 4033 1667 4047
rect 2353 4033 2367 4047
rect 1613 3993 1627 4007
rect 2473 4033 2487 4047
rect 2833 4033 2847 4047
rect 2933 4033 2947 4047
rect 3133 4073 3147 4087
rect 3253 4073 3267 4087
rect 3293 4073 3307 4087
rect 4993 4073 5007 4087
rect 5073 4073 5087 4087
rect 3093 4053 3107 4067
rect 3133 4052 3147 4066
rect 3193 4053 3207 4067
rect 3313 4052 3327 4066
rect 3533 4053 3547 4067
rect 2413 3993 2427 4007
rect 2513 3993 2527 4007
rect 2793 3993 2807 4007
rect 2933 3993 2947 4007
rect 3253 4033 3267 4047
rect 3393 4033 3407 4047
rect 4713 4053 4727 4067
rect 4833 4053 4847 4067
rect 5027 4053 5041 4067
rect 5093 4053 5107 4067
rect 3113 3993 3127 4007
rect 3193 3993 3207 4007
rect 3353 3993 3367 4007
rect 3773 4033 3787 4047
rect 3893 4033 3907 4047
rect 3993 4033 4007 4047
rect 4173 4033 4187 4047
rect 4433 4033 4447 4047
rect 4613 4033 4627 4047
rect 5593 4033 5607 4047
rect 3633 3993 3647 4007
rect 3733 3993 3747 4007
rect 3853 3993 3867 4007
rect 3993 3993 4007 4007
rect 4133 3993 4147 4007
rect 4433 3993 4447 4007
rect 4653 3993 4667 4007
rect 5633 3993 5647 4007
rect 1233 3973 1247 3987
rect 4593 3973 4607 3987
rect 4633 3959 4647 3973
rect 3173 3871 3187 3885
rect 273 3853 287 3867
rect 293 3853 307 3867
rect 1753 3833 1767 3847
rect 1813 3833 1827 3847
rect 393 3813 407 3827
rect 1093 3813 1107 3827
rect 1593 3813 1607 3827
rect 1633 3813 1647 3827
rect 2933 3813 2947 3827
rect 433 3773 447 3787
rect 1093 3773 1107 3787
rect 2933 3773 2947 3787
rect 633 3753 647 3767
rect 713 3753 727 3767
rect 4473 3833 4487 3847
rect 4533 3833 4547 3847
rect 3353 3813 3367 3827
rect 4173 3813 4187 3827
rect 3353 3773 3367 3787
rect 4653 3813 4667 3827
rect 5013 3813 5027 3827
rect 4613 3773 4627 3787
rect 5193 3813 5207 3827
rect 5733 3813 5747 3827
rect 5053 3773 5067 3787
rect 5153 3773 5167 3787
rect 5733 3773 5747 3787
rect 3253 3751 3267 3765
rect 4153 3751 4167 3765
rect 4893 3753 4907 3767
rect 4973 3753 4987 3767
rect 5553 3753 5567 3767
rect 5653 3753 5667 3767
rect 5573 3733 5587 3747
rect 5633 3733 5647 3747
rect 233 3533 247 3547
rect 313 3533 327 3547
rect 1413 3533 1427 3547
rect 1473 3534 1487 3548
rect 2333 3533 2347 3547
rect 3573 3533 3587 3547
rect 1533 3513 1547 3527
rect 1533 3473 1547 3487
rect 2433 3513 2447 3527
rect 4193 3532 4207 3546
rect 4233 3533 4247 3547
rect 3813 3513 3827 3527
rect 4553 3513 4567 3527
rect 3773 3492 3787 3506
rect 2433 3473 2447 3487
rect 3613 3473 3627 3487
rect 4553 3473 4567 3487
rect 4973 3513 4987 3527
rect 5153 3533 5167 3547
rect 5433 3533 5447 3547
rect 5513 3533 5527 3547
rect 5253 3513 5267 3527
rect 5393 3513 5407 3527
rect 5533 3513 5547 3527
rect 5673 3513 5687 3527
rect 5113 3473 5127 3487
rect 5213 3473 5227 3487
rect 5393 3473 5407 3487
rect 5493 3473 5507 3487
rect 5673 3473 5687 3487
rect 2313 3453 2327 3467
rect 3093 3453 3107 3467
rect 3133 3453 3147 3467
rect 4973 3453 4987 3467
rect 1073 3333 1087 3347
rect 1113 3333 1127 3347
rect 1293 3333 1307 3347
rect 1353 3333 1367 3347
rect 1473 3313 1487 3327
rect 1113 3293 1127 3307
rect 3353 3313 3367 3327
rect 4513 3313 4527 3327
rect 1113 3253 1127 3267
rect 1073 3233 1087 3247
rect 1153 3233 1167 3247
rect 2873 3293 2887 3307
rect 2993 3293 3007 3307
rect 2833 3253 2847 3267
rect 3533 3293 3547 3307
rect 3753 3293 3767 3307
rect 4433 3293 4447 3307
rect 1553 3233 1567 3247
rect 2973 3233 2987 3247
rect 3013 3233 3027 3247
rect 3493 3253 3507 3267
rect 4893 3313 4907 3327
rect 5273 3313 5287 3327
rect 5333 3313 5347 3327
rect 3793 3253 3807 3267
rect 4473 3253 4487 3267
rect 4573 3253 4587 3267
rect 4753 3293 4767 3307
rect 5133 3293 5147 3307
rect 4893 3253 4907 3267
rect 5133 3253 5147 3267
rect 5713 3293 5727 3307
rect 5713 3253 5727 3267
rect 3433 3231 3447 3245
rect 3613 3233 3627 3247
rect 3693 3233 3707 3247
rect 4553 3233 4567 3247
rect 4673 3233 4687 3247
rect 4753 3233 4767 3247
rect 4813 3233 4827 3247
rect 5633 3233 5647 3247
rect 5673 3233 5687 3247
rect 2973 3212 2987 3226
rect 1273 3013 1287 3027
rect 1333 3013 1347 3027
rect 3353 3013 3367 3027
rect 3393 3013 3407 3027
rect 1493 2993 1507 3007
rect 1493 2953 1507 2967
rect 2773 2993 2787 3007
rect 3453 3013 3467 3027
rect 3993 3013 4007 3027
rect 4053 3013 4067 3027
rect 4133 3013 4147 3027
rect 4213 3014 4227 3028
rect 3513 2993 3527 3007
rect 2773 2953 2787 2967
rect 3373 2953 3387 2967
rect 3513 2953 3527 2967
rect 4173 2993 4187 3007
rect 4853 2993 4867 3007
rect 5493 2993 5507 3007
rect 4873 2972 4887 2986
rect 5513 2953 5527 2967
rect 293 2933 307 2947
rect 353 2933 367 2947
rect 4133 2933 4147 2947
rect 673 2913 687 2927
rect 713 2893 727 2907
rect 393 2792 407 2806
rect 433 2793 447 2807
rect 1213 2793 1227 2807
rect 1253 2793 1267 2807
rect 4393 2793 4407 2807
rect 4433 2793 4447 2807
rect 5033 2793 5047 2807
rect 5113 2793 5127 2807
rect 633 2773 647 2787
rect 4793 2773 4807 2787
rect 4833 2773 4847 2787
rect 4973 2773 4987 2787
rect 5073 2773 5087 2787
rect 5473 2773 5487 2787
rect 5573 2773 5587 2787
rect 633 2733 647 2747
rect 4933 2733 4947 2747
rect 5033 2733 5047 2747
rect 5473 2733 5487 2747
rect 5573 2733 5587 2747
rect 893 2713 907 2727
rect 1013 2711 1027 2725
rect 3653 2713 3667 2727
rect 3693 2713 3707 2727
rect 5433 2713 5447 2727
rect 5533 2713 5547 2727
rect 5613 2713 5627 2727
rect 5673 2713 5687 2727
rect 333 2493 347 2507
rect 373 2494 387 2508
rect 1553 2493 1567 2507
rect 1593 2493 1607 2507
rect 5713 2473 5727 2487
rect 5773 2473 5787 2487
rect 5713 2433 5727 2447
rect 5773 2433 5787 2447
rect 2073 2372 2087 2386
rect 2093 2373 2107 2387
rect 1733 2273 1747 2287
rect 773 2193 787 2207
rect 813 2193 827 2207
rect 1373 2193 1387 2207
rect 1433 2193 1447 2207
rect 3353 2253 3367 2267
rect 4233 2253 4247 2267
rect 3393 2213 3407 2227
rect 1733 2192 1747 2206
rect 4253 2192 4267 2206
rect 833 1953 847 1967
rect 953 1953 967 1967
rect 2873 1953 2887 1967
rect 3113 1953 3127 1967
rect 5433 1953 5447 1967
rect 873 1913 887 1927
rect 953 1913 967 1927
rect 2933 1913 2947 1927
rect 3153 1913 3167 1927
rect 4513 1893 4527 1907
rect 4573 1893 4587 1907
rect 5473 1893 5487 1907
rect 873 1753 887 1767
rect 913 1753 927 1767
rect 1453 1753 1467 1767
rect 1493 1753 1507 1767
rect 413 1733 427 1747
rect 4173 1733 4187 1747
rect 4313 1733 4327 1747
rect 373 1713 387 1727
rect 4213 1693 4227 1707
rect 4933 1733 4947 1747
rect 1073 1673 1087 1687
rect 1153 1673 1167 1687
rect 2213 1673 2227 1687
rect 2293 1673 2307 1687
rect 4273 1673 4287 1687
rect 4893 1693 4907 1707
rect 2953 1453 2967 1467
rect 1273 1433 1287 1447
rect 5113 1452 5127 1466
rect 5173 1453 5187 1467
rect 5233 1433 5247 1447
rect 1233 1393 1247 1407
rect 2993 1393 3007 1407
rect 5233 1393 5247 1407
rect 1493 1373 1507 1387
rect 1553 1373 1567 1387
rect 353 1253 367 1267
rect 393 1253 407 1267
rect 3293 1233 3307 1247
rect 3333 1233 3347 1247
rect 253 1213 267 1227
rect 1553 1213 1567 1227
rect 2773 1213 2787 1227
rect 3633 1213 3647 1227
rect 293 1173 307 1187
rect 1513 1173 1527 1187
rect 4293 1213 4307 1227
rect 5113 1213 5127 1227
rect 3673 1173 3687 1187
rect 4293 1173 4307 1187
rect 5113 1173 5127 1187
rect 2793 1153 2807 1167
rect 3473 933 3487 947
rect 273 913 287 927
rect 313 913 327 927
rect 3553 933 3567 947
rect 4213 933 4227 947
rect 4333 933 4347 947
rect 3913 913 3927 927
rect 4153 913 4167 927
rect 3493 873 3507 887
rect 3873 873 3887 887
rect 4113 873 4127 887
rect 1913 693 1927 707
rect 2033 693 2047 707
rect 5393 693 5407 707
rect 5433 693 5447 707
rect 613 633 627 647
rect 673 633 687 647
rect 1953 633 1967 647
rect 2053 633 2067 647
rect 2113 633 2127 647
rect 3653 633 3667 647
rect 3713 633 3727 647
rect 4293 633 4307 647
rect 4373 633 4387 647
rect 4573 633 4587 647
rect 4633 633 4647 647
rect 2053 612 2067 626
rect 1233 413 1247 427
rect 1273 413 1287 427
rect 3293 413 3307 427
rect 3333 413 3347 427
rect 4053 413 4067 427
rect 4133 413 4147 427
rect 2053 393 2067 407
rect 2273 393 2287 407
rect 2773 393 2787 407
rect 3193 393 3207 407
rect 2793 372 2807 386
rect 2053 353 2067 367
rect 2313 353 2327 367
rect 3193 353 3207 367
rect 853 333 867 347
rect 933 333 947 347
rect 2173 333 2187 347
rect 2213 333 2227 347
rect 4433 193 4447 207
rect 4493 194 4507 208
rect 3193 173 3207 187
rect 3213 152 3227 166
rect 4733 73 4747 87
rect 4773 72 4787 86
<< metal2 >>
rect 116 5376 123 5413
rect 256 5376 263 5413
rect 296 5387 303 5413
rect 416 5387 423 5413
rect 76 5076 83 5153
rect 96 5127 103 5343
rect 136 5340 163 5343
rect 136 5336 167 5340
rect 153 5327 167 5336
rect 176 5088 183 5373
rect 236 5287 243 5343
rect 316 5223 323 5373
rect 436 5346 443 5413
rect 536 5376 583 5383
rect 616 5376 623 5413
rect 396 5307 403 5343
rect 476 5307 483 5343
rect 516 5267 523 5343
rect 576 5327 583 5376
rect 736 5376 743 5413
rect 896 5376 903 5453
rect 1036 5376 1043 5413
rect 1176 5376 1183 5433
rect 1316 5388 1323 5453
rect 1496 5407 1503 5433
rect 316 5216 343 5223
rect 256 5107 263 5153
rect 276 5076 283 5193
rect 16 4287 23 4613
rect 36 4267 43 4893
rect 76 4856 83 4893
rect 96 4887 103 5043
rect 116 4856 123 4913
rect 156 4867 163 4953
rect 256 4927 263 5043
rect 256 4883 263 4913
rect 236 4876 263 4883
rect 56 4568 63 4813
rect 96 4707 103 4823
rect 136 4556 143 4613
rect 176 4587 183 4873
rect 236 4856 243 4876
rect 216 4707 223 4823
rect 296 4767 303 4813
rect 316 4807 323 5193
rect 336 5147 343 5216
rect 376 5107 383 5153
rect 376 5076 383 5093
rect 513 5088 527 5093
rect 356 4967 363 5043
rect 396 4947 403 5043
rect 353 4860 367 4873
rect 356 4856 363 4860
rect 396 4856 403 4893
rect 436 4867 443 4933
rect 456 4907 463 5074
rect 536 5040 543 5043
rect 533 5027 547 5040
rect 536 4856 543 4933
rect 576 4867 583 4893
rect 376 4820 383 4823
rect 373 4807 387 4820
rect 176 4526 183 4573
rect 256 4556 263 4753
rect 296 4568 303 4713
rect 456 4587 463 4853
rect 516 4787 523 4823
rect 596 4747 603 5293
rect 636 5187 643 5343
rect 696 5307 703 5374
rect 756 5340 763 5343
rect 753 5327 767 5340
rect 836 5343 843 5374
rect 836 5336 883 5343
rect 633 5080 647 5093
rect 636 5076 643 5080
rect 676 5076 683 5173
rect 776 5147 783 5273
rect 656 5027 663 5043
rect 656 4987 663 5013
rect 636 4856 643 4933
rect 676 4868 683 5013
rect 696 4887 703 5043
rect 736 4987 743 5133
rect 776 5076 783 5133
rect 816 5076 823 5173
rect 856 5087 863 5133
rect 876 5046 883 5313
rect 936 5076 943 5253
rect 976 5088 983 5113
rect 1116 5083 1123 5332
rect 1116 5076 1133 5083
rect 736 4867 743 4973
rect 756 4947 763 5033
rect 756 4867 763 4933
rect 796 4907 803 5043
rect 836 5007 843 5043
rect 836 4856 843 4993
rect 700 4823 713 4827
rect 656 4820 663 4823
rect 373 4560 387 4573
rect 413 4560 427 4573
rect 476 4567 483 4693
rect 536 4587 543 4613
rect 376 4556 383 4560
rect 416 4556 423 4560
rect 56 4347 63 4513
rect 76 4487 83 4523
rect 116 4363 123 4512
rect 96 4356 123 4363
rect 96 4336 103 4356
rect 133 4340 147 4353
rect 136 4336 143 4340
rect 116 4300 123 4303
rect 113 4287 127 4300
rect 56 3947 63 4053
rect 133 4040 147 4053
rect 176 4048 183 4512
rect 196 4347 203 4473
rect 236 4407 243 4523
rect 276 4487 283 4523
rect 213 4340 227 4353
rect 253 4340 267 4353
rect 216 4336 223 4340
rect 256 4336 263 4340
rect 136 4036 143 4040
rect 196 4027 203 4293
rect 236 4267 243 4303
rect 276 4036 283 4113
rect 156 3883 163 4003
rect 256 3947 263 4003
rect 156 3876 183 3883
rect 56 3647 63 3873
rect 96 3816 103 3873
rect 16 3527 23 3553
rect 16 3407 23 3473
rect 16 3327 23 3353
rect 36 3308 43 3593
rect 56 3523 63 3633
rect 76 3607 83 3783
rect 96 3567 103 3613
rect 56 3516 83 3523
rect 113 3520 127 3533
rect 116 3516 123 3520
rect 156 3347 163 3853
rect 176 3786 183 3876
rect 267 3853 273 3867
rect 213 3820 227 3833
rect 216 3816 223 3820
rect 176 3567 183 3772
rect 233 3547 247 3553
rect 236 3516 243 3533
rect 276 3528 283 3832
rect 296 3823 303 3853
rect 316 3847 323 4393
rect 336 4348 343 4553
rect 476 4523 483 4553
rect 396 4347 403 4523
rect 436 4516 483 4523
rect 536 4520 543 4523
rect 533 4507 547 4520
rect 576 4507 583 4573
rect 596 4407 603 4653
rect 616 4487 623 4813
rect 653 4807 667 4820
rect 696 4816 713 4823
rect 700 4813 713 4816
rect 736 4627 743 4832
rect 773 4807 787 4812
rect 816 4807 823 4823
rect 796 4796 813 4803
rect 756 4587 763 4773
rect 736 4556 763 4563
rect 736 4427 743 4493
rect 756 4467 763 4556
rect 396 4063 403 4293
rect 416 4067 423 4353
rect 453 4340 467 4353
rect 456 4336 463 4340
rect 556 4306 563 4393
rect 776 4387 783 4613
rect 796 4547 803 4796
rect 816 4587 823 4733
rect 836 4727 843 4793
rect 876 4667 883 4853
rect 896 4807 903 5033
rect 956 4947 963 5043
rect 1016 5007 1023 5073
rect 1096 5036 1123 5043
rect 1057 5013 1064 5032
rect 1057 5006 1103 5013
rect 1096 4896 1103 5006
rect 1116 4987 1123 5036
rect 1136 4947 1143 5074
rect 1196 4987 1203 5043
rect 1236 5040 1263 5043
rect 1236 5036 1267 5040
rect 1253 5027 1267 5036
rect 1276 5007 1283 5074
rect 996 4823 1003 4873
rect 1047 4856 1063 4863
rect 916 4687 923 4823
rect 976 4816 1003 4823
rect 1036 4727 1043 4854
rect 1176 4823 1183 4873
rect 1256 4856 1263 4933
rect 1296 4867 1303 5153
rect 1316 5087 1323 5374
rect 1516 5376 1523 5413
rect 1536 5407 1543 5433
rect 1656 5376 1663 5413
rect 1736 5387 1743 5433
rect 1456 5346 1463 5373
rect 1376 5323 1383 5343
rect 1367 5316 1383 5323
rect 1356 5076 1363 5313
rect 1416 5127 1423 5332
rect 1496 5287 1503 5332
rect 1336 4967 1343 5043
rect 1156 4816 1183 4823
rect 1196 4807 1203 4853
rect 1316 4826 1323 4913
rect 1376 4887 1383 5043
rect 1416 5027 1423 5113
rect 1456 5088 1463 5213
rect 1516 5167 1523 5313
rect 1536 5247 1543 5343
rect 1576 5207 1583 5333
rect 1536 5047 1543 5193
rect 1576 5076 1583 5193
rect 1596 5103 1603 5373
rect 1756 5346 1763 5413
rect 1773 5388 1787 5393
rect 1816 5376 1823 5453
rect 1856 5376 1863 5413
rect 1936 5388 1943 5433
rect 2036 5346 2043 5453
rect 2096 5376 2103 5433
rect 2256 5376 2263 5413
rect 2396 5376 2403 5413
rect 2576 5387 2583 5453
rect 1636 5247 1643 5343
rect 1676 5287 1683 5343
rect 1836 5287 1843 5343
rect 1956 5323 1963 5343
rect 2056 5343 2063 5373
rect 2196 5346 2203 5373
rect 2056 5336 2083 5343
rect 1936 5320 1963 5323
rect 1936 5316 1967 5320
rect 1936 5267 1943 5316
rect 1953 5307 1967 5316
rect 1596 5096 1623 5103
rect 1616 5076 1623 5096
rect 1656 5087 1663 5173
rect 1476 5040 1483 5043
rect 1376 4856 1383 4873
rect 1236 4767 1243 4823
rect 1356 4787 1363 4823
rect 1256 4747 1263 4773
rect 916 4556 943 4563
rect 796 4516 823 4523
rect 796 4427 803 4516
rect 936 4487 943 4556
rect 996 4556 1003 4593
rect 1053 4587 1067 4593
rect 956 4443 963 4554
rect 1056 4520 1063 4523
rect 1053 4507 1067 4520
rect 916 4436 963 4443
rect 673 4347 687 4353
rect 476 4267 483 4303
rect 376 4056 403 4063
rect 376 4036 383 4056
rect 436 4043 443 4113
rect 496 4063 503 4273
rect 556 4087 563 4292
rect 616 4267 623 4303
rect 696 4306 703 4373
rect 916 4348 923 4436
rect 956 4367 963 4413
rect 616 4147 623 4253
rect 496 4056 523 4063
rect 416 4036 463 4043
rect 516 4036 523 4056
rect 553 4040 567 4052
rect 556 4036 563 4040
rect 356 3887 363 4003
rect 396 3967 403 3992
rect 296 3816 323 3823
rect 396 3827 403 3913
rect 436 3828 443 3993
rect 456 3927 463 4036
rect 496 3967 503 4003
rect 536 4000 543 4003
rect 533 3987 547 4000
rect 416 3816 433 3823
rect 376 3776 403 3783
rect 313 3520 327 3533
rect 316 3516 323 3520
rect 356 3516 363 3633
rect 216 3447 223 3483
rect 16 3127 23 3273
rect 36 3103 43 3233
rect 16 3096 43 3103
rect 16 2627 23 3096
rect 56 3087 63 3333
rect 196 3263 203 3333
rect 176 3256 203 3263
rect 216 3107 223 3393
rect 256 3347 263 3433
rect 256 3296 263 3333
rect 336 3303 343 3483
rect 396 3467 403 3776
rect 416 3587 423 3816
rect 487 3818 523 3825
rect 447 3783 460 3787
rect 447 3776 463 3783
rect 496 3780 503 3783
rect 447 3773 460 3776
rect 493 3767 507 3780
rect 476 3528 483 3573
rect 336 3296 363 3303
rect 76 2996 83 3033
rect 96 2827 103 2963
rect 136 2927 143 2963
rect 156 2827 163 2953
rect 136 2787 143 2813
rect 176 2783 183 3073
rect 213 3023 227 3033
rect 236 3023 243 3073
rect 213 3020 243 3023
rect 216 3016 243 3020
rect 216 3008 223 3016
rect 256 2996 263 3133
rect 276 3008 283 3263
rect 236 2927 243 2963
rect 296 2947 303 3033
rect 336 2996 343 3193
rect 376 3047 383 3263
rect 436 3207 443 3453
rect 456 3308 463 3483
rect 516 3308 523 3818
rect 536 3786 543 3853
rect 576 3816 583 3913
rect 596 3887 603 4073
rect 616 3867 623 4073
rect 656 4036 663 4133
rect 676 4087 683 4293
rect 696 4107 703 4292
rect 756 4283 763 4303
rect 756 4276 783 4283
rect 716 4067 723 4233
rect 776 4227 783 4276
rect 796 4187 803 4303
rect 836 4203 843 4334
rect 836 4196 863 4203
rect 676 3867 683 4003
rect 716 3816 723 4053
rect 776 4036 783 4093
rect 756 4000 763 4003
rect 753 3987 767 4000
rect 796 3967 803 4003
rect 796 3887 803 3953
rect 756 3827 763 3873
rect 836 3867 843 3993
rect 856 3927 863 4196
rect 876 4107 883 4273
rect 896 4227 903 4303
rect 896 4127 903 4213
rect 916 4187 923 4213
rect 876 4047 883 4093
rect 936 4063 943 4293
rect 956 4187 963 4353
rect 1013 4340 1027 4353
rect 1016 4336 1023 4340
rect 1056 4336 1063 4373
rect 1096 4343 1103 4573
rect 1116 4527 1123 4573
rect 1156 4568 1163 4713
rect 1196 4556 1203 4593
rect 1156 4348 1163 4473
rect 1216 4447 1223 4523
rect 1256 4503 1263 4633
rect 1293 4560 1307 4573
rect 1296 4556 1303 4560
rect 1356 4567 1363 4752
rect 1436 4687 1443 5033
rect 1473 5027 1487 5040
rect 1516 4947 1523 5033
rect 1676 5043 1683 5133
rect 1716 5076 1723 5133
rect 1876 5076 1883 5113
rect 1916 5087 1923 5133
rect 1676 5036 1703 5043
rect 1736 5040 1743 5043
rect 1576 4907 1583 4953
rect 1596 4827 1603 4993
rect 1456 4747 1463 4812
rect 1256 4496 1303 4503
rect 1096 4336 1123 4343
rect 1036 4247 1043 4303
rect 1076 4300 1083 4303
rect 1073 4287 1087 4300
rect 1036 4147 1043 4212
rect 927 4056 943 4063
rect 913 4040 927 4053
rect 953 4040 967 4053
rect 976 4047 983 4113
rect 916 4036 923 4040
rect 956 4036 963 4040
rect 936 3967 943 4003
rect 856 3816 863 3873
rect 636 3780 643 3783
rect 633 3767 647 3780
rect 676 3767 683 3793
rect 736 3767 743 3783
rect 776 3767 783 3813
rect 916 3787 923 3913
rect 956 3828 963 3853
rect 976 3843 983 3993
rect 996 3947 1003 4053
rect 1013 4047 1027 4053
rect 1036 4036 1043 4133
rect 1116 4067 1123 4336
rect 1196 4336 1203 4373
rect 1256 4306 1263 4453
rect 1296 4363 1303 4496
rect 1336 4387 1343 4493
rect 1356 4487 1363 4513
rect 1376 4367 1383 4673
rect 1396 4587 1403 4673
rect 1456 4556 1463 4733
rect 1476 4627 1483 4823
rect 1556 4787 1563 4823
rect 1476 4568 1483 4613
rect 1432 4527 1446 4532
rect 1396 4487 1403 4513
rect 1427 4505 1440 4507
rect 1427 4493 1433 4505
rect 1496 4467 1503 4653
rect 1296 4356 1323 4363
rect 1316 4348 1323 4356
rect 1353 4340 1367 4353
rect 1356 4336 1363 4340
rect 1133 4287 1147 4293
rect 1176 4227 1183 4303
rect 1296 4300 1303 4303
rect 1293 4287 1307 4300
rect 1236 4183 1243 4253
rect 1236 4176 1263 4183
rect 1153 4040 1167 4053
rect 1156 4036 1163 4040
rect 1236 4003 1243 4133
rect 1256 4127 1263 4176
rect 1256 4047 1263 4113
rect 1316 4063 1323 4253
rect 1336 4227 1343 4303
rect 1376 4296 1403 4303
rect 1356 4187 1363 4233
rect 1316 4056 1343 4063
rect 1293 4040 1307 4053
rect 1296 4036 1303 4040
rect 1336 4036 1343 4056
rect 976 3836 1003 3843
rect 996 3816 1003 3836
rect 727 3756 743 3767
rect 727 3753 740 3756
rect 576 3567 583 3613
rect 553 3520 567 3533
rect 556 3516 563 3520
rect 596 3516 603 3593
rect 636 3567 643 3593
rect 656 3487 663 3514
rect 676 3447 683 3553
rect 776 3516 783 3553
rect 456 3047 463 3294
rect 476 3243 483 3263
rect 476 3236 503 3243
rect 476 3087 483 3213
rect 496 3147 503 3236
rect 536 3227 543 3263
rect 476 2996 483 3073
rect 496 3023 503 3133
rect 496 3016 523 3023
rect 516 2996 523 3016
rect 356 2960 363 2963
rect 236 2867 243 2913
rect 236 2783 243 2853
rect 156 2776 183 2783
rect 216 2776 243 2783
rect 16 2187 23 2333
rect 36 2307 43 2773
rect 76 2707 83 2743
rect 56 2696 73 2703
rect 56 2487 63 2696
rect 156 2483 163 2776
rect 256 2743 263 2933
rect 316 2887 323 2953
rect 353 2947 367 2960
rect 356 2776 363 2873
rect 396 2827 403 2963
rect 496 2927 503 2963
rect 507 2916 523 2923
rect 236 2736 263 2743
rect 236 2647 243 2736
rect 336 2667 343 2743
rect 136 2476 163 2483
rect 196 2476 203 2513
rect 236 2476 243 2633
rect 333 2507 347 2513
rect 376 2508 383 2733
rect 116 2256 123 2293
rect 136 2287 143 2476
rect 333 2480 347 2493
rect 336 2476 343 2480
rect 396 2483 403 2792
rect 416 2787 423 2853
rect 447 2803 460 2807
rect 447 2793 463 2803
rect 456 2776 463 2793
rect 496 2787 503 2813
rect 516 2707 523 2916
rect 536 2787 543 2893
rect 576 2847 583 3333
rect 596 3266 603 3293
rect 676 3227 683 3252
rect 596 2803 603 2873
rect 636 2807 643 2952
rect 673 2907 687 2913
rect 696 2887 703 2993
rect 716 2907 723 3483
rect 736 3227 743 3433
rect 756 3387 763 3483
rect 816 3482 823 3533
rect 856 3516 863 3553
rect 876 3547 883 3772
rect 976 3687 983 3783
rect 1056 3567 1063 3873
rect 1096 3827 1103 3993
rect 1176 3947 1183 4003
rect 1216 3996 1243 4003
rect 1173 3820 1187 3833
rect 1176 3816 1183 3820
rect 996 3516 1003 3553
rect 1076 3523 1083 3813
rect 1107 3783 1120 3787
rect 1107 3776 1123 3783
rect 1107 3773 1120 3776
rect 1156 3727 1163 3783
rect 1216 3687 1223 3996
rect 1236 3827 1243 3973
rect 1316 3907 1323 4003
rect 1273 3820 1287 3833
rect 1276 3816 1283 3820
rect 1356 3786 1363 3913
rect 1376 3827 1383 4273
rect 1396 4227 1403 4296
rect 1416 4163 1423 4353
rect 1436 4343 1443 4413
rect 1496 4407 1503 4453
rect 1453 4367 1467 4373
rect 1436 4336 1463 4343
rect 1516 4347 1523 4773
rect 1536 4307 1543 4693
rect 1616 4563 1623 4933
rect 1656 4907 1663 5013
rect 1676 4868 1683 4973
rect 1696 4967 1703 5036
rect 1733 5027 1747 5040
rect 1796 4987 1803 5074
rect 1936 5047 1943 5253
rect 1956 5087 1963 5173
rect 2076 5147 2083 5336
rect 2116 5307 2123 5343
rect 2136 5223 2143 5313
rect 2156 5307 2163 5343
rect 2236 5327 2243 5343
rect 2156 5247 2163 5293
rect 2136 5216 2163 5223
rect 2087 5136 2103 5143
rect 2067 5093 2073 5107
rect 1993 5080 2007 5093
rect 1996 5076 2003 5080
rect 2096 5083 2103 5136
rect 2076 5076 2103 5083
rect 2113 5080 2127 5093
rect 2156 5087 2163 5216
rect 2116 5076 2123 5080
rect 1816 4963 1823 5033
rect 1796 4956 1823 4963
rect 1636 4787 1643 4823
rect 1716 4823 1723 4913
rect 1796 4856 1803 4956
rect 1836 4868 1843 4953
rect 1856 4887 1863 5043
rect 2076 5046 2083 5076
rect 1936 4856 1943 5012
rect 1976 4947 1983 5043
rect 1707 4816 1723 4823
rect 1736 4707 1743 4853
rect 1656 4587 1663 4633
rect 1616 4556 1643 4563
rect 1556 4447 1563 4493
rect 1576 4447 1583 4523
rect 1636 4467 1643 4556
rect 1656 4527 1663 4573
rect 1676 4443 1683 4613
rect 1696 4556 1703 4653
rect 1756 4587 1763 4753
rect 1816 4747 1823 4823
rect 1796 4587 1803 4653
rect 1816 4607 1823 4733
rect 1836 4568 1843 4613
rect 1876 4587 1883 4854
rect 1896 4607 1903 4653
rect 1916 4587 1923 4823
rect 1936 4647 1943 4773
rect 1956 4623 1963 4812
rect 1996 4787 2003 5013
rect 2016 4707 2023 4993
rect 2116 4823 2123 4993
rect 2176 4923 2183 5273
rect 2236 5187 2243 5313
rect 2216 5076 2223 5133
rect 2336 5107 2343 5373
rect 2416 5340 2423 5343
rect 2413 5327 2427 5340
rect 2456 5307 2463 5333
rect 2476 5267 2483 5373
rect 2516 5227 2523 5343
rect 2556 5287 2563 5343
rect 2356 5088 2363 5193
rect 2396 5076 2403 5133
rect 2496 5127 2503 5193
rect 2556 5167 2563 5213
rect 2176 4916 2203 4923
rect 2096 4816 2123 4823
rect 2116 4687 2123 4773
rect 2136 4627 2143 4913
rect 1936 4616 1963 4623
rect 1756 4556 1783 4563
rect 1716 4527 1730 4532
rect 1776 4507 1783 4556
rect 1873 4560 1887 4573
rect 1876 4556 1883 4560
rect 1796 4527 1803 4552
rect 1916 4527 1923 4573
rect 1936 4567 1943 4616
rect 1976 4556 1983 4613
rect 2013 4560 2027 4573
rect 2016 4556 2023 4560
rect 1796 4516 1813 4527
rect 1800 4513 1813 4516
rect 1707 4503 1720 4507
rect 1707 4493 1723 4503
rect 1716 4447 1723 4493
rect 1676 4436 1703 4443
rect 1576 4387 1583 4433
rect 1653 4423 1667 4433
rect 1653 4420 1683 4423
rect 1656 4416 1683 4420
rect 1596 4336 1603 4373
rect 1436 4207 1443 4253
rect 1476 4247 1483 4303
rect 1396 4156 1423 4163
rect 1396 3887 1403 4156
rect 1436 4127 1443 4172
rect 1473 4103 1487 4113
rect 1516 4103 1523 4293
rect 1576 4247 1583 4303
rect 1536 4107 1543 4213
rect 1456 4100 1487 4103
rect 1453 4096 1483 4100
rect 1496 4096 1523 4103
rect 1453 4087 1467 4096
rect 1413 4040 1427 4053
rect 1473 4040 1487 4053
rect 1496 4048 1503 4096
rect 1416 4036 1423 4040
rect 1476 4036 1483 4040
rect 1456 4000 1463 4003
rect 1453 3987 1467 4000
rect 1467 3976 1483 3983
rect 1416 3816 1423 3973
rect 1256 3747 1263 3783
rect 1336 3776 1353 3783
rect 1296 3627 1303 3772
rect 1336 3528 1343 3776
rect 1436 3747 1443 3772
rect 1076 3516 1103 3523
rect 1256 3516 1283 3523
rect 816 3475 873 3482
rect 836 3263 843 3333
rect 916 3323 923 3483
rect 1016 3480 1023 3483
rect 1013 3467 1027 3480
rect 1056 3347 1063 3483
rect 1056 3336 1073 3347
rect 1060 3333 1073 3336
rect 916 3316 943 3323
rect 936 3308 943 3316
rect 1096 3308 1103 3516
rect 1116 3447 1123 3493
rect 1276 3487 1283 3516
rect 1376 3516 1383 3553
rect 1476 3548 1483 3976
rect 1496 3827 1503 4034
rect 1516 4007 1523 4053
rect 1556 4036 1563 4173
rect 1596 4127 1603 4253
rect 1616 4147 1623 4303
rect 1596 4036 1603 4073
rect 1636 4006 1643 4273
rect 1656 4047 1663 4293
rect 1676 4087 1683 4416
rect 1696 4347 1703 4436
rect 1736 4336 1743 4493
rect 1833 4487 1847 4493
rect 1776 4347 1783 4453
rect 1716 4247 1723 4303
rect 1756 4127 1763 4303
rect 1796 4267 1803 4473
rect 1820 4443 1833 4447
rect 1816 4433 1833 4443
rect 1816 4367 1823 4433
rect 1856 4336 1863 4373
rect 1896 4336 1903 4513
rect 2016 4447 2023 4493
rect 2036 4467 2043 4513
rect 2056 4447 2063 4573
rect 1916 4387 1923 4413
rect 1916 4347 1923 4373
rect 1816 4187 1823 4293
rect 1876 4283 1883 4303
rect 1876 4276 1903 4283
rect 1673 4040 1687 4052
rect 1676 4036 1683 4040
rect 1836 4036 1843 4193
rect 1856 4087 1863 4153
rect 1876 4048 1883 4193
rect 1616 3927 1623 3993
rect 1696 3907 1703 4003
rect 1516 3816 1523 3853
rect 1696 3848 1703 3893
rect 1556 3840 1603 3843
rect 1556 3836 1607 3840
rect 1556 3816 1563 3836
rect 1593 3827 1607 3836
rect 1716 3843 1723 3873
rect 1736 3867 1743 3992
rect 1776 3927 1783 4033
rect 1896 4007 1903 4276
rect 1916 4047 1923 4293
rect 1936 4247 1943 4393
rect 1976 4336 1983 4373
rect 1996 4367 2003 4393
rect 2016 4348 2023 4433
rect 2096 4383 2103 4433
rect 2116 4407 2123 4523
rect 2156 4467 2163 4873
rect 2176 4867 2183 4893
rect 2196 4887 2203 4916
rect 2216 4856 2223 5013
rect 2276 4927 2283 5043
rect 2236 4787 2243 4823
rect 2176 4443 2183 4633
rect 2216 4556 2223 4593
rect 2256 4568 2263 4793
rect 2296 4607 2303 5033
rect 2316 5007 2323 5074
rect 2376 5007 2383 5043
rect 2396 4967 2403 5013
rect 2416 4967 2423 5043
rect 2456 5027 2463 5093
rect 2516 5076 2523 5153
rect 2553 5080 2567 5093
rect 2576 5087 2583 5153
rect 2556 5076 2563 5080
rect 2456 5016 2473 5027
rect 2460 5013 2473 5016
rect 2496 5007 2503 5043
rect 2536 5040 2543 5043
rect 2533 5027 2547 5040
rect 2573 5023 2587 5033
rect 2556 5020 2587 5023
rect 2556 5016 2583 5020
rect 2356 4856 2363 4913
rect 2416 4907 2423 4932
rect 2433 4883 2447 4893
rect 2396 4880 2447 4883
rect 2396 4876 2443 4880
rect 2396 4856 2403 4876
rect 2456 4867 2463 4993
rect 2496 4856 2503 4913
rect 2556 4907 2563 5016
rect 2376 4727 2383 4823
rect 2413 4807 2427 4813
rect 2396 4747 2403 4793
rect 2336 4568 2343 4633
rect 2396 4556 2403 4673
rect 2416 4647 2423 4753
rect 2436 4687 2443 4853
rect 2456 4816 2483 4823
rect 2456 4727 2463 4816
rect 2176 4436 2203 4443
rect 2096 4376 2123 4383
rect 2027 4336 2043 4343
rect 1996 4247 2003 4303
rect 1936 4067 1943 4113
rect 1933 4040 1947 4053
rect 1936 4036 1943 4040
rect 1976 4036 1983 4193
rect 2016 4043 2023 4133
rect 2036 4063 2043 4336
rect 2116 4336 2123 4376
rect 2096 4147 2103 4303
rect 2176 4167 2183 4413
rect 2196 4267 2203 4436
rect 2236 4367 2243 4523
rect 2276 4447 2283 4513
rect 2296 4487 2303 4553
rect 2416 4526 2423 4633
rect 2256 4336 2263 4393
rect 2296 4347 2303 4473
rect 2316 4347 2323 4493
rect 2336 4447 2343 4473
rect 2336 4347 2343 4433
rect 2396 4336 2403 4413
rect 2236 4247 2243 4303
rect 2036 4056 2063 4063
rect 2016 4036 2043 4043
rect 1716 3836 1743 3843
rect 1736 3816 1743 3836
rect 1753 3827 1767 3833
rect 1496 3647 1503 3773
rect 1536 3727 1543 3783
rect 1136 3476 1163 3483
rect 1136 3407 1143 3476
rect 1116 3307 1123 3333
rect 816 3256 843 3263
rect 836 2996 863 3003
rect 916 2996 923 3263
rect 996 3003 1003 3293
rect 1096 3266 1103 3294
rect 1127 3296 1143 3303
rect 1176 3296 1183 3333
rect 1276 3327 1283 3473
rect 1296 3347 1303 3513
rect 1356 3480 1363 3483
rect 1353 3467 1367 3480
rect 1416 3447 1423 3533
rect 1536 3527 1543 3713
rect 1456 3447 1463 3483
rect 1533 3467 1547 3473
rect 1396 3436 1413 3443
rect 1056 3247 1063 3263
rect 1156 3260 1163 3263
rect 1056 3236 1073 3247
rect 1060 3233 1073 3236
rect 976 2996 1003 3003
rect 856 2927 863 2996
rect 976 2966 983 2996
rect 1096 3003 1103 3252
rect 1116 3008 1123 3253
rect 1153 3247 1167 3260
rect 1236 3087 1243 3313
rect 1256 3067 1263 3213
rect 1076 2996 1103 3003
rect 576 2796 603 2803
rect 576 2776 583 2796
rect 616 2773 633 2787
rect 696 2776 703 2833
rect 876 2827 883 2952
rect 616 2768 626 2773
rect 656 2746 663 2773
rect 796 2767 803 2793
rect 816 2787 823 2813
rect 833 2780 847 2793
rect 836 2776 843 2780
rect 956 2787 963 2813
rect 996 2776 1003 2913
rect 1016 2827 1023 2963
rect 1136 2867 1143 3033
rect 1336 3027 1343 3293
rect 1356 3147 1363 3333
rect 1396 3296 1403 3436
rect 1473 3300 1487 3313
rect 1496 3307 1503 3451
rect 1476 3296 1483 3300
rect 1416 3243 1423 3263
rect 1416 3240 1443 3243
rect 1416 3236 1447 3240
rect 1433 3227 1447 3236
rect 1276 2963 1283 3013
rect 1336 2996 1343 3013
rect 1376 3008 1383 3033
rect 1256 2956 1283 2963
rect 1216 2807 1223 2913
rect 1356 2883 1363 2963
rect 1336 2876 1363 2883
rect 1253 2780 1267 2793
rect 1256 2776 1263 2780
rect 1296 2776 1303 2813
rect 556 2667 563 2732
rect 636 2507 643 2733
rect 756 2707 763 2743
rect 896 2740 903 2743
rect 893 2727 907 2740
rect 893 2707 907 2713
rect 936 2547 943 2773
rect 1196 2747 1203 2774
rect 1013 2707 1027 2711
rect 1136 2707 1143 2743
rect 1013 2700 1033 2707
rect 1016 2696 1033 2700
rect 1020 2693 1033 2696
rect 996 2647 1003 2693
rect 1336 2667 1343 2876
rect 1356 2783 1363 2853
rect 1416 2847 1423 3193
rect 1456 3087 1463 3263
rect 1496 3007 1503 3253
rect 1516 3008 1523 3313
rect 1536 3303 1543 3393
rect 1556 3327 1563 3633
rect 1596 3567 1603 3733
rect 1616 3687 1623 3793
rect 1636 3786 1643 3813
rect 1596 3516 1603 3553
rect 1636 3516 1643 3633
rect 1616 3467 1623 3483
rect 1676 3467 1683 3533
rect 1696 3523 1703 3713
rect 1716 3687 1723 3772
rect 1776 3543 1783 3913
rect 1796 3827 1803 3853
rect 1816 3847 1823 3992
rect 1856 3947 1863 4003
rect 1836 3816 1843 3893
rect 1856 3887 1863 3933
rect 1896 3823 1903 3953
rect 1996 3947 2003 4003
rect 2036 3907 2043 4036
rect 2056 3903 2063 4056
rect 2073 4040 2087 4053
rect 2076 4036 2083 4040
rect 2136 4036 2143 4133
rect 2096 3967 2103 4003
rect 2156 3983 2163 4034
rect 2136 3976 2163 3983
rect 2056 3900 2083 3903
rect 2056 3896 2087 3900
rect 2073 3887 2087 3896
rect 1876 3816 1903 3823
rect 1916 3816 1923 3853
rect 1936 3847 1943 3873
rect 1816 3747 1823 3783
rect 1756 3536 1783 3543
rect 1696 3516 1723 3523
rect 1756 3516 1763 3536
rect 1796 3527 1803 3713
rect 1856 3623 1863 3773
rect 1876 3747 1883 3816
rect 1976 3747 1983 3783
rect 2016 3767 2023 3783
rect 1876 3667 1883 3733
rect 1856 3616 1883 3623
rect 1616 3383 1623 3453
rect 1616 3376 1643 3383
rect 1536 3296 1563 3303
rect 1536 3227 1543 3253
rect 1576 3247 1583 3263
rect 1567 3236 1583 3247
rect 1567 3233 1580 3236
rect 1556 3127 1563 3193
rect 1616 3167 1623 3353
rect 1636 3307 1643 3376
rect 1716 3308 1723 3433
rect 1776 3407 1783 3472
rect 1876 3467 1883 3616
rect 1896 3507 1903 3613
rect 1916 3527 1923 3733
rect 1933 3520 1947 3533
rect 1936 3516 1943 3520
rect 2016 3523 2023 3753
rect 2116 3727 2123 3893
rect 2007 3516 2023 3523
rect 1736 3363 1743 3393
rect 1767 3376 1793 3383
rect 1856 3363 1863 3393
rect 1876 3387 1883 3432
rect 1916 3387 1923 3473
rect 1736 3356 1763 3363
rect 1856 3360 1883 3363
rect 1856 3356 1887 3360
rect 1756 3287 1763 3356
rect 1873 3347 1887 3356
rect 1833 3300 1847 3313
rect 1836 3296 1843 3300
rect 1496 2807 1503 2953
rect 1516 2927 1523 2994
rect 1536 2966 1543 3073
rect 1556 2996 1563 3033
rect 1576 3027 1583 3133
rect 1676 3003 1683 3233
rect 1696 3227 1703 3263
rect 1616 2996 1643 3003
rect 1536 2907 1543 2952
rect 1356 2776 1383 2783
rect 1516 2746 1523 2833
rect 1636 2783 1643 2996
rect 1656 2996 1683 3003
rect 1693 3000 1707 3013
rect 1736 3007 1743 3253
rect 1856 3227 1863 3253
rect 1696 2996 1703 3000
rect 1656 2966 1663 2996
rect 1756 2947 1763 3093
rect 1816 2996 1823 3173
rect 1856 2996 1863 3113
rect 1876 3087 1883 3333
rect 1956 3296 1963 3333
rect 1936 3127 1943 3263
rect 1996 3187 2003 3413
rect 2016 3147 2023 3473
rect 2036 3327 2043 3633
rect 2116 3587 2123 3713
rect 2136 3647 2143 3976
rect 2176 3967 2183 4153
rect 2236 4048 2243 4153
rect 2276 3947 2283 4133
rect 2296 4047 2303 4293
rect 2316 4087 2323 4312
rect 2316 4036 2323 4073
rect 2356 4047 2363 4292
rect 2336 3947 2343 4003
rect 2176 3907 2183 3932
rect 2196 3847 2203 3933
rect 2336 3907 2343 3933
rect 2196 3816 2203 3833
rect 2256 3780 2263 3783
rect 2253 3767 2267 3780
rect 2316 3763 2323 3783
rect 2316 3756 2343 3763
rect 2056 3467 2063 3553
rect 2076 3527 2083 3573
rect 2113 3520 2127 3533
rect 2116 3516 2123 3520
rect 2076 3427 2083 3473
rect 2096 3407 2103 3483
rect 2136 3480 2143 3483
rect 2133 3467 2147 3480
rect 2076 3296 2083 3373
rect 2096 3327 2103 3393
rect 2136 3267 2143 3373
rect 2156 3308 2163 3353
rect 2176 3343 2183 3473
rect 2196 3367 2203 3673
rect 2296 3516 2303 3553
rect 2336 3547 2343 3756
rect 2356 3687 2363 3833
rect 2376 3828 2383 4073
rect 2396 4006 2403 4193
rect 2436 4067 2443 4593
rect 2476 4568 2483 4773
rect 2516 4767 2523 4812
rect 2516 4556 2523 4732
rect 2576 4727 2583 4993
rect 2596 4867 2603 5523
rect 2956 5487 2963 5523
rect 2636 5388 2643 5433
rect 2936 5427 2943 5453
rect 2756 5387 2763 5413
rect 2796 5376 2803 5413
rect 2953 5380 2967 5393
rect 2956 5376 2963 5380
rect 2700 5343 2713 5347
rect 2613 5327 2627 5333
rect 2616 5087 2623 5173
rect 2656 5147 2663 5343
rect 2696 5336 2713 5343
rect 2700 5333 2713 5336
rect 2736 5327 2743 5373
rect 2776 5340 2783 5343
rect 2773 5327 2787 5340
rect 2876 5336 2893 5343
rect 2756 5316 2773 5323
rect 2727 5273 2733 5287
rect 2676 5127 2683 5213
rect 2636 5076 2643 5113
rect 2756 5107 2763 5316
rect 2816 5283 2823 5311
rect 2787 5276 2823 5283
rect 2876 5267 2883 5336
rect 2787 5196 2813 5203
rect 2816 5127 2823 5153
rect 2856 5127 2863 5173
rect 2876 5127 2883 5232
rect 2896 5187 2903 5293
rect 2916 5287 2923 5313
rect 2673 5088 2687 5092
rect 2760 5086 2780 5087
rect 2767 5083 2780 5086
rect 2767 5076 2783 5083
rect 2767 5073 2780 5076
rect 2916 5076 2923 5213
rect 2976 5187 2983 5343
rect 2956 5076 2963 5113
rect 2613 5027 2627 5032
rect 2676 4887 2683 4993
rect 2696 4947 2703 5043
rect 2713 5027 2727 5033
rect 2736 4967 2743 5053
rect 2756 4947 2763 5033
rect 2796 4967 2803 5043
rect 2696 4907 2703 4933
rect 2716 4883 2723 4933
rect 2696 4880 2723 4883
rect 2693 4876 2723 4880
rect 2693 4867 2707 4876
rect 2736 4856 2743 4893
rect 2576 4526 2583 4593
rect 2496 4467 2503 4523
rect 2536 4487 2543 4523
rect 2576 4427 2583 4453
rect 2533 4340 2547 4353
rect 2536 4336 2543 4340
rect 2456 4163 2463 4333
rect 2516 4283 2523 4303
rect 2496 4276 2523 4283
rect 2496 4227 2503 4276
rect 2596 4247 2603 4813
rect 2616 4767 2623 4823
rect 2676 4787 2683 4833
rect 2716 4747 2723 4812
rect 2636 4660 2683 4663
rect 2633 4656 2683 4660
rect 2633 4647 2647 4656
rect 2646 4640 2647 4647
rect 2616 4556 2623 4593
rect 2656 4587 2663 4633
rect 2676 4587 2683 4656
rect 2696 4583 2703 4733
rect 2736 4607 2743 4793
rect 2756 4787 2763 4823
rect 2796 4707 2803 4813
rect 2816 4627 2823 5013
rect 2836 4887 2843 5043
rect 2876 4856 2883 4893
rect 2896 4887 2903 4953
rect 2936 4947 2943 5043
rect 2976 5023 2983 5032
rect 3016 5027 3023 5473
rect 3036 5387 3043 5523
rect 3636 5516 3644 5523
rect 3476 5476 3523 5483
rect 3067 5460 3103 5463
rect 3067 5456 3107 5460
rect 3093 5447 3107 5456
rect 3133 5447 3147 5453
rect 3076 5388 3083 5433
rect 3047 5346 3060 5347
rect 3047 5333 3053 5346
rect 3093 5327 3107 5332
rect 3116 5307 3123 5433
rect 3196 5407 3203 5433
rect 3133 5387 3147 5393
rect 3216 5376 3223 5433
rect 3056 5267 3063 5293
rect 3076 5227 3083 5293
rect 3156 5247 3163 5343
rect 3233 5327 3247 5333
rect 3256 5323 3263 5453
rect 3356 5376 3363 5413
rect 3476 5407 3483 5476
rect 3496 5376 3503 5453
rect 3516 5388 3523 5476
rect 3636 5407 3643 5516
rect 3673 5447 3687 5453
rect 3713 5447 3727 5453
rect 3396 5347 3403 5374
rect 3247 5316 3263 5323
rect 3296 5307 3303 5332
rect 3236 5247 3243 5292
rect 3167 5236 3183 5243
rect 3096 5187 3103 5233
rect 3076 5076 3083 5113
rect 3116 5088 3123 5173
rect 2956 5016 2983 5023
rect 2916 4856 2923 4893
rect 2936 4867 2943 4912
rect 2856 4787 2863 4812
rect 2896 4747 2903 4823
rect 2916 4767 2923 4793
rect 2936 4687 2943 4813
rect 2836 4647 2843 4673
rect 2696 4576 2723 4583
rect 2676 4556 2703 4563
rect 2616 4347 2623 4413
rect 2656 4363 2663 4493
rect 2696 4487 2703 4556
rect 2636 4356 2663 4363
rect 2636 4336 2643 4356
rect 2676 4336 2683 4373
rect 2696 4367 2703 4473
rect 2716 4447 2723 4576
rect 2736 4306 2743 4572
rect 2813 4560 2827 4573
rect 2816 4556 2823 4560
rect 2856 4547 2863 4613
rect 2792 4528 2806 4532
rect 2756 4427 2763 4513
rect 2787 4503 2800 4507
rect 2787 4493 2803 4503
rect 2796 4407 2803 4493
rect 2836 4467 2843 4513
rect 2876 4523 2883 4673
rect 2896 4587 2903 4633
rect 2956 4627 2963 5016
rect 3096 4927 3103 5043
rect 2976 4867 2983 4893
rect 2976 4687 2983 4813
rect 3056 4820 3063 4823
rect 3053 4807 3067 4820
rect 2947 4596 2973 4603
rect 2933 4560 2947 4572
rect 2936 4556 2943 4560
rect 2876 4516 2923 4523
rect 2856 4427 2863 4512
rect 2896 4447 2903 4493
rect 2956 4447 2963 4523
rect 2996 4447 3003 4513
rect 2796 4336 2803 4372
rect 2473 4163 2487 4173
rect 2456 4160 2487 4163
rect 2456 4156 2483 4160
rect 2456 4036 2463 4133
rect 2476 4047 2483 4156
rect 2413 3987 2427 3993
rect 2436 3967 2443 4003
rect 2476 3883 2483 3993
rect 2496 3927 2503 4213
rect 2556 4067 2563 4113
rect 2656 4103 2663 4233
rect 2676 4147 2683 4273
rect 2716 4147 2723 4213
rect 2796 4187 2803 4273
rect 2656 4096 2683 4103
rect 2553 4040 2567 4053
rect 2556 4036 2563 4040
rect 2676 4036 2683 4096
rect 2780 4083 2793 4087
rect 2776 4073 2793 4083
rect 2776 4036 2783 4073
rect 2516 3967 2523 3993
rect 2476 3876 2503 3883
rect 2476 3828 2483 3853
rect 2356 3523 2363 3633
rect 2416 3528 2423 3593
rect 2476 3583 2483 3814
rect 2496 3767 2503 3876
rect 2516 3647 2523 3932
rect 2536 3927 2543 4003
rect 2576 3867 2583 3973
rect 2596 3967 2603 4034
rect 2716 4007 2723 4034
rect 2596 3816 2603 3873
rect 2576 3780 2583 3783
rect 2616 3780 2623 3783
rect 2573 3767 2587 3780
rect 2613 3767 2627 3780
rect 2656 3647 2663 3953
rect 2736 3687 2743 3783
rect 2776 3767 2783 3813
rect 2796 3747 2803 3993
rect 2816 3967 2823 4303
rect 2836 4047 2843 4213
rect 2856 4107 2863 4293
rect 2876 4167 2883 4333
rect 2896 4287 2903 4373
rect 2916 4347 2923 4433
rect 2953 4340 2967 4353
rect 2956 4336 2963 4340
rect 2980 4303 2993 4307
rect 2936 4267 2943 4303
rect 2976 4296 2993 4303
rect 2980 4293 2993 4296
rect 3016 4167 3023 4673
rect 3036 4567 3043 4793
rect 3096 4767 3103 4854
rect 3116 4826 3123 4873
rect 3136 4863 3143 4993
rect 3156 4887 3163 5153
rect 3176 5087 3183 5236
rect 3276 5243 3283 5273
rect 3276 5236 3303 5243
rect 3196 5076 3203 5193
rect 3236 5076 3243 5133
rect 3256 5107 3263 5193
rect 3296 5187 3303 5236
rect 3316 5227 3323 5313
rect 3336 5207 3343 5343
rect 3376 5267 3383 5333
rect 3436 5267 3443 5332
rect 3476 5307 3483 5343
rect 3536 5343 3543 5393
rect 3636 5376 3643 5393
rect 3696 5346 3703 5433
rect 3756 5376 3763 5413
rect 3776 5407 3783 5473
rect 3536 5336 3563 5343
rect 3456 5276 3493 5283
rect 3456 5227 3463 5276
rect 3353 5167 3367 5173
rect 3296 5083 3303 5133
rect 3276 5076 3303 5083
rect 3176 4883 3183 5033
rect 3216 4987 3223 5043
rect 3256 5040 3263 5043
rect 3253 5027 3267 5040
rect 3176 4876 3203 4883
rect 3136 4856 3163 4863
rect 3196 4856 3203 4876
rect 3256 4826 3263 4992
rect 3296 4947 3303 5033
rect 3316 5027 3323 5073
rect 3336 5047 3343 5093
rect 3356 5087 3363 5113
rect 3373 5080 3387 5093
rect 3376 5076 3383 5080
rect 3356 5007 3363 5033
rect 3396 5007 3403 5043
rect 3436 5040 3443 5043
rect 3433 5027 3447 5040
rect 3456 4967 3463 5033
rect 3476 5027 3483 5253
rect 3516 5207 3523 5333
rect 3496 5196 3513 5203
rect 3496 5087 3503 5196
rect 3536 5167 3543 5313
rect 3556 5307 3563 5336
rect 3576 5283 3583 5343
rect 3556 5280 3583 5283
rect 3553 5276 3583 5280
rect 3553 5267 3567 5276
rect 3616 5247 3623 5343
rect 3656 5340 3663 5343
rect 3653 5327 3667 5340
rect 3573 5227 3587 5233
rect 3573 5220 3593 5227
rect 3576 5216 3593 5220
rect 3580 5213 3593 5216
rect 3636 5207 3643 5293
rect 3716 5287 3723 5313
rect 3776 5307 3783 5343
rect 3547 5113 3553 5127
rect 3533 5080 3547 5092
rect 3576 5088 3583 5133
rect 3536 5076 3543 5080
rect 3636 5087 3643 5113
rect 3696 5088 3703 5253
rect 3716 5107 3723 5173
rect 3647 5083 3660 5087
rect 3647 5076 3663 5083
rect 3647 5073 3660 5076
rect 3556 5023 3563 5043
rect 3556 5020 3583 5023
rect 3556 5016 3587 5020
rect 3573 5007 3587 5016
rect 3333 4883 3347 4893
rect 3316 4880 3347 4883
rect 3316 4876 3343 4880
rect 3316 4856 3323 4876
rect 3176 4820 3183 4823
rect 3173 4807 3187 4820
rect 3296 4787 3303 4823
rect 3376 4787 3383 4853
rect 3396 4807 3403 4913
rect 3536 4823 3543 4993
rect 3596 4967 3603 5033
rect 3587 4956 3603 4967
rect 3587 4953 3600 4956
rect 3596 4856 3603 4933
rect 3056 4647 3063 4673
rect 3036 4516 3063 4523
rect 3036 4367 3043 4516
rect 3056 4336 3063 4373
rect 3096 4336 3103 4513
rect 3116 4427 3123 4613
rect 3147 4563 3160 4567
rect 3147 4556 3163 4563
rect 3196 4556 3203 4613
rect 3147 4553 3160 4556
rect 3296 4556 3303 4613
rect 3336 4568 3343 4773
rect 3256 4526 3263 4553
rect 3376 4527 3383 4733
rect 3416 4687 3423 4812
rect 3476 4767 3483 4823
rect 3536 4816 3563 4823
rect 3396 4567 3403 4633
rect 3436 4556 3443 4593
rect 3236 4407 3243 4493
rect 3293 4487 3307 4493
rect 3256 4387 3263 4473
rect 3156 4347 3163 4373
rect 3253 4347 3267 4352
rect 2887 4073 2893 4087
rect 2936 4047 2943 4153
rect 2816 3816 2823 3873
rect 2836 3847 2843 3993
rect 2876 3983 2883 4003
rect 2933 3983 2947 3993
rect 2876 3976 2903 3983
rect 2856 3747 2863 3783
rect 2876 3727 2883 3953
rect 2896 3907 2903 3976
rect 2916 3980 2947 3983
rect 2916 3976 2943 3980
rect 2896 3687 2903 3853
rect 2467 3576 2483 3583
rect 2336 3516 2363 3523
rect 2216 3387 2223 3473
rect 2236 3447 2243 3483
rect 2313 3467 2327 3472
rect 2336 3447 2343 3516
rect 2436 3527 2443 3553
rect 2433 3467 2447 3473
rect 2176 3336 2203 3343
rect 2196 3296 2203 3336
rect 1976 3067 1983 3113
rect 1636 2776 1653 2783
rect 1713 2780 1727 2793
rect 1716 2776 1723 2780
rect 1656 2743 1663 2774
rect 1776 2767 1783 2893
rect 1796 2867 1803 2952
rect 1796 2787 1803 2832
rect 1836 2776 1843 2963
rect 1896 2927 1903 2963
rect 1956 2927 1963 3033
rect 1996 3023 2003 3113
rect 2056 3087 2063 3263
rect 2096 3260 2103 3263
rect 2093 3247 2107 3260
rect 2216 3256 2243 3263
rect 1996 3016 2023 3023
rect 1976 2887 1983 3013
rect 2016 2996 2023 3016
rect 2076 2996 2083 3133
rect 2096 3007 2103 3073
rect 1996 2783 2003 2953
rect 1976 2776 2003 2783
rect 2016 2746 2023 2793
rect 2036 2787 2043 2833
rect 2096 2807 2103 2953
rect 2116 2947 2123 3053
rect 2136 2827 2143 3113
rect 2176 3008 2183 3252
rect 2236 3187 2243 3256
rect 2216 3127 2223 3153
rect 2256 3147 2263 3263
rect 2316 3243 2323 3263
rect 2316 3236 2343 3243
rect 2216 2996 2223 3113
rect 2156 2803 2163 2953
rect 2256 2847 2263 3073
rect 2336 3067 2343 3236
rect 2356 3087 2363 3353
rect 2376 3107 2383 3433
rect 2456 3327 2463 3573
rect 2536 3516 2543 3573
rect 2756 3516 2763 3573
rect 2476 3266 2483 3333
rect 2356 2867 2363 2963
rect 2376 2903 2383 2952
rect 2396 2927 2403 3053
rect 2436 2996 2443 3113
rect 2476 2996 2483 3153
rect 2496 3127 2503 3393
rect 2516 3347 2523 3483
rect 2576 3427 2583 3514
rect 2516 3247 2523 3312
rect 2536 3244 2543 3263
rect 2527 3237 2543 3244
rect 2536 3167 2543 3237
rect 2596 3003 2603 3333
rect 2616 3227 2623 3433
rect 2636 3367 2643 3483
rect 2676 3480 2683 3483
rect 2673 3467 2687 3480
rect 2716 3447 2723 3514
rect 2776 3427 2783 3483
rect 2836 3383 2843 3633
rect 2916 3587 2923 3976
rect 2936 3867 2943 3953
rect 2956 3947 2963 4093
rect 2976 4047 2983 4153
rect 3016 4048 3023 4132
rect 3036 4067 3043 4113
rect 3056 4036 3063 4093
rect 3076 4047 3083 4303
rect 3116 4300 3123 4303
rect 3113 4287 3127 4300
rect 3096 4167 3103 4253
rect 3156 4243 3163 4312
rect 3136 4236 3163 4243
rect 3176 4243 3183 4293
rect 3196 4267 3203 4303
rect 3236 4300 3243 4303
rect 3233 4287 3247 4300
rect 3253 4287 3267 4293
rect 3276 4287 3283 4393
rect 3296 4347 3303 4413
rect 3376 4347 3383 4393
rect 3396 4303 3403 4473
rect 3440 4363 3453 4367
rect 3436 4353 3453 4363
rect 3436 4348 3447 4353
rect 3476 4348 3483 4554
rect 3496 4427 3503 4713
rect 3516 4556 3523 4633
rect 3576 4523 3583 4633
rect 3556 4516 3583 4523
rect 3556 4387 3563 4493
rect 3513 4348 3527 4353
rect 3176 4236 3213 4243
rect 3108 4087 3115 4133
rect 3136 4087 3143 4236
rect 3176 4107 3183 4193
rect 3216 4147 3223 4193
rect 3096 4003 3103 4053
rect 3133 4040 3147 4052
rect 3136 4036 3143 4040
rect 3176 4036 3183 4072
rect 3193 4047 3207 4053
rect 2976 3923 2983 3993
rect 2996 3947 3003 4003
rect 2956 3916 2983 3923
rect 2956 3843 2963 3916
rect 2936 3840 2963 3843
rect 2933 3836 2963 3840
rect 2933 3827 2947 3836
rect 2976 3816 2983 3893
rect 3036 3887 3043 4003
rect 3076 3996 3103 4003
rect 2996 3847 3003 3873
rect 2956 3780 2963 3783
rect 2936 3627 2943 3773
rect 2953 3767 2967 3780
rect 2996 3727 3003 3783
rect 3036 3727 3043 3773
rect 2876 3528 2883 3573
rect 2936 3523 2943 3613
rect 2916 3516 2943 3523
rect 2896 3480 2903 3483
rect 2893 3467 2907 3480
rect 2896 3427 2903 3453
rect 2956 3447 2963 3493
rect 2976 3486 2983 3613
rect 2996 3587 3003 3713
rect 3016 3607 3023 3673
rect 3036 3623 3043 3673
rect 3056 3647 3063 3973
rect 3076 3763 3083 3996
rect 3113 3987 3127 3993
rect 3176 3885 3183 3973
rect 3176 3847 3183 3871
rect 3113 3820 3127 3833
rect 3116 3816 3123 3820
rect 3096 3780 3103 3783
rect 3093 3767 3107 3780
rect 3076 3756 3093 3763
rect 3036 3616 3063 3623
rect 3056 3516 3063 3616
rect 2836 3376 2853 3383
rect 2676 3296 2683 3333
rect 2713 3300 2727 3313
rect 2716 3296 2723 3300
rect 2796 3296 2803 3373
rect 2836 3307 2843 3333
rect 2576 2996 2603 3003
rect 2633 3000 2647 3013
rect 2696 3008 2703 3133
rect 2636 2996 2643 3000
rect 2376 2896 2403 2903
rect 2136 2796 2163 2803
rect 396 2476 423 2483
rect 156 2267 163 2413
rect 176 2347 183 2443
rect 276 2427 283 2473
rect 416 2446 423 2476
rect 493 2480 507 2493
rect 496 2476 503 2480
rect 556 2446 563 2473
rect 316 2343 323 2443
rect 316 2336 343 2343
rect 56 1963 63 2213
rect 96 2187 103 2223
rect 176 1968 183 2273
rect 336 2123 343 2336
rect 476 2263 483 2443
rect 476 2256 503 2263
rect 356 2227 363 2254
rect 316 2116 343 2123
rect 56 1956 83 1963
rect 116 1956 163 1963
rect 96 1767 103 1923
rect 156 1887 163 1956
rect 316 1963 323 2116
rect 296 1956 323 1963
rect 336 1956 343 2093
rect 356 2047 363 2213
rect 376 1956 383 1993
rect 196 1847 203 1923
rect 236 1743 243 1923
rect 296 1743 303 1956
rect 236 1736 263 1743
rect 36 1167 43 1703
rect 256 1647 263 1736
rect 276 1736 303 1743
rect 336 1736 343 1873
rect 56 1436 83 1443
rect 56 1227 63 1436
rect 176 1287 183 1453
rect 216 1436 223 1593
rect 256 1436 263 1553
rect 276 1467 283 1736
rect 316 1487 323 1692
rect 376 1607 383 1713
rect 396 1706 403 1833
rect 416 1767 423 2033
rect 456 2027 463 2223
rect 496 2187 503 2256
rect 516 2226 523 2293
rect 596 2256 603 2293
rect 676 2287 683 2473
rect 707 2443 720 2447
rect 796 2446 803 2533
rect 836 2476 843 2533
rect 876 2476 883 2513
rect 956 2476 983 2483
rect 1036 2476 1043 2573
rect 936 2446 943 2473
rect 707 2436 723 2443
rect 707 2433 720 2436
rect 633 2260 647 2273
rect 696 2263 703 2293
rect 716 2268 723 2413
rect 636 2256 643 2260
rect 676 2256 703 2263
rect 616 2187 623 2223
rect 676 2167 683 2256
rect 756 2256 763 2293
rect 736 2203 743 2223
rect 776 2220 783 2223
rect 716 2196 743 2203
rect 773 2207 787 2220
rect 816 2207 823 2353
rect 896 2347 903 2443
rect 836 2267 843 2333
rect 956 2307 963 2476
rect 1176 2476 1183 2573
rect 1236 2487 1243 2553
rect 1276 2476 1283 2513
rect 1336 2483 1343 2653
rect 1316 2476 1343 2483
rect 996 2440 1003 2443
rect 993 2427 1007 2440
rect 1136 2407 1143 2443
rect 1296 2407 1303 2443
rect 1356 2427 1363 2473
rect 1336 2416 1353 2423
rect 876 2256 883 2293
rect 907 2276 933 2283
rect 973 2260 987 2273
rect 976 2256 983 2260
rect 847 2223 860 2227
rect 847 2216 863 2223
rect 847 2213 860 2216
rect 413 1747 427 1753
rect 436 1748 443 1913
rect 476 1887 483 1923
rect 516 1887 523 1923
rect 576 1847 583 2093
rect 473 1740 487 1753
rect 596 1747 603 2013
rect 616 1983 623 2152
rect 616 1976 643 1983
rect 636 1956 643 1976
rect 696 1956 703 2013
rect 716 1987 723 2196
rect 936 2167 943 2223
rect 736 1748 743 1993
rect 816 1967 823 2153
rect 956 2147 963 2213
rect 956 2107 963 2133
rect 1036 2087 1043 2273
rect 1056 2226 1063 2253
rect 1236 2226 1243 2313
rect 1296 2256 1303 2353
rect 1336 2267 1343 2416
rect 816 1956 833 1967
rect 820 1953 833 1956
rect 856 1927 863 2073
rect 1156 2027 1163 2223
rect 1356 2187 1363 2293
rect 1376 2207 1383 2673
rect 1576 2527 1583 2743
rect 1656 2736 1683 2743
rect 1736 2567 1743 2732
rect 1816 2667 1823 2743
rect 1876 2587 1883 2743
rect 2096 2740 2103 2743
rect 2016 2627 2023 2732
rect 2093 2727 2107 2740
rect 2136 2727 2143 2796
rect 2216 2776 2223 2813
rect 2156 2746 2163 2773
rect 2396 2747 2403 2896
rect 2516 2887 2523 2963
rect 2453 2863 2467 2873
rect 2576 2867 2583 2996
rect 2736 2963 2743 3193
rect 2716 2956 2743 2963
rect 2453 2860 2483 2863
rect 2456 2856 2483 2860
rect 2416 2827 2423 2853
rect 2476 2776 2483 2856
rect 2236 2727 2243 2743
rect 2296 2740 2303 2743
rect 2293 2727 2307 2740
rect 2636 2743 2643 2853
rect 2716 2776 2723 2956
rect 2756 2788 2763 3273
rect 2787 3003 2800 3007
rect 2787 2996 2803 3003
rect 2836 2996 2843 3253
rect 2856 3207 2863 3373
rect 3076 3367 3083 3693
rect 3096 3467 3103 3633
rect 3116 3527 3123 3593
rect 3136 3516 3143 3613
rect 3156 3607 3163 3783
rect 3176 3707 3183 3812
rect 3196 3763 3203 3993
rect 3216 3987 3223 4053
rect 3236 3967 3243 4153
rect 3256 4127 3263 4173
rect 3276 4107 3283 4153
rect 3296 4147 3303 4293
rect 3296 4087 3303 4133
rect 3316 4087 3323 4303
rect 3336 4187 3343 4273
rect 3356 4147 3363 4303
rect 3396 4296 3423 4303
rect 3256 4047 3263 4073
rect 3313 4040 3327 4052
rect 3316 4036 3323 4040
rect 3376 4007 3383 4273
rect 3396 4103 3403 4273
rect 3416 4167 3423 4296
rect 3436 4167 3443 4233
rect 3456 4187 3463 4303
rect 3496 4300 3503 4303
rect 3493 4287 3507 4300
rect 3496 4247 3503 4273
rect 3536 4263 3543 4353
rect 3576 4336 3583 4413
rect 3596 4387 3603 4593
rect 3616 4567 3623 5073
rect 3636 5007 3643 5033
rect 3736 5007 3743 5053
rect 3756 5027 3763 5193
rect 3816 5076 3823 5333
rect 3836 5127 3843 5473
rect 4127 5456 4163 5463
rect 4013 5380 4027 5393
rect 4053 5387 4067 5393
rect 4016 5376 4023 5380
rect 4076 5367 4083 5413
rect 4136 5388 4143 5433
rect 4156 5427 4163 5456
rect 4316 5376 4323 5413
rect 3856 5088 3863 5333
rect 3876 5227 3883 5273
rect 3896 5147 3903 5343
rect 4076 5307 4083 5332
rect 4156 5287 4163 5343
rect 3996 5147 4003 5253
rect 4216 5187 4223 5373
rect 4236 5167 4243 5333
rect 4256 5287 4263 5343
rect 4296 5247 4303 5343
rect 4356 5327 4363 5522
rect 4396 5376 4403 5413
rect 4496 5346 4503 5413
rect 4656 5403 4663 5523
rect 4636 5396 4663 5403
rect 3876 5087 3883 5113
rect 3896 5047 3903 5093
rect 3956 5076 3963 5133
rect 3993 5080 4007 5093
rect 3996 5076 4003 5080
rect 3716 4856 3723 4913
rect 3656 4627 3663 4813
rect 3696 4787 3703 4823
rect 3653 4560 3667 4573
rect 3656 4556 3663 4560
rect 3736 4526 3743 4812
rect 3776 4607 3783 4993
rect 3796 4987 3803 5043
rect 3836 5040 3843 5043
rect 3833 5027 3847 5040
rect 4036 5046 4043 5153
rect 3796 4907 3803 4973
rect 3916 4927 3923 5033
rect 4056 4967 4063 5093
rect 4113 5080 4127 5093
rect 4116 5076 4123 5080
rect 4236 5076 4243 5153
rect 4273 5080 4287 5093
rect 4316 5087 4323 5313
rect 4416 5247 4423 5343
rect 4456 5307 4463 5332
rect 4356 5088 4363 5113
rect 4416 5107 4423 5133
rect 4276 5076 4283 5080
rect 4336 5076 4353 5083
rect 4196 5046 4203 5073
rect 3896 4867 3903 4893
rect 3936 4867 3943 4953
rect 3996 4868 4003 4893
rect 3836 4747 3843 4823
rect 3896 4767 3903 4813
rect 3916 4787 3923 4853
rect 4020 4823 4033 4827
rect 3976 4820 3983 4823
rect 3973 4807 3987 4820
rect 4016 4813 4033 4823
rect 3996 4727 4003 4753
rect 4016 4747 4023 4813
rect 3767 4583 3780 4587
rect 3767 4573 3783 4583
rect 3776 4556 3783 4573
rect 3896 4556 3903 4613
rect 3836 4526 3843 4553
rect 3936 4526 3943 4593
rect 3996 4556 4003 4613
rect 4036 4556 4043 4673
rect 4056 4567 4063 4932
rect 4096 4883 4103 5043
rect 4076 4880 4123 4883
rect 4073 4876 4123 4880
rect 4073 4867 4087 4876
rect 4116 4856 4123 4876
rect 4160 4863 4173 4867
rect 4156 4856 4173 4863
rect 4160 4853 4173 4856
rect 4160 4848 4166 4853
rect 4092 4829 4106 4834
rect 4087 4793 4093 4807
rect 4076 4667 4083 4713
rect 4176 4687 4183 4813
rect 4196 4767 4203 4953
rect 4256 4856 4263 4993
rect 4296 4868 4303 5043
rect 4316 4967 4323 5033
rect 4336 4987 4343 5076
rect 4456 5087 4463 5173
rect 4356 4907 4363 4953
rect 4376 4883 4383 5043
rect 4413 5027 4427 5032
rect 4336 4876 4383 4883
rect 3616 4487 3623 4513
rect 3636 4447 3643 4523
rect 3676 4427 3683 4523
rect 3656 4347 3663 4413
rect 3596 4300 3603 4303
rect 3553 4287 3567 4293
rect 3593 4287 3607 4300
rect 3676 4287 3683 4413
rect 3736 4348 3743 4512
rect 3716 4300 3723 4303
rect 3713 4287 3727 4300
rect 3536 4256 3563 4263
rect 3516 4223 3523 4253
rect 3487 4216 3523 4223
rect 3396 4096 3413 4103
rect 3393 4047 3407 4053
rect 3416 4036 3423 4093
rect 3456 4047 3463 4133
rect 3476 4027 3483 4192
rect 3516 4067 3523 4173
rect 3536 4107 3543 4213
rect 3556 4147 3563 4256
rect 3533 4040 3547 4053
rect 3536 4036 3543 4040
rect 3576 4036 3583 4093
rect 3596 4047 3603 4133
rect 3616 4107 3623 4253
rect 3236 3828 3243 3932
rect 3256 3847 3263 3913
rect 3276 3816 3283 3973
rect 3336 3847 3343 3953
rect 3196 3756 3213 3763
rect 3216 3627 3223 3753
rect 3176 3516 3183 3593
rect 2876 3307 2883 3353
rect 2993 3307 3007 3313
rect 2856 3147 2863 3193
rect 2896 3187 2903 3263
rect 2916 3107 2923 3153
rect 2936 3107 2943 3252
rect 2976 3247 2983 3293
rect 3016 3260 3023 3263
rect 3013 3247 3027 3260
rect 3056 3227 3063 3263
rect 3116 3247 3123 3473
rect 3136 3263 3143 3453
rect 3156 3447 3163 3483
rect 3176 3367 3183 3433
rect 3196 3347 3203 3393
rect 3216 3303 3223 3613
rect 3236 3363 3243 3713
rect 3256 3528 3263 3751
rect 3336 3647 3343 3833
rect 3356 3827 3363 3993
rect 3436 3963 3443 3992
rect 3496 3967 3503 3993
rect 3416 3960 3443 3963
rect 3413 3956 3443 3960
rect 3413 3947 3427 3956
rect 3516 3923 3523 4003
rect 3516 3916 3543 3923
rect 3436 3827 3443 3873
rect 3456 3847 3463 3893
rect 3516 3816 3523 3893
rect 3536 3867 3543 3916
rect 3376 3780 3383 3783
rect 3296 3516 3303 3573
rect 3356 3523 3363 3773
rect 3373 3767 3387 3780
rect 3416 3763 3423 3783
rect 3396 3756 3423 3763
rect 3336 3516 3363 3523
rect 3376 3487 3383 3732
rect 3396 3647 3403 3756
rect 3496 3747 3503 3783
rect 3436 3607 3443 3633
rect 3456 3528 3463 3573
rect 3276 3407 3283 3483
rect 3396 3447 3403 3473
rect 3436 3407 3443 3483
rect 3236 3356 3253 3363
rect 3216 3296 3233 3303
rect 3236 3267 3243 3294
rect 3136 3256 3163 3263
rect 2956 3187 2963 3213
rect 2787 2993 2800 2996
rect 2976 3003 2983 3212
rect 2956 2996 2983 3003
rect 2816 2960 2823 2963
rect 2773 2947 2787 2953
rect 2813 2947 2827 2960
rect 2856 2847 2863 2963
rect 2596 2736 2643 2743
rect 2236 2567 2243 2713
rect 1553 2480 1567 2493
rect 1556 2476 1563 2480
rect 1436 2387 1443 2443
rect 1536 2347 1543 2443
rect 1596 2407 1603 2493
rect 1636 2476 1663 2483
rect 1776 2476 1783 2513
rect 1456 2256 1463 2293
rect 1616 2226 1623 2293
rect 1436 2220 1443 2223
rect 1396 2147 1403 2213
rect 1433 2207 1447 2220
rect 1516 2220 1523 2223
rect 1513 2207 1527 2220
rect 1576 2216 1603 2223
rect 1596 2187 1603 2216
rect 1636 2207 1643 2476
rect 2016 2476 2063 2483
rect 1836 2407 1843 2443
rect 1916 2387 1923 2474
rect 2056 2427 2063 2476
rect 2153 2480 2167 2493
rect 2156 2476 2163 2480
rect 2376 2476 2403 2483
rect 2076 2407 2083 2473
rect 2196 2447 2203 2474
rect 2256 2387 2263 2443
rect 2356 2403 2363 2474
rect 2376 2427 2383 2476
rect 2513 2480 2527 2493
rect 2516 2476 2523 2480
rect 2356 2396 2383 2403
rect 2067 2386 2080 2387
rect 2067 2373 2073 2386
rect 2107 2373 2113 2387
rect 1736 2287 1743 2333
rect 1816 2256 1823 2293
rect 1876 2268 1883 2313
rect 1736 2227 1743 2252
rect 913 1960 927 1973
rect 953 1967 967 1973
rect 916 1956 923 1960
rect 476 1736 483 1740
rect 747 1736 763 1743
rect 416 1567 423 1693
rect 456 1507 463 1703
rect 576 1696 603 1703
rect 596 1647 603 1696
rect 476 1463 483 1533
rect 456 1456 483 1463
rect 456 1436 463 1456
rect 496 1436 503 1513
rect 67 1216 83 1223
rect 256 1227 263 1273
rect 136 1187 143 1214
rect 296 1223 303 1433
rect 356 1347 363 1403
rect 396 1287 403 1433
rect 536 1406 543 1493
rect 616 1447 623 1513
rect 676 1436 683 1473
rect 393 1267 407 1273
rect 276 1216 303 1223
rect 313 1220 327 1233
rect 316 1216 323 1220
rect 356 1216 363 1253
rect 36 567 43 1153
rect 56 927 63 1173
rect 276 1186 283 1216
rect 436 1216 443 1403
rect 476 1347 483 1392
rect 636 1367 643 1413
rect 136 886 143 1173
rect 196 1163 203 1183
rect 196 1156 223 1163
rect 216 928 223 1156
rect 260 923 273 927
rect 256 916 273 923
rect 260 913 273 916
rect 56 703 63 873
rect 76 787 83 883
rect 56 696 83 703
rect 116 696 123 773
rect 236 747 243 883
rect 156 666 163 733
rect 296 727 303 1173
rect 396 1007 403 1213
rect 396 947 403 993
rect 353 920 367 933
rect 356 916 363 920
rect 416 916 423 973
rect 316 847 323 913
rect 456 907 463 933
rect 476 923 483 993
rect 496 947 503 1273
rect 596 1216 603 1253
rect 696 1243 703 1403
rect 756 1307 763 1736
rect 836 1736 843 1773
rect 876 1767 883 1913
rect 956 1787 963 1913
rect 976 1763 983 1954
rect 1256 1956 1263 2013
rect 913 1740 927 1753
rect 956 1756 983 1763
rect 916 1736 923 1740
rect 956 1736 963 1756
rect 976 1743 983 1756
rect 1096 1748 1103 1773
rect 1136 1748 1143 1793
rect 1156 1783 1163 1953
rect 1316 1916 1424 1923
rect 1156 1776 1183 1783
rect 976 1736 1003 1743
rect 776 1547 783 1693
rect 816 1527 823 1703
rect 996 1687 1003 1736
rect 1176 1736 1183 1776
rect 1236 1736 1243 1773
rect 1056 1667 1063 1703
rect 1073 1687 1087 1693
rect 1056 1587 1063 1653
rect 776 1447 783 1473
rect 813 1440 827 1453
rect 816 1436 823 1440
rect 836 1367 843 1403
rect 836 1327 843 1353
rect 876 1303 883 1453
rect 936 1448 943 1513
rect 916 1367 923 1403
rect 856 1296 883 1303
rect 676 1236 703 1243
rect 676 1216 683 1236
rect 816 1223 823 1293
rect 816 1216 843 1223
rect 536 967 543 1183
rect 476 916 503 923
rect 447 893 463 907
rect 456 886 463 893
rect 256 627 263 663
rect 296 567 303 663
rect 216 396 223 453
rect 96 188 103 363
rect 196 267 203 352
rect 236 183 243 363
rect 296 323 303 553
rect 356 396 363 433
rect 396 408 403 713
rect 416 467 423 833
rect 536 747 543 853
rect 596 787 603 953
rect 636 916 643 973
rect 696 947 703 1183
rect 736 1180 743 1183
rect 733 1167 747 1180
rect 736 1107 743 1153
rect 716 916 723 973
rect 516 627 523 693
rect 616 660 623 663
rect 576 587 583 652
rect 613 647 627 660
rect 416 366 423 432
rect 556 396 563 433
rect 593 400 607 413
rect 596 396 603 400
rect 276 316 303 323
rect 236 176 263 183
rect 256 146 263 176
rect 216 47 223 143
rect 276 47 283 316
rect 336 207 343 363
rect 376 356 403 363
rect 396 327 403 356
rect 636 347 643 393
rect 356 176 363 213
rect 396 147 403 313
rect 656 307 663 773
rect 696 747 703 883
rect 676 736 693 743
rect 676 647 683 736
rect 756 727 763 933
rect 796 916 803 973
rect 836 928 843 1216
rect 816 863 823 883
rect 796 856 823 863
rect 713 700 727 713
rect 776 703 783 753
rect 716 696 723 700
rect 756 696 783 703
rect 796 696 803 856
rect 836 787 843 873
rect 856 767 863 1296
rect 916 1267 923 1353
rect 976 1347 983 1573
rect 1096 1443 1103 1734
rect 1296 1706 1303 1813
rect 1156 1700 1163 1703
rect 1116 1507 1123 1693
rect 1153 1687 1167 1700
rect 1316 1647 1323 1916
rect 1456 1703 1463 1753
rect 1416 1696 1463 1703
rect 1096 1436 1113 1443
rect 1196 1436 1203 1513
rect 1236 1447 1243 1633
rect 1476 1627 1483 1954
rect 1496 1767 1503 2013
rect 1596 1968 1603 2013
rect 1636 1968 1643 2193
rect 1736 2027 1743 2192
rect 1596 1807 1603 1873
rect 1656 1803 1663 2013
rect 1713 1960 1727 1973
rect 1753 1960 1767 1973
rect 1796 1963 1803 2212
rect 1836 2147 1843 2223
rect 1716 1956 1723 1960
rect 1756 1956 1763 1960
rect 1796 1956 1823 1963
rect 1836 1956 1843 2133
rect 1956 2087 1963 2353
rect 2096 2226 2103 2293
rect 2296 2256 2303 2293
rect 2116 2227 2123 2254
rect 2056 2187 2063 2223
rect 2196 2220 2203 2223
rect 2193 2207 2207 2220
rect 1696 1887 1703 1923
rect 1796 1887 1803 1933
rect 1816 1807 1823 1956
rect 1876 1916 1903 1923
rect 1636 1796 1663 1803
rect 1596 1736 1603 1793
rect 1496 1707 1503 1732
rect 1536 1667 1543 1703
rect 1576 1700 1583 1703
rect 1573 1687 1587 1700
rect 1636 1667 1643 1796
rect 996 1223 1003 1433
rect 1116 1407 1123 1434
rect 1216 1407 1226 1413
rect 1216 1393 1233 1407
rect 976 1216 1003 1223
rect 976 1186 983 1216
rect 1116 1216 1123 1253
rect 1193 1220 1207 1233
rect 1196 1216 1203 1220
rect 1036 1147 1043 1183
rect 1236 1147 1243 1233
rect 1256 1227 1263 1493
rect 1276 1447 1283 1473
rect 1356 1436 1363 1613
rect 1476 1436 1483 1473
rect 1576 1436 1583 1513
rect 1396 1407 1403 1434
rect 1276 1367 1283 1393
rect 1296 1347 1303 1403
rect 1656 1406 1663 1773
rect 1716 1736 1723 1793
rect 1756 1703 1763 1734
rect 1776 1706 1783 1793
rect 1836 1736 1843 1773
rect 1676 1436 1683 1703
rect 1736 1696 1763 1703
rect 1896 1667 1903 1916
rect 1916 1747 1923 1923
rect 1976 1887 1983 1973
rect 2096 1956 2103 2173
rect 2236 2087 2243 2254
rect 2316 2220 2323 2223
rect 2313 2207 2327 2220
rect 2376 2203 2383 2396
rect 2436 2256 2443 2474
rect 2456 2387 2463 2432
rect 2556 2287 2563 2553
rect 2576 2507 2583 2653
rect 2456 2220 2463 2223
rect 2376 2196 2393 2203
rect 2156 2047 2163 2073
rect 1996 1867 2003 1933
rect 2156 1926 2163 2033
rect 1996 1567 2003 1793
rect 2016 1787 2023 1913
rect 2036 1736 2043 1853
rect 2156 1807 2163 1912
rect 2176 1867 2183 1953
rect 2336 1887 2343 1923
rect 2076 1736 2083 1773
rect 2136 1706 2143 1733
rect 2156 1696 2183 1703
rect 2216 1700 2223 1703
rect 1736 1436 1743 1473
rect 1956 1436 2003 1443
rect 1296 1216 1303 1253
rect 1316 1247 1323 1353
rect 1336 1216 1343 1333
rect 1456 1267 1463 1403
rect 1556 1400 1563 1403
rect 1553 1387 1567 1400
rect 1496 1327 1503 1373
rect 1553 1367 1567 1373
rect 1636 1396 1653 1403
rect 1396 1186 1403 1253
rect 1476 1216 1483 1273
rect 1500 1183 1513 1187
rect 1496 1176 1513 1183
rect 1500 1173 1513 1176
rect 1356 1107 1363 1133
rect 1053 920 1067 933
rect 1056 916 1063 920
rect 876 867 883 913
rect 996 887 1003 914
rect 936 847 943 883
rect 1036 880 1043 883
rect 716 396 723 493
rect 736 427 743 663
rect 856 396 863 713
rect 876 666 883 773
rect 996 707 1003 873
rect 1033 867 1047 880
rect 1156 847 1163 883
rect 1027 836 1053 843
rect 1216 767 1223 913
rect 1336 883 1343 933
rect 1413 920 1427 933
rect 1416 916 1423 920
rect 1296 876 1343 883
rect 1476 886 1483 993
rect 1536 947 1543 1313
rect 1553 1267 1567 1273
rect 1553 1260 1573 1267
rect 1556 1256 1573 1260
rect 1560 1253 1573 1256
rect 1553 1227 1567 1233
rect 1636 1227 1643 1396
rect 1776 1367 1783 1403
rect 1996 1307 2003 1436
rect 1496 916 1523 923
rect 1356 847 1363 873
rect 1396 787 1403 883
rect 1496 847 1503 916
rect 1507 836 1523 843
rect 976 567 983 663
rect 893 400 907 413
rect 896 396 903 400
rect 796 363 803 394
rect 936 363 943 453
rect 1016 447 1023 653
rect 1036 567 1043 663
rect 1096 656 1123 663
rect 1116 607 1123 656
rect 1256 527 1263 673
rect 1276 647 1283 773
rect 1316 696 1323 753
rect 1336 567 1343 663
rect 1376 607 1383 694
rect 1436 660 1443 663
rect 1433 647 1447 660
rect 736 307 743 363
rect 796 356 843 363
rect 847 333 853 347
rect 876 327 883 363
rect 916 356 943 363
rect 956 363 963 413
rect 956 356 983 363
rect 916 283 923 356
rect 947 333 953 347
rect 907 276 923 283
rect 436 176 443 253
rect 576 176 583 213
rect 616 176 623 213
rect 896 176 903 273
rect 516 146 523 173
rect 696 147 703 174
rect 996 146 1003 233
rect 1096 188 1103 433
rect 1116 327 1123 413
rect 1236 366 1243 413
rect 1256 407 1263 513
rect 1287 423 1300 427
rect 1287 413 1303 423
rect 1296 396 1303 413
rect 1156 307 1163 363
rect 1256 307 1263 333
rect 1316 307 1323 363
rect 1356 327 1363 593
rect 1516 427 1523 836
rect 1576 827 1583 1172
rect 1616 1107 1623 1183
rect 1756 1186 1763 1253
rect 1636 1007 1643 1173
rect 1656 1147 1663 1183
rect 1776 1107 1783 1214
rect 1996 1186 2003 1253
rect 1896 1107 1903 1183
rect 1636 916 1643 993
rect 1676 916 1683 953
rect 1816 928 1823 953
rect 1596 847 1603 893
rect 1876 886 1883 1013
rect 2016 1007 2023 1473
rect 2076 1436 2083 1513
rect 2056 1307 2063 1403
rect 2136 1307 2143 1373
rect 2116 1107 2123 1273
rect 2156 1223 2163 1696
rect 2213 1687 2227 1700
rect 2176 1403 2183 1553
rect 2176 1396 2203 1403
rect 2196 1327 2203 1396
rect 2256 1387 2263 1853
rect 2396 1827 2403 2193
rect 2416 1968 2423 2212
rect 2453 2207 2467 2220
rect 2456 1956 2463 1993
rect 2316 1736 2323 1813
rect 2376 1736 2383 1793
rect 2296 1687 2303 1703
rect 2276 1363 2283 1653
rect 2296 1447 2303 1673
rect 2336 1647 2343 1703
rect 2436 1547 2443 1912
rect 2476 1887 2483 1923
rect 2576 1923 2583 2493
rect 2636 2347 2643 2443
rect 2676 2367 2683 2443
rect 2596 2267 2603 2333
rect 2716 2226 2723 2413
rect 2816 2307 2823 2773
rect 2876 2747 2883 2953
rect 2836 2707 2843 2732
rect 2956 2667 2963 2743
rect 2996 2667 3003 3073
rect 3016 2947 3023 3033
rect 3116 2887 3123 3233
rect 3136 2847 3143 3093
rect 3156 3087 3163 3256
rect 3176 3227 3183 3263
rect 3256 3227 3263 3353
rect 3353 3307 3367 3313
rect 3287 3256 3303 3263
rect 3276 3207 3283 3253
rect 3196 2996 3203 3153
rect 3136 2743 3143 2833
rect 3176 2747 3183 2963
rect 3216 2927 3223 2963
rect 3276 2947 3283 3193
rect 3336 3107 3343 3252
rect 3376 3147 3383 3333
rect 3456 3296 3463 3333
rect 3496 3307 3503 3553
rect 3556 3516 3563 3593
rect 3576 3547 3583 3773
rect 3596 3567 3603 3993
rect 3616 3783 3623 4072
rect 3676 4067 3683 4133
rect 3736 4087 3743 4273
rect 3756 4167 3763 4253
rect 3673 4040 3687 4053
rect 3676 4036 3683 4040
rect 3776 4047 3783 4253
rect 3636 3887 3643 3993
rect 3656 3967 3663 4003
rect 3696 4000 3703 4003
rect 3693 3987 3707 4000
rect 3656 3816 3663 3913
rect 3616 3780 3643 3783
rect 3616 3776 3647 3780
rect 3633 3767 3647 3776
rect 3536 3307 3543 3483
rect 3576 3480 3583 3483
rect 3573 3467 3587 3480
rect 3616 3407 3623 3473
rect 3636 3467 3643 3673
rect 3676 3567 3683 3633
rect 3696 3627 3703 3783
rect 3716 3567 3723 3853
rect 3676 3516 3683 3553
rect 3736 3543 3743 3993
rect 3756 3947 3763 4034
rect 3796 4036 3803 4173
rect 3816 4067 3823 4373
rect 3916 4367 3923 4493
rect 3876 4300 3883 4303
rect 3873 4287 3887 4300
rect 3836 4207 3843 4253
rect 3916 4167 3923 4303
rect 3936 4207 3943 4293
rect 3896 4156 3913 4163
rect 3856 4107 3863 4153
rect 3836 4036 3843 4073
rect 3816 3967 3823 4003
rect 3876 4006 3883 4133
rect 3896 4047 3903 4156
rect 3956 4163 3963 4453
rect 3976 4287 3983 4523
rect 4016 4487 4023 4512
rect 4036 4467 4043 4493
rect 4056 4343 4063 4513
rect 4076 4507 4083 4573
rect 4096 4547 4103 4633
rect 4176 4583 4183 4673
rect 4216 4667 4223 4813
rect 4236 4787 4243 4823
rect 4336 4826 4343 4876
rect 4436 4863 4443 4973
rect 4476 4868 4483 5133
rect 4496 5107 4503 5173
rect 4516 5103 4523 5373
rect 4536 5307 4543 5343
rect 4536 5207 4543 5293
rect 4596 5207 4603 5343
rect 4616 5267 4623 5353
rect 4616 5187 4623 5213
rect 4516 5096 4543 5103
rect 4536 5088 4543 5096
rect 4576 5076 4583 5113
rect 4516 4967 4523 5043
rect 4560 5003 4573 5007
rect 4556 5000 4573 5003
rect 4553 4993 4573 5000
rect 4636 5003 4643 5396
rect 4696 5376 4703 5433
rect 4856 5376 4863 5413
rect 4776 5343 4783 5373
rect 4676 5307 4683 5343
rect 4716 5340 4723 5343
rect 4713 5327 4727 5340
rect 4776 5336 4803 5343
rect 4776 5083 4783 5313
rect 4796 5147 4803 5336
rect 4836 5323 4843 5343
rect 4876 5340 4883 5343
rect 4873 5327 4887 5340
rect 4916 5327 4923 5433
rect 4936 5395 4943 5523
rect 4936 5388 4983 5395
rect 4836 5316 4863 5323
rect 4836 5088 4843 5173
rect 4696 5076 4723 5083
rect 4716 5046 4723 5076
rect 4756 5076 4783 5083
rect 4656 5007 4663 5043
rect 4636 4996 4653 5003
rect 4553 4987 4567 4993
rect 4756 4927 4763 5076
rect 4856 5067 4863 5316
rect 4936 5107 4943 5388
rect 4976 5371 4983 5388
rect 4956 5287 4963 5353
rect 4996 5207 5003 5293
rect 5016 5267 5023 5332
rect 4416 4856 4443 4863
rect 4156 4576 4183 4583
rect 4156 4556 4163 4576
rect 4196 4556 4203 4613
rect 4216 4568 4223 4653
rect 4036 4336 4063 4343
rect 4076 4323 4083 4453
rect 4136 4387 4143 4523
rect 4176 4487 4183 4523
rect 4056 4316 4083 4323
rect 3996 4267 4003 4303
rect 3936 4156 3963 4163
rect 3936 4036 3943 4156
rect 3976 4036 3983 4093
rect 3996 4047 4003 4213
rect 4056 4167 4063 4316
rect 4076 4267 4083 4293
rect 4076 4207 4083 4232
rect 4096 4187 4103 4373
rect 4153 4340 4167 4353
rect 4156 4336 4163 4340
rect 4116 4267 4123 4303
rect 4113 4247 4127 4253
rect 4136 4127 4143 4173
rect 4076 4087 4083 4113
rect 4096 4036 4103 4073
rect 3796 3847 3803 3913
rect 3856 3816 3863 3993
rect 3876 3903 3883 3953
rect 3996 3927 4003 3993
rect 4016 3967 4023 4034
rect 4136 3967 4143 3993
rect 3876 3896 3903 3903
rect 3896 3883 3903 3896
rect 3896 3876 3923 3883
rect 3876 3827 3883 3873
rect 3716 3536 3743 3543
rect 3716 3516 3723 3536
rect 3776 3527 3783 3773
rect 3796 3763 3803 3783
rect 3796 3756 3823 3763
rect 3773 3487 3787 3492
rect 3747 3476 3763 3483
rect 3556 3296 3563 3353
rect 3596 3296 3603 3333
rect 3356 3027 3363 3133
rect 3396 3127 3403 3233
rect 3476 3243 3483 3263
rect 3447 3236 3483 3243
rect 3313 3000 3327 3013
rect 3316 2996 3323 3000
rect 3356 2996 3363 3013
rect 3373 2943 3387 2953
rect 3356 2940 3387 2943
rect 3356 2936 3383 2940
rect 3356 2827 3363 2936
rect 3116 2736 3143 2743
rect 3247 2736 3263 2743
rect 3156 2527 3163 2613
rect 3256 2607 3263 2736
rect 3276 2707 3283 2743
rect 3336 2736 3363 2743
rect 2836 2407 2843 2474
rect 2936 2446 2943 2513
rect 3156 2476 3163 2513
rect 2736 2127 2743 2253
rect 2576 1916 2603 1923
rect 2456 1706 2463 1753
rect 2476 1747 2483 1873
rect 2556 1700 2563 1703
rect 2553 1687 2567 1700
rect 2356 1436 2363 1533
rect 2396 1387 2403 1403
rect 2456 1387 2463 1633
rect 2576 1436 2583 1673
rect 2596 1547 2603 1916
rect 2256 1356 2283 1363
rect 2196 1287 2203 1313
rect 2187 1256 2243 1263
rect 2156 1216 2173 1223
rect 2213 1220 2227 1233
rect 2236 1227 2243 1256
rect 2216 1216 2223 1220
rect 1536 747 1543 813
rect 1413 400 1427 413
rect 1536 408 1543 733
rect 1576 696 1583 733
rect 1616 696 1623 773
rect 1636 707 1643 853
rect 1656 666 1663 883
rect 1696 787 1703 872
rect 1796 763 1803 883
rect 1836 763 1843 872
rect 1916 807 1923 872
rect 1796 756 1823 763
rect 1836 756 1863 763
rect 1753 740 1767 753
rect 1756 736 1763 740
rect 1596 627 1603 663
rect 1556 547 1563 573
rect 1576 487 1583 593
rect 1676 567 1683 733
rect 1816 723 1823 756
rect 1816 716 1843 723
rect 1796 696 1823 703
rect 1796 547 1803 593
rect 1816 567 1823 696
rect 1416 396 1423 400
rect 1576 396 1583 473
rect 1496 367 1503 394
rect 1436 327 1443 363
rect 1716 363 1723 493
rect 1696 356 1723 363
rect 1456 207 1463 253
rect 1453 180 1467 193
rect 1456 176 1463 180
rect 1356 147 1363 174
rect 1556 176 1563 233
rect 556 107 563 132
rect 796 47 803 143
rect 916 107 923 143
rect 1056 140 1063 143
rect 1053 127 1067 140
rect 1276 47 1283 143
rect 1396 87 1403 143
rect 1436 107 1443 143
rect 1496 87 1503 173
rect 1616 143 1623 233
rect 1736 207 1743 413
rect 1773 400 1787 413
rect 1776 396 1783 400
rect 1816 396 1823 513
rect 1836 427 1843 716
rect 1856 707 1863 756
rect 1916 707 1923 753
rect 1896 607 1903 633
rect 1936 543 1943 733
rect 1976 708 1983 993
rect 2016 916 2023 972
rect 2016 696 2023 793
rect 2036 707 2043 883
rect 2096 747 2103 1053
rect 2136 916 2143 1113
rect 2256 1067 2263 1356
rect 2156 827 2163 883
rect 2216 847 2223 883
rect 2276 847 2283 1273
rect 2353 1220 2367 1233
rect 2396 1227 2403 1373
rect 2356 1216 2363 1220
rect 2416 1183 2423 1233
rect 2376 1007 2383 1183
rect 2416 1176 2443 1183
rect 2333 920 2347 933
rect 2396 928 2403 1093
rect 2336 916 2343 920
rect 2296 847 2303 914
rect 1953 647 1967 653
rect 1916 536 1943 543
rect 1916 507 1923 536
rect 1796 283 1803 363
rect 1836 307 1843 352
rect 1796 276 1853 283
rect 1736 146 1743 193
rect 1876 146 1883 253
rect 1536 140 1543 143
rect 1533 127 1547 140
rect 1576 136 1623 143
rect 1696 107 1703 143
rect 1796 47 1803 143
rect 1896 47 1903 413
rect 1916 327 1923 433
rect 1936 396 1943 513
rect 1996 447 2003 663
rect 2066 653 2067 660
rect 2296 666 2303 733
rect 2396 707 2403 733
rect 2116 660 2123 663
rect 2053 647 2067 653
rect 1986 433 1987 440
rect 1973 423 1987 433
rect 1973 420 2003 423
rect 1976 416 2003 420
rect 1996 396 2003 416
rect 2016 267 2023 593
rect 2056 507 2063 612
rect 2076 587 2083 653
rect 2113 647 2127 660
rect 2196 607 2203 663
rect 2256 656 2283 663
rect 2276 627 2283 656
rect 2316 627 2323 693
rect 2416 607 2423 873
rect 2436 807 2443 1176
rect 2496 1180 2503 1183
rect 2493 1167 2507 1180
rect 2536 1167 2543 1313
rect 2596 1216 2603 1393
rect 2616 1327 2623 1813
rect 2736 1787 2743 2073
rect 2653 1740 2667 1753
rect 2656 1736 2663 1740
rect 2696 1736 2703 1773
rect 2636 1247 2643 1693
rect 2676 1667 2683 1703
rect 2656 1223 2663 1613
rect 2716 1436 2723 1692
rect 2736 1323 2743 1593
rect 2756 1406 2763 2293
rect 2816 2187 2823 2223
rect 2856 2220 2863 2223
rect 2853 2207 2867 2220
rect 2956 2187 2963 2453
rect 2976 2347 2983 2432
rect 3056 2407 3063 2443
rect 3116 2407 3123 2474
rect 3256 2446 3263 2593
rect 3356 2587 3363 2736
rect 3376 2567 3383 2913
rect 3396 2847 3403 3013
rect 3416 3007 3423 3093
rect 3496 3067 3503 3253
rect 3453 3000 3467 3013
rect 3456 2996 3463 3000
rect 3516 3007 3523 3293
rect 3616 3256 3643 3263
rect 3613 3227 3627 3233
rect 3476 2887 3483 2963
rect 3396 2447 3403 2573
rect 3456 2476 3463 2653
rect 3496 2607 3503 2774
rect 3496 2476 3503 2593
rect 3516 2587 3523 2953
rect 3536 2787 3543 3013
rect 3556 3008 3563 3193
rect 3616 3167 3623 3213
rect 3636 3207 3643 3256
rect 3576 2996 3583 3093
rect 3616 2996 3623 3153
rect 3656 3067 3663 3333
rect 3676 3307 3683 3433
rect 3696 3387 3703 3472
rect 3756 3307 3763 3476
rect 3796 3467 3803 3593
rect 3816 3527 3823 3756
rect 3896 3607 3903 3853
rect 3916 3786 3923 3876
rect 3927 3776 3943 3783
rect 4036 3627 4043 3693
rect 4056 3667 4063 3833
rect 4076 3786 4083 3953
rect 4156 3847 4163 4273
rect 4176 4107 4183 4303
rect 4216 4107 4223 4453
rect 4236 4287 4243 4713
rect 4316 4556 4323 4813
rect 4356 4563 4363 4853
rect 4376 4743 4383 4823
rect 4436 4807 4443 4856
rect 4556 4867 4563 4893
rect 4496 4787 4503 4823
rect 4427 4783 4440 4787
rect 4427 4773 4443 4783
rect 4376 4736 4403 4743
rect 4376 4687 4383 4713
rect 4396 4607 4403 4736
rect 4436 4727 4443 4773
rect 4356 4556 4383 4563
rect 4376 4527 4383 4556
rect 4396 4547 4403 4593
rect 4476 4587 4483 4733
rect 4496 4687 4503 4773
rect 4416 4556 4443 4563
rect 4416 4527 4423 4556
rect 4296 4427 4303 4523
rect 4376 4407 4383 4492
rect 4416 4367 4423 4473
rect 4456 4368 4463 4393
rect 4476 4367 4483 4433
rect 4416 4336 4423 4353
rect 4496 4347 4503 4553
rect 4516 4527 4523 4793
rect 4536 4567 4543 4823
rect 4556 4787 4563 4813
rect 4576 4647 4583 4913
rect 4596 4867 4603 4893
rect 4776 4856 4783 4953
rect 4876 4947 4883 5093
rect 4996 5076 5003 5193
rect 5016 5167 5023 5253
rect 5016 5087 5023 5153
rect 5056 5107 5063 5373
rect 5096 5307 5103 5343
rect 5113 5107 5127 5113
rect 5176 5107 5183 5393
rect 5353 5380 5367 5393
rect 5356 5376 5363 5380
rect 4936 5027 4943 5043
rect 4876 4883 4883 4933
rect 4856 4880 4883 4883
rect 4853 4876 4883 4880
rect 4636 4820 4643 4823
rect 4596 4627 4603 4813
rect 4633 4807 4647 4820
rect 4676 4767 4683 4823
rect 4556 4588 4563 4613
rect 4636 4587 4643 4693
rect 4627 4576 4643 4587
rect 4653 4587 4667 4593
rect 4627 4573 4640 4576
rect 4593 4560 4607 4573
rect 4596 4556 4603 4560
rect 4676 4556 4683 4732
rect 4716 4727 4723 4853
rect 4836 4826 4843 4873
rect 4853 4867 4867 4876
rect 4866 4860 4867 4867
rect 4716 4567 4723 4633
rect 4236 4147 4243 4193
rect 4216 4096 4233 4107
rect 4220 4093 4233 4096
rect 4176 4047 4183 4093
rect 4187 4036 4203 4043
rect 4233 4040 4247 4053
rect 4256 4047 4263 4293
rect 4276 4267 4283 4303
rect 4316 4300 4323 4303
rect 4313 4287 4327 4300
rect 4236 4036 4243 4040
rect 4176 3827 4183 3993
rect 4216 3983 4223 4003
rect 4216 3976 4243 3983
rect 4196 3887 4203 3913
rect 4196 3763 4203 3813
rect 4176 3760 4203 3763
rect 4173 3756 4203 3760
rect 4016 3516 4023 3573
rect 4056 3516 4063 3653
rect 3936 3476 3963 3483
rect 3796 3323 3803 3373
rect 3836 3323 3843 3453
rect 3956 3427 3963 3476
rect 3976 3323 3983 3513
rect 3996 3387 4003 3413
rect 4013 3323 4027 3333
rect 4036 3327 4043 3483
rect 3796 3316 3823 3323
rect 3836 3316 3863 3323
rect 3816 3296 3823 3316
rect 3856 3296 3863 3316
rect 3956 3316 3983 3323
rect 3996 3320 4027 3323
rect 3996 3316 4023 3320
rect 3956 3308 3963 3316
rect 3996 3296 4003 3316
rect 3696 3260 3703 3263
rect 3693 3247 3707 3260
rect 3747 3256 3763 3263
rect 3636 2783 3643 2833
rect 3656 2807 3663 3032
rect 3696 3008 3703 3093
rect 3733 3023 3747 3033
rect 3756 3023 3763 3256
rect 3776 3207 3783 3293
rect 3896 3266 3903 3293
rect 3796 3187 3803 3253
rect 3733 3020 3763 3023
rect 3736 3016 3763 3020
rect 3736 2996 3743 3016
rect 3716 2907 3723 2963
rect 3696 2816 3763 2823
rect 3696 2803 3703 2816
rect 3676 2800 3703 2803
rect 3673 2796 3703 2800
rect 3673 2787 3687 2796
rect 3636 2776 3663 2783
rect 3596 2667 3603 2743
rect 3636 2627 3643 2733
rect 3656 2727 3663 2776
rect 3713 2780 3727 2793
rect 3716 2776 3723 2780
rect 3756 2776 3763 2816
rect 3776 2783 3783 3033
rect 3796 3027 3803 3173
rect 3836 3047 3843 3263
rect 3856 3107 3863 3173
rect 3936 3167 3943 3263
rect 3976 3243 3983 3263
rect 3976 3236 4003 3243
rect 3816 2927 3823 2963
rect 3776 2776 3803 2783
rect 3856 2776 3863 2833
rect 3876 2807 3883 3013
rect 3916 2996 3923 3053
rect 3956 2996 3963 3233
rect 3996 3127 4003 3236
rect 4016 3207 4023 3263
rect 4036 3143 4043 3253
rect 4056 3167 4063 3373
rect 4096 3323 4103 3733
rect 4156 3647 4163 3751
rect 4173 3747 4187 3756
rect 4186 3740 4187 3747
rect 4196 3567 4203 3733
rect 4216 3603 4223 3953
rect 4236 3867 4243 3976
rect 4256 3828 4263 3993
rect 4276 3967 4283 4253
rect 4336 4227 4343 4253
rect 4356 4227 4363 4333
rect 4454 4328 4468 4333
rect 4396 4147 4403 4292
rect 4436 4147 4443 4303
rect 4296 3947 4303 4053
rect 4316 4036 4323 4133
rect 4393 4127 4407 4133
rect 4496 4127 4503 4213
rect 4516 4207 4523 4413
rect 4536 4407 4543 4513
rect 4556 4367 4563 4493
rect 4576 4423 4583 4523
rect 4636 4507 4643 4553
rect 4736 4526 4743 4593
rect 4756 4567 4763 4812
rect 4796 4707 4803 4823
rect 4776 4556 4783 4593
rect 4656 4467 4663 4513
rect 4756 4503 4763 4532
rect 4756 4496 4803 4503
rect 4613 4447 4627 4453
rect 4607 4440 4627 4447
rect 4607 4436 4623 4440
rect 4607 4433 4620 4436
rect 4576 4416 4603 4423
rect 4576 4336 4583 4393
rect 4596 4367 4603 4416
rect 4396 4006 4403 4092
rect 4296 3707 4303 3772
rect 4316 3627 4323 3653
rect 4216 3596 4233 3603
rect 4116 3347 4123 3553
rect 4156 3516 4163 3553
rect 4236 3547 4243 3593
rect 4193 3520 4207 3532
rect 4196 3516 4203 3520
rect 4176 3447 4183 3483
rect 4076 3320 4103 3323
rect 4073 3316 4103 3320
rect 4073 3307 4087 3316
rect 4153 3300 4167 3313
rect 4176 3307 4183 3333
rect 4156 3296 4163 3300
rect 4016 3136 4043 3143
rect 4016 3027 4023 3136
rect 3993 3007 4007 3013
rect 3976 2847 3983 2963
rect 4016 2927 4023 3013
rect 4036 3007 4043 3113
rect 4053 3000 4067 3013
rect 4056 2996 4063 3000
rect 4096 2996 4103 3213
rect 4136 3127 4143 3263
rect 4176 3187 4183 3253
rect 4127 3013 4133 3027
rect 4116 2960 4123 2963
rect 4113 2947 4127 2960
rect 4133 2947 4147 2952
rect 4156 2947 4163 3153
rect 4196 3107 4203 3413
rect 4216 3343 4223 3433
rect 4236 3387 4243 3533
rect 4296 3516 4303 3553
rect 4336 3527 4343 3813
rect 4356 3707 4363 3853
rect 4416 3847 4423 4073
rect 4436 4047 4443 4112
rect 4516 4067 4523 4172
rect 4436 3843 4443 3993
rect 4476 3947 4483 4003
rect 4536 3847 4543 4293
rect 4556 4267 4563 4303
rect 4596 4287 4603 4303
rect 4556 4207 4563 4253
rect 4596 4247 4603 4273
rect 4576 4036 4583 4173
rect 4616 4047 4623 4293
rect 4636 4247 4643 4453
rect 4656 4307 4663 4353
rect 4756 4303 4763 4473
rect 4676 4207 4683 4303
rect 4736 4296 4763 4303
rect 4596 4000 4603 4003
rect 4593 3987 4607 4000
rect 4436 3840 4463 3843
rect 4436 3836 4467 3840
rect 4413 3820 4427 3833
rect 4453 3827 4467 3836
rect 4416 3816 4423 3820
rect 4316 3447 4323 3483
rect 4356 3347 4363 3633
rect 4376 3527 4383 3673
rect 4436 3627 4443 3783
rect 4476 3747 4483 3833
rect 4536 3816 4543 3833
rect 4576 3816 4583 3973
rect 4616 3927 4623 3993
rect 4636 3987 4643 4133
rect 4656 4048 4663 4113
rect 4676 4036 4683 4093
rect 4696 4087 4703 4233
rect 4716 4187 4723 4253
rect 4736 4067 4743 4213
rect 4713 4040 4727 4053
rect 4756 4047 4763 4153
rect 4716 4036 4723 4040
rect 4456 3347 4463 3513
rect 4476 3367 4483 3693
rect 4516 3607 4523 3783
rect 4536 3647 4543 3753
rect 4556 3747 4563 3783
rect 4567 3736 4583 3743
rect 4540 3523 4553 3527
rect 4536 3516 4553 3523
rect 4540 3513 4553 3516
rect 4576 3486 4583 3736
rect 4616 3687 4623 3773
rect 4636 3607 4643 3833
rect 4656 3827 4663 3993
rect 4696 3887 4703 4003
rect 4673 3820 4687 3833
rect 4676 3816 4683 3820
rect 4716 3816 4723 3853
rect 4696 3747 4703 3783
rect 4736 3707 4743 3783
rect 4776 3707 4783 4453
rect 4796 4347 4803 4496
rect 4836 4467 4843 4633
rect 4856 4526 4863 4813
rect 4876 4747 4883 4773
rect 4876 4567 4883 4653
rect 4896 4583 4903 4823
rect 4916 4767 4923 4813
rect 4936 4707 4943 5013
rect 4976 4856 4983 4893
rect 5016 4856 5023 4913
rect 5036 4887 5043 5093
rect 5073 5080 5087 5093
rect 5113 5080 5127 5093
rect 5076 5076 5083 5080
rect 5116 5076 5123 5080
rect 5236 5076 5243 5343
rect 5096 5040 5103 5043
rect 5093 5027 5107 5040
rect 5136 4987 5143 5043
rect 5176 5043 5183 5072
rect 5167 5036 5183 5043
rect 5156 4963 5163 5032
rect 5196 4967 5203 5033
rect 5127 4956 5163 4963
rect 5076 4827 5083 4953
rect 5156 4856 5163 4913
rect 5236 4867 5243 5013
rect 5256 5007 5263 5043
rect 5296 5046 5303 5153
rect 5316 5087 5323 5374
rect 5700 5383 5713 5387
rect 5696 5376 5713 5383
rect 5700 5373 5713 5376
rect 5376 5340 5383 5343
rect 5373 5327 5387 5340
rect 5496 5340 5503 5343
rect 5536 5340 5543 5343
rect 5413 5327 5427 5332
rect 5493 5327 5507 5340
rect 5533 5327 5547 5340
rect 5336 5076 5343 5293
rect 5273 5027 5287 5033
rect 5436 5007 5443 5113
rect 5556 5076 5563 5133
rect 5456 4987 5463 5074
rect 5596 5067 5603 5373
rect 5700 5368 5706 5373
rect 5616 5087 5623 5333
rect 5636 5307 5643 5343
rect 5676 5287 5683 5343
rect 5736 5267 5743 5374
rect 5796 5340 5803 5343
rect 5753 5323 5767 5333
rect 5793 5327 5807 5340
rect 5753 5320 5783 5323
rect 5756 5316 5783 5320
rect 5696 5147 5703 5253
rect 5647 5083 5660 5087
rect 5647 5076 5663 5083
rect 5696 5076 5703 5133
rect 5647 5073 5660 5076
rect 5600 5046 5613 5047
rect 4956 4607 4963 4813
rect 4996 4747 5003 4823
rect 5036 4820 5043 4823
rect 5033 4807 5047 4820
rect 5067 4816 5083 4827
rect 5067 4813 5080 4816
rect 4896 4576 4923 4583
rect 4916 4556 4923 4576
rect 4936 4467 4943 4523
rect 4976 4487 4983 4513
rect 4836 4367 4843 4413
rect 4856 4336 4863 4373
rect 4796 4127 4803 4293
rect 4836 4067 4843 4303
rect 4896 4287 4903 4373
rect 4996 4363 5003 4733
rect 5056 4556 5063 4773
rect 5076 4763 5083 4793
rect 5096 4787 5103 4813
rect 5136 4783 5143 4812
rect 5116 4776 5143 4783
rect 5116 4763 5123 4776
rect 5076 4756 5123 4763
rect 5156 4683 5163 4753
rect 5176 4747 5183 4823
rect 5156 4676 5183 4683
rect 5096 4568 5103 4593
rect 5136 4527 5143 4593
rect 5176 4568 5183 4676
rect 5196 4607 5203 4813
rect 5216 4747 5223 4854
rect 5296 4867 5303 4913
rect 5316 4868 5323 4953
rect 5496 4927 5503 5043
rect 5607 5033 5613 5046
rect 5476 4867 5483 4893
rect 5316 4827 5323 4854
rect 5516 4856 5523 4893
rect 5556 4856 5563 4893
rect 5276 4807 5283 4823
rect 5347 4823 5360 4827
rect 5347 4816 5363 4823
rect 5347 4813 5360 4816
rect 5393 4807 5407 4812
rect 5276 4796 5293 4807
rect 5280 4793 5293 4796
rect 5316 4568 5323 4593
rect 5016 4387 5023 4513
rect 5036 4367 5043 4523
rect 5196 4487 5203 4523
rect 5236 4427 5243 4523
rect 5276 4467 5283 4553
rect 5376 4467 5383 4523
rect 5396 4487 5403 4513
rect 5056 4367 5063 4393
rect 4976 4356 5003 4363
rect 4976 4336 4983 4356
rect 5013 4340 5027 4352
rect 5016 4336 5023 4340
rect 4956 4300 4963 4303
rect 4953 4287 4967 4300
rect 4836 4036 4843 4053
rect 4873 4040 4887 4053
rect 4876 4036 4883 4040
rect 4856 3947 4863 4003
rect 4916 3987 4923 4253
rect 4996 4147 5003 4303
rect 5056 4107 5063 4353
rect 5116 4336 5123 4393
rect 5236 4363 5243 4413
rect 5216 4356 5243 4363
rect 5216 4336 5223 4356
rect 5316 4347 5323 4373
rect 5256 4336 5303 4343
rect 4987 4073 4993 4087
rect 5013 4040 5027 4053
rect 5016 4036 5023 4040
rect 4796 3907 4803 3933
rect 4876 3827 4883 3873
rect 4816 3647 4823 3783
rect 4636 3516 4643 3553
rect 4676 3528 4683 3593
rect 4856 3587 4863 3783
rect 4876 3727 4883 3773
rect 4896 3767 4903 3853
rect 4956 3828 4963 4003
rect 4996 3816 5003 3853
rect 5016 3827 5023 3933
rect 4973 3767 4987 3772
rect 4796 3516 4803 3573
rect 4556 3427 4563 3473
rect 4656 3480 4663 3483
rect 4653 3467 4667 3480
rect 4216 3336 4243 3343
rect 4236 3296 4243 3336
rect 4467 3336 4483 3343
rect 4176 3007 4183 3053
rect 4216 3043 4223 3253
rect 4256 3227 4263 3263
rect 4267 3216 4283 3223
rect 4256 3127 4263 3173
rect 4196 3040 4223 3043
rect 4193 3036 4223 3040
rect 4193 3027 4207 3036
rect 4227 3016 4263 3023
rect 4256 2996 4263 3016
rect 4276 3007 4283 3216
rect 3696 2740 3703 2743
rect 3596 2476 3603 2613
rect 2816 1956 2823 1993
rect 2876 1967 2883 2073
rect 2860 1963 2873 1967
rect 2856 1956 2873 1963
rect 2860 1953 2873 1956
rect 2836 1887 2843 1923
rect 2796 1748 2803 1833
rect 2836 1736 2843 1793
rect 2816 1667 2823 1703
rect 2796 1436 2803 1513
rect 2833 1440 2847 1453
rect 2836 1436 2843 1440
rect 2756 1347 2763 1392
rect 2736 1316 2763 1323
rect 2636 1216 2683 1223
rect 2713 1220 2727 1233
rect 2756 1227 2763 1316
rect 2876 1247 2883 1693
rect 2896 1647 2903 2113
rect 2976 2087 2983 2333
rect 3033 2260 3047 2273
rect 3036 2256 3043 2260
rect 3076 2167 3083 2273
rect 3096 2268 3103 2373
rect 3096 2123 3103 2254
rect 3156 2187 3163 2223
rect 3236 2207 3243 2393
rect 3296 2288 3303 2432
rect 3336 2303 3343 2443
rect 3476 2347 3483 2443
rect 3336 2296 3363 2303
rect 3333 2260 3347 2273
rect 3356 2267 3363 2296
rect 3336 2256 3343 2260
rect 3496 2267 3503 2413
rect 3556 2367 3563 2473
rect 3676 2347 3683 2733
rect 3693 2727 3707 2740
rect 3696 2647 3703 2713
rect 3796 2707 3803 2776
rect 3916 2746 3923 2793
rect 3936 2783 3943 2833
rect 3936 2776 3963 2783
rect 3996 2776 4003 2813
rect 3716 2447 3723 2513
rect 3787 2476 3803 2483
rect 3096 2116 3123 2123
rect 3076 1956 3083 2113
rect 3116 1967 3123 2116
rect 2916 1747 2923 1933
rect 2936 1887 2943 1913
rect 3016 1923 3023 1954
rect 2996 1916 3023 1923
rect 2936 1547 2943 1703
rect 2956 1527 2963 1793
rect 2976 1667 2983 1773
rect 2996 1607 3003 1916
rect 3136 1923 3143 2093
rect 3156 2027 3163 2173
rect 3196 1968 3203 2191
rect 3276 2167 3283 2223
rect 3316 2220 3323 2223
rect 3313 2207 3327 2220
rect 3276 2007 3283 2153
rect 3356 2107 3363 2213
rect 3376 2187 3383 2253
rect 3407 2223 3420 2227
rect 3407 2216 3423 2223
rect 3407 2213 3420 2216
rect 3336 2027 3343 2073
rect 3396 2047 3403 2153
rect 3456 2087 3463 2223
rect 3576 2220 3583 2223
rect 3573 2207 3587 2220
rect 3336 1956 3343 2013
rect 3456 1956 3463 1993
rect 3496 1956 3503 2013
rect 3596 1956 3603 2013
rect 3636 1956 3643 2333
rect 3696 2268 3703 2353
rect 3736 2167 3743 2443
rect 3796 2287 3803 2476
rect 3816 2347 3823 2573
rect 3836 2487 3843 2732
rect 3976 2707 3983 2743
rect 4016 2740 4023 2743
rect 4013 2727 4027 2740
rect 4056 2607 4063 2633
rect 3856 2476 3863 2513
rect 3896 2476 3903 2533
rect 3820 2283 3833 2287
rect 3816 2273 3833 2283
rect 3756 2207 3763 2273
rect 3816 2256 3823 2273
rect 3856 2267 3863 2413
rect 3876 2407 3883 2443
rect 4056 2407 4063 2473
rect 3836 2220 3843 2223
rect 3833 2207 3847 2220
rect 3736 2127 3743 2153
rect 3756 2027 3763 2193
rect 3976 2187 3983 2273
rect 3996 2207 4003 2333
rect 4076 2263 4083 2773
rect 4096 2667 4103 2873
rect 4116 2787 4123 2813
rect 4196 2807 4203 2833
rect 4136 2707 4143 2743
rect 4176 2736 4203 2743
rect 4176 2367 4183 2713
rect 4196 2607 4203 2736
rect 4216 2707 4223 2933
rect 4236 2923 4243 2963
rect 4236 2916 4263 2923
rect 4236 2783 4243 2893
rect 4256 2847 4263 2916
rect 4296 2907 4303 3253
rect 4316 3247 4323 3333
rect 4433 3307 4447 3313
rect 4476 3307 4483 3336
rect 4500 3323 4513 3327
rect 4496 3313 4513 3323
rect 4556 3323 4563 3413
rect 4536 3316 4563 3323
rect 4496 3296 4503 3313
rect 4536 3296 4543 3316
rect 4576 3307 4583 3353
rect 4376 3260 4383 3263
rect 4373 3247 4387 3260
rect 4416 3243 4423 3263
rect 4396 3240 4423 3243
rect 4396 3236 4427 3240
rect 4316 3008 4323 3233
rect 4396 3127 4403 3236
rect 4413 3227 4427 3236
rect 4456 3207 4463 3273
rect 4416 3047 4423 3153
rect 4416 2996 4423 3033
rect 4356 2960 4363 2963
rect 4353 2947 4367 2960
rect 4456 2947 4463 3193
rect 4476 3008 4483 3253
rect 4596 3266 4603 3333
rect 4656 3296 4663 3413
rect 4716 3347 4723 3514
rect 4553 3247 4567 3252
rect 4576 3207 4583 3253
rect 4736 3263 4743 3393
rect 4756 3307 4763 3453
rect 4776 3427 4783 3483
rect 4856 3303 4863 3573
rect 4916 3516 4923 3573
rect 4896 3407 4903 3483
rect 4956 3447 4963 3693
rect 4976 3527 4983 3613
rect 5036 3567 5043 3953
rect 5056 3907 5063 4034
rect 5076 3887 5083 4073
rect 5096 4067 5103 4303
rect 5236 4267 5243 4303
rect 5116 4036 5123 4093
rect 5176 3967 5183 4003
rect 5096 3867 5103 3893
rect 5136 3816 5143 3853
rect 5056 3627 5063 3773
rect 5176 3786 5183 3913
rect 5196 3827 5203 3933
rect 5216 3847 5223 4093
rect 5296 4063 5303 4336
rect 5356 4336 5363 4413
rect 5416 4347 5423 4713
rect 5436 4607 5443 4813
rect 5456 4587 5463 4853
rect 5596 4826 5603 4973
rect 5616 4867 5623 4993
rect 5636 4987 5643 5013
rect 5676 4967 5683 5043
rect 5716 4907 5723 5043
rect 5716 4863 5723 4893
rect 5696 4856 5723 4863
rect 5516 4556 5523 4613
rect 5456 4367 5463 4523
rect 5376 4267 5383 4303
rect 5276 4056 5303 4063
rect 5276 4036 5283 4056
rect 5316 4048 5323 4233
rect 5236 3816 5243 3933
rect 5256 3847 5263 4003
rect 5296 4000 5303 4003
rect 5293 3987 5307 4000
rect 5356 3987 5363 4153
rect 5376 4003 5383 4253
rect 5436 4247 5443 4334
rect 5516 4336 5523 4413
rect 5556 4336 5563 4793
rect 5636 4747 5643 4823
rect 5596 4568 5603 4673
rect 5636 4556 5643 4613
rect 5456 4167 5463 4332
rect 5456 4107 5463 4153
rect 5376 3996 5403 4003
rect 5276 3828 5283 3893
rect 4996 3516 5003 3553
rect 4973 3467 4987 3472
rect 5096 3467 5103 3553
rect 5136 3516 5143 3613
rect 5156 3547 5163 3773
rect 5200 3487 5206 3492
rect 5200 3483 5213 3487
rect 5156 3480 5163 3483
rect 4893 3307 4907 3313
rect 4856 3296 4883 3303
rect 4676 3260 4683 3263
rect 4673 3247 4687 3260
rect 4716 3256 4743 3263
rect 4496 2996 4503 3073
rect 4656 2996 4663 3033
rect 4696 2996 4703 3113
rect 4716 3087 4723 3256
rect 4736 3127 4743 3233
rect 4756 3063 4763 3233
rect 4776 3227 4783 3263
rect 4813 3247 4827 3252
rect 4736 3056 4763 3063
rect 4736 2966 4743 3056
rect 4813 3000 4827 3013
rect 4853 3007 4867 3013
rect 4876 3007 4883 3296
rect 4933 3300 4947 3313
rect 4936 3296 4943 3300
rect 5056 3296 5063 3393
rect 5116 3327 5123 3473
rect 5153 3467 5167 3480
rect 5196 3476 5213 3483
rect 5200 3473 5213 3476
rect 5136 3307 5143 3433
rect 5236 3367 5243 3753
rect 5256 3567 5263 3783
rect 5316 3767 5323 3853
rect 5356 3816 5363 3913
rect 5396 3816 5403 3996
rect 5476 4003 5483 4173
rect 5536 4087 5543 4303
rect 5576 4036 5583 4153
rect 5596 4047 5603 4453
rect 5656 4387 5663 4523
rect 5616 4347 5623 4373
rect 5676 4363 5683 4513
rect 5696 4507 5703 4573
rect 5716 4567 5723 4813
rect 5736 4687 5743 4853
rect 5756 4727 5763 5293
rect 5776 4587 5783 5316
rect 5796 4827 5803 5273
rect 5766 4573 5767 4580
rect 5753 4560 5767 4573
rect 5756 4556 5763 4560
rect 5796 4556 5803 4653
rect 5656 4356 5683 4363
rect 5656 4336 5663 4356
rect 5696 4336 5703 4453
rect 5636 4267 5643 4303
rect 5616 4048 5623 4073
rect 5676 4063 5683 4292
rect 5736 4187 5743 4523
rect 5676 4056 5703 4063
rect 5696 4036 5703 4056
rect 5456 3996 5483 4003
rect 5416 3847 5423 3992
rect 5336 3727 5343 3773
rect 5416 3780 5423 3783
rect 5413 3767 5427 3780
rect 5256 3527 5263 3553
rect 5376 3486 5383 3533
rect 5396 3527 5403 3573
rect 5416 3547 5423 3753
rect 5456 3587 5463 3996
rect 5496 3816 5503 3913
rect 5516 3887 5523 4003
rect 5516 3547 5523 3783
rect 5556 3767 5563 3992
rect 5616 3987 5623 4034
rect 5576 3747 5583 3973
rect 5636 3967 5643 3993
rect 5756 4003 5763 4493
rect 5776 4447 5783 4523
rect 5716 3967 5723 4003
rect 5736 3996 5763 4003
rect 5633 3863 5647 3873
rect 5616 3860 5647 3863
rect 5616 3856 5643 3860
rect 5616 3843 5623 3856
rect 5596 3840 5623 3843
rect 5593 3836 5623 3840
rect 5593 3827 5607 3836
rect 5633 3820 5647 3833
rect 5636 3816 5643 3820
rect 5736 3827 5743 3996
rect 5776 3907 5783 4213
rect 5796 3887 5803 4493
rect 5816 3847 5823 4433
rect 5433 3528 5447 3533
rect 5276 3327 5283 3483
rect 5396 3447 5403 3473
rect 5287 3316 5303 3323
rect 5016 3266 5023 3293
rect 4896 3187 4903 3253
rect 4956 3227 4963 3263
rect 5116 3187 5123 3263
rect 5156 3266 5163 3313
rect 4816 2996 4823 3000
rect 4476 2927 4483 2953
rect 4556 2847 4563 2963
rect 4796 2960 4803 2963
rect 4793 2947 4807 2960
rect 4787 2916 4813 2923
rect 4236 2776 4253 2783
rect 4196 2307 4203 2513
rect 4236 2476 4243 2533
rect 4376 2527 4383 2813
rect 4396 2767 4403 2793
rect 4433 2780 4447 2793
rect 4436 2776 4443 2780
rect 4516 2746 4523 2833
rect 4573 2780 4587 2793
rect 4576 2776 4583 2780
rect 4616 2776 4623 2813
rect 4713 2780 4727 2793
rect 4716 2776 4723 2780
rect 4796 2787 4803 2813
rect 4456 2740 4463 2743
rect 4453 2727 4467 2740
rect 4596 2740 4603 2743
rect 4696 2740 4703 2743
rect 4593 2727 4607 2740
rect 4693 2727 4707 2740
rect 4256 2347 4263 2432
rect 4416 2407 4423 2473
rect 4536 2447 4543 2533
rect 4576 2476 4583 2513
rect 4616 2476 4623 2593
rect 4756 2476 4763 2533
rect 4476 2367 4483 2443
rect 4076 2256 4103 2263
rect 3673 1960 3687 1973
rect 3676 1956 3683 1960
rect 3096 1907 3103 1923
rect 3116 1916 3143 1923
rect 3016 1627 3023 1793
rect 2953 1440 2967 1453
rect 2996 1447 3003 1473
rect 2956 1436 2963 1440
rect 2936 1383 2943 1403
rect 2936 1376 2963 1383
rect 2716 1216 2723 1220
rect 2756 1216 2773 1227
rect 2676 1187 2683 1216
rect 2760 1213 2773 1216
rect 2616 1167 2623 1183
rect 2436 647 2443 733
rect 2456 727 2463 953
rect 2496 916 2503 953
rect 2536 916 2543 1093
rect 2616 1003 2623 1153
rect 2736 1107 2743 1183
rect 2796 1183 2803 1233
rect 2896 1216 2903 1293
rect 2796 1176 2843 1183
rect 2596 996 2623 1003
rect 2596 887 2603 996
rect 2616 927 2623 953
rect 2516 880 2523 883
rect 2513 867 2527 880
rect 2636 880 2643 883
rect 2633 867 2647 880
rect 2687 883 2700 887
rect 2687 873 2703 883
rect 2553 700 2567 713
rect 2556 696 2563 700
rect 2476 587 2483 663
rect 2036 366 2043 433
rect 2056 407 2063 433
rect 2076 427 2083 513
rect 2256 396 2263 573
rect 2276 407 2283 433
rect 2056 287 2063 353
rect 2116 263 2123 363
rect 2176 347 2183 394
rect 2393 400 2407 413
rect 2416 403 2423 513
rect 2436 467 2443 493
rect 2476 487 2483 513
rect 2516 487 2523 652
rect 2396 396 2403 400
rect 2416 396 2443 403
rect 2096 256 2123 263
rect 2096 146 2103 256
rect 2196 227 2203 353
rect 2236 347 2243 363
rect 2227 336 2243 347
rect 2227 333 2240 336
rect 2276 267 2283 353
rect 2296 327 2303 394
rect 2327 363 2340 367
rect 2327 356 2343 363
rect 2327 353 2340 356
rect 2536 287 2543 433
rect 2296 243 2303 273
rect 2276 240 2303 243
rect 2273 236 2303 240
rect 2273 227 2287 236
rect 2196 188 2203 213
rect 2293 180 2307 193
rect 2296 176 2303 180
rect 1916 27 1923 143
rect 2216 107 2223 173
rect 2416 146 2423 213
rect 2556 167 2563 593
rect 2616 507 2623 793
rect 2636 547 2643 853
rect 2696 787 2703 873
rect 2676 660 2683 663
rect 2673 647 2687 660
rect 2736 607 2743 663
rect 2616 176 2623 213
rect 2656 207 2663 493
rect 2676 366 2683 413
rect 2716 396 2723 573
rect 2736 447 2743 553
rect 2753 400 2767 413
rect 2776 407 2783 1173
rect 2796 923 2803 1153
rect 2936 987 2943 1353
rect 2956 1327 2963 1376
rect 2996 1287 3003 1393
rect 3016 1263 3023 1493
rect 3036 1367 3043 1653
rect 3076 1607 3083 1873
rect 3096 1847 3103 1893
rect 3116 1807 3123 1916
rect 3176 1920 3183 1923
rect 3216 1920 3223 1923
rect 3156 1827 3163 1913
rect 3173 1907 3187 1920
rect 3213 1907 3227 1920
rect 3276 1887 3283 1953
rect 3056 1436 3063 1493
rect 3116 1443 3123 1692
rect 3116 1436 3143 1443
rect 3056 1327 3063 1373
rect 3096 1347 3103 1403
rect 3236 1327 3243 1813
rect 3316 1787 3323 1923
rect 3416 1907 3423 1954
rect 3536 1927 3543 1954
rect 3356 1707 3363 1853
rect 3456 1703 3463 1793
rect 3476 1747 3483 1923
rect 3576 1807 3583 1923
rect 3616 1867 3623 1923
rect 3776 1827 3783 1954
rect 3456 1696 3472 1703
rect 3256 1323 3263 1593
rect 3316 1367 3323 1403
rect 3256 1316 3283 1323
rect 3016 1256 3043 1263
rect 2973 1220 2987 1233
rect 3013 1220 3027 1233
rect 3036 1227 3043 1256
rect 2976 1216 2983 1220
rect 3016 1216 3023 1220
rect 3053 1220 3067 1233
rect 3056 1216 3063 1220
rect 3116 1186 3123 1293
rect 2796 916 2813 923
rect 2876 916 2883 953
rect 2927 883 2940 887
rect 2927 876 2943 883
rect 2927 873 2940 876
rect 2796 407 2803 793
rect 2996 787 3003 1093
rect 2836 696 2843 733
rect 2876 708 2883 773
rect 3016 767 3023 1073
rect 3036 923 3043 1173
rect 3136 1147 3143 1233
rect 3236 1107 3243 1183
rect 3276 1127 3283 1316
rect 3036 916 3053 923
rect 3116 916 3123 1013
rect 2976 696 2983 753
rect 2856 527 2863 663
rect 2916 647 2923 693
rect 2756 396 2763 400
rect 2873 400 2887 413
rect 2916 407 2923 533
rect 2876 396 2883 400
rect 2653 180 2667 193
rect 2656 176 2663 180
rect 2276 107 2283 143
rect 2636 107 2643 143
rect 2676 67 2683 143
rect 2716 67 2723 313
rect 2736 267 2743 363
rect 2796 327 2803 372
rect 2936 367 2943 413
rect 2976 396 2983 453
rect 3016 396 3023 473
rect 3036 467 3043 653
rect 3056 627 3063 773
rect 3056 447 3063 613
rect 2856 287 2863 363
rect 3036 360 3043 363
rect 3033 347 3047 360
rect 3076 307 3083 793
rect 3156 703 3163 1053
rect 3176 807 3183 1073
rect 3236 1027 3243 1093
rect 3216 916 3223 973
rect 3236 827 3243 883
rect 3196 703 3203 813
rect 3136 696 3163 703
rect 3176 696 3203 703
rect 3236 696 3243 773
rect 3276 703 3283 953
rect 3296 947 3303 1233
rect 3316 1227 3323 1273
rect 3356 1247 3363 1633
rect 3416 1367 3423 1403
rect 3476 1403 3483 1692
rect 3536 1647 3543 1703
rect 3596 1700 3603 1703
rect 3593 1687 3607 1700
rect 3696 1687 3703 1813
rect 3776 1736 3783 1773
rect 3796 1767 3803 2113
rect 3996 1963 4003 2073
rect 4096 1987 4103 2256
rect 4153 2260 4167 2273
rect 4156 2256 4163 2260
rect 4236 2267 4243 2293
rect 4116 2226 4123 2253
rect 4256 2227 4263 2253
rect 4176 2220 4183 2223
rect 4173 2207 4187 2220
rect 3976 1956 4003 1963
rect 3856 1827 3863 1912
rect 3516 1436 3523 1493
rect 3596 1443 3603 1673
rect 3716 1483 3723 1734
rect 3716 1476 3733 1483
rect 3596 1436 3623 1443
rect 3673 1440 3687 1453
rect 3676 1436 3683 1440
rect 3716 1407 3723 1452
rect 3476 1396 3503 1403
rect 3456 1287 3463 1393
rect 3347 1236 3363 1247
rect 3456 1216 3463 1273
rect 3496 1228 3503 1396
rect 3536 1327 3543 1403
rect 3316 916 3323 973
rect 3336 747 3343 883
rect 3376 827 3383 873
rect 3396 747 3403 1113
rect 3416 987 3423 1213
rect 3476 947 3483 1183
rect 3536 1087 3543 1313
rect 3593 1220 3607 1233
rect 3736 1243 3743 1473
rect 3836 1367 3843 1753
rect 3876 1736 3883 1773
rect 3936 1706 3943 1733
rect 3996 1700 4003 1703
rect 3896 1647 3903 1692
rect 3993 1687 4007 1700
rect 4036 1647 4043 1703
rect 3856 1387 3863 1513
rect 4056 1467 4063 1693
rect 4076 1687 4083 1793
rect 4096 1747 4103 1813
rect 4136 1807 4143 1973
rect 4193 1960 4207 1973
rect 4196 1956 4203 1960
rect 4256 1847 4263 2192
rect 4336 2047 4343 2223
rect 4376 2087 4383 2353
rect 4416 2256 4423 2333
rect 4476 2267 4483 2332
rect 4496 2287 4503 2432
rect 4596 2407 4603 2443
rect 4676 2367 4683 2474
rect 4796 2447 4803 2513
rect 4276 1956 4303 1963
rect 4276 1827 4283 1956
rect 4276 1787 4283 1813
rect 4173 1747 4187 1753
rect 4293 1740 4307 1753
rect 4316 1747 4323 1833
rect 4296 1736 4303 1740
rect 4116 1683 4123 1703
rect 4116 1676 4143 1683
rect 3936 1400 3943 1403
rect 3896 1347 3903 1392
rect 3933 1387 3947 1400
rect 3736 1236 3763 1243
rect 3633 1227 3647 1233
rect 3756 1228 3763 1236
rect 3596 1216 3603 1220
rect 4076 1223 4083 1363
rect 4136 1247 4143 1676
rect 4156 1607 4163 1703
rect 4196 1687 4203 1734
rect 4356 1743 4363 1883
rect 4336 1736 4363 1743
rect 4396 1736 4403 1793
rect 4416 1767 4423 2033
rect 4436 2027 4443 2223
rect 4496 2047 4503 2273
rect 4553 2260 4567 2273
rect 4556 2256 4563 2260
rect 4596 1983 4603 2013
rect 4616 2007 4623 2273
rect 4653 2260 4667 2273
rect 4696 2267 4703 2413
rect 4656 2256 4663 2260
rect 4596 1976 4623 1983
rect 4616 1956 4623 1976
rect 4656 1956 4663 1993
rect 4676 1963 4683 2223
rect 4676 1956 4703 1963
rect 4496 1907 4503 1923
rect 4576 1920 4603 1923
rect 4573 1916 4603 1920
rect 4496 1896 4513 1907
rect 4500 1893 4513 1896
rect 4536 1827 4543 1913
rect 4573 1907 4587 1916
rect 4227 1703 4240 1707
rect 4227 1696 4243 1703
rect 4276 1700 4283 1703
rect 4227 1693 4240 1696
rect 4273 1687 4287 1700
rect 4176 1507 4183 1533
rect 4056 1216 4083 1223
rect 3576 1147 3583 1183
rect 3656 1167 3663 1214
rect 3687 1183 3700 1187
rect 3687 1176 3703 1183
rect 3687 1173 3700 1176
rect 3736 1087 3743 1183
rect 3796 1147 3803 1183
rect 3856 1180 3863 1183
rect 3853 1167 3867 1180
rect 3756 1107 3763 1133
rect 3480 883 3493 887
rect 3476 876 3493 883
rect 3480 873 3493 876
rect 3516 787 3523 933
rect 3553 920 3567 933
rect 3556 916 3563 920
rect 3636 886 3643 973
rect 3576 847 3583 883
rect 3687 836 3713 843
rect 3276 696 3303 703
rect 3096 587 3103 652
rect 3136 396 3143 493
rect 3176 463 3183 696
rect 3256 587 3263 663
rect 3196 527 3203 553
rect 3216 467 3223 493
rect 3176 456 3203 463
rect 3176 396 3183 433
rect 3196 407 3203 456
rect 3256 427 3263 453
rect 3296 427 3303 696
rect 3373 700 3387 713
rect 3416 707 3423 773
rect 3656 747 3663 813
rect 3756 807 3763 1093
rect 4056 1027 4063 1216
rect 4133 1220 4147 1233
rect 4136 1216 4143 1220
rect 4116 987 4123 1183
rect 3793 920 3807 933
rect 3796 916 3803 920
rect 3836 916 3843 973
rect 4176 947 4183 1493
rect 4236 1436 4243 1513
rect 4196 1367 4203 1403
rect 4256 1323 4263 1673
rect 4336 1467 4343 1736
rect 4416 1527 4423 1692
rect 4356 1436 4363 1513
rect 4276 1347 4283 1434
rect 4396 1406 4403 1453
rect 4256 1316 4283 1323
rect 4276 1207 4283 1316
rect 4336 1267 4343 1403
rect 4416 1327 4423 1513
rect 4436 1263 4443 1633
rect 4456 1607 4463 1753
rect 4476 1587 4483 1793
rect 4513 1743 4527 1753
rect 4496 1740 4527 1743
rect 4496 1736 4523 1740
rect 4496 1707 4503 1736
rect 4636 1743 4643 1923
rect 4696 1867 4703 1956
rect 4716 1923 4723 2013
rect 4816 1967 4823 2853
rect 4836 2827 4843 2963
rect 4876 2927 4883 2972
rect 4936 2927 4943 2963
rect 5016 2927 5023 3113
rect 5036 2967 5043 3033
rect 5116 3007 5123 3173
rect 4847 2783 4860 2787
rect 4847 2776 4863 2783
rect 4896 2776 4903 2853
rect 4847 2773 4860 2776
rect 4920 2743 4933 2747
rect 4916 2733 4933 2743
rect 4916 2487 4923 2733
rect 4956 2607 4963 2893
rect 4976 2787 4983 2913
rect 5136 2867 5143 3253
rect 5196 3207 5203 3263
rect 5296 3207 5303 3316
rect 5416 3323 5423 3483
rect 5516 3486 5523 3533
rect 5536 3527 5543 3633
rect 5596 3607 5603 3773
rect 5616 3727 5623 3783
rect 5656 3780 5663 3783
rect 5653 3767 5667 3780
rect 5596 3516 5603 3553
rect 5636 3527 5643 3733
rect 5696 3683 5703 3773
rect 5676 3676 5703 3683
rect 5676 3647 5683 3676
rect 5716 3663 5723 3813
rect 5736 3687 5743 3773
rect 5696 3656 5723 3663
rect 5676 3527 5683 3593
rect 5696 3528 5703 3656
rect 5716 3547 5723 3633
rect 5736 3516 5743 3593
rect 5756 3527 5763 3713
rect 5333 3300 5347 3313
rect 5396 3316 5423 3323
rect 5336 3296 5343 3300
rect 5216 2996 5223 3173
rect 5033 2807 5047 2813
rect 5056 2807 5063 2833
rect 5056 2746 5063 2793
rect 5076 2787 5083 2853
rect 5113 2807 5127 2813
rect 5113 2780 5127 2793
rect 5116 2776 5123 2780
rect 5176 2783 5183 2963
rect 5236 2927 5243 2993
rect 5256 2887 5263 3053
rect 5296 2996 5303 3033
rect 5356 3023 5363 3263
rect 5376 3127 5383 3233
rect 5336 3016 5363 3023
rect 5336 2996 5343 3016
rect 5396 2966 5403 3316
rect 5416 3296 5443 3303
rect 5416 3147 5423 3296
rect 5476 3207 5483 3263
rect 5476 3007 5483 3133
rect 5496 3067 5503 3473
rect 5516 3027 5523 3293
rect 5536 3247 5543 3433
rect 5636 3347 5643 3453
rect 5656 3323 5663 3513
rect 5636 3316 5663 3323
rect 5636 3296 5643 3316
rect 5676 3307 5683 3473
rect 5716 3343 5723 3483
rect 5696 3336 5723 3343
rect 5576 3147 5583 3263
rect 5616 3107 5623 3263
rect 5633 3227 5647 3233
rect 5476 2996 5493 3007
rect 5480 2993 5493 2996
rect 5536 2996 5563 3003
rect 5536 2967 5543 2996
rect 5316 2827 5323 2963
rect 5216 2787 5223 2813
rect 5176 2776 5203 2783
rect 4996 2476 5003 2613
rect 4836 2127 4843 2443
rect 4916 2387 4923 2473
rect 5036 2447 5043 2733
rect 5136 2740 5143 2743
rect 5133 2727 5147 2740
rect 5116 2476 5123 2553
rect 5176 2483 5183 2733
rect 5196 2667 5203 2776
rect 5253 2780 5267 2793
rect 5256 2776 5263 2780
rect 5236 2740 5243 2743
rect 5233 2727 5247 2740
rect 5216 2587 5223 2673
rect 5156 2476 5183 2483
rect 5156 2446 5163 2476
rect 5253 2480 5267 2493
rect 5256 2476 5263 2480
rect 5316 2476 5323 2593
rect 5336 2567 5343 2773
rect 5356 2746 5363 2913
rect 5416 2727 5423 2743
rect 5416 2716 5433 2727
rect 5420 2713 5433 2716
rect 5456 2583 5463 2873
rect 5516 2867 5523 2953
rect 5473 2787 5487 2793
rect 5516 2776 5523 2813
rect 5576 2787 5583 2893
rect 5616 2887 5623 2923
rect 5676 2907 5683 3233
rect 5696 2966 5703 3336
rect 5756 3323 5763 3473
rect 5713 3307 5727 3313
rect 5736 3316 5763 3323
rect 5736 3296 5743 3316
rect 5776 3307 5783 3783
rect 5596 2787 5603 2853
rect 5656 2776 5663 2813
rect 5716 2783 5723 3253
rect 5776 3207 5783 3233
rect 5756 2787 5763 2933
rect 5776 2807 5783 2963
rect 5796 2788 5803 3753
rect 5816 3707 5823 3773
rect 5816 2947 5823 3672
rect 5716 2776 5743 2783
rect 5476 2587 5483 2733
rect 5533 2727 5547 2732
rect 5436 2576 5463 2583
rect 5416 2446 5423 2473
rect 5436 2446 5443 2576
rect 4956 2227 4963 2273
rect 5013 2260 5027 2273
rect 5016 2256 5023 2260
rect 5056 2256 5063 2373
rect 5276 2327 5283 2443
rect 5536 2387 5543 2493
rect 4996 2187 5003 2223
rect 4876 1956 4883 2033
rect 4716 1916 4763 1923
rect 4616 1736 4643 1743
rect 4556 1687 4563 1703
rect 4456 1448 4463 1513
rect 4516 1507 4523 1593
rect 4556 1387 4563 1673
rect 4576 1447 4583 1693
rect 4596 1436 4603 1733
rect 4616 1667 4623 1736
rect 4676 1667 4683 1703
rect 4756 1527 4763 1893
rect 4796 1867 4803 1923
rect 4836 1736 4843 1793
rect 4873 1740 4887 1753
rect 4876 1736 4883 1740
rect 4776 1706 4783 1733
rect 4816 1587 4823 1703
rect 4856 1567 4863 1703
rect 4896 1487 4903 1693
rect 4916 1687 4923 1923
rect 4936 1747 4943 1953
rect 5016 1736 5023 1773
rect 4956 1667 4963 1703
rect 4636 1436 4683 1443
rect 4733 1440 4747 1453
rect 4736 1436 4743 1440
rect 4436 1256 4453 1263
rect 4296 1227 4303 1253
rect 4216 1127 4223 1183
rect 4216 1087 4223 1113
rect 4213 928 4227 933
rect 3927 923 3940 927
rect 3927 916 3943 923
rect 3976 916 4023 923
rect 3927 913 3940 916
rect 3816 863 3823 883
rect 3896 886 3903 913
rect 3873 863 3887 873
rect 3816 860 3887 863
rect 3816 856 3883 860
rect 3847 836 3873 843
rect 3516 707 3523 733
rect 3376 696 3383 700
rect 3416 656 3443 663
rect 3496 660 3503 663
rect 3116 360 3123 363
rect 3113 347 3127 360
rect 3156 267 3163 363
rect 2753 180 2767 193
rect 2796 188 2803 233
rect 2756 176 2763 180
rect 3196 187 3203 353
rect 3216 187 3223 393
rect 3296 327 3303 363
rect 3236 207 3243 293
rect 2916 146 2923 173
rect 2776 107 2783 143
rect 3136 107 3143 143
rect 3216 -24 3223 152
rect 3236 146 3243 193
rect 3336 146 3343 413
rect 3356 407 3363 553
rect 3416 547 3423 656
rect 3493 647 3507 660
rect 3376 423 3383 533
rect 3376 416 3403 423
rect 3396 396 3403 416
rect 3436 408 3443 613
rect 3516 527 3523 653
rect 3536 647 3543 713
rect 3556 587 3563 694
rect 3656 647 3663 733
rect 3676 647 3683 773
rect 3716 660 3723 663
rect 3713 647 3727 660
rect 3756 567 3763 663
rect 3796 660 3803 663
rect 3793 647 3807 660
rect 3796 587 3803 633
rect 3896 607 3903 793
rect 3956 787 3963 883
rect 4016 847 4023 916
rect 4167 923 4180 927
rect 4167 916 4183 923
rect 4167 913 4180 916
rect 4136 886 4143 913
rect 4276 907 4283 1113
rect 4296 987 4303 1173
rect 4336 947 4343 1183
rect 4436 1147 4443 1213
rect 4353 920 4367 933
rect 4356 916 4363 920
rect 4116 847 4123 873
rect 4273 883 4287 893
rect 4236 880 4287 883
rect 4236 876 4283 880
rect 3396 267 3403 293
rect 3416 247 3423 363
rect 3476 327 3483 413
rect 3513 400 3527 413
rect 3516 396 3523 400
rect 3676 396 3683 553
rect 3816 547 3823 593
rect 3916 547 3923 733
rect 4056 667 4063 694
rect 3956 660 3963 663
rect 3953 647 3967 660
rect 4016 607 4023 663
rect 4076 647 4083 733
rect 4196 666 4203 693
rect 4156 660 4163 663
rect 4153 647 4167 660
rect 3496 307 3503 353
rect 3476 227 3483 292
rect 3576 247 3583 394
rect 3616 307 3623 363
rect 3656 247 3663 363
rect 3436 147 3443 193
rect 3276 140 3283 143
rect 3273 127 3287 140
rect 3296 67 3303 93
rect 3336 27 3343 132
rect 3456 -24 3463 173
rect 3516 107 3523 143
rect 3556 87 3563 213
rect 3716 176 3723 493
rect 3756 396 3763 513
rect 3876 396 3883 453
rect 3916 396 3923 493
rect 3756 176 3763 213
rect 3776 207 3783 363
rect 3816 287 3823 394
rect 3856 327 3863 363
rect 3896 307 3903 363
rect 3876 176 3883 233
rect 3656 -24 3663 133
rect 3736 87 3743 143
rect 3756 -24 3763 113
rect 3776 87 3783 143
rect 3916 -17 3923 143
rect 3956 107 3963 533
rect 4053 400 4067 413
rect 4056 396 4063 400
rect 3996 327 4003 363
rect 4036 227 4043 363
rect 4096 247 4103 413
rect 4116 366 4123 453
rect 4136 427 4143 473
rect 4156 447 4163 533
rect 4216 507 4223 773
rect 4276 696 4283 733
rect 4356 667 4363 694
rect 4296 660 4303 663
rect 4293 647 4307 660
rect 4376 647 4383 1133
rect 4436 1067 4443 1093
rect 4416 727 4423 1013
rect 4436 787 4443 1053
rect 4456 1047 4463 1253
rect 4476 1227 4483 1273
rect 4556 1147 4563 1183
rect 4476 923 4483 1133
rect 4596 1107 4603 1373
rect 4516 987 4523 1053
rect 4616 1007 4623 1403
rect 4676 1403 4683 1436
rect 4676 1396 4723 1403
rect 4656 1228 4663 1393
rect 4636 1216 4653 1223
rect 4636 1167 4643 1216
rect 4696 1216 4703 1253
rect 4676 1180 4683 1183
rect 4673 1167 4687 1180
rect 4756 1107 4763 1313
rect 4816 1267 4823 1473
rect 4936 1406 4943 1433
rect 4896 1327 4903 1403
rect 5036 1327 5043 1692
rect 5056 1607 5063 1953
rect 5096 1926 5103 2293
rect 5256 2256 5263 2293
rect 5316 2267 5323 2353
rect 5196 2207 5203 2254
rect 5316 2226 5323 2253
rect 5436 2226 5443 2373
rect 5536 2256 5543 2293
rect 5556 2283 5563 2573
rect 5576 2407 5583 2733
rect 5596 2527 5603 2773
rect 5636 2740 5643 2743
rect 5676 2740 5683 2743
rect 5613 2727 5627 2733
rect 5633 2727 5647 2740
rect 5673 2727 5687 2740
rect 5716 2687 5723 2733
rect 5656 2476 5663 2513
rect 5636 2423 5643 2443
rect 5616 2416 5643 2423
rect 5616 2323 5623 2416
rect 5596 2316 5623 2323
rect 5556 2276 5583 2283
rect 5576 2256 5583 2276
rect 5596 2267 5603 2316
rect 5236 2220 5243 2223
rect 5233 2207 5247 2220
rect 5356 2220 5363 2223
rect 5353 2207 5367 2220
rect 5416 2007 5423 2223
rect 5456 2207 5463 2254
rect 5133 1960 5147 1973
rect 5136 1956 5143 1960
rect 5296 1956 5303 1993
rect 5420 1963 5433 1967
rect 5416 1956 5433 1963
rect 5420 1953 5433 1956
rect 5096 1667 5103 1912
rect 5136 1736 5143 1773
rect 5116 1487 5123 1703
rect 5127 1476 5143 1483
rect 5113 1440 5127 1452
rect 5136 1447 5143 1476
rect 5116 1436 5123 1440
rect 4656 967 4663 993
rect 4476 916 4503 923
rect 4436 696 4443 773
rect 4236 547 4243 573
rect 4156 396 4163 433
rect 4196 396 4203 493
rect 4236 396 4243 533
rect 4456 527 4463 733
rect 4336 396 4343 493
rect 3993 180 4007 193
rect 3996 176 4003 180
rect 4116 176 4123 293
rect 4176 187 4183 363
rect 4276 327 4283 394
rect 4236 176 4243 213
rect 3916 -24 3924 -17
rect 4036 -24 4043 143
rect 4156 -17 4163 143
rect 4276 -17 4283 143
rect 4316 127 4323 352
rect 4356 247 4363 363
rect 4376 176 4383 313
rect 4416 187 4423 363
rect 4476 227 4483 713
rect 4496 707 4503 916
rect 4516 863 4523 914
rect 4536 887 4543 953
rect 4696 927 4703 953
rect 4667 923 4680 927
rect 4667 914 4683 923
rect 4660 913 4683 914
rect 4716 916 4723 1033
rect 4756 928 4763 1093
rect 4676 887 4683 913
rect 4516 856 4543 863
rect 4536 696 4543 856
rect 4596 747 4603 883
rect 4656 720 4703 723
rect 4656 716 4707 720
rect 4656 696 4663 716
rect 4693 708 4707 716
rect 4496 208 4503 533
rect 4556 507 4563 663
rect 4573 647 4587 653
rect 4596 647 4603 693
rect 4636 660 4643 663
rect 4633 647 4647 660
rect 4596 607 4603 633
rect 4516 408 4523 433
rect 4533 400 4547 413
rect 4536 396 4543 400
rect 4596 396 4603 593
rect 4636 366 4643 633
rect 4656 366 4663 493
rect 4716 447 4723 773
rect 4796 747 4803 1013
rect 4816 967 4823 1183
rect 4836 916 4843 1053
rect 4876 1027 4883 1253
rect 4976 1228 4983 1313
rect 5016 1186 5023 1233
rect 5076 1216 5083 1273
rect 5096 1247 5103 1403
rect 5116 1227 5123 1313
rect 5156 1223 5163 1653
rect 5196 1467 5203 1953
rect 5216 1707 5223 1793
rect 5336 1748 5343 1953
rect 5396 1787 5403 1923
rect 5256 1567 5263 1703
rect 5256 1507 5263 1553
rect 5296 1547 5303 1703
rect 5396 1523 5403 1733
rect 5416 1543 5423 1893
rect 5456 1827 5463 2033
rect 5496 1968 5503 2193
rect 5616 1967 5623 2293
rect 5473 1907 5487 1912
rect 5636 1767 5643 2393
rect 5696 2367 5703 2593
rect 5736 2503 5743 2776
rect 5716 2500 5743 2503
rect 5713 2496 5743 2500
rect 5713 2487 5727 2496
rect 5776 2487 5783 2732
rect 5676 2256 5683 2313
rect 5716 2287 5723 2433
rect 5776 2407 5783 2433
rect 5736 2263 5743 2393
rect 5716 2256 5743 2263
rect 5696 2047 5703 2223
rect 5756 1983 5763 2353
rect 5747 1976 5763 1983
rect 5733 1960 5747 1973
rect 5736 1956 5743 1960
rect 5516 1667 5523 1703
rect 5576 1667 5583 1703
rect 5416 1536 5433 1543
rect 5376 1516 5403 1523
rect 5173 1443 5187 1453
rect 5233 1447 5247 1453
rect 5173 1440 5203 1443
rect 5176 1436 5203 1440
rect 5296 1436 5303 1473
rect 5216 1367 5223 1403
rect 5236 1267 5243 1393
rect 5256 1367 5263 1434
rect 5316 1327 5323 1403
rect 5376 1363 5383 1516
rect 5396 1447 5403 1493
rect 5436 1436 5443 1533
rect 5556 1436 5563 1473
rect 5676 1443 5683 1773
rect 5696 1527 5703 1813
rect 5776 1787 5783 2273
rect 5796 1748 5803 2713
rect 5816 2327 5823 2474
rect 5816 1667 5823 1973
rect 5656 1436 5683 1443
rect 5696 1436 5703 1473
rect 5376 1356 5403 1363
rect 5236 1228 5243 1253
rect 5136 1216 5163 1223
rect 4916 1180 4923 1183
rect 4913 1167 4927 1180
rect 4956 1147 4963 1183
rect 5100 1183 5113 1187
rect 5096 1176 5113 1183
rect 5100 1173 5113 1176
rect 5136 1167 5143 1216
rect 5296 1127 5303 1183
rect 5336 1087 5343 1183
rect 5096 916 5103 993
rect 5216 923 5223 993
rect 5216 916 5243 923
rect 4936 887 4943 914
rect 4856 807 4863 883
rect 4736 666 4743 733
rect 4976 727 4983 883
rect 5016 787 5023 872
rect 5116 827 5123 883
rect 4976 666 4983 713
rect 4756 627 4763 663
rect 4856 660 4863 663
rect 4916 660 4923 663
rect 4853 647 4867 660
rect 4913 647 4927 660
rect 5196 663 5203 914
rect 5376 887 5383 1333
rect 5396 1223 5403 1356
rect 5416 1247 5423 1392
rect 5456 1228 5463 1403
rect 5496 1327 5503 1393
rect 5516 1347 5523 1434
rect 5656 1406 5663 1436
rect 5576 1367 5583 1403
rect 5716 1400 5723 1403
rect 5656 1287 5663 1392
rect 5713 1387 5727 1400
rect 5756 1387 5763 1513
rect 5396 1216 5423 1223
rect 5516 1216 5523 1253
rect 5756 1216 5763 1373
rect 5796 1216 5803 1273
rect 5816 1227 5823 1653
rect 5396 967 5403 1173
rect 5456 916 5463 953
rect 5336 876 5363 883
rect 5276 836 5303 843
rect 5216 667 5223 793
rect 5276 767 5283 836
rect 5356 827 5363 876
rect 5536 886 5543 1183
rect 5676 1127 5683 1183
rect 5296 736 5303 813
rect 5176 656 5203 663
rect 4856 547 4863 633
rect 4736 396 4743 473
rect 4776 396 4783 533
rect 4916 403 4923 513
rect 4916 396 4943 403
rect 4996 396 5003 533
rect 4356 140 4363 143
rect 4353 127 4367 140
rect 4436 143 4443 193
rect 4536 176 4543 273
rect 4494 167 4508 173
rect 4436 136 4483 143
rect 4516 87 4523 143
rect 4556 140 4563 143
rect 4553 127 4567 140
rect 4596 127 4603 213
rect 4616 187 4623 233
rect 4636 176 4643 352
rect 4716 327 4723 363
rect 5076 363 5083 433
rect 5133 400 5147 413
rect 5136 396 5143 400
rect 5176 367 5183 656
rect 5376 663 5383 694
rect 5356 656 5383 663
rect 5216 408 5223 453
rect 5253 400 5267 413
rect 5256 396 5263 400
rect 5076 356 5103 363
rect 5356 366 5363 413
rect 5396 403 5403 693
rect 5416 663 5423 773
rect 5436 707 5443 883
rect 5676 883 5683 953
rect 5656 876 5683 883
rect 5716 883 5723 1073
rect 5776 967 5783 1183
rect 5716 876 5743 883
rect 5616 703 5623 843
rect 5596 696 5623 703
rect 5416 656 5463 663
rect 5396 396 5423 403
rect 5476 396 5483 633
rect 5596 423 5603 696
rect 5696 660 5703 663
rect 5693 647 5707 660
rect 5596 416 5623 423
rect 5616 396 5623 416
rect 5736 396 5743 753
rect 5816 647 5823 1173
rect 5376 363 5383 394
rect 5376 356 5403 363
rect 5096 247 5103 313
rect 4856 207 4863 233
rect 4673 180 4687 193
rect 4676 176 4683 180
rect 4656 140 4663 143
rect 4653 127 4667 140
rect 4736 87 4743 193
rect 4853 180 4867 193
rect 4856 176 4863 180
rect 4776 107 4783 143
rect 4836 87 4843 132
rect 4916 107 4923 193
rect 5096 176 5103 233
rect 5356 183 5363 352
rect 5347 176 5363 183
rect 5396 176 5403 356
rect 5456 207 5463 273
rect 5596 267 5603 363
rect 5636 327 5643 352
rect 5453 180 5467 193
rect 5456 176 5463 180
rect 5336 146 5343 173
rect 4780 86 4793 87
rect 4787 73 4793 86
rect 5036 47 5043 143
rect 5216 140 5223 143
rect 5213 127 5227 140
rect 5276 47 5283 143
rect 5376 107 5383 143
rect 5516 107 5523 193
rect 5556 187 5563 253
rect 5636 87 5643 143
rect 5676 127 5683 353
rect 5716 327 5723 363
rect 5796 327 5803 353
rect 5696 147 5703 233
rect 5716 187 5723 313
rect 5756 176 5763 313
rect 5816 87 5823 633
rect 5636 47 5643 73
rect 4156 -24 4164 -17
rect 4276 -24 4284 -17
<< m3contact >>
rect 893 5453 907 5467
rect 1313 5453 1327 5467
rect 1813 5453 1827 5467
rect 2033 5453 2047 5467
rect 2573 5453 2587 5467
rect 113 5413 127 5427
rect 253 5413 267 5427
rect 293 5413 307 5427
rect 412 5413 426 5427
rect 433 5413 447 5427
rect 613 5413 627 5427
rect 733 5413 747 5427
rect 173 5373 187 5387
rect 213 5374 227 5388
rect 292 5373 306 5387
rect 313 5373 327 5387
rect 373 5374 387 5388
rect 413 5373 427 5387
rect 73 5153 87 5167
rect 153 5313 167 5327
rect 93 5113 107 5127
rect 273 5332 287 5346
rect 233 5273 247 5287
rect 493 5374 507 5388
rect 353 5332 367 5346
rect 433 5332 447 5346
rect 393 5293 407 5307
rect 473 5293 487 5307
rect 653 5374 667 5388
rect 693 5374 707 5388
rect 773 5374 787 5388
rect 833 5374 847 5388
rect 1173 5433 1187 5447
rect 1033 5413 1047 5427
rect 993 5374 1007 5388
rect 1133 5374 1147 5388
rect 1493 5433 1507 5447
rect 1533 5433 1547 5447
rect 1733 5433 1747 5447
rect 1513 5413 1527 5427
rect 1253 5374 1267 5388
rect 1313 5374 1327 5388
rect 1353 5374 1367 5388
rect 1393 5374 1407 5388
rect 573 5313 587 5327
rect 593 5293 607 5307
rect 513 5253 527 5267
rect 273 5193 287 5207
rect 313 5193 327 5207
rect 253 5153 267 5167
rect 253 5093 267 5107
rect 113 5074 127 5088
rect 173 5074 187 5088
rect 233 5074 247 5088
rect 33 4893 47 4907
rect 73 4893 87 4907
rect 13 4613 27 4627
rect 133 5032 147 5046
rect 213 5032 227 5046
rect 153 4953 167 4967
rect 113 4913 127 4927
rect 93 4873 107 4887
rect 253 4913 267 4927
rect 173 4873 187 4887
rect 153 4853 167 4867
rect 53 4813 67 4827
rect 133 4812 147 4826
rect 93 4693 107 4707
rect 133 4613 147 4627
rect 53 4554 67 4568
rect 93 4554 107 4568
rect 273 4854 287 4868
rect 253 4812 267 4826
rect 293 4813 307 4827
rect 373 5153 387 5167
rect 333 5133 347 5147
rect 373 5093 387 5107
rect 413 5074 427 5088
rect 453 5074 467 5088
rect 513 5074 527 5088
rect 553 5074 567 5088
rect 353 4953 367 4967
rect 393 4933 407 4947
rect 433 4933 447 4947
rect 393 4893 407 4907
rect 353 4873 367 4887
rect 493 5032 507 5046
rect 533 4933 547 4947
rect 453 4893 467 4907
rect 432 4853 446 4867
rect 453 4853 467 4867
rect 493 4854 507 4868
rect 573 4893 587 4907
rect 573 4853 587 4867
rect 413 4812 427 4826
rect 313 4793 327 4807
rect 373 4793 387 4807
rect 253 4753 267 4767
rect 293 4753 307 4767
rect 213 4693 227 4707
rect 173 4573 187 4587
rect 53 4513 67 4527
rect 293 4713 307 4727
rect 553 4812 567 4826
rect 513 4773 527 4787
rect 793 5332 807 5346
rect 973 5332 987 5346
rect 1013 5332 1027 5346
rect 1113 5332 1127 5346
rect 1153 5332 1167 5346
rect 1273 5332 1287 5346
rect 753 5313 767 5327
rect 873 5313 887 5327
rect 693 5293 707 5307
rect 773 5273 787 5287
rect 633 5173 647 5187
rect 673 5173 687 5187
rect 813 5173 827 5187
rect 733 5133 747 5147
rect 773 5133 787 5147
rect 673 5013 687 5027
rect 653 4973 667 4987
rect 633 4933 647 4947
rect 853 5133 867 5147
rect 753 5033 767 5047
rect 933 5253 947 5267
rect 973 5113 987 5127
rect 973 5074 987 5088
rect 1013 5073 1027 5087
rect 1073 5074 1087 5088
rect 1293 5153 1307 5167
rect 1133 5074 1147 5088
rect 1173 5074 1187 5088
rect 1213 5074 1227 5088
rect 1273 5074 1287 5088
rect 733 4973 747 4987
rect 693 4873 707 4887
rect 673 4854 687 4868
rect 753 4933 767 4947
rect 873 5032 887 5046
rect 833 4993 847 5007
rect 793 4893 807 4907
rect 753 4853 767 4867
rect 793 4854 807 4868
rect 873 4853 887 4867
rect 733 4832 747 4846
rect 613 4813 627 4827
rect 593 4733 607 4747
rect 473 4693 487 4707
rect 373 4573 387 4587
rect 293 4554 307 4568
rect 333 4553 347 4567
rect 593 4653 607 4667
rect 533 4613 547 4627
rect 533 4573 547 4587
rect 573 4573 587 4587
rect 473 4553 487 4567
rect 513 4554 527 4568
rect 113 4512 127 4526
rect 173 4512 187 4526
rect 73 4473 87 4487
rect 53 4333 67 4347
rect 133 4353 147 4367
rect 73 4292 87 4306
rect 33 4253 47 4267
rect 93 4034 107 4048
rect 193 4473 207 4487
rect 273 4473 287 4487
rect 233 4393 247 4407
rect 313 4393 327 4407
rect 213 4353 227 4367
rect 193 4333 207 4347
rect 253 4353 267 4367
rect 193 4293 207 4307
rect 173 4034 187 4048
rect 273 4292 287 4306
rect 233 4253 247 4267
rect 273 4113 287 4127
rect 233 4034 247 4048
rect 193 4013 207 4027
rect 113 3992 127 4006
rect 53 3933 67 3947
rect 53 3873 67 3887
rect 93 3873 107 3887
rect 253 3933 267 3947
rect 153 3853 167 3867
rect 53 3633 67 3647
rect 33 3593 47 3607
rect 13 3553 27 3567
rect 13 3513 27 3527
rect 13 3473 27 3487
rect 13 3393 27 3407
rect 13 3353 27 3367
rect 13 3313 27 3327
rect 133 3772 147 3786
rect 93 3613 107 3627
rect 73 3593 87 3607
rect 93 3553 107 3567
rect 113 3533 127 3547
rect 93 3472 107 3486
rect 253 3853 267 3867
rect 213 3833 227 3847
rect 273 3832 287 3846
rect 173 3772 187 3786
rect 233 3772 247 3786
rect 173 3553 187 3567
rect 233 3553 247 3567
rect 193 3514 207 3528
rect 333 4334 347 4348
rect 372 4334 386 4348
rect 533 4493 547 4507
rect 573 4493 587 4507
rect 773 4812 787 4826
rect 753 4773 767 4787
rect 733 4613 747 4627
rect 773 4613 787 4627
rect 753 4573 767 4587
rect 633 4512 647 4526
rect 733 4493 747 4507
rect 613 4473 627 4487
rect 673 4473 687 4487
rect 753 4453 767 4467
rect 733 4413 747 4427
rect 553 4393 567 4407
rect 593 4393 607 4407
rect 413 4353 427 4367
rect 453 4353 467 4367
rect 393 4333 407 4347
rect 353 4292 367 4306
rect 393 4293 407 4307
rect 493 4334 507 4348
rect 833 4793 847 4807
rect 813 4733 827 4747
rect 833 4713 847 4727
rect 913 5032 927 5046
rect 1053 5032 1067 5046
rect 1013 4993 1027 5007
rect 953 4933 967 4947
rect 1113 4973 1127 4987
rect 1253 5013 1267 5027
rect 1273 4993 1287 5007
rect 1193 4973 1207 4987
rect 1133 4933 1147 4947
rect 1253 4933 1267 4947
rect 993 4873 1007 4887
rect 1173 4873 1187 4887
rect 953 4854 967 4868
rect 1033 4854 1047 4868
rect 1193 4853 1207 4867
rect 1453 5373 1467 5387
rect 1653 5413 1667 5427
rect 1553 5374 1567 5388
rect 1593 5373 1607 5387
rect 1693 5374 1707 5388
rect 1753 5413 1767 5427
rect 1353 5313 1367 5327
rect 1413 5332 1427 5346
rect 1453 5332 1467 5346
rect 1493 5332 1507 5346
rect 1313 5073 1327 5087
rect 1513 5313 1527 5327
rect 1493 5273 1507 5287
rect 1453 5213 1467 5227
rect 1413 5113 1427 5127
rect 1333 4953 1347 4967
rect 1313 4913 1327 4927
rect 1293 4853 1307 4867
rect 1573 5333 1587 5347
rect 1533 5233 1547 5247
rect 1533 5193 1547 5207
rect 1573 5193 1587 5207
rect 1513 5153 1527 5167
rect 1453 5074 1467 5088
rect 1493 5074 1507 5088
rect 1773 5374 1787 5388
rect 1933 5433 1947 5447
rect 1853 5413 1867 5427
rect 1933 5374 1947 5388
rect 1973 5374 1987 5388
rect 2093 5433 2107 5447
rect 2053 5373 2067 5387
rect 2253 5413 2267 5427
rect 2393 5413 2407 5427
rect 2133 5374 2147 5388
rect 2193 5373 2207 5387
rect 2293 5374 2307 5388
rect 2333 5373 2347 5387
rect 2433 5374 2447 5388
rect 2473 5373 2487 5387
rect 2533 5374 2547 5388
rect 1753 5332 1767 5346
rect 1793 5332 1807 5346
rect 1993 5332 2007 5346
rect 2033 5332 2047 5346
rect 1673 5273 1687 5287
rect 1833 5273 1847 5287
rect 1953 5293 1967 5307
rect 1933 5253 1947 5267
rect 1633 5233 1647 5247
rect 1653 5173 1667 5187
rect 1673 5133 1687 5147
rect 1713 5133 1727 5147
rect 1913 5133 1927 5147
rect 1653 5073 1667 5087
rect 1433 5033 1447 5047
rect 1413 5013 1427 5027
rect 1373 4873 1387 4887
rect 1193 4793 1207 4807
rect 1273 4812 1287 4826
rect 1313 4812 1327 4826
rect 1393 4812 1407 4826
rect 1253 4773 1267 4787
rect 1353 4773 1367 4787
rect 1233 4753 1247 4767
rect 1353 4752 1367 4766
rect 1253 4733 1267 4747
rect 1033 4713 1047 4727
rect 1153 4713 1167 4727
rect 913 4673 927 4687
rect 873 4653 887 4667
rect 993 4593 1007 4607
rect 1053 4593 1067 4607
rect 813 4573 827 4587
rect 793 4533 807 4547
rect 953 4554 967 4568
rect 1093 4573 1107 4587
rect 1033 4554 1047 4568
rect 853 4473 867 4487
rect 933 4473 947 4487
rect 1013 4512 1027 4526
rect 1053 4493 1067 4507
rect 793 4413 807 4427
rect 693 4373 707 4387
rect 773 4373 787 4387
rect 673 4353 687 4367
rect 593 4334 607 4348
rect 633 4334 647 4348
rect 513 4292 527 4306
rect 553 4292 567 4306
rect 493 4273 507 4287
rect 473 4253 487 4267
rect 433 4113 447 4127
rect 413 4053 427 4067
rect 653 4292 667 4306
rect 953 4413 967 4427
rect 1053 4373 1067 4387
rect 733 4334 747 4348
rect 773 4334 787 4348
rect 833 4334 847 4348
rect 873 4334 887 4348
rect 913 4334 927 4348
rect 613 4253 627 4267
rect 613 4133 627 4147
rect 653 4133 667 4147
rect 613 4073 627 4087
rect 553 4052 567 4066
rect 393 3992 407 4006
rect 433 3993 447 4007
rect 393 3953 407 3967
rect 393 3913 407 3927
rect 353 3873 367 3887
rect 313 3833 327 3847
rect 353 3814 367 3828
rect 533 3973 547 3987
rect 493 3953 507 3967
rect 453 3913 467 3927
rect 573 3913 587 3927
rect 533 3853 547 3867
rect 333 3772 347 3786
rect 353 3633 367 3647
rect 273 3514 287 3528
rect 213 3433 227 3447
rect 253 3433 267 3447
rect 213 3393 227 3407
rect 53 3333 67 3347
rect 113 3333 127 3347
rect 153 3333 167 3347
rect 193 3333 207 3347
rect 33 3294 47 3308
rect 13 3273 27 3287
rect 33 3233 47 3247
rect 13 3113 27 3127
rect 73 3294 87 3308
rect 253 3333 267 3347
rect 433 3814 447 3828
rect 473 3814 487 3828
rect 493 3753 507 3767
rect 413 3573 427 3587
rect 473 3573 487 3587
rect 433 3514 447 3528
rect 473 3514 487 3528
rect 393 3453 407 3467
rect 433 3453 447 3467
rect 393 3294 407 3308
rect 253 3133 267 3147
rect 213 3093 227 3107
rect 53 3073 67 3087
rect 173 3073 187 3087
rect 233 3073 247 3087
rect 73 3033 87 3047
rect 113 2994 127 3008
rect 153 2953 167 2967
rect 133 2913 147 2927
rect 93 2813 107 2827
rect 132 2813 146 2827
rect 153 2813 167 2827
rect 33 2773 47 2787
rect 93 2774 107 2788
rect 133 2773 147 2787
rect 213 3033 227 3047
rect 213 2994 227 3008
rect 333 3193 347 3207
rect 293 3033 307 3047
rect 273 2994 287 3008
rect 593 3873 607 3887
rect 693 4292 707 4306
rect 713 4233 727 4247
rect 693 4093 707 4107
rect 673 4073 687 4087
rect 773 4213 787 4227
rect 873 4273 887 4287
rect 793 4173 807 4187
rect 773 4093 787 4107
rect 713 4053 727 4067
rect 613 3853 627 3867
rect 673 3853 687 3867
rect 613 3814 627 3828
rect 813 4034 827 4048
rect 753 3973 767 3987
rect 833 3993 847 4007
rect 793 3953 807 3967
rect 753 3873 767 3887
rect 793 3873 807 3887
rect 933 4293 947 4307
rect 892 4213 906 4227
rect 913 4213 927 4227
rect 913 4173 927 4187
rect 893 4113 907 4127
rect 873 4093 887 4107
rect 913 4053 927 4067
rect 1253 4633 1267 4647
rect 1193 4593 1207 4607
rect 1153 4554 1167 4568
rect 1113 4513 1127 4527
rect 1173 4512 1187 4526
rect 1153 4473 1167 4487
rect 1293 4573 1307 4587
rect 1333 4554 1347 4568
rect 1512 5033 1526 5047
rect 1533 5033 1547 5047
rect 1473 5013 1487 5027
rect 1593 5032 1607 5046
rect 1633 5032 1647 5046
rect 1873 5113 1887 5127
rect 1753 5074 1767 5088
rect 1793 5074 1807 5088
rect 1833 5074 1847 5088
rect 1653 5013 1667 5027
rect 1593 4993 1607 5007
rect 1573 4953 1587 4967
rect 1513 4933 1527 4947
rect 1573 4893 1587 4907
rect 1493 4854 1507 4868
rect 1533 4854 1547 4868
rect 1613 4933 1627 4947
rect 1453 4812 1467 4826
rect 1453 4733 1467 4747
rect 1372 4673 1386 4687
rect 1393 4673 1407 4687
rect 1433 4673 1447 4687
rect 1313 4512 1327 4526
rect 1353 4513 1367 4527
rect 1253 4453 1267 4467
rect 1213 4433 1227 4447
rect 1193 4373 1207 4387
rect 993 4292 1007 4306
rect 1033 4233 1047 4247
rect 1033 4212 1047 4226
rect 953 4173 967 4187
rect 1033 4133 1047 4147
rect 973 4113 987 4127
rect 873 4033 887 4047
rect 993 4053 1007 4067
rect 973 4033 987 4047
rect 893 3992 907 4006
rect 973 3993 987 4007
rect 933 3953 947 3967
rect 853 3913 867 3927
rect 913 3913 927 3927
rect 853 3873 867 3887
rect 833 3853 847 3867
rect 752 3813 766 3827
rect 773 3813 787 3827
rect 813 3814 827 3828
rect 673 3793 687 3807
rect 533 3772 547 3786
rect 593 3772 607 3786
rect 953 3853 967 3867
rect 1013 4033 1027 4047
rect 1153 4334 1167 4348
rect 1133 4293 1147 4307
rect 1353 4473 1367 4487
rect 1333 4373 1347 4387
rect 1393 4573 1407 4587
rect 1413 4554 1427 4568
rect 1513 4812 1527 4826
rect 1593 4813 1607 4827
rect 1513 4773 1527 4787
rect 1553 4773 1567 4787
rect 1493 4653 1507 4667
rect 1473 4613 1487 4627
rect 1473 4554 1487 4568
rect 1432 4513 1446 4527
rect 1433 4491 1447 4505
rect 1393 4473 1407 4487
rect 1493 4453 1507 4467
rect 1433 4413 1447 4427
rect 1373 4353 1387 4367
rect 1413 4353 1427 4367
rect 1313 4334 1327 4348
rect 1213 4292 1227 4306
rect 1253 4292 1267 4306
rect 1313 4253 1327 4267
rect 1173 4213 1187 4227
rect 1233 4133 1247 4147
rect 1073 4034 1087 4048
rect 1193 4034 1207 4048
rect 1053 3992 1067 4006
rect 1093 3993 1107 4007
rect 1253 4113 1267 4127
rect 1293 4053 1307 4067
rect 1373 4273 1387 4287
rect 1353 4233 1367 4247
rect 1333 4213 1347 4227
rect 1353 4173 1367 4187
rect 993 3933 1007 3947
rect 1053 3873 1067 3887
rect 953 3814 967 3828
rect 833 3772 847 3786
rect 873 3772 887 3786
rect 913 3773 927 3787
rect 673 3753 687 3767
rect 773 3753 787 3767
rect 573 3613 587 3627
rect 593 3593 607 3607
rect 633 3593 647 3607
rect 573 3553 587 3567
rect 553 3533 567 3547
rect 633 3553 647 3567
rect 673 3553 687 3567
rect 773 3553 787 3567
rect 853 3553 867 3567
rect 653 3514 667 3528
rect 573 3472 587 3486
rect 613 3472 627 3486
rect 653 3473 667 3487
rect 733 3514 747 3528
rect 813 3533 827 3547
rect 673 3433 687 3447
rect 573 3333 587 3347
rect 453 3294 467 3308
rect 513 3294 527 3308
rect 433 3193 447 3207
rect 473 3213 487 3227
rect 533 3213 547 3227
rect 493 3133 507 3147
rect 473 3073 487 3087
rect 373 3033 387 3047
rect 453 3033 467 3047
rect 373 2994 387 3008
rect 313 2953 327 2967
rect 253 2933 267 2947
rect 233 2913 247 2927
rect 233 2853 247 2867
rect 13 2613 27 2627
rect 13 2333 27 2347
rect 113 2732 127 2746
rect 73 2693 87 2707
rect 53 2473 67 2487
rect 93 2474 107 2488
rect 193 2732 207 2746
rect 313 2873 327 2887
rect 353 2873 367 2887
rect 313 2774 327 2788
rect 533 2952 547 2966
rect 493 2913 507 2927
rect 413 2853 427 2867
rect 393 2813 407 2827
rect 293 2732 307 2746
rect 373 2733 387 2747
rect 333 2653 347 2667
rect 233 2633 247 2647
rect 193 2513 207 2527
rect 333 2513 347 2527
rect 73 2432 87 2446
rect 33 2293 47 2307
rect 113 2293 127 2307
rect 73 2254 87 2268
rect 273 2473 287 2487
rect 373 2473 387 2487
rect 493 2813 507 2827
rect 413 2773 427 2787
rect 493 2773 507 2787
rect 433 2732 447 2746
rect 473 2732 487 2746
rect 533 2893 547 2907
rect 593 3293 607 3307
rect 653 3294 667 3308
rect 593 3252 607 3266
rect 633 3252 647 3266
rect 673 3252 687 3266
rect 673 3213 687 3227
rect 613 2994 627 3008
rect 693 2993 707 3007
rect 633 2952 647 2966
rect 593 2873 607 2887
rect 573 2833 587 2847
rect 673 2893 687 2907
rect 733 3433 747 3447
rect 1013 3772 1027 3786
rect 973 3673 987 3687
rect 1173 3933 1187 3947
rect 1173 3833 1187 3847
rect 1073 3813 1087 3827
rect 1133 3814 1147 3828
rect 993 3553 1007 3567
rect 1053 3553 1067 3567
rect 873 3533 887 3547
rect 893 3514 907 3528
rect 1033 3514 1047 3528
rect 1093 3773 1107 3774
rect 1093 3760 1107 3773
rect 1153 3713 1167 3727
rect 1273 3992 1287 4006
rect 1353 3913 1367 3927
rect 1313 3893 1327 3907
rect 1273 3833 1287 3847
rect 1233 3813 1247 3827
rect 1393 4213 1407 4227
rect 1493 4393 1507 4407
rect 1453 4373 1467 4387
rect 1493 4334 1507 4348
rect 1533 4693 1547 4707
rect 1553 4554 1567 4568
rect 1673 4973 1687 4987
rect 1653 4893 1667 4907
rect 1733 5013 1747 5027
rect 1913 5073 1927 5087
rect 1953 5173 1967 5187
rect 2133 5313 2147 5327
rect 2113 5293 2127 5307
rect 2193 5332 2207 5346
rect 2273 5332 2287 5346
rect 2233 5313 2247 5327
rect 2153 5293 2167 5307
rect 2173 5273 2187 5287
rect 2153 5233 2167 5247
rect 2073 5133 2087 5147
rect 2073 5093 2087 5107
rect 2033 5074 2047 5088
rect 2113 5093 2127 5107
rect 1813 5033 1827 5047
rect 1793 4973 1807 4987
rect 1693 4953 1707 4967
rect 1713 4913 1727 4927
rect 1673 4854 1687 4868
rect 1693 4812 1707 4826
rect 1733 4853 1747 4867
rect 1833 4953 1847 4967
rect 1893 5032 1907 5046
rect 1933 5033 1947 5047
rect 1853 4873 1867 4887
rect 1833 4854 1847 4868
rect 1873 4854 1887 4868
rect 2013 5032 2027 5046
rect 2073 5032 2087 5046
rect 2133 5032 2147 5046
rect 1993 5013 2007 5027
rect 1973 4933 1987 4947
rect 1633 4773 1647 4787
rect 1773 4812 1787 4826
rect 1753 4753 1767 4767
rect 1733 4693 1747 4707
rect 1693 4653 1707 4667
rect 1653 4633 1667 4647
rect 1673 4613 1687 4627
rect 1653 4573 1667 4587
rect 1553 4493 1567 4507
rect 1653 4513 1667 4527
rect 1633 4453 1647 4467
rect 1552 4433 1566 4447
rect 1573 4433 1587 4447
rect 1653 4433 1667 4447
rect 1813 4733 1827 4747
rect 1793 4653 1807 4667
rect 1833 4613 1847 4627
rect 1813 4593 1827 4607
rect 1793 4573 1807 4587
rect 1893 4653 1907 4667
rect 1893 4593 1907 4607
rect 1953 4812 1967 4826
rect 1933 4773 1947 4787
rect 1933 4633 1947 4647
rect 2013 4993 2027 5007
rect 2113 4993 2127 5007
rect 1993 4773 2007 4787
rect 2073 4854 2087 4868
rect 2033 4812 2047 4826
rect 2133 4913 2147 4927
rect 2233 5173 2247 5187
rect 2213 5133 2227 5147
rect 2373 5332 2387 5346
rect 2453 5333 2467 5347
rect 2413 5313 2427 5327
rect 2453 5293 2467 5307
rect 2473 5253 2487 5267
rect 2553 5273 2567 5287
rect 2513 5213 2527 5227
rect 2553 5213 2567 5227
rect 2353 5193 2367 5207
rect 2493 5193 2507 5207
rect 2333 5093 2347 5107
rect 2393 5133 2407 5147
rect 2253 5074 2267 5088
rect 2313 5074 2327 5088
rect 2353 5074 2367 5088
rect 2513 5153 2527 5167
rect 2552 5153 2566 5167
rect 2573 5153 2587 5167
rect 2493 5113 2507 5127
rect 2453 5093 2467 5107
rect 2233 5032 2247 5046
rect 2113 4773 2127 4787
rect 2013 4693 2027 4707
rect 2113 4673 2127 4687
rect 2173 4893 2187 4907
rect 2153 4873 2167 4887
rect 1716 4513 1730 4527
rect 1833 4554 1847 4568
rect 1973 4613 1987 4627
rect 2133 4613 2147 4627
rect 2013 4573 2027 4587
rect 2053 4573 2067 4587
rect 1813 4513 1827 4527
rect 1853 4512 1867 4526
rect 1913 4513 1927 4527
rect 1693 4493 1707 4507
rect 1733 4493 1747 4507
rect 1572 4373 1586 4387
rect 1593 4373 1607 4387
rect 1633 4334 1647 4348
rect 1433 4253 1447 4267
rect 1533 4293 1547 4307
rect 1473 4233 1487 4247
rect 1433 4193 1447 4207
rect 1433 4172 1447 4186
rect 1433 4113 1447 4127
rect 1473 4113 1487 4127
rect 1593 4253 1607 4267
rect 1573 4233 1587 4247
rect 1533 4213 1547 4227
rect 1553 4173 1567 4187
rect 1453 4073 1467 4087
rect 1413 4053 1427 4067
rect 1473 4053 1487 4067
rect 1533 4093 1547 4107
rect 1513 4053 1527 4067
rect 1493 4034 1507 4048
rect 1413 3973 1427 3987
rect 1453 3973 1467 3987
rect 1393 3873 1407 3887
rect 1373 3813 1387 3827
rect 1293 3772 1307 3786
rect 1253 3733 1267 3747
rect 1213 3673 1227 3687
rect 1293 3613 1307 3627
rect 1353 3772 1367 3786
rect 1393 3772 1407 3786
rect 1433 3772 1447 3786
rect 1433 3733 1447 3747
rect 1373 3553 1387 3567
rect 873 3472 887 3486
rect 753 3373 767 3387
rect 833 3333 847 3347
rect 773 3294 787 3308
rect 753 3252 767 3266
rect 1013 3453 1027 3467
rect 1113 3493 1127 3507
rect 1293 3513 1307 3527
rect 1333 3514 1347 3528
rect 1633 4273 1647 4287
rect 1613 4133 1627 4147
rect 1593 4113 1607 4127
rect 1593 4073 1607 4087
rect 1513 3993 1527 4007
rect 1573 3992 1587 4006
rect 1713 4433 1727 4447
rect 1793 4473 1807 4487
rect 1833 4473 1847 4487
rect 1773 4453 1787 4467
rect 1713 4233 1727 4247
rect 1833 4433 1847 4447
rect 1853 4373 1867 4387
rect 1813 4353 1827 4367
rect 1953 4512 1967 4526
rect 1993 4512 2007 4526
rect 2033 4513 2047 4527
rect 2013 4493 2027 4507
rect 2033 4453 2047 4467
rect 2093 4554 2107 4568
rect 2013 4433 2027 4447
rect 2053 4433 2067 4447
rect 2093 4433 2107 4447
rect 1913 4413 1927 4427
rect 1933 4393 1947 4407
rect 1993 4393 2007 4407
rect 1913 4373 1927 4387
rect 1913 4333 1927 4347
rect 1793 4253 1807 4267
rect 1833 4292 1847 4306
rect 1913 4293 1927 4307
rect 1833 4193 1847 4207
rect 1873 4193 1887 4207
rect 1813 4173 1827 4187
rect 1753 4113 1767 4127
rect 1673 4073 1687 4087
rect 1673 4052 1687 4066
rect 1713 4034 1727 4048
rect 1773 4033 1787 4047
rect 1853 4153 1867 4167
rect 1853 4073 1867 4087
rect 1873 4034 1887 4048
rect 1633 3992 1647 4006
rect 1613 3913 1627 3927
rect 1733 3992 1747 4006
rect 1693 3893 1707 3907
rect 1513 3853 1527 3867
rect 1493 3813 1507 3827
rect 1713 3873 1727 3887
rect 1693 3834 1707 3848
rect 1973 4373 1987 4387
rect 1993 4353 2007 4367
rect 2193 4873 2207 4887
rect 2173 4853 2187 4867
rect 2293 5033 2307 5047
rect 2273 4913 2287 4927
rect 2253 4854 2267 4868
rect 2193 4812 2207 4826
rect 2253 4793 2267 4807
rect 2233 4773 2247 4787
rect 2173 4633 2187 4647
rect 2153 4453 2167 4467
rect 2213 4593 2227 4607
rect 2393 5013 2407 5027
rect 2313 4993 2327 5007
rect 2373 4993 2387 5007
rect 2573 5073 2587 5087
rect 2473 5013 2487 5027
rect 2519 5013 2533 5027
rect 2453 4993 2467 5007
rect 2493 4993 2507 5007
rect 2392 4953 2406 4967
rect 2413 4953 2427 4967
rect 2413 4932 2427 4946
rect 2353 4913 2367 4927
rect 2412 4893 2426 4907
rect 2433 4893 2447 4907
rect 2493 4913 2507 4927
rect 2433 4853 2447 4867
rect 2573 4993 2587 5007
rect 2553 4893 2567 4907
rect 2533 4854 2547 4868
rect 2333 4812 2347 4826
rect 2413 4813 2427 4827
rect 2393 4793 2407 4807
rect 2413 4753 2427 4767
rect 2393 4733 2407 4747
rect 2373 4713 2387 4727
rect 2393 4673 2407 4687
rect 2333 4633 2347 4647
rect 2293 4593 2307 4607
rect 2253 4554 2267 4568
rect 2293 4553 2307 4567
rect 2333 4554 2347 4568
rect 2513 4812 2527 4826
rect 2473 4773 2487 4787
rect 2453 4713 2467 4727
rect 2433 4673 2447 4687
rect 2413 4633 2427 4647
rect 2173 4413 2187 4427
rect 2113 4393 2127 4407
rect 2013 4334 2027 4348
rect 1933 4233 1947 4247
rect 1993 4233 2007 4247
rect 1973 4193 1987 4207
rect 1933 4113 1947 4127
rect 1933 4053 1947 4067
rect 1913 4033 1927 4047
rect 2013 4133 2027 4147
rect 2073 4334 2087 4348
rect 2133 4292 2147 4306
rect 2273 4513 2287 4527
rect 2433 4593 2447 4607
rect 2353 4512 2367 4526
rect 2413 4512 2427 4526
rect 2313 4493 2327 4507
rect 2293 4473 2307 4487
rect 2273 4433 2287 4447
rect 2253 4393 2267 4407
rect 2233 4353 2247 4367
rect 2333 4473 2347 4487
rect 2333 4433 2347 4447
rect 2393 4413 2407 4427
rect 2313 4333 2327 4347
rect 2193 4253 2207 4267
rect 2273 4292 2287 4306
rect 2233 4233 2247 4247
rect 2173 4153 2187 4167
rect 2233 4153 2247 4167
rect 2093 4133 2107 4147
rect 2133 4133 2147 4147
rect 1813 3992 1827 4006
rect 1773 3913 1787 3927
rect 1733 3853 1747 3867
rect 1693 3813 1707 3827
rect 1753 3813 1767 3827
rect 1613 3793 1627 3807
rect 1493 3773 1507 3787
rect 1573 3772 1587 3786
rect 1593 3733 1607 3747
rect 1533 3713 1547 3727
rect 1493 3633 1507 3647
rect 1113 3433 1127 3447
rect 1273 3473 1287 3487
rect 1193 3433 1207 3447
rect 1133 3393 1147 3407
rect 1173 3333 1187 3347
rect 893 3294 907 3308
rect 933 3294 947 3308
rect 993 3293 1007 3307
rect 1033 3294 1047 3308
rect 1093 3294 1107 3308
rect 733 3213 747 3227
rect 953 3252 967 3266
rect 1353 3453 1367 3467
rect 1473 3513 1487 3527
rect 1513 3514 1527 3528
rect 1553 3633 1567 3647
rect 1493 3472 1507 3486
rect 1493 3451 1507 3465
rect 1533 3453 1547 3467
rect 1233 3313 1247 3327
rect 1273 3313 1287 3327
rect 1093 3252 1107 3266
rect 733 2952 747 2966
rect 1033 2994 1047 3008
rect 1193 3252 1207 3266
rect 1293 3294 1307 3308
rect 1333 3293 1347 3307
rect 1273 3252 1287 3266
rect 1253 3213 1267 3227
rect 1233 3073 1247 3087
rect 1253 3053 1267 3067
rect 1133 3033 1147 3047
rect 1113 2994 1127 3008
rect 873 2952 887 2966
rect 933 2952 947 2966
rect 973 2952 987 2966
rect 773 2913 787 2927
rect 853 2913 867 2927
rect 693 2873 707 2887
rect 693 2833 707 2847
rect 533 2773 547 2787
rect 633 2793 647 2807
rect 653 2773 667 2787
rect 993 2913 1007 2927
rect 813 2813 827 2827
rect 873 2813 887 2827
rect 953 2813 967 2827
rect 793 2793 807 2807
rect 733 2774 747 2788
rect 553 2732 567 2746
rect 593 2732 607 2746
rect 833 2793 847 2807
rect 813 2773 827 2787
rect 873 2774 887 2788
rect 932 2773 946 2787
rect 953 2773 967 2787
rect 1053 2952 1067 2966
rect 1413 3433 1427 3447
rect 1453 3433 1467 3447
rect 1433 3294 1447 3308
rect 1533 3393 1547 3407
rect 1513 3313 1527 3327
rect 1493 3293 1507 3307
rect 1433 3213 1447 3227
rect 1413 3193 1427 3207
rect 1353 3133 1367 3147
rect 1373 3033 1387 3047
rect 1153 2994 1167 3008
rect 1373 2994 1387 3008
rect 1213 2913 1227 2927
rect 1133 2853 1147 2867
rect 1013 2813 1027 2827
rect 1293 2813 1307 2827
rect 1033 2774 1047 2788
rect 1113 2774 1127 2788
rect 1153 2774 1167 2788
rect 1193 2774 1207 2788
rect 793 2753 807 2767
rect 513 2693 527 2707
rect 553 2653 567 2667
rect 653 2732 667 2746
rect 713 2732 727 2746
rect 853 2732 867 2746
rect 753 2693 767 2707
rect 893 2693 907 2707
rect 973 2732 987 2746
rect 1013 2732 1027 2746
rect 1193 2733 1207 2747
rect 1273 2732 1287 2746
rect 993 2693 1007 2707
rect 1033 2693 1047 2707
rect 1133 2693 1147 2707
rect 1353 2853 1367 2867
rect 1493 3253 1507 3267
rect 1453 3073 1467 3087
rect 1473 2994 1487 3008
rect 1633 3772 1647 3786
rect 1673 3772 1687 3786
rect 1713 3772 1727 3786
rect 1693 3713 1707 3727
rect 1613 3673 1627 3687
rect 1633 3633 1647 3647
rect 1593 3553 1607 3567
rect 1673 3533 1687 3547
rect 1713 3673 1727 3687
rect 1793 3853 1807 3867
rect 1893 3993 1907 4007
rect 1953 3992 1967 4006
rect 1893 3953 1907 3967
rect 1853 3933 1867 3947
rect 1833 3893 1847 3907
rect 1793 3813 1807 3827
rect 1853 3873 1867 3887
rect 1993 3933 2007 3947
rect 2033 3893 2047 3907
rect 2073 4053 2087 4067
rect 2153 4034 2167 4048
rect 2093 3953 2107 3967
rect 2113 3893 2127 3907
rect 1933 3873 1947 3887
rect 2073 3873 2087 3887
rect 1913 3853 1927 3867
rect 1933 3833 1947 3847
rect 1853 3773 1867 3787
rect 1813 3733 1827 3747
rect 1793 3713 1807 3727
rect 1953 3814 1967 3828
rect 1933 3772 1947 3786
rect 2073 3772 2087 3786
rect 2013 3753 2027 3767
rect 1873 3733 1887 3747
rect 1913 3733 1927 3747
rect 1973 3733 1987 3747
rect 1873 3653 1887 3667
rect 1793 3513 1807 3527
rect 1733 3472 1747 3486
rect 1773 3472 1787 3486
rect 1813 3472 1827 3486
rect 1613 3453 1627 3467
rect 1673 3453 1687 3467
rect 1713 3433 1727 3447
rect 1613 3353 1627 3367
rect 1553 3313 1567 3327
rect 1533 3253 1547 3267
rect 1533 3213 1547 3227
rect 1553 3193 1567 3207
rect 1893 3613 1907 3627
rect 1933 3533 1947 3547
rect 1913 3513 1927 3527
rect 1993 3514 2007 3528
rect 2113 3713 2127 3727
rect 2033 3633 2047 3647
rect 1893 3493 1907 3507
rect 1913 3473 1927 3487
rect 2013 3473 2027 3487
rect 1873 3453 1887 3467
rect 1873 3432 1887 3446
rect 1733 3393 1747 3407
rect 1773 3393 1787 3407
rect 1853 3393 1867 3407
rect 1753 3373 1767 3387
rect 1793 3373 1807 3387
rect 1993 3413 2007 3427
rect 1873 3373 1887 3387
rect 1913 3373 1927 3387
rect 1633 3293 1647 3307
rect 1673 3294 1687 3308
rect 1713 3294 1727 3308
rect 1873 3333 1887 3347
rect 1953 3333 1967 3347
rect 1833 3313 1847 3327
rect 1793 3294 1807 3308
rect 1753 3273 1767 3287
rect 1653 3252 1667 3266
rect 1673 3233 1687 3247
rect 1613 3153 1627 3167
rect 1573 3133 1587 3147
rect 1553 3113 1567 3127
rect 1533 3073 1547 3087
rect 1513 2994 1527 3008
rect 1453 2952 1467 2966
rect 1413 2833 1427 2847
rect 1413 2812 1427 2826
rect 1553 3033 1567 3047
rect 1573 3013 1587 3027
rect 1733 3253 1747 3267
rect 1693 3213 1707 3227
rect 1533 2952 1547 2966
rect 1573 2952 1587 2966
rect 1513 2913 1527 2927
rect 1533 2893 1547 2907
rect 1513 2833 1527 2847
rect 1493 2793 1507 2807
rect 1593 2774 1607 2788
rect 1693 3013 1707 3027
rect 1813 3252 1827 3266
rect 1853 3253 1867 3267
rect 1853 3213 1867 3227
rect 1813 3173 1827 3187
rect 1753 3093 1767 3107
rect 1733 2993 1747 3007
rect 1653 2952 1667 2966
rect 1713 2952 1727 2966
rect 1853 3113 1867 3127
rect 1913 3294 1927 3308
rect 1993 3173 2007 3187
rect 2273 4133 2287 4147
rect 2233 4034 2247 4048
rect 2213 3992 2227 4006
rect 2173 3953 2187 3967
rect 2353 4292 2367 4306
rect 2413 4292 2427 4306
rect 2313 4073 2327 4087
rect 2293 4033 2307 4047
rect 2393 4193 2407 4207
rect 2373 4073 2387 4087
rect 2172 3932 2186 3946
rect 2193 3933 2207 3947
rect 2273 3933 2287 3947
rect 2333 3933 2347 3947
rect 2173 3893 2187 3907
rect 2333 3893 2347 3907
rect 2193 3833 2207 3847
rect 2353 3833 2367 3847
rect 2253 3753 2267 3767
rect 2193 3673 2207 3687
rect 2133 3633 2147 3647
rect 2073 3573 2087 3587
rect 2113 3573 2127 3587
rect 2053 3553 2067 3567
rect 2113 3533 2127 3547
rect 2073 3513 2087 3527
rect 2153 3514 2167 3528
rect 2073 3473 2087 3487
rect 2053 3453 2067 3467
rect 2073 3413 2087 3427
rect 2173 3473 2187 3487
rect 2133 3453 2147 3467
rect 2093 3393 2107 3407
rect 2073 3373 2087 3387
rect 2033 3313 2047 3327
rect 2133 3373 2147 3387
rect 2093 3313 2107 3327
rect 2153 3353 2167 3367
rect 2293 3553 2307 3567
rect 2253 3514 2267 3528
rect 2513 4753 2527 4767
rect 2513 4732 2527 4746
rect 2473 4554 2487 4568
rect 2953 5473 2967 5487
rect 3013 5473 3027 5487
rect 2933 5453 2947 5467
rect 2633 5433 2647 5447
rect 2753 5413 2767 5427
rect 2793 5413 2807 5427
rect 2933 5413 2947 5427
rect 2633 5374 2647 5388
rect 2673 5374 2687 5388
rect 2733 5373 2747 5387
rect 2913 5374 2927 5388
rect 2613 5313 2627 5327
rect 2613 5173 2627 5187
rect 2813 5332 2827 5346
rect 2713 5273 2727 5287
rect 2673 5213 2687 5227
rect 2653 5133 2667 5147
rect 2893 5332 2907 5346
rect 2933 5332 2947 5346
rect 2893 5293 2907 5307
rect 2873 5253 2887 5267
rect 2873 5232 2887 5246
rect 2773 5193 2787 5207
rect 2813 5193 2827 5207
rect 2813 5153 2827 5167
rect 2913 5273 2927 5287
rect 2913 5213 2927 5227
rect 2813 5113 2827 5127
rect 2852 5113 2866 5127
rect 2873 5113 2887 5127
rect 2753 5093 2767 5107
rect 2673 5074 2687 5088
rect 2813 5074 2827 5088
rect 2973 5173 2987 5187
rect 2953 5113 2967 5127
rect 2733 5053 2747 5067
rect 2613 5032 2627 5046
rect 2653 5032 2667 5046
rect 2673 4993 2687 5007
rect 2713 5013 2727 5027
rect 2753 5033 2767 5047
rect 2733 4953 2747 4967
rect 2813 5013 2827 5027
rect 2793 4953 2807 4967
rect 2692 4933 2706 4947
rect 2713 4933 2727 4947
rect 2753 4933 2767 4947
rect 2693 4893 2707 4907
rect 2673 4873 2687 4887
rect 2733 4893 2747 4907
rect 2593 4853 2607 4867
rect 2633 4854 2647 4868
rect 2773 4854 2787 4868
rect 2593 4813 2607 4827
rect 2573 4713 2587 4727
rect 2573 4593 2587 4607
rect 2573 4512 2587 4526
rect 2533 4473 2547 4487
rect 2493 4453 2507 4467
rect 2573 4453 2587 4467
rect 2573 4413 2587 4427
rect 2533 4353 2547 4367
rect 2453 4333 2467 4347
rect 2493 4334 2507 4348
rect 2553 4292 2567 4306
rect 2713 4812 2727 4826
rect 2673 4773 2687 4787
rect 2613 4753 2627 4767
rect 2733 4793 2747 4807
rect 2692 4733 2706 4747
rect 2713 4733 2727 4747
rect 2632 4633 2646 4647
rect 2653 4633 2667 4647
rect 2613 4593 2627 4607
rect 2653 4573 2667 4587
rect 2793 4813 2807 4827
rect 2753 4773 2767 4787
rect 2793 4693 2807 4707
rect 2893 4953 2907 4967
rect 2873 4893 2887 4907
rect 2833 4873 2847 4887
rect 2973 5032 2987 5046
rect 3053 5453 3067 5467
rect 3133 5453 3147 5467
rect 3253 5453 3267 5467
rect 3073 5433 3087 5447
rect 3113 5433 3127 5447
rect 3192 5433 3206 5447
rect 3213 5433 3227 5447
rect 3033 5373 3047 5387
rect 3073 5374 3087 5388
rect 3053 5332 3067 5346
rect 3093 5332 3107 5346
rect 3133 5393 3147 5407
rect 3193 5393 3207 5407
rect 3173 5374 3187 5388
rect 3053 5293 3067 5307
rect 3053 5253 3067 5267
rect 3193 5332 3207 5346
rect 3233 5333 3247 5347
rect 3353 5413 3367 5427
rect 3313 5374 3327 5388
rect 3493 5453 3507 5467
rect 3393 5374 3407 5388
rect 3453 5374 3467 5388
rect 3773 5473 3787 5487
rect 3833 5473 3847 5487
rect 3673 5453 3687 5467
rect 3713 5453 3727 5467
rect 3693 5433 3707 5447
rect 3533 5393 3547 5407
rect 3513 5374 3527 5388
rect 3293 5332 3307 5346
rect 3233 5292 3247 5306
rect 3293 5293 3307 5307
rect 3273 5273 3287 5287
rect 3093 5233 3107 5247
rect 3153 5233 3167 5247
rect 3073 5213 3087 5227
rect 3092 5173 3106 5187
rect 3113 5173 3127 5187
rect 3073 5113 3087 5127
rect 3153 5153 3167 5167
rect 3113 5074 3127 5088
rect 3053 5032 3067 5046
rect 2933 4933 2947 4947
rect 2933 4912 2947 4926
rect 2913 4893 2927 4907
rect 2893 4873 2907 4887
rect 2933 4853 2947 4867
rect 2853 4812 2867 4826
rect 2853 4773 2867 4787
rect 2913 4793 2927 4807
rect 2913 4753 2927 4767
rect 2893 4733 2907 4747
rect 2833 4673 2847 4687
rect 2873 4673 2887 4687
rect 2933 4673 2947 4687
rect 2733 4593 2747 4607
rect 2633 4512 2647 4526
rect 2653 4493 2667 4507
rect 2613 4413 2627 4427
rect 2693 4473 2707 4487
rect 2673 4373 2687 4387
rect 2613 4333 2627 4347
rect 2733 4572 2747 4586
rect 2813 4573 2827 4587
rect 2713 4433 2727 4447
rect 2693 4353 2707 4367
rect 2773 4554 2787 4568
rect 2753 4513 2767 4527
rect 2792 4514 2806 4528
rect 2753 4413 2767 4427
rect 2853 4512 2867 4526
rect 3013 5013 3027 5027
rect 3133 4993 3147 5007
rect 3093 4913 3107 4927
rect 2973 4893 2987 4907
rect 3113 4873 3127 4887
rect 2993 4854 3007 4868
rect 3033 4854 3047 4868
rect 3093 4854 3107 4868
rect 2973 4813 2987 4827
rect 3013 4812 3027 4826
rect 3053 4793 3067 4807
rect 2973 4673 2987 4687
rect 3013 4673 3027 4687
rect 2953 4613 2967 4627
rect 2933 4593 2947 4607
rect 2973 4593 2987 4607
rect 2973 4554 2987 4568
rect 2833 4453 2847 4467
rect 2893 4493 2907 4507
rect 2993 4513 3007 4527
rect 2892 4433 2906 4447
rect 2913 4433 2927 4447
rect 2953 4433 2967 4447
rect 2993 4433 3007 4447
rect 2853 4413 2867 4427
rect 2793 4393 2807 4407
rect 2793 4372 2807 4386
rect 2893 4373 2907 4387
rect 2833 4334 2847 4348
rect 2873 4333 2887 4347
rect 2653 4292 2667 4306
rect 2693 4292 2707 4306
rect 2733 4292 2747 4306
rect 2773 4292 2787 4306
rect 2673 4273 2687 4287
rect 2793 4273 2807 4287
rect 2593 4233 2607 4247
rect 2653 4233 2667 4247
rect 2493 4213 2507 4227
rect 2473 4173 2487 4187
rect 2453 4133 2467 4147
rect 2433 4053 2447 4067
rect 2393 3992 2407 4006
rect 2413 3973 2427 3987
rect 2473 3993 2487 4007
rect 2433 3953 2447 3967
rect 2553 4113 2567 4127
rect 2713 4213 2727 4227
rect 2793 4173 2807 4187
rect 2673 4133 2687 4147
rect 2713 4133 2727 4147
rect 2553 4053 2567 4067
rect 2593 4034 2607 4048
rect 2633 4034 2647 4048
rect 2713 4034 2727 4048
rect 2513 3953 2527 3967
rect 2513 3932 2527 3946
rect 2493 3913 2507 3927
rect 2473 3853 2487 3867
rect 2373 3814 2387 3828
rect 2433 3814 2447 3828
rect 2473 3814 2487 3828
rect 2353 3673 2367 3687
rect 2353 3633 2367 3647
rect 2413 3593 2427 3607
rect 2453 3573 2467 3587
rect 2493 3753 2507 3767
rect 2573 3973 2587 3987
rect 2533 3913 2547 3927
rect 2653 3992 2667 4006
rect 2713 3993 2727 4007
rect 2753 3992 2767 4006
rect 2593 3953 2607 3967
rect 2653 3953 2667 3967
rect 2593 3873 2607 3887
rect 2573 3853 2587 3867
rect 2553 3814 2567 3828
rect 2573 3753 2587 3767
rect 2613 3753 2627 3767
rect 2713 3814 2727 3828
rect 2773 3813 2787 3827
rect 2693 3772 2707 3786
rect 2773 3753 2787 3767
rect 2853 4293 2867 4307
rect 2833 4213 2847 4227
rect 2953 4353 2967 4367
rect 2913 4333 2927 4347
rect 2893 4273 2907 4287
rect 2993 4293 3007 4307
rect 2933 4253 2947 4267
rect 3233 5233 3247 5247
rect 3193 5193 3207 5207
rect 3253 5193 3267 5207
rect 3173 5073 3187 5087
rect 3233 5133 3247 5147
rect 3313 5213 3327 5227
rect 3393 5333 3407 5347
rect 3433 5332 3447 5346
rect 3513 5333 3527 5347
rect 3593 5374 3607 5388
rect 3753 5413 3767 5427
rect 3793 5374 3807 5388
rect 3473 5293 3487 5307
rect 3373 5253 3387 5267
rect 3433 5253 3447 5267
rect 3493 5273 3507 5287
rect 3473 5253 3487 5267
rect 3453 5213 3467 5227
rect 3333 5193 3347 5207
rect 3353 5153 3367 5167
rect 3293 5133 3307 5147
rect 3353 5113 3367 5127
rect 3333 5093 3347 5107
rect 3313 5073 3327 5087
rect 3173 5033 3187 5047
rect 3153 4873 3167 4887
rect 3293 5033 3307 5047
rect 3253 4992 3267 5006
rect 3213 4973 3227 4987
rect 3353 5073 3367 5087
rect 3413 5074 3427 5088
rect 3332 5033 3346 5047
rect 3353 5033 3367 5047
rect 3453 5033 3467 5047
rect 3433 5013 3447 5027
rect 3353 4993 3367 5007
rect 3393 4993 3407 5007
rect 3533 5313 3547 5327
rect 3513 5193 3527 5207
rect 3553 5293 3567 5307
rect 3553 5253 3567 5267
rect 3693 5332 3707 5346
rect 3733 5332 3747 5346
rect 3653 5313 3667 5327
rect 3713 5313 3727 5327
rect 3633 5293 3647 5307
rect 3573 5233 3587 5247
rect 3613 5233 3627 5247
rect 3593 5213 3607 5227
rect 3813 5333 3827 5347
rect 3773 5293 3787 5307
rect 3713 5273 3727 5287
rect 3693 5253 3707 5267
rect 3633 5193 3647 5207
rect 3533 5153 3547 5167
rect 3573 5133 3587 5147
rect 3533 5113 3547 5127
rect 3533 5092 3547 5106
rect 3493 5073 3507 5087
rect 3573 5074 3587 5088
rect 3753 5193 3767 5207
rect 3713 5173 3727 5187
rect 3713 5093 3727 5107
rect 3613 5073 3627 5087
rect 3693 5074 3707 5088
rect 3513 5032 3527 5046
rect 3473 5013 3487 5027
rect 3593 5033 3607 5047
rect 3533 4993 3547 5007
rect 3573 4993 3587 5007
rect 3453 4953 3467 4967
rect 3293 4933 3307 4947
rect 3393 4913 3407 4927
rect 3333 4893 3347 4907
rect 3373 4853 3387 4867
rect 3113 4812 3127 4826
rect 3213 4812 3227 4826
rect 3253 4812 3267 4826
rect 3333 4812 3347 4826
rect 3453 4854 3467 4868
rect 3413 4812 3427 4826
rect 3573 4953 3587 4967
rect 3593 4933 3607 4947
rect 3393 4793 3407 4807
rect 3293 4773 3307 4787
rect 3333 4773 3347 4787
rect 3373 4773 3387 4787
rect 3093 4753 3107 4767
rect 3053 4673 3067 4687
rect 3053 4633 3067 4647
rect 3113 4613 3127 4627
rect 3193 4613 3207 4627
rect 3293 4613 3307 4627
rect 3033 4553 3047 4567
rect 3073 4554 3087 4568
rect 3053 4373 3067 4387
rect 3033 4353 3047 4367
rect 3253 4553 3267 4567
rect 3373 4733 3387 4747
rect 3333 4554 3347 4568
rect 3473 4753 3487 4767
rect 3493 4713 3507 4727
rect 3413 4673 3427 4687
rect 3393 4633 3407 4647
rect 3433 4593 3447 4607
rect 3393 4553 3407 4567
rect 3473 4554 3487 4568
rect 3173 4512 3187 4526
rect 3213 4512 3227 4526
rect 3253 4512 3267 4526
rect 3313 4512 3327 4526
rect 3373 4513 3387 4527
rect 3413 4512 3427 4526
rect 3113 4413 3127 4427
rect 3253 4473 3267 4487
rect 3293 4473 3307 4487
rect 3393 4473 3407 4487
rect 3233 4393 3247 4407
rect 3293 4413 3307 4427
rect 3273 4393 3287 4407
rect 3153 4373 3167 4387
rect 3253 4373 3267 4387
rect 3253 4352 3267 4366
rect 3213 4334 3227 4348
rect 3153 4312 3167 4326
rect 2873 4153 2887 4167
rect 2933 4153 2947 4167
rect 2973 4153 2987 4167
rect 3013 4153 3027 4167
rect 2853 4093 2867 4107
rect 2893 4073 2907 4087
rect 2853 4034 2867 4048
rect 2893 4034 2907 4048
rect 2953 4093 2967 4107
rect 2833 3993 2847 4007
rect 2813 3953 2827 3967
rect 2813 3873 2827 3887
rect 2913 3992 2927 4006
rect 2873 3953 2887 3967
rect 2833 3833 2847 3847
rect 2793 3733 2807 3747
rect 2853 3733 2867 3747
rect 2893 3893 2907 3907
rect 2893 3853 2907 3867
rect 2873 3713 2887 3727
rect 2733 3673 2747 3687
rect 2893 3673 2907 3687
rect 2513 3633 2527 3647
rect 2653 3633 2667 3647
rect 2833 3633 2847 3647
rect 2533 3573 2547 3587
rect 2753 3573 2767 3587
rect 2433 3553 2447 3567
rect 2213 3473 2227 3487
rect 2273 3472 2287 3486
rect 2313 3472 2327 3486
rect 2373 3514 2387 3528
rect 2413 3514 2427 3528
rect 2393 3472 2407 3486
rect 2433 3453 2447 3467
rect 2233 3433 2247 3447
rect 2333 3433 2347 3447
rect 2373 3433 2387 3447
rect 2213 3373 2227 3387
rect 2193 3353 2207 3367
rect 2353 3353 2367 3367
rect 2153 3294 2167 3308
rect 2013 3133 2027 3147
rect 1933 3113 1947 3127
rect 1972 3113 1986 3127
rect 1993 3113 2007 3127
rect 1873 3073 1887 3087
rect 1973 3053 1987 3067
rect 1953 3033 1967 3047
rect 1793 2952 1807 2966
rect 1753 2933 1767 2947
rect 1773 2893 1787 2907
rect 1713 2793 1727 2807
rect 1653 2774 1667 2788
rect 1473 2732 1487 2746
rect 1513 2732 1527 2746
rect 1793 2853 1807 2867
rect 1793 2832 1807 2846
rect 1793 2773 1807 2787
rect 1973 3013 1987 3027
rect 2133 3253 2147 3267
rect 2173 3252 2187 3266
rect 2093 3233 2107 3247
rect 2073 3133 2087 3147
rect 2053 3073 2067 3087
rect 1893 2913 1907 2927
rect 1953 2913 1967 2927
rect 2133 3113 2147 3127
rect 2093 3073 2107 3087
rect 2113 3053 2127 3067
rect 2093 2993 2107 3007
rect 1993 2953 2007 2967
rect 2093 2953 2107 2967
rect 1973 2873 1987 2887
rect 2033 2833 2047 2847
rect 2013 2793 2027 2807
rect 1773 2753 1787 2767
rect 2113 2933 2127 2947
rect 2233 3173 2247 3187
rect 2213 3153 2227 3167
rect 2253 3133 2267 3147
rect 2213 3113 2227 3127
rect 2173 2994 2187 3008
rect 2253 3073 2267 3087
rect 2153 2953 2167 2967
rect 2133 2813 2147 2827
rect 2093 2793 2107 2807
rect 2193 2952 2207 2966
rect 2493 3514 2507 3528
rect 2573 3514 2587 3528
rect 2613 3514 2627 3528
rect 2653 3514 2667 3528
rect 2713 3514 2727 3528
rect 2793 3514 2807 3528
rect 2493 3393 2507 3407
rect 2473 3333 2487 3347
rect 2453 3313 2467 3327
rect 2433 3294 2447 3308
rect 2473 3252 2487 3266
rect 2473 3153 2487 3167
rect 2433 3113 2447 3127
rect 2373 3093 2387 3107
rect 2353 3073 2367 3087
rect 2333 3053 2347 3067
rect 2393 3053 2407 3067
rect 2293 2994 2307 3008
rect 2333 2994 2347 3008
rect 2313 2952 2327 2966
rect 2373 2952 2387 2966
rect 2613 3433 2627 3447
rect 2573 3413 2587 3427
rect 2513 3333 2527 3347
rect 2593 3333 2607 3347
rect 2513 3312 2527 3326
rect 2573 3294 2587 3308
rect 2513 3233 2527 3247
rect 2533 3153 2547 3167
rect 2493 3113 2507 3127
rect 2673 3453 2687 3467
rect 2713 3433 2727 3447
rect 2773 3413 2787 3427
rect 2793 3373 2807 3387
rect 2933 3953 2947 3967
rect 3013 4132 3027 4146
rect 3033 4113 3047 4127
rect 3053 4093 3067 4107
rect 3033 4053 3047 4067
rect 2973 4033 2987 4047
rect 3013 4034 3027 4048
rect 3113 4273 3127 4287
rect 3093 4253 3107 4267
rect 3373 4393 3387 4407
rect 3293 4333 3307 4347
rect 3333 4334 3347 4348
rect 3293 4293 3307 4307
rect 3453 4353 3467 4367
rect 3513 4633 3527 4647
rect 3573 4633 3587 4647
rect 3593 4593 3607 4607
rect 3553 4493 3567 4507
rect 3493 4413 3507 4427
rect 3573 4413 3587 4427
rect 3553 4373 3567 4387
rect 3533 4353 3547 4367
rect 3433 4334 3447 4348
rect 3473 4334 3487 4348
rect 3513 4334 3527 4348
rect 3253 4273 3267 4287
rect 3193 4253 3207 4267
rect 3093 4153 3107 4167
rect 3104 4133 3118 4147
rect 3213 4233 3227 4247
rect 3173 4193 3187 4207
rect 3213 4193 3227 4207
rect 3253 4173 3267 4187
rect 3233 4153 3247 4167
rect 3213 4133 3227 4147
rect 3104 4073 3118 4087
rect 3173 4072 3187 4086
rect 3073 4033 3087 4047
rect 2973 3993 2987 4007
rect 3213 4053 3227 4067
rect 3193 4033 3207 4047
rect 2953 3933 2967 3947
rect 2993 3933 3007 3947
rect 2933 3853 2947 3867
rect 2973 3893 2987 3907
rect 3053 3973 3067 3987
rect 2993 3873 3007 3887
rect 3033 3873 3047 3887
rect 2993 3833 3007 3847
rect 3013 3814 3027 3828
rect 2953 3753 2967 3767
rect 3033 3773 3047 3787
rect 2993 3713 3007 3727
rect 3033 3713 3047 3727
rect 2933 3613 2947 3627
rect 2973 3613 2987 3627
rect 2873 3573 2887 3587
rect 2913 3573 2927 3587
rect 2873 3514 2887 3528
rect 2953 3493 2967 3507
rect 2893 3453 2907 3467
rect 3012 3673 3026 3687
rect 3033 3673 3047 3687
rect 3153 3992 3167 4006
rect 3113 3973 3127 3987
rect 3173 3973 3187 3987
rect 3113 3833 3127 3847
rect 3173 3833 3187 3847
rect 3173 3812 3187 3826
rect 3093 3753 3107 3767
rect 3073 3693 3087 3707
rect 3053 3633 3067 3647
rect 3013 3593 3027 3607
rect 2993 3573 3007 3587
rect 2993 3514 3007 3528
rect 2973 3472 2987 3486
rect 3033 3472 3047 3486
rect 2953 3433 2967 3447
rect 2893 3413 2907 3427
rect 2853 3373 2867 3387
rect 2633 3353 2647 3367
rect 2673 3333 2687 3347
rect 2713 3313 2727 3327
rect 2833 3333 2847 3347
rect 2833 3293 2847 3307
rect 2753 3273 2767 3287
rect 2653 3252 2667 3266
rect 2693 3252 2707 3266
rect 2613 3213 2627 3227
rect 2733 3193 2747 3207
rect 2693 3133 2707 3147
rect 2633 3013 2647 3027
rect 2453 2952 2467 2966
rect 2393 2913 2407 2927
rect 2353 2853 2367 2867
rect 2253 2833 2267 2847
rect 2213 2813 2227 2827
rect 2033 2773 2047 2787
rect 2073 2774 2087 2788
rect 1373 2673 1387 2687
rect 1333 2653 1347 2667
rect 993 2633 1007 2647
rect 1033 2573 1047 2587
rect 1173 2573 1187 2587
rect 793 2533 807 2547
rect 833 2533 847 2547
rect 933 2533 947 2547
rect 493 2493 507 2507
rect 633 2493 647 2507
rect 153 2413 167 2427
rect 133 2273 147 2287
rect 213 2432 227 2446
rect 453 2474 467 2488
rect 553 2473 567 2487
rect 613 2474 627 2488
rect 673 2473 687 2487
rect 733 2474 747 2488
rect 273 2413 287 2427
rect 173 2333 187 2347
rect 353 2432 367 2446
rect 413 2432 427 2446
rect 173 2273 187 2287
rect 153 2253 167 2267
rect 53 2213 67 2227
rect 13 2173 27 2187
rect 133 2212 147 2226
rect 93 2173 107 2187
rect 233 2254 247 2268
rect 273 2254 287 2268
rect 213 2212 227 2226
rect 353 2254 367 2268
rect 513 2432 527 2446
rect 553 2432 567 2446
rect 633 2432 647 2446
rect 513 2293 527 2307
rect 593 2293 607 2307
rect 353 2213 367 2227
rect 173 1954 187 1968
rect 213 1954 227 1968
rect 253 1954 267 1968
rect 333 2093 347 2107
rect 393 2212 407 2226
rect 353 2033 367 2047
rect 413 2033 427 2047
rect 373 1993 387 2007
rect 153 1873 167 1887
rect 193 1833 207 1847
rect 93 1753 107 1767
rect 213 1734 227 1748
rect 353 1912 367 1926
rect 333 1873 347 1887
rect 93 1692 107 1706
rect 393 1833 407 1847
rect 253 1633 267 1647
rect 213 1593 227 1607
rect 173 1453 187 1467
rect 133 1434 147 1448
rect 93 1392 107 1406
rect 253 1553 267 1567
rect 313 1692 327 1706
rect 353 1692 367 1706
rect 553 2254 567 2268
rect 693 2433 707 2447
rect 873 2513 887 2527
rect 933 2473 947 2487
rect 753 2432 767 2446
rect 793 2432 807 2446
rect 853 2432 867 2446
rect 713 2413 727 2427
rect 693 2293 707 2307
rect 633 2273 647 2287
rect 673 2273 687 2287
rect 813 2353 827 2367
rect 753 2293 767 2307
rect 513 2212 527 2226
rect 573 2212 587 2226
rect 493 2173 507 2187
rect 613 2173 627 2187
rect 713 2254 727 2268
rect 933 2432 947 2446
rect 833 2333 847 2347
rect 893 2333 907 2347
rect 1113 2474 1127 2488
rect 1233 2553 1247 2567
rect 1273 2513 1287 2527
rect 1233 2473 1247 2487
rect 1353 2473 1367 2487
rect 993 2413 1007 2427
rect 1253 2432 1267 2446
rect 1133 2393 1147 2407
rect 1293 2393 1307 2407
rect 1293 2353 1307 2367
rect 1233 2313 1247 2327
rect 873 2293 887 2307
rect 953 2293 967 2307
rect 833 2253 847 2267
rect 893 2273 907 2287
rect 933 2273 947 2287
rect 973 2273 987 2287
rect 1033 2273 1047 2287
rect 913 2254 927 2268
rect 833 2213 847 2227
rect 893 2212 907 2226
rect 613 2152 627 2166
rect 673 2153 687 2167
rect 573 2093 587 2107
rect 453 2013 467 2027
rect 453 1954 467 1968
rect 433 1913 447 1927
rect 413 1753 427 1767
rect 473 1873 487 1887
rect 513 1873 527 1887
rect 593 2013 607 2027
rect 573 1833 587 1847
rect 473 1753 487 1767
rect 433 1734 447 1748
rect 693 2013 707 2027
rect 953 2213 967 2227
rect 813 2153 827 2167
rect 933 2153 947 2167
rect 733 1993 747 2007
rect 713 1973 727 1987
rect 953 2133 967 2147
rect 953 2093 967 2107
rect 1053 2253 1067 2267
rect 1353 2413 1367 2427
rect 1353 2293 1367 2307
rect 1333 2253 1347 2267
rect 1053 2212 1067 2226
rect 1093 2212 1107 2226
rect 853 2073 867 2087
rect 1033 2073 1047 2087
rect 1233 2212 1247 2226
rect 1273 2212 1287 2226
rect 1313 2212 1327 2226
rect 1733 2732 1747 2746
rect 1813 2653 1827 2667
rect 1953 2732 1967 2746
rect 2013 2732 2027 2746
rect 2053 2732 2067 2746
rect 2153 2773 2167 2787
rect 2253 2774 2267 2788
rect 2453 2873 2467 2887
rect 2513 2873 2527 2887
rect 2413 2853 2427 2867
rect 2693 2994 2707 3008
rect 2413 2813 2427 2827
rect 2573 2853 2587 2867
rect 2633 2853 2647 2867
rect 2153 2732 2167 2746
rect 2193 2732 2207 2746
rect 2353 2732 2367 2746
rect 2393 2733 2407 2747
rect 2533 2732 2547 2746
rect 2813 3252 2827 3266
rect 3093 3633 3107 3647
rect 3133 3613 3147 3627
rect 3113 3593 3127 3607
rect 3113 3513 3127 3527
rect 3213 3973 3227 3987
rect 3273 4153 3287 4167
rect 3253 4113 3267 4127
rect 3293 4133 3307 4147
rect 3333 4273 3347 4287
rect 3333 4173 3347 4187
rect 3373 4273 3387 4287
rect 3353 4133 3367 4147
rect 3313 4073 3327 4087
rect 3273 4034 3287 4048
rect 3433 4233 3447 4247
rect 3493 4273 3507 4287
rect 3513 4253 3527 4267
rect 3733 5053 3747 5067
rect 3673 5032 3687 5046
rect 4113 5453 4127 5467
rect 4133 5433 4147 5447
rect 4073 5413 4087 5427
rect 4013 5393 4027 5407
rect 3873 5374 3887 5388
rect 3973 5374 3987 5388
rect 4053 5393 4067 5407
rect 4153 5413 4167 5427
rect 4313 5413 4327 5427
rect 4133 5374 4147 5388
rect 4173 5374 4187 5388
rect 4213 5373 4227 5387
rect 4273 5374 4287 5388
rect 4073 5353 4087 5367
rect 3853 5333 3867 5347
rect 3833 5113 3847 5127
rect 3873 5273 3887 5287
rect 3873 5213 3887 5227
rect 3993 5332 4007 5346
rect 4033 5332 4047 5346
rect 4113 5332 4127 5346
rect 4073 5293 4087 5307
rect 4153 5273 4167 5287
rect 3993 5253 4007 5267
rect 4233 5333 4247 5347
rect 4213 5173 4227 5187
rect 4253 5273 4267 5287
rect 4393 5413 4407 5427
rect 4493 5413 4507 5427
rect 4433 5374 4447 5388
rect 4693 5433 4707 5447
rect 4913 5433 4927 5447
rect 4513 5373 4527 5387
rect 4553 5374 4567 5388
rect 4313 5313 4327 5327
rect 4353 5313 4367 5327
rect 4293 5233 4307 5247
rect 4033 5153 4047 5167
rect 4233 5153 4247 5167
rect 3893 5133 3907 5147
rect 3953 5133 3967 5147
rect 3993 5133 4007 5147
rect 3873 5113 3887 5127
rect 3853 5074 3867 5088
rect 3893 5093 3907 5107
rect 3993 5093 4007 5107
rect 3753 5013 3767 5027
rect 3633 4993 3647 5007
rect 3733 4993 3747 5007
rect 3773 4993 3787 5007
rect 3713 4913 3727 4927
rect 3673 4854 3687 4868
rect 3653 4813 3667 4827
rect 3733 4812 3747 4826
rect 3693 4773 3707 4787
rect 3653 4613 3667 4627
rect 3693 4554 3707 4568
rect 3893 5033 3907 5047
rect 4053 5093 4067 5107
rect 4113 5093 4127 5107
rect 3833 5013 3847 5027
rect 3793 4973 3807 4987
rect 3933 5032 3947 5046
rect 3973 5032 3987 5046
rect 4033 5032 4047 5046
rect 4153 5074 4167 5088
rect 4193 5073 4207 5087
rect 4453 5332 4467 5346
rect 4493 5332 4507 5346
rect 4453 5293 4467 5307
rect 4413 5233 4427 5247
rect 4453 5173 4467 5187
rect 4493 5173 4507 5187
rect 4413 5133 4427 5147
rect 4353 5113 4367 5127
rect 3933 4953 3947 4967
rect 4053 4953 4067 4967
rect 3913 4913 3927 4927
rect 3793 4893 3807 4907
rect 3893 4893 3907 4907
rect 3813 4854 3827 4868
rect 3853 4854 3867 4868
rect 4053 4932 4067 4946
rect 3993 4893 4007 4907
rect 3892 4853 3906 4867
rect 3913 4853 3927 4867
rect 3953 4854 3967 4868
rect 3993 4854 4007 4868
rect 3873 4812 3887 4826
rect 3973 4793 3987 4807
rect 3913 4773 3927 4787
rect 3893 4753 3907 4767
rect 3993 4753 4007 4767
rect 3833 4733 3847 4747
rect 4013 4733 4027 4747
rect 3993 4713 4007 4727
rect 4033 4673 4047 4687
rect 3893 4613 3907 4627
rect 3993 4613 4007 4627
rect 3773 4593 3787 4607
rect 3833 4553 3847 4567
rect 3933 4593 3947 4607
rect 4133 5032 4147 5046
rect 4193 5032 4207 5046
rect 4253 5032 4267 5046
rect 4253 4993 4267 5007
rect 4193 4953 4207 4967
rect 4092 4815 4106 4829
rect 4133 4812 4147 4826
rect 4093 4793 4107 4807
rect 4073 4713 4087 4727
rect 4353 5074 4367 5088
rect 4393 5074 4407 5088
rect 4433 5074 4447 5088
rect 4473 5133 4487 5147
rect 4333 4973 4347 4987
rect 4313 4953 4327 4967
rect 4353 4953 4367 4967
rect 4353 4893 4367 4907
rect 4413 5032 4427 5046
rect 4433 4973 4447 4987
rect 4293 4854 4307 4868
rect 4213 4813 4227 4827
rect 4193 4753 4207 4767
rect 4173 4673 4187 4687
rect 4073 4653 4087 4667
rect 4093 4633 4107 4647
rect 4073 4573 4087 4587
rect 4053 4553 4067 4567
rect 3613 4473 3627 4487
rect 3633 4433 3647 4447
rect 3733 4512 3747 4526
rect 3793 4512 3807 4526
rect 3833 4512 3847 4526
rect 3873 4512 3887 4526
rect 3933 4512 3947 4526
rect 3652 4413 3666 4427
rect 3673 4413 3687 4427
rect 3593 4373 3607 4387
rect 3613 4334 3627 4348
rect 3553 4273 3567 4287
rect 3633 4292 3647 4306
rect 3913 4493 3927 4507
rect 3813 4373 3827 4387
rect 3733 4334 3747 4348
rect 3773 4334 3787 4348
rect 3753 4292 3767 4306
rect 3673 4273 3687 4287
rect 3713 4273 3727 4287
rect 3493 4233 3507 4247
rect 3473 4213 3487 4227
rect 3533 4213 3547 4227
rect 3473 4192 3487 4206
rect 3453 4173 3467 4187
rect 3412 4153 3426 4167
rect 3433 4153 3447 4167
rect 3453 4133 3467 4147
rect 3413 4093 3427 4107
rect 3393 4053 3407 4067
rect 3453 4033 3467 4047
rect 3513 4173 3527 4187
rect 3553 4133 3567 4147
rect 3593 4133 3607 4147
rect 3533 4093 3547 4107
rect 3513 4053 3527 4067
rect 3673 4133 3687 4147
rect 3613 4072 3627 4086
rect 3593 4033 3607 4047
rect 3473 4013 3487 4027
rect 3293 3992 3307 4006
rect 3333 3992 3347 4006
rect 3373 3993 3387 4007
rect 3273 3973 3287 3987
rect 3233 3953 3247 3967
rect 3233 3932 3247 3946
rect 3253 3913 3267 3927
rect 3253 3833 3267 3847
rect 3233 3814 3247 3828
rect 3333 3953 3347 3967
rect 3333 3833 3347 3847
rect 3253 3772 3267 3786
rect 3293 3772 3307 3786
rect 3213 3753 3227 3767
rect 3173 3693 3187 3707
rect 3233 3713 3247 3727
rect 3213 3613 3227 3627
rect 3152 3593 3166 3607
rect 3173 3593 3187 3607
rect 3113 3473 3127 3487
rect 2873 3353 2887 3367
rect 3073 3353 3087 3367
rect 2993 3313 3007 3327
rect 2913 3294 2927 3308
rect 2972 3293 2986 3307
rect 3033 3294 3047 3308
rect 3073 3294 3087 3308
rect 2853 3193 2867 3207
rect 2933 3252 2947 3266
rect 2893 3173 2907 3187
rect 2913 3153 2927 3167
rect 2853 3133 2867 3147
rect 3152 3433 3166 3447
rect 3173 3433 3187 3447
rect 3193 3393 3207 3407
rect 3173 3353 3187 3367
rect 3193 3333 3207 3347
rect 3193 3294 3207 3308
rect 3433 3992 3447 4006
rect 3493 3993 3507 4007
rect 3493 3953 3507 3967
rect 3413 3933 3427 3947
rect 3553 3992 3567 4006
rect 3593 3993 3607 4007
rect 3453 3893 3467 3907
rect 3513 3893 3527 3907
rect 3433 3873 3447 3887
rect 3393 3814 3407 3828
rect 3453 3833 3467 3847
rect 3433 3813 3447 3827
rect 3533 3853 3547 3867
rect 3553 3814 3567 3828
rect 3333 3633 3347 3647
rect 3293 3573 3307 3587
rect 3253 3514 3267 3528
rect 3373 3753 3387 3767
rect 3373 3732 3387 3746
rect 3533 3772 3547 3786
rect 3573 3773 3587 3787
rect 3493 3733 3507 3747
rect 3393 3633 3407 3647
rect 3433 3633 3447 3647
rect 3433 3593 3447 3607
rect 3553 3593 3567 3607
rect 3453 3573 3467 3587
rect 3493 3553 3507 3567
rect 3413 3514 3427 3528
rect 3453 3514 3467 3528
rect 3313 3472 3327 3486
rect 3372 3473 3386 3487
rect 3393 3473 3407 3487
rect 3393 3433 3407 3447
rect 3273 3393 3287 3407
rect 3433 3393 3447 3407
rect 3253 3353 3267 3367
rect 3233 3294 3247 3308
rect 3113 3233 3127 3247
rect 2953 3213 2967 3227
rect 3053 3213 3067 3227
rect 2953 3173 2967 3187
rect 2912 3093 2926 3107
rect 2933 3093 2947 3107
rect 2893 2994 2907 3008
rect 2993 3073 3007 3087
rect 2773 2933 2787 2947
rect 2813 2933 2827 2947
rect 2873 2953 2887 2967
rect 2853 2833 2867 2847
rect 2753 2774 2767 2788
rect 2813 2773 2827 2787
rect 2093 2713 2107 2727
rect 2133 2713 2147 2727
rect 2233 2713 2247 2727
rect 2293 2713 2307 2727
rect 2013 2613 2027 2627
rect 1873 2573 1887 2587
rect 2573 2653 2587 2667
rect 1733 2553 1747 2567
rect 2233 2553 2247 2567
rect 2553 2553 2567 2567
rect 1573 2513 1587 2527
rect 1773 2513 1787 2527
rect 1393 2474 1407 2488
rect 1513 2474 1527 2488
rect 1433 2373 1447 2387
rect 2153 2493 2167 2507
rect 1593 2393 1607 2407
rect 1533 2333 1547 2347
rect 1453 2293 1467 2307
rect 1613 2293 1627 2307
rect 1413 2254 1427 2268
rect 1393 2213 1407 2227
rect 1353 2173 1367 2187
rect 1473 2212 1487 2226
rect 1513 2193 1527 2207
rect 1613 2212 1627 2226
rect 1913 2474 1927 2488
rect 1953 2474 1967 2488
rect 1833 2393 1847 2407
rect 2073 2473 2087 2487
rect 2113 2474 2127 2488
rect 2513 2493 2527 2507
rect 2193 2474 2207 2488
rect 2233 2474 2247 2488
rect 2273 2474 2287 2488
rect 2353 2474 2367 2488
rect 2053 2413 2067 2427
rect 2133 2432 2147 2446
rect 2193 2433 2207 2447
rect 2073 2393 2087 2407
rect 2293 2432 2307 2446
rect 2433 2474 2447 2488
rect 2373 2413 2387 2427
rect 1913 2373 1927 2387
rect 2053 2373 2067 2387
rect 2113 2373 2127 2387
rect 2253 2373 2267 2387
rect 1953 2353 1967 2367
rect 1733 2333 1747 2347
rect 1873 2313 1887 2327
rect 1813 2293 1827 2307
rect 1693 2254 1707 2268
rect 1733 2252 1747 2266
rect 1873 2254 1887 2268
rect 1733 2213 1747 2227
rect 1793 2212 1807 2226
rect 1633 2193 1647 2207
rect 1593 2173 1607 2187
rect 1393 2133 1407 2147
rect 1153 2013 1167 2027
rect 1253 2013 1267 2027
rect 1493 2013 1507 2027
rect 1593 2013 1607 2027
rect 913 1973 927 1987
rect 953 1973 967 1987
rect 973 1954 987 1968
rect 1013 1954 1027 1968
rect 793 1912 807 1926
rect 853 1913 867 1927
rect 833 1773 847 1787
rect 593 1733 607 1747
rect 693 1734 707 1748
rect 733 1734 747 1748
rect 392 1692 406 1706
rect 413 1693 427 1707
rect 373 1593 387 1607
rect 413 1553 427 1567
rect 513 1692 527 1706
rect 593 1633 607 1647
rect 473 1533 487 1547
rect 453 1493 467 1507
rect 313 1473 327 1487
rect 273 1453 287 1467
rect 493 1513 507 1527
rect 613 1513 627 1527
rect 293 1433 307 1447
rect 333 1434 347 1448
rect 393 1433 407 1447
rect 533 1493 547 1507
rect 233 1392 247 1406
rect 173 1273 187 1287
rect 253 1273 267 1287
rect 53 1213 67 1227
rect 133 1214 147 1228
rect 173 1214 187 1228
rect 213 1214 227 1228
rect 353 1333 367 1347
rect 573 1434 587 1448
rect 673 1473 687 1487
rect 613 1433 627 1447
rect 713 1434 727 1448
rect 633 1413 647 1427
rect 393 1273 407 1287
rect 313 1233 327 1247
rect 53 1173 67 1187
rect 33 1153 47 1167
rect 93 1172 107 1186
rect 133 1173 147 1187
rect 393 1213 407 1227
rect 473 1392 487 1406
rect 533 1392 547 1406
rect 593 1392 607 1406
rect 633 1353 647 1367
rect 473 1333 487 1347
rect 493 1273 507 1287
rect 53 913 67 927
rect 93 914 107 928
rect 53 873 67 887
rect 233 1172 247 1186
rect 273 1172 287 1186
rect 213 914 227 928
rect 133 872 147 886
rect 193 872 207 886
rect 73 773 87 787
rect 113 773 127 787
rect 153 733 167 747
rect 233 733 247 747
rect 333 1172 347 1186
rect 453 1172 467 1186
rect 393 993 407 1007
rect 473 993 487 1007
rect 413 973 427 987
rect 353 933 367 947
rect 393 933 407 947
rect 453 933 467 947
rect 593 1253 607 1267
rect 553 1214 567 1228
rect 793 1734 807 1748
rect 893 1912 907 1926
rect 933 1912 947 1926
rect 953 1773 967 1787
rect 1153 1953 1167 1967
rect 1193 1954 1207 1968
rect 1353 1954 1367 1968
rect 1473 1954 1487 1968
rect 1033 1912 1047 1926
rect 1073 1912 1087 1926
rect 1133 1793 1147 1807
rect 1093 1773 1107 1787
rect 1293 1813 1307 1827
rect 773 1693 787 1707
rect 773 1533 787 1547
rect 933 1692 947 1706
rect 1033 1734 1047 1748
rect 1093 1734 1107 1748
rect 1133 1734 1147 1748
rect 1233 1773 1247 1787
rect 993 1673 1007 1687
rect 1073 1693 1087 1707
rect 1053 1653 1067 1667
rect 973 1573 987 1587
rect 1053 1573 1067 1587
rect 813 1513 827 1527
rect 933 1513 947 1527
rect 773 1473 787 1487
rect 813 1453 827 1467
rect 873 1453 887 1467
rect 773 1433 787 1447
rect 793 1392 807 1406
rect 833 1353 847 1367
rect 833 1313 847 1327
rect 753 1293 767 1307
rect 813 1293 827 1307
rect 933 1434 947 1448
rect 913 1353 927 1367
rect 573 1172 587 1186
rect 633 973 647 987
rect 533 953 547 967
rect 593 953 607 967
rect 493 933 507 947
rect 533 914 547 928
rect 433 893 447 907
rect 373 872 387 886
rect 453 872 467 886
rect 513 872 527 886
rect 553 872 567 886
rect 533 853 547 867
rect 313 833 327 847
rect 413 833 427 847
rect 293 713 307 727
rect 393 713 407 727
rect 193 694 207 708
rect 233 694 247 708
rect 93 652 107 666
rect 153 652 167 666
rect 213 652 227 666
rect 253 613 267 627
rect 353 652 367 666
rect 33 553 47 567
rect 293 553 307 567
rect 213 453 227 467
rect 113 394 127 408
rect 253 394 267 408
rect 193 352 207 366
rect 193 253 207 267
rect 33 174 47 188
rect 93 174 107 188
rect 353 433 367 447
rect 793 1172 807 1186
rect 733 1153 747 1167
rect 733 1093 747 1107
rect 713 973 727 987
rect 793 973 807 987
rect 693 933 707 947
rect 673 914 687 928
rect 753 933 767 947
rect 653 872 667 886
rect 593 773 607 787
rect 653 773 667 787
rect 533 733 547 747
rect 473 694 487 708
rect 513 693 527 707
rect 593 694 607 708
rect 573 652 587 666
rect 513 613 527 627
rect 573 573 587 587
rect 413 453 427 467
rect 413 432 427 446
rect 553 433 567 447
rect 393 394 407 408
rect 473 394 487 408
rect 593 413 607 427
rect 633 393 647 407
rect 153 132 167 146
rect 253 132 267 146
rect 413 352 427 366
rect 453 352 467 366
rect 573 352 587 366
rect 633 333 647 347
rect 393 313 407 327
rect 353 213 367 227
rect 333 193 347 207
rect 313 174 327 188
rect 693 733 707 747
rect 833 914 847 928
rect 833 873 847 887
rect 773 753 787 767
rect 713 713 727 727
rect 753 713 767 727
rect 833 773 847 787
rect 993 1433 1007 1447
rect 1053 1434 1067 1448
rect 1113 1693 1127 1707
rect 1193 1692 1207 1706
rect 1293 1692 1307 1706
rect 1353 1692 1367 1706
rect 1233 1633 1247 1647
rect 1313 1633 1327 1647
rect 1193 1513 1207 1527
rect 1113 1493 1127 1507
rect 1113 1434 1127 1448
rect 1153 1434 1167 1448
rect 1653 2013 1667 2027
rect 1733 2013 1747 2027
rect 1533 1954 1547 1968
rect 1593 1954 1607 1968
rect 1633 1954 1647 1968
rect 1593 1873 1607 1887
rect 1593 1793 1607 1807
rect 1713 1973 1727 1987
rect 1753 1973 1767 1987
rect 1833 2133 1847 2147
rect 2093 2293 2107 2307
rect 2293 2293 2307 2307
rect 2113 2254 2127 2268
rect 2173 2254 2187 2268
rect 2233 2254 2247 2268
rect 2333 2254 2347 2268
rect 1993 2212 2007 2226
rect 2092 2212 2106 2226
rect 2113 2213 2127 2227
rect 2153 2212 2167 2226
rect 2193 2193 2207 2207
rect 2053 2173 2067 2187
rect 2093 2173 2107 2187
rect 1953 2073 1967 2087
rect 1973 1973 1987 1987
rect 1793 1933 1807 1947
rect 1733 1912 1747 1926
rect 1693 1873 1707 1887
rect 1793 1873 1807 1887
rect 1493 1732 1507 1746
rect 1553 1734 1567 1748
rect 1493 1693 1507 1707
rect 1573 1673 1587 1687
rect 1713 1793 1727 1807
rect 1773 1793 1787 1807
rect 1813 1793 1827 1807
rect 1653 1773 1667 1787
rect 1533 1653 1547 1667
rect 1633 1653 1647 1667
rect 1353 1613 1367 1627
rect 1473 1613 1487 1627
rect 1253 1493 1267 1507
rect 973 1333 987 1347
rect 913 1253 927 1267
rect 913 1214 927 1228
rect 1233 1433 1247 1447
rect 1033 1392 1047 1406
rect 1073 1392 1087 1406
rect 1113 1393 1127 1407
rect 1173 1392 1187 1406
rect 1113 1253 1127 1267
rect 1013 1214 1027 1228
rect 1193 1233 1207 1247
rect 1233 1233 1247 1247
rect 1153 1214 1167 1228
rect 973 1172 987 1186
rect 1133 1172 1147 1186
rect 1173 1172 1187 1186
rect 1273 1473 1287 1487
rect 1313 1434 1327 1448
rect 1573 1513 1587 1527
rect 1473 1473 1487 1487
rect 1393 1434 1407 1448
rect 1433 1434 1447 1448
rect 1273 1393 1287 1407
rect 1273 1353 1287 1367
rect 1333 1392 1347 1406
rect 1393 1393 1407 1407
rect 1753 1734 1767 1748
rect 1833 1773 1847 1787
rect 1773 1692 1787 1706
rect 1813 1692 1827 1706
rect 1853 1692 1867 1706
rect 2033 1954 2047 1968
rect 2273 2212 2287 2226
rect 2313 2193 2327 2207
rect 2453 2432 2467 2446
rect 2453 2373 2467 2387
rect 2573 2493 2587 2507
rect 2553 2273 2567 2287
rect 2493 2254 2507 2268
rect 2413 2212 2427 2226
rect 2393 2193 2407 2207
rect 2153 2073 2167 2087
rect 2233 2073 2247 2087
rect 2153 2033 2167 2047
rect 1993 1933 2007 1947
rect 1973 1873 1987 1887
rect 2013 1913 2027 1927
rect 2173 1953 2187 1967
rect 2233 1954 2247 1968
rect 2313 1954 2327 1968
rect 2353 1954 2367 1968
rect 1993 1853 2007 1867
rect 1993 1793 2007 1807
rect 1913 1733 1927 1747
rect 1933 1734 1947 1748
rect 1953 1692 1967 1706
rect 1893 1653 1907 1667
rect 2153 1912 2167 1926
rect 2033 1853 2047 1867
rect 2013 1773 2027 1787
rect 2193 1912 2207 1926
rect 2333 1873 2347 1887
rect 2173 1853 2187 1867
rect 2253 1853 2267 1867
rect 2153 1793 2167 1807
rect 2073 1773 2087 1787
rect 2133 1733 2147 1747
rect 2193 1734 2207 1748
rect 2053 1692 2067 1706
rect 2093 1692 2107 1706
rect 2133 1692 2147 1706
rect 1993 1553 2007 1567
rect 2073 1513 2087 1527
rect 1733 1473 1747 1487
rect 2013 1473 2027 1487
rect 1893 1434 1907 1448
rect 1313 1353 1327 1367
rect 1293 1333 1307 1347
rect 1293 1253 1307 1267
rect 1253 1213 1267 1227
rect 1333 1333 1347 1347
rect 1313 1233 1327 1247
rect 1553 1353 1567 1367
rect 1493 1313 1507 1327
rect 1533 1313 1547 1327
rect 1473 1273 1487 1287
rect 1393 1253 1407 1267
rect 1453 1253 1467 1267
rect 1433 1214 1447 1228
rect 1273 1172 1287 1186
rect 1313 1172 1327 1186
rect 1393 1172 1407 1186
rect 1453 1172 1467 1186
rect 1033 1133 1047 1147
rect 1233 1133 1247 1147
rect 1353 1133 1367 1147
rect 1353 1093 1367 1107
rect 1473 993 1487 1007
rect 1053 933 1067 947
rect 1333 933 1347 947
rect 1413 933 1427 947
rect 873 913 887 927
rect 913 914 927 928
rect 953 914 967 928
rect 993 914 1007 928
rect 1173 914 1187 928
rect 1213 913 1227 927
rect 1273 914 1287 928
rect 873 853 887 867
rect 993 873 1007 887
rect 933 833 947 847
rect 873 773 887 787
rect 853 753 867 767
rect 853 713 867 727
rect 713 493 727 507
rect 733 413 747 427
rect 753 394 767 408
rect 793 394 807 408
rect 1073 872 1087 886
rect 1033 853 1047 867
rect 1013 833 1027 847
rect 1053 833 1067 847
rect 1153 833 1167 847
rect 1253 872 1267 886
rect 1373 914 1387 928
rect 1353 873 1367 887
rect 1553 1273 1567 1287
rect 1573 1253 1587 1267
rect 1553 1233 1567 1247
rect 1593 1214 1607 1228
rect 1653 1392 1667 1406
rect 1713 1392 1727 1406
rect 1773 1353 1787 1367
rect 1993 1293 2007 1307
rect 1753 1253 1767 1267
rect 1993 1253 2007 1267
rect 1633 1213 1647 1227
rect 1573 1172 1587 1186
rect 1533 933 1547 947
rect 1353 833 1367 847
rect 1433 872 1447 886
rect 1473 872 1487 886
rect 1553 872 1567 886
rect 1493 833 1507 847
rect 1273 773 1287 787
rect 1393 773 1407 787
rect 1213 753 1227 767
rect 993 693 1007 707
rect 1213 694 1227 708
rect 1253 673 1267 687
rect 873 652 887 666
rect 913 652 927 666
rect 1013 653 1027 667
rect 973 553 987 567
rect 933 453 947 467
rect 893 413 907 427
rect 693 352 707 366
rect 1113 593 1127 607
rect 1033 553 1047 567
rect 1313 753 1327 767
rect 1373 694 1387 708
rect 1413 694 1427 708
rect 1453 694 1467 708
rect 1273 633 1287 647
rect 1473 652 1487 666
rect 1433 633 1447 647
rect 1352 593 1366 607
rect 1373 593 1387 607
rect 1333 553 1347 567
rect 1253 513 1267 527
rect 1013 433 1027 447
rect 1093 433 1107 447
rect 953 413 967 427
rect 833 333 847 347
rect 1073 394 1087 408
rect 873 313 887 327
rect 653 293 667 307
rect 733 293 747 307
rect 893 273 907 287
rect 953 333 967 347
rect 1013 313 1027 327
rect 433 253 447 267
rect 573 213 587 227
rect 613 213 627 227
rect 473 174 487 188
rect 513 173 527 187
rect 693 174 707 188
rect 993 233 1007 247
rect 933 174 947 188
rect 333 132 347 146
rect 393 133 407 147
rect 453 132 467 146
rect 513 132 527 146
rect 553 132 567 146
rect 693 133 707 147
rect 1113 413 1127 427
rect 1173 394 1187 408
rect 1253 393 1267 407
rect 1113 313 1127 327
rect 1193 352 1207 366
rect 1233 352 1247 366
rect 1273 352 1287 366
rect 1253 333 1267 347
rect 1633 1173 1647 1187
rect 1773 1214 1787 1228
rect 1833 1214 1847 1228
rect 1613 1093 1627 1107
rect 1713 1172 1727 1186
rect 1753 1172 1767 1186
rect 1653 1133 1667 1147
rect 1953 1172 1967 1186
rect 1993 1172 2007 1186
rect 1773 1093 1787 1107
rect 1893 1093 1907 1107
rect 1873 1013 1887 1027
rect 1633 993 1647 1007
rect 1673 953 1687 967
rect 1813 953 1827 967
rect 1773 914 1787 928
rect 1813 914 1827 928
rect 1593 893 1607 907
rect 2113 1434 2127 1448
rect 2093 1392 2107 1406
rect 2133 1373 2147 1387
rect 2053 1293 2067 1307
rect 2133 1293 2147 1307
rect 2113 1273 2127 1287
rect 2073 1214 2087 1228
rect 2173 1553 2187 1567
rect 2233 1434 2247 1448
rect 2453 2193 2467 2207
rect 2453 1993 2467 2007
rect 2413 1954 2427 1968
rect 2433 1912 2447 1926
rect 2313 1813 2327 1827
rect 2393 1813 2407 1827
rect 2373 1793 2387 1807
rect 2273 1653 2287 1667
rect 2253 1373 2267 1387
rect 2333 1633 2347 1647
rect 2513 1912 2527 1926
rect 2613 2474 2627 2488
rect 2653 2474 2667 2488
rect 2713 2474 2727 2488
rect 2773 2474 2787 2488
rect 2713 2413 2727 2427
rect 2673 2353 2687 2367
rect 2593 2333 2607 2347
rect 2633 2333 2647 2347
rect 2593 2253 2607 2267
rect 2833 2732 2847 2746
rect 2873 2733 2887 2747
rect 2833 2693 2847 2707
rect 3013 3033 3027 3047
rect 3073 2952 3087 2966
rect 3013 2933 3027 2947
rect 3133 3093 3147 3107
rect 3113 2873 3127 2887
rect 3233 3253 3247 3267
rect 3373 3333 3387 3347
rect 3453 3333 3467 3347
rect 3313 3294 3327 3308
rect 3353 3293 3367 3307
rect 3273 3253 3287 3267
rect 3173 3213 3187 3227
rect 3253 3213 3267 3227
rect 3333 3252 3347 3266
rect 3273 3193 3287 3207
rect 3193 3153 3207 3167
rect 3153 3073 3167 3087
rect 3233 2994 3247 3008
rect 3133 2833 3147 2847
rect 3073 2774 3087 2788
rect 3413 3294 3427 3308
rect 3752 4253 3766 4267
rect 3773 4253 3787 4267
rect 3753 4153 3767 4167
rect 3733 4073 3747 4087
rect 3673 4053 3687 4067
rect 3713 4034 3727 4048
rect 3753 4034 3767 4048
rect 3793 4173 3807 4187
rect 3693 3973 3707 3987
rect 3653 3953 3667 3967
rect 3653 3913 3667 3927
rect 3633 3873 3647 3887
rect 3713 3853 3727 3867
rect 3633 3753 3647 3767
rect 3633 3673 3647 3687
rect 3593 3553 3607 3567
rect 3593 3514 3607 3528
rect 3573 3453 3587 3467
rect 3673 3633 3687 3647
rect 3693 3613 3707 3627
rect 3673 3553 3687 3567
rect 3713 3553 3727 3567
rect 3953 4453 3967 4467
rect 3913 4353 3927 4367
rect 3853 4334 3867 4348
rect 3893 4334 3907 4348
rect 3873 4273 3887 4287
rect 3833 4253 3847 4267
rect 3833 4193 3847 4207
rect 3933 4293 3947 4307
rect 3933 4193 3947 4207
rect 3853 4153 3867 4167
rect 3873 4133 3887 4147
rect 3853 4093 3867 4107
rect 3833 4073 3847 4087
rect 3813 4053 3827 4067
rect 3913 4153 3927 4167
rect 4013 4512 4027 4526
rect 4053 4513 4067 4527
rect 4013 4473 4027 4487
rect 4033 4453 4047 4467
rect 4273 4812 4287 4826
rect 4313 4813 4327 4827
rect 4353 4853 4367 4867
rect 4613 5353 4627 5367
rect 4533 5293 4547 5307
rect 4613 5253 4627 5267
rect 4613 5213 4627 5227
rect 4533 5193 4547 5207
rect 4593 5193 4607 5207
rect 4613 5173 4627 5187
rect 4573 5113 4587 5127
rect 4533 5074 4547 5088
rect 4553 5032 4567 5046
rect 4573 4993 4587 5007
rect 4853 5413 4867 5427
rect 4773 5373 4787 5387
rect 4813 5374 4827 5388
rect 4673 5293 4687 5307
rect 5173 5393 5187 5407
rect 5353 5393 5367 5407
rect 4833 5173 4847 5187
rect 4793 5133 4807 5147
rect 4713 5032 4727 5046
rect 4653 4993 4667 5007
rect 4553 4973 4567 4987
rect 4513 4953 4527 4967
rect 4833 5074 4847 5088
rect 4873 5313 4887 5327
rect 4913 5313 4927 5327
rect 5053 5373 5067 5387
rect 5113 5374 5127 5388
rect 4953 5353 4967 5367
rect 5013 5332 5027 5346
rect 4993 5293 5007 5307
rect 4953 5273 4967 5287
rect 5013 5253 5027 5267
rect 4993 5193 5007 5207
rect 4853 5053 4867 5067
rect 4793 5032 4807 5046
rect 4773 4953 4787 4967
rect 4573 4913 4587 4927
rect 4753 4913 4767 4927
rect 4553 4893 4567 4907
rect 4233 4773 4247 4787
rect 4233 4713 4247 4727
rect 4213 4653 4227 4667
rect 4193 4613 4207 4627
rect 4213 4554 4227 4568
rect 4093 4533 4107 4547
rect 4073 4453 4087 4467
rect 4173 4473 4187 4487
rect 4213 4453 4227 4467
rect 4093 4373 4107 4387
rect 4133 4373 4147 4387
rect 3973 4273 3987 4287
rect 3993 4253 4007 4267
rect 3993 4213 4007 4227
rect 3973 4093 3987 4107
rect 4073 4293 4087 4307
rect 4073 4253 4087 4267
rect 4073 4193 4087 4207
rect 4153 4353 4167 4367
rect 4153 4273 4167 4287
rect 4113 4253 4127 4267
rect 4093 4173 4107 4187
rect 4133 4173 4147 4187
rect 4053 4153 4067 4167
rect 4073 4113 4087 4127
rect 4133 4113 4147 4127
rect 4072 4073 4086 4087
rect 4093 4073 4107 4087
rect 4013 4034 4027 4048
rect 4053 4034 4067 4048
rect 3813 3953 3827 3967
rect 3753 3933 3767 3947
rect 3793 3913 3807 3927
rect 3793 3833 3807 3847
rect 3813 3814 3827 3828
rect 3873 3992 3887 4006
rect 3913 3992 3927 4006
rect 3953 3992 3967 4006
rect 3873 3953 3887 3967
rect 4073 3992 4087 4006
rect 4113 3992 4127 4006
rect 4013 3953 4027 3967
rect 4073 3953 4087 3967
rect 4133 3953 4147 3967
rect 3993 3913 4007 3927
rect 3873 3873 3887 3887
rect 3893 3853 3907 3867
rect 3873 3813 3887 3827
rect 3773 3773 3787 3787
rect 3833 3772 3847 3786
rect 3793 3593 3807 3607
rect 3773 3513 3787 3527
rect 3693 3472 3707 3486
rect 3733 3472 3747 3486
rect 3633 3453 3647 3467
rect 3673 3433 3687 3447
rect 3613 3393 3627 3407
rect 3553 3353 3567 3367
rect 3492 3293 3506 3307
rect 3513 3293 3527 3307
rect 3593 3333 3607 3347
rect 3653 3333 3667 3347
rect 3433 3252 3447 3266
rect 3393 3233 3407 3247
rect 3352 3133 3366 3147
rect 3373 3133 3387 3147
rect 3333 3093 3347 3107
rect 3393 3113 3407 3127
rect 3413 3093 3427 3107
rect 3313 3013 3327 3027
rect 3333 2952 3347 2966
rect 3273 2933 3287 2947
rect 3213 2913 3227 2927
rect 3373 2913 3387 2927
rect 3353 2813 3367 2827
rect 3193 2774 3207 2788
rect 3173 2733 3187 2747
rect 3233 2732 3247 2746
rect 2953 2653 2967 2667
rect 2993 2653 3007 2667
rect 3153 2613 3167 2627
rect 3273 2693 3287 2707
rect 3253 2593 3267 2607
rect 2933 2513 2947 2527
rect 3153 2513 3167 2527
rect 2833 2474 2847 2488
rect 3033 2474 3047 2488
rect 3073 2474 3087 2488
rect 3113 2474 3127 2488
rect 3193 2474 3207 2488
rect 2953 2453 2967 2467
rect 2893 2432 2907 2446
rect 2933 2432 2947 2446
rect 2833 2393 2847 2407
rect 2753 2293 2767 2307
rect 2813 2293 2827 2307
rect 2733 2253 2747 2267
rect 2613 2212 2627 2226
rect 2673 2212 2687 2226
rect 2713 2212 2727 2226
rect 2733 2113 2747 2127
rect 2733 2073 2747 2087
rect 2633 1954 2647 1968
rect 2693 1954 2707 1968
rect 2473 1873 2487 1887
rect 2453 1753 2467 1767
rect 2473 1733 2487 1747
rect 2453 1692 2467 1706
rect 2493 1692 2507 1706
rect 2553 1673 2567 1687
rect 2573 1673 2587 1687
rect 2453 1633 2467 1647
rect 2353 1533 2367 1547
rect 2433 1533 2447 1547
rect 2293 1433 2307 1447
rect 2313 1434 2327 1448
rect 2333 1392 2347 1406
rect 2513 1434 2527 1448
rect 2613 1813 2627 1827
rect 2593 1533 2607 1547
rect 2593 1393 2607 1407
rect 2393 1373 2407 1387
rect 2453 1373 2467 1387
rect 2193 1313 2207 1327
rect 2193 1273 2207 1287
rect 2173 1253 2187 1267
rect 2213 1233 2227 1247
rect 2173 1214 2187 1228
rect 2233 1213 2247 1227
rect 2193 1172 2207 1186
rect 2133 1113 2147 1127
rect 2113 1093 2127 1107
rect 2093 1053 2107 1067
rect 1973 993 1987 1007
rect 2013 993 2027 1007
rect 1933 914 1947 928
rect 1633 853 1647 867
rect 1593 833 1607 847
rect 1533 813 1547 827
rect 1573 813 1587 827
rect 1613 773 1627 787
rect 1533 733 1547 747
rect 1573 733 1587 747
rect 1413 413 1427 427
rect 1513 413 1527 427
rect 1633 693 1647 707
rect 1693 872 1707 886
rect 1693 773 1707 787
rect 1753 753 1767 767
rect 1833 872 1847 886
rect 1873 872 1887 886
rect 1913 872 1927 886
rect 1913 793 1927 807
rect 1673 733 1687 747
rect 1653 652 1667 666
rect 1593 613 1607 627
rect 1573 593 1587 607
rect 1553 573 1567 587
rect 1553 533 1567 547
rect 1693 652 1707 666
rect 1793 593 1807 607
rect 1673 553 1687 567
rect 1813 553 1827 567
rect 1793 533 1807 547
rect 1813 513 1827 527
rect 1713 493 1727 507
rect 1573 473 1587 487
rect 1453 394 1467 408
rect 1493 394 1507 408
rect 1533 394 1547 408
rect 1653 394 1667 408
rect 1393 352 1407 366
rect 1493 353 1507 367
rect 1553 352 1567 366
rect 1733 413 1747 427
rect 1773 413 1787 427
rect 1353 313 1367 327
rect 1433 313 1447 327
rect 1153 293 1167 307
rect 1253 293 1267 307
rect 1313 293 1327 307
rect 1453 253 1467 267
rect 1553 233 1567 247
rect 1613 233 1627 247
rect 1453 193 1467 207
rect 1033 174 1047 188
rect 1093 174 1107 188
rect 1353 174 1367 188
rect 1413 174 1427 188
rect 1493 173 1507 187
rect 733 132 747 146
rect 553 93 567 107
rect 953 132 967 146
rect 993 132 1007 146
rect 1213 132 1227 146
rect 1053 113 1067 127
rect 913 93 927 107
rect 1353 133 1367 147
rect 1433 93 1447 107
rect 1913 753 1927 767
rect 1853 693 1867 707
rect 1893 694 1907 708
rect 1933 733 1947 747
rect 1873 652 1887 666
rect 1893 633 1907 647
rect 1893 593 1907 607
rect 2013 972 2027 986
rect 2053 914 2067 928
rect 2013 793 2027 807
rect 1973 694 1987 708
rect 2273 1273 2287 1287
rect 2253 1053 2267 1067
rect 2173 914 2187 928
rect 2353 1233 2367 1247
rect 2313 1214 2327 1228
rect 2533 1313 2547 1327
rect 2413 1233 2427 1247
rect 2393 1213 2407 1227
rect 2333 1172 2347 1186
rect 2473 1214 2487 1228
rect 2393 1093 2407 1107
rect 2373 993 2387 1007
rect 2333 933 2347 947
rect 2293 914 2307 928
rect 2393 914 2407 928
rect 2413 873 2427 887
rect 2213 833 2227 847
rect 2272 833 2286 847
rect 2293 833 2307 847
rect 2153 813 2167 827
rect 2093 733 2107 747
rect 2293 733 2307 747
rect 2393 733 2407 747
rect 2093 694 2107 708
rect 2133 694 2147 708
rect 1953 653 1967 667
rect 1933 513 1947 527
rect 1913 493 1927 507
rect 1913 433 1927 447
rect 1833 413 1847 427
rect 1893 413 1907 427
rect 1833 352 1847 366
rect 1833 293 1847 307
rect 1853 273 1867 287
rect 1873 253 1887 267
rect 1733 193 1747 207
rect 1673 174 1687 188
rect 1653 132 1667 146
rect 1533 113 1547 127
rect 1733 132 1747 146
rect 1693 93 1707 107
rect 1393 73 1407 87
rect 1493 73 1507 87
rect 1873 132 1887 146
rect 2052 653 2066 667
rect 2073 653 2087 667
rect 2313 693 2327 707
rect 2372 694 2386 708
rect 2393 693 2407 707
rect 2013 593 2027 607
rect 1972 433 1986 447
rect 1993 433 2007 447
rect 1973 352 1987 366
rect 1913 313 1927 327
rect 2153 652 2167 666
rect 2293 652 2307 666
rect 2273 613 2287 627
rect 2313 613 2327 627
rect 2453 1172 2467 1186
rect 2693 1773 2707 1787
rect 2733 1773 2747 1787
rect 2653 1753 2667 1767
rect 2633 1693 2647 1707
rect 2613 1313 2627 1327
rect 2713 1692 2727 1706
rect 2673 1653 2687 1667
rect 2653 1613 2667 1627
rect 2633 1233 2647 1247
rect 2733 1593 2747 1607
rect 2673 1392 2687 1406
rect 2793 2254 2807 2268
rect 2913 2212 2927 2226
rect 2853 2193 2867 2207
rect 2973 2432 2987 2446
rect 3013 2432 3027 2446
rect 3353 2573 3367 2587
rect 3493 3053 3507 3067
rect 3413 2993 3427 3007
rect 3493 2994 3507 3008
rect 3573 3252 3587 3266
rect 3613 3213 3627 3227
rect 3553 3193 3567 3207
rect 3533 3013 3547 3027
rect 3433 2952 3447 2966
rect 3473 2873 3487 2887
rect 3393 2833 3407 2847
rect 3453 2774 3467 2788
rect 3493 2774 3507 2788
rect 3453 2653 3467 2667
rect 3393 2573 3407 2587
rect 3373 2553 3387 2567
rect 3313 2474 3327 2488
rect 3353 2474 3367 2488
rect 3493 2593 3507 2607
rect 3633 3193 3647 3207
rect 3613 3153 3627 3167
rect 3573 3093 3587 3107
rect 3553 2994 3567 3008
rect 3693 3373 3707 3387
rect 3673 3293 3687 3307
rect 3713 3294 3727 3308
rect 3773 3473 3787 3487
rect 3993 3853 4007 3867
rect 4053 3833 4067 3847
rect 4033 3814 4047 3828
rect 3913 3772 3927 3786
rect 4033 3693 4047 3707
rect 4273 4554 4287 4568
rect 4333 4812 4347 4826
rect 4473 4854 4487 4868
rect 4513 4854 4527 4868
rect 4553 4853 4567 4867
rect 4433 4793 4447 4807
rect 4513 4793 4527 4807
rect 4413 4773 4427 4787
rect 4493 4773 4507 4787
rect 4373 4713 4387 4727
rect 4373 4673 4387 4687
rect 4473 4733 4487 4747
rect 4433 4713 4447 4727
rect 4393 4593 4407 4607
rect 4493 4673 4507 4687
rect 4473 4573 4487 4587
rect 4493 4553 4507 4567
rect 4333 4512 4347 4526
rect 4373 4513 4387 4527
rect 4473 4512 4487 4526
rect 4293 4413 4307 4427
rect 4373 4393 4387 4407
rect 4473 4433 4487 4447
rect 4453 4393 4467 4407
rect 4413 4353 4427 4367
rect 4473 4353 4487 4367
rect 4293 4334 4307 4348
rect 4353 4333 4367 4347
rect 4553 4813 4567 4827
rect 4553 4773 4567 4787
rect 4593 4893 4607 4907
rect 4613 4854 4627 4868
rect 4653 4854 4667 4868
rect 4713 4853 4727 4867
rect 4913 5074 4927 5088
rect 4953 5074 4967 5088
rect 5013 5153 5027 5167
rect 5133 5332 5147 5346
rect 5093 5293 5107 5307
rect 5113 5113 5127 5127
rect 5213 5374 5227 5388
rect 5253 5374 5267 5388
rect 5313 5374 5327 5388
rect 5393 5374 5407 5388
rect 5513 5374 5527 5388
rect 5553 5374 5567 5388
rect 5033 5093 5047 5107
rect 5073 5093 5087 5107
rect 5013 5073 5027 5087
rect 4973 5032 4987 5046
rect 4933 5013 4947 5027
rect 4873 4933 4887 4947
rect 4833 4873 4847 4887
rect 4593 4813 4607 4827
rect 4573 4633 4587 4647
rect 4673 4753 4687 4767
rect 4673 4732 4687 4746
rect 4633 4693 4647 4707
rect 4553 4613 4567 4627
rect 4593 4613 4607 4627
rect 4613 4573 4627 4587
rect 4653 4593 4667 4607
rect 4533 4553 4547 4567
rect 4553 4553 4567 4567
rect 4633 4553 4647 4567
rect 4852 4853 4866 4867
rect 4873 4854 4887 4868
rect 4753 4812 4767 4826
rect 4713 4713 4727 4727
rect 4713 4633 4727 4647
rect 4733 4593 4747 4607
rect 4513 4513 4527 4527
rect 4513 4413 4527 4427
rect 4454 4333 4468 4347
rect 4493 4333 4507 4347
rect 4253 4293 4267 4307
rect 4233 4273 4247 4287
rect 4233 4193 4247 4207
rect 4233 4133 4247 4147
rect 4173 4093 4187 4107
rect 4233 4093 4247 4107
rect 4233 4053 4247 4067
rect 4313 4273 4327 4287
rect 4273 4253 4287 4267
rect 4333 4253 4347 4267
rect 4253 4033 4267 4047
rect 4173 3993 4187 4007
rect 4153 3833 4167 3847
rect 4133 3814 4147 3828
rect 4253 3993 4267 4007
rect 4213 3953 4227 3967
rect 4193 3913 4207 3927
rect 4193 3873 4207 3887
rect 4193 3813 4207 3827
rect 4073 3772 4087 3786
rect 4113 3772 4127 3786
rect 4153 3772 4167 3786
rect 4093 3733 4107 3747
rect 4053 3653 4067 3667
rect 4033 3613 4047 3627
rect 3893 3593 3907 3607
rect 4013 3573 4027 3587
rect 3833 3514 3847 3528
rect 3973 3513 3987 3527
rect 3793 3453 3807 3467
rect 3833 3453 3847 3467
rect 3793 3373 3807 3387
rect 3893 3433 3907 3447
rect 3953 3413 3967 3427
rect 3993 3413 4007 3427
rect 3993 3373 4007 3387
rect 4013 3333 4027 3347
rect 4053 3373 4067 3387
rect 3773 3293 3787 3307
rect 3893 3293 3907 3307
rect 3953 3294 3967 3308
rect 4033 3313 4047 3327
rect 3733 3252 3747 3266
rect 3693 3093 3707 3107
rect 3653 3053 3667 3067
rect 3653 3032 3667 3046
rect 3593 2952 3607 2966
rect 3633 2833 3647 2847
rect 3533 2773 3547 2787
rect 3573 2774 3587 2788
rect 3613 2774 3627 2788
rect 3733 3033 3747 3047
rect 3773 3193 3787 3207
rect 3793 3173 3807 3187
rect 3773 3033 3787 3047
rect 3693 2994 3707 3008
rect 3713 2893 3727 2907
rect 3653 2793 3667 2807
rect 3633 2733 3647 2747
rect 3593 2653 3607 2667
rect 3673 2773 3687 2787
rect 3713 2793 3727 2807
rect 3893 3252 3907 3266
rect 3853 3173 3867 3187
rect 3953 3233 3967 3247
rect 3933 3153 3947 3167
rect 3853 3093 3867 3107
rect 3913 3053 3927 3067
rect 3833 3033 3847 3047
rect 3793 3013 3807 3027
rect 3873 3013 3887 3027
rect 3833 2994 3847 3008
rect 3813 2913 3827 2927
rect 3853 2833 3867 2847
rect 4033 3253 4047 3267
rect 4013 3193 4027 3207
rect 4172 3733 4186 3747
rect 4193 3733 4207 3747
rect 4153 3633 4167 3647
rect 4233 3853 4247 3867
rect 4393 4292 4407 4306
rect 4332 4213 4346 4227
rect 4353 4213 4367 4227
rect 4473 4292 4487 4306
rect 4493 4213 4507 4227
rect 4313 4133 4327 4147
rect 4393 4133 4407 4147
rect 4433 4133 4447 4147
rect 4293 4053 4307 4067
rect 4273 3953 4287 3967
rect 4553 4493 4567 4507
rect 4533 4393 4547 4407
rect 4653 4513 4667 4527
rect 4832 4812 4846 4826
rect 4853 4813 4867 4827
rect 4793 4693 4807 4707
rect 4833 4633 4847 4647
rect 4773 4593 4787 4607
rect 4753 4553 4767 4567
rect 4633 4493 4647 4507
rect 4693 4512 4707 4526
rect 4733 4512 4747 4526
rect 4813 4512 4827 4526
rect 4753 4473 4767 4487
rect 4633 4453 4647 4467
rect 4593 4433 4607 4447
rect 4573 4393 4587 4407
rect 4553 4353 4567 4367
rect 4593 4353 4607 4367
rect 4513 4193 4527 4207
rect 4513 4172 4527 4186
rect 4493 4113 4507 4127
rect 4393 4092 4407 4106
rect 4373 4034 4387 4048
rect 4413 4073 4427 4087
rect 4353 3992 4367 4006
rect 4393 3992 4407 4006
rect 4293 3933 4307 3947
rect 4353 3853 4367 3867
rect 4253 3814 4267 3828
rect 4333 3813 4347 3827
rect 4233 3772 4247 3786
rect 4293 3772 4307 3786
rect 4293 3693 4307 3707
rect 4313 3653 4327 3667
rect 4313 3613 4327 3627
rect 4233 3593 4247 3607
rect 4113 3553 4127 3567
rect 4153 3553 4167 3567
rect 4193 3553 4207 3567
rect 4293 3553 4307 3567
rect 4173 3433 4187 3447
rect 4213 3433 4227 3447
rect 4193 3413 4207 3427
rect 4113 3333 4127 3347
rect 4173 3333 4187 3347
rect 4153 3313 4167 3327
rect 4073 3293 4087 3307
rect 4113 3294 4127 3308
rect 4173 3293 4187 3307
rect 4093 3252 4107 3266
rect 4093 3213 4107 3227
rect 4053 3153 4067 3167
rect 3993 3113 4007 3127
rect 4033 3113 4047 3127
rect 4013 3013 4027 3027
rect 3993 2993 4007 3007
rect 3933 2952 3947 2966
rect 4033 2993 4047 3007
rect 4173 3253 4187 3267
rect 4173 3173 4187 3187
rect 4153 3153 4167 3167
rect 4133 3113 4147 3127
rect 4113 3013 4127 3027
rect 4073 2952 4087 2966
rect 4113 2933 4127 2947
rect 4133 2952 4147 2966
rect 4513 4053 4527 4067
rect 4453 4034 4467 4048
rect 4493 4034 4507 4048
rect 4413 3833 4427 3847
rect 4473 3933 4487 3947
rect 4613 4293 4627 4307
rect 4593 4273 4607 4287
rect 4553 4253 4567 4267
rect 4593 4233 4607 4247
rect 4553 4193 4567 4207
rect 4573 4173 4587 4187
rect 4653 4353 4667 4367
rect 4713 4334 4727 4348
rect 4653 4293 4667 4307
rect 4773 4453 4787 4467
rect 4633 4233 4647 4247
rect 4713 4253 4727 4267
rect 4693 4233 4707 4247
rect 4673 4193 4687 4207
rect 4633 4133 4647 4147
rect 4613 3993 4627 4007
rect 4573 3973 4587 3987
rect 4453 3813 4467 3827
rect 4393 3772 4407 3786
rect 4353 3693 4367 3707
rect 4373 3673 4387 3687
rect 4353 3633 4367 3647
rect 4333 3513 4347 3527
rect 4273 3472 4287 3486
rect 4313 3433 4327 3447
rect 4233 3373 4247 3387
rect 4653 4113 4667 4127
rect 4673 4093 4687 4107
rect 4653 4034 4667 4048
rect 4733 4213 4747 4227
rect 4713 4173 4727 4187
rect 4693 4073 4707 4087
rect 4753 4153 4767 4167
rect 4733 4053 4747 4067
rect 4753 4033 4767 4047
rect 4633 3973 4647 3987
rect 4613 3913 4627 3927
rect 4633 3833 4647 3847
rect 4473 3733 4487 3747
rect 4473 3693 4487 3707
rect 4433 3613 4447 3627
rect 4373 3513 4387 3527
rect 4413 3514 4427 3528
rect 4453 3513 4467 3527
rect 4393 3472 4407 3486
rect 4533 3753 4547 3767
rect 4593 3772 4607 3786
rect 4553 3733 4567 3747
rect 4533 3633 4547 3647
rect 4513 3593 4527 3607
rect 4513 3472 4527 3486
rect 4613 3673 4627 3687
rect 4733 3992 4747 4006
rect 4693 3873 4707 3887
rect 4713 3853 4727 3867
rect 4673 3833 4687 3847
rect 4693 3733 4707 3747
rect 4873 4773 4887 4787
rect 4873 4733 4887 4747
rect 4873 4653 4887 4667
rect 4913 4813 4927 4827
rect 4913 4753 4927 4767
rect 5013 4913 5027 4927
rect 4973 4893 4987 4907
rect 5173 5072 5187 5086
rect 5273 5332 5287 5346
rect 5293 5153 5307 5167
rect 5093 5013 5107 5027
rect 5153 5032 5167 5046
rect 5133 4973 5147 4987
rect 5073 4953 5087 4967
rect 5113 4953 5127 4967
rect 5213 5032 5227 5046
rect 5233 5013 5247 5027
rect 5193 4953 5207 4967
rect 5033 4873 5047 4887
rect 5153 4913 5167 4927
rect 5113 4854 5127 4868
rect 5213 4854 5227 4868
rect 5593 5373 5607 5387
rect 5653 5374 5667 5388
rect 5733 5374 5747 5388
rect 5773 5374 5787 5388
rect 5373 5313 5387 5327
rect 5413 5332 5427 5346
rect 5493 5313 5507 5327
rect 5533 5313 5547 5327
rect 5333 5293 5347 5307
rect 5553 5133 5567 5147
rect 5433 5113 5447 5127
rect 5373 5074 5387 5088
rect 5293 5032 5307 5046
rect 5353 5032 5367 5046
rect 5393 5032 5407 5046
rect 5273 5013 5287 5027
rect 5453 5074 5467 5088
rect 5513 5074 5527 5088
rect 5253 4993 5267 5007
rect 5433 4993 5447 5007
rect 5613 5333 5627 5347
rect 5633 5293 5647 5307
rect 5673 5273 5687 5287
rect 5753 5293 5767 5307
rect 5693 5253 5707 5267
rect 5733 5253 5747 5267
rect 5693 5133 5707 5147
rect 5613 5073 5627 5087
rect 5453 4973 5467 4987
rect 5313 4953 5327 4967
rect 5293 4913 5307 4927
rect 4953 4813 4967 4827
rect 4933 4693 4947 4707
rect 5053 4813 5067 4827
rect 5093 4813 5107 4827
rect 5053 4773 5067 4787
rect 4993 4733 5007 4747
rect 4953 4593 4967 4607
rect 4873 4553 4887 4567
rect 4953 4554 4967 4568
rect 4853 4512 4867 4526
rect 4893 4512 4907 4526
rect 4973 4513 4987 4527
rect 4973 4473 4987 4487
rect 4833 4453 4847 4467
rect 4933 4453 4947 4467
rect 4833 4413 4847 4427
rect 4853 4373 4867 4387
rect 4893 4373 4907 4387
rect 4833 4353 4847 4367
rect 4813 4334 4827 4348
rect 4793 4113 4807 4127
rect 5133 4812 5147 4826
rect 5093 4773 5107 4787
rect 5153 4753 5167 4767
rect 5173 4733 5187 4747
rect 5093 4593 5107 4607
rect 5133 4593 5147 4607
rect 5093 4554 5107 4568
rect 5253 4854 5267 4868
rect 5533 5032 5547 5046
rect 5593 5032 5607 5046
rect 5613 4993 5627 5007
rect 5493 4913 5507 4927
rect 5473 4893 5487 4907
rect 5513 4893 5527 4907
rect 5553 4893 5567 4907
rect 5313 4854 5327 4868
rect 5373 4854 5387 4868
rect 5413 4854 5427 4868
rect 5453 4853 5467 4867
rect 5313 4813 5327 4827
rect 5393 4812 5407 4826
rect 5213 4733 5227 4747
rect 5413 4713 5427 4727
rect 5193 4593 5207 4607
rect 5313 4593 5327 4607
rect 5173 4554 5187 4568
rect 5213 4554 5227 4568
rect 5273 4553 5287 4567
rect 5313 4554 5327 4568
rect 5353 4554 5367 4568
rect 5013 4513 5027 4527
rect 5013 4373 5027 4387
rect 5073 4512 5087 4526
rect 5133 4513 5147 4527
rect 5193 4473 5207 4487
rect 5333 4512 5347 4526
rect 5393 4513 5407 4527
rect 5393 4473 5407 4487
rect 5273 4453 5287 4467
rect 5373 4453 5387 4467
rect 5233 4413 5247 4427
rect 5353 4413 5367 4427
rect 5053 4393 5067 4407
rect 5113 4393 5127 4407
rect 4933 4334 4947 4348
rect 5033 4353 5047 4367
rect 4893 4273 4907 4287
rect 4953 4273 4967 4287
rect 4913 4253 4927 4267
rect 4873 4053 4887 4067
rect 4813 3992 4827 4006
rect 4993 4133 5007 4147
rect 5313 4373 5327 4387
rect 5053 4093 5067 4107
rect 4973 4073 4987 4087
rect 5013 4053 5027 4067
rect 4973 4034 4987 4048
rect 5053 4034 5067 4048
rect 4913 3973 4927 3987
rect 4793 3933 4807 3947
rect 4853 3933 4867 3947
rect 4793 3893 4807 3907
rect 4873 3873 4887 3887
rect 4833 3814 4847 3828
rect 4893 3853 4907 3867
rect 4873 3813 4887 3827
rect 4733 3693 4747 3707
rect 4773 3693 4787 3707
rect 4813 3633 4827 3647
rect 4633 3593 4647 3607
rect 4673 3593 4687 3607
rect 4633 3553 4647 3567
rect 4873 3773 4887 3787
rect 4993 3992 5007 4006
rect 5033 3953 5047 3967
rect 5013 3933 5027 3947
rect 4993 3853 5007 3867
rect 4953 3814 4967 3828
rect 4933 3772 4947 3786
rect 4973 3772 4987 3786
rect 4873 3713 4887 3727
rect 4953 3693 4967 3707
rect 4793 3573 4807 3587
rect 4853 3573 4867 3587
rect 4913 3573 4927 3587
rect 4673 3514 4687 3528
rect 4713 3514 4727 3528
rect 4753 3514 4767 3528
rect 4573 3472 4587 3486
rect 4613 3472 4627 3486
rect 4653 3453 4667 3467
rect 4553 3413 4567 3427
rect 4653 3413 4667 3427
rect 4473 3353 4487 3367
rect 4313 3333 4327 3347
rect 4353 3333 4367 3347
rect 4453 3333 4467 3347
rect 4273 3294 4287 3308
rect 4213 3253 4227 3267
rect 4193 3093 4207 3107
rect 4173 3053 4187 3067
rect 4293 3253 4307 3267
rect 4253 3213 4267 3227
rect 4253 3173 4267 3187
rect 4253 3113 4267 3127
rect 4193 3013 4207 3027
rect 4213 2993 4227 3007
rect 4273 2993 4287 3007
rect 4193 2952 4207 2966
rect 4153 2933 4167 2947
rect 4213 2933 4227 2947
rect 4013 2913 4027 2927
rect 4093 2873 4107 2887
rect 3933 2833 3947 2847
rect 3973 2833 3987 2847
rect 3873 2793 3887 2807
rect 3913 2793 3927 2807
rect 3673 2733 3687 2747
rect 3593 2613 3607 2627
rect 3633 2613 3647 2627
rect 3513 2573 3527 2587
rect 3553 2473 3567 2487
rect 3633 2474 3647 2488
rect 3173 2432 3187 2446
rect 3213 2432 3227 2446
rect 3253 2432 3267 2446
rect 3293 2432 3307 2446
rect 3053 2393 3067 2407
rect 3113 2393 3127 2407
rect 3233 2393 3247 2407
rect 3093 2373 3107 2387
rect 2973 2333 2987 2347
rect 2813 2173 2827 2187
rect 2953 2173 2967 2187
rect 2893 2113 2907 2127
rect 2873 2073 2887 2087
rect 2813 1993 2827 2007
rect 2793 1912 2807 1926
rect 2833 1873 2847 1887
rect 2793 1833 2807 1847
rect 2833 1793 2847 1807
rect 2793 1734 2807 1748
rect 2873 1693 2887 1707
rect 2813 1653 2827 1667
rect 2793 1513 2807 1527
rect 2833 1453 2847 1467
rect 2753 1392 2767 1406
rect 2813 1392 2827 1406
rect 2753 1333 2767 1347
rect 2713 1233 2727 1247
rect 3033 2273 3047 2287
rect 3073 2273 3087 2287
rect 3093 2254 3107 2268
rect 3133 2254 3147 2268
rect 3173 2254 3187 2268
rect 3073 2153 3087 2167
rect 3073 2113 3087 2127
rect 3193 2212 3207 2226
rect 3393 2433 3407 2447
rect 3433 2432 3447 2446
rect 3493 2413 3507 2427
rect 3473 2333 3487 2347
rect 3293 2274 3307 2288
rect 3333 2273 3347 2287
rect 3293 2253 3307 2267
rect 3373 2253 3387 2267
rect 3433 2254 3447 2268
rect 3472 2254 3486 2268
rect 3613 2432 3627 2446
rect 3553 2353 3567 2367
rect 3733 2732 3747 2746
rect 3993 2813 4007 2827
rect 4033 2774 4047 2788
rect 4073 2773 4087 2787
rect 3833 2732 3847 2746
rect 3873 2732 3887 2746
rect 3913 2732 3927 2746
rect 3793 2693 3807 2707
rect 3693 2633 3707 2647
rect 3813 2573 3827 2587
rect 3713 2513 3727 2527
rect 3773 2474 3787 2488
rect 3713 2433 3727 2447
rect 3693 2353 3707 2367
rect 3633 2333 3647 2347
rect 3673 2333 3687 2347
rect 3493 2253 3507 2267
rect 3193 2191 3207 2205
rect 3233 2193 3247 2207
rect 3153 2173 3167 2187
rect 2973 2073 2987 2087
rect 2953 1954 2967 1968
rect 3013 1954 3027 1968
rect 3133 2093 3147 2107
rect 2913 1933 2927 1947
rect 2973 1912 2987 1926
rect 2933 1873 2947 1887
rect 2953 1793 2967 1807
rect 2913 1733 2927 1747
rect 2893 1633 2907 1647
rect 2933 1533 2947 1547
rect 2973 1773 2987 1787
rect 2973 1653 2987 1667
rect 3053 1912 3067 1926
rect 3153 2013 3167 2027
rect 3353 2213 3367 2227
rect 3313 2193 3327 2207
rect 3273 2153 3287 2167
rect 3373 2173 3387 2187
rect 3393 2153 3407 2167
rect 3353 2093 3367 2107
rect 3333 2073 3347 2087
rect 3513 2212 3527 2226
rect 3573 2193 3587 2207
rect 3453 2073 3467 2087
rect 3393 2033 3407 2047
rect 3333 2013 3347 2027
rect 3493 2013 3507 2027
rect 3593 2013 3607 2027
rect 3273 1993 3287 2007
rect 3193 1954 3207 1968
rect 3233 1954 3247 1968
rect 3273 1953 3287 1967
rect 3453 1993 3467 2007
rect 3373 1954 3387 1968
rect 3413 1954 3427 1968
rect 3533 1954 3547 1968
rect 3693 2254 3707 2268
rect 4013 2713 4027 2727
rect 3973 2693 3987 2707
rect 4053 2633 4067 2647
rect 4053 2593 4067 2607
rect 3893 2533 3907 2547
rect 3853 2513 3867 2527
rect 3833 2473 3847 2487
rect 3953 2474 3967 2488
rect 4013 2474 4027 2488
rect 4053 2473 4067 2487
rect 3853 2413 3867 2427
rect 3813 2333 3827 2347
rect 3753 2273 3767 2287
rect 3793 2273 3807 2287
rect 3833 2273 3847 2287
rect 3913 2432 3927 2446
rect 3873 2393 3887 2407
rect 4053 2393 4067 2407
rect 3993 2333 4007 2347
rect 3973 2273 3987 2287
rect 3853 2253 3867 2267
rect 3793 2212 3807 2226
rect 3873 2212 3887 2226
rect 3933 2212 3947 2226
rect 3753 2193 3767 2207
rect 3833 2193 3847 2207
rect 3733 2153 3747 2167
rect 3733 2113 3747 2127
rect 4053 2254 4067 2268
rect 4193 2833 4207 2847
rect 4113 2813 4127 2827
rect 4193 2793 4207 2807
rect 4113 2773 4127 2787
rect 4153 2774 4167 2788
rect 4173 2713 4187 2727
rect 4133 2693 4147 2707
rect 4093 2653 4107 2667
rect 4133 2432 4147 2446
rect 4233 2893 4247 2907
rect 4433 3313 4447 3327
rect 4353 3294 4367 3308
rect 4393 3294 4407 3308
rect 4573 3353 4587 3367
rect 4473 3293 4487 3307
rect 4593 3333 4607 3347
rect 4573 3293 4587 3307
rect 4453 3273 4467 3287
rect 4313 3233 4327 3247
rect 4373 3233 4387 3247
rect 4413 3213 4427 3227
rect 4453 3193 4467 3207
rect 4413 3153 4427 3167
rect 4393 3113 4407 3127
rect 4413 3033 4427 3047
rect 4313 2994 4327 3008
rect 4373 2994 4387 3008
rect 4393 2952 4407 2966
rect 4513 3252 4527 3266
rect 4553 3252 4567 3266
rect 4753 3453 4767 3467
rect 4733 3393 4747 3407
rect 4713 3333 4727 3347
rect 4693 3294 4707 3308
rect 4593 3252 4607 3266
rect 4633 3252 4647 3266
rect 4813 3472 4827 3486
rect 4773 3413 4787 3427
rect 4793 3294 4807 3308
rect 4833 3294 4847 3308
rect 4973 3613 4987 3627
rect 5053 3893 5067 3907
rect 5193 4292 5207 4306
rect 5233 4253 5247 4267
rect 5113 4093 5127 4107
rect 5213 4093 5227 4107
rect 5153 4034 5167 4048
rect 5133 3992 5147 4006
rect 5173 3953 5187 3967
rect 5193 3933 5207 3947
rect 5173 3913 5187 3927
rect 5093 3893 5107 3907
rect 5073 3873 5087 3887
rect 5093 3853 5107 3867
rect 5133 3853 5147 3867
rect 5093 3814 5107 3828
rect 5073 3772 5087 3786
rect 5113 3772 5127 3786
rect 5313 4333 5327 4347
rect 5393 4334 5407 4348
rect 5433 4593 5447 4607
rect 5673 4953 5687 4967
rect 5713 4893 5727 4907
rect 5653 4854 5667 4868
rect 5733 4853 5747 4867
rect 5493 4812 5507 4826
rect 5533 4812 5547 4826
rect 5593 4812 5607 4826
rect 5513 4613 5527 4627
rect 5453 4573 5467 4587
rect 5473 4554 5487 4568
rect 5493 4512 5507 4526
rect 5513 4413 5527 4427
rect 5453 4353 5467 4367
rect 5433 4334 5447 4348
rect 5333 4292 5347 4306
rect 5373 4253 5387 4267
rect 5313 4233 5327 4247
rect 5353 4153 5367 4167
rect 5313 4034 5327 4048
rect 5233 3933 5247 3947
rect 5213 3833 5227 3847
rect 5673 4812 5687 4826
rect 5713 4813 5727 4827
rect 5633 4733 5647 4747
rect 5593 4673 5607 4687
rect 5633 4613 5647 4627
rect 5593 4554 5607 4568
rect 5693 4573 5707 4587
rect 5613 4512 5627 4526
rect 5593 4453 5607 4467
rect 5433 4233 5447 4247
rect 5493 4292 5507 4306
rect 5473 4173 5487 4187
rect 5453 4153 5467 4167
rect 5453 4093 5467 4107
rect 5433 4034 5447 4048
rect 5293 3973 5307 3987
rect 5353 3973 5367 3987
rect 5353 3913 5367 3927
rect 5273 3893 5287 3907
rect 5253 3833 5267 3847
rect 5313 3853 5327 3867
rect 5273 3814 5287 3828
rect 5053 3613 5067 3627
rect 5133 3613 5147 3627
rect 4993 3553 5007 3567
rect 5033 3553 5047 3567
rect 5093 3553 5107 3567
rect 5033 3514 5047 3528
rect 4973 3472 4987 3486
rect 5013 3472 5027 3486
rect 5053 3472 5067 3486
rect 5173 3772 5187 3786
rect 5213 3772 5227 3786
rect 5233 3753 5247 3767
rect 5173 3514 5187 3528
rect 5093 3453 5107 3467
rect 4953 3433 4967 3447
rect 4893 3393 4907 3407
rect 5053 3393 5067 3407
rect 4573 3193 4587 3207
rect 4693 3113 4707 3127
rect 4493 3073 4507 3087
rect 4473 2994 4487 3008
rect 4653 3033 4667 3047
rect 4533 2994 4547 3008
rect 4733 3233 4747 3247
rect 4733 3113 4747 3127
rect 4713 3073 4727 3087
rect 4813 3252 4827 3266
rect 4773 3213 4787 3227
rect 4473 2953 4487 2967
rect 4813 3013 4827 3027
rect 4773 2994 4787 3008
rect 4853 3013 4867 3027
rect 4893 3293 4907 3307
rect 4933 3313 4947 3327
rect 4973 3294 4987 3308
rect 5013 3293 5027 3307
rect 5153 3453 5167 3467
rect 5133 3433 5147 3447
rect 5113 3313 5127 3327
rect 5093 3294 5107 3308
rect 5413 3992 5427 4006
rect 5573 4153 5587 4167
rect 5533 4073 5547 4087
rect 5533 4034 5547 4048
rect 5673 4513 5687 4527
rect 5613 4373 5627 4387
rect 5653 4373 5667 4387
rect 5753 4713 5767 4727
rect 5733 4673 5747 4687
rect 5793 5313 5807 5327
rect 5793 5273 5807 5287
rect 5793 4813 5807 4827
rect 5793 4653 5807 4667
rect 5752 4573 5766 4587
rect 5773 4573 5787 4587
rect 5713 4553 5727 4567
rect 5693 4493 5707 4507
rect 5693 4453 5707 4467
rect 5613 4333 5627 4347
rect 5673 4292 5687 4306
rect 5633 4253 5647 4267
rect 5613 4073 5627 4087
rect 5753 4493 5767 4507
rect 5733 4173 5747 4187
rect 5613 4034 5627 4048
rect 5653 4034 5667 4048
rect 5413 3833 5427 3847
rect 5333 3773 5347 3787
rect 5313 3753 5327 3767
rect 5373 3772 5387 3786
rect 5413 3753 5427 3767
rect 5333 3713 5347 3727
rect 5393 3573 5407 3587
rect 5253 3553 5267 3567
rect 5373 3533 5387 3547
rect 5293 3514 5307 3528
rect 5333 3514 5347 3528
rect 5493 3913 5507 3927
rect 5553 3992 5567 4006
rect 5513 3873 5527 3887
rect 5453 3573 5467 3587
rect 5573 3973 5587 3987
rect 5613 3973 5627 3987
rect 5673 3992 5687 4006
rect 5793 4493 5807 4507
rect 5773 4433 5787 4447
rect 5773 4213 5787 4227
rect 5633 3953 5647 3967
rect 5713 3953 5727 3967
rect 5633 3873 5647 3887
rect 5593 3813 5607 3827
rect 5633 3833 5647 3847
rect 5673 3814 5687 3828
rect 5773 3893 5787 3907
rect 5813 4433 5827 4447
rect 5793 3873 5807 3887
rect 5813 3833 5827 3847
rect 5713 3813 5727 3827
rect 5753 3814 5767 3828
rect 5793 3814 5807 3828
rect 5593 3773 5607 3787
rect 5533 3633 5547 3647
rect 5413 3533 5427 3547
rect 5433 3514 5447 3528
rect 5473 3514 5487 3528
rect 5233 3353 5247 3367
rect 5313 3472 5327 3486
rect 5373 3472 5387 3486
rect 5393 3433 5407 3447
rect 5153 3313 5167 3327
rect 4913 3252 4927 3266
rect 5013 3252 5027 3266
rect 5073 3252 5087 3266
rect 4953 3213 4967 3227
rect 5213 3294 5227 3308
rect 5253 3294 5267 3308
rect 4893 3173 4907 3187
rect 5113 3173 5127 3187
rect 5013 3113 5027 3127
rect 4873 2993 4887 3007
rect 4913 2994 4927 3008
rect 4953 2994 4967 3008
rect 4353 2933 4367 2947
rect 4453 2933 4467 2947
rect 4513 2952 4527 2966
rect 4473 2913 4487 2927
rect 4293 2893 4307 2907
rect 4633 2952 4647 2966
rect 4673 2952 4687 2966
rect 4733 2952 4747 2966
rect 4793 2933 4807 2947
rect 4773 2913 4787 2927
rect 4813 2913 4827 2927
rect 4813 2853 4827 2867
rect 4253 2833 4267 2847
rect 4513 2833 4527 2847
rect 4553 2833 4567 2847
rect 4293 2813 4307 2827
rect 4373 2813 4387 2827
rect 4253 2774 4267 2788
rect 4353 2732 4367 2746
rect 4213 2693 4227 2707
rect 4193 2593 4207 2607
rect 4233 2533 4247 2547
rect 4193 2513 4207 2527
rect 4173 2353 4187 2367
rect 4473 2774 4487 2788
rect 4393 2753 4407 2767
rect 4613 2813 4627 2827
rect 4793 2813 4807 2827
rect 4573 2793 4587 2807
rect 4713 2793 4727 2807
rect 4753 2774 4767 2788
rect 4513 2732 4527 2746
rect 4553 2732 4567 2746
rect 4453 2713 4467 2727
rect 4593 2713 4607 2727
rect 4733 2732 4747 2746
rect 4693 2713 4707 2727
rect 4613 2593 4627 2607
rect 4533 2533 4547 2547
rect 4373 2513 4387 2527
rect 4293 2474 4307 2488
rect 4353 2474 4367 2488
rect 4413 2473 4427 2487
rect 4253 2432 4267 2446
rect 4573 2513 4587 2527
rect 4753 2533 4767 2547
rect 4673 2474 4687 2488
rect 4713 2474 4727 2488
rect 4793 2513 4807 2527
rect 4413 2393 4427 2407
rect 4493 2432 4507 2446
rect 4533 2433 4547 2447
rect 4373 2353 4387 2367
rect 4473 2353 4487 2367
rect 4253 2333 4267 2347
rect 4193 2293 4207 2307
rect 4233 2293 4247 2307
rect 4153 2273 4167 2287
rect 3993 2193 4007 2207
rect 3973 2173 3987 2187
rect 3793 2113 3807 2127
rect 3753 2013 3767 2027
rect 3673 1973 3687 1987
rect 3733 1954 3747 1968
rect 3773 1954 3787 1968
rect 3093 1893 3107 1907
rect 3073 1873 3087 1887
rect 3013 1793 3027 1807
rect 3053 1692 3067 1706
rect 3033 1653 3047 1667
rect 3013 1613 3027 1627
rect 2993 1593 3007 1607
rect 2953 1513 2967 1527
rect 3013 1493 3027 1507
rect 2993 1473 3007 1487
rect 2913 1434 2927 1448
rect 2993 1433 3007 1447
rect 2973 1392 2987 1406
rect 2933 1353 2947 1367
rect 2893 1293 2907 1307
rect 2793 1233 2807 1247
rect 2873 1233 2887 1247
rect 2573 1172 2587 1186
rect 2673 1173 2687 1187
rect 2493 1153 2507 1167
rect 2533 1153 2547 1167
rect 2613 1153 2627 1167
rect 2533 1093 2547 1107
rect 2453 953 2467 967
rect 2493 953 2507 967
rect 2433 793 2447 807
rect 2433 733 2447 747
rect 2773 1173 2787 1187
rect 2853 1214 2867 1228
rect 2733 1093 2747 1107
rect 2613 953 2627 967
rect 2613 913 2627 927
rect 2653 914 2667 928
rect 2553 872 2567 886
rect 2593 873 2607 887
rect 2513 853 2527 867
rect 2673 873 2687 887
rect 2633 853 2647 867
rect 2613 793 2627 807
rect 2453 713 2467 727
rect 2553 713 2567 727
rect 2493 694 2507 708
rect 2433 633 2447 647
rect 2193 593 2207 607
rect 2413 593 2427 607
rect 2513 652 2527 666
rect 2073 573 2087 587
rect 2253 573 2267 587
rect 2473 573 2487 587
rect 2073 513 2087 527
rect 2053 493 2067 507
rect 2032 433 2046 447
rect 2053 433 2067 447
rect 2073 413 2087 427
rect 2093 394 2107 408
rect 2133 394 2147 408
rect 2173 394 2187 408
rect 2213 394 2227 408
rect 2413 513 2427 527
rect 2473 513 2487 527
rect 2273 433 2287 447
rect 2393 413 2407 427
rect 2033 352 2047 366
rect 2073 352 2087 366
rect 2053 273 2067 287
rect 2013 253 2027 267
rect 2293 394 2307 408
rect 2353 394 2367 408
rect 2433 493 2447 507
rect 2553 593 2567 607
rect 2473 473 2487 487
rect 2513 473 2527 487
rect 2433 453 2447 467
rect 2533 433 2547 447
rect 2493 394 2507 408
rect 2193 353 2207 367
rect 2273 353 2287 367
rect 2373 352 2387 366
rect 2293 313 2307 327
rect 2293 273 2307 287
rect 2533 273 2547 287
rect 2273 253 2287 267
rect 2193 213 2207 227
rect 2273 213 2287 227
rect 2413 213 2427 227
rect 2293 193 2307 207
rect 2153 174 2167 188
rect 2192 174 2206 188
rect 2213 173 2227 187
rect 2253 174 2267 188
rect 2333 174 2347 188
rect 213 33 227 47
rect 273 33 287 47
rect 793 33 807 47
rect 1273 33 1287 47
rect 1793 33 1807 47
rect 1893 33 1907 47
rect 1973 132 1987 146
rect 2033 132 2047 146
rect 2093 132 2107 146
rect 2693 773 2707 787
rect 2673 633 2687 647
rect 2733 593 2747 607
rect 2713 573 2727 587
rect 2633 533 2647 547
rect 2613 493 2627 507
rect 2653 493 2667 507
rect 2613 352 2627 366
rect 2613 213 2627 227
rect 2673 413 2687 427
rect 2733 553 2747 567
rect 2733 433 2747 447
rect 2753 413 2767 427
rect 2873 1172 2887 1186
rect 2953 1313 2967 1327
rect 2993 1273 3007 1287
rect 3093 1833 3107 1847
rect 3173 1893 3187 1907
rect 3213 1893 3227 1907
rect 3273 1873 3287 1887
rect 3153 1813 3167 1827
rect 3233 1813 3247 1827
rect 3113 1793 3127 1807
rect 3113 1692 3127 1706
rect 3173 1692 3187 1706
rect 3073 1593 3087 1607
rect 3053 1493 3067 1507
rect 3193 1434 3207 1448
rect 3053 1373 3067 1387
rect 3033 1353 3047 1367
rect 3093 1333 3107 1347
rect 3353 1912 3367 1926
rect 3413 1893 3427 1907
rect 3353 1853 3367 1867
rect 3313 1773 3327 1787
rect 3293 1734 3307 1748
rect 3453 1793 3467 1807
rect 3393 1734 3407 1748
rect 3353 1693 3367 1707
rect 3413 1692 3427 1706
rect 3533 1913 3547 1927
rect 3613 1853 3627 1867
rect 3693 1813 3707 1827
rect 3773 1813 3787 1827
rect 3573 1793 3587 1807
rect 3473 1733 3487 1747
rect 3513 1734 3527 1748
rect 3553 1734 3567 1748
rect 3472 1692 3486 1706
rect 3493 1692 3507 1706
rect 3353 1633 3367 1647
rect 3253 1593 3267 1607
rect 3053 1313 3067 1327
rect 3233 1313 3247 1327
rect 3313 1353 3327 1367
rect 3113 1293 3127 1307
rect 2973 1233 2987 1247
rect 3013 1233 3027 1247
rect 3053 1233 3067 1247
rect 3033 1213 3047 1227
rect 2993 1172 3007 1186
rect 3033 1173 3047 1187
rect 3133 1233 3147 1247
rect 2993 1093 3007 1107
rect 2933 973 2947 987
rect 2873 953 2887 967
rect 2813 914 2827 928
rect 2913 873 2927 887
rect 2793 793 2807 807
rect 3013 1073 3027 1087
rect 2873 773 2887 787
rect 2993 773 3007 787
rect 2833 733 2847 747
rect 3113 1172 3127 1186
rect 3173 1172 3187 1186
rect 3133 1133 3147 1147
rect 3313 1273 3327 1287
rect 3273 1113 3287 1127
rect 3233 1093 3247 1107
rect 3173 1073 3187 1087
rect 3153 1053 3167 1067
rect 3113 1013 3127 1027
rect 3053 914 3067 928
rect 3073 793 3087 807
rect 3053 773 3067 787
rect 2973 753 2987 767
rect 3013 753 3027 767
rect 2873 694 2887 708
rect 2913 693 2927 707
rect 3013 694 3027 708
rect 2993 652 3007 666
rect 3033 653 3047 667
rect 2913 633 2927 647
rect 2913 533 2927 547
rect 2853 513 2867 527
rect 2873 413 2887 427
rect 2793 393 2807 407
rect 2833 394 2847 408
rect 3013 473 3027 487
rect 2973 453 2987 467
rect 2933 413 2947 427
rect 2913 393 2927 407
rect 2673 352 2687 366
rect 2713 313 2727 327
rect 2653 193 2667 207
rect 2553 153 2567 167
rect 2413 132 2427 146
rect 2453 132 2467 146
rect 2513 132 2527 146
rect 2213 93 2227 107
rect 2273 93 2287 107
rect 2633 93 2647 107
rect 3053 613 3067 627
rect 3033 453 3047 467
rect 3053 433 3067 447
rect 2793 313 2807 327
rect 2893 352 2907 366
rect 2933 353 2947 367
rect 2993 352 3007 366
rect 3033 333 3047 347
rect 3233 1013 3247 1027
rect 3213 973 3227 987
rect 3273 953 3287 967
rect 3193 813 3207 827
rect 3233 813 3247 827
rect 3173 793 3187 807
rect 3233 773 3247 787
rect 3433 1434 3447 1448
rect 3453 1393 3467 1407
rect 3653 1692 3667 1706
rect 3773 1773 3787 1787
rect 3713 1734 3727 1748
rect 3993 2073 4007 2087
rect 3913 1954 3927 1968
rect 4113 2253 4127 2267
rect 4193 2254 4207 2268
rect 4253 2253 4267 2267
rect 4313 2254 4327 2268
rect 4113 2212 4127 2226
rect 4213 2212 4227 2226
rect 4253 2213 4267 2227
rect 4293 2212 4307 2226
rect 4173 2193 4187 2207
rect 4093 1973 4107 1987
rect 4133 1973 4147 1987
rect 4193 1973 4207 1987
rect 3853 1912 3867 1926
rect 4093 1912 4107 1926
rect 3853 1813 3867 1827
rect 4093 1813 4107 1827
rect 4073 1793 4087 1807
rect 3873 1773 3887 1787
rect 3793 1753 3807 1767
rect 3833 1753 3847 1767
rect 3593 1673 3607 1687
rect 3693 1673 3707 1687
rect 3533 1633 3547 1647
rect 3513 1493 3527 1507
rect 3553 1434 3567 1448
rect 3733 1473 3747 1487
rect 3673 1453 3687 1467
rect 3713 1452 3727 1466
rect 3413 1353 3427 1367
rect 3453 1273 3467 1287
rect 3313 1213 3327 1227
rect 3353 1214 3367 1228
rect 3413 1213 3427 1227
rect 3573 1392 3587 1406
rect 3713 1393 3727 1407
rect 3533 1313 3547 1327
rect 3493 1214 3507 1228
rect 3333 1172 3347 1186
rect 3373 1172 3387 1186
rect 3393 1113 3407 1127
rect 3313 973 3327 987
rect 3293 933 3307 947
rect 3353 914 3367 928
rect 3373 873 3387 887
rect 3373 813 3387 827
rect 3413 973 3427 987
rect 3593 1233 3607 1247
rect 3633 1233 3647 1247
rect 3793 1392 3807 1406
rect 3933 1733 3947 1747
rect 3973 1734 3987 1748
rect 4013 1734 4027 1748
rect 3893 1692 3907 1706
rect 3933 1692 3947 1706
rect 3993 1673 4007 1687
rect 4053 1693 4067 1707
rect 3893 1633 3907 1647
rect 4033 1633 4047 1647
rect 3853 1513 3867 1527
rect 4213 1912 4227 1926
rect 4413 2333 4427 2347
rect 4473 2332 4487 2346
rect 4452 2254 4466 2268
rect 4633 2432 4647 2446
rect 4593 2393 4607 2407
rect 4733 2432 4747 2446
rect 4793 2433 4807 2447
rect 4693 2413 4707 2427
rect 4673 2353 4687 2367
rect 4493 2273 4507 2287
rect 4553 2273 4567 2287
rect 4613 2273 4627 2287
rect 4653 2273 4667 2287
rect 4473 2253 4487 2267
rect 4373 2073 4387 2087
rect 4333 2033 4347 2047
rect 4413 2033 4427 2047
rect 4253 1833 4267 1847
rect 4393 1912 4407 1926
rect 4313 1833 4327 1847
rect 4273 1813 4287 1827
rect 4133 1793 4147 1807
rect 4273 1773 4287 1787
rect 4173 1753 4187 1767
rect 4093 1733 4107 1747
rect 4133 1734 4147 1748
rect 4293 1753 4307 1767
rect 4193 1734 4207 1748
rect 4253 1734 4267 1748
rect 4073 1673 4087 1687
rect 4053 1453 4067 1467
rect 3913 1434 3927 1448
rect 4013 1434 4027 1448
rect 3893 1392 3907 1406
rect 3853 1373 3867 1387
rect 3833 1353 3847 1367
rect 4113 1392 4127 1406
rect 3933 1373 3947 1387
rect 3893 1333 3907 1347
rect 3653 1214 3667 1228
rect 3713 1214 3727 1228
rect 3753 1214 3767 1228
rect 3973 1214 3987 1228
rect 4393 1793 4407 1807
rect 4533 2212 4547 2226
rect 4573 2212 4587 2226
rect 4493 2033 4507 2047
rect 4433 2013 4447 2027
rect 4593 2013 4607 2027
rect 4693 2253 4707 2267
rect 4613 1993 4627 2007
rect 4653 1993 4667 2007
rect 4473 1954 4487 1968
rect 4513 1954 4527 1968
rect 4713 2212 4727 2226
rect 4773 2212 4787 2226
rect 4713 2013 4727 2027
rect 4533 1913 4547 1927
rect 4533 1813 4547 1827
rect 4473 1793 4487 1807
rect 4413 1753 4427 1767
rect 4453 1753 4467 1767
rect 4193 1673 4207 1687
rect 4253 1673 4267 1687
rect 4153 1593 4167 1607
rect 4173 1533 4187 1547
rect 4233 1513 4247 1527
rect 4173 1493 4187 1507
rect 4133 1233 4147 1247
rect 3613 1172 3627 1186
rect 3653 1153 3667 1167
rect 3573 1133 3587 1147
rect 3853 1153 3867 1167
rect 3753 1133 3767 1147
rect 3793 1133 3807 1147
rect 3753 1093 3767 1107
rect 3533 1073 3547 1087
rect 3733 1073 3747 1087
rect 3633 973 3647 987
rect 3513 933 3527 947
rect 3453 914 3467 928
rect 3593 914 3607 928
rect 3693 914 3707 928
rect 3633 872 3647 886
rect 3673 872 3687 886
rect 3713 872 3727 886
rect 3573 833 3587 847
rect 3673 833 3687 847
rect 3713 833 3727 847
rect 3653 813 3667 827
rect 3413 773 3427 787
rect 3513 773 3527 787
rect 3333 733 3347 747
rect 3393 733 3407 747
rect 3373 713 3387 727
rect 3093 652 3107 666
rect 3093 573 3107 587
rect 3133 493 3147 507
rect 3213 652 3227 666
rect 3253 573 3267 587
rect 3193 553 3207 567
rect 3193 513 3207 527
rect 3213 493 3227 507
rect 3173 433 3187 447
rect 3213 453 3227 467
rect 3253 453 3267 467
rect 3333 694 3347 708
rect 4093 1214 4107 1228
rect 4053 1013 4067 1027
rect 3833 973 3847 987
rect 4113 973 4127 987
rect 3793 933 3807 947
rect 4193 1353 4207 1367
rect 4373 1692 4387 1706
rect 4413 1692 4427 1706
rect 4433 1633 4447 1647
rect 4353 1513 4367 1527
rect 4413 1513 4427 1527
rect 4333 1453 4347 1467
rect 4273 1434 4287 1448
rect 4313 1434 4327 1448
rect 4393 1453 4407 1467
rect 4273 1333 4287 1347
rect 4233 1214 4247 1228
rect 4393 1392 4407 1406
rect 4413 1313 4427 1327
rect 4293 1253 4307 1267
rect 4333 1253 4347 1267
rect 4453 1593 4467 1607
rect 4513 1753 4527 1767
rect 4593 1733 4607 1747
rect 4773 1954 4787 1968
rect 4973 2952 4987 2966
rect 5033 3033 5047 3047
rect 5073 2994 5087 3008
rect 5113 2993 5127 3007
rect 5033 2953 5047 2967
rect 5093 2952 5107 2966
rect 4873 2913 4887 2927
rect 4933 2913 4947 2927
rect 4973 2913 4987 2927
rect 5013 2913 5027 2927
rect 4953 2893 4967 2907
rect 4893 2853 4907 2867
rect 4833 2813 4847 2827
rect 4873 2732 4887 2746
rect 4873 2474 4887 2488
rect 5153 3252 5167 3266
rect 5233 3252 5247 3266
rect 5453 3472 5467 3486
rect 5693 3773 5707 3787
rect 5613 3713 5627 3727
rect 5593 3593 5607 3607
rect 5593 3553 5607 3567
rect 5553 3514 5567 3528
rect 5753 3713 5767 3727
rect 5733 3673 5747 3687
rect 5673 3633 5687 3647
rect 5673 3593 5687 3607
rect 5713 3633 5727 3647
rect 5733 3593 5747 3607
rect 5713 3533 5727 3547
rect 5632 3513 5646 3527
rect 5653 3513 5667 3527
rect 5693 3514 5707 3528
rect 5753 3513 5767 3527
rect 5193 3193 5207 3207
rect 5293 3193 5307 3207
rect 5213 3173 5227 3187
rect 5253 3053 5267 3067
rect 5233 2993 5247 3007
rect 5073 2853 5087 2867
rect 5133 2853 5147 2867
rect 5053 2833 5067 2847
rect 5033 2813 5047 2827
rect 5053 2793 5067 2807
rect 5013 2774 5027 2788
rect 4993 2732 5007 2746
rect 5113 2813 5127 2827
rect 5153 2774 5167 2788
rect 5233 2913 5247 2927
rect 5293 3033 5307 3047
rect 5373 3233 5387 3247
rect 5373 3113 5387 3127
rect 5473 3193 5487 3207
rect 5413 3133 5427 3147
rect 5473 3133 5487 3147
rect 5433 2994 5447 3008
rect 5513 3472 5527 3486
rect 5573 3472 5587 3486
rect 5613 3472 5627 3486
rect 5633 3453 5647 3467
rect 5533 3433 5547 3447
rect 5513 3293 5527 3307
rect 5493 3053 5507 3067
rect 5633 3333 5647 3347
rect 5593 3294 5607 3308
rect 5753 3473 5767 3487
rect 5673 3293 5687 3307
rect 5533 3233 5547 3247
rect 5573 3133 5587 3147
rect 5653 3252 5667 3266
rect 5633 3213 5647 3227
rect 5613 3093 5627 3107
rect 5513 3013 5527 3027
rect 5253 2873 5267 2887
rect 5353 2952 5367 2966
rect 5393 2952 5407 2966
rect 5453 2952 5467 2966
rect 5533 2953 5547 2967
rect 5353 2913 5367 2927
rect 5213 2813 5227 2827
rect 5313 2813 5327 2827
rect 5253 2793 5267 2807
rect 4993 2613 5007 2627
rect 4953 2593 4967 2607
rect 4913 2473 4927 2487
rect 4953 2474 4967 2488
rect 5053 2732 5067 2746
rect 5093 2732 5107 2746
rect 5173 2733 5187 2747
rect 5133 2713 5147 2727
rect 5113 2553 5127 2567
rect 5073 2474 5087 2488
rect 5213 2773 5227 2787
rect 5293 2774 5307 2788
rect 5333 2773 5347 2787
rect 5273 2732 5287 2746
rect 5233 2713 5247 2727
rect 5213 2673 5227 2687
rect 5193 2653 5207 2667
rect 5313 2593 5327 2607
rect 5213 2573 5227 2587
rect 5253 2493 5267 2507
rect 4973 2432 4987 2446
rect 5033 2433 5047 2447
rect 5213 2474 5227 2488
rect 5453 2873 5467 2887
rect 5393 2774 5407 2788
rect 5353 2732 5367 2746
rect 5653 2952 5667 2966
rect 5573 2893 5587 2907
rect 5513 2853 5527 2867
rect 5513 2813 5527 2827
rect 5473 2793 5487 2807
rect 5553 2774 5567 2788
rect 5713 3313 5727 3327
rect 5813 3773 5827 3787
rect 5793 3753 5807 3767
rect 5773 3293 5787 3307
rect 5693 2952 5707 2966
rect 5673 2893 5687 2907
rect 5613 2873 5627 2887
rect 5593 2853 5607 2867
rect 5653 2813 5667 2827
rect 5593 2773 5607 2787
rect 5693 2774 5707 2788
rect 5753 3252 5767 3266
rect 5773 3233 5787 3247
rect 5773 3193 5787 3207
rect 5733 2994 5747 3008
rect 5753 2933 5767 2947
rect 5773 2793 5787 2807
rect 5813 3693 5827 3707
rect 5813 3672 5827 3686
rect 5813 2933 5827 2947
rect 5493 2732 5507 2746
rect 5533 2732 5547 2746
rect 5333 2553 5347 2567
rect 5373 2474 5387 2488
rect 5413 2473 5427 2487
rect 5473 2573 5487 2587
rect 5553 2573 5567 2587
rect 5533 2493 5547 2507
rect 5093 2432 5107 2446
rect 5153 2432 5167 2446
rect 5193 2432 5207 2446
rect 5233 2432 5247 2446
rect 4913 2373 4927 2387
rect 5053 2373 5067 2387
rect 4953 2273 4967 2287
rect 5013 2273 5027 2287
rect 4893 2254 4907 2268
rect 5412 2432 5426 2446
rect 5433 2432 5447 2446
rect 5493 2432 5507 2446
rect 5433 2373 5447 2387
rect 5533 2373 5547 2387
rect 5313 2353 5327 2367
rect 5273 2313 5287 2327
rect 5093 2293 5107 2307
rect 5253 2293 5267 2307
rect 4953 2213 4967 2227
rect 5033 2212 5047 2226
rect 4993 2173 5007 2187
rect 4833 2113 4847 2127
rect 4873 2033 4887 2047
rect 4813 1953 4827 1967
rect 4933 1953 4947 1967
rect 5013 1954 5027 1968
rect 5053 1953 5067 1967
rect 4753 1893 4767 1907
rect 4693 1853 4707 1867
rect 4493 1693 4507 1707
rect 4573 1693 4587 1707
rect 4553 1673 4567 1687
rect 4513 1593 4527 1607
rect 4473 1573 4487 1587
rect 4453 1513 4467 1527
rect 4513 1493 4527 1507
rect 4453 1434 4467 1448
rect 4513 1434 4527 1448
rect 4493 1392 4507 1406
rect 4573 1433 4587 1447
rect 4653 1734 4667 1748
rect 4693 1734 4707 1748
rect 4713 1692 4727 1706
rect 4613 1653 4627 1667
rect 4673 1653 4687 1667
rect 4793 1853 4807 1867
rect 4833 1793 4847 1807
rect 4773 1733 4787 1747
rect 4873 1753 4887 1767
rect 4773 1692 4787 1706
rect 4813 1573 4827 1587
rect 4853 1553 4867 1567
rect 4753 1513 4767 1527
rect 5013 1773 5027 1787
rect 4973 1734 4987 1748
rect 4913 1673 4927 1687
rect 4993 1692 5007 1706
rect 5033 1692 5047 1706
rect 4953 1653 4967 1667
rect 4813 1473 4827 1487
rect 4893 1473 4907 1487
rect 4733 1453 4747 1467
rect 4553 1373 4567 1387
rect 4593 1373 4607 1387
rect 4473 1273 4487 1287
rect 4453 1253 4467 1267
rect 4313 1214 4327 1228
rect 4373 1214 4387 1228
rect 4433 1213 4447 1227
rect 4273 1193 4287 1207
rect 4213 1113 4227 1127
rect 4273 1113 4287 1127
rect 4213 1073 4227 1087
rect 4173 933 4187 947
rect 3893 913 3907 927
rect 3853 872 3867 886
rect 3893 872 3907 886
rect 3833 833 3847 847
rect 3873 833 3887 847
rect 3753 793 3767 807
rect 3893 793 3907 807
rect 3673 773 3687 787
rect 3513 733 3527 747
rect 3653 733 3667 747
rect 3533 713 3547 727
rect 3413 693 3427 707
rect 3513 693 3527 707
rect 3353 652 3367 666
rect 3393 652 3407 666
rect 3353 553 3367 567
rect 3253 413 3267 427
rect 3213 393 3227 407
rect 3273 394 3287 408
rect 3113 333 3127 347
rect 3073 293 3087 307
rect 2853 273 2867 287
rect 2733 253 2747 267
rect 3153 253 3167 267
rect 2793 233 2807 247
rect 2753 193 2767 207
rect 2793 174 2807 188
rect 2833 174 2847 188
rect 2913 173 2927 187
rect 3113 174 3127 188
rect 3153 174 3167 188
rect 3253 352 3267 366
rect 3293 313 3307 327
rect 3233 293 3247 307
rect 3233 193 3247 207
rect 3213 173 3227 187
rect 2913 132 2927 146
rect 2953 132 2967 146
rect 3013 132 3027 146
rect 3173 132 3187 146
rect 2773 93 2787 107
rect 3133 93 3147 107
rect 2673 53 2687 67
rect 2713 53 2727 67
rect 1913 13 1927 27
rect 3513 653 3527 667
rect 3493 633 3507 647
rect 3433 613 3447 627
rect 3373 533 3387 547
rect 3413 533 3427 547
rect 3353 393 3367 407
rect 3553 694 3567 708
rect 3613 694 3627 708
rect 3533 633 3547 647
rect 3733 694 3747 708
rect 3773 694 3787 708
rect 3833 694 3847 708
rect 3673 633 3687 647
rect 3553 573 3567 587
rect 3793 633 3807 647
rect 4073 914 4087 928
rect 4133 913 4147 927
rect 4213 914 4227 928
rect 4053 872 4067 886
rect 4093 872 4107 886
rect 4293 973 4307 987
rect 4373 1133 4387 1147
rect 4433 1133 4447 1147
rect 4353 933 4367 947
rect 4273 893 4287 907
rect 4133 872 4147 886
rect 4193 872 4207 886
rect 4013 833 4027 847
rect 4113 833 4127 847
rect 3953 773 3967 787
rect 4213 773 4227 787
rect 3913 733 3927 747
rect 4073 733 4087 747
rect 3813 593 3827 607
rect 3893 593 3907 607
rect 3793 573 3807 587
rect 3673 553 3687 567
rect 3753 553 3767 567
rect 3513 513 3527 527
rect 3473 413 3487 427
rect 3513 413 3527 427
rect 3433 394 3447 408
rect 3373 352 3387 366
rect 3393 293 3407 307
rect 3393 253 3407 267
rect 3573 394 3587 408
rect 3633 394 3647 408
rect 4053 694 4067 708
rect 3953 633 3967 647
rect 4053 653 4067 667
rect 4133 694 4147 708
rect 4193 693 4207 707
rect 4113 652 4127 666
rect 4193 652 4207 666
rect 4073 633 4087 647
rect 4153 633 4167 647
rect 4013 593 4027 607
rect 3813 533 3827 547
rect 3913 533 3927 547
rect 3953 533 3967 547
rect 4153 533 4167 547
rect 3753 513 3767 527
rect 3713 493 3727 507
rect 3493 353 3507 367
rect 3473 313 3487 327
rect 3533 352 3547 366
rect 3472 292 3486 306
rect 3493 293 3507 307
rect 3413 233 3427 247
rect 3613 293 3627 307
rect 3573 233 3587 247
rect 3653 233 3667 247
rect 3473 213 3487 227
rect 3553 213 3567 227
rect 3433 193 3447 207
rect 3453 173 3467 187
rect 3493 174 3507 188
rect 3233 132 3247 146
rect 3333 132 3347 146
rect 3393 132 3407 146
rect 3433 133 3447 147
rect 3273 113 3287 127
rect 3293 93 3307 107
rect 3293 53 3307 67
rect 3333 13 3347 27
rect 3513 93 3527 107
rect 3633 174 3647 188
rect 3913 493 3927 507
rect 3873 453 3887 467
rect 3813 394 3827 408
rect 3753 213 3767 227
rect 3853 313 3867 327
rect 3893 293 3907 307
rect 3813 273 3827 287
rect 3873 233 3887 247
rect 3773 193 3787 207
rect 3613 132 3627 146
rect 3653 133 3667 147
rect 3553 73 3567 87
rect 3753 113 3767 127
rect 3733 73 3747 87
rect 3773 73 3787 87
rect 4133 473 4147 487
rect 4113 453 4127 467
rect 4093 413 4107 427
rect 4013 394 4027 408
rect 3993 313 4007 327
rect 4273 733 4287 747
rect 4313 694 4327 708
rect 4353 694 4367 708
rect 4253 652 4267 666
rect 4353 653 4367 667
rect 4433 1093 4447 1107
rect 4433 1053 4447 1067
rect 4413 1013 4427 1027
rect 4473 1213 4487 1227
rect 4493 1172 4507 1186
rect 4473 1133 4487 1147
rect 4553 1133 4567 1147
rect 4453 1033 4467 1047
rect 4593 1093 4607 1107
rect 4513 1053 4527 1067
rect 4653 1393 4667 1407
rect 4773 1434 4787 1448
rect 4753 1392 4767 1406
rect 4753 1313 4767 1327
rect 4693 1253 4707 1267
rect 4653 1214 4667 1228
rect 4713 1172 4727 1186
rect 4633 1153 4647 1167
rect 4673 1153 4687 1167
rect 4873 1434 4887 1448
rect 4933 1433 4947 1447
rect 4993 1434 5007 1448
rect 4853 1392 4867 1406
rect 4933 1392 4947 1406
rect 4973 1392 4987 1406
rect 5153 2254 5167 2268
rect 5193 2254 5207 2268
rect 5133 2212 5147 2226
rect 5313 2253 5327 2267
rect 5373 2254 5387 2268
rect 5533 2293 5547 2307
rect 5453 2254 5467 2268
rect 5493 2254 5507 2268
rect 5613 2733 5627 2747
rect 5633 2713 5647 2727
rect 5713 2733 5727 2747
rect 5713 2673 5727 2687
rect 5693 2593 5707 2607
rect 5593 2513 5607 2527
rect 5653 2513 5667 2527
rect 5613 2474 5627 2488
rect 5573 2393 5587 2407
rect 5633 2393 5647 2407
rect 5613 2293 5627 2307
rect 5273 2212 5287 2226
rect 5313 2212 5327 2226
rect 5193 2193 5207 2207
rect 5233 2193 5247 2207
rect 5353 2193 5367 2207
rect 5433 2212 5447 2226
rect 5593 2253 5607 2267
rect 5513 2212 5527 2226
rect 5553 2212 5567 2226
rect 5453 2193 5467 2207
rect 5493 2193 5507 2207
rect 5453 2033 5467 2047
rect 5293 1993 5307 2007
rect 5413 1993 5427 2007
rect 5133 1973 5147 1987
rect 5193 1953 5207 1967
rect 5233 1954 5247 1968
rect 5333 1953 5347 1967
rect 5373 1954 5387 1968
rect 5093 1912 5107 1926
rect 5133 1773 5147 1787
rect 5093 1653 5107 1667
rect 5053 1593 5067 1607
rect 5173 1692 5187 1706
rect 5153 1653 5167 1667
rect 5113 1473 5127 1487
rect 5073 1434 5087 1448
rect 5133 1433 5147 1447
rect 4893 1313 4907 1327
rect 4973 1313 4987 1327
rect 5033 1313 5047 1327
rect 4813 1253 4827 1267
rect 4873 1253 4887 1267
rect 4793 1214 4807 1228
rect 4833 1214 4847 1228
rect 4753 1093 4767 1107
rect 4713 1033 4727 1047
rect 4613 993 4627 1007
rect 4653 993 4667 1007
rect 4513 973 4527 987
rect 4533 953 4547 967
rect 4653 953 4667 967
rect 4693 953 4707 967
rect 4433 773 4447 787
rect 4413 713 4427 727
rect 4453 733 4467 747
rect 4393 652 4407 666
rect 4233 573 4247 587
rect 4233 533 4247 547
rect 4192 493 4206 507
rect 4213 493 4227 507
rect 4153 433 4167 447
rect 4473 713 4487 727
rect 4453 513 4467 527
rect 4333 493 4347 507
rect 4273 394 4287 408
rect 4373 394 4387 408
rect 4113 352 4127 366
rect 4113 293 4127 307
rect 4093 233 4107 247
rect 4033 213 4047 227
rect 3993 193 4007 207
rect 4213 352 4227 366
rect 4313 352 4327 366
rect 4273 313 4287 327
rect 4233 213 4247 227
rect 4173 173 4187 187
rect 3953 93 3967 107
rect 4373 313 4387 327
rect 4353 233 4367 247
rect 4513 914 4527 928
rect 4573 914 4587 928
rect 4613 914 4627 928
rect 4653 914 4667 928
rect 4693 913 4707 927
rect 4793 1013 4807 1027
rect 4753 914 4767 928
rect 4533 873 4547 887
rect 4493 693 4507 707
rect 4633 872 4647 886
rect 4673 873 4687 887
rect 4733 872 4747 886
rect 4713 773 4727 787
rect 4593 733 4607 747
rect 4593 693 4607 707
rect 4693 694 4707 708
rect 4513 652 4527 666
rect 4493 533 4507 547
rect 4473 213 4487 227
rect 4573 653 4587 667
rect 4673 652 4687 666
rect 4593 633 4607 647
rect 4593 593 4607 607
rect 4553 493 4567 507
rect 4513 433 4527 447
rect 4533 413 4547 427
rect 4513 394 4527 408
rect 4653 493 4667 507
rect 4833 1053 4847 1067
rect 4813 953 4827 967
rect 5073 1273 5087 1287
rect 5013 1233 5027 1247
rect 4933 1214 4947 1228
rect 4973 1214 4987 1228
rect 5113 1313 5127 1327
rect 5093 1233 5107 1247
rect 5253 1912 5267 1926
rect 5213 1793 5227 1807
rect 5413 1893 5427 1907
rect 5393 1773 5407 1787
rect 5273 1734 5287 1748
rect 5333 1734 5347 1748
rect 5393 1733 5407 1747
rect 5213 1693 5227 1707
rect 5253 1553 5267 1567
rect 5293 1533 5307 1547
rect 5493 1954 5507 1968
rect 5613 1953 5627 1967
rect 5473 1912 5487 1926
rect 5513 1912 5527 1926
rect 5553 1912 5567 1926
rect 5453 1813 5467 1827
rect 5753 2773 5767 2787
rect 5793 2774 5807 2788
rect 5773 2732 5787 2746
rect 5733 2474 5747 2488
rect 5793 2713 5807 2727
rect 5693 2353 5707 2367
rect 5673 2313 5687 2327
rect 5753 2432 5767 2446
rect 5733 2393 5747 2407
rect 5773 2393 5787 2407
rect 5713 2273 5727 2287
rect 5753 2353 5767 2367
rect 5693 2033 5707 2047
rect 5733 1973 5747 1987
rect 5773 2273 5787 2287
rect 5673 1954 5687 1968
rect 5693 1813 5707 1827
rect 5673 1773 5687 1787
rect 5633 1753 5647 1767
rect 5453 1692 5467 1706
rect 5633 1692 5647 1706
rect 5513 1653 5527 1667
rect 5573 1653 5587 1667
rect 5433 1533 5447 1547
rect 5253 1493 5267 1507
rect 5293 1473 5307 1487
rect 5193 1453 5207 1467
rect 5233 1453 5247 1467
rect 5253 1434 5267 1448
rect 5333 1434 5347 1448
rect 5213 1353 5227 1367
rect 5253 1353 5267 1367
rect 5393 1493 5407 1507
rect 5393 1433 5407 1447
rect 5553 1473 5567 1487
rect 5473 1434 5487 1448
rect 5513 1434 5527 1448
rect 5593 1434 5607 1448
rect 5773 1773 5787 1787
rect 5813 2474 5827 2488
rect 5813 2313 5827 2327
rect 5813 1973 5827 1987
rect 5753 1734 5767 1748
rect 5793 1734 5807 1748
rect 5813 1653 5827 1667
rect 5693 1513 5707 1527
rect 5753 1513 5767 1527
rect 5693 1473 5707 1487
rect 5413 1392 5427 1406
rect 5373 1333 5387 1347
rect 5313 1313 5327 1327
rect 5233 1253 5247 1267
rect 4913 1153 4927 1167
rect 5013 1172 5027 1186
rect 5053 1172 5067 1186
rect 5193 1214 5207 1228
rect 5233 1214 5247 1228
rect 5273 1214 5287 1228
rect 5313 1214 5327 1228
rect 5173 1172 5187 1186
rect 5133 1153 5147 1167
rect 4953 1133 4967 1147
rect 5293 1113 5307 1127
rect 5333 1073 5347 1087
rect 4873 1013 4887 1027
rect 5093 993 5107 1007
rect 5213 993 5227 1007
rect 4873 914 4887 928
rect 4933 914 4947 928
rect 4993 914 5007 928
rect 5133 914 5147 928
rect 5193 914 5207 928
rect 4893 872 4907 886
rect 4933 873 4947 887
rect 4853 793 4867 807
rect 4733 733 4747 747
rect 4793 733 4807 747
rect 5013 872 5027 886
rect 5153 872 5167 886
rect 5113 813 5127 827
rect 5013 773 5027 787
rect 4973 713 4987 727
rect 4773 694 4787 708
rect 5033 694 5047 708
rect 5153 694 5167 708
rect 4733 652 4747 666
rect 4813 652 4827 666
rect 4853 633 4867 647
rect 4973 652 4987 666
rect 5133 652 5147 666
rect 5413 1233 5427 1247
rect 5493 1393 5507 1407
rect 5613 1392 5627 1406
rect 5653 1392 5667 1406
rect 5573 1353 5587 1367
rect 5513 1333 5527 1347
rect 5493 1313 5507 1327
rect 5713 1373 5727 1387
rect 5753 1373 5767 1387
rect 5653 1273 5667 1287
rect 5513 1253 5527 1267
rect 5453 1214 5467 1228
rect 5553 1214 5567 1228
rect 5653 1214 5667 1228
rect 5793 1273 5807 1287
rect 5813 1213 5827 1227
rect 5393 1173 5407 1187
rect 5433 1172 5447 1186
rect 5393 953 5407 967
rect 5453 953 5467 967
rect 5413 914 5427 928
rect 5213 793 5227 807
rect 5373 873 5387 887
rect 5673 1113 5687 1127
rect 5713 1073 5727 1087
rect 5673 953 5687 967
rect 5553 914 5567 928
rect 5293 813 5307 827
rect 5353 813 5367 827
rect 5273 753 5287 767
rect 5413 773 5427 787
rect 5253 694 5267 708
rect 5373 694 5387 708
rect 4913 633 4927 647
rect 4753 613 4767 627
rect 4773 533 4787 547
rect 4853 533 4867 547
rect 4993 533 5007 547
rect 4733 473 4747 487
rect 4713 433 4727 447
rect 4693 394 4707 408
rect 4913 513 4927 527
rect 5073 433 5087 447
rect 4632 352 4646 366
rect 4653 352 4667 366
rect 4533 273 4547 287
rect 4413 173 4427 187
rect 4393 132 4407 146
rect 4494 173 4508 187
rect 4613 233 4627 247
rect 4593 213 4607 227
rect 4313 113 4327 127
rect 4353 113 4367 127
rect 4613 173 4627 187
rect 4753 352 4767 366
rect 4813 352 4827 366
rect 5133 413 5147 427
rect 5213 653 5227 667
rect 5213 453 5227 467
rect 5253 413 5267 427
rect 5353 413 5367 427
rect 5213 394 5227 408
rect 5173 353 5187 367
rect 5373 394 5387 408
rect 5473 872 5487 886
rect 5533 872 5547 886
rect 5813 1173 5827 1187
rect 5773 953 5787 967
rect 5773 914 5787 928
rect 5473 694 5487 708
rect 5513 694 5527 708
rect 5733 753 5747 767
rect 5473 633 5487 647
rect 5633 652 5647 666
rect 5693 633 5707 647
rect 5573 394 5587 408
rect 5813 633 5827 647
rect 5773 394 5787 408
rect 5233 352 5247 366
rect 5293 352 5307 366
rect 5353 352 5367 366
rect 4713 313 4727 327
rect 5093 313 5107 327
rect 4853 233 4867 247
rect 5093 233 5107 247
rect 4673 193 4687 207
rect 4733 193 4747 207
rect 4853 193 4867 207
rect 4913 193 4927 207
rect 4693 132 4707 146
rect 4553 113 4567 127
rect 4593 113 4607 127
rect 4653 113 4667 127
rect 4793 174 4807 188
rect 4812 132 4826 146
rect 4833 132 4847 146
rect 4773 93 4787 107
rect 5333 173 5347 187
rect 5453 273 5467 287
rect 5633 352 5647 366
rect 5673 353 5687 367
rect 5633 313 5647 327
rect 5553 253 5567 267
rect 5593 253 5607 267
rect 5453 193 5467 207
rect 5513 193 5527 207
rect 4973 132 4987 146
rect 4913 93 4927 107
rect 4513 73 4527 87
rect 4793 73 4807 87
rect 4833 73 4847 87
rect 5213 113 5227 127
rect 5333 132 5347 146
rect 5413 132 5427 146
rect 5553 173 5567 187
rect 5573 132 5587 146
rect 5373 93 5387 107
rect 5513 93 5527 107
rect 5753 352 5767 366
rect 5793 353 5807 367
rect 5713 313 5727 327
rect 5753 313 5767 327
rect 5793 313 5807 327
rect 5693 233 5707 247
rect 5713 173 5727 187
rect 5693 133 5707 147
rect 5733 132 5747 146
rect 5773 132 5787 146
rect 5673 113 5687 127
rect 5633 73 5647 87
rect 5813 73 5827 87
rect 5033 33 5047 47
rect 5273 33 5287 47
rect 5633 33 5647 47
<< metal3 >>
rect 2967 5476 3013 5484
rect 3787 5476 3833 5484
rect 907 5456 1313 5464
rect 1827 5456 2033 5464
rect 2047 5456 2573 5464
rect 2947 5456 3053 5464
rect 3147 5456 3253 5464
rect 3507 5456 3673 5464
rect 3727 5456 4113 5464
rect 1187 5436 1493 5444
rect 1547 5436 1733 5444
rect 1947 5436 2093 5444
rect 2647 5436 3073 5444
rect 3127 5436 3192 5444
rect 3227 5436 3693 5444
rect 3707 5436 4133 5444
rect 4707 5436 4913 5444
rect 127 5416 253 5424
rect 307 5416 412 5424
rect 447 5416 613 5424
rect 627 5416 733 5424
rect 1047 5416 1513 5424
rect 1527 5416 1653 5424
rect 1667 5416 1753 5424
rect 1867 5416 2253 5424
rect 2267 5416 2393 5424
rect 2767 5416 2793 5424
rect 2807 5416 2933 5424
rect 3367 5416 3753 5424
rect 3767 5416 4073 5424
rect 4167 5416 4313 5424
rect 4327 5416 4393 5424
rect 4507 5416 4853 5424
rect 3207 5396 3533 5404
rect 4027 5396 4053 5404
rect 5187 5396 5353 5404
rect 187 5376 213 5384
rect 280 5384 292 5387
rect 276 5373 292 5384
rect 327 5376 373 5384
rect 427 5376 493 5384
rect 667 5377 693 5385
rect 787 5377 833 5385
rect 847 5376 993 5384
rect 1007 5376 1133 5384
rect 1327 5377 1353 5385
rect 1407 5376 1453 5384
rect 276 5346 284 5373
rect 1256 5364 1264 5374
rect 1567 5376 1593 5384
rect 1676 5376 1693 5384
rect 1676 5364 1684 5376
rect 1787 5377 1933 5385
rect 1987 5376 2053 5384
rect 2147 5376 2193 5384
rect 2307 5376 2333 5384
rect 2447 5376 2473 5384
rect 2547 5376 2633 5384
rect 2656 5376 2673 5384
rect 2656 5364 2664 5376
rect 2747 5376 2913 5384
rect 3133 5384 3147 5393
rect 3133 5380 3173 5384
rect 3136 5376 3173 5380
rect 3327 5377 3393 5385
rect 3467 5376 3484 5384
rect 796 5356 1144 5364
rect 1256 5356 1304 5364
rect 796 5346 804 5356
rect 976 5346 984 5356
rect 367 5335 433 5343
rect 1027 5336 1113 5344
rect 1136 5344 1144 5356
rect 1136 5336 1153 5344
rect 1167 5336 1273 5344
rect 1296 5344 1304 5356
rect 1636 5356 1684 5364
rect 2496 5356 2664 5364
rect 2676 5356 2924 5364
rect 1296 5336 1413 5344
rect 1467 5335 1493 5343
rect 1636 5344 1644 5356
rect 1587 5336 1644 5344
rect 1767 5335 1793 5343
rect 2007 5335 2033 5343
rect 2207 5335 2273 5343
rect 2287 5336 2373 5344
rect 2496 5344 2504 5356
rect 2676 5344 2684 5356
rect 2467 5336 2504 5344
rect 2616 5340 2684 5344
rect 2613 5336 2684 5340
rect 355 5324 363 5332
rect 2613 5327 2627 5336
rect 2827 5336 2893 5344
rect 2916 5344 2924 5356
rect 2916 5336 2933 5344
rect 167 5316 363 5324
rect 587 5316 753 5324
rect 767 5316 873 5324
rect 887 5316 1353 5324
rect 1527 5316 2133 5324
rect 2247 5316 2413 5324
rect 407 5296 473 5304
rect 487 5296 593 5304
rect 607 5296 693 5304
rect 1967 5296 2113 5304
rect 2167 5296 2453 5304
rect 3036 5304 3044 5373
rect 3076 5364 3084 5374
rect 3076 5356 3264 5364
rect 3067 5335 3093 5343
rect 3207 5336 3233 5344
rect 3256 5344 3264 5356
rect 3256 5336 3293 5344
rect 3407 5336 3433 5344
rect 3476 5344 3484 5376
rect 3527 5377 3593 5385
rect 3807 5376 3824 5384
rect 3816 5347 3824 5376
rect 3856 5376 3873 5384
rect 3856 5347 3864 5376
rect 3887 5376 3973 5384
rect 3996 5376 4133 5384
rect 3476 5336 3513 5344
rect 3707 5335 3733 5343
rect 3996 5346 4004 5376
rect 4187 5376 4213 5384
rect 4236 5376 4273 5384
rect 4073 5344 4087 5353
rect 4236 5347 4244 5376
rect 4447 5376 4513 5384
rect 4556 5364 4564 5374
rect 4787 5376 4813 5384
rect 5067 5376 5113 5384
rect 5267 5377 5313 5385
rect 5327 5376 5393 5384
rect 5407 5376 5513 5384
rect 5567 5376 5593 5384
rect 4556 5356 4613 5364
rect 5216 5364 5224 5374
rect 5747 5377 5773 5385
rect 4967 5356 5224 5364
rect 4047 5336 4113 5344
rect 4467 5335 4493 5343
rect 5027 5336 5133 5344
rect 5287 5336 5413 5344
rect 5656 5344 5664 5374
rect 5627 5336 5664 5344
rect 3547 5316 3653 5324
rect 3667 5316 3713 5324
rect 4327 5316 4353 5324
rect 4887 5316 4913 5324
rect 4927 5316 5373 5324
rect 5387 5316 5493 5324
rect 5547 5316 5793 5324
rect 2907 5296 3044 5304
rect 3067 5296 3233 5304
rect 3307 5296 3473 5304
rect 3567 5296 3633 5304
rect 3787 5296 4073 5304
rect 4087 5296 4453 5304
rect 4547 5296 4673 5304
rect 5007 5296 5093 5304
rect 5107 5296 5333 5304
rect 5647 5296 5753 5304
rect 247 5276 773 5284
rect 1507 5276 1673 5284
rect 1687 5276 1833 5284
rect 2187 5276 2553 5284
rect 2567 5276 2713 5284
rect 2927 5276 3273 5284
rect 3507 5276 3544 5284
rect 3536 5267 3544 5276
rect 3727 5276 3873 5284
rect 4167 5276 4253 5284
rect 4267 5276 4953 5284
rect 5687 5276 5793 5284
rect 527 5256 933 5264
rect 947 5256 1933 5264
rect 2487 5256 2604 5264
rect 1547 5236 1633 5244
rect 1647 5236 2153 5244
rect 2596 5244 2604 5256
rect 2887 5256 3053 5264
rect 3156 5256 3373 5264
rect 3156 5247 3164 5256
rect 3447 5256 3473 5264
rect 3536 5256 3553 5267
rect 3540 5253 3553 5256
rect 3707 5256 3993 5264
rect 4627 5256 5013 5264
rect 5707 5256 5733 5264
rect 2596 5236 2873 5244
rect 3107 5236 3153 5244
rect 3247 5236 3573 5244
rect 3627 5236 4293 5244
rect 4307 5236 4413 5244
rect 1467 5216 2513 5224
rect 2567 5216 2673 5224
rect 2687 5216 2913 5224
rect 2927 5216 3073 5224
rect 3327 5216 3453 5224
rect 3607 5216 3864 5224
rect 287 5196 313 5204
rect 327 5196 1533 5204
rect 1587 5196 2353 5204
rect 2507 5196 2773 5204
rect 2827 5196 3193 5204
rect 3207 5196 3253 5204
rect 3347 5196 3513 5204
rect 3647 5196 3753 5204
rect 3856 5204 3864 5216
rect 3887 5216 4613 5224
rect 3856 5196 4533 5204
rect 4607 5196 4993 5204
rect 647 5176 673 5184
rect 687 5176 813 5184
rect 1667 5176 1953 5184
rect 1967 5176 2233 5184
rect 2627 5176 2964 5184
rect 87 5156 253 5164
rect 387 5156 884 5164
rect 347 5136 733 5144
rect 787 5136 853 5144
rect 876 5144 884 5156
rect 1307 5156 1513 5164
rect 2527 5156 2552 5164
rect 2587 5156 2813 5164
rect 2956 5164 2964 5176
rect 2987 5176 3092 5184
rect 3127 5176 3713 5184
rect 4227 5176 4453 5184
rect 4596 5184 4604 5193
rect 4507 5176 4604 5184
rect 4627 5176 4833 5184
rect 2956 5156 3153 5164
rect 3367 5156 3533 5164
rect 4047 5156 4233 5164
rect 5027 5156 5293 5164
rect 876 5136 1673 5144
rect 1727 5136 1913 5144
rect 2087 5136 2213 5144
rect 2227 5136 2393 5144
rect 2667 5136 3233 5144
rect 3307 5136 3573 5144
rect 3907 5136 3953 5144
rect 4007 5136 4413 5144
rect 4487 5136 4793 5144
rect 4807 5136 5553 5144
rect 5567 5136 5693 5144
rect 107 5116 973 5124
rect 1427 5116 1873 5124
rect 1916 5124 1924 5133
rect 1916 5116 2493 5124
rect 2827 5116 2852 5124
rect 2887 5116 2953 5124
rect 2967 5116 3073 5124
rect 3367 5116 3533 5124
rect 3847 5116 3873 5124
rect 4367 5116 4573 5124
rect 5127 5116 5433 5124
rect 267 5096 373 5104
rect 2087 5096 2113 5104
rect 2347 5096 2453 5104
rect 3347 5096 3533 5104
rect 127 5076 173 5084
rect 187 5077 233 5085
rect 427 5077 453 5085
rect 567 5076 584 5084
rect 147 5036 213 5044
rect 227 5036 493 5044
rect 516 5024 524 5074
rect 576 5044 584 5076
rect 576 5036 753 5044
rect 887 5035 913 5043
rect 976 5044 984 5074
rect 1027 5076 1073 5084
rect 1147 5077 1173 5085
rect 1227 5077 1273 5085
rect 1287 5076 1313 5084
rect 1640 5084 1653 5087
rect 1456 5047 1464 5074
rect 976 5036 1053 5044
rect 1447 5036 1464 5047
rect 1496 5047 1504 5074
rect 1636 5073 1653 5084
rect 1767 5077 1793 5085
rect 1496 5036 1512 5047
rect 1447 5033 1460 5036
rect 1500 5033 1512 5036
rect 1636 5046 1644 5073
rect 1836 5047 1844 5074
rect 2047 5076 2253 5084
rect 2267 5077 2313 5085
rect 2336 5076 2353 5084
rect 1913 5064 1927 5073
rect 2336 5064 2344 5076
rect 2687 5076 2704 5084
rect 2573 5064 2587 5073
rect 1913 5060 1964 5064
rect 1916 5056 1964 5060
rect 1547 5036 1593 5044
rect 1827 5036 1844 5047
rect 1827 5033 1840 5036
rect 1907 5036 1933 5044
rect 516 5016 673 5024
rect 1267 5016 1413 5024
rect 1427 5016 1473 5024
rect 1667 5016 1733 5024
rect 1956 5024 1964 5056
rect 2256 5056 2344 5064
rect 2436 5060 2587 5064
rect 2696 5064 2704 5076
rect 2436 5056 2584 5060
rect 2696 5056 2733 5064
rect 2027 5035 2073 5043
rect 2147 5036 2233 5044
rect 2256 5044 2264 5056
rect 2247 5036 2264 5044
rect 2436 5044 2444 5056
rect 2756 5047 2764 5093
rect 3727 5096 3893 5104
rect 4007 5096 4053 5104
rect 4067 5096 4113 5104
rect 4916 5096 5033 5104
rect 4916 5088 4924 5096
rect 5047 5096 5073 5104
rect 2827 5076 3113 5084
rect 3327 5076 3353 5084
rect 3176 5047 3184 5073
rect 3416 5064 3424 5074
rect 3507 5084 3520 5087
rect 3507 5073 3524 5084
rect 3587 5076 3613 5084
rect 3627 5076 3693 5084
rect 3867 5076 4153 5084
rect 4167 5076 4193 5084
rect 4367 5077 4393 5085
rect 4447 5076 4533 5084
rect 4847 5076 4913 5084
rect 4936 5076 4953 5084
rect 3356 5060 3464 5064
rect 3353 5056 3467 5060
rect 3353 5047 3367 5056
rect 2307 5036 2444 5044
rect 2456 5036 2604 5044
rect 1956 5016 1993 5024
rect 2456 5024 2464 5036
rect 2407 5016 2464 5024
rect 2487 5016 2519 5024
rect 2596 5024 2604 5036
rect 2627 5035 2653 5043
rect 2667 5040 2724 5044
rect 2667 5036 2727 5040
rect 2713 5027 2727 5036
rect 2987 5036 3053 5044
rect 3307 5036 3332 5044
rect 3453 5047 3467 5056
rect 3516 5046 3524 5073
rect 3747 5056 4724 5064
rect 3607 5036 3673 5044
rect 4716 5046 4724 5056
rect 4936 5064 4944 5076
rect 4976 5076 5013 5084
rect 4867 5056 4944 5064
rect 4976 5046 4984 5076
rect 5187 5077 5373 5085
rect 5467 5077 5513 5085
rect 5613 5064 5627 5073
rect 5613 5060 5644 5064
rect 5616 5056 5644 5060
rect 3907 5036 3933 5044
rect 3987 5035 4033 5043
rect 4047 5036 4133 5044
rect 4207 5035 4253 5043
rect 4427 5036 4553 5044
rect 4727 5035 4793 5043
rect 5167 5035 5213 5043
rect 5307 5035 5353 5043
rect 5407 5036 5533 5044
rect 5547 5036 5593 5044
rect 2596 5016 2704 5024
rect 847 4996 1013 5004
rect 1287 4996 1593 5004
rect 1736 5004 1744 5013
rect 1736 4996 2013 5004
rect 2127 4996 2313 5004
rect 2327 4996 2373 5004
rect 2467 4996 2493 5004
rect 2587 4996 2673 5004
rect 2696 5004 2704 5016
rect 2827 5016 3013 5024
rect 3447 5016 3473 5024
rect 3767 5016 3833 5024
rect 4947 5016 5093 5024
rect 5247 5016 5273 5024
rect 5636 5007 5644 5056
rect 2696 4996 3133 5004
rect 3267 4996 3353 5004
rect 3407 4996 3533 5004
rect 3587 4996 3633 5004
rect 3647 4996 3733 5004
rect 3787 4996 4253 5004
rect 4587 4996 4653 5004
rect 5267 4996 5433 5004
rect 5627 4996 5644 5007
rect 5627 4993 5640 4996
rect 667 4976 733 4984
rect 1127 4976 1193 4984
rect 1687 4976 1793 4984
rect 1807 4976 3213 4984
rect 3396 4984 3404 4993
rect 3227 4976 3404 4984
rect 3807 4976 4333 4984
rect 4447 4976 4553 4984
rect 5147 4976 5453 4984
rect 5467 4976 5604 4984
rect 167 4956 353 4964
rect 1347 4956 1573 4964
rect 1707 4956 1784 4964
rect 407 4936 433 4944
rect 447 4936 533 4944
rect 547 4936 633 4944
rect 767 4936 953 4944
rect 1147 4936 1253 4944
rect 1527 4936 1613 4944
rect 1776 4944 1784 4956
rect 1847 4956 2392 4964
rect 2427 4956 2733 4964
rect 2747 4956 2793 4964
rect 2907 4956 3204 4964
rect 1776 4936 1973 4944
rect 2427 4936 2692 4944
rect 2727 4936 2753 4944
rect 2920 4944 2933 4947
rect 2916 4933 2933 4944
rect 3196 4944 3204 4956
rect 3467 4956 3573 4964
rect 3947 4956 4053 4964
rect 4207 4956 4313 4964
rect 4367 4956 4513 4964
rect 4787 4956 5073 4964
rect 5087 4956 5113 4964
rect 5207 4956 5313 4964
rect 5596 4964 5604 4976
rect 5596 4956 5673 4964
rect 3196 4936 3293 4944
rect 3607 4936 4053 4944
rect 127 4916 253 4924
rect 1327 4916 1713 4924
rect 2147 4916 2273 4924
rect 2367 4916 2493 4924
rect 2916 4924 2924 4933
rect 4067 4936 4873 4944
rect 2507 4916 2924 4924
rect 2947 4916 3093 4924
rect 3407 4916 3713 4924
rect 3927 4916 4444 4924
rect 47 4896 73 4904
rect 407 4896 453 4904
rect 467 4896 573 4904
rect 587 4896 793 4904
rect 1587 4896 1653 4904
rect 2187 4896 2412 4904
rect 2447 4896 2553 4904
rect 2707 4896 2733 4904
rect 2747 4896 2873 4904
rect 2927 4896 2973 4904
rect 3347 4896 3793 4904
rect 3907 4896 3993 4904
rect 4007 4896 4353 4904
rect 4436 4904 4444 4916
rect 4587 4916 4753 4924
rect 5027 4916 5153 4924
rect 5167 4916 5293 4924
rect 5307 4916 5493 4924
rect 4436 4896 4553 4904
rect 4607 4896 4973 4904
rect 5487 4896 5513 4904
rect 5567 4896 5713 4904
rect 56 4876 93 4884
rect 56 4827 64 4876
rect 187 4876 353 4884
rect 707 4884 720 4887
rect 707 4873 724 4884
rect 1007 4876 1173 4884
rect 1187 4876 1373 4884
rect 1867 4876 2153 4884
rect 2207 4876 2244 4884
rect 140 4864 153 4867
rect 136 4853 153 4864
rect 420 4864 432 4867
rect 287 4856 304 4864
rect 136 4826 144 4853
rect 296 4827 304 4856
rect 416 4853 432 4864
rect 467 4856 493 4864
rect 560 4864 573 4867
rect 556 4853 573 4864
rect 147 4816 253 4824
rect 416 4826 424 4853
rect 556 4826 564 4853
rect 676 4844 684 4854
rect 616 4840 684 4844
rect 613 4836 684 4840
rect 716 4847 724 4873
rect 767 4864 780 4867
rect 767 4853 784 4864
rect 807 4856 873 4864
rect 967 4857 1033 4865
rect 1207 4856 1293 4864
rect 1547 4856 1673 4864
rect 716 4846 740 4847
rect 716 4836 733 4846
rect 613 4827 627 4836
rect 720 4833 733 4836
rect 776 4826 784 4853
rect 1287 4815 1313 4823
rect 1407 4815 1453 4823
rect 1496 4824 1504 4854
rect 1747 4856 1833 4864
rect 1887 4857 2073 4865
rect 2187 4864 2200 4867
rect 2187 4853 2204 4864
rect 1467 4816 1504 4824
rect 1527 4816 1593 4824
rect 2196 4826 2204 4853
rect 1707 4816 1773 4824
rect 1967 4816 2033 4824
rect 2236 4824 2244 4876
rect 2687 4876 2833 4884
rect 3127 4876 3153 4884
rect 4847 4876 5033 4884
rect 2256 4844 2264 4854
rect 2447 4856 2533 4864
rect 2893 4864 2907 4873
rect 2920 4864 2933 4867
rect 2836 4860 2907 4864
rect 2836 4856 2904 4860
rect 2256 4836 2444 4844
rect 2336 4826 2344 4836
rect 2236 4820 2264 4824
rect 2236 4816 2267 4820
rect 2253 4807 2267 4816
rect 2356 4816 2413 4824
rect 327 4796 373 4804
rect 847 4796 1193 4804
rect 376 4784 384 4793
rect 376 4776 513 4784
rect 767 4776 1253 4784
rect 1367 4776 1513 4784
rect 1527 4776 1553 4784
rect 1567 4776 1633 4784
rect 1947 4776 1993 4784
rect 2007 4776 2113 4784
rect 2356 4784 2364 4816
rect 2436 4824 2444 4836
rect 2596 4827 2604 4853
rect 2436 4816 2513 4824
rect 2636 4824 2644 4854
rect 2636 4816 2713 4824
rect 2407 4796 2733 4804
rect 2776 4804 2784 4854
rect 2836 4824 2844 4856
rect 2916 4853 2933 4864
rect 2976 4856 2993 4864
rect 2916 4844 2924 4853
rect 2856 4836 2924 4844
rect 2856 4826 2864 4836
rect 2976 4827 2984 4856
rect 3047 4857 3093 4865
rect 3387 4856 3453 4864
rect 3736 4856 3813 4864
rect 3676 4827 3684 4854
rect 2807 4816 2844 4824
rect 3027 4815 3113 4823
rect 3227 4815 3253 4823
rect 3347 4816 3413 4824
rect 3667 4816 3684 4827
rect 3736 4826 3744 4856
rect 3667 4813 3680 4816
rect 2776 4796 2913 4804
rect 3067 4796 3393 4804
rect 3856 4804 3864 4854
rect 3927 4856 3953 4864
rect 4007 4856 4104 4864
rect 3896 4824 3904 4853
rect 4096 4829 4104 4856
rect 4307 4856 4353 4864
rect 4487 4857 4513 4865
rect 4596 4856 4613 4864
rect 3887 4816 3904 4824
rect 4556 4827 4564 4853
rect 4596 4827 4604 4856
rect 4667 4856 4713 4864
rect 5227 4857 5253 4865
rect 5327 4857 5373 4865
rect 5427 4856 5453 4864
rect 4856 4827 4864 4853
rect 4147 4816 4213 4824
rect 4287 4815 4313 4823
rect 4327 4815 4333 4823
rect 4767 4815 4832 4823
rect 4876 4824 4884 4854
rect 5116 4827 5124 4854
rect 5667 4856 5733 4864
rect 4876 4816 4913 4824
rect 4967 4816 5053 4824
rect 5107 4816 5124 4827
rect 5107 4813 5120 4816
rect 5147 4816 5313 4824
rect 5407 4816 5493 4824
rect 5547 4815 5593 4823
rect 5607 4816 5673 4824
rect 5727 4816 5793 4824
rect 3856 4796 3973 4804
rect 4107 4796 4224 4804
rect 2247 4776 2364 4784
rect 2487 4776 2673 4784
rect 2767 4776 2853 4784
rect 3307 4776 3333 4784
rect 3347 4776 3373 4784
rect 3707 4776 3913 4784
rect 4216 4784 4224 4796
rect 4447 4796 4513 4804
rect 4216 4776 4233 4784
rect 4247 4776 4413 4784
rect 4507 4776 4553 4784
rect 4887 4776 5053 4784
rect 267 4756 293 4764
rect 1247 4756 1353 4764
rect 1396 4756 1753 4764
rect 607 4736 813 4744
rect 1396 4744 1404 4756
rect 1776 4756 2413 4764
rect 1267 4736 1404 4744
rect 1776 4744 1784 4756
rect 2527 4756 2613 4764
rect 2927 4756 3093 4764
rect 3487 4756 3893 4764
rect 4007 4756 4193 4764
rect 4687 4756 4913 4764
rect 5093 4764 5107 4773
rect 4927 4756 5153 4764
rect 1467 4736 1784 4744
rect 1827 4736 2393 4744
rect 2527 4736 2692 4744
rect 2727 4736 2893 4744
rect 2907 4736 3373 4744
rect 3847 4736 4013 4744
rect 4487 4736 4673 4744
rect 4687 4736 4873 4744
rect 5007 4736 5173 4744
rect 5187 4736 5213 4744
rect 5227 4736 5633 4744
rect 307 4716 833 4724
rect 1047 4716 1153 4724
rect 2387 4716 2453 4724
rect 2467 4716 2573 4724
rect 3507 4716 3993 4724
rect 4087 4716 4233 4724
rect 4247 4716 4373 4724
rect 4447 4716 4713 4724
rect 5427 4716 5753 4724
rect 107 4696 213 4704
rect 227 4696 473 4704
rect 1547 4696 1733 4704
rect 2027 4696 2793 4704
rect 4647 4696 4793 4704
rect 4807 4696 4933 4704
rect 927 4676 1372 4684
rect 1407 4676 1433 4684
rect 1447 4676 1964 4684
rect 607 4656 873 4664
rect 1507 4656 1693 4664
rect 1807 4656 1893 4664
rect 1956 4664 1964 4676
rect 2127 4676 2393 4684
rect 2447 4676 2833 4684
rect 2887 4676 2933 4684
rect 2987 4676 3013 4684
rect 3067 4676 3413 4684
rect 4047 4676 4173 4684
rect 4387 4676 4493 4684
rect 5607 4676 5733 4684
rect 1956 4656 4073 4664
rect 4227 4656 4873 4664
rect 5616 4656 5793 4664
rect 1267 4636 1653 4644
rect 1796 4636 1933 4644
rect 27 4616 133 4624
rect 147 4616 533 4624
rect 747 4616 773 4624
rect 1487 4616 1673 4624
rect 1796 4624 1804 4636
rect 2187 4636 2333 4644
rect 2427 4636 2632 4644
rect 2667 4636 3053 4644
rect 3407 4636 3513 4644
rect 3587 4636 4093 4644
rect 4587 4636 4713 4644
rect 5616 4644 5624 4656
rect 4847 4636 5624 4644
rect 1687 4616 1804 4624
rect 1847 4616 1973 4624
rect 2147 4616 2953 4624
rect 3127 4616 3193 4624
rect 3207 4616 3293 4624
rect 3667 4616 3893 4624
rect 3907 4616 3993 4624
rect 4007 4616 4193 4624
rect 4567 4616 4593 4624
rect 4607 4616 5513 4624
rect 5527 4616 5633 4624
rect 1007 4596 1053 4604
rect 1207 4596 1813 4604
rect 1907 4596 2213 4604
rect 2227 4596 2293 4604
rect 2307 4596 2433 4604
rect 2447 4596 2573 4604
rect 2627 4596 2724 4604
rect 187 4576 373 4584
rect 547 4576 573 4584
rect 587 4576 753 4584
rect 1107 4576 1293 4584
rect 1307 4576 1393 4584
rect 1667 4576 1793 4584
rect 2027 4576 2053 4584
rect 2716 4584 2724 4596
rect 2747 4596 2933 4604
rect 2987 4596 3433 4604
rect 3447 4596 3593 4604
rect 3787 4596 3933 4604
rect 4407 4600 4624 4604
rect 4407 4596 4627 4600
rect 4613 4587 4627 4596
rect 4667 4596 4733 4604
rect 4747 4596 4773 4604
rect 4967 4596 5093 4604
rect 5147 4596 5193 4604
rect 5327 4596 5433 4604
rect 2716 4576 2733 4584
rect 67 4557 93 4565
rect 307 4556 333 4564
rect 56 4527 64 4554
rect 487 4556 513 4564
rect 813 4564 827 4573
rect 813 4560 844 4564
rect 816 4556 844 4560
rect 127 4515 173 4523
rect 647 4520 744 4524
rect 647 4516 747 4520
rect 733 4507 747 4516
rect 547 4496 573 4504
rect 87 4476 193 4484
rect 207 4476 273 4484
rect 627 4476 673 4484
rect 796 4484 804 4533
rect 836 4524 844 4556
rect 967 4557 1033 4565
rect 1347 4556 1413 4564
rect 1427 4557 1473 4565
rect 1496 4556 1553 4564
rect 1156 4544 1164 4554
rect 1496 4544 1504 4556
rect 2036 4556 2093 4564
rect 1836 4544 1844 4554
rect 2036 4544 2044 4556
rect 2267 4556 2293 4564
rect 2347 4556 2473 4564
rect 1156 4536 1264 4544
rect 836 4516 1013 4524
rect 1127 4516 1173 4524
rect 1256 4524 1264 4536
rect 1456 4536 1504 4544
rect 1796 4536 1844 4544
rect 1996 4536 2044 4544
rect 1256 4516 1313 4524
rect 1367 4516 1432 4524
rect 1456 4507 1464 4536
rect 1667 4516 1716 4524
rect 1796 4524 1804 4536
rect 1776 4516 1804 4524
rect 1440 4505 1464 4507
rect 1067 4496 1284 4504
rect 796 4476 853 4484
rect 947 4476 1153 4484
rect 1276 4484 1284 4496
rect 1447 4496 1464 4505
rect 1447 4493 1460 4496
rect 1567 4496 1693 4504
rect 1776 4504 1784 4516
rect 1827 4516 1853 4524
rect 1996 4526 2004 4536
rect 1927 4516 1953 4524
rect 2047 4516 2273 4524
rect 2367 4515 2413 4523
rect 2587 4515 2633 4523
rect 2656 4507 2664 4573
rect 2747 4576 2813 4584
rect 4087 4576 4473 4584
rect 5707 4576 5752 4584
rect 5787 4584 5800 4587
rect 5787 4573 5804 4584
rect 2776 4544 2784 4554
rect 2756 4540 2784 4544
rect 2753 4536 2784 4540
rect 2753 4527 2767 4536
rect 2976 4527 2984 4554
rect 3087 4556 3184 4564
rect 2806 4515 2853 4523
rect 2976 4516 2993 4527
rect 2980 4513 2993 4516
rect 1747 4496 1784 4504
rect 2027 4496 2313 4504
rect 3036 4504 3044 4553
rect 3176 4526 3184 4556
rect 3267 4556 3333 4564
rect 3487 4557 3693 4565
rect 3707 4556 3833 4564
rect 4227 4557 4273 4565
rect 4507 4556 4533 4564
rect 4547 4556 4553 4564
rect 4647 4556 4753 4564
rect 4887 4564 4900 4567
rect 4887 4553 4904 4564
rect 5016 4556 5093 4564
rect 3227 4515 3253 4523
rect 3327 4516 3373 4524
rect 3396 4524 3404 4553
rect 4056 4527 4064 4553
rect 4107 4536 4404 4544
rect 3396 4516 3413 4524
rect 3396 4504 3404 4516
rect 3747 4515 3793 4523
rect 3847 4515 3873 4523
rect 3947 4515 4013 4523
rect 4347 4515 4373 4523
rect 4396 4524 4404 4536
rect 4396 4516 4473 4524
rect 4487 4516 4513 4524
rect 4896 4526 4904 4553
rect 4956 4527 4964 4554
rect 5016 4527 5024 4556
rect 5187 4556 5204 4564
rect 5196 4544 5204 4556
rect 5227 4556 5273 4564
rect 5287 4556 5313 4564
rect 5196 4536 5344 4544
rect 4667 4516 4693 4524
rect 4707 4515 4733 4523
rect 4827 4515 4853 4523
rect 4956 4516 4973 4527
rect 4960 4513 4973 4516
rect 5087 4516 5133 4524
rect 5336 4526 5344 4536
rect 5356 4524 5364 4554
rect 5456 4544 5464 4573
rect 5487 4556 5593 4564
rect 5713 4544 5727 4553
rect 5456 4536 5504 4544
rect 5676 4540 5727 4544
rect 5356 4516 5393 4524
rect 5496 4526 5504 4536
rect 5673 4536 5724 4540
rect 5673 4527 5687 4536
rect 5507 4516 5613 4524
rect 5796 4507 5804 4573
rect 2907 4496 3044 4504
rect 3296 4500 3404 4504
rect 3293 4496 3404 4500
rect 3293 4487 3307 4496
rect 3567 4496 3913 4504
rect 4567 4496 4633 4504
rect 5707 4496 5753 4504
rect 1276 4476 1353 4484
rect 1407 4476 1793 4484
rect 1847 4476 2293 4484
rect 2347 4476 2533 4484
rect 2707 4476 3253 4484
rect 3407 4476 3613 4484
rect 4027 4476 4173 4484
rect 4196 4476 4504 4484
rect 936 4464 944 4473
rect 767 4456 944 4464
rect 1267 4456 1493 4464
rect 1647 4456 1773 4464
rect 1796 4456 2033 4464
rect 1227 4436 1552 4444
rect 1587 4436 1653 4444
rect 1796 4444 1804 4456
rect 2167 4456 2493 4464
rect 2587 4456 2833 4464
rect 2896 4456 3953 4464
rect 2896 4447 2904 4456
rect 3967 4456 4033 4464
rect 4196 4464 4204 4476
rect 4087 4456 4204 4464
rect 4496 4464 4504 4476
rect 4767 4476 4973 4484
rect 4987 4476 5193 4484
rect 5207 4476 5393 4484
rect 4227 4456 4484 4464
rect 4496 4456 4633 4464
rect 4476 4447 4484 4456
rect 4787 4456 4833 4464
rect 4947 4456 5273 4464
rect 5387 4456 5593 4464
rect 5607 4456 5693 4464
rect 1727 4436 1804 4444
rect 1847 4436 2013 4444
rect 2067 4436 2093 4444
rect 2287 4436 2333 4444
rect 2727 4436 2892 4444
rect 2927 4436 2953 4444
rect 3007 4436 3633 4444
rect 4487 4436 4593 4444
rect 5787 4436 5813 4444
rect 747 4416 793 4424
rect 807 4416 953 4424
rect 1447 4416 1913 4424
rect 2187 4416 2393 4424
rect 2407 4416 2573 4424
rect 2627 4416 2753 4424
rect 2867 4416 3113 4424
rect 3307 4416 3493 4424
rect 3587 4416 3652 4424
rect 3687 4416 4293 4424
rect 4527 4416 4833 4424
rect 5247 4416 5353 4424
rect 5367 4416 5513 4424
rect 247 4396 313 4404
rect 567 4396 593 4404
rect 1507 4396 1933 4404
rect 2007 4396 2113 4404
rect 2127 4396 2253 4404
rect 2807 4396 3233 4404
rect 3287 4396 3373 4404
rect 4387 4396 4453 4404
rect 4547 4396 4573 4404
rect 5067 4396 5113 4404
rect 707 4376 773 4384
rect 1067 4376 1193 4384
rect 1207 4376 1333 4384
rect 1467 4376 1572 4384
rect 1607 4376 1853 4384
rect 1927 4376 1973 4384
rect 2687 4376 2793 4384
rect 2907 4376 3053 4384
rect 3067 4376 3153 4384
rect 3267 4376 3553 4384
rect 3607 4376 3813 4384
rect 4107 4376 4133 4384
rect 4867 4376 4893 4384
rect 4907 4376 5013 4384
rect 5327 4376 5464 4384
rect 5456 4367 5464 4376
rect 5627 4376 5653 4384
rect 147 4356 213 4364
rect 267 4356 413 4364
rect 467 4356 604 4364
rect 596 4348 604 4356
rect 1387 4356 1413 4364
rect 1776 4356 1813 4364
rect 67 4344 80 4347
rect 67 4333 84 4344
rect 347 4337 372 4345
rect 673 4344 687 4353
rect 647 4340 687 4344
rect 647 4336 684 4340
rect 696 4336 733 4344
rect 76 4306 84 4333
rect 196 4307 204 4333
rect 396 4307 404 4333
rect 287 4296 353 4304
rect 496 4287 504 4334
rect 596 4324 604 4334
rect 696 4324 704 4336
rect 787 4337 833 4345
rect 1056 4336 1153 4344
rect 596 4316 704 4324
rect 527 4295 553 4303
rect 667 4295 693 4303
rect 876 4287 884 4334
rect 916 4307 924 4334
rect 1056 4324 1064 4336
rect 1507 4336 1633 4344
rect 1776 4344 1784 4356
rect 1836 4356 1993 4364
rect 1647 4336 1784 4344
rect 996 4316 1064 4324
rect 1316 4324 1324 4334
rect 1316 4316 1384 4324
rect 916 4296 933 4307
rect 920 4293 933 4296
rect 996 4306 1004 4316
rect 1147 4296 1213 4304
rect 1227 4295 1253 4303
rect 1376 4287 1384 4316
rect 1836 4306 1844 4356
rect 2136 4356 2233 4364
rect 2027 4337 2073 4345
rect 1916 4307 1924 4333
rect 1547 4300 1644 4304
rect 1547 4296 1647 4300
rect 1633 4287 1647 4296
rect 2136 4306 2144 4356
rect 2547 4356 2664 4364
rect 2327 4337 2453 4345
rect 2467 4337 2493 4345
rect 2287 4296 2353 4304
rect 2427 4296 2553 4304
rect 2616 4304 2624 4333
rect 2656 4306 2664 4356
rect 2736 4356 2953 4364
rect 2696 4324 2704 4353
rect 2736 4324 2744 4356
rect 2967 4356 3033 4364
rect 3467 4356 3533 4364
rect 3927 4356 4124 4364
rect 2676 4316 2704 4324
rect 2716 4316 2744 4324
rect 2567 4296 2624 4304
rect 2676 4287 2684 4316
rect 2716 4304 2724 4316
rect 2836 4307 2844 4334
rect 2887 4336 2913 4344
rect 3253 4344 3267 4352
rect 3227 4340 3267 4344
rect 3227 4336 3264 4340
rect 3347 4336 3433 4344
rect 3487 4337 3513 4345
rect 3627 4336 3733 4344
rect 3787 4336 3853 4344
rect 4116 4344 4124 4356
rect 4167 4356 4413 4364
rect 4460 4364 4473 4367
rect 4456 4353 4473 4364
rect 4516 4356 4553 4364
rect 3907 4336 3944 4344
rect 4116 4336 4284 4344
rect 3293 4324 3307 4333
rect 3167 4320 3307 4324
rect 3167 4316 3304 4320
rect 3936 4307 3944 4336
rect 4276 4324 4284 4336
rect 4456 4347 4464 4353
rect 4307 4336 4353 4344
rect 4493 4324 4507 4333
rect 4276 4320 4507 4324
rect 4276 4316 4504 4320
rect 2707 4296 2724 4304
rect 2747 4295 2773 4303
rect 2836 4296 2853 4307
rect 2840 4293 2853 4296
rect 3007 4296 3293 4304
rect 3556 4300 3633 4304
rect 3553 4296 3633 4300
rect 3553 4287 3567 4296
rect 3647 4296 3753 4304
rect 4087 4296 4253 4304
rect 4396 4306 4404 4316
rect 4516 4304 4524 4356
rect 4607 4356 4653 4364
rect 4667 4356 4824 4364
rect 4816 4348 4824 4356
rect 4847 4356 5033 4364
rect 5467 4356 5504 4364
rect 4827 4336 4933 4344
rect 4487 4296 4524 4304
rect 4627 4296 4653 4304
rect 2807 4276 2893 4284
rect 3127 4276 3253 4284
rect 3267 4276 3333 4284
rect 3387 4276 3493 4284
rect 3687 4276 3713 4284
rect 3887 4276 3973 4284
rect 4167 4276 4233 4284
rect 4247 4276 4313 4284
rect 4716 4284 4724 4334
rect 5327 4344 5340 4347
rect 5327 4333 5344 4344
rect 5407 4337 5433 4345
rect 5336 4306 5344 4333
rect 5496 4306 5504 4356
rect 5627 4336 5684 4344
rect 5676 4306 5684 4336
rect 5207 4296 5333 4304
rect 4607 4276 4724 4284
rect 4907 4276 4953 4284
rect 47 4256 233 4264
rect 487 4256 613 4264
rect 1327 4256 1433 4264
rect 1607 4256 1793 4264
rect 1807 4256 2193 4264
rect 2656 4256 2933 4264
rect 2656 4247 2664 4256
rect 3107 4256 3193 4264
rect 3527 4256 3752 4264
rect 3787 4256 3833 4264
rect 4007 4256 4073 4264
rect 4127 4256 4273 4264
rect 4347 4256 4553 4264
rect 4727 4256 4913 4264
rect 5247 4256 5373 4264
rect 5387 4256 5633 4264
rect 727 4236 1033 4244
rect 1367 4236 1473 4244
rect 1587 4236 1713 4244
rect 1727 4236 1933 4244
rect 2007 4236 2233 4244
rect 2247 4236 2593 4244
rect 2607 4236 2653 4244
rect 3227 4236 3433 4244
rect 3507 4236 4593 4244
rect 4647 4236 4693 4244
rect 5327 4236 5433 4244
rect 787 4216 892 4224
rect 927 4216 1033 4224
rect 1187 4216 1333 4224
rect 1407 4216 1533 4224
rect 2507 4216 2713 4224
rect 2847 4216 3473 4224
rect 3547 4216 3964 4224
rect 1447 4196 1833 4204
rect 1887 4196 1973 4204
rect 2407 4196 3173 4204
rect 3227 4196 3473 4204
rect 807 4176 913 4184
rect 967 4176 1353 4184
rect 1447 4176 1553 4184
rect 1567 4176 1813 4184
rect 2396 4184 2404 4193
rect 3847 4196 3933 4204
rect 3956 4204 3964 4216
rect 4007 4216 4332 4224
rect 4367 4216 4493 4224
rect 4747 4216 5773 4224
rect 3956 4196 4073 4204
rect 4247 4196 4513 4204
rect 4567 4196 4673 4204
rect 1827 4176 2404 4184
rect 2487 4176 2793 4184
rect 2836 4176 3253 4184
rect 1867 4156 2173 4164
rect 2836 4164 2844 4176
rect 3347 4176 3453 4184
rect 3527 4176 3793 4184
rect 3807 4176 4093 4184
rect 4147 4176 4513 4184
rect 4587 4176 4713 4184
rect 5487 4176 5733 4184
rect 2247 4156 2844 4164
rect 2887 4156 2933 4164
rect 2987 4156 3013 4164
rect 3107 4156 3233 4164
rect 3287 4156 3412 4164
rect 3447 4156 3744 4164
rect 627 4136 653 4144
rect 1047 4136 1233 4144
rect 1627 4136 2013 4144
rect 2027 4136 2093 4144
rect 2147 4136 2273 4144
rect 2287 4136 2453 4144
rect 2467 4136 2673 4144
rect 2727 4136 3013 4144
rect 3118 4136 3213 4144
rect 3307 4136 3353 4144
rect 3467 4136 3553 4144
rect 3607 4136 3673 4144
rect 3736 4144 3744 4156
rect 3767 4156 3853 4164
rect 3927 4156 4053 4164
rect 4767 4156 5353 4164
rect 5467 4156 5573 4164
rect 3736 4136 3873 4144
rect 4056 4136 4233 4144
rect 287 4116 433 4124
rect 907 4116 973 4124
rect 1267 4116 1433 4124
rect 1487 4116 1593 4124
rect 1767 4116 1933 4124
rect 2567 4116 3033 4124
rect 4056 4124 4064 4136
rect 4327 4136 4393 4144
rect 4447 4136 4633 4144
rect 4647 4136 4993 4144
rect 3267 4116 4064 4124
rect 4087 4116 4133 4124
rect 4507 4116 4624 4124
rect 707 4096 773 4104
rect 887 4096 1224 4104
rect 627 4076 673 4084
rect 1216 4084 1224 4096
rect 1547 4096 1904 4104
rect 1216 4076 1453 4084
rect 1607 4076 1673 4084
rect 1687 4076 1853 4084
rect 1896 4084 1904 4096
rect 2867 4096 2953 4104
rect 3067 4096 3344 4104
rect 1896 4076 2313 4084
rect 2327 4076 2373 4084
rect 2907 4076 3104 4084
rect 3173 4086 3187 4096
rect 3336 4084 3344 4096
rect 3427 4096 3533 4104
rect 3867 4096 3944 4104
rect 3336 4076 3613 4084
rect 427 4064 440 4067
rect 427 4053 444 4064
rect 107 4037 173 4045
rect 116 4016 193 4024
rect 116 4006 124 4016
rect 236 4004 244 4034
rect 436 4007 444 4053
rect 567 4056 713 4064
rect 927 4056 993 4064
rect 1307 4056 1413 4064
rect 1487 4056 1513 4064
rect 1527 4056 1673 4064
rect 1947 4056 2073 4064
rect 2447 4056 2553 4064
rect 3047 4056 3213 4064
rect 3313 4064 3327 4073
rect 3747 4076 3833 4084
rect 3936 4084 3944 4096
rect 3987 4096 4173 4104
rect 4247 4096 4393 4104
rect 4616 4104 4624 4116
rect 4667 4116 4793 4124
rect 4616 4096 4673 4104
rect 4687 4096 5053 4104
rect 5067 4096 5113 4104
rect 5227 4096 5453 4104
rect 3936 4076 4072 4084
rect 4107 4076 4413 4084
rect 4707 4076 4973 4084
rect 5547 4076 5613 4084
rect 3227 4060 3327 4064
rect 3227 4056 3324 4060
rect 816 4007 824 4034
rect 887 4044 900 4047
rect 887 4033 904 4044
rect 1207 4037 1493 4045
rect 1727 4037 1773 4045
rect 236 3996 393 4004
rect 816 3996 833 4007
rect 820 3993 833 3996
rect 896 4006 904 4033
rect 976 4007 984 4033
rect 1016 4004 1024 4033
rect 1016 3996 1053 4004
rect 1076 4004 1084 4034
rect 1787 4037 1873 4045
rect 1900 4044 1913 4047
rect 1896 4033 1913 4044
rect 2167 4037 2233 4045
rect 2307 4036 2484 4044
rect 1896 4024 1904 4033
rect 1816 4016 1904 4024
rect 1076 3996 1093 4004
rect 1107 3996 1273 4004
rect 1816 4006 1824 4016
rect 2476 4007 2484 4036
rect 2607 4037 2633 4045
rect 2727 4037 2853 4045
rect 1527 3996 1573 4004
rect 1647 3995 1733 4003
rect 1907 3996 1953 4004
rect 2227 3995 2393 4003
rect 2667 3996 2713 4004
rect 2727 3996 2753 4004
rect 2896 4004 2904 4034
rect 3027 4036 3073 4044
rect 3180 4044 3193 4047
rect 3176 4033 3193 4044
rect 3393 4044 3407 4053
rect 3687 4056 3813 4064
rect 4247 4056 4293 4064
rect 4307 4056 4383 4064
rect 3393 4040 3453 4044
rect 3396 4036 3453 4040
rect 2976 4007 2984 4033
rect 2847 3996 2904 4004
rect 2927 3996 2944 4004
rect 547 3976 753 3984
rect 1427 3976 1453 3984
rect 2427 3976 2573 3984
rect 2936 3967 2944 3996
rect 3176 4004 3184 4033
rect 3167 3996 3184 4004
rect 3276 3987 3284 4034
rect 3513 4044 3527 4053
rect 4375 4048 4383 4056
rect 4527 4056 4733 4064
rect 4887 4056 5013 4064
rect 3513 4040 3564 4044
rect 3516 4036 3564 4040
rect 3296 4016 3473 4024
rect 3296 4006 3304 4016
rect 3347 3996 3373 4004
rect 3447 3996 3493 4004
rect 3556 4006 3564 4036
rect 3727 4037 3753 4045
rect 4027 4037 4053 4045
rect 4387 4036 4453 4044
rect 4507 4037 4653 4045
rect 4987 4037 5053 4045
rect 5067 4036 5153 4044
rect 5447 4036 5533 4044
rect 5627 4037 5653 4045
rect 3596 4007 3604 4033
rect 4256 4007 4264 4033
rect 4753 4024 4767 4033
rect 4696 4020 4767 4024
rect 4696 4016 4764 4020
rect 3887 3995 3913 4003
rect 3967 3996 4073 4004
rect 4127 3996 4173 4004
rect 4367 3995 4393 4003
rect 4696 4004 4704 4016
rect 4627 3996 4704 4004
rect 4716 3996 4733 4004
rect 3067 3976 3113 3984
rect 3187 3976 3213 3984
rect 4396 3984 4404 3992
rect 3707 3976 3904 3984
rect 4396 3976 4573 3984
rect 407 3956 493 3964
rect 807 3956 933 3964
rect 1907 3956 2093 3964
rect 2107 3956 2173 3964
rect 2447 3956 2513 3964
rect 2607 3956 2653 3964
rect 2827 3956 2873 3964
rect 3247 3956 3333 3964
rect 3507 3956 3653 3964
rect 3827 3956 3873 3964
rect 3896 3964 3904 3976
rect 4716 3984 4724 3996
rect 4747 3996 4813 4004
rect 5007 3996 5133 4004
rect 5316 4004 5324 4034
rect 5316 3996 5413 4004
rect 5567 3996 5673 4004
rect 4647 3976 4724 3984
rect 4996 3984 5004 3992
rect 4927 3976 5004 3984
rect 5307 3976 5353 3984
rect 5587 3976 5613 3984
rect 3896 3956 4013 3964
rect 4087 3956 4133 3964
rect 4227 3956 4273 3964
rect 5047 3956 5173 3964
rect 5647 3956 5713 3964
rect 67 3936 253 3944
rect 1007 3936 1173 3944
rect 1867 3936 1993 3944
rect 2007 3936 2172 3944
rect 2207 3936 2273 3944
rect 2347 3936 2513 3944
rect 2967 3936 2993 3944
rect 3007 3936 3233 3944
rect 3247 3936 3413 3944
rect 3767 3936 4293 3944
rect 4487 3936 4793 3944
rect 4867 3936 5013 3944
rect 5207 3936 5233 3944
rect 407 3916 453 3924
rect 467 3916 573 3924
rect 867 3916 913 3924
rect 1367 3916 1613 3924
rect 1787 3916 2493 3924
rect 2507 3916 2533 3924
rect 2547 3916 3253 3924
rect 3496 3916 3653 3924
rect 1327 3896 1693 3904
rect 1847 3896 2033 3904
rect 2047 3896 2113 3904
rect 2187 3896 2333 3904
rect 2907 3896 2973 3904
rect 3496 3904 3504 3916
rect 3807 3916 3993 3924
rect 4207 3916 4613 3924
rect 4636 3916 5173 3924
rect 3467 3896 3504 3904
rect 4636 3904 4644 3916
rect 5187 3916 5353 3924
rect 5367 3916 5493 3924
rect 3527 3896 4644 3904
rect 4807 3896 5053 3904
rect 5107 3896 5273 3904
rect 5787 3896 5894 3904
rect 67 3876 93 3884
rect 107 3876 353 3884
rect 607 3876 753 3884
rect 807 3876 853 3884
rect 1067 3876 1393 3884
rect 1727 3876 1853 3884
rect 1947 3876 2073 3884
rect 2607 3876 2813 3884
rect 3007 3876 3033 3884
rect 3316 3876 3433 3884
rect 167 3856 253 3864
rect 547 3856 613 3864
rect 687 3856 833 3864
rect 847 3856 953 3864
rect 1276 3856 1513 3864
rect 1276 3847 1284 3856
rect 1747 3856 1793 3864
rect 1927 3856 2473 3864
rect 2587 3856 2893 3864
rect 3316 3864 3324 3876
rect 3647 3876 3873 3884
rect 3887 3876 4193 3884
rect 4707 3876 4873 3884
rect 5087 3876 5513 3884
rect 5647 3876 5793 3884
rect 2947 3856 3324 3864
rect 3547 3856 3713 3864
rect 3907 3856 3993 3864
rect 4247 3856 4353 3864
rect 4727 3856 4893 3864
rect 5007 3856 5093 3864
rect 5147 3856 5313 3864
rect 227 3836 273 3844
rect 287 3836 313 3844
rect 1187 3836 1273 3844
rect 1576 3836 1693 3844
rect 367 3817 433 3825
rect 616 3804 624 3814
rect 766 3813 767 3820
rect 787 3816 813 3824
rect 876 3816 953 3824
rect 616 3796 673 3804
rect 753 3804 767 3813
rect 753 3800 844 3804
rect 756 3796 844 3800
rect 836 3786 844 3796
rect 876 3786 884 3816
rect 1087 3816 1133 3824
rect 1247 3824 1260 3827
rect 1247 3813 1264 3824
rect 1387 3816 1444 3824
rect 1256 3804 1264 3813
rect 1256 3796 1304 3804
rect 147 3775 173 3783
rect 247 3776 333 3784
rect 547 3775 593 3783
rect 1296 3786 1304 3796
rect 1436 3786 1444 3816
rect 1496 3787 1504 3813
rect 927 3776 1013 3784
rect 507 3756 673 3764
rect 687 3756 773 3764
rect 1013 3764 1093 3772
rect 1367 3775 1393 3783
rect 1576 3786 1584 3836
rect 2207 3836 2353 3844
rect 2847 3836 2993 3844
rect 3127 3836 3173 3844
rect 3347 3836 3453 3844
rect 3536 3836 3793 3844
rect 1616 3820 1693 3824
rect 1613 3816 1693 3820
rect 1613 3807 1627 3816
rect 1716 3816 1753 3824
rect 1716 3786 1724 3816
rect 1807 3816 1864 3824
rect 1856 3787 1864 3816
rect 1647 3775 1673 3783
rect 1936 3786 1944 3833
rect 1967 3816 2084 3824
rect 2076 3786 2084 3816
rect 2387 3817 2433 3825
rect 2487 3817 2553 3825
rect 2567 3816 2664 3824
rect 2656 3804 2664 3816
rect 2727 3816 2773 3824
rect 2656 3796 2704 3804
rect 2696 3786 2704 3796
rect 3016 3787 3024 3814
rect 3187 3817 3233 3825
rect 3016 3776 3033 3787
rect 3020 3773 3033 3776
rect 3256 3786 3264 3833
rect 3296 3816 3393 3824
rect 3296 3804 3304 3816
rect 3536 3824 3544 3836
rect 4067 3836 4153 3844
rect 4427 3836 4633 3844
rect 4647 3836 4673 3844
rect 5427 3836 5633 3844
rect 5827 3844 5840 3847
rect 5827 3833 5844 3844
rect 3447 3816 3544 3824
rect 3776 3816 3813 3824
rect 3556 3804 3564 3814
rect 3296 3796 3544 3804
rect 3556 3800 3584 3804
rect 3556 3796 3587 3800
rect 3296 3786 3304 3796
rect 3536 3786 3544 3796
rect 3573 3787 3587 3796
rect 3776 3787 3784 3816
rect 3887 3816 4033 3824
rect 4147 3816 4193 3824
rect 4267 3816 4333 3824
rect 4467 3816 4604 3824
rect 4596 3786 4604 3816
rect 4847 3816 4864 3824
rect 4856 3787 4864 3816
rect 4887 3816 4944 3824
rect 4936 3804 4944 3816
rect 4967 3816 5093 3824
rect 5213 3824 5227 3833
rect 5213 3820 5244 3824
rect 5216 3816 5244 3820
rect 4936 3796 5124 3804
rect 3847 3775 3913 3783
rect 4087 3775 4113 3783
rect 4167 3776 4233 3784
rect 4307 3776 4393 3784
rect 4856 3776 4873 3787
rect 4860 3773 4873 3776
rect 4936 3786 4944 3796
rect 5116 3786 5124 3796
rect 4987 3776 5073 3784
rect 5187 3775 5213 3783
rect 5236 3767 5244 3816
rect 5256 3804 5264 3833
rect 5287 3816 5384 3824
rect 5256 3800 5344 3804
rect 5256 3796 5347 3800
rect 5333 3787 5347 3796
rect 5376 3786 5384 3816
rect 5687 3816 5713 3824
rect 5736 3816 5753 3824
rect 5596 3787 5604 3813
rect 5736 3804 5744 3816
rect 5696 3800 5744 3804
rect 5693 3796 5744 3800
rect 5693 3787 5707 3796
rect 5796 3767 5804 3814
rect 5836 3787 5844 3833
rect 5827 3776 5844 3787
rect 5827 3773 5840 3776
rect 2027 3756 2253 3764
rect 2507 3756 2573 3764
rect 2627 3756 2773 3764
rect 2967 3756 3093 3764
rect 3227 3756 3373 3764
rect 3647 3756 4533 3764
rect 5327 3756 5413 3764
rect 1267 3736 1433 3744
rect 1607 3736 1813 3744
rect 1827 3736 1873 3744
rect 1927 3736 1973 3744
rect 2496 3744 2504 3753
rect 1996 3736 2504 3744
rect 1167 3716 1533 3724
rect 1547 3716 1693 3724
rect 1996 3724 2004 3736
rect 2807 3736 2853 3744
rect 3387 3736 3493 3744
rect 4107 3736 4172 3744
rect 4207 3736 4473 3744
rect 4567 3736 4693 3744
rect 1807 3716 2004 3724
rect 2127 3716 2784 3724
rect 2776 3704 2784 3716
rect 2887 3716 2993 3724
rect 3047 3716 3233 3724
rect 4887 3716 5333 3724
rect 5347 3716 5613 3724
rect 5627 3716 5753 3724
rect 2876 3704 2884 3713
rect 2776 3696 2884 3704
rect 3087 3696 3173 3704
rect 4047 3696 4293 3704
rect 4367 3696 4473 3704
rect 4487 3696 4733 3704
rect 4787 3696 4953 3704
rect 5827 3704 5840 3707
rect 5827 3693 5844 3704
rect 987 3676 1213 3684
rect 1227 3676 1613 3684
rect 1727 3676 2193 3684
rect 2367 3676 2733 3684
rect 2907 3676 3012 3684
rect 3047 3676 3633 3684
rect 4387 3676 4613 3684
rect 5747 3676 5813 3684
rect 1887 3656 3244 3664
rect 67 3636 353 3644
rect 1507 3636 1553 3644
rect 1567 3636 1633 3644
rect 2047 3636 2133 3644
rect 2367 3636 2513 3644
rect 2667 3636 2833 3644
rect 3067 3636 3093 3644
rect 3236 3644 3244 3656
rect 4067 3656 4313 3664
rect 3236 3636 3333 3644
rect 3347 3636 3393 3644
rect 3447 3636 3673 3644
rect 4167 3636 4353 3644
rect 4547 3636 4813 3644
rect 5547 3636 5673 3644
rect 5836 3644 5844 3693
rect 5727 3636 5844 3644
rect 107 3616 573 3624
rect 1307 3616 1893 3624
rect 2947 3616 2973 3624
rect 2987 3616 3133 3624
rect 3227 3616 3693 3624
rect 3707 3616 4033 3624
rect 4327 3616 4433 3624
rect 4987 3616 5053 3624
rect 5067 3616 5133 3624
rect 47 3596 73 3604
rect 87 3596 593 3604
rect 647 3596 2413 3604
rect 3027 3596 3113 3604
rect 3127 3596 3152 3604
rect 3187 3596 3433 3604
rect 3567 3596 3793 3604
rect 3807 3596 3893 3604
rect 4247 3596 4513 3604
rect 4647 3596 4673 3604
rect 5607 3596 5673 3604
rect 5687 3596 5733 3604
rect 427 3576 473 3584
rect 2087 3576 2113 3584
rect 2467 3576 2533 3584
rect 2767 3576 2873 3584
rect 2887 3576 2913 3584
rect 3007 3576 3293 3584
rect 3467 3576 4013 3584
rect 4636 3576 4793 3584
rect 4636 3567 4644 3576
rect 4867 3576 4913 3584
rect 5407 3576 5453 3584
rect 27 3556 93 3564
rect 187 3556 233 3564
rect 587 3556 633 3564
rect 687 3556 773 3564
rect 867 3556 993 3564
rect 1007 3556 1053 3564
rect 1387 3556 1593 3564
rect 1976 3556 2053 3564
rect 127 3536 284 3544
rect 276 3528 284 3536
rect 436 3536 553 3544
rect 436 3528 444 3536
rect 827 3536 873 3544
rect 1476 3536 1673 3544
rect -74 3516 13 3524
rect 287 3517 433 3525
rect 487 3516 524 3524
rect -74 3476 13 3484
rect 196 3484 204 3514
rect 107 3476 204 3484
rect 516 3484 524 3516
rect 667 3517 733 3525
rect 907 3516 1033 3524
rect 1036 3504 1044 3514
rect 1307 3516 1333 3524
rect 1476 3527 1484 3536
rect 1976 3544 1984 3556
rect 2307 3556 2433 3564
rect 3507 3556 3593 3564
rect 3687 3556 3713 3564
rect 4127 3556 4153 3564
rect 4167 3556 4193 3564
rect 4307 3556 4633 3564
rect 5007 3556 5033 3564
rect 5047 3556 5093 3564
rect 5267 3556 5593 3564
rect 1947 3536 1984 3544
rect 2127 3536 2184 3544
rect 1780 3524 1793 3527
rect 1036 3496 1113 3504
rect 516 3476 573 3484
rect 627 3476 653 3484
rect 1287 3476 1493 3484
rect 1516 3484 1524 3514
rect 1776 3513 1793 3524
rect 1776 3486 1784 3513
rect 1816 3496 1893 3504
rect 1816 3486 1824 3496
rect 1916 3487 1924 3513
rect 1996 3487 2004 3514
rect 2176 3524 2184 3536
rect 5387 3536 5413 3544
rect 5727 3544 5740 3547
rect 5727 3533 5744 3544
rect 2176 3516 2253 3524
rect 2267 3516 2373 3524
rect 2427 3516 2493 3524
rect 2587 3517 2613 3525
rect 2667 3517 2713 3525
rect 2887 3516 2993 3524
rect 2076 3487 2084 3513
rect 2156 3487 2164 3514
rect 2256 3504 2264 3514
rect 2236 3496 2264 3504
rect 2796 3504 2804 3514
rect 3267 3517 3413 3525
rect 2796 3496 2953 3504
rect 2236 3487 2244 3496
rect 3116 3487 3124 3513
rect 1516 3476 1733 3484
rect 1996 3476 2013 3487
rect 2000 3473 2013 3476
rect 2156 3476 2173 3487
rect 2160 3473 2173 3476
rect 2227 3476 2244 3487
rect 2227 3473 2240 3476
rect 2287 3475 2313 3483
rect 2407 3480 2444 3484
rect 2407 3476 2447 3480
rect 407 3456 433 3464
rect 876 3464 884 3472
rect 2433 3467 2447 3476
rect 2987 3475 3033 3483
rect 3327 3476 3372 3484
rect 3456 3484 3464 3514
rect 3596 3504 3604 3514
rect 3787 3517 3833 3525
rect 3987 3516 4333 3524
rect 4360 3524 4373 3527
rect 4356 3513 4373 3524
rect 4427 3516 4453 3524
rect 4476 3516 4673 3524
rect 4356 3504 4364 3513
rect 4476 3504 4484 3516
rect 4727 3517 4753 3525
rect 4856 3516 5033 3524
rect 3596 3496 3664 3504
rect 3407 3476 3464 3484
rect 3656 3484 3664 3496
rect 4276 3496 4364 3504
rect 4396 3496 4484 3504
rect 3656 3476 3693 3484
rect 3747 3476 3773 3484
rect 4276 3486 4284 3496
rect 4396 3486 4404 3496
rect 4527 3476 4573 3484
rect 4587 3475 4613 3483
rect 4856 3484 4864 3516
rect 5047 3516 5173 3524
rect 5347 3516 5433 3524
rect 5296 3504 5304 3514
rect 5476 3504 5484 3514
rect 5556 3504 5564 3514
rect 5646 3513 5647 3520
rect 5667 3516 5693 3524
rect 5633 3504 5647 3513
rect 5736 3504 5744 3533
rect 5276 3496 5564 3504
rect 5616 3500 5647 3504
rect 5616 3496 5643 3500
rect 5716 3496 5744 3504
rect 4827 3476 4864 3484
rect 4987 3475 5013 3483
rect 5276 3484 5284 3496
rect 5616 3486 5624 3496
rect 5067 3476 5284 3484
rect 5327 3475 5373 3483
rect 5387 3476 5453 3484
rect 5527 3475 5573 3483
rect 876 3456 1013 3464
rect 1367 3456 1493 3464
rect 1507 3456 1533 3464
rect 1627 3456 1673 3464
rect 1836 3456 1873 3464
rect 227 3436 253 3444
rect 687 3436 733 3444
rect 1127 3436 1193 3444
rect 1427 3436 1453 3444
rect 1836 3444 1844 3456
rect 2067 3456 2133 3464
rect 2687 3456 2893 3464
rect 3587 3456 3633 3464
rect 3807 3456 3833 3464
rect 4667 3456 4753 3464
rect 5107 3456 5153 3464
rect 5716 3464 5724 3496
rect 5756 3487 5764 3513
rect 5647 3456 5724 3464
rect 1727 3436 1844 3444
rect 1887 3436 2144 3444
rect 2007 3416 2073 3424
rect 2136 3424 2144 3436
rect 2247 3436 2333 3444
rect 2347 3436 2373 3444
rect 2627 3436 2713 3444
rect 2967 3436 3152 3444
rect 3187 3436 3393 3444
rect 3687 3436 3893 3444
rect 4187 3436 4213 3444
rect 4227 3436 4313 3444
rect 4967 3436 5133 3444
rect 5407 3436 5533 3444
rect 2136 3416 2573 3424
rect 2587 3416 2773 3424
rect 2907 3416 3953 3424
rect 4007 3416 4193 3424
rect 4567 3416 4653 3424
rect 4667 3416 4773 3424
rect 27 3396 213 3404
rect 1147 3396 1533 3404
rect 1547 3396 1733 3404
rect 1787 3396 1853 3404
rect 2107 3396 2493 3404
rect 3207 3396 3273 3404
rect 3447 3396 3613 3404
rect 3627 3396 4733 3404
rect 4747 3396 4893 3404
rect 4907 3396 5053 3404
rect 767 3376 1753 3384
rect 1807 3376 1873 3384
rect 1927 3376 2073 3384
rect 2147 3376 2213 3384
rect 2807 3376 2853 3384
rect 2867 3376 3144 3384
rect 27 3356 1613 3364
rect 2167 3356 2193 3364
rect 2367 3356 2633 3364
rect 2887 3356 3073 3364
rect 3136 3364 3144 3376
rect 3707 3376 3793 3384
rect 3807 3376 3993 3384
rect 4067 3376 4233 3384
rect 3136 3356 3173 3364
rect 3267 3356 3553 3364
rect 4487 3356 4573 3364
rect 5247 3356 5704 3364
rect 67 3336 113 3344
rect 167 3336 193 3344
rect 267 3336 573 3344
rect 847 3336 1173 3344
rect 1887 3336 1953 3344
rect 2487 3336 2513 3344
rect 2607 3336 2673 3344
rect 2847 3336 3193 3344
rect 3387 3336 3453 3344
rect 3607 3336 3653 3344
rect 4027 3336 4113 3344
rect 4127 3336 4173 3344
rect 4327 3336 4353 3344
rect 4467 3336 4593 3344
rect 4607 3336 4713 3344
rect -74 3316 13 3324
rect 1247 3316 1273 3324
rect 1527 3316 1553 3324
rect 1847 3316 2033 3324
rect 2047 3316 2093 3324
rect 2467 3316 2513 3324
rect 2527 3316 2713 3324
rect 4047 3316 4153 3324
rect 47 3297 73 3305
rect 407 3297 453 3305
rect 527 3296 593 3304
rect 787 3296 893 3304
rect 947 3296 993 3304
rect -74 3276 13 3284
rect 607 3255 633 3263
rect -74 3236 33 3244
rect 656 3244 664 3294
rect 1007 3296 1033 3304
rect 1107 3297 1293 3305
rect 1347 3296 1433 3304
rect 1727 3296 1744 3304
rect 1496 3267 1504 3293
rect 1633 3284 1647 3293
rect 1633 3280 1664 3284
rect 1636 3276 1664 3280
rect 687 3256 753 3264
rect 967 3255 1093 3263
rect 1207 3256 1273 3264
rect 1656 3266 1664 3276
rect 1547 3256 1653 3264
rect 1676 3247 1684 3294
rect 1736 3267 1744 3296
rect 1807 3296 1913 3304
rect 1767 3284 1780 3287
rect 1767 3273 1784 3284
rect 1776 3264 1784 3273
rect 1856 3267 1864 3296
rect 1927 3297 2153 3305
rect 2476 3296 2573 3304
rect 2436 3284 2444 3294
rect 2476 3284 2484 3296
rect 2927 3296 2972 3304
rect 2993 3304 3007 3313
rect 2993 3300 3033 3304
rect 2996 3296 3033 3300
rect 3207 3297 3233 3305
rect 3327 3296 3353 3304
rect 2436 3276 2753 3284
rect 1776 3256 1813 3264
rect 2147 3256 2173 3264
rect 2487 3255 2653 3263
rect 2707 3256 2813 3264
rect 2836 3264 2844 3293
rect 2827 3256 2844 3264
rect 3076 3264 3084 3294
rect 2947 3256 3084 3264
rect 3247 3256 3273 3264
rect 3416 3264 3424 3294
rect 3506 3293 3507 3300
rect 3527 3296 3673 3304
rect 3727 3296 3773 3304
rect 3907 3296 3953 3304
rect 3493 3284 3507 3293
rect 3493 3280 3584 3284
rect 3496 3276 3584 3280
rect 3576 3266 3584 3276
rect 4036 3267 4044 3313
rect 4127 3296 4164 3304
rect 3347 3256 3424 3264
rect 3747 3255 3893 3263
rect 4076 3264 4084 3293
rect 4156 3267 4164 3296
rect 4187 3296 4224 3304
rect 4216 3267 4224 3296
rect 4433 3304 4447 3313
rect 4797 3316 4933 3324
rect 4797 3308 4805 3316
rect 5127 3316 5153 3324
rect 4407 3300 4447 3304
rect 4407 3296 4444 3300
rect 4276 3284 4284 3294
rect 4356 3284 4364 3294
rect 4560 3304 4573 3307
rect 4487 3296 4524 3304
rect 4276 3280 4304 3284
rect 4276 3276 4307 3280
rect 4356 3276 4453 3284
rect 4293 3267 4307 3276
rect 4076 3256 4093 3264
rect 496 3236 664 3244
rect 496 3227 504 3236
rect 2107 3236 2513 3244
rect 3127 3236 3384 3244
rect 487 3216 504 3227
rect 487 3213 500 3216
rect 547 3216 673 3224
rect 747 3216 1253 3224
rect 1447 3216 1533 3224
rect 1707 3216 1853 3224
rect 2627 3216 2953 3224
rect 3067 3216 3173 3224
rect 3187 3216 3253 3224
rect 3376 3224 3384 3236
rect 3436 3244 3444 3252
rect 3407 3236 3444 3244
rect 4076 3244 4084 3256
rect 4156 3256 4173 3267
rect 4160 3253 4173 3256
rect 4516 3266 4524 3296
rect 4556 3293 4573 3304
rect 4707 3296 4793 3304
rect 4556 3266 4564 3293
rect 4607 3255 4633 3263
rect 4736 3247 4744 3296
rect 4847 3296 4893 3304
rect 4987 3296 5013 3304
rect 5107 3296 5213 3304
rect 5267 3296 5513 3304
rect 5527 3296 5593 3304
rect 5636 3284 5644 3333
rect 5660 3304 5673 3307
rect 5616 3276 5644 3284
rect 5656 3293 5673 3304
rect 4827 3256 4913 3264
rect 5027 3255 5073 3263
rect 5167 3255 5233 3263
rect 3967 3236 4084 3244
rect 4327 3236 4373 3244
rect 5387 3236 5533 3244
rect 5616 3244 5624 3276
rect 5656 3266 5664 3293
rect 5696 3284 5704 3356
rect 5713 3304 5727 3313
rect 5713 3300 5773 3304
rect 5716 3296 5773 3300
rect 5696 3276 5764 3284
rect 5756 3266 5764 3276
rect 5616 3240 5644 3244
rect 5616 3236 5647 3240
rect 5633 3227 5647 3236
rect 5787 3236 5894 3244
rect 3376 3216 3613 3224
rect 4107 3216 4253 3224
rect 4427 3216 4773 3224
rect 4787 3216 4953 3224
rect 347 3196 433 3204
rect 447 3196 1413 3204
rect 1567 3196 2244 3204
rect 2236 3187 2244 3196
rect 2747 3196 2853 3204
rect 3287 3196 3553 3204
rect 3647 3196 3773 3204
rect 3916 3196 4013 3204
rect 1827 3176 1993 3184
rect 2247 3176 2893 3184
rect 2967 3176 3793 3184
rect 3916 3184 3924 3196
rect 4467 3196 4573 3204
rect 5207 3196 5293 3204
rect 5487 3196 5773 3204
rect 3867 3176 3924 3184
rect 4187 3176 4253 3184
rect 4907 3176 5113 3184
rect 5227 3176 5894 3184
rect 1627 3156 2213 3164
rect 2487 3156 2533 3164
rect 2927 3156 3193 3164
rect 3627 3156 3933 3164
rect 3947 3156 4053 3164
rect 4167 3156 4413 3164
rect 267 3136 493 3144
rect 1367 3136 1573 3144
rect 2027 3136 2073 3144
rect 2087 3136 2253 3144
rect 2267 3136 2693 3144
rect 2867 3136 3352 3144
rect 3387 3136 5413 3144
rect 5487 3136 5573 3144
rect 27 3116 1553 3124
rect 1867 3116 1933 3124
rect 1947 3116 1972 3124
rect 2007 3116 2133 3124
rect 2227 3116 2433 3124
rect 2507 3116 3393 3124
rect 4007 3116 4033 3124
rect 4047 3116 4133 3124
rect 4267 3116 4393 3124
rect 4707 3116 4733 3124
rect 5027 3116 5373 3124
rect 227 3096 1753 3104
rect 2387 3096 2912 3104
rect 2947 3096 3133 3104
rect 3147 3096 3333 3104
rect 3347 3096 3413 3104
rect 3427 3096 3573 3104
rect 3707 3096 3853 3104
rect 4207 3096 5613 3104
rect 67 3076 173 3084
rect 247 3076 473 3084
rect 1247 3076 1453 3084
rect 1547 3076 1873 3084
rect 2067 3076 2093 3084
rect 2267 3076 2353 3084
rect 3007 3076 3153 3084
rect 4507 3076 4713 3084
rect 1267 3056 1724 3064
rect 87 3036 213 3044
rect 307 3036 373 3044
rect 467 3036 1133 3044
rect 1387 3036 1553 3044
rect 1716 3044 1724 3056
rect 1987 3064 2000 3067
rect 1987 3053 2004 3064
rect 2127 3056 2333 3064
rect 2407 3056 3493 3064
rect 3667 3056 3913 3064
rect 3927 3056 4173 3064
rect 5267 3056 5493 3064
rect 1716 3036 1953 3044
rect 1587 3016 1693 3024
rect 1707 3016 1973 3024
rect 287 2997 373 3005
rect 116 2964 124 2994
rect 216 2984 224 2994
rect 216 2976 244 2984
rect 116 2956 153 2964
rect 236 2947 244 2976
rect 316 2967 324 2997
rect 627 2996 693 3004
rect 1047 2997 1113 3005
rect 1167 2996 1373 3004
rect 1487 2997 1513 3005
rect 1036 2984 1044 2994
rect 936 2976 1044 2984
rect 936 2966 944 2976
rect 547 2956 633 2964
rect 747 2955 873 2963
rect 987 2955 1053 2963
rect 1467 2955 1533 2963
rect 1587 2955 1653 2963
rect 1736 2964 1744 2993
rect 1996 2967 2004 3053
rect 2636 3040 3013 3044
rect 2633 3036 3013 3040
rect 2633 3027 2647 3036
rect 3667 3036 3733 3044
rect 3787 3036 3833 3044
rect 4427 3036 4653 3044
rect 5047 3036 5293 3044
rect 2176 3016 2324 3024
rect 2176 3008 2184 3016
rect 2316 3004 2324 3016
rect 3327 3016 3533 3024
rect 3807 3016 3873 3024
rect 4027 3016 4113 3024
rect 4827 3016 4853 3024
rect 5436 3016 5513 3024
rect 2316 2996 2333 3004
rect 2707 2996 2893 3004
rect 2096 2967 2104 2993
rect 2176 2967 2184 2994
rect 1727 2956 1793 2964
rect 2167 2956 2184 2967
rect 2167 2953 2180 2956
rect 2296 2964 2304 2994
rect 2896 2967 2904 2994
rect 3236 2984 3244 2994
rect 3427 3004 3440 3007
rect 3427 2993 3444 3004
rect 3567 2997 3693 3005
rect 3847 2996 3944 3004
rect 3236 2976 3264 2984
rect 2207 2956 2304 2964
rect 2327 2955 2373 2963
rect 2467 2960 2784 2964
rect 2467 2956 2787 2960
rect 2773 2947 2787 2956
rect 2887 2956 2904 2967
rect 2887 2953 2900 2956
rect 3256 2964 3264 2976
rect 3436 2966 3444 2993
rect 3087 2956 3244 2964
rect 3256 2956 3333 2964
rect 236 2936 253 2947
rect 240 2933 253 2936
rect 1767 2936 2113 2944
rect 2827 2936 3013 2944
rect 3236 2944 3244 2956
rect 3496 2964 3504 2994
rect 3936 2984 3944 2996
rect 4047 2996 4104 3004
rect 3993 2984 4007 2993
rect 3936 2980 4007 2984
rect 4096 2984 4104 2996
rect 4196 2984 4204 3013
rect 5436 3008 5444 3016
rect 4227 2996 4273 3004
rect 4327 2997 4373 3005
rect 4487 2997 4533 3005
rect 4787 2996 4873 3004
rect 4887 2997 4913 3005
rect 4967 2996 5073 3004
rect 5100 3004 5113 3007
rect 5096 2993 5113 3004
rect 5247 2996 5433 3004
rect 5747 2996 5894 3004
rect 3936 2976 4004 2980
rect 4096 2976 4184 2984
rect 4196 2976 4224 2984
rect 3936 2966 3944 2976
rect 3496 2956 3593 2964
rect 4087 2955 4133 2963
rect 4176 2964 4184 2976
rect 4176 2956 4193 2964
rect 4216 2947 4224 2976
rect 4407 2956 4473 2964
rect 4527 2956 4633 2964
rect 4687 2955 4733 2963
rect 4987 2956 5033 2964
rect 5096 2966 5104 2993
rect 5367 2955 5393 2963
rect 5467 2956 5533 2964
rect 5667 2955 5693 2963
rect 3236 2936 3273 2944
rect 4127 2936 4153 2944
rect 4367 2936 4453 2944
rect 5093 2944 5107 2952
rect 4807 2936 5107 2944
rect 5767 2936 5813 2944
rect 147 2916 233 2924
rect 507 2916 773 2924
rect 867 2916 993 2924
rect 1007 2916 1213 2924
rect 1527 2916 1893 2924
rect 1967 2916 2393 2924
rect 3227 2916 3373 2924
rect 3827 2916 4013 2924
rect 4487 2916 4773 2924
rect 4827 2916 4873 2924
rect 4887 2916 4933 2924
rect 4987 2916 5013 2924
rect 5247 2916 5353 2924
rect 547 2896 673 2904
rect 1547 2896 1773 2904
rect 3727 2896 4233 2904
rect 4247 2896 4293 2904
rect 4967 2896 5484 2904
rect 327 2876 353 2884
rect 607 2876 693 2884
rect 1987 2876 2453 2884
rect 2527 2876 3113 2884
rect 3487 2876 4093 2884
rect 5267 2876 5453 2884
rect 5476 2884 5484 2896
rect 5587 2896 5673 2904
rect 5476 2876 5613 2884
rect 247 2856 413 2864
rect 1147 2856 1353 2864
rect 1807 2856 2353 2864
rect 2367 2856 2413 2864
rect 2587 2856 2633 2864
rect 4827 2856 4893 2864
rect 5087 2856 5133 2864
rect 5527 2856 5593 2864
rect 587 2836 693 2844
rect 1427 2836 1513 2844
rect 1527 2836 1793 2844
rect 2047 2836 2253 2844
rect 2867 2836 3133 2844
rect 3407 2836 3633 2844
rect 3867 2836 3933 2844
rect 3987 2836 4193 2844
rect 4267 2836 4513 2844
rect 4567 2836 5053 2844
rect 107 2816 132 2824
rect 167 2816 393 2824
rect 407 2816 493 2824
rect 507 2816 813 2824
rect 887 2816 953 2824
rect 967 2816 1013 2824
rect 1027 2816 1293 2824
rect 1376 2816 1413 2824
rect 647 2796 793 2804
rect 807 2796 833 2804
rect 47 2776 93 2784
rect 120 2784 133 2787
rect 116 2773 133 2784
rect 327 2776 384 2784
rect 116 2746 124 2773
rect 376 2747 384 2776
rect 427 2784 440 2787
rect 480 2784 493 2787
rect 427 2773 444 2784
rect 207 2736 293 2744
rect 436 2746 444 2773
rect 476 2773 493 2784
rect 667 2776 733 2784
rect 827 2776 864 2784
rect 476 2746 484 2773
rect 533 2764 547 2773
rect 533 2760 564 2764
rect 536 2756 564 2760
rect 556 2746 564 2756
rect 716 2756 793 2764
rect 716 2746 724 2756
rect 856 2746 864 2776
rect 887 2776 932 2784
rect 967 2784 980 2787
rect 967 2773 984 2784
rect 1047 2776 1113 2784
rect 1167 2777 1193 2785
rect 976 2746 984 2773
rect 607 2735 653 2743
rect 1207 2736 1273 2744
rect 1016 2707 1024 2732
rect 87 2696 513 2704
rect 767 2696 893 2704
rect 1007 2696 1024 2707
rect 1007 2693 1020 2696
rect 1047 2696 1133 2704
rect 1376 2687 1384 2816
rect 2147 2816 2213 2824
rect 2427 2816 3353 2824
rect 4007 2816 4113 2824
rect 4307 2816 4373 2824
rect 4627 2816 4793 2824
rect 4847 2816 5033 2824
rect 5127 2816 5213 2824
rect 5327 2816 5513 2824
rect 5527 2816 5653 2824
rect 1507 2796 1713 2804
rect 2027 2796 2093 2804
rect 3667 2796 3713 2804
rect 3887 2796 3913 2804
rect 4207 2796 4573 2804
rect 4587 2796 4713 2804
rect 5067 2796 5253 2804
rect 1607 2777 1653 2785
rect 1807 2776 2033 2784
rect 2087 2776 2153 2784
rect 2767 2777 2813 2785
rect 2256 2764 2264 2774
rect 2827 2777 3073 2785
rect 3087 2776 3193 2784
rect 3507 2777 3533 2785
rect 1787 2756 2264 2764
rect 3456 2764 3464 2774
rect 3547 2777 3573 2785
rect 3596 2776 3613 2784
rect 3596 2764 3604 2776
rect 4047 2776 4073 2784
rect 4167 2776 4244 2784
rect 3456 2760 3644 2764
rect 3456 2756 3647 2760
rect 3633 2747 3647 2756
rect 3676 2747 3684 2773
rect 4113 2764 4127 2773
rect 4236 2764 4244 2776
rect 4267 2776 4473 2784
rect 4767 2776 5013 2784
rect 5167 2776 5184 2784
rect 4113 2760 4184 2764
rect 4116 2756 4184 2760
rect 4236 2756 4393 2764
rect 1487 2735 1513 2743
rect 1747 2736 1953 2744
rect 2027 2735 2053 2743
rect 2167 2735 2193 2743
rect 2367 2736 2393 2744
rect 2547 2736 2833 2744
rect 2847 2736 2873 2744
rect 3187 2736 3233 2744
rect 3747 2736 3833 2744
rect 3887 2735 3913 2743
rect 2107 2716 2133 2724
rect 2147 2716 2233 2724
rect 2536 2724 2544 2732
rect 2307 2716 2544 2724
rect 3836 2724 3844 2732
rect 4176 2727 4184 2756
rect 4356 2746 4364 2756
rect 4516 2756 4744 2764
rect 4516 2746 4524 2756
rect 4736 2746 4744 2756
rect 5176 2747 5184 2776
rect 5227 2776 5284 2784
rect 4527 2735 4553 2743
rect 4887 2736 4993 2744
rect 5067 2735 5093 2743
rect 5276 2746 5284 2776
rect 5307 2776 5333 2784
rect 5347 2776 5393 2784
rect 5473 2784 5487 2793
rect 5736 2796 5773 2804
rect 5473 2780 5553 2784
rect 5476 2776 5553 2780
rect 5607 2776 5693 2784
rect 5736 2764 5744 2796
rect 5716 2760 5744 2764
rect 5713 2756 5744 2760
rect 5713 2747 5727 2756
rect 5367 2735 5493 2743
rect 5547 2736 5613 2744
rect 5756 2744 5764 2773
rect 5756 2736 5773 2744
rect 3836 2716 4013 2724
rect 4467 2716 4593 2724
rect 4607 2716 4693 2724
rect 4996 2724 5004 2732
rect 4996 2716 5133 2724
rect 5147 2716 5233 2724
rect 5496 2724 5504 2732
rect 5796 2727 5804 2774
rect 5496 2716 5633 2724
rect 2847 2696 3273 2704
rect 3807 2696 3973 2704
rect 4147 2696 4213 2704
rect 5227 2676 5713 2684
rect 347 2656 553 2664
rect 1347 2656 1813 2664
rect 2587 2656 2953 2664
rect 2967 2656 2993 2664
rect 3467 2656 3593 2664
rect 4107 2656 5193 2664
rect 247 2636 993 2644
rect 3707 2636 4053 2644
rect 27 2616 2013 2624
rect 3167 2616 3593 2624
rect 3647 2616 4993 2624
rect 3267 2596 3493 2604
rect 4067 2596 4193 2604
rect 4627 2596 4953 2604
rect 5327 2596 5693 2604
rect 1047 2576 1173 2584
rect 1187 2576 1873 2584
rect 3367 2576 3393 2584
rect 3527 2576 3813 2584
rect 4216 2576 5213 2584
rect 1247 2556 1733 2564
rect 2247 2556 2553 2564
rect 4216 2564 4224 2576
rect 5487 2576 5553 2584
rect 3387 2556 4224 2564
rect 5127 2556 5333 2564
rect 807 2536 833 2544
rect 847 2536 933 2544
rect 3907 2536 4233 2544
rect 4547 2536 4753 2544
rect 207 2516 333 2524
rect 887 2516 1273 2524
rect 1287 2516 1573 2524
rect 1787 2516 2524 2524
rect 2516 2507 2524 2516
rect 2947 2516 3153 2524
rect 3727 2516 3853 2524
rect 4207 2516 4373 2524
rect 4587 2516 4793 2524
rect 5607 2516 5653 2524
rect 507 2496 633 2504
rect 2167 2496 2284 2504
rect 2276 2488 2284 2496
rect 2527 2496 2573 2504
rect 5076 2496 5253 2504
rect 5076 2488 5084 2496
rect 5267 2496 5533 2504
rect 5547 2496 5604 2504
rect 67 2484 80 2487
rect 67 2473 84 2484
rect 107 2476 224 2484
rect 76 2446 84 2473
rect 216 2446 224 2476
rect 287 2476 373 2484
rect 387 2476 453 2484
rect 567 2476 613 2484
rect 687 2476 733 2484
rect 947 2476 1113 2484
rect 1247 2484 1260 2487
rect 1247 2473 1264 2484
rect 1367 2476 1393 2484
rect 1407 2476 1513 2484
rect 1927 2477 1953 2485
rect 2087 2476 2113 2484
rect 2207 2477 2233 2485
rect 2287 2477 2353 2485
rect 2447 2477 2613 2485
rect 2787 2477 2833 2485
rect 3127 2477 3193 2485
rect 3207 2476 3313 2484
rect 3367 2476 3553 2484
rect 636 2456 824 2464
rect 636 2446 644 2456
rect 367 2435 413 2443
rect 527 2435 553 2443
rect 647 2436 693 2444
rect 767 2435 793 2443
rect 816 2444 824 2456
rect 1256 2446 1264 2473
rect 2356 2464 2364 2474
rect 2656 2464 2664 2474
rect 2356 2456 2664 2464
rect 816 2436 853 2444
rect 867 2435 933 2443
rect 2147 2436 2193 2444
rect 2307 2435 2453 2443
rect 2716 2427 2724 2474
rect 3036 2464 3044 2474
rect 2967 2456 3044 2464
rect 2907 2435 2933 2443
rect 2987 2435 3013 2443
rect 3076 2444 3084 2474
rect 3647 2476 3773 2484
rect 3787 2476 3833 2484
rect 3847 2476 3924 2484
rect 3076 2436 3173 2444
rect 3227 2436 3253 2444
rect 3267 2435 3293 2443
rect 3407 2436 3433 2444
rect 3627 2436 3713 2444
rect 3916 2446 3924 2476
rect 4027 2476 4053 2484
rect 3956 2464 3964 2474
rect 4367 2476 4413 2484
rect 4296 2464 4304 2474
rect 4687 2477 4713 2485
rect 4887 2476 4913 2484
rect 4927 2476 4953 2484
rect 4967 2476 5073 2484
rect 5176 2476 5213 2484
rect 5176 2464 5184 2476
rect 5387 2476 5413 2484
rect 5596 2484 5604 2496
rect 5596 2476 5613 2484
rect 5747 2477 5813 2485
rect 3956 2456 4304 2464
rect 5136 2456 5184 2464
rect 167 2416 273 2424
rect 287 2416 713 2424
rect 727 2416 993 2424
rect 1007 2416 1353 2424
rect 2067 2416 2373 2424
rect 2387 2416 2713 2424
rect 2727 2416 3493 2424
rect 3507 2416 3853 2424
rect 3956 2424 3964 2456
rect 4147 2436 4253 2444
rect 4507 2435 4533 2443
rect 4547 2435 4633 2443
rect 4747 2436 4793 2444
rect 4987 2436 5033 2444
rect 5136 2444 5144 2456
rect 5107 2436 5144 2444
rect 5167 2435 5193 2443
rect 5247 2435 5412 2443
rect 5447 2435 5493 2443
rect 5507 2436 5753 2444
rect 3867 2416 4693 2424
rect 1147 2396 1293 2404
rect 1607 2396 1833 2404
rect 1847 2396 2073 2404
rect 2847 2396 3053 2404
rect 3127 2396 3233 2404
rect 3887 2396 4053 2404
rect 4427 2396 4593 2404
rect 5587 2396 5633 2404
rect 5747 2396 5773 2404
rect 1447 2376 1784 2384
rect 827 2356 1293 2364
rect 1776 2364 1784 2376
rect 1927 2376 2053 2384
rect 2127 2376 2253 2384
rect 2467 2376 3093 2384
rect 4927 2376 5053 2384
rect 5447 2376 5533 2384
rect 1776 2356 1953 2364
rect 2687 2356 2984 2364
rect 2976 2347 2984 2356
rect 3567 2356 3693 2364
rect 4187 2356 4373 2364
rect 4487 2356 4673 2364
rect 4687 2356 5313 2364
rect 5707 2356 5753 2364
rect 27 2336 173 2344
rect 847 2336 893 2344
rect 1547 2336 1733 2344
rect 2607 2336 2633 2344
rect 2987 2336 3473 2344
rect 3647 2336 3673 2344
rect 3827 2336 3993 2344
rect 4267 2336 4413 2344
rect 4427 2336 4473 2344
rect 1247 2316 1873 2324
rect 5287 2316 5673 2324
rect 5687 2316 5813 2324
rect 47 2296 113 2304
rect 527 2296 593 2304
rect 707 2296 753 2304
rect 887 2296 953 2304
rect 1367 2296 1453 2304
rect 1627 2296 1813 2304
rect 2107 2296 2293 2304
rect 2767 2296 2813 2304
rect 4207 2296 4233 2304
rect 5107 2296 5253 2304
rect 5547 2296 5613 2304
rect 147 2276 173 2284
rect 647 2276 673 2284
rect 880 2284 893 2287
rect 876 2273 893 2284
rect 947 2284 960 2287
rect 947 2273 964 2284
rect 987 2276 1033 2284
rect 2567 2276 2744 2284
rect 56 2256 73 2264
rect 56 2227 64 2256
rect 140 2264 153 2267
rect 136 2253 153 2264
rect 247 2256 273 2264
rect 367 2257 553 2265
rect 576 2256 713 2264
rect 136 2226 144 2253
rect 227 2216 353 2224
rect 576 2226 584 2256
rect 836 2227 844 2253
rect 407 2215 513 2223
rect 876 2224 884 2273
rect 956 2264 964 2273
rect 956 2256 1053 2264
rect 916 2244 924 2254
rect 1320 2264 1333 2267
rect 1316 2253 1333 2264
rect 1707 2257 1733 2265
rect 916 2240 964 2244
rect 916 2236 967 2240
rect 953 2227 967 2236
rect 876 2216 893 2224
rect 1316 2226 1324 2253
rect 1416 2227 1424 2254
rect 1887 2257 2113 2265
rect 2187 2256 2224 2264
rect 2216 2244 2224 2256
rect 2247 2257 2333 2265
rect 2736 2267 2744 2276
rect 3047 2276 3073 2284
rect 3307 2276 3333 2284
rect 3767 2276 3793 2284
rect 3847 2276 3973 2284
rect 4167 2276 4493 2284
rect 4567 2276 4613 2284
rect 4627 2276 4653 2284
rect 4967 2276 5013 2284
rect 5727 2276 5773 2284
rect 2216 2236 2284 2244
rect 1067 2215 1093 2223
rect 1247 2215 1273 2223
rect 1407 2216 1424 2227
rect 1407 2213 1420 2216
rect 1487 2215 1613 2223
rect 1747 2216 1793 2224
rect 2007 2215 2092 2223
rect 2276 2226 2284 2236
rect 2127 2216 2153 2224
rect 2496 2224 2504 2254
rect 2607 2264 2620 2267
rect 2607 2253 2624 2264
rect 2747 2256 2793 2264
rect 3107 2257 3133 2265
rect 3156 2256 3173 2264
rect 2616 2226 2624 2253
rect 3156 2244 3164 2256
rect 3196 2256 3293 2264
rect 2916 2236 3164 2244
rect 2916 2226 2924 2236
rect 3196 2226 3204 2256
rect 3387 2256 3433 2264
rect 2427 2216 2504 2224
rect 2687 2215 2713 2223
rect 3476 2224 3484 2254
rect 3507 2264 3520 2267
rect 3507 2253 3524 2264
rect 3707 2256 3804 2264
rect 3516 2226 3524 2253
rect 3796 2226 3804 2256
rect 3867 2264 3880 2267
rect 3867 2253 3884 2264
rect 3876 2226 3884 2253
rect 4056 2244 4064 2254
rect 4127 2256 4193 2264
rect 4267 2256 4313 2264
rect 4456 2244 4464 2254
rect 4487 2256 4584 2264
rect 4056 2236 4464 2244
rect 3367 2216 3484 2224
rect 3947 2215 4113 2223
rect 4227 2215 4253 2223
rect 4456 2224 4464 2236
rect 4576 2226 4584 2256
rect 4707 2264 4720 2267
rect 4707 2253 4724 2264
rect 4907 2256 5153 2264
rect 5167 2257 5193 2265
rect 5327 2256 5373 2264
rect 5467 2257 5493 2265
rect 5556 2256 5593 2264
rect 4716 2226 4724 2253
rect 4307 2216 4533 2224
rect 4787 2216 4953 2224
rect 5556 2226 5564 2256
rect 5047 2216 5133 2224
rect 5287 2215 5313 2223
rect 5447 2215 5513 2223
rect 1527 2196 1633 2204
rect 2207 2196 2313 2204
rect 2327 2196 2393 2204
rect 2407 2196 2453 2204
rect 2716 2204 2724 2212
rect 2716 2196 2853 2204
rect 27 2176 93 2184
rect 507 2176 613 2184
rect 1367 2176 1593 2184
rect 1636 2184 1644 2193
rect 3207 2196 3233 2204
rect 3247 2196 3313 2204
rect 3767 2196 3833 2204
rect 4007 2196 4173 2204
rect 5207 2196 5233 2204
rect 5247 2196 5353 2204
rect 5467 2196 5493 2204
rect 1636 2176 2053 2184
rect 2067 2176 2093 2184
rect 2827 2176 2953 2184
rect 2967 2176 3153 2184
rect 3573 2184 3587 2193
rect 3387 2180 3587 2184
rect 3387 2176 3584 2180
rect 3987 2176 4993 2184
rect 627 2156 673 2164
rect 827 2156 933 2164
rect 3087 2156 3273 2164
rect 3407 2156 3733 2164
rect 967 2136 1393 2144
rect 1407 2136 1833 2144
rect 2747 2116 2893 2124
rect 2907 2116 3073 2124
rect 3747 2116 3793 2124
rect 3807 2116 4833 2124
rect 347 2096 573 2104
rect 587 2096 953 2104
rect 3147 2096 3353 2104
rect 867 2076 1033 2084
rect 1967 2076 2153 2084
rect 2247 2076 2733 2084
rect 2887 2076 2973 2084
rect 3347 2076 3453 2084
rect 4007 2076 4373 2084
rect 367 2036 413 2044
rect 2167 2036 3393 2044
rect 4347 2036 4413 2044
rect 4427 2036 4493 2044
rect 4507 2036 4873 2044
rect 5467 2036 5693 2044
rect 467 2016 593 2024
rect 607 2016 693 2024
rect 707 2016 1153 2024
rect 1167 2016 1253 2024
rect 1267 2016 1493 2024
rect 1507 2016 1593 2024
rect 1667 2016 1733 2024
rect 3167 2016 3333 2024
rect 3507 2016 3593 2024
rect 3607 2016 3753 2024
rect 4447 2016 4593 2024
rect 4607 2016 4713 2024
rect 387 1996 733 2004
rect 2467 1996 2813 2004
rect 3287 1996 3453 2004
rect 4627 1996 4653 2004
rect 5307 1996 5413 2004
rect 456 1976 713 1984
rect 456 1968 464 1976
rect 927 1976 953 1984
rect 1476 1976 1713 1984
rect 1476 1968 1484 1976
rect 1767 1976 1973 1984
rect 3687 1976 3784 1984
rect 3776 1968 3784 1976
rect 4107 1976 4133 1984
rect 4147 1976 4193 1984
rect 5147 1976 5733 1984
rect 5747 1976 5813 1984
rect 187 1957 213 1965
rect 987 1957 1013 1965
rect 256 1924 264 1954
rect 456 1927 464 1954
rect 1167 1956 1193 1964
rect 1367 1957 1473 1965
rect 1547 1956 1584 1964
rect 1576 1944 1584 1956
rect 1607 1957 1633 1965
rect 2016 1956 2033 1964
rect 1576 1936 1644 1944
rect 256 1916 353 1924
rect 447 1916 464 1927
rect 447 1913 460 1916
rect 807 1916 853 1924
rect 867 1916 893 1924
rect 947 1916 1033 1924
rect 1047 1916 1073 1924
rect 1636 1924 1644 1936
rect 1807 1936 1993 1944
rect 2016 1927 2024 1956
rect 2187 1956 2233 1964
rect 2247 1956 2313 1964
rect 2367 1957 2413 1965
rect 2967 1957 3013 1965
rect 3056 1956 3193 1964
rect 1636 1916 1733 1924
rect 2167 1915 2193 1923
rect 2447 1916 2513 1924
rect 2636 1924 2644 1954
rect 2696 1944 2704 1954
rect 2696 1936 2913 1944
rect 3056 1926 3064 1956
rect 3247 1956 3273 1964
rect 3387 1957 3413 1965
rect 3547 1957 3733 1965
rect 3787 1957 3913 1965
rect 4756 1956 4773 1964
rect 2636 1916 2793 1924
rect 2987 1916 3053 1924
rect 3367 1916 3533 1924
rect 3736 1916 3853 1924
rect 3107 1896 3173 1904
rect 3227 1896 3413 1904
rect 3736 1904 3744 1916
rect 4107 1916 4213 1924
rect 4227 1916 4393 1924
rect 4476 1924 4484 1954
rect 4407 1916 4484 1924
rect 4516 1927 4524 1954
rect 4516 1916 4533 1927
rect 4520 1913 4533 1916
rect 4756 1907 4764 1956
rect 4827 1956 4933 1964
rect 5027 1956 5053 1964
rect 5207 1956 5233 1964
rect 5347 1956 5373 1964
rect 5496 1944 5504 1954
rect 5627 1956 5673 1964
rect 5456 1936 5504 1944
rect 5107 1915 5253 1923
rect 5456 1924 5464 1936
rect 5416 1920 5464 1924
rect 5413 1916 5464 1920
rect 5413 1907 5427 1916
rect 5487 1915 5513 1923
rect 5527 1916 5553 1924
rect 3596 1896 3744 1904
rect 167 1876 333 1884
rect 487 1876 513 1884
rect 1607 1876 1693 1884
rect 1707 1876 1793 1884
rect 1987 1876 2333 1884
rect 2487 1876 2833 1884
rect 2947 1876 3073 1884
rect 3596 1884 3604 1896
rect 3287 1876 3604 1884
rect 2007 1856 2033 1864
rect 2047 1856 2173 1864
rect 2187 1856 2253 1864
rect 3367 1856 3613 1864
rect 4707 1856 4793 1864
rect 207 1836 393 1844
rect 407 1836 573 1844
rect 2807 1836 3093 1844
rect 4267 1836 4313 1844
rect 1307 1816 2313 1824
rect 2407 1816 2613 1824
rect 3167 1816 3233 1824
rect 3707 1816 3773 1824
rect 3867 1816 4093 1824
rect 4287 1816 4533 1824
rect 5467 1816 5693 1824
rect 1147 1796 1593 1804
rect 1727 1796 1773 1804
rect 1787 1796 1813 1804
rect 2007 1796 2153 1804
rect 2387 1796 2833 1804
rect 2847 1796 2953 1804
rect 3027 1796 3113 1804
rect 3467 1796 3573 1804
rect 4087 1796 4133 1804
rect 4407 1796 4473 1804
rect 4847 1796 5213 1804
rect 847 1776 953 1784
rect 1107 1776 1233 1784
rect 1667 1776 1833 1784
rect 2027 1776 2073 1784
rect 2707 1776 2733 1784
rect 2747 1776 2973 1784
rect 3276 1776 3313 1784
rect 427 1756 473 1764
rect 2467 1756 2653 1764
rect 2976 1764 2984 1773
rect 3276 1764 3284 1776
rect 3787 1776 3873 1784
rect 3887 1776 4273 1784
rect 5027 1776 5133 1784
rect 5147 1776 5393 1784
rect 5687 1776 5773 1784
rect 2976 1756 3284 1764
rect 3807 1756 3833 1764
rect 4307 1756 4413 1764
rect 4427 1756 4453 1764
rect 4527 1756 4873 1764
rect 96 1706 104 1753
rect 516 1736 593 1744
rect 216 1704 224 1734
rect 436 1707 444 1734
rect 216 1696 313 1704
rect 367 1695 392 1703
rect 427 1696 444 1707
rect 516 1706 524 1736
rect 707 1737 733 1745
rect 1047 1737 1093 1745
rect 1116 1736 1133 1744
rect 796 1707 804 1734
rect 1116 1707 1124 1736
rect 1507 1737 1553 1745
rect 1767 1737 1913 1745
rect 427 1693 440 1696
rect 787 1704 804 1707
rect 787 1696 933 1704
rect 787 1693 800 1696
rect 1073 1684 1087 1693
rect 1207 1695 1293 1703
rect 1367 1696 1493 1704
rect 1856 1706 1864 1737
rect 1927 1737 1933 1745
rect 2147 1736 2193 1744
rect 2473 1724 2487 1733
rect 2473 1720 2604 1724
rect 2476 1716 2604 1720
rect 1787 1695 1813 1703
rect 1967 1696 2053 1704
rect 2107 1695 2133 1703
rect 2467 1695 2493 1703
rect 2596 1704 2604 1716
rect 2596 1696 2633 1704
rect 2796 1704 2804 1734
rect 3307 1736 3393 1744
rect 3567 1737 3713 1745
rect 2727 1696 2873 1704
rect 2916 1704 2924 1733
rect 3473 1724 3487 1733
rect 3473 1720 3504 1724
rect 3476 1716 3504 1720
rect 2916 1696 3053 1704
rect 3067 1696 3113 1704
rect 3187 1696 3353 1704
rect 3496 1706 3504 1716
rect 3427 1695 3472 1703
rect 3516 1704 3524 1734
rect 3947 1736 3973 1744
rect 4027 1736 4064 1744
rect 4056 1707 4064 1736
rect 4173 1744 4187 1753
rect 4147 1740 4187 1744
rect 4147 1736 4184 1740
rect 4207 1737 4253 1745
rect 4607 1736 4653 1744
rect 4093 1724 4107 1733
rect 4093 1720 4244 1724
rect 4096 1716 4244 1720
rect 3516 1696 3653 1704
rect 3907 1695 3933 1703
rect 4236 1704 4244 1716
rect 4236 1696 4373 1704
rect 4427 1696 4493 1704
rect 4696 1704 4704 1734
rect 4787 1736 4973 1744
rect 5176 1736 5273 1744
rect 5176 1706 5184 1736
rect 5347 1736 5393 1744
rect 4587 1696 4704 1704
rect 4727 1695 4773 1703
rect 5007 1695 5033 1703
rect 5636 1706 5644 1753
rect 5767 1737 5793 1745
rect 5227 1696 5453 1704
rect 1007 1680 1087 1684
rect 1007 1676 1084 1680
rect 1496 1676 1573 1684
rect 1496 1664 1504 1676
rect 2567 1676 2573 1684
rect 3116 1684 3124 1692
rect 2587 1676 3593 1684
rect 3607 1676 3693 1684
rect 4007 1676 4073 1684
rect 4207 1676 4253 1684
rect 4567 1676 4913 1684
rect 1067 1656 1504 1664
rect 1547 1656 1633 1664
rect 1907 1656 2273 1664
rect 2687 1656 2813 1664
rect 2987 1656 3033 1664
rect 4627 1656 4673 1664
rect 4967 1656 5093 1664
rect 5107 1656 5153 1664
rect 5527 1656 5573 1664
rect 5587 1656 5813 1664
rect 267 1636 593 1644
rect 1247 1636 1313 1644
rect 2347 1636 2453 1644
rect 2907 1636 3353 1644
rect 3547 1636 3893 1644
rect 4047 1636 4433 1644
rect 1367 1616 1473 1624
rect 2667 1616 3013 1624
rect 227 1596 373 1604
rect 2747 1596 2993 1604
rect 3087 1596 3253 1604
rect 4167 1596 4453 1604
rect 4527 1596 5053 1604
rect 987 1576 1053 1584
rect 4487 1576 4813 1584
rect 267 1556 413 1564
rect 2007 1556 2173 1564
rect 4867 1556 5253 1564
rect 487 1536 773 1544
rect 2367 1536 2433 1544
rect 2607 1536 2933 1544
rect 2947 1536 4173 1544
rect 5307 1536 5433 1544
rect 507 1516 613 1524
rect 627 1516 813 1524
rect 947 1516 1193 1524
rect 1587 1516 2073 1524
rect 2807 1516 2953 1524
rect 3516 1516 3853 1524
rect 3516 1507 3524 1516
rect 4247 1516 4353 1524
rect 4367 1516 4413 1524
rect 4467 1516 4753 1524
rect 5707 1516 5753 1524
rect 467 1496 533 1504
rect 1127 1496 1253 1504
rect 3027 1496 3053 1504
rect 3067 1496 3513 1504
rect 4187 1496 4513 1504
rect 5267 1496 5393 1504
rect 327 1476 673 1484
rect 687 1476 773 1484
rect 1287 1476 1473 1484
rect 1747 1476 2013 1484
rect 2836 1476 2993 1484
rect 2836 1467 2844 1476
rect 3007 1476 3733 1484
rect 4827 1476 4893 1484
rect 5127 1476 5293 1484
rect 5567 1476 5693 1484
rect 187 1456 273 1464
rect 827 1456 873 1464
rect 2316 1456 2833 1464
rect 2316 1448 2324 1456
rect 3687 1456 3713 1464
rect 4016 1456 4053 1464
rect 4016 1448 4024 1456
rect 4347 1456 4393 1464
rect 4747 1456 5164 1464
rect 147 1436 293 1444
rect 307 1436 333 1444
rect 407 1436 573 1444
rect 600 1444 613 1447
rect 596 1433 613 1444
rect 676 1436 713 1444
rect 596 1406 604 1433
rect 676 1424 684 1436
rect 787 1444 800 1447
rect 787 1433 804 1444
rect 947 1436 984 1444
rect 647 1416 684 1424
rect 796 1406 804 1433
rect 976 1424 984 1436
rect 1007 1436 1053 1444
rect 1127 1437 1153 1445
rect 1407 1437 1433 1445
rect 1907 1436 1964 1444
rect 976 1416 1044 1424
rect 1036 1406 1044 1416
rect 107 1396 233 1404
rect 487 1395 533 1403
rect 1087 1396 1113 1404
rect 1236 1404 1244 1433
rect 1187 1396 1244 1404
rect 1316 1404 1324 1434
rect 1956 1424 1964 1436
rect 2247 1436 2293 1444
rect 1956 1416 2104 1424
rect 1287 1396 1324 1404
rect 1347 1396 1393 1404
rect 2096 1406 2104 1416
rect 1667 1395 1713 1403
rect 2116 1404 2124 1434
rect 2307 1436 2313 1444
rect 2980 1444 2993 1447
rect 2116 1396 2333 1404
rect 2516 1404 2524 1434
rect 2516 1396 2593 1404
rect 2687 1395 2753 1403
rect 2916 1404 2924 1434
rect 2976 1433 2993 1444
rect 3056 1436 3193 1444
rect 2976 1406 2984 1433
rect 2827 1396 2924 1404
rect 3056 1387 3064 1436
rect 3567 1436 3913 1444
rect 4287 1437 4313 1445
rect 4336 1436 4453 1444
rect 3436 1407 3444 1434
rect 4336 1424 4344 1436
rect 4527 1436 4573 1444
rect 4587 1436 4744 1444
rect 4136 1416 4344 1424
rect 4736 1424 4744 1436
rect 4787 1436 4873 1444
rect 4947 1436 4993 1444
rect 5007 1436 5073 1444
rect 5096 1436 5133 1444
rect 5096 1424 5104 1436
rect 5156 1444 5164 1456
rect 5207 1456 5233 1464
rect 5156 1436 5253 1444
rect 5267 1437 5333 1445
rect 5407 1444 5420 1447
rect 5407 1433 5424 1444
rect 5527 1437 5593 1445
rect 4736 1416 4764 1424
rect 3436 1396 3453 1407
rect 3440 1393 3453 1396
rect 3587 1396 3713 1404
rect 3807 1396 3893 1404
rect 4136 1404 4144 1416
rect 4127 1396 4144 1404
rect 4407 1395 4493 1403
rect 4507 1396 4653 1404
rect 4756 1406 4764 1416
rect 4996 1416 5104 1424
rect 4867 1395 4933 1403
rect 4996 1404 5004 1416
rect 5416 1406 5424 1433
rect 5476 1407 5484 1434
rect 4987 1396 5004 1404
rect 5476 1396 5493 1407
rect 5480 1393 5493 1396
rect 5627 1395 5653 1403
rect 2147 1376 2253 1384
rect 2407 1376 2453 1384
rect 3867 1376 3933 1384
rect 4567 1376 4593 1384
rect 5727 1376 5753 1384
rect 647 1356 833 1364
rect 927 1356 1273 1364
rect 1287 1356 1313 1364
rect 1567 1356 1773 1364
rect 2947 1356 3033 1364
rect 3327 1356 3413 1364
rect 3847 1356 4193 1364
rect 5227 1356 5253 1364
rect 5267 1356 5573 1364
rect 367 1336 473 1344
rect 987 1336 1293 1344
rect 1307 1336 1333 1344
rect 2767 1336 3093 1344
rect 3907 1336 4273 1344
rect 5387 1336 5513 1344
rect 847 1316 1493 1324
rect 1547 1316 2193 1324
rect 2547 1316 2613 1324
rect 2967 1316 3053 1324
rect 3247 1316 3533 1324
rect 4427 1316 4753 1324
rect 4907 1316 4973 1324
rect 4987 1316 5033 1324
rect 5127 1316 5313 1324
rect 5327 1316 5493 1324
rect 767 1296 813 1304
rect 2007 1296 2044 1304
rect 187 1276 253 1284
rect 407 1276 493 1284
rect 1487 1276 1553 1284
rect 2036 1284 2044 1296
rect 2067 1296 2133 1304
rect 2907 1296 3113 1304
rect 2036 1276 2113 1284
rect 2207 1276 2273 1284
rect 3007 1276 3313 1284
rect 3327 1276 3453 1284
rect 4487 1276 5073 1284
rect 5667 1276 5793 1284
rect 607 1256 913 1264
rect 1127 1256 1293 1264
rect 1407 1256 1453 1264
rect 1587 1256 1753 1264
rect 2007 1256 2173 1264
rect 4307 1256 4333 1264
rect 4467 1256 4693 1264
rect 4827 1256 4873 1264
rect 5247 1256 5513 1264
rect 176 1236 313 1244
rect 176 1228 184 1236
rect 1207 1236 1233 1244
rect 2227 1236 2353 1244
rect 2367 1236 2413 1244
rect 2427 1236 2633 1244
rect 2727 1236 2793 1244
rect 2807 1236 2873 1244
rect 2887 1236 2973 1244
rect 3027 1236 3053 1244
rect 3067 1236 3133 1244
rect 3607 1236 3633 1244
rect 4147 1236 4324 1244
rect 147 1217 173 1225
rect 227 1216 393 1224
rect 476 1216 553 1224
rect 56 1187 64 1213
rect 476 1204 484 1216
rect 927 1216 1013 1224
rect 1036 1216 1153 1224
rect 1036 1204 1044 1216
rect 1267 1224 1280 1227
rect 1267 1213 1284 1224
rect 436 1196 484 1204
rect 796 1196 1044 1204
rect 107 1176 133 1184
rect 247 1175 273 1183
rect 436 1184 444 1196
rect 796 1186 804 1196
rect 1276 1186 1284 1213
rect 1316 1186 1324 1233
rect 1553 1224 1567 1233
rect 4316 1228 4324 1236
rect 5027 1236 5093 1244
rect 1553 1220 1593 1224
rect 1556 1216 1593 1220
rect 1436 1204 1444 1214
rect 1787 1217 1833 1225
rect 2087 1216 2173 1224
rect 2247 1216 2313 1224
rect 2487 1216 2584 1224
rect 1436 1196 1484 1204
rect 347 1176 444 1184
rect 467 1176 573 1184
rect 987 1175 1133 1183
rect 1187 1176 1273 1184
rect 1407 1175 1453 1183
rect 1476 1184 1484 1196
rect 1636 1187 1644 1213
rect 1476 1176 1573 1184
rect 1727 1175 1753 1183
rect 1967 1175 1993 1183
rect 2207 1176 2333 1184
rect 2396 1184 2404 1213
rect 2576 1186 2584 1216
rect 2396 1176 2453 1184
rect 2687 1176 2773 1184
rect 2856 1184 2864 1214
rect 3367 1216 3413 1224
rect 3436 1216 3493 1224
rect 3036 1187 3044 1213
rect 3313 1204 3327 1213
rect 3436 1204 3444 1216
rect 3667 1217 3713 1225
rect 3736 1216 3753 1224
rect 3736 1204 3744 1216
rect 3987 1216 4093 1224
rect 4107 1216 4233 1224
rect 4327 1216 4373 1224
rect 4447 1216 4473 1224
rect 4667 1217 4793 1225
rect 4816 1216 4833 1224
rect 3313 1200 3344 1204
rect 3316 1196 3344 1200
rect 2787 1176 2864 1184
rect 2887 1176 2993 1184
rect 3336 1186 3344 1196
rect 3376 1196 3444 1204
rect 3616 1196 3744 1204
rect 3376 1186 3384 1196
rect 3616 1186 3624 1196
rect 4287 1204 4300 1207
rect 4816 1204 4824 1216
rect 4847 1216 4933 1224
rect 5207 1217 5233 1225
rect 5413 1224 5427 1233
rect 5327 1216 5404 1224
rect 5413 1220 5444 1224
rect 5416 1216 5444 1220
rect 4287 1193 4304 1204
rect 3127 1175 3173 1183
rect 4296 1184 4304 1193
rect 4716 1196 4824 1204
rect 4976 1204 4984 1214
rect 5276 1204 5284 1214
rect 4976 1196 5284 1204
rect 4716 1186 4724 1196
rect 4296 1176 4493 1184
rect 5027 1175 5053 1183
rect 5276 1184 5284 1196
rect 5396 1187 5404 1216
rect 5187 1176 5284 1184
rect 5436 1186 5444 1216
rect 5467 1217 5553 1225
rect 5567 1216 5653 1224
rect 5816 1187 5824 1213
rect 47 1156 733 1164
rect 2507 1156 2533 1164
rect 2547 1156 2613 1164
rect 3667 1156 3853 1164
rect 4647 1156 4673 1164
rect 4927 1156 5133 1164
rect 1047 1136 1233 1144
rect 1367 1136 1653 1144
rect 3147 1136 3573 1144
rect 3767 1136 3793 1144
rect 4387 1136 4433 1144
rect 4487 1136 4553 1144
rect 4967 1136 5244 1144
rect 1236 1124 1244 1133
rect 1236 1116 2133 1124
rect 3287 1116 3393 1124
rect 4227 1116 4273 1124
rect 5236 1124 5244 1136
rect 5236 1116 5293 1124
rect 5307 1116 5673 1124
rect 747 1096 1353 1104
rect 1627 1096 1773 1104
rect 1907 1096 2113 1104
rect 2127 1096 2393 1104
rect 2547 1096 2733 1104
rect 2747 1096 2993 1104
rect 3247 1096 3753 1104
rect 4447 1096 4593 1104
rect 4767 1096 5224 1104
rect 1776 1084 1784 1093
rect 1776 1076 3013 1084
rect 3187 1076 3533 1084
rect 3747 1076 4213 1084
rect 5216 1084 5224 1096
rect 5216 1076 5333 1084
rect 5347 1076 5713 1084
rect 2107 1056 2253 1064
rect 2267 1056 3153 1064
rect 3167 1056 4433 1064
rect 4527 1056 4833 1064
rect 4467 1036 4713 1044
rect 1887 1016 2404 1024
rect 407 996 473 1004
rect 1487 996 1633 1004
rect 1987 996 2013 1004
rect 2396 1004 2404 1016
rect 3127 1016 3233 1024
rect 4067 1016 4413 1024
rect 4807 1016 4873 1024
rect 2396 996 4613 1004
rect 4667 996 5093 1004
rect 5107 996 5213 1004
rect 427 976 633 984
rect 727 976 793 984
rect 807 976 2013 984
rect 2373 984 2387 993
rect 2373 980 2933 984
rect 2376 976 2933 980
rect 2947 976 3213 984
rect 3327 976 3413 984
rect 3647 976 3833 984
rect 3847 976 4113 984
rect 4307 976 4513 984
rect 547 956 593 964
rect 1687 956 1813 964
rect 2336 960 2453 964
rect 2333 956 2453 960
rect 2333 947 2347 956
rect 2467 956 2493 964
rect 2627 956 2873 964
rect 3287 956 4184 964
rect 4176 947 4184 956
rect 4547 956 4653 964
rect 4707 956 4813 964
rect 5407 956 5453 964
rect 5687 956 5773 964
rect 367 936 393 944
rect 467 936 493 944
rect 707 936 753 944
rect 1067 936 1333 944
rect 1347 936 1413 944
rect 1547 944 1560 947
rect 1547 933 1564 944
rect 3307 936 3513 944
rect 3576 936 3793 944
rect 107 916 213 924
rect 687 916 824 924
rect 56 887 64 913
rect 376 896 433 904
rect 376 886 384 896
rect 147 875 193 883
rect 467 875 513 883
rect 536 867 544 914
rect 816 887 824 916
rect 847 917 873 925
rect 887 917 913 925
rect 967 917 993 925
rect 1187 916 1204 924
rect 1196 904 1204 916
rect 1227 916 1273 924
rect 1196 896 1224 904
rect 567 876 653 884
rect 816 876 833 887
rect 820 873 833 876
rect 1007 876 1073 884
rect 1216 884 1224 896
rect 1376 887 1384 914
rect 1216 876 1253 884
rect 1367 876 1384 887
rect 1556 886 1564 933
rect 1827 916 1933 924
rect 2067 916 2173 924
rect 2187 917 2293 925
rect 2407 916 2613 924
rect 1776 904 1784 914
rect 1607 896 1784 904
rect 2416 887 2424 916
rect 3067 916 3264 924
rect 2656 887 2664 914
rect 1367 873 1380 876
rect 1447 875 1473 883
rect 1707 876 1833 884
rect 1887 875 1913 883
rect 2567 876 2593 884
rect 2656 876 2673 887
rect 2660 873 2673 876
rect 2816 884 2824 914
rect 3256 904 3264 916
rect 3367 916 3453 924
rect 3576 924 3584 936
rect 4187 936 4353 944
rect 3467 916 3584 924
rect 3607 916 3693 924
rect 3907 916 4073 924
rect 4147 916 4213 924
rect 4527 917 4573 925
rect 4627 917 4653 925
rect 4680 924 4693 927
rect 4676 913 4693 924
rect 4767 916 4864 924
rect 3256 896 3344 904
rect 2816 876 2913 884
rect 3336 884 3344 896
rect 4076 896 4273 904
rect 3336 876 3373 884
rect 3647 875 3673 883
rect 3727 876 3853 884
rect 3867 875 3893 883
rect 4076 884 4084 896
rect 4676 904 4684 913
rect 4636 896 4684 904
rect 4856 904 4864 916
rect 4887 917 4933 925
rect 5007 916 5133 924
rect 5207 917 5413 925
rect 5787 916 5894 924
rect 5556 904 5564 914
rect 4856 896 4904 904
rect 4067 876 4084 884
rect 4107 875 4133 883
rect 4207 876 4533 884
rect 4636 886 4644 896
rect 4896 886 4904 896
rect 5456 896 5564 904
rect 4687 876 4733 884
rect 4947 876 5013 884
rect 5167 876 5373 884
rect 5456 884 5464 896
rect 5387 876 5464 884
rect 5487 875 5533 883
rect 887 856 1033 864
rect 1876 864 1884 872
rect 1647 856 1884 864
rect 2527 856 2633 864
rect 327 836 413 844
rect 947 836 1013 844
rect 1067 836 1153 844
rect 1167 836 1353 844
rect 1507 836 1593 844
rect 2227 836 2272 844
rect 2516 844 2524 853
rect 2307 836 2524 844
rect 3587 836 3673 844
rect 3727 836 3833 844
rect 3887 836 4013 844
rect 4027 836 4113 844
rect 1547 816 1573 824
rect 2167 816 2764 824
rect 1927 796 2013 804
rect 2447 796 2613 804
rect 2756 804 2764 816
rect 3207 816 3233 824
rect 3387 816 3653 824
rect 5127 816 5293 824
rect 5307 816 5353 824
rect 2756 796 2793 804
rect 3087 796 3173 804
rect 3767 796 3893 804
rect 4867 796 5213 804
rect 87 776 113 784
rect 127 776 593 784
rect 607 776 653 784
rect 847 776 873 784
rect 1287 776 1393 784
rect 1627 776 1693 784
rect 2707 776 2873 784
rect 3007 776 3053 784
rect 3247 776 3413 784
rect 3527 776 3673 784
rect 3967 776 4213 784
rect 4447 776 4713 784
rect 5027 776 5413 784
rect 787 756 853 764
rect 1227 756 1313 764
rect 1767 756 1913 764
rect 2987 756 3013 764
rect 5287 756 5733 764
rect 167 736 233 744
rect 547 736 693 744
rect 707 736 1533 744
rect 1587 736 1673 744
rect 1947 736 2093 744
rect 2307 736 2393 744
rect 2447 736 2833 744
rect 3347 744 3360 747
rect 3347 733 3364 744
rect 3407 736 3513 744
rect 3667 736 3913 744
rect 4087 736 4273 744
rect 4467 736 4593 744
rect 4747 736 4793 744
rect 307 716 393 724
rect 727 716 753 724
rect 767 716 853 724
rect 2467 716 2553 724
rect 247 696 364 704
rect 196 684 204 694
rect 136 676 204 684
rect 136 664 144 676
rect 356 666 364 696
rect 107 656 144 664
rect 167 655 213 663
rect 476 664 484 694
rect 527 696 593 704
rect 1007 704 1020 707
rect 1007 693 1024 704
rect 1227 697 1373 705
rect 1396 696 1413 704
rect 1016 667 1024 693
rect 1396 684 1404 696
rect 1476 696 1633 704
rect 1267 676 1404 684
rect 476 656 573 664
rect 887 655 913 663
rect 1287 636 1433 644
rect 267 616 513 624
rect 1456 624 1464 694
rect 1476 666 1484 696
rect 1907 696 1973 704
rect 2147 696 2313 704
rect 1667 655 1693 663
rect 1856 664 1864 693
rect 2096 667 2104 694
rect 1856 656 1873 664
rect 1967 656 2052 664
rect 2087 656 2104 667
rect 2087 653 2100 656
rect 2167 655 2293 663
rect 2376 664 2384 694
rect 2407 696 2493 704
rect 2887 696 2913 704
rect 2927 696 3013 704
rect 2376 656 2513 664
rect 3007 656 3033 664
rect 3107 656 3213 664
rect 3336 664 3344 694
rect 3356 666 3364 733
rect 3387 716 3533 724
rect 4427 716 4473 724
rect 4676 716 4973 724
rect 3400 704 3413 707
rect 3396 693 3413 704
rect 3567 697 3613 705
rect 3627 696 3733 704
rect 3787 696 3833 704
rect 3847 697 4053 705
rect 4147 696 4193 704
rect 4327 697 4353 705
rect 4507 696 4593 704
rect 3396 666 3404 693
rect 3516 667 3524 693
rect 3227 656 3344 664
rect 4067 656 4113 664
rect 4207 655 4253 663
rect 4367 656 4393 664
rect 1907 636 2433 644
rect 2687 636 2913 644
rect 3507 636 3533 644
rect 3687 636 3793 644
rect 3967 636 4073 644
rect 4356 644 4364 653
rect 4407 656 4513 664
rect 4527 656 4573 664
rect 4676 666 4684 716
rect 4707 697 4773 705
rect 5047 696 5153 704
rect 5167 696 5253 704
rect 5387 697 5473 705
rect 5487 696 5513 704
rect 4747 655 4813 663
rect 4987 655 5133 663
rect 5227 656 5633 664
rect 4167 636 4364 644
rect 4607 636 4853 644
rect 4900 644 4913 647
rect 4896 633 4913 644
rect 5487 636 5693 644
rect 5707 636 5813 644
rect 1456 616 1593 624
rect 2287 616 2313 624
rect 3067 616 3433 624
rect 4896 624 4904 633
rect 4767 616 4904 624
rect 1127 596 1352 604
rect 1387 596 1573 604
rect 1807 596 1893 604
rect 2027 596 2193 604
rect 2207 596 2413 604
rect 2427 596 2553 604
rect 2567 596 2733 604
rect 3827 596 3893 604
rect 3907 596 4013 604
rect 4027 596 4593 604
rect 587 576 1553 584
rect 2087 576 2253 584
rect 2267 576 2473 584
rect 2487 576 2713 584
rect 2727 576 3093 584
rect 3267 576 3553 584
rect 3807 576 4233 584
rect 47 556 293 564
rect 307 556 973 564
rect 987 556 1033 564
rect 1347 556 1673 564
rect 1687 556 1813 564
rect 2747 556 3084 564
rect 1567 536 1793 544
rect 2647 536 2913 544
rect 3076 544 3084 556
rect 3207 556 3353 564
rect 3687 556 3753 564
rect 3076 536 3373 544
rect 3427 536 3813 544
rect 3927 536 3953 544
rect 3967 536 4153 544
rect 4247 536 4493 544
rect 4507 536 4773 544
rect 4867 536 4993 544
rect 1267 516 1813 524
rect 1827 516 1933 524
rect 2087 516 2413 524
rect 2487 516 2844 524
rect 1256 504 1264 513
rect 727 496 1264 504
rect 1727 496 1913 504
rect 2067 496 2433 504
rect 2627 496 2653 504
rect 2836 504 2844 516
rect 2867 516 3193 524
rect 3527 516 3753 524
rect 4467 516 4913 524
rect 2836 496 3133 504
rect 3227 496 3713 504
rect 3927 496 4192 504
rect 4227 496 4333 504
rect 4567 496 4653 504
rect 1587 476 2473 484
rect 2527 476 3013 484
rect 4147 476 4733 484
rect 227 456 413 464
rect 427 456 933 464
rect 2447 456 2973 464
rect 3047 456 3213 464
rect 3267 456 3873 464
rect 4127 456 5213 464
rect 367 436 413 444
rect 427 436 553 444
rect 1027 436 1093 444
rect 1927 436 1972 444
rect 2007 436 2032 444
rect 2067 436 2273 444
rect 2547 436 2733 444
rect 3067 436 3173 444
rect 4167 436 4513 444
rect 4727 436 5073 444
rect 607 416 733 424
rect 747 416 893 424
rect 907 416 953 424
rect 1127 416 1413 424
rect 1527 416 1733 424
rect 1747 416 1773 424
rect 1907 416 2073 424
rect 2276 416 2393 424
rect 267 397 393 405
rect 487 396 633 404
rect 116 364 124 394
rect 767 397 793 405
rect 1087 396 1173 404
rect 1267 404 1280 407
rect 1267 393 1284 404
rect 1467 397 1493 405
rect 1516 396 1533 404
rect 1276 366 1284 393
rect 1516 384 1524 396
rect 1547 396 1653 404
rect 1833 404 1847 413
rect 1833 400 2093 404
rect 1836 396 2093 400
rect 2147 397 2173 405
rect 2196 396 2213 404
rect 1416 376 1524 384
rect 116 356 193 364
rect 427 355 453 363
rect 587 356 693 364
rect 1207 355 1233 363
rect 1416 364 1424 376
rect 2196 367 2204 396
rect 2276 367 2284 416
rect 2687 416 2753 424
rect 2767 416 2873 424
rect 2947 416 3253 424
rect 3487 416 3513 424
rect 4107 416 4533 424
rect 5147 416 5253 424
rect 5267 416 5353 424
rect 2307 397 2353 405
rect 1407 356 1424 364
rect 1507 356 1553 364
rect 1847 356 1973 364
rect 2047 355 2073 363
rect 2496 364 2504 394
rect 2807 397 2833 405
rect 2900 404 2913 407
rect 2896 393 2913 404
rect 3227 396 3273 404
rect 3367 396 3424 404
rect 2896 366 2904 393
rect 3416 384 3424 396
rect 3447 396 3544 404
rect 3416 380 3504 384
rect 3416 376 3507 380
rect 3493 367 3507 376
rect 2387 356 2504 364
rect 2627 355 2673 363
rect 2947 356 2993 364
rect 3267 356 3373 364
rect 3536 366 3544 396
rect 3587 397 3633 405
rect 3827 397 4013 405
rect 4287 397 4373 405
rect 4527 397 4693 405
rect 5227 396 5304 404
rect 4127 355 4213 363
rect 4327 355 4632 363
rect 4667 355 4753 363
rect 4767 356 4813 364
rect 5296 366 5304 396
rect 5387 397 5573 405
rect 5776 367 5784 394
rect 5187 356 5233 364
rect 5367 355 5633 363
rect 5687 356 5753 364
rect 5776 356 5793 367
rect 5780 353 5793 356
rect 647 336 833 344
rect 967 336 1253 344
rect 2896 344 2904 352
rect 2896 336 3033 344
rect 3047 336 3113 344
rect 3256 344 3264 352
rect 3127 336 3264 344
rect 407 316 873 324
rect 1027 316 1113 324
rect 1367 316 1433 324
rect 1927 316 2293 324
rect 2727 316 2793 324
rect 3307 316 3473 324
rect 3487 316 3853 324
rect 3867 316 3993 324
rect 4287 316 4373 324
rect 4727 316 5093 324
rect 5647 316 5713 324
rect 5767 316 5793 324
rect 667 296 733 304
rect 876 304 884 313
rect 876 296 1153 304
rect 1267 296 1313 304
rect 1327 296 1833 304
rect 3087 296 3233 304
rect 3407 296 3472 304
rect 3507 296 3613 304
rect 3907 296 4113 304
rect 907 276 1024 284
rect 207 256 433 264
rect 1016 264 1024 276
rect 1867 276 2053 284
rect 2307 276 2533 284
rect 2867 276 3813 284
rect 4547 276 5453 284
rect 1016 256 1453 264
rect 1887 256 2013 264
rect 2287 256 2733 264
rect 3167 256 3393 264
rect 5567 256 5593 264
rect 1007 236 1553 244
rect 1627 236 2793 244
rect 3427 236 3573 244
rect 3667 236 3873 244
rect 4107 236 4353 244
rect 4627 236 4853 244
rect 5107 236 5693 244
rect 367 216 573 224
rect 587 216 613 224
rect 2207 216 2273 224
rect 2427 216 2613 224
rect 3487 216 3553 224
rect 3767 216 3804 224
rect 1467 196 1733 204
rect 2307 196 2653 204
rect 2667 196 2753 204
rect 2767 196 3164 204
rect 47 177 93 185
rect 107 176 313 184
rect 336 146 344 193
rect 3156 188 3164 196
rect 3247 196 3433 204
rect 3760 204 3773 207
rect 3756 193 3773 204
rect 3796 204 3804 216
rect 4047 216 4233 224
rect 4487 216 4593 224
rect 3796 196 3993 204
rect 4687 196 4733 204
rect 4867 196 4913 204
rect 5467 196 5513 204
rect 487 176 513 184
rect 707 177 933 185
rect 1047 176 1093 184
rect 1367 177 1413 185
rect 1507 176 1673 184
rect 2167 177 2192 185
rect 2227 176 2253 184
rect 2267 176 2333 184
rect 2807 176 2833 184
rect 2927 176 3113 184
rect 3167 177 3213 185
rect 3467 176 3493 184
rect 3647 176 3664 184
rect 2516 156 2553 164
rect 167 135 253 143
rect 407 136 453 144
rect 527 135 553 143
rect 707 136 733 144
rect 967 135 993 143
rect 1227 136 1353 144
rect 2516 146 2524 156
rect 2567 156 2984 164
rect 1596 136 1653 144
rect 1067 116 1204 124
rect 567 96 913 104
rect 1196 104 1204 116
rect 1596 124 1604 136
rect 1667 135 1733 143
rect 1887 135 1973 143
rect 2047 135 2093 143
rect 2427 135 2453 143
rect 2927 135 2953 143
rect 2976 144 2984 156
rect 3656 147 3664 176
rect 2976 136 3013 144
rect 3187 135 3233 143
rect 3347 135 3393 143
rect 3447 136 3613 144
rect 1547 116 1604 124
rect 3016 124 3024 132
rect 3756 127 3764 193
rect 4187 176 4413 184
rect 4508 176 4613 184
rect 4696 176 4793 184
rect 4416 144 4424 173
rect 4696 146 4704 176
rect 4876 176 5333 184
rect 4876 164 4884 176
rect 5567 184 5580 187
rect 5567 173 5584 184
rect 5727 176 5784 184
rect 4816 156 4884 164
rect 4816 146 4824 156
rect 5576 146 5584 173
rect 4407 136 4424 144
rect 4847 135 4973 143
rect 5347 135 5413 143
rect 5776 146 5784 176
rect 5707 136 5733 144
rect 3016 116 3273 124
rect 4327 116 4353 124
rect 4496 116 4553 124
rect 1196 96 1433 104
rect 1707 96 2213 104
rect 2287 96 2633 104
rect 2787 96 3133 104
rect 3307 96 3513 104
rect 4496 104 4504 116
rect 4607 116 4653 124
rect 5227 116 5673 124
rect 3967 96 4504 104
rect 4787 96 4913 104
rect 5387 96 5513 104
rect 1407 76 1493 84
rect 3567 76 3733 84
rect 3787 76 4513 84
rect 4807 76 4833 84
rect 5647 76 5813 84
rect 2687 56 2713 64
rect 2727 56 3293 64
rect 227 36 273 44
rect 287 36 793 44
rect 807 36 1273 44
rect 1287 36 1793 44
rect 1807 36 1893 44
rect 5047 36 5273 44
rect 5287 36 5633 44
rect 1927 16 3333 24
use NOR2X1  _723_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform -1 0 2890 0 -1 790
box -12 -8 74 272
use INVX2  _724_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform -1 0 2670 0 1 790
box -12 -8 52 272
use NOR2X1  _725_
timestamp 1701862152
transform -1 0 2770 0 -1 1310
box -12 -8 74 272
use OAI21X1  _726_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform 1 0 3370 0 1 270
box -12 -8 92 272
use INVX2  _727_
timestamp 1701862152
transform 1 0 2950 0 1 1830
box -12 -8 52 272
use NOR2X1  _728_
timestamp 1701862152
transform -1 0 3110 0 1 1830
box -12 -8 74 272
use AOI22X1  _729_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform 1 0 3710 0 -1 790
box -14 -8 114 272
use OAI21X1  _730_
timestamp 1702508443
transform 1 0 3610 0 1 270
box -12 -8 92 272
use INVX1  _731_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform -1 0 3550 0 1 270
box -12 -8 52 272
use INVX1  _732_
timestamp 1701862152
transform -1 0 830 0 1 790
box -12 -8 52 272
use NAND2X1  _733_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform -1 0 2070 0 1 790
box -12 -8 72 272
use OAI21X1  _734_
timestamp 1702508443
transform -1 0 3050 0 1 270
box -12 -8 92 272
use AOI22X1  _735_
timestamp 1701862152
transform 1 0 4150 0 1 270
box -14 -8 114 272
use OAI21X1  _736_
timestamp 1702508443
transform 1 0 3850 0 1 270
box -12 -8 92 272
use INVX1  _737_
timestamp 1701862152
transform 1 0 1010 0 -1 1310
box -12 -8 52 272
use NAND2X1  _738_
timestamp 1702508443
transform -1 0 2190 0 1 790
box -12 -8 72 272
use OAI21X1  _739_
timestamp 1702508443
transform -1 0 2910 0 1 270
box -12 -8 92 272
use AOI22X1  _740_
timestamp 1701862152
transform 1 0 4690 0 1 270
box -14 -8 114 272
use OAI21X1  _741_
timestamp 1702508443
transform 1 0 3990 0 1 270
box -12 -8 92 272
use NOR2X1  _742_
timestamp 1701862152
transform -1 0 3030 0 -1 790
box -12 -8 74 272
use OAI21X1  _743_
timestamp 1702508443
transform 1 0 3110 0 1 270
box -12 -8 92 272
use AOI22X1  _744_
timestamp 1701862152
transform -1 0 4570 0 -1 270
box -14 -8 114 272
use OAI21X1  _745_
timestamp 1702508443
transform 1 0 3710 0 -1 270
box -12 -8 92 272
use INVX2  _746_
timestamp 1701862152
transform 1 0 2310 0 1 3910
box -12 -8 52 272
use NAND2X1  _747_
timestamp 1702508443
transform 1 0 3310 0 1 2870
box -12 -8 72 272
use OAI21X1  _748_
timestamp 1702508443
transform 1 0 3170 0 1 2870
box -12 -8 92 272
use INVX1  _749_
timestamp 1701862152
transform 1 0 2210 0 1 3910
box -12 -8 52 272
use NAND2X1  _750_
timestamp 1702508443
transform -1 0 3350 0 -1 3390
box -12 -8 72 272
use OAI21X1  _751_
timestamp 1702508443
transform 1 0 3410 0 -1 3390
box -12 -8 92 272
use INVX2  _752_
timestamp 1701862152
transform 1 0 1690 0 1 2870
box -12 -8 52 272
use NAND2X1  _753_
timestamp 1702508443
transform 1 0 3570 0 1 2870
box -12 -8 72 272
use OAI21X1  _754_
timestamp 1702508443
transform 1 0 3430 0 1 2870
box -12 -8 92 272
use INVX2  _755_
timestamp 1701862152
transform -1 0 1490 0 1 2870
box -12 -8 52 272
use NAND2X1  _756_
timestamp 1702508443
transform 1 0 2690 0 -1 3910
box -12 -8 72 272
use OAI21X1  _757_
timestamp 1702508443
transform 1 0 2550 0 -1 3910
box -12 -8 92 272
use NAND2X1  _758_
timestamp 1702508443
transform -1 0 2430 0 1 3390
box -12 -8 72 272
use OAI21X1  _759_
timestamp 1702508443
transform 1 0 2230 0 1 3390
box -12 -8 92 272
use NAND2X1  _760_
timestamp 1702508443
transform -1 0 2230 0 -1 3390
box -12 -8 72 272
use OAI21X1  _761_
timestamp 1702508443
transform 1 0 2090 0 1 3390
box -12 -8 92 272
use NAND2X1  _762_
timestamp 1702508443
transform -1 0 2230 0 1 2870
box -12 -8 72 272
use OAI21X1  _763_
timestamp 1702508443
transform -1 0 2370 0 1 2870
box -12 -8 92 272
use NAND2X1  _764_
timestamp 1702508443
transform 1 0 2050 0 -1 2870
box -12 -8 72 272
use OAI21X1  _765_
timestamp 1702508443
transform -1 0 2270 0 -1 2870
box -12 -8 92 272
use INVX1  _766_
timestamp 1701862152
transform 1 0 3410 0 1 1310
box -12 -8 52 272
use NAND2X1  _767_
timestamp 1702508443
transform 1 0 2790 0 1 1310
box -12 -8 72 272
use OAI21X1  _768_
timestamp 1702508443
transform -1 0 2990 0 1 1310
box -12 -8 92 272
use INVX1  _769_
timestamp 1701862152
transform -1 0 4250 0 -1 1310
box -12 -8 52 272
use NAND2X1  _770_
timestamp 1702508443
transform -1 0 3630 0 -1 1310
box -12 -8 72 272
use OAI21X1  _771_
timestamp 1702508443
transform -1 0 3770 0 -1 1310
box -12 -8 92 272
use INVX1  _772_
timestamp 1701862152
transform -1 0 5490 0 -1 790
box -12 -8 52 272
use NAND2X1  _773_
timestamp 1702508443
transform -1 0 4370 0 1 1310
box -12 -8 72 272
use OAI21X1  _774_
timestamp 1702508443
transform -1 0 4910 0 1 790
box -12 -8 92 272
use INVX1  _775_
timestamp 1701862152
transform -1 0 5810 0 -1 2870
box -12 -8 52 272
use NAND2X1  _776_
timestamp 1702508443
transform 1 0 4950 0 1 2350
box -12 -8 72 272
use OAI21X1  _777_
timestamp 1702508443
transform 1 0 5730 0 1 4430
box -12 -8 92 272
use INVX1  _778_
timestamp 1701862152
transform 1 0 5410 0 -1 1310
box -12 -8 52 272
use NAND2X1  _779_
timestamp 1702508443
transform -1 0 4430 0 -1 1830
box -12 -8 72 272
use OAI21X1  _780_
timestamp 1702508443
transform -1 0 4890 0 -1 1830
box -12 -8 92 272
use INVX1  _781_
timestamp 1701862152
transform -1 0 5170 0 -1 2350
box -12 -8 52 272
use NAND2X1  _782_
timestamp 1702508443
transform -1 0 3850 0 -1 2350
box -12 -8 72 272
use OAI21X1  _783_
timestamp 1702508443
transform -1 0 5070 0 -1 2350
box -12 -8 92 272
use INVX1  _784_
timestamp 1701862152
transform 1 0 3870 0 -1 1830
box -12 -8 52 272
use NAND2X1  _785_
timestamp 1702508443
transform -1 0 3510 0 1 1830
box -12 -8 72 272
use OAI21X1  _786_
timestamp 1702508443
transform -1 0 3570 0 -1 1830
box -12 -8 92 272
use INVX1  _787_
timestamp 1701862152
transform -1 0 4270 0 1 2350
box -12 -8 52 272
use NAND2X1  _788_
timestamp 1702508443
transform -1 0 3650 0 1 2350
box -12 -8 72 272
use OAI21X1  _789_
timestamp 1702508443
transform -1 0 3930 0 1 2350
box -12 -8 92 272
use INVX1  _790_
timestamp 1701862152
transform 1 0 1930 0 -1 1830
box -12 -8 52 272
use NAND2X1  _791_
timestamp 1702508443
transform -1 0 2230 0 -1 1830
box -12 -8 72 272
use OAI21X1  _792_
timestamp 1702508443
transform 1 0 2030 0 -1 1830
box -12 -8 92 272
use INVX1  _793_
timestamp 1701862152
transform 1 0 1030 0 -1 270
box -12 -8 52 272
use NAND2X1  _794_
timestamp 1702508443
transform 1 0 1650 0 -1 270
box -12 -8 72 272
use OAI21X1  _795_
timestamp 1702508443
transform -1 0 1470 0 -1 270
box -12 -8 92 272
use INVX1  _796_
timestamp 1701862152
transform -1 0 590 0 -1 270
box -12 -8 52 272
use NAND2X1  _797_
timestamp 1702508443
transform 1 0 1530 0 -1 270
box -12 -8 72 272
use OAI21X1  _798_
timestamp 1702508443
transform 1 0 890 0 -1 270
box -12 -8 92 272
use INVX1  _799_
timestamp 1701862152
transform 1 0 1550 0 1 1310
box -12 -8 52 272
use NAND2X1  _800_
timestamp 1702508443
transform 1 0 2310 0 1 1310
box -12 -8 72 272
use OAI21X1  _801_
timestamp 1702508443
transform 1 0 2050 0 1 1310
box -12 -8 92 272
use INVX1  _802_
timestamp 1701862152
transform -1 0 490 0 1 1830
box -12 -8 52 272
use NAND2X1  _803_
timestamp 1702508443
transform -1 0 1330 0 -1 2350
box -12 -8 72 272
use OAI21X1  _804_
timestamp 1702508443
transform 1 0 710 0 -1 2350
box -12 -8 92 272
use INVX1  _805_
timestamp 1701862152
transform -1 0 1050 0 1 1830
box -12 -8 52 272
use NAND2X1  _806_
timestamp 1702508443
transform 1 0 2290 0 -1 1830
box -12 -8 72 272
use OAI21X1  _807_
timestamp 1702508443
transform 1 0 1130 0 -1 1830
box -12 -8 92 272
use INVX1  _808_
timestamp 1701862152
transform 1 0 1030 0 -1 1830
box -12 -8 52 272
use NAND2X1  _809_
timestamp 1702508443
transform 1 0 1510 0 1 2350
box -12 -8 72 272
use OAI21X1  _810_
timestamp 1702508443
transform -1 0 1610 0 -1 1830
box -12 -8 92 272
use INVX1  _811_
timestamp 1701862152
transform -1 0 1390 0 1 1830
box -12 -8 52 272
use NAND2X1  _812_
timestamp 1702508443
transform 1 0 2310 0 1 1830
box -12 -8 72 272
use OAI21X1  _813_
timestamp 1702508443
transform 1 0 1690 0 1 1830
box -12 -8 92 272
use INVX1  _814_
timestamp 1701862152
transform 1 0 3390 0 -1 1830
box -12 -8 52 272
use NAND3X1  _815_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform 1 0 3690 0 -1 2870
box -12 -8 92 272
use OAI21X1  _816_
timestamp 1702508443
transform 1 0 3570 0 1 1830
box -12 -8 92 272
use INVX8  _817_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform 1 0 4490 0 -1 1830
box -12 -8 114 272
use NAND2X1  _818_
timestamp 1702508443
transform -1 0 4190 0 -1 2870
box -12 -8 72 272
use NAND2X1  _819_
timestamp 1702508443
transform 1 0 3690 0 1 2870
box -12 -8 72 272
use XNOR2X1  _820_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform -1 0 4370 0 -1 2870
box -12 -8 132 272
use NAND2X1  _821_
timestamp 1702508443
transform 1 0 4110 0 -1 1830
box -12 -8 72 272
use OAI21X1  _822_
timestamp 1702508443
transform -1 0 4310 0 -1 1830
box -12 -8 92 272
use NOR2X1  _823_
timestamp 1701862152
transform 1 0 4430 0 -1 2870
box -12 -8 74 272
use NAND2X1  _824_
timestamp 1702508443
transform 1 0 4010 0 1 3390
box -12 -8 72 272
use NAND2X1  _825_
timestamp 1702508443
transform -1 0 4210 0 1 3390
box -12 -8 72 272
use NOR2X1  _826_
timestamp 1701862152
transform -1 0 4290 0 -1 3390
box -12 -8 74 272
use AOI22X1  _827_
timestamp 1701862152
transform -1 0 4030 0 -1 3390
box -14 -8 114 272
use OAI21X1  _828_
timestamp 1702508443
transform 1 0 4190 0 1 2870
box -12 -8 92 272
use INVX1  _829_
timestamp 1701862152
transform 1 0 3810 0 1 2870
box -12 -8 52 272
use AND2X2  _830_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform -1 0 4310 0 -1 3910
box -12 -8 94 272
use AND2X2  _831_
timestamp 1701862152
transform 1 0 4110 0 -1 4430
box -12 -8 94 272
use NAND2X1  _832_
timestamp 1702508443
transform -1 0 4170 0 -1 3910
box -12 -8 72 272
use INVX1  _833_
timestamp 1701862152
transform -1 0 3210 0 -1 3390
box -12 -8 52 272
use INVX1  _834_
timestamp 1701862152
transform 1 0 3410 0 1 4430
box -12 -8 52 272
use NAND2X1  _835_
timestamp 1702508443
transform 1 0 3690 0 -1 3390
box -12 -8 72 272
use OAI21X1  _836_
timestamp 1702508443
transform 1 0 3550 0 -1 3390
box -12 -8 92 272
use NAND3X1  _837_
timestamp 1702508443
transform 1 0 3910 0 1 2870
box -12 -8 92 272
use NAND3X1  _838_
timestamp 1702508443
transform 1 0 4690 0 -1 2870
box -12 -8 92 272
use INVX1  _839_
timestamp 1701862152
transform -1 0 5030 0 -1 2870
box -12 -8 52 272
use AOI21X1  _840_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform 1 0 4550 0 -1 2870
box -12 -8 92 272
use OAI21X1  _841_
timestamp 1702508443
transform 1 0 4850 0 -1 2870
box -12 -8 92 272
use INVX1  _842_
timestamp 1701862152
transform -1 0 5170 0 -1 790
box -12 -8 52 272
use NAND2X1  _843_
timestamp 1702508443
transform -1 0 4690 0 -1 790
box -12 -8 72 272
use AND2X2  _844_
timestamp 1701862152
transform -1 0 4830 0 -1 790
box -12 -8 94 272
use INVX1  _845_
timestamp 1701862152
transform -1 0 5770 0 1 2350
box -12 -8 52 272
use NAND2X1  _846_
timestamp 1702508443
transform -1 0 3470 0 1 3390
box -12 -8 72 272
use AOI21X1  _847_
timestamp 1702508443
transform 1 0 4050 0 1 2870
box -12 -8 92 272
use NAND2X1  _848_
timestamp 1702508443
transform 1 0 4390 0 -1 3910
box -12 -8 72 272
use NAND2X1  _849_
timestamp 1702508443
transform 1 0 4550 0 1 4430
box -12 -8 72 272
use NOR2X1  _850_
timestamp 1701862152
transform -1 0 4330 0 1 3390
box -12 -8 74 272
use AOI22X1  _851_
timestamp 1701862152
transform 1 0 4510 0 -1 3910
box -14 -8 114 272
use OAI21X1  _852_
timestamp 1702508443
transform 1 0 4610 0 1 3390
box -12 -8 92 272
use INVX1  _853_
timestamp 1701862152
transform 1 0 4390 0 1 3390
box -12 -8 52 272
use AND2X2  _854_
timestamp 1701862152
transform 1 0 4310 0 1 3910
box -12 -8 94 272
use NAND2X1  _855_
timestamp 1702508443
transform 1 0 4190 0 1 3910
box -12 -8 72 272
use INVX1  _856_
timestamp 1701862152
transform 1 0 4510 0 1 3390
box -12 -8 52 272
use NAND3X1  _857_
timestamp 1702508443
transform 1 0 4630 0 -1 3390
box -12 -8 92 272
use NAND3X1  _858_
timestamp 1702508443
transform -1 0 4710 0 1 2870
box -12 -8 92 272
use OAI21X1  _859_
timestamp 1702508443
transform -1 0 4170 0 -1 3390
box -12 -8 92 272
use AOI21X1  _860_
timestamp 1702508443
transform -1 0 4570 0 -1 3390
box -12 -8 92 272
use INVX2  _861_
timestamp 1701862152
transform 1 0 3410 0 1 3910
box -12 -8 52 272
use OAI21X1  _862_
timestamp 1702508443
transform 1 0 3650 0 1 3910
box -12 -8 92 272
use INVX2  _863_
timestamp 1701862152
transform -1 0 2470 0 1 3910
box -12 -8 52 272
use INVX1  _864_
timestamp 1701862152
transform -1 0 4710 0 1 4430
box -12 -8 52 272
use OAI21X1  _865_
timestamp 1702508443
transform 1 0 3910 0 1 3910
box -12 -8 92 272
use AOI21X1  _866_
timestamp 1702508443
transform 1 0 4050 0 1 3910
box -12 -8 92 272
use OAI21X1  _867_
timestamp 1702508443
transform 1 0 4350 0 -1 3390
box -12 -8 92 272
use NAND3X1  _868_
timestamp 1702508443
transform 1 0 4490 0 1 2870
box -12 -8 92 272
use INVX1  _869_
timestamp 1701862152
transform 1 0 4890 0 1 3390
box -12 -8 52 272
use NAND3X1  _870_
timestamp 1702508443
transform 1 0 4770 0 -1 3390
box -12 -8 92 272
use OAI21X1  _871_
timestamp 1702508443
transform 1 0 4350 0 1 2870
box -12 -8 92 272
use NAND3X1  _872_
timestamp 1702508443
transform 1 0 4770 0 1 2870
box -12 -8 92 272
use AOI21X1  _873_
timestamp 1702508443
transform 1 0 5090 0 -1 2870
box -12 -8 92 272
use NAND3X1  _874_
timestamp 1702508443
transform 1 0 5230 0 -1 2870
box -12 -8 92 272
use NAND2X1  _875_
timestamp 1702508443
transform 1 0 5070 0 1 2350
box -12 -8 72 272
use OAI22X1  _876_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform -1 0 5290 0 1 2350
box -12 -8 112 272
use INVX1  _877_
timestamp 1701862152
transform -1 0 5530 0 1 1830
box -12 -8 52 272
use INVX1  _878_
timestamp 1701862152
transform 1 0 5390 0 -1 2870
box -12 -8 52 272
use AOI21X1  _879_
timestamp 1702508443
transform 1 0 4910 0 -1 3390
box -12 -8 92 272
use OAI21X1  _880_
timestamp 1702508443
transform 1 0 5050 0 -1 3390
box -12 -8 92 272
use OAI21X1  _881_
timestamp 1702508443
transform 1 0 4670 0 -1 3910
box -12 -8 92 272
use AND2X2  _882_
timestamp 1701862152
transform -1 0 4850 0 1 4950
box -12 -8 94 272
use NAND2X1  _883_
timestamp 1702508443
transform 1 0 4450 0 1 3910
box -12 -8 72 272
use AOI22X1  _884_
timestamp 1701862152
transform -1 0 4490 0 -1 4430
box -14 -8 114 272
use INVX1  _885_
timestamp 1701862152
transform -1 0 4610 0 1 3910
box -12 -8 52 272
use NAND2X1  _886_
timestamp 1702508443
transform 1 0 4270 0 -1 4430
box -12 -8 72 272
use INVX1  _887_
timestamp 1701862152
transform -1 0 5130 0 -1 4430
box -12 -8 52 272
use NAND3X1  _888_
timestamp 1702508443
transform -1 0 5030 0 1 3910
box -12 -8 92 272
use NAND2X1  _889_
timestamp 1702508443
transform 1 0 4750 0 -1 4950
box -12 -8 72 272
use NOR2X1  _890_
timestamp 1701862152
transform 1 0 4810 0 -1 4430
box -12 -8 74 272
use OAI21X1  _891_
timestamp 1702508443
transform -1 0 4750 0 1 3910
box -12 -8 92 272
use AOI21X1  _892_
timestamp 1702508443
transform 1 0 4930 0 -1 3910
box -12 -8 92 272
use AOI21X1  _893_
timestamp 1702508443
transform 1 0 4750 0 1 3390
box -12 -8 92 272
use NAND3X1  _894_
timestamp 1702508443
transform 1 0 5110 0 1 3910
box -12 -8 92 272
use OAI21X1  _895_
timestamp 1702508443
transform 1 0 4810 0 1 3910
box -12 -8 92 272
use AOI21X1  _896_
timestamp 1702508443
transform 1 0 5130 0 1 3390
box -12 -8 92 272
use NAND2X1  _897_
timestamp 1702508443
transform 1 0 3370 0 -1 3910
box -12 -8 72 272
use INVX1  _898_
timestamp 1701862152
transform 1 0 2790 0 -1 3390
box -12 -8 52 272
use INVX2  _899_
timestamp 1701862152
transform 1 0 1810 0 -1 3910
box -12 -8 52 272
use NAND2X1  _900_
timestamp 1702508443
transform -1 0 3370 0 -1 4430
box -12 -8 72 272
use OAI21X1  _901_
timestamp 1702508443
transform 1 0 3270 0 1 3390
box -12 -8 92 272
use OAI21X1  _902_
timestamp 1702508443
transform -1 0 3570 0 -1 3910
box -12 -8 92 272
use OAI21X1  _903_
timestamp 1702508443
transform -1 0 5290 0 -1 3910
box -12 -8 92 272
use NAND3X1  _904_
timestamp 1702508443
transform 1 0 4990 0 1 3390
box -12 -8 92 272
use NAND3X1  _905_
timestamp 1702508443
transform 1 0 5070 0 -1 3910
box -12 -8 92 272
use INVX1  _906_
timestamp 1701862152
transform 1 0 5490 0 -1 3910
box -12 -8 52 272
use NAND3X1  _907_
timestamp 1702508443
transform -1 0 5350 0 1 3390
box -12 -8 92 272
use NAND3X1  _908_
timestamp 1702508443
transform 1 0 5190 0 -1 3390
box -12 -8 92 272
use INVX1  _909_
timestamp 1701862152
transform -1 0 5110 0 1 2870
box -12 -8 52 272
use AOI21X1  _910_
timestamp 1702508443
transform 1 0 4910 0 1 2870
box -12 -8 92 272
use AOI21X1  _911_
timestamp 1702508443
transform -1 0 5490 0 1 3390
box -12 -8 92 272
use INVX1  _912_
timestamp 1701862152
transform 1 0 5330 0 -1 3390
box -12 -8 52 272
use OAI21X1  _913_
timestamp 1702508443
transform -1 0 5370 0 1 2870
box -12 -8 92 272
use AOI21X1  _914_
timestamp 1702508443
transform 1 0 5490 0 -1 2870
box -12 -8 92 272
use NAND3X1  _915_
timestamp 1702508443
transform 1 0 5630 0 -1 2870
box -12 -8 92 272
use NAND2X1  _916_
timestamp 1702508443
transform 1 0 5610 0 1 2350
box -12 -8 72 272
use OAI22X1  _917_
timestamp 1701862152
transform 1 0 5490 0 -1 2350
box -12 -8 112 272
use AND2X2  _918_
timestamp 1701862152
transform -1 0 3710 0 -1 3910
box -12 -8 94 272
use NAND2X1  _919_
timestamp 1702508443
transform 1 0 4810 0 -1 3910
box -12 -8 72 272
use INVX1  _920_
timestamp 1701862152
transform 1 0 5730 0 -1 3390
box -12 -8 52 272
use AOI21X1  _921_
timestamp 1702508443
transform 1 0 5550 0 1 3390
box -12 -8 92 272
use NAND2X1  _922_
timestamp 1702508443
transform 1 0 2630 0 1 3910
box -12 -8 72 272
use AND2X2  _923_
timestamp 1701862152
transform -1 0 3170 0 -1 3910
box -12 -8 94 272
use OAI21X1  _924_
timestamp 1702508443
transform -1 0 3030 0 -1 3910
box -12 -8 92 272
use INVX2  _925_
timestamp 1701862152
transform -1 0 2570 0 1 3910
box -12 -8 52 272
use OAI21X1  _926_
timestamp 1702508443
transform 1 0 2990 0 1 3910
box -12 -8 92 272
use NAND3X1  _927_
timestamp 1702508443
transform 1 0 2850 0 1 3910
box -12 -8 92 272
use INVX1  _928_
timestamp 1701862152
transform 1 0 2750 0 1 3910
box -12 -8 52 272
use NAND2X1  _929_
timestamp 1702508443
transform -1 0 3190 0 1 3910
box -12 -8 72 272
use OAI21X1  _930_
timestamp 1702508443
transform 1 0 3230 0 -1 3910
box -12 -8 92 272
use NAND3X1  _931_
timestamp 1702508443
transform 1 0 3270 0 1 3910
box -12 -8 92 272
use NAND2X1  _932_
timestamp 1702508443
transform -1 0 4610 0 -1 4430
box -12 -8 72 272
use OAI22X1  _933_
timestamp 1701862152
transform 1 0 4930 0 -1 4430
box -12 -8 112 272
use INVX1  _934_
timestamp 1701862152
transform 1 0 5250 0 -1 4950
box -12 -8 52 272
use NAND2X1  _935_
timestamp 1702508443
transform -1 0 4550 0 -1 4950
box -12 -8 72 272
use NAND3X1  _936_
timestamp 1702508443
transform 1 0 5330 0 1 4950
box -12 -8 92 272
use NAND2X1  _937_
timestamp 1702508443
transform 1 0 5090 0 -1 5470
box -12 -8 72 272
use NAND3X1  _938_
timestamp 1702508443
transform 1 0 5070 0 1 4950
box -12 -8 92 272
use NAND3X1  _939_
timestamp 1702508443
transform -1 0 5570 0 1 4950
box -12 -8 92 272
use INVX1  _940_
timestamp 1701862152
transform 1 0 5770 0 -1 5470
box -12 -8 52 272
use AND2X2  _941_
timestamp 1701862152
transform -1 0 4610 0 -1 5470
box -12 -8 94 272
use NAND2X1  _942_
timestamp 1702508443
transform -1 0 4730 0 -1 5470
box -12 -8 72 272
use OAI21X1  _943_
timestamp 1702508443
transform 1 0 5030 0 1 4430
box -12 -8 92 272
use NAND3X1  _944_
timestamp 1702508443
transform -1 0 5430 0 -1 5470
box -12 -8 92 272
use NAND3X1  _945_
timestamp 1702508443
transform 1 0 5350 0 -1 4950
box -12 -8 92 272
use AOI21X1  _946_
timestamp 1702508443
transform 1 0 5490 0 -1 5470
box -12 -8 92 272
use AOI21X1  _947_
timestamp 1702508443
transform 1 0 5650 0 1 4950
box -12 -8 92 272
use OAI21X1  _948_
timestamp 1702508443
transform -1 0 5710 0 -1 4950
box -12 -8 92 272
use NAND3X1  _949_
timestamp 1702508443
transform -1 0 5530 0 1 4430
box -12 -8 92 272
use AND2X2  _950_
timestamp 1701862152
transform 1 0 4670 0 -1 4430
box -12 -8 94 272
use NAND3X1  _951_
timestamp 1702508443
transform -1 0 5190 0 -1 4950
box -12 -8 92 272
use OAI21X1  _952_
timestamp 1702508443
transform -1 0 5570 0 -1 4950
box -12 -8 92 272
use NAND3X1  _953_
timestamp 1702508443
transform 1 0 5170 0 1 4430
box -12 -8 92 272
use NAND3X1  _954_
timestamp 1702508443
transform 1 0 5490 0 -1 4430
box -12 -8 92 272
use OAI21X1  _955_
timestamp 1702508443
transform 1 0 5350 0 -1 3910
box -12 -8 92 272
use AOI21X1  _956_
timestamp 1702508443
transform 1 0 5310 0 1 4430
box -12 -8 92 272
use AOI21X1  _957_
timestamp 1702508443
transform 1 0 5590 0 1 4430
box -12 -8 92 272
use OAI21X1  _958_
timestamp 1702508443
transform -1 0 5710 0 -1 4430
box -12 -8 92 272
use NAND3X1  _959_
timestamp 1702508443
transform 1 0 5630 0 -1 5470
box -12 -8 92 272
use NAND3X1  _960_
timestamp 1702508443
transform 1 0 5330 0 -1 4430
box -12 -8 92 272
use OAI21X1  _961_
timestamp 1702508443
transform -1 0 5730 0 1 3910
box -12 -8 92 272
use NAND3X1  _962_
timestamp 1702508443
transform 1 0 5610 0 -1 3910
box -12 -8 92 272
use NAND2X1  _963_
timestamp 1702508443
transform -1 0 5750 0 1 3390
box -12 -8 72 272
use NAND2X1  _964_
timestamp 1702508443
transform 1 0 5430 0 1 2870
box -12 -8 72 272
use XNOR2X1  _965_
timestamp 1702508443
transform 1 0 5550 0 1 2870
box -12 -8 132 272
use NAND2X1  _966_
timestamp 1702508443
transform 1 0 4710 0 1 2350
box -12 -8 72 272
use OAI21X1  _967_
timestamp 1702508443
transform -1 0 4650 0 1 2350
box -12 -8 92 272
use INVX1  _968_
timestamp 1701862152
transform -1 0 4230 0 1 1830
box -12 -8 52 272
use AOI22X1  _969_
timestamp 1701862152
transform -1 0 5670 0 -1 3390
box -14 -8 114 272
use AOI21X1  _970_
timestamp 1702508443
transform 1 0 5190 0 -1 4430
box -12 -8 92 272
use OAI21X1  _971_
timestamp 1702508443
transform 1 0 5250 0 1 3910
box -12 -8 92 272
use NAND2X1  _972_
timestamp 1702508443
transform -1 0 3250 0 -1 4430
box -12 -8 72 272
use OAI21X1  _973_
timestamp 1702508443
transform 1 0 3430 0 -1 4430
box -12 -8 92 272
use INVX1  _974_
timestamp 1701862152
transform 1 0 3870 0 1 4430
box -12 -8 52 272
use INVX1  _975_
timestamp 1701862152
transform 1 0 4870 0 -1 4950
box -12 -8 52 272
use AOI21X1  _976_
timestamp 1702508443
transform -1 0 4970 0 1 4430
box -12 -8 92 272
use NAND2X1  _977_
timestamp 1702508443
transform -1 0 2990 0 -1 4430
box -12 -8 72 272
use AND2X2  _978_
timestamp 1701862152
transform -1 0 2690 0 1 4430
box -12 -8 94 272
use OAI21X1  _979_
timestamp 1702508443
transform -1 0 2850 0 -1 4430
box -12 -8 92 272
use AND2X2  _980_
timestamp 1701862152
transform 1 0 2350 0 -1 4430
box -12 -8 94 272
use OAI21X1  _981_
timestamp 1702508443
transform 1 0 2490 0 -1 4430
box -12 -8 92 272
use NAND3X1  _982_
timestamp 1702508443
transform -1 0 2710 0 -1 4430
box -12 -8 92 272
use INVX1  _983_
timestamp 1701862152
transform 1 0 3050 0 1 4430
box -12 -8 52 272
use NAND2X1  _984_
timestamp 1702508443
transform 1 0 2770 0 1 4430
box -12 -8 72 272
use OAI21X1  _985_
timestamp 1702508443
transform 1 0 3050 0 -1 4430
box -12 -8 92 272
use NAND3X1  _986_
timestamp 1702508443
transform 1 0 3150 0 1 4430
box -12 -8 92 272
use NAND2X1  _987_
timestamp 1702508443
transform 1 0 3290 0 -1 4950
box -12 -8 72 272
use NOR2X1  _988_
timestamp 1701862152
transform 1 0 5210 0 1 4950
box -12 -8 74 272
use AOI21X1  _989_
timestamp 1702508443
transform -1 0 5290 0 -1 5470
box -12 -8 92 272
use NAND2X1  _990_
timestamp 1702508443
transform -1 0 2570 0 -1 5470
box -12 -8 72 272
use NAND2X1  _991_
timestamp 1702508443
transform -1 0 3710 0 1 4950
box -12 -8 72 272
use NAND3X1  _992_
timestamp 1702508443
transform 1 0 3370 0 1 4950
box -12 -8 92 272
use NAND2X1  _993_
timestamp 1702508443
transform 1 0 1710 0 1 4950
box -12 -8 72 272
use NAND3X1  _994_
timestamp 1702508443
transform -1 0 3590 0 1 4950
box -12 -8 92 272
use NAND3X1  _995_
timestamp 1702508443
transform 1 0 3290 0 -1 5470
box -12 -8 92 272
use INVX1  _996_
timestamp 1701862152
transform -1 0 3090 0 -1 5470
box -12 -8 52 272
use AND2X2  _997_
timestamp 1701862152
transform -1 0 2410 0 1 4430
box -12 -8 94 272
use NAND2X1  _998_
timestamp 1702508443
transform -1 0 2830 0 -1 5470
box -12 -8 72 272
use OAI21X1  _999_
timestamp 1702508443
transform 1 0 3150 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1000_
timestamp 1702508443
transform 1 0 3150 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1001_
timestamp 1702508443
transform 1 0 4110 0 -1 5470
box -12 -8 92 272
use AOI22X1  _1002_
timestamp 1701862152
transform 1 0 4910 0 1 4950
box -14 -8 114 272
use OAI21X1  _1003_
timestamp 1702508443
transform 1 0 4810 0 -1 5470
box -12 -8 92 272
use AOI22X1  _1004_
timestamp 1701862152
transform -1 0 3670 0 -1 5470
box -14 -8 114 272
use AOI21X1  _1005_
timestamp 1702508443
transform 1 0 3430 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1006_
timestamp 1702508443
transform 1 0 4390 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1007_
timestamp 1702508443
transform -1 0 4590 0 1 4950
box -12 -8 92 272
use AND2X2  _1008_
timestamp 1701862152
transform 1 0 3410 0 -1 4950
box -12 -8 94 272
use NAND3X1  _1009_
timestamp 1702508443
transform -1 0 4050 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1010_
timestamp 1702508443
transform -1 0 4330 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1011_
timestamp 1702508443
transform -1 0 4170 0 1 4950
box -12 -8 92 272
use NAND3X1  _1012_
timestamp 1702508443
transform 1 0 4090 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1013_
timestamp 1702508443
transform -1 0 5050 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1014_
timestamp 1702508443
transform 1 0 4610 0 -1 4950
box -12 -8 92 272
use AOI21X1  _1015_
timestamp 1702508443
transform 1 0 4230 0 1 4950
box -12 -8 92 272
use AOI21X1  _1016_
timestamp 1702508443
transform -1 0 4450 0 1 4950
box -12 -8 92 272
use OAI21X1  _1017_
timestamp 1702508443
transform -1 0 4310 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1018_
timestamp 1702508443
transform -1 0 4210 0 1 4430
box -12 -8 92 272
use NAND3X1  _1019_
timestamp 1702508443
transform -1 0 3890 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1020_
timestamp 1702508443
transform -1 0 4350 0 1 4430
box -12 -8 92 272
use NAND3X1  _1021_
timestamp 1702508443
transform -1 0 3650 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1022_
timestamp 1702508443
transform -1 0 3850 0 1 3910
box -12 -8 72 272
use XNOR2X1  _1023_
timestamp 1702508443
transform 1 0 3930 0 -1 3910
box -12 -8 132 272
use NOR2X1  _1024_
timestamp 1701862152
transform 1 0 3810 0 -1 3390
box -12 -8 74 272
use NAND3X1  _1025_
timestamp 1702508443
transform -1 0 3590 0 1 3910
box -12 -8 92 272
use INVX1  _1026_
timestamp 1701862152
transform 1 0 5410 0 1 3910
box -12 -8 52 272
use AOI21X1  _1027_
timestamp 1702508443
transform -1 0 5590 0 1 3910
box -12 -8 92 272
use AOI21X1  _1028_
timestamp 1702508443
transform 1 0 3710 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1029_
timestamp 1702508443
transform -1 0 4050 0 1 4430
box -12 -8 92 272
use OAI21X1  _1030_
timestamp 1702508443
transform 1 0 3850 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1031_
timestamp 1702508443
transform 1 0 3670 0 1 3390
box -12 -8 92 272
use NAND2X1  _1032_
timestamp 1702508443
transform 1 0 3830 0 -1 2870
box -12 -8 72 272
use OAI22X1  _1033_
timestamp 1701862152
transform -1 0 4050 0 -1 2870
box -12 -8 112 272
use OAI21X1  _1034_
timestamp 1702508443
transform -1 0 3870 0 -1 3910
box -12 -8 92 272
use INVX1  _1035_
timestamp 1701862152
transform -1 0 3810 0 1 4430
box -12 -8 52 272
use AOI21X1  _1036_
timestamp 1702508443
transform -1 0 3710 0 1 4430
box -12 -8 92 272
use NAND2X1  _1037_
timestamp 1702508443
transform 1 0 3290 0 1 4430
box -12 -8 72 272
use INVX1  _1038_
timestamp 1701862152
transform -1 0 2650 0 -1 4950
box -12 -8 52 272
use INVX1  _1039_
timestamp 1701862152
transform 1 0 3870 0 -1 5470
box -12 -8 52 272
use AOI21X1  _1040_
timestamp 1702508443
transform -1 0 4010 0 1 4950
box -12 -8 92 272
use NAND2X1  _1041_
timestamp 1702508443
transform -1 0 2290 0 -1 4430
box -12 -8 72 272
use AND2X2  _1042_
timestamp 1701862152
transform -1 0 1770 0 1 4430
box -12 -8 94 272
use OAI21X1  _1043_
timestamp 1702508443
transform -1 0 1650 0 -1 4430
box -12 -8 92 272
use AND2X2  _1044_
timestamp 1701862152
transform -1 0 2150 0 1 3910
box -12 -8 94 272
use OAI21X1  _1045_
timestamp 1702508443
transform -1 0 2010 0 1 3910
box -12 -8 92 272
use NAND3X1  _1046_
timestamp 1702508443
transform 1 0 1830 0 -1 4430
box -12 -8 92 272
use INVX1  _1047_
timestamp 1701862152
transform -1 0 2130 0 1 4430
box -12 -8 52 272
use NAND2X1  _1048_
timestamp 1702508443
transform -1 0 1770 0 -1 4430
box -12 -8 72 272
use NAND2X1  _1049_
timestamp 1702508443
transform -1 0 2270 0 1 4430
box -12 -8 72 272
use OAI21X1  _1050_
timestamp 1702508443
transform 1 0 2070 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1051_
timestamp 1702508443
transform -1 0 2030 0 1 4430
box -12 -8 92 272
use NAND2X1  _1052_
timestamp 1702508443
transform 1 0 1910 0 -1 4950
box -12 -8 72 272
use AOI22X1  _1053_
timestamp 1701862152
transform 1 0 2890 0 -1 5470
box -14 -8 114 272
use NAND2X1  _1054_
timestamp 1702508443
transform -1 0 1510 0 1 4950
box -12 -8 72 272
use NAND2X1  _1055_
timestamp 1702508443
transform 1 0 1350 0 -1 4950
box -12 -8 72 272
use NOR2X1  _1056_
timestamp 1701862152
transform 1 0 1330 0 1 4950
box -12 -8 74 272
use AOI22X1  _1057_
timestamp 1701862152
transform 1 0 1470 0 -1 4950
box -14 -8 114 272
use OAI21X1  _1058_
timestamp 1702508443
transform 1 0 1350 0 -1 5470
box -12 -8 92 272
use INVX1  _1059_
timestamp 1701862152
transform 1 0 1250 0 -1 5470
box -12 -8 52 272
use AND2X2  _1060_
timestamp 1701862152
transform 1 0 1630 0 -1 4950
box -12 -8 94 272
use NAND2X1  _1061_
timestamp 1702508443
transform 1 0 1230 0 -1 4950
box -12 -8 72 272
use INVX1  _1062_
timestamp 1701862152
transform -1 0 910 0 -1 5470
box -12 -8 52 272
use NAND3X1  _1063_
timestamp 1702508443
transform 1 0 970 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1064_
timestamp 1702508443
transform 1 0 1790 0 -1 5470
box -12 -8 92 272
use AOI22X1  _1065_
timestamp 1701862152
transform -1 0 3290 0 1 4950
box -14 -8 114 272
use OAI21X1  _1066_
timestamp 1702508443
transform 1 0 2630 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1067_
timestamp 1702508443
transform 1 0 1110 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1068_
timestamp 1702508443
transform -1 0 1850 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1069_
timestamp 1702508443
transform -1 0 2550 0 1 4430
box -12 -8 92 272
use AOI21X1  _1070_
timestamp 1702508443
transform 1 0 1830 0 1 4950
box -12 -8 92 272
use OAI21X1  _1071_
timestamp 1702508443
transform 1 0 2090 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1072_
timestamp 1702508443
transform 1 0 2230 0 -1 5470
box -12 -8 92 272
use AND2X2  _1073_
timestamp 1701862152
transform 1 0 2030 0 -1 4950
box -12 -8 94 272
use NAND3X1  _1074_
timestamp 1702508443
transform 1 0 1630 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1075_
timestamp 1702508443
transform 1 0 1930 0 -1 5470
box -12 -8 92 272
use NAND3X1  _1076_
timestamp 1702508443
transform 1 0 2350 0 1 4950
box -12 -8 92 272
use NAND3X1  _1077_
timestamp 1702508443
transform 1 0 2770 0 1 4950
box -12 -8 92 272
use AOI21X1  _1078_
timestamp 1702508443
transform 1 0 3730 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1079_
timestamp 1702508443
transform 1 0 3790 0 1 4950
box -12 -8 92 272
use AOI21X1  _1080_
timestamp 1702508443
transform 1 0 2210 0 1 4950
box -12 -8 92 272
use AOI21X1  _1081_
timestamp 1702508443
transform 1 0 2370 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1082_
timestamp 1702508443
transform -1 0 2990 0 1 4950
box -12 -8 92 272
use AOI21X1  _1083_
timestamp 1702508443
transform 1 0 2470 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1084_
timestamp 1702508443
transform 1 0 2630 0 1 4950
box -12 -8 92 272
use OAI21X1  _1085_
timestamp 1702508443
transform 1 0 3050 0 1 4950
box -12 -8 92 272
use AOI21X1  _1086_
timestamp 1702508443
transform 1 0 2850 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1087_
timestamp 1702508443
transform 1 0 2910 0 1 4430
box -12 -8 92 272
use AOI21X1  _1088_
timestamp 1702508443
transform -1 0 4030 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1089_
timestamp 1702508443
transform 1 0 3670 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1090_
timestamp 1702508443
transform 1 0 2710 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1091_
timestamp 1702508443
transform 1 0 2330 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1092_
timestamp 1702508443
transform -1 0 3070 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1093_
timestamp 1702508443
transform -1 0 2930 0 1 3390
box -12 -8 72 272
use XOR2X1  _1094_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform 1 0 3830 0 1 3390
box -12 -8 132 272
use NAND2X1  _1095_
timestamp 1702508443
transform 1 0 4290 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1096_
timestamp 1702508443
transform 1 0 4150 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1097_
timestamp 1702508443
transform 1 0 1790 0 -1 2350
box -12 -8 72 272
use NAND2X1  _1098_
timestamp 1702508443
transform 1 0 3130 0 1 3390
box -12 -8 72 272
use NAND2X1  _1099_
timestamp 1702508443
transform 1 0 2750 0 1 3390
box -12 -8 72 272
use OAI21X1  _1100_
timestamp 1702508443
transform -1 0 2690 0 1 3390
box -12 -8 92 272
use AOI21X1  _1101_
timestamp 1702508443
transform -1 0 2570 0 1 4950
box -12 -8 92 272
use OAI21X1  _1102_
timestamp 1702508443
transform -1 0 2270 0 -1 4950
box -12 -8 92 272
use NAND2X1  _1103_
timestamp 1702508443
transform 1 0 1830 0 1 4430
box -12 -8 72 272
use INVX1  _1104_
timestamp 1701862152
transform -1 0 550 0 1 4430
box -12 -8 52 272
use INVX1  _1105_
timestamp 1701862152
transform -1 0 2150 0 1 4950
box -12 -8 52 272
use AOI21X1  _1106_
timestamp 1702508443
transform -1 0 2050 0 1 4950
box -12 -8 92 272
use INVX2  _1107_
timestamp 1701862152
transform -1 0 2010 0 -1 4430
box -12 -8 52 272
use NOR2X1  _1108_
timestamp 1701862152
transform -1 0 1510 0 -1 4430
box -12 -8 74 272
use AND2X2  _1109_
timestamp 1701862152
transform -1 0 1630 0 1 4430
box -12 -8 94 272
use AOI22X1  _1110_
timestamp 1701862152
transform -1 0 1390 0 -1 4430
box -14 -8 114 272
use AOI21X1  _1111_
timestamp 1702508443
transform -1 0 1230 0 -1 4430
box -12 -8 92 272
use XNOR2X1  _1112_
timestamp 1702508443
transform -1 0 930 0 1 4430
box -12 -8 132 272
use AOI21X1  _1113_
timestamp 1702508443
transform -1 0 810 0 -1 5470
box -12 -8 92 272
use NAND2X1  _1114_
timestamp 1702508443
transform 1 0 1410 0 1 4430
box -12 -8 72 272
use NAND2X1  _1115_
timestamp 1702508443
transform -1 0 1210 0 1 3910
box -12 -8 72 272
use NAND2X1  _1116_
timestamp 1702508443
transform -1 0 1350 0 1 4430
box -12 -8 72 272
use OAI21X1  _1117_
timestamp 1702508443
transform -1 0 1230 0 1 4430
box -12 -8 92 272
use OAI21X1  _1118_
timestamp 1702508443
transform -1 0 1070 0 1 4430
box -12 -8 92 272
use NOR2X1  _1119_
timestamp 1701862152
transform -1 0 670 0 -1 5470
box -12 -8 74 272
use OAI21X1  _1120_
timestamp 1702508443
transform -1 0 1250 0 1 4950
box -12 -8 92 272
use XOR2X1  _1121_
timestamp 1702508443
transform -1 0 1170 0 -1 4950
box -12 -8 132 272
use NOR2X1  _1122_
timestamp 1701862152
transform -1 0 1110 0 1 4950
box -12 -8 74 272
use OAI21X1  _1123_
timestamp 1702508443
transform -1 0 850 0 1 4950
box -12 -8 92 272
use XOR2X1  _1124_
timestamp 1702508443
transform -1 0 750 0 1 4430
box -12 -8 132 272
use OAI21X1  _1125_
timestamp 1702508443
transform 1 0 910 0 1 4950
box -12 -8 92 272
use NAND2X1  _1126_
timestamp 1702508443
transform -1 0 410 0 -1 5470
box -12 -8 72 272
use NAND3X1  _1127_
timestamp 1702508443
transform -1 0 710 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1128_
timestamp 1702508443
transform -1 0 430 0 1 4950
box -12 -8 92 272
use AOI21X1  _1129_
timestamp 1702508443
transform 1 0 1490 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1130_
timestamp 1702508443
transform -1 0 1650 0 1 4950
box -12 -8 92 272
use AOI21X1  _1131_
timestamp 1702508443
transform -1 0 570 0 1 4950
box -12 -8 92 272
use NAND2X1  _1132_
timestamp 1702508443
transform 1 0 90 0 -1 5470
box -12 -8 72 272
use OAI21X1  _1133_
timestamp 1702508443
transform -1 0 550 0 -1 5470
box -12 -8 92 272
use AOI21X1  _1134_
timestamp 1702508443
transform -1 0 290 0 -1 5470
box -12 -8 92 272
use OAI21X1  _1135_
timestamp 1702508443
transform 1 0 210 0 1 4950
box -12 -8 92 272
use NAND3X1  _1136_
timestamp 1702508443
transform 1 0 210 0 -1 4950
box -12 -8 92 272
use NAND3X1  _1137_
timestamp 1702508443
transform -1 0 430 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1138_
timestamp 1702508443
transform -1 0 150 0 1 4950
box -12 -8 92 272
use NAND3X1  _1139_
timestamp 1702508443
transform -1 0 150 0 1 4430
box -12 -8 92 272
use NAND3X1  _1140_
timestamp 1702508443
transform -1 0 310 0 1 4430
box -12 -8 92 272
use INVX1  _1141_
timestamp 1701862152
transform -1 0 390 0 -1 4430
box -12 -8 52 272
use AOI21X1  _1142_
timestamp 1702508443
transform 1 0 70 0 -1 4430
box -12 -8 92 272
use AOI21X1  _1143_
timestamp 1702508443
transform -1 0 150 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1144_
timestamp 1702508443
transform 1 0 210 0 -1 4430
box -12 -8 92 272
use NAND2X1  _1145_
timestamp 1702508443
transform 1 0 430 0 1 3390
box -12 -8 72 272
use XOR2X1  _1146_
timestamp 1702508443
transform -1 0 1490 0 -1 2870
box -12 -8 132 272
use OAI21X1  _1147_
timestamp 1702508443
transform 1 0 1410 0 -1 2350
box -12 -8 92 272
use INVX1  _1148_
timestamp 1701862152
transform 1 0 210 0 -1 3910
box -12 -8 52 272
use AOI21X1  _1149_
timestamp 1702508443
transform -1 0 390 0 -1 3910
box -12 -8 92 272
use AOI22X1  _1150_
timestamp 1701862152
transform -1 0 1090 0 -1 4430
box -14 -8 114 272
use INVX1  _1151_
timestamp 1701862152
transform 1 0 710 0 -1 3910
box -12 -8 52 272
use OAI21X1  _1152_
timestamp 1702508443
transform -1 0 850 0 -1 4950
box -12 -8 92 272
use NOR2X1  _1153_
timestamp 1701862152
transform -1 0 1870 0 1 3910
box -12 -8 74 272
use NAND2X1  _1154_
timestamp 1702508443
transform 1 0 1550 0 1 3910
box -12 -8 72 272
use NAND2X1  _1155_
timestamp 1702508443
transform 1 0 1390 0 -1 3910
box -12 -8 72 272
use OR2X2  _1156_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform -1 0 1490 0 1 3910
box -12 -8 92 272
use OAI21X1  _1157_
timestamp 1702508443
transform -1 0 1750 0 1 3910
box -12 -8 92 272
use NAND3X1  _1158_
timestamp 1702508443
transform -1 0 1350 0 1 3910
box -12 -8 92 272
use NAND2X1  _1159_
timestamp 1702508443
transform -1 0 1310 0 -1 3910
box -12 -8 72 272
use NAND2X1  _1160_
timestamp 1702508443
transform 1 0 1330 0 1 3390
box -12 -8 72 272
use OAI21X1  _1161_
timestamp 1702508443
transform 1 0 1510 0 -1 3910
box -12 -8 92 272
use OAI21X1  _1162_
timestamp 1702508443
transform -1 0 1750 0 -1 3910
box -12 -8 92 272
use NAND2X1  _1163_
timestamp 1702508443
transform -1 0 1090 0 1 3910
box -12 -8 72 272
use OAI21X1  _1164_
timestamp 1702508443
transform 1 0 890 0 1 3910
box -12 -8 92 272
use NOR2X1  _1165_
timestamp 1701862152
transform -1 0 930 0 -1 4430
box -12 -8 74 272
use NAND3X1  _1166_
timestamp 1702508443
transform -1 0 1030 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1167_
timestamp 1702508443
transform -1 0 890 0 -1 3910
box -12 -8 92 272
use AOI21X1  _1168_
timestamp 1702508443
transform 1 0 630 0 1 4950
box -12 -8 92 272
use AOI21X1  _1169_
timestamp 1702508443
transform -1 0 810 0 -1 4430
box -12 -8 92 272
use INVX1  _1170_
timestamp 1701862152
transform -1 0 690 0 1 3910
box -12 -8 52 272
use OAI21X1  _1171_
timestamp 1702508443
transform 1 0 590 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1172_
timestamp 1702508443
transform -1 0 650 0 -1 3910
box -12 -8 92 272
use NAND3X1  _1173_
timestamp 1702508443
transform -1 0 830 0 1 3910
box -12 -8 92 272
use OAI21X1  _1174_
timestamp 1702508443
transform 1 0 450 0 -1 4430
box -12 -8 92 272
use NAND3X1  _1175_
timestamp 1702508443
transform -1 0 570 0 1 3910
box -12 -8 92 272
use NAND2X1  _1176_
timestamp 1702508443
transform -1 0 290 0 1 3910
box -12 -8 72 272
use NAND3X1  _1177_
timestamp 1702508443
transform 1 0 90 0 1 3910
box -12 -8 92 272
use AOI21X1  _1178_
timestamp 1702508443
transform -1 0 570 0 -1 4950
box -12 -8 92 272
use OAI21X1  _1179_
timestamp 1702508443
transform -1 0 450 0 1 4430
box -12 -8 92 272
use NAND3X1  _1180_
timestamp 1702508443
transform -1 0 430 0 1 3910
box -12 -8 92 272
use AND2X2  _1181_
timestamp 1701862152
transform -1 0 150 0 -1 3910
box -12 -8 94 272
use XOR2X1  _1182_
timestamp 1702508443
transform -1 0 190 0 -1 3390
box -12 -8 132 272
use NAND2X1  _1183_
timestamp 1702508443
transform -1 0 390 0 1 1830
box -12 -8 72 272
use OAI21X1  _1184_
timestamp 1702508443
transform 1 0 190 0 1 1830
box -12 -8 92 272
use INVX1  _1185_
timestamp 1701862152
transform 1 0 90 0 1 270
box -12 -8 52 272
use NAND2X1  _1186_
timestamp 1702508443
transform -1 0 370 0 1 3390
box -12 -8 72 272
use NOR2X1  _1187_
timestamp 1701862152
transform 1 0 350 0 -1 3390
box -12 -8 74 272
use NAND2X1  _1188_
timestamp 1702508443
transform 1 0 70 0 1 3390
box -12 -8 72 272
use NAND2X1  _1189_
timestamp 1702508443
transform -1 0 250 0 1 3390
box -12 -8 72 272
use INVX1  _1190_
timestamp 1701862152
transform 1 0 250 0 -1 3390
box -12 -8 52 272
use AOI21X1  _1191_
timestamp 1702508443
transform 1 0 330 0 1 2870
box -12 -8 92 272
use NAND2X1  _1192_
timestamp 1702508443
transform -1 0 510 0 -1 3910
box -12 -8 72 272
use OAI21X1  _1193_
timestamp 1702508443
transform -1 0 1190 0 -1 3910
box -12 -8 92 272
use INVX1  _1194_
timestamp 1701862152
transform -1 0 1310 0 -1 3390
box -12 -8 52 272
use OR2X2  _1195_
timestamp 1702508443
transform -1 0 990 0 -1 4950
box -12 -8 92 272
use NOR2X1  _1196_
timestamp 1701862152
transform -1 0 1850 0 -1 3390
box -12 -8 74 272
use OAI21X1  _1197_
timestamp 1702508443
transform -1 0 1790 0 1 3390
box -12 -8 92 272
use NAND2X1  _1198_
timestamp 1702508443
transform -1 0 1650 0 1 3390
box -12 -8 72 272
use OAI21X1  _1199_
timestamp 1702508443
transform 1 0 1450 0 1 3390
box -12 -8 92 272
use XOR2X1  _1200_
timestamp 1702508443
transform -1 0 1270 0 1 3390
box -12 -8 132 272
use AOI21X1  _1201_
timestamp 1702508443
transform 1 0 990 0 1 3390
box -12 -8 92 272
use NAND3X1  _1202_
timestamp 1702508443
transform 1 0 850 0 1 3390
box -12 -8 92 272
use INVX1  _1203_
timestamp 1701862152
transform 1 0 1030 0 -1 3390
box -12 -8 52 272
use OAI21X1  _1204_
timestamp 1702508443
transform 1 0 1130 0 -1 3390
box -12 -8 92 272
use INVX1  _1205_
timestamp 1701862152
transform -1 0 950 0 1 2870
box -12 -8 52 272
use NAND3X1  _1206_
timestamp 1702508443
transform -1 0 970 0 -1 3390
box -12 -8 92 272
use AND2X2  _1207_
timestamp 1701862152
transform -1 0 830 0 -1 3390
box -12 -8 94 272
use NAND2X1  _1208_
timestamp 1702508443
transform 1 0 630 0 -1 3390
box -12 -8 72 272
use OR2X2  _1209_
timestamp 1702508443
transform -1 0 550 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1210_
timestamp 1702508443
transform 1 0 210 0 1 2870
box -12 -8 72 272
use NAND2X1  _1211_
timestamp 1702508443
transform 1 0 430 0 -1 2870
box -12 -8 72 272
use AND2X2  _1212_
timestamp 1701862152
transform 1 0 2990 0 1 3390
box -12 -8 94 272
use NAND3X1  _1213_
timestamp 1702508443
transform -1 0 3610 0 1 3390
box -12 -8 92 272
use NAND3X1  _1214_
timestamp 1702508443
transform 1 0 550 0 1 3390
box -12 -8 92 272
use AOI21X1  _1215_
timestamp 1702508443
transform -1 0 790 0 1 3390
box -12 -8 92 272
use INVX1  _1216_
timestamp 1701862152
transform -1 0 230 0 -1 2870
box -12 -8 52 272
use OAI21X1  _1217_
timestamp 1702508443
transform -1 0 370 0 -1 2870
box -12 -8 92 272
use NAND3X1  _1218_
timestamp 1702508443
transform -1 0 390 0 1 2350
box -12 -8 92 272
use OAI21X1  _1219_
timestamp 1702508443
transform 1 0 190 0 1 270
box -12 -8 92 272
use NAND2X1  _1220_
timestamp 1702508443
transform 1 0 310 0 -1 1830
box -12 -8 72 272
use AOI21X1  _1221_
timestamp 1702508443
transform -1 0 1090 0 1 2870
box -12 -8 92 272
use INVX1  _1222_
timestamp 1701862152
transform 1 0 1550 0 -1 3390
box -12 -8 52 272
use OAI22X1  _1223_
timestamp 1701862152
transform 1 0 1390 0 -1 3390
box -12 -8 112 272
use OAI21X1  _1224_
timestamp 1702508443
transform -1 0 1730 0 -1 3390
box -12 -8 92 272
use NOR2X1  _1225_
timestamp 1701862152
transform -1 0 1970 0 -1 3390
box -12 -8 74 272
use INVX1  _1226_
timestamp 1701862152
transform -1 0 1990 0 -1 2870
box -12 -8 52 272
use OR2X2  _1227_
timestamp 1702508443
transform -1 0 1750 0 -1 2870
box -12 -8 92 272
use AND2X2  _1228_
timestamp 1701862152
transform -1 0 1630 0 1 2870
box -12 -8 94 272
use XNOR2X1  _1229_
timestamp 1702508443
transform 1 0 1150 0 1 2870
box -12 -8 132 272
use XOR2X1  _1230_
timestamp 1702508443
transform -1 0 850 0 1 2870
box -12 -8 132 272
use INVX1  _1231_
timestamp 1701862152
transform 1 0 70 0 1 2350
box -12 -8 52 272
use NAND3X1  _1232_
timestamp 1702508443
transform -1 0 250 0 1 2350
box -12 -8 92 272
use OAI21X1  _1233_
timestamp 1702508443
transform -1 0 150 0 1 2870
box -12 -8 92 272
use NAND2X1  _1234_
timestamp 1702508443
transform 1 0 70 0 -1 2870
box -12 -8 72 272
use NAND3X1  _1235_
timestamp 1702508443
transform -1 0 150 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1236_
timestamp 1702508443
transform -1 0 130 0 1 1830
box -12 -8 72 272
use INVX1  _1237_
timestamp 1701862152
transform -1 0 250 0 -1 2350
box -12 -8 52 272
use NOR2X1  _1238_
timestamp 1701862152
transform -1 0 1310 0 -1 2870
box -12 -8 74 272
use AOI21X1  _1239_
timestamp 1702508443
transform 1 0 970 0 -1 2870
box -12 -8 92 272
use NOR2X1  _1240_
timestamp 1701862152
transform -1 0 1170 0 -1 2870
box -12 -8 74 272
use NAND3X1  _1241_
timestamp 1702508443
transform 1 0 470 0 1 2870
box -12 -8 92 272
use OAI21X1  _1242_
timestamp 1702508443
transform 1 0 830 0 -1 2870
box -12 -8 92 272
use NAND2X1  _1243_
timestamp 1702508443
transform 1 0 1330 0 1 2870
box -12 -8 72 272
use OAI21X1  _1244_
timestamp 1702508443
transform 1 0 1790 0 1 2870
box -12 -8 92 272
use OR2X2  _1245_
timestamp 1702508443
transform 1 0 1810 0 -1 2870
box -12 -8 92 272
use INVX1  _1246_
timestamp 1701862152
transform -1 0 1610 0 -1 2870
box -12 -8 52 272
use OAI21X1  _1247_
timestamp 1702508443
transform 1 0 1250 0 1 2350
box -12 -8 92 272
use AND2X2  _1248_
timestamp 1701862152
transform -1 0 1190 0 1 2350
box -12 -8 94 272
use NOR2X1  _1249_
timestamp 1701862152
transform 1 0 710 0 1 2350
box -12 -8 74 272
use INVX1  _1250_
timestamp 1701862152
transform -1 0 650 0 1 2870
box -12 -8 52 272
use OAI21X1  _1251_
timestamp 1702508443
transform 1 0 690 0 -1 2870
box -12 -8 92 272
use AOI21X1  _1252_
timestamp 1702508443
transform 1 0 550 0 -1 2870
box -12 -8 92 272
use INVX1  _1253_
timestamp 1701862152
transform -1 0 650 0 1 2350
box -12 -8 52 272
use OAI21X1  _1254_
timestamp 1702508443
transform -1 0 530 0 1 2350
box -12 -8 92 272
use OAI22X1  _1255_
timestamp 1701862152
transform 1 0 550 0 -1 2350
box -12 -8 112 272
use INVX1  _1256_
timestamp 1701862152
transform 1 0 790 0 1 1830
box -12 -8 52 272
use AOI21X1  _1257_
timestamp 1702508443
transform 1 0 830 0 1 2350
box -12 -8 92 272
use AND2X2  _1258_
timestamp 1701862152
transform -1 0 1050 0 1 2350
box -12 -8 94 272
use AOI22X1  _1259_
timestamp 1701862152
transform -1 0 950 0 -1 2350
box -14 -8 114 272
use NOR2X1  _1260_
timestamp 1701862152
transform 1 0 3450 0 -1 1310
box -12 -8 74 272
use INVX1  _1261_
timestamp 1701862152
transform -1 0 3490 0 1 790
box -12 -8 52 272
use NAND2X1  _1262_
timestamp 1702508443
transform 1 0 3330 0 -1 1310
box -12 -8 72 272
use NAND2X1  _1263_
timestamp 1702508443
transform 1 0 3310 0 1 790
box -12 -8 72 272
use NAND2X1  _1264_
timestamp 1702508443
transform -1 0 3270 0 -1 790
box -12 -8 72 272
use OAI21X1  _1265_
timestamp 1702508443
transform 1 0 3330 0 -1 790
box -12 -8 92 272
use INVX1  _1266_
timestamp 1701862152
transform 1 0 4310 0 -1 1310
box -12 -8 52 272
use NOR2X1  _1267_
timestamp 1701862152
transform 1 0 4050 0 1 790
box -12 -8 74 272
use NOR2X1  _1268_
timestamp 1701862152
transform 1 0 4090 0 -1 1310
box -12 -8 74 272
use NOR2X1  _1269_
timestamp 1701862152
transform 1 0 3670 0 1 790
box -12 -8 74 272
use NAND2X1  _1270_
timestamp 1702508443
transform 1 0 3550 0 1 790
box -12 -8 72 272
use OAI21X1  _1271_
timestamp 1702508443
transform -1 0 3870 0 1 790
box -12 -8 92 272
use NAND2X1  _1272_
timestamp 1702508443
transform 1 0 3930 0 1 790
box -12 -8 72 272
use NAND2X1  _1273_
timestamp 1702508443
transform -1 0 4410 0 -1 270
box -12 -8 72 272
use OAI21X1  _1274_
timestamp 1702508443
transform 1 0 4310 0 1 270
box -12 -8 92 272
use OAI21X1  _1275_
timestamp 1702508443
transform -1 0 4250 0 1 790
box -12 -8 92 272
use XOR2X1  _1276_
timestamp 1702508443
transform -1 0 5370 0 -1 790
box -12 -8 132 272
use XNOR2X1  _1277_
timestamp 1702508443
transform 1 0 5230 0 1 790
box -12 -8 132 272
use NAND2X1  _1278_
timestamp 1702508443
transform 1 0 5730 0 -1 270
box -12 -8 72 272
use OAI21X1  _1279_
timestamp 1702508443
transform 1 0 5710 0 1 270
box -12 -8 92 272
use NOR2X1  _1280_
timestamp 1701862152
transform -1 0 5030 0 1 790
box -12 -8 74 272
use AOI21X1  _1281_
timestamp 1702508443
transform 1 0 5090 0 1 790
box -12 -8 92 272
use NOR2X1  _1282_
timestamp 1701862152
transform -1 0 5810 0 -1 3910
box -12 -8 74 272
use NOR2X1  _1283_
timestamp 1701862152
transform -1 0 5730 0 -1 2350
box -12 -8 74 272
use NOR2X1  _1284_
timestamp 1701862152
transform -1 0 5810 0 -1 1310
box -12 -8 74 272
use XOR2X1  _1285_
timestamp 1702508443
transform 1 0 5550 0 1 790
box -12 -8 132 272
use NAND2X1  _1286_
timestamp 1702508443
transform 1 0 5370 0 -1 270
box -12 -8 72 272
use OAI21X1  _1287_
timestamp 1702508443
transform -1 0 5650 0 1 270
box -12 -8 92 272
use NAND2X1  _1288_
timestamp 1702508443
transform 1 0 4110 0 -1 790
box -12 -8 72 272
use NAND2X1  _1289_
timestamp 1702508443
transform 1 0 5250 0 -1 1830
box -12 -8 72 272
use NAND2X1  _1290_
timestamp 1702508443
transform 1 0 5370 0 1 1830
box -12 -8 72 272
use AND2X2  _1291_
timestamp 1701862152
transform -1 0 5190 0 -1 1830
box -12 -8 94 272
use INVX1  _1292_
timestamp 1701862152
transform 1 0 4970 0 1 1310
box -12 -8 52 272
use INVX1  _1293_
timestamp 1701862152
transform -1 0 5730 0 1 1310
box -12 -8 52 272
use OAI21X1  _1294_
timestamp 1702508443
transform -1 0 5630 0 1 1310
box -12 -8 92 272
use INVX1  _1295_
timestamp 1701862152
transform -1 0 5230 0 1 1310
box -12 -8 52 272
use NAND2X1  _1296_
timestamp 1702508443
transform 1 0 5070 0 1 1310
box -12 -8 72 272
use NAND2X1  _1297_
timestamp 1702508443
transform 1 0 5290 0 1 1310
box -12 -8 72 272
use NAND2X1  _1298_
timestamp 1702508443
transform -1 0 5110 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1299_
timestamp 1702508443
transform -1 0 4330 0 -1 790
box -12 -8 92 272
use NAND2X1  _1300_
timestamp 1702508443
transform 1 0 5210 0 1 270
box -12 -8 72 272
use OAI21X1  _1301_
timestamp 1702508443
transform 1 0 5410 0 1 1310
box -12 -8 92 272
use OR2X2  _1302_
timestamp 1702508443
transform 1 0 5350 0 -1 2350
box -12 -8 92 272
use NAND2X1  _1303_
timestamp 1702508443
transform 1 0 5230 0 -1 2350
box -12 -8 72 272
use AND2X2  _1304_
timestamp 1701862152
transform -1 0 5310 0 1 1830
box -12 -8 94 272
use NOR2X1  _1305_
timestamp 1701862152
transform 1 0 5510 0 -1 1310
box -12 -8 74 272
use INVX1  _1306_
timestamp 1701862152
transform 1 0 5650 0 -1 1310
box -12 -8 52 272
use INVX1  _1307_
timestamp 1701862152
transform -1 0 5210 0 -1 1310
box -12 -8 52 272
use OAI21X1  _1308_
timestamp 1702508443
transform 1 0 5270 0 -1 1310
box -12 -8 92 272
use OAI21X1  _1309_
timestamp 1702508443
transform -1 0 5490 0 1 790
box -12 -8 92 272
use NAND2X1  _1310_
timestamp 1702508443
transform -1 0 4570 0 -1 790
box -12 -8 72 272
use OAI21X1  _1311_
timestamp 1702508443
transform -1 0 4990 0 -1 1310
box -12 -8 92 272
use XOR2X1  _1312_
timestamp 1702508443
transform 1 0 4290 0 1 1830
box -12 -8 132 272
use NOR2X1  _1313_
timestamp 1701862152
transform 1 0 4790 0 -1 1310
box -12 -8 74 272
use NAND2X1  _1314_
timestamp 1702508443
transform 1 0 4670 0 -1 1310
box -12 -8 72 272
use NAND2X1  _1315_
timestamp 1702508443
transform -1 0 4770 0 1 790
box -12 -8 72 272
use OAI21X1  _1316_
timestamp 1702508443
transform -1 0 4650 0 1 790
box -12 -8 92 272
use OAI21X1  _1317_
timestamp 1702508443
transform 1 0 3970 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1318_
timestamp 1701862152
transform 1 0 4410 0 -1 2350
box -12 -8 74 272
use NAND2X1  _1319_
timestamp 1702508443
transform -1 0 4590 0 -1 2350
box -12 -8 72 272
use INVX1  _1320_
timestamp 1701862152
transform 1 0 4650 0 -1 2350
box -12 -8 52 272
use NOR2X1  _1321_
timestamp 1701862152
transform 1 0 4750 0 1 1830
box -12 -8 74 272
use XNOR2X1  _1322_
timestamp 1702508443
transform 1 0 4010 0 1 1310
box -12 -8 132 272
use NAND2X1  _1323_
timestamp 1702508443
transform 1 0 4770 0 -1 270
box -12 -8 72 272
use OAI21X1  _1324_
timestamp 1702508443
transform 1 0 4630 0 -1 270
box -12 -8 92 272
use NAND2X1  _1325_
timestamp 1702508443
transform 1 0 2210 0 1 270
box -12 -8 72 272
use OAI21X1  _1326_
timestamp 1702508443
transform -1 0 5030 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1327_
timestamp 1702508443
transform -1 0 4530 0 1 1830
box -12 -8 72 272
use OAI21X1  _1328_
timestamp 1702508443
transform 1 0 4590 0 1 1830
box -12 -8 92 272
use AND2X2  _1329_
timestamp 1701862152
transform 1 0 4450 0 1 1310
box -12 -8 94 272
use AOI21X1  _1330_
timestamp 1702508443
transform -1 0 4730 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1331_
timestamp 1701862152
transform -1 0 4910 0 1 1310
box -12 -8 74 272
use NAND3X1  _1332_
timestamp 1702508443
transform -1 0 4790 0 1 1310
box -12 -8 92 272
use NAND2X1  _1333_
timestamp 1702508443
transform 1 0 4590 0 1 1310
box -12 -8 72 272
use OR2X2  _1334_
timestamp 1702508443
transform -1 0 1750 0 -1 1830
box -12 -8 92 272
use NAND2X1  _1335_
timestamp 1702508443
transform -1 0 1870 0 -1 1830
box -12 -8 72 272
use AND2X2  _1336_
timestamp 1701862152
transform 1 0 1670 0 1 1310
box -12 -8 94 272
use NOR2X1  _1337_
timestamp 1701862152
transform 1 0 1970 0 -1 790
box -12 -8 74 272
use INVX1  _1338_
timestamp 1701862152
transform 1 0 1910 0 1 790
box -12 -8 52 272
use INVX1  _1339_
timestamp 1701862152
transform -1 0 1910 0 -1 790
box -12 -8 52 272
use OAI21X1  _1340_
timestamp 1702508443
transform -1 0 1850 0 1 790
box -12 -8 92 272
use OAI21X1  _1341_
timestamp 1702508443
transform 1 0 2070 0 1 270
box -12 -8 92 272
use OAI21X1  _1342_
timestamp 1702508443
transform -1 0 1710 0 1 790
box -12 -8 92 272
use NOR2X1  _1343_
timestamp 1701862152
transform -1 0 1090 0 1 790
box -12 -8 74 272
use NAND2X1  _1344_
timestamp 1702508443
transform -1 0 970 0 1 790
box -12 -8 72 272
use INVX1  _1345_
timestamp 1701862152
transform 1 0 1150 0 1 790
box -12 -8 52 272
use NOR2X1  _1346_
timestamp 1701862152
transform -1 0 1310 0 1 790
box -12 -8 74 272
use INVX1  _1347_
timestamp 1701862152
transform 1 0 1310 0 -1 790
box -12 -8 52 272
use XOR2X1  _1348_
timestamp 1702508443
transform 1 0 1690 0 -1 790
box -12 -8 132 272
use NAND2X1  _1349_
timestamp 1702508443
transform -1 0 2530 0 -1 790
box -12 -8 72 272
use OAI21X1  _1350_
timestamp 1702508443
transform 1 0 2090 0 -1 790
box -12 -8 92 272
use NAND2X1  _1351_
timestamp 1702508443
transform -1 0 2770 0 1 270
box -12 -8 72 272
use NOR2X1  _1352_
timestamp 1701862152
transform 1 0 1570 0 -1 790
box -12 -8 74 272
use OAI21X1  _1353_
timestamp 1702508443
transform -1 0 1450 0 1 790
box -12 -8 92 272
use AOI21X1  _1354_
timestamp 1702508443
transform -1 0 1490 0 -1 790
box -12 -8 92 272
use NOR2X1  _1355_
timestamp 1701862152
transform -1 0 370 0 -1 270
box -12 -8 74 272
use NOR2X1  _1356_
timestamp 1701862152
transform -1 0 490 0 -1 270
box -12 -8 74 272
use NOR2X1  _1357_
timestamp 1701862152
transform 1 0 330 0 1 270
box -12 -8 74 272
use INVX1  _1358_
timestamp 1701862152
transform 1 0 450 0 1 270
box -12 -8 52 272
use AND2X2  _1359_
timestamp 1701862152
transform 1 0 1930 0 1 270
box -12 -8 94 272
use OAI21X1  _1360_
timestamp 1702508443
transform -1 0 1850 0 1 270
box -12 -8 92 272
use OAI21X1  _1361_
timestamp 1702508443
transform 1 0 2330 0 1 270
box -12 -8 92 272
use NOR2X1  _1362_
timestamp 1701862152
transform -1 0 1330 0 1 270
box -12 -8 74 272
use NOR2X1  _1363_
timestamp 1701862152
transform 1 0 1150 0 1 270
box -12 -8 74 272
use NOR2X1  _1364_
timestamp 1701862152
transform -1 0 850 0 1 1310
box -12 -8 74 272
use NAND2X1  _1365_
timestamp 1702508443
transform -1 0 730 0 1 1310
box -12 -8 72 272
use INVX1  _1366_
timestamp 1701862152
transform 1 0 670 0 -1 1310
box -12 -8 52 272
use NOR2X1  _1367_
timestamp 1701862152
transform -1 0 770 0 -1 790
box -12 -8 74 272
use XOR2X1  _1368_
timestamp 1702508443
transform -1 0 1090 0 1 270
box -12 -8 132 272
use NAND2X1  _1369_
timestamp 1702508443
transform -1 0 1590 0 1 270
box -12 -8 72 272
use OAI21X1  _1370_
timestamp 1702508443
transform 1 0 1390 0 1 270
box -12 -8 92 272
use NAND2X1  _1371_
timestamp 1702508443
transform 1 0 570 0 -1 790
box -12 -8 72 272
use AOI21X1  _1372_
timestamp 1702508443
transform -1 0 910 0 1 270
box -12 -8 92 272
use NAND2X1  _1373_
timestamp 1702508443
transform -1 0 610 0 1 270
box -12 -8 72 272
use OAI21X1  _1374_
timestamp 1702508443
transform 1 0 690 0 1 270
box -12 -8 92 272
use NAND2X1  _1375_
timestamp 1702508443
transform -1 0 270 0 1 1310
box -12 -8 72 272
use NOR2X1  _1376_
timestamp 1701862152
transform 1 0 430 0 -1 1830
box -12 -8 74 272
use INVX1  _1377_
timestamp 1701862152
transform -1 0 370 0 1 1310
box -12 -8 52 272
use AND2X2  _1378_
timestamp 1701862152
transform -1 0 150 0 1 1310
box -12 -8 94 272
use NOR2X1  _1379_
timestamp 1701862152
transform 1 0 70 0 -1 790
box -12 -8 74 272
use INVX1  _1380_
timestamp 1701862152
transform 1 0 70 0 1 790
box -12 -8 52 272
use INVX1  _1381_
timestamp 1701862152
transform 1 0 70 0 -1 1310
box -12 -8 52 272
use OAI21X1  _1382_
timestamp 1702508443
transform 1 0 190 0 1 790
box -12 -8 92 272
use OAI21X1  _1383_
timestamp 1702508443
transform 1 0 190 0 -1 790
box -12 -8 92 272
use OAI21X1  _1384_
timestamp 1702508443
transform 1 0 170 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1385_
timestamp 1701862152
transform -1 0 950 0 1 1830
box -12 -8 74 272
use NOR2X1  _1386_
timestamp 1701862152
transform -1 0 970 0 -1 1830
box -12 -8 74 272
use NOR2X1  _1387_
timestamp 1701862152
transform -1 0 850 0 -1 1830
box -12 -8 74 272
use INVX1  _1388_
timestamp 1701862152
transform -1 0 610 0 1 1310
box -12 -8 52 272
use OR2X2  _1389_
timestamp 1702508443
transform 1 0 350 0 1 790
box -12 -8 92 272
use AOI21X1  _1390_
timestamp 1702508443
transform 1 0 490 0 1 790
box -12 -8 92 272
use AOI22X1  _1391_
timestamp 1701862152
transform -1 0 730 0 1 790
box -14 -8 114 272
use AOI21X1  _1392_
timestamp 1702508443
transform -1 0 510 0 1 1310
box -12 -8 92 272
use INVX1  _1393_
timestamp 1701862152
transform 1 0 430 0 -1 1310
box -12 -8 52 272
use NOR2X1  _1394_
timestamp 1701862152
transform -1 0 370 0 -1 1310
box -12 -8 74 272
use AOI21X1  _1395_
timestamp 1702508443
transform 1 0 530 0 -1 1310
box -12 -8 92 272
use INVX1  _1396_
timestamp 1701862152
transform 1 0 910 0 1 1310
box -12 -8 52 272
use NOR2X1  _1397_
timestamp 1701862152
transform -1 0 1090 0 1 1310
box -12 -8 74 272
use OAI21X1  _1398_
timestamp 1702508443
transform -1 0 1350 0 -1 1310
box -12 -8 92 272
use OAI22X1  _1399_
timestamp 1701862152
transform -1 0 1210 0 -1 1310
box -12 -8 112 272
use NAND2X1  _1400_
timestamp 1702508443
transform -1 0 1630 0 -1 1310
box -12 -8 72 272
use NAND3X1  _1401_
timestamp 1702508443
transform 1 0 1150 0 1 1310
box -12 -8 92 272
use OAI21X1  _1402_
timestamp 1702508443
transform 1 0 1290 0 1 1310
box -12 -8 92 272
use NAND2X1  _1403_
timestamp 1702508443
transform 1 0 1430 0 1 1310
box -12 -8 72 272
use OAI21X1  _1404_
timestamp 1702508443
transform 1 0 1430 0 -1 1310
box -12 -8 92 272
use INVX1  _1405_
timestamp 1701862152
transform -1 0 3250 0 1 790
box -12 -8 52 272
use NAND3X1  _1406_
timestamp 1702508443
transform 1 0 2490 0 1 790
box -12 -8 92 272
use NAND2X1  _1407_
timestamp 1702508443
transform 1 0 2150 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1408_
timestamp 1702508443
transform -1 0 2350 0 -1 2350
box -12 -8 92 272
use INVX1  _1409_
timestamp 1701862152
transform 1 0 3490 0 -1 270
box -12 -8 52 272
use NAND2X1  _1410_
timestamp 1702508443
transform 1 0 2450 0 -1 1310
box -12 -8 72 272
use OAI21X1  _1411_
timestamp 1702508443
transform -1 0 2650 0 -1 1310
box -12 -8 92 272
use INVX1  _1412_
timestamp 1701862152
transform -1 0 3650 0 -1 270
box -12 -8 52 272
use NAND2X1  _1413_
timestamp 1702508443
transform 1 0 2110 0 1 2350
box -12 -8 72 272
use OAI21X1  _1414_
timestamp 1702508443
transform -1 0 2310 0 1 2350
box -12 -8 92 272
use INVX1  _1415_
timestamp 1701862152
transform -1 0 3790 0 1 270
box -12 -8 52 272
use NAND2X1  _1416_
timestamp 1702508443
transform 1 0 2410 0 -1 2350
box -12 -8 72 272
use OAI21X1  _1417_
timestamp 1702508443
transform -1 0 2690 0 1 2350
box -12 -8 92 272
use NOR2X1  _1418_
timestamp 1701862152
transform 1 0 3250 0 1 270
box -12 -8 74 272
use NOR2X1  _1419_
timestamp 1701862152
transform 1 0 2170 0 -1 1310
box -12 -8 74 272
use AOI21X1  _1420_
timestamp 1702508443
transform -1 0 2390 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1421_
timestamp 1701862152
transform 1 0 2250 0 -1 270
box -12 -8 74 272
use AOI21X1  _1422_
timestamp 1702508443
transform -1 0 2690 0 -1 270
box -12 -8 92 272
use NOR2X1  _1423_
timestamp 1701862152
transform -1 0 2810 0 -1 270
box -12 -8 74 272
use AOI21X1  _1424_
timestamp 1702508443
transform -1 0 3190 0 -1 270
box -12 -8 92 272
use NOR2X1  _1425_
timestamp 1701862152
transform 1 0 2430 0 1 1830
box -12 -8 74 272
use AOI21X1  _1426_
timestamp 1702508443
transform -1 0 2870 0 1 1830
box -12 -8 92 272
use INVX1  _1427_
timestamp 1701862152
transform 1 0 2790 0 -1 2350
box -12 -8 52 272
use OAI21X1  _1428_
timestamp 1702508443
transform 1 0 3170 0 1 1830
box -12 -8 92 272
use OAI21X1  _1429_
timestamp 1702508443
transform 1 0 3310 0 1 1830
box -12 -8 92 272
use OAI21X1  _1430_
timestamp 1702508443
transform 1 0 3290 0 1 2350
box -12 -8 92 272
use OAI21X1  _1431_
timestamp 1702508443
transform -1 0 3490 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1432_
timestamp 1702508443
transform -1 0 3350 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1433_
timestamp 1702508443
transform 1 0 3130 0 -1 2350
box -12 -8 92 272
use OAI21X1  _1434_
timestamp 1702508443
transform -1 0 3230 0 1 2350
box -12 -8 92 272
use OAI21X1  _1435_
timestamp 1702508443
transform 1 0 3010 0 1 2350
box -12 -8 92 272
use NOR2X1  _1436_
timestamp 1701862152
transform 1 0 2790 0 -1 1830
box -12 -8 74 272
use AOI21X1  _1437_
timestamp 1702508443
transform -1 0 2730 0 -1 1830
box -12 -8 92 272
use NOR2X1  _1438_
timestamp 1701862152
transform 1 0 2970 0 -1 1310
box -12 -8 74 272
use AOI21X1  _1439_
timestamp 1702508443
transform 1 0 2830 0 -1 1310
box -12 -8 92 272
use NOR2X1  _1440_
timestamp 1701862152
transform -1 0 3950 0 1 1310
box -12 -8 74 272
use AOI21X1  _1441_
timestamp 1702508443
transform 1 0 3510 0 1 1310
box -12 -8 92 272
use NOR2X1  _1442_
timestamp 1701862152
transform 1 0 3570 0 -1 2870
box -12 -8 74 272
use AOI21X1  _1443_
timestamp 1702508443
transform -1 0 3510 0 1 2350
box -12 -8 92 272
use NAND2X1  _1444_
timestamp 1702508443
transform -1 0 2550 0 1 3390
box -12 -8 72 272
use OAI21X1  _1445_
timestamp 1702508443
transform -1 0 2730 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1446_
timestamp 1702508443
transform -1 0 2950 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1447_
timestamp 1702508443
transform -1 0 3090 0 -1 3390
box -12 -8 92 272
use NAND2X1  _1448_
timestamp 1702508443
transform -1 0 2490 0 1 2870
box -12 -8 72 272
use OAI21X1  _1449_
timestamp 1702508443
transform -1 0 2870 0 1 2870
box -12 -8 92 272
use NAND2X1  _1450_
timestamp 1702508443
transform -1 0 2110 0 -1 3390
box -12 -8 72 272
use OAI21X1  _1451_
timestamp 1702508443
transform 1 0 1910 0 -1 3910
box -12 -8 92 272
use DFFPOSX1  _1452_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform 1 0 2230 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1453_
timestamp 1702508443
transform -1 0 2030 0 1 3390
box -13 -8 253 272
use DFFPOSX1  _1454_
timestamp 1702508443
transform 1 0 2270 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1455_
timestamp 1702508443
transform -1 0 2110 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1456_
timestamp 1702508443
transform 1 0 3110 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1457_
timestamp 1702508443
transform 1 0 3770 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1458_
timestamp 1702508443
transform -1 0 5730 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1459_
timestamp 1702508443
transform 1 0 5550 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1460_
timestamp 1702508443
transform -1 0 5550 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1461_
timestamp 1702508443
transform 1 0 4690 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1462_
timestamp 1702508443
transform 1 0 3570 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1463_
timestamp 1702508443
transform 1 0 3930 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1464_
timestamp 1702508443
transform -1 0 2130 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1465_
timestamp 1702508443
transform -1 0 1310 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1466_
timestamp 1702508443
transform -1 0 830 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1467_
timestamp 1702508443
transform -1 0 1990 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1468_
timestamp 1702508443
transform -1 0 730 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1469_
timestamp 1702508443
transform -1 0 1290 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1470_
timestamp 1702508443
transform -1 0 1450 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1471_
timestamp 1702508443
transform -1 0 1630 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1472_
timestamp 1702508443
transform 1 0 3090 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1473_
timestamp 1702508443
transform -1 0 4590 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1474_
timestamp 1702508443
transform 1 0 4830 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1475_
timestamp 1702508443
transform 1 0 5290 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1476_
timestamp 1702508443
transform -1 0 5770 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1477_
timestamp 1702508443
transform 1 0 4270 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1478_
timestamp 1702508443
transform 1 0 3890 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1479_
timestamp 1702508443
transform 1 0 3850 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1480_
timestamp 1702508443
transform 1 0 1490 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1481_
timestamp 1702508443
transform 1 0 490 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1482_
timestamp 1702508443
transform -1 0 250 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1483_
timestamp 1702508443
transform 1 0 10 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1484_
timestamp 1702508443
transform -1 0 490 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1485_
timestamp 1702508443
transform -1 0 1190 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1486_
timestamp 1702508443
transform 1 0 3410 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1487_
timestamp 1702508443
transform -1 0 4630 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1488_
timestamp 1702508443
transform -1 0 5310 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1489_
timestamp 1702508443
transform -1 0 5670 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1490_
timestamp 1702508443
transform -1 0 4050 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1491_
timestamp 1702508443
transform -1 0 5510 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1492_
timestamp 1702508443
transform -1 0 5030 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1493_
timestamp 1702508443
transform -1 0 5070 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1494_
timestamp 1702508443
transform 1 0 1950 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1495_
timestamp 1702508443
transform 1 0 2170 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1496_
timestamp 1702508443
transform 1 0 2410 0 1 270
box -13 -8 253 272
use DFFPOSX1  _1497_
timestamp 1702508443
transform 1 0 1010 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1498_
timestamp 1702508443
transform 1 0 270 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1499_
timestamp 1702508443
transform -1 0 1010 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1500_
timestamp 1702508443
transform 1 0 710 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1501_
timestamp 1702508443
transform 1 0 1630 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1502_
timestamp 1702508443
transform -1 0 2090 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1503_
timestamp 1702508443
transform -1 0 2610 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1504_
timestamp 1702508443
transform -1 0 2050 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1505_
timestamp 1702508443
transform -1 0 2710 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1506_
timestamp 1702508443
transform 1 0 1870 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1507_
timestamp 1702508443
transform -1 0 2550 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1508_
timestamp 1702508443
transform -1 0 3050 0 -1 270
box -13 -8 253 272
use DFFPOSX1  _1509_
timestamp 1702508443
transform -1 0 2730 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1510_
timestamp 1702508443
transform 1 0 3650 0 1 1830
box -13 -8 253 272
use DFFPOSX1  _1511_
timestamp 1702508443
transform 1 0 3490 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1512_
timestamp 1702508443
transform 1 0 2830 0 -1 2350
box -13 -8 253 272
use DFFPOSX1  _1513_
timestamp 1702508443
transform 1 0 2690 0 1 2350
box -13 -8 253 272
use DFFPOSX1  _1514_
timestamp 1702508443
transform -1 0 2590 0 -1 1830
box -13 -8 253 272
use DFFPOSX1  _1515_
timestamp 1702508443
transform -1 0 3270 0 -1 1310
box -13 -8 253 272
use DFFPOSX1  _1516_
timestamp 1702508443
transform 1 0 3590 0 1 1310
box -13 -8 253 272
use DFFPOSX1  _1517_
timestamp 1702508443
transform 1 0 3250 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1518_
timestamp 1702508443
transform 1 0 2510 0 -1 2870
box -13 -8 253 272
use DFFPOSX1  _1519_
timestamp 1702508443
transform 1 0 2870 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1520_
timestamp 1702508443
transform -1 0 2730 0 1 2870
box -13 -8 253 272
use DFFPOSX1  _1521_
timestamp 1702508443
transform 1 0 1990 0 -1 3910
box -13 -8 253 272
use DFFPOSX1  _1522_
timestamp 1702508443
transform 1 0 2230 0 -1 3390
box -13 -8 253 272
use DFFPOSX1  _1523_
timestamp 1702508443
transform -1 0 3150 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1524_
timestamp 1702508443
transform -1 0 2910 0 1 790
box -13 -8 253 272
use DFFPOSX1  _1525_
timestamp 1702508443
transform -1 0 2770 0 -1 790
box -13 -8 253 272
use DFFPOSX1  _1526_
timestamp 1702508443
transform -1 0 2430 0 1 790
box -13 -8 253 272
use BUFX2  _1527_ ~/ETRI050_DesignKit/digital_ETRI
timestamp 1702508443
transform 1 0 5730 0 1 790
box -12 -8 72 272
use BUFX2  _1528_
timestamp 1702508443
transform -1 0 5790 0 1 2870
box -12 -8 72 272
use BUFX2  _1529_
timestamp 1702508443
transform 1 0 5430 0 -1 3390
box -12 -8 72 272
use BUFX2  _1530_
timestamp 1702508443
transform 1 0 5170 0 1 2870
box -12 -8 72 272
use BUFX2  _1531_
timestamp 1702508443
transform 1 0 2810 0 -1 3910
box -12 -8 72 272
use BUFX2  _1532_
timestamp 1702508443
transform 1 0 3870 0 -1 270
box -12 -8 72 272
use BUFX2  _1533_
timestamp 1702508443
transform 1 0 4110 0 -1 270
box -12 -8 72 272
use BUFX2  _1534_
timestamp 1702508443
transform 1 0 4230 0 -1 270
box -12 -8 72 272
use BUFX2  _1535_
timestamp 1702508443
transform 1 0 3990 0 -1 270
box -12 -8 72 272
use BUFX2  BUFX2_insert0
timestamp 1702508443
transform -1 0 1570 0 1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert1
timestamp 1702508443
transform 1 0 2190 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert2
timestamp 1702508443
transform 1 0 4830 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert3
timestamp 1702508443
transform 1 0 3730 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert4
timestamp 1702508443
transform 1 0 2190 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert5
timestamp 1702508443
transform 1 0 4190 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert6
timestamp 1702508443
transform -1 0 1450 0 1 2350
box -12 -8 72 272
use BUFX2  BUFX2_insert15
timestamp 1702508443
transform -1 0 4830 0 1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert16
timestamp 1702508443
transform -1 0 3610 0 -1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert17
timestamp 1702508443
transform -1 0 4050 0 -1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert18
timestamp 1702508443
transform 1 0 4970 0 -1 5470
box -12 -8 72 272
use BUFX2  BUFX2_insert19
timestamp 1702508443
transform -1 0 1710 0 1 270
box -12 -8 72 272
use BUFX2  BUFX2_insert20
timestamp 1702508443
transform -1 0 4450 0 -1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert21
timestamp 1702508443
transform -1 0 1890 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert22
timestamp 1702508443
transform -1 0 4930 0 1 1830
box -12 -8 72 272
use BUFX2  BUFX2_insert23
timestamp 1702508443
transform -1 0 3150 0 -1 790
box -12 -8 72 272
use BUFX2  BUFX2_insert24
timestamp 1702508443
transform 1 0 5090 0 1 270
box -12 -8 72 272
use BUFX2  BUFX2_insert25
timestamp 1702508443
transform -1 0 3110 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert26
timestamp 1702508443
transform 1 0 3070 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert27
timestamp 1702508443
transform 1 0 3190 0 -1 2870
box -12 -8 72 272
use BUFX2  BUFX2_insert28
timestamp 1702508443
transform 1 0 2670 0 1 1310
box -12 -8 72 272
use BUFX2  BUFX2_insert29
timestamp 1702508443
transform -1 0 2590 0 -1 3390
box -12 -8 72 272
use BUFX2  BUFX2_insert30
timestamp 1702508443
transform -1 0 4430 0 -1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert31
timestamp 1702508443
transform -1 0 3570 0 1 4430
box -12 -8 72 272
use BUFX2  BUFX2_insert32
timestamp 1702508443
transform 1 0 4650 0 1 4950
box -12 -8 72 272
use BUFX2  BUFX2_insert33
timestamp 1702508443
transform -1 0 4490 0 1 4430
box -12 -8 72 272
use CLKBUF1  CLKBUF1_insert7 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701862152
transform -1 0 2990 0 -1 2870
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert8
timestamp 1701862152
transform -1 0 1810 0 1 2350
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert9
timestamp 1701862152
transform -1 0 1950 0 -1 270
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert10
timestamp 1701862152
transform -1 0 2550 0 1 2350
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert11
timestamp 1701862152
transform 1 0 4330 0 1 790
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert12
timestamp 1701862152
transform -1 0 3430 0 -1 270
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert13
timestamp 1701862152
transform 1 0 2910 0 -1 1830
box -12 -8 192 272
use CLKBUF1  CLKBUF1_insert14
timestamp 1701862152
transform 1 0 4990 0 1 1830
box -12 -8 192 272
use FILL  FILL85650x62550 ~/ETRI050_DesignKit/digital_ETRI
timestamp 1701859473
transform -1 0 5730 0 -1 4430
box -12 -8 32 272
use FILL  FILL85650x70350
timestamp 1701859473
transform -1 0 5730 0 -1 4950
box -12 -8 32 272
use FILL  FILL85950x7950
timestamp 1701859473
transform -1 0 5750 0 -1 790
box -12 -8 32 272
use FILL  FILL85950x19650
timestamp 1701859473
transform 1 0 5730 0 1 1310
box -12 -8 32 272
use FILL  FILL85950x31350
timestamp 1701859473
transform -1 0 5750 0 -1 2350
box -12 -8 32 272
use FILL  FILL85950x58650
timestamp 1701859473
transform 1 0 5730 0 1 3910
box -12 -8 32 272
use FILL  FILL85950x62550
timestamp 1701859473
transform -1 0 5750 0 -1 4430
box -12 -8 32 272
use FILL  FILL85950x70350
timestamp 1701859473
transform -1 0 5750 0 -1 4950
box -12 -8 32 272
use FILL  FILL85950x74250
timestamp 1701859473
transform 1 0 5730 0 1 4950
box -12 -8 32 272
use FILL  FILL86250x7950
timestamp 1701859473
transform -1 0 5770 0 -1 790
box -12 -8 32 272
use FILL  FILL86250x19650
timestamp 1701859473
transform 1 0 5750 0 1 1310
box -12 -8 32 272
use FILL  FILL86250x31350
timestamp 1701859473
transform -1 0 5770 0 -1 2350
box -12 -8 32 272
use FILL  FILL86250x50850
timestamp 1701859473
transform 1 0 5750 0 1 3390
box -12 -8 32 272
use FILL  FILL86250x58650
timestamp 1701859473
transform 1 0 5750 0 1 3910
box -12 -8 32 272
use FILL  FILL86250x62550
timestamp 1701859473
transform -1 0 5770 0 -1 4430
box -12 -8 32 272
use FILL  FILL86250x70350
timestamp 1701859473
transform -1 0 5770 0 -1 4950
box -12 -8 32 272
use FILL  FILL86250x74250
timestamp 1701859473
transform 1 0 5750 0 1 4950
box -12 -8 32 272
use FILL  FILL86550x7950
timestamp 1701859473
transform -1 0 5790 0 -1 790
box -12 -8 32 272
use FILL  FILL86550x19650
timestamp 1701859473
transform 1 0 5770 0 1 1310
box -12 -8 32 272
use FILL  FILL86550x27450
timestamp 1701859473
transform 1 0 5770 0 1 1830
box -12 -8 32 272
use FILL  FILL86550x31350
timestamp 1701859473
transform -1 0 5790 0 -1 2350
box -12 -8 32 272
use FILL  FILL86550x35250
timestamp 1701859473
transform 1 0 5770 0 1 2350
box -12 -8 32 272
use FILL  FILL86550x46950
timestamp 1701859473
transform -1 0 5790 0 -1 3390
box -12 -8 32 272
use FILL  FILL86550x50850
timestamp 1701859473
transform 1 0 5770 0 1 3390
box -12 -8 32 272
use FILL  FILL86550x58650
timestamp 1701859473
transform 1 0 5770 0 1 3910
box -12 -8 32 272
use FILL  FILL86550x62550
timestamp 1701859473
transform -1 0 5790 0 -1 4430
box -12 -8 32 272
use FILL  FILL86550x70350
timestamp 1701859473
transform -1 0 5790 0 -1 4950
box -12 -8 32 272
use FILL  FILL86550x74250
timestamp 1701859473
transform 1 0 5770 0 1 4950
box -12 -8 32 272
use FILL  FILL86850x150
timestamp 1701859473
transform -1 0 5810 0 -1 270
box -12 -8 32 272
use FILL  FILL86850x4050
timestamp 1701859473
transform 1 0 5790 0 1 270
box -12 -8 32 272
use FILL  FILL86850x7950
timestamp 1701859473
transform -1 0 5810 0 -1 790
box -12 -8 32 272
use FILL  FILL86850x11850
timestamp 1701859473
transform 1 0 5790 0 1 790
box -12 -8 32 272
use FILL  FILL86850x19650
timestamp 1701859473
transform 1 0 5790 0 1 1310
box -12 -8 32 272
use FILL  FILL86850x23550
timestamp 1701859473
transform -1 0 5810 0 -1 1830
box -12 -8 32 272
use FILL  FILL86850x27450
timestamp 1701859473
transform 1 0 5790 0 1 1830
box -12 -8 32 272
use FILL  FILL86850x31350
timestamp 1701859473
transform -1 0 5810 0 -1 2350
box -12 -8 32 272
use FILL  FILL86850x35250
timestamp 1701859473
transform 1 0 5790 0 1 2350
box -12 -8 32 272
use FILL  FILL86850x43050
timestamp 1701859473
transform 1 0 5790 0 1 2870
box -12 -8 32 272
use FILL  FILL86850x46950
timestamp 1701859473
transform -1 0 5810 0 -1 3390
box -12 -8 32 272
use FILL  FILL86850x50850
timestamp 1701859473
transform 1 0 5790 0 1 3390
box -12 -8 32 272
use FILL  FILL86850x58650
timestamp 1701859473
transform 1 0 5790 0 1 3910
box -12 -8 32 272
use FILL  FILL86850x62550
timestamp 1701859473
transform -1 0 5810 0 -1 4430
box -12 -8 32 272
use FILL  FILL86850x70350
timestamp 1701859473
transform -1 0 5810 0 -1 4950
box -12 -8 32 272
use FILL  FILL86850x74250
timestamp 1701859473
transform 1 0 5790 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__723_
timestamp 1701859473
transform -1 0 2790 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__724_
timestamp 1701859473
transform -1 0 2590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__725_
timestamp 1701859473
transform -1 0 2670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__726_
timestamp 1701859473
transform 1 0 3310 0 1 270
box -12 -8 32 272
use FILL  FILL_0__727_
timestamp 1701859473
transform 1 0 2870 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__728_
timestamp 1701859473
transform -1 0 3010 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__729_
timestamp 1701859473
transform 1 0 3650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__730_
timestamp 1701859473
transform 1 0 3550 0 1 270
box -12 -8 32 272
use FILL  FILL_0__731_
timestamp 1701859473
transform -1 0 3470 0 1 270
box -12 -8 32 272
use FILL  FILL_0__732_
timestamp 1701859473
transform -1 0 750 0 1 790
box -12 -8 32 272
use FILL  FILL_0__733_
timestamp 1701859473
transform -1 0 1970 0 1 790
box -12 -8 32 272
use FILL  FILL_0__734_
timestamp 1701859473
transform -1 0 2930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__735_
timestamp 1701859473
transform 1 0 4070 0 1 270
box -12 -8 32 272
use FILL  FILL_0__736_
timestamp 1701859473
transform 1 0 3790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__737_
timestamp 1701859473
transform 1 0 950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__738_
timestamp 1701859473
transform -1 0 2090 0 1 790
box -12 -8 32 272
use FILL  FILL_0__739_
timestamp 1701859473
transform -1 0 2790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__740_
timestamp 1701859473
transform 1 0 4630 0 1 270
box -12 -8 32 272
use FILL  FILL_0__741_
timestamp 1701859473
transform 1 0 3930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__742_
timestamp 1701859473
transform -1 0 2910 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__743_
timestamp 1701859473
transform 1 0 3050 0 1 270
box -12 -8 32 272
use FILL  FILL_0__744_
timestamp 1701859473
transform -1 0 4430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__745_
timestamp 1701859473
transform 1 0 3650 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__746_
timestamp 1701859473
transform 1 0 2250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__747_
timestamp 1701859473
transform 1 0 3250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__748_
timestamp 1701859473
transform 1 0 3110 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__749_
timestamp 1701859473
transform 1 0 2150 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__750_
timestamp 1701859473
transform -1 0 3230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__751_
timestamp 1701859473
transform 1 0 3350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__752_
timestamp 1701859473
transform 1 0 1630 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__753_
timestamp 1701859473
transform 1 0 3510 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__754_
timestamp 1701859473
transform 1 0 3370 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__755_
timestamp 1701859473
transform -1 0 1410 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__756_
timestamp 1701859473
transform 1 0 2630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__757_
timestamp 1701859473
transform 1 0 2470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__758_
timestamp 1701859473
transform -1 0 2330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__759_
timestamp 1701859473
transform 1 0 2170 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__760_
timestamp 1701859473
transform -1 0 2130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__761_
timestamp 1701859473
transform 1 0 2030 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__762_
timestamp 1701859473
transform -1 0 2130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__763_
timestamp 1701859473
transform -1 0 2250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__764_
timestamp 1701859473
transform 1 0 1990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__765_
timestamp 1701859473
transform -1 0 2130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__766_
timestamp 1701859473
transform 1 0 3350 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__767_
timestamp 1701859473
transform 1 0 2730 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__768_
timestamp 1701859473
transform -1 0 2870 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__769_
timestamp 1701859473
transform -1 0 4170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__770_
timestamp 1701859473
transform -1 0 3530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__771_
timestamp 1701859473
transform -1 0 3650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__772_
timestamp 1701859473
transform -1 0 5390 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__773_
timestamp 1701859473
transform -1 0 4270 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__774_
timestamp 1701859473
transform -1 0 4790 0 1 790
box -12 -8 32 272
use FILL  FILL_0__775_
timestamp 1701859473
transform -1 0 5730 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__776_
timestamp 1701859473
transform 1 0 4890 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__777_
timestamp 1701859473
transform 1 0 5670 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__778_
timestamp 1701859473
transform 1 0 5350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__779_
timestamp 1701859473
transform -1 0 4330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__780_
timestamp 1701859473
transform -1 0 4750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__781_
timestamp 1701859473
transform -1 0 5090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__782_
timestamp 1701859473
transform -1 0 3750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__783_
timestamp 1701859473
transform -1 0 4950 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__784_
timestamp 1701859473
transform 1 0 3810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__785_
timestamp 1701859473
transform -1 0 3410 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__786_
timestamp 1701859473
transform -1 0 3450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__787_
timestamp 1701859473
transform -1 0 4190 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__788_
timestamp 1701859473
transform -1 0 3530 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__789_
timestamp 1701859473
transform -1 0 3810 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__790_
timestamp 1701859473
transform 1 0 1870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__791_
timestamp 1701859473
transform -1 0 2130 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__792_
timestamp 1701859473
transform 1 0 1970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__793_
timestamp 1701859473
transform 1 0 970 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__794_
timestamp 1701859473
transform 1 0 1590 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__795_
timestamp 1701859473
transform -1 0 1330 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__796_
timestamp 1701859473
transform -1 0 510 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__797_
timestamp 1701859473
transform 1 0 1470 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__798_
timestamp 1701859473
transform 1 0 830 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__799_
timestamp 1701859473
transform 1 0 1490 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__800_
timestamp 1701859473
transform 1 0 2250 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__801_
timestamp 1701859473
transform 1 0 1990 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__802_
timestamp 1701859473
transform -1 0 410 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__803_
timestamp 1701859473
transform -1 0 1210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__804_
timestamp 1701859473
transform 1 0 650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__805_
timestamp 1701859473
transform -1 0 970 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__806_
timestamp 1701859473
transform 1 0 2230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__807_
timestamp 1701859473
transform 1 0 1070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__808_
timestamp 1701859473
transform 1 0 970 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__809_
timestamp 1701859473
transform 1 0 1450 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__810_
timestamp 1701859473
transform -1 0 1470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__811_
timestamp 1701859473
transform -1 0 1310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__812_
timestamp 1701859473
transform 1 0 2250 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__813_
timestamp 1701859473
transform 1 0 1630 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__814_
timestamp 1701859473
transform 1 0 3330 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__815_
timestamp 1701859473
transform 1 0 3630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__816_
timestamp 1701859473
transform 1 0 3510 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__817_
timestamp 1701859473
transform 1 0 4430 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__818_
timestamp 1701859473
transform -1 0 4070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__819_
timestamp 1701859473
transform 1 0 3630 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__820_
timestamp 1701859473
transform -1 0 4210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__821_
timestamp 1701859473
transform 1 0 4050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__822_
timestamp 1701859473
transform -1 0 4190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__823_
timestamp 1701859473
transform 1 0 4370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__824_
timestamp 1701859473
transform 1 0 3950 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__825_
timestamp 1701859473
transform -1 0 4090 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__826_
timestamp 1701859473
transform -1 0 4190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__827_
timestamp 1701859473
transform -1 0 3890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__828_
timestamp 1701859473
transform 1 0 4130 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__829_
timestamp 1701859473
transform 1 0 3750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__830_
timestamp 1701859473
transform -1 0 4190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__831_
timestamp 1701859473
transform 1 0 4050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__832_
timestamp 1701859473
transform -1 0 4070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__833_
timestamp 1701859473
transform -1 0 3110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__834_
timestamp 1701859473
transform 1 0 3350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__835_
timestamp 1701859473
transform 1 0 3630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__836_
timestamp 1701859473
transform 1 0 3490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__837_
timestamp 1701859473
transform 1 0 3850 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__838_
timestamp 1701859473
transform 1 0 4630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__839_
timestamp 1701859473
transform -1 0 4950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__840_
timestamp 1701859473
transform 1 0 4490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__841_
timestamp 1701859473
transform 1 0 4770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__842_
timestamp 1701859473
transform -1 0 5090 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__843_
timestamp 1701859473
transform -1 0 4590 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__844_
timestamp 1701859473
transform -1 0 4710 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__845_
timestamp 1701859473
transform -1 0 5690 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__846_
timestamp 1701859473
transform -1 0 3370 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__847_
timestamp 1701859473
transform 1 0 3990 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__848_
timestamp 1701859473
transform 1 0 4310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__849_
timestamp 1701859473
transform 1 0 4490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__850_
timestamp 1701859473
transform -1 0 4230 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__851_
timestamp 1701859473
transform 1 0 4450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__852_
timestamp 1701859473
transform 1 0 4550 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__853_
timestamp 1701859473
transform 1 0 4330 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__854_
timestamp 1701859473
transform 1 0 4250 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__855_
timestamp 1701859473
transform 1 0 4130 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__856_
timestamp 1701859473
transform 1 0 4430 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__857_
timestamp 1701859473
transform 1 0 4570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__858_
timestamp 1701859473
transform -1 0 4590 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__859_
timestamp 1701859473
transform -1 0 4050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__860_
timestamp 1701859473
transform -1 0 4450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__861_
timestamp 1701859473
transform 1 0 3350 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__862_
timestamp 1701859473
transform 1 0 3590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__863_
timestamp 1701859473
transform -1 0 2370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__864_
timestamp 1701859473
transform -1 0 4630 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__865_
timestamp 1701859473
transform 1 0 3850 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__866_
timestamp 1701859473
transform 1 0 3990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__867_
timestamp 1701859473
transform 1 0 4290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__868_
timestamp 1701859473
transform 1 0 4430 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__869_
timestamp 1701859473
transform 1 0 4830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__870_
timestamp 1701859473
transform 1 0 4710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__871_
timestamp 1701859473
transform 1 0 4270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__872_
timestamp 1701859473
transform 1 0 4710 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__873_
timestamp 1701859473
transform 1 0 5030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__874_
timestamp 1701859473
transform 1 0 5170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__875_
timestamp 1701859473
transform 1 0 5010 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__876_
timestamp 1701859473
transform -1 0 5150 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__877_
timestamp 1701859473
transform -1 0 5450 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__878_
timestamp 1701859473
transform 1 0 5310 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__879_
timestamp 1701859473
transform 1 0 4850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__880_
timestamp 1701859473
transform 1 0 4990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__881_
timestamp 1701859473
transform 1 0 4610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__882_
timestamp 1701859473
transform -1 0 4730 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__883_
timestamp 1701859473
transform 1 0 4390 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__884_
timestamp 1701859473
transform -1 0 4350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__885_
timestamp 1701859473
transform -1 0 4530 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__886_
timestamp 1701859473
transform 1 0 4190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__887_
timestamp 1701859473
transform -1 0 5050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__888_
timestamp 1701859473
transform -1 0 4910 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__889_
timestamp 1701859473
transform 1 0 4690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__890_
timestamp 1701859473
transform 1 0 4750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__891_
timestamp 1701859473
transform -1 0 4630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__892_
timestamp 1701859473
transform 1 0 4870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__893_
timestamp 1701859473
transform 1 0 4690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__894_
timestamp 1701859473
transform 1 0 5030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__895_
timestamp 1701859473
transform 1 0 4750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__896_
timestamp 1701859473
transform 1 0 5070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__897_
timestamp 1701859473
transform 1 0 3310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__898_
timestamp 1701859473
transform 1 0 2730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__899_
timestamp 1701859473
transform 1 0 1750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__900_
timestamp 1701859473
transform -1 0 3270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__901_
timestamp 1701859473
transform 1 0 3190 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__902_
timestamp 1701859473
transform -1 0 3450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__903_
timestamp 1701859473
transform -1 0 5170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__904_
timestamp 1701859473
transform 1 0 4930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__905_
timestamp 1701859473
transform 1 0 5010 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__906_
timestamp 1701859473
transform 1 0 5430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__907_
timestamp 1701859473
transform -1 0 5230 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__908_
timestamp 1701859473
transform 1 0 5130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__909_
timestamp 1701859473
transform -1 0 5010 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__910_
timestamp 1701859473
transform 1 0 4850 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__911_
timestamp 1701859473
transform -1 0 5370 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__912_
timestamp 1701859473
transform 1 0 5270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__913_
timestamp 1701859473
transform -1 0 5250 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__914_
timestamp 1701859473
transform 1 0 5430 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__915_
timestamp 1701859473
transform 1 0 5570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__916_
timestamp 1701859473
transform 1 0 5530 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__917_
timestamp 1701859473
transform 1 0 5430 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__918_
timestamp 1701859473
transform -1 0 3590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__919_
timestamp 1701859473
transform 1 0 4750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__920_
timestamp 1701859473
transform 1 0 5670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__921_
timestamp 1701859473
transform 1 0 5490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__922_
timestamp 1701859473
transform 1 0 2570 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__923_
timestamp 1701859473
transform -1 0 3050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__924_
timestamp 1701859473
transform -1 0 2890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__925_
timestamp 1701859473
transform -1 0 2490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__926_
timestamp 1701859473
transform 1 0 2930 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__927_
timestamp 1701859473
transform 1 0 2790 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__928_
timestamp 1701859473
transform 1 0 2690 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__929_
timestamp 1701859473
transform -1 0 3090 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__930_
timestamp 1701859473
transform 1 0 3170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__931_
timestamp 1701859473
transform 1 0 3190 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__932_
timestamp 1701859473
transform -1 0 4510 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__933_
timestamp 1701859473
transform 1 0 4870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__934_
timestamp 1701859473
transform 1 0 5190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__935_
timestamp 1701859473
transform -1 0 4450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__936_
timestamp 1701859473
transform 1 0 5270 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__937_
timestamp 1701859473
transform 1 0 5030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__938_
timestamp 1701859473
transform 1 0 5010 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__939_
timestamp 1701859473
transform -1 0 5430 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__940_
timestamp 1701859473
transform 1 0 5710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__941_
timestamp 1701859473
transform -1 0 4490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__942_
timestamp 1701859473
transform -1 0 4630 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__943_
timestamp 1701859473
transform 1 0 4970 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__944_
timestamp 1701859473
transform -1 0 5310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__945_
timestamp 1701859473
transform 1 0 5290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__946_
timestamp 1701859473
transform 1 0 5430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__947_
timestamp 1701859473
transform 1 0 5570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__948_
timestamp 1701859473
transform -1 0 5590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__949_
timestamp 1701859473
transform -1 0 5410 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__950_
timestamp 1701859473
transform 1 0 4610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__951_
timestamp 1701859473
transform -1 0 5070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__952_
timestamp 1701859473
transform -1 0 5450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__953_
timestamp 1701859473
transform 1 0 5110 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__954_
timestamp 1701859473
transform 1 0 5410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__955_
timestamp 1701859473
transform 1 0 5290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__956_
timestamp 1701859473
transform 1 0 5250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__957_
timestamp 1701859473
transform 1 0 5530 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__958_
timestamp 1701859473
transform -1 0 5590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__959_
timestamp 1701859473
transform 1 0 5570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__960_
timestamp 1701859473
transform 1 0 5270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__961_
timestamp 1701859473
transform -1 0 5610 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__962_
timestamp 1701859473
transform 1 0 5530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__963_
timestamp 1701859473
transform -1 0 5650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__964_
timestamp 1701859473
transform 1 0 5370 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__965_
timestamp 1701859473
transform 1 0 5490 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__966_
timestamp 1701859473
transform 1 0 4650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__967_
timestamp 1701859473
transform -1 0 4530 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__968_
timestamp 1701859473
transform -1 0 4150 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__969_
timestamp 1701859473
transform -1 0 5510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__970_
timestamp 1701859473
transform 1 0 5130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__971_
timestamp 1701859473
transform 1 0 5190 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__972_
timestamp 1701859473
transform -1 0 3150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__973_
timestamp 1701859473
transform 1 0 3370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__974_
timestamp 1701859473
transform 1 0 3810 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__975_
timestamp 1701859473
transform 1 0 4810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__976_
timestamp 1701859473
transform -1 0 4850 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__977_
timestamp 1701859473
transform -1 0 2870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__978_
timestamp 1701859473
transform -1 0 2570 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__979_
timestamp 1701859473
transform -1 0 2730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__980_
timestamp 1701859473
transform 1 0 2290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__981_
timestamp 1701859473
transform 1 0 2430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__982_
timestamp 1701859473
transform -1 0 2590 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__983_
timestamp 1701859473
transform 1 0 2990 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__984_
timestamp 1701859473
transform 1 0 2690 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__985_
timestamp 1701859473
transform 1 0 2990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__986_
timestamp 1701859473
transform 1 0 3090 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__987_
timestamp 1701859473
transform 1 0 3230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__988_
timestamp 1701859473
transform 1 0 5150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__989_
timestamp 1701859473
transform -1 0 5170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__990_
timestamp 1701859473
transform -1 0 2470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__991_
timestamp 1701859473
transform -1 0 3610 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__992_
timestamp 1701859473
transform 1 0 3290 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__993_
timestamp 1701859473
transform 1 0 1650 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__994_
timestamp 1701859473
transform -1 0 3470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__995_
timestamp 1701859473
transform 1 0 3230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__996_
timestamp 1701859473
transform -1 0 3010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__997_
timestamp 1701859473
transform -1 0 2290 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__998_
timestamp 1701859473
transform -1 0 2730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__999_
timestamp 1701859473
transform 1 0 3070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1000_
timestamp 1701859473
transform 1 0 3090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1001_
timestamp 1701859473
transform 1 0 4050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1002_
timestamp 1701859473
transform 1 0 4850 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1003_
timestamp 1701859473
transform 1 0 4730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1004_
timestamp 1701859473
transform -1 0 3530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1005_
timestamp 1701859473
transform 1 0 3370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1006_
timestamp 1701859473
transform 1 0 4330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1007_
timestamp 1701859473
transform -1 0 4470 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1008_
timestamp 1701859473
transform 1 0 3350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1009_
timestamp 1701859473
transform -1 0 3930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1010_
timestamp 1701859473
transform -1 0 4210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1011_
timestamp 1701859473
transform -1 0 4030 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1012_
timestamp 1701859473
transform 1 0 4030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1013_
timestamp 1701859473
transform -1 0 4930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1014_
timestamp 1701859473
transform 1 0 4550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1015_
timestamp 1701859473
transform 1 0 4170 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1016_
timestamp 1701859473
transform -1 0 4330 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1017_
timestamp 1701859473
transform -1 0 4190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1018_
timestamp 1701859473
transform -1 0 4070 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1019_
timestamp 1701859473
transform -1 0 3770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1020_
timestamp 1701859473
transform -1 0 4230 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1021_
timestamp 1701859473
transform -1 0 3530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1022_
timestamp 1701859473
transform -1 0 3750 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1023_
timestamp 1701859473
transform 1 0 3870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1024_
timestamp 1701859473
transform 1 0 3750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1025_
timestamp 1701859473
transform -1 0 3470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1026_
timestamp 1701859473
transform 1 0 5330 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1027_
timestamp 1701859473
transform -1 0 5470 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1028_
timestamp 1701859473
transform 1 0 3650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1029_
timestamp 1701859473
transform -1 0 3930 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1030_
timestamp 1701859473
transform 1 0 3790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1031_
timestamp 1701859473
transform 1 0 3610 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1032_
timestamp 1701859473
transform 1 0 3770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1033_
timestamp 1701859473
transform -1 0 3910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1034_
timestamp 1701859473
transform -1 0 3730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1035_
timestamp 1701859473
transform -1 0 3730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1036_
timestamp 1701859473
transform -1 0 3590 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1037_
timestamp 1701859473
transform 1 0 3230 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1038_
timestamp 1701859473
transform -1 0 2570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1039_
timestamp 1701859473
transform 1 0 3810 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1040_
timestamp 1701859473
transform -1 0 3890 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1041_
timestamp 1701859473
transform -1 0 2170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1042_
timestamp 1701859473
transform -1 0 1650 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1043_
timestamp 1701859473
transform -1 0 1530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1044_
timestamp 1701859473
transform -1 0 2030 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1045_
timestamp 1701859473
transform -1 0 1890 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1046_
timestamp 1701859473
transform 1 0 1770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1047_
timestamp 1701859473
transform -1 0 2050 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1048_
timestamp 1701859473
transform -1 0 1670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1049_
timestamp 1701859473
transform -1 0 2150 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1050_
timestamp 1701859473
transform 1 0 2010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1051_
timestamp 1701859473
transform -1 0 1910 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1052_
timestamp 1701859473
transform 1 0 1850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1053_
timestamp 1701859473
transform 1 0 2830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1054_
timestamp 1701859473
transform -1 0 1410 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1055_
timestamp 1701859473
transform 1 0 1290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1056_
timestamp 1701859473
transform 1 0 1250 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1057_
timestamp 1701859473
transform 1 0 1410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1058_
timestamp 1701859473
transform 1 0 1290 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1059_
timestamp 1701859473
transform 1 0 1190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1060_
timestamp 1701859473
transform 1 0 1570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1061_
timestamp 1701859473
transform 1 0 1170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1062_
timestamp 1701859473
transform -1 0 830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1063_
timestamp 1701859473
transform 1 0 910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1064_
timestamp 1701859473
transform 1 0 1710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1065_
timestamp 1701859473
transform -1 0 3150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1066_
timestamp 1701859473
transform 1 0 2570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1067_
timestamp 1701859473
transform 1 0 1050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1068_
timestamp 1701859473
transform -1 0 1730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1069_
timestamp 1701859473
transform -1 0 2430 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1070_
timestamp 1701859473
transform 1 0 1770 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1071_
timestamp 1701859473
transform 1 0 2010 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1072_
timestamp 1701859473
transform 1 0 2170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1073_
timestamp 1701859473
transform 1 0 1970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1074_
timestamp 1701859473
transform 1 0 1570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1075_
timestamp 1701859473
transform 1 0 1870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1076_
timestamp 1701859473
transform 1 0 2290 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1077_
timestamp 1701859473
transform 1 0 2710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1078_
timestamp 1701859473
transform 1 0 3670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1079_
timestamp 1701859473
transform 1 0 3710 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1080_
timestamp 1701859473
transform 1 0 2150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1081_
timestamp 1701859473
transform 1 0 2310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1082_
timestamp 1701859473
transform -1 0 2870 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1083_
timestamp 1701859473
transform 1 0 2410 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1084_
timestamp 1701859473
transform 1 0 2570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1085_
timestamp 1701859473
transform 1 0 2990 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1086_
timestamp 1701859473
transform 1 0 2790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1087_
timestamp 1701859473
transform 1 0 2830 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1088_
timestamp 1701859473
transform -1 0 3910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1089_
timestamp 1701859473
transform 1 0 3610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1090_
timestamp 1701859473
transform 1 0 2650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1091_
timestamp 1701859473
transform 1 0 2270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1092_
timestamp 1701859473
transform -1 0 2950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1093_
timestamp 1701859473
transform -1 0 2830 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1094_
timestamp 1701859473
transform 1 0 3750 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1095_
timestamp 1701859473
transform 1 0 4230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1096_
timestamp 1701859473
transform 1 0 4090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1097_
timestamp 1701859473
transform 1 0 1730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1098_
timestamp 1701859473
transform 1 0 3070 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1099_
timestamp 1701859473
transform 1 0 2690 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1100_
timestamp 1701859473
transform -1 0 2570 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1101_
timestamp 1701859473
transform -1 0 2450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1102_
timestamp 1701859473
transform -1 0 2130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1103_
timestamp 1701859473
transform 1 0 1770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1104_
timestamp 1701859473
transform -1 0 470 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1105_
timestamp 1701859473
transform -1 0 2070 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1106_
timestamp 1701859473
transform -1 0 1930 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1107_
timestamp 1701859473
transform -1 0 1930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1108_
timestamp 1701859473
transform -1 0 1410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1109_
timestamp 1701859473
transform -1 0 1490 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1110_
timestamp 1701859473
transform -1 0 1250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1111_
timestamp 1701859473
transform -1 0 1110 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1112_
timestamp 1701859473
transform -1 0 770 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1113_
timestamp 1701859473
transform -1 0 690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1114_
timestamp 1701859473
transform 1 0 1350 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1115_
timestamp 1701859473
transform -1 0 1110 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1116_
timestamp 1701859473
transform -1 0 1250 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1117_
timestamp 1701859473
transform -1 0 1090 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1118_
timestamp 1701859473
transform -1 0 950 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1119_
timestamp 1701859473
transform -1 0 570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1120_
timestamp 1701859473
transform -1 0 1130 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1121_
timestamp 1701859473
transform -1 0 1010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1122_
timestamp 1701859473
transform -1 0 1010 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1123_
timestamp 1701859473
transform -1 0 730 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1124_
timestamp 1701859473
transform -1 0 570 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1125_
timestamp 1701859473
transform 1 0 850 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1126_
timestamp 1701859473
transform -1 0 310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1127_
timestamp 1701859473
transform -1 0 590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1128_
timestamp 1701859473
transform -1 0 310 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1129_
timestamp 1701859473
transform 1 0 1430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1130_
timestamp 1701859473
transform -1 0 1530 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1131_
timestamp 1701859473
transform -1 0 450 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1132_
timestamp 1701859473
transform 1 0 10 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1133_
timestamp 1701859473
transform -1 0 430 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1134_
timestamp 1701859473
transform -1 0 170 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0__1135_
timestamp 1701859473
transform 1 0 150 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1136_
timestamp 1701859473
transform 1 0 150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1137_
timestamp 1701859473
transform -1 0 310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1138_
timestamp 1701859473
transform -1 0 30 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1139_
timestamp 1701859473
transform -1 0 30 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1140_
timestamp 1701859473
transform -1 0 170 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1141_
timestamp 1701859473
transform -1 0 310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1142_
timestamp 1701859473
transform 1 0 10 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1143_
timestamp 1701859473
transform -1 0 30 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1144_
timestamp 1701859473
transform 1 0 150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1145_
timestamp 1701859473
transform 1 0 370 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1146_
timestamp 1701859473
transform -1 0 1330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1147_
timestamp 1701859473
transform 1 0 1330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1148_
timestamp 1701859473
transform 1 0 150 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1149_
timestamp 1701859473
transform -1 0 270 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1150_
timestamp 1701859473
transform -1 0 950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1151_
timestamp 1701859473
transform 1 0 650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1152_
timestamp 1701859473
transform -1 0 730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1153_
timestamp 1701859473
transform -1 0 1770 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1154_
timestamp 1701859473
transform 1 0 1490 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1155_
timestamp 1701859473
transform 1 0 1310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1156_
timestamp 1701859473
transform -1 0 1370 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1157_
timestamp 1701859473
transform -1 0 1630 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1158_
timestamp 1701859473
transform -1 0 1230 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1159_
timestamp 1701859473
transform -1 0 1210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1160_
timestamp 1701859473
transform 1 0 1270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1161_
timestamp 1701859473
transform 1 0 1450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1162_
timestamp 1701859473
transform -1 0 1610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1163_
timestamp 1701859473
transform -1 0 990 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1164_
timestamp 1701859473
transform 1 0 830 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1165_
timestamp 1701859473
transform -1 0 830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1166_
timestamp 1701859473
transform -1 0 910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1167_
timestamp 1701859473
transform -1 0 770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1168_
timestamp 1701859473
transform 1 0 570 0 1 4950
box -12 -8 32 272
use FILL  FILL_0__1169_
timestamp 1701859473
transform -1 0 690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1170_
timestamp 1701859473
transform -1 0 590 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1171_
timestamp 1701859473
transform 1 0 530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1172_
timestamp 1701859473
transform -1 0 530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1173_
timestamp 1701859473
transform -1 0 710 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1174_
timestamp 1701859473
transform 1 0 390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0__1175_
timestamp 1701859473
transform -1 0 450 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1176_
timestamp 1701859473
transform -1 0 190 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1177_
timestamp 1701859473
transform 1 0 10 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1178_
timestamp 1701859473
transform -1 0 450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1179_
timestamp 1701859473
transform -1 0 330 0 1 4430
box -12 -8 32 272
use FILL  FILL_0__1180_
timestamp 1701859473
transform -1 0 310 0 1 3910
box -12 -8 32 272
use FILL  FILL_0__1181_
timestamp 1701859473
transform -1 0 30 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1182_
timestamp 1701859473
transform -1 0 30 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1183_
timestamp 1701859473
transform -1 0 290 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1184_
timestamp 1701859473
transform 1 0 130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1185_
timestamp 1701859473
transform 1 0 10 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1186_
timestamp 1701859473
transform -1 0 270 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1187_
timestamp 1701859473
transform 1 0 290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1188_
timestamp 1701859473
transform 1 0 10 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1189_
timestamp 1701859473
transform -1 0 150 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1190_
timestamp 1701859473
transform 1 0 190 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1191_
timestamp 1701859473
transform 1 0 270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1192_
timestamp 1701859473
transform -1 0 410 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1193_
timestamp 1701859473
transform -1 0 1050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1194_
timestamp 1701859473
transform -1 0 1230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1195_
timestamp 1701859473
transform -1 0 870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0__1196_
timestamp 1701859473
transform -1 0 1750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1197_
timestamp 1701859473
transform -1 0 1670 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1198_
timestamp 1701859473
transform -1 0 1550 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1199_
timestamp 1701859473
transform 1 0 1390 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1200_
timestamp 1701859473
transform -1 0 1090 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1201_
timestamp 1701859473
transform 1 0 930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1202_
timestamp 1701859473
transform 1 0 790 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1203_
timestamp 1701859473
transform 1 0 970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1204_
timestamp 1701859473
transform 1 0 1070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1205_
timestamp 1701859473
transform -1 0 870 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1206_
timestamp 1701859473
transform -1 0 850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1207_
timestamp 1701859473
transform -1 0 710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1208_
timestamp 1701859473
transform 1 0 550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1209_
timestamp 1701859473
transform -1 0 430 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1210_
timestamp 1701859473
transform 1 0 150 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1211_
timestamp 1701859473
transform 1 0 370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1212_
timestamp 1701859473
transform 1 0 2930 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1213_
timestamp 1701859473
transform -1 0 3490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1214_
timestamp 1701859473
transform 1 0 490 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1215_
timestamp 1701859473
transform -1 0 650 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1216_
timestamp 1701859473
transform -1 0 150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1217_
timestamp 1701859473
transform -1 0 250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1218_
timestamp 1701859473
transform -1 0 270 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1219_
timestamp 1701859473
transform 1 0 130 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1220_
timestamp 1701859473
transform 1 0 250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1221_
timestamp 1701859473
transform -1 0 970 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1222_
timestamp 1701859473
transform 1 0 1490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1223_
timestamp 1701859473
transform 1 0 1310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1224_
timestamp 1701859473
transform -1 0 1610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1225_
timestamp 1701859473
transform -1 0 1870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1226_
timestamp 1701859473
transform -1 0 1910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1227_
timestamp 1701859473
transform -1 0 1630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1228_
timestamp 1701859473
transform -1 0 1510 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1229_
timestamp 1701859473
transform 1 0 1090 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1230_
timestamp 1701859473
transform -1 0 670 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1231_
timestamp 1701859473
transform 1 0 10 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1232_
timestamp 1701859473
transform -1 0 130 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1233_
timestamp 1701859473
transform -1 0 30 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1234_
timestamp 1701859473
transform 1 0 10 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1235_
timestamp 1701859473
transform -1 0 30 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1236_
timestamp 1701859473
transform -1 0 30 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1237_
timestamp 1701859473
transform -1 0 170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1238_
timestamp 1701859473
transform -1 0 1190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1239_
timestamp 1701859473
transform 1 0 910 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1240_
timestamp 1701859473
transform -1 0 1070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1241_
timestamp 1701859473
transform 1 0 410 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1242_
timestamp 1701859473
transform 1 0 770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1243_
timestamp 1701859473
transform 1 0 1270 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1244_
timestamp 1701859473
transform 1 0 1730 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1245_
timestamp 1701859473
transform 1 0 1750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1246_
timestamp 1701859473
transform -1 0 1510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1247_
timestamp 1701859473
transform 1 0 1190 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1248_
timestamp 1701859473
transform -1 0 1070 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1249_
timestamp 1701859473
transform 1 0 650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1250_
timestamp 1701859473
transform -1 0 570 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1251_
timestamp 1701859473
transform 1 0 630 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1252_
timestamp 1701859473
transform 1 0 490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1253_
timestamp 1701859473
transform -1 0 550 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1254_
timestamp 1701859473
transform -1 0 410 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1255_
timestamp 1701859473
transform 1 0 490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1256_
timestamp 1701859473
transform 1 0 730 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1257_
timestamp 1701859473
transform 1 0 770 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1258_
timestamp 1701859473
transform -1 0 930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1259_
timestamp 1701859473
transform -1 0 810 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1260_
timestamp 1701859473
transform 1 0 3390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1261_
timestamp 1701859473
transform -1 0 3390 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1262_
timestamp 1701859473
transform 1 0 3270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1263_
timestamp 1701859473
transform 1 0 3250 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1264_
timestamp 1701859473
transform -1 0 3170 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1265_
timestamp 1701859473
transform 1 0 3270 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1266_
timestamp 1701859473
transform 1 0 4250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1267_
timestamp 1701859473
transform 1 0 3990 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1268_
timestamp 1701859473
transform 1 0 4010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1269_
timestamp 1701859473
transform 1 0 3610 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1270_
timestamp 1701859473
transform 1 0 3490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1271_
timestamp 1701859473
transform -1 0 3750 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1272_
timestamp 1701859473
transform 1 0 3870 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1273_
timestamp 1701859473
transform -1 0 4310 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1274_
timestamp 1701859473
transform 1 0 4250 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1275_
timestamp 1701859473
transform -1 0 4130 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1276_
timestamp 1701859473
transform -1 0 5190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1277_
timestamp 1701859473
transform 1 0 5170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1278_
timestamp 1701859473
transform 1 0 5670 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1279_
timestamp 1701859473
transform 1 0 5650 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1280_
timestamp 1701859473
transform -1 0 4930 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1281_
timestamp 1701859473
transform 1 0 5030 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1282_
timestamp 1701859473
transform -1 0 5710 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1283_
timestamp 1701859473
transform -1 0 5610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1284_
timestamp 1701859473
transform -1 0 5710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1285_
timestamp 1701859473
transform 1 0 5490 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1286_
timestamp 1701859473
transform 1 0 5310 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1287_
timestamp 1701859473
transform -1 0 5530 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1288_
timestamp 1701859473
transform 1 0 4050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1289_
timestamp 1701859473
transform 1 0 5190 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1290_
timestamp 1701859473
transform 1 0 5310 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1291_
timestamp 1701859473
transform -1 0 5050 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1292_
timestamp 1701859473
transform 1 0 4910 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1293_
timestamp 1701859473
transform -1 0 5650 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1294_
timestamp 1701859473
transform -1 0 5510 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1295_
timestamp 1701859473
transform -1 0 5150 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1296_
timestamp 1701859473
transform 1 0 5010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1297_
timestamp 1701859473
transform 1 0 5230 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1298_
timestamp 1701859473
transform -1 0 5010 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1299_
timestamp 1701859473
transform -1 0 4190 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1300_
timestamp 1701859473
transform 1 0 5150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1301_
timestamp 1701859473
transform 1 0 5350 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1302_
timestamp 1701859473
transform 1 0 5290 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1303_
timestamp 1701859473
transform 1 0 5170 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1304_
timestamp 1701859473
transform -1 0 5190 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1305_
timestamp 1701859473
transform 1 0 5450 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1306_
timestamp 1701859473
transform 1 0 5570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1307_
timestamp 1701859473
transform -1 0 5130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1308_
timestamp 1701859473
transform 1 0 5210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1309_
timestamp 1701859473
transform -1 0 5370 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1310_
timestamp 1701859473
transform -1 0 4470 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1311_
timestamp 1701859473
transform -1 0 4870 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1312_
timestamp 1701859473
transform 1 0 4230 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1313_
timestamp 1701859473
transform 1 0 4730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1314_
timestamp 1701859473
transform 1 0 4590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1315_
timestamp 1701859473
transform -1 0 4670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1316_
timestamp 1701859473
transform -1 0 4530 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1317_
timestamp 1701859473
transform 1 0 3910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1318_
timestamp 1701859473
transform 1 0 4350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1319_
timestamp 1701859473
transform -1 0 4490 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1320_
timestamp 1701859473
transform 1 0 4590 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1321_
timestamp 1701859473
transform 1 0 4670 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1322_
timestamp 1701859473
transform 1 0 3950 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1323_
timestamp 1701859473
transform 1 0 4710 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1324_
timestamp 1701859473
transform 1 0 4570 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1325_
timestamp 1701859473
transform 1 0 2150 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1326_
timestamp 1701859473
transform -1 0 4910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1327_
timestamp 1701859473
transform -1 0 4430 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1328_
timestamp 1701859473
transform 1 0 4530 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1329_
timestamp 1701859473
transform 1 0 4370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1330_
timestamp 1701859473
transform -1 0 4610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1331_
timestamp 1701859473
transform -1 0 4810 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1332_
timestamp 1701859473
transform -1 0 4670 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1333_
timestamp 1701859473
transform 1 0 4530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1334_
timestamp 1701859473
transform -1 0 1630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1335_
timestamp 1701859473
transform -1 0 1770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1336_
timestamp 1701859473
transform 1 0 1590 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1337_
timestamp 1701859473
transform 1 0 1910 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1338_
timestamp 1701859473
transform 1 0 1850 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1339_
timestamp 1701859473
transform -1 0 1830 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1340_
timestamp 1701859473
transform -1 0 1730 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1341_
timestamp 1701859473
transform 1 0 2010 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1342_
timestamp 1701859473
transform -1 0 1590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1343_
timestamp 1701859473
transform -1 0 990 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1344_
timestamp 1701859473
transform -1 0 850 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1345_
timestamp 1701859473
transform 1 0 1090 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1346_
timestamp 1701859473
transform -1 0 1210 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1347_
timestamp 1701859473
transform 1 0 1250 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1348_
timestamp 1701859473
transform 1 0 1630 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1349_
timestamp 1701859473
transform -1 0 2430 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1350_
timestamp 1701859473
transform 1 0 2030 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1351_
timestamp 1701859473
transform -1 0 2670 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1352_
timestamp 1701859473
transform 1 0 1490 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1353_
timestamp 1701859473
transform -1 0 1330 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1354_
timestamp 1701859473
transform -1 0 1370 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1355_
timestamp 1701859473
transform -1 0 270 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1356_
timestamp 1701859473
transform -1 0 390 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1357_
timestamp 1701859473
transform 1 0 270 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1358_
timestamp 1701859473
transform 1 0 390 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1359_
timestamp 1701859473
transform 1 0 1850 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1360_
timestamp 1701859473
transform -1 0 1730 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1361_
timestamp 1701859473
transform 1 0 2270 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1362_
timestamp 1701859473
transform -1 0 1230 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1363_
timestamp 1701859473
transform 1 0 1090 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1364_
timestamp 1701859473
transform -1 0 750 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1365_
timestamp 1701859473
transform -1 0 630 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1366_
timestamp 1701859473
transform 1 0 610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1367_
timestamp 1701859473
transform -1 0 650 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1368_
timestamp 1701859473
transform -1 0 930 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1369_
timestamp 1701859473
transform -1 0 1490 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1370_
timestamp 1701859473
transform 1 0 1330 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1371_
timestamp 1701859473
transform 1 0 510 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1372_
timestamp 1701859473
transform -1 0 790 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1373_
timestamp 1701859473
transform -1 0 510 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1374_
timestamp 1701859473
transform 1 0 610 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1375_
timestamp 1701859473
transform -1 0 170 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1376_
timestamp 1701859473
transform 1 0 370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1377_
timestamp 1701859473
transform -1 0 290 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1378_
timestamp 1701859473
transform -1 0 30 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1379_
timestamp 1701859473
transform 1 0 10 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1380_
timestamp 1701859473
transform 1 0 10 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1381_
timestamp 1701859473
transform 1 0 10 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1382_
timestamp 1701859473
transform 1 0 110 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1383_
timestamp 1701859473
transform 1 0 130 0 -1 790
box -12 -8 32 272
use FILL  FILL_0__1384_
timestamp 1701859473
transform 1 0 110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1385_
timestamp 1701859473
transform -1 0 850 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1386_
timestamp 1701859473
transform -1 0 870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1387_
timestamp 1701859473
transform -1 0 750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1388_
timestamp 1701859473
transform -1 0 530 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1389_
timestamp 1701859473
transform 1 0 270 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1390_
timestamp 1701859473
transform 1 0 430 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1391_
timestamp 1701859473
transform -1 0 590 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1392_
timestamp 1701859473
transform -1 0 390 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1393_
timestamp 1701859473
transform 1 0 370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1394_
timestamp 1701859473
transform -1 0 270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1395_
timestamp 1701859473
transform 1 0 470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1396_
timestamp 1701859473
transform 1 0 850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1397_
timestamp 1701859473
transform -1 0 970 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1398_
timestamp 1701859473
transform -1 0 1230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1399_
timestamp 1701859473
transform -1 0 1070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1400_
timestamp 1701859473
transform -1 0 1530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1401_
timestamp 1701859473
transform 1 0 1090 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1402_
timestamp 1701859473
transform 1 0 1230 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1403_
timestamp 1701859473
transform 1 0 1370 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1404_
timestamp 1701859473
transform 1 0 1350 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1405_
timestamp 1701859473
transform -1 0 3170 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1406_
timestamp 1701859473
transform 1 0 2430 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1407_
timestamp 1701859473
transform 1 0 2090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1408_
timestamp 1701859473
transform -1 0 2230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1409_
timestamp 1701859473
transform 1 0 3430 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1410_
timestamp 1701859473
transform 1 0 2390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1411_
timestamp 1701859473
transform -1 0 2530 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1412_
timestamp 1701859473
transform -1 0 3550 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1413_
timestamp 1701859473
transform 1 0 2050 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1414_
timestamp 1701859473
transform -1 0 2190 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1415_
timestamp 1701859473
transform -1 0 3710 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1416_
timestamp 1701859473
transform 1 0 2350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1417_
timestamp 1701859473
transform -1 0 2570 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1418_
timestamp 1701859473
transform 1 0 3190 0 1 270
box -12 -8 32 272
use FILL  FILL_0__1419_
timestamp 1701859473
transform 1 0 2110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1420_
timestamp 1701859473
transform -1 0 2250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1421_
timestamp 1701859473
transform 1 0 2190 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1422_
timestamp 1701859473
transform -1 0 2570 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1423_
timestamp 1701859473
transform -1 0 2710 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1424_
timestamp 1701859473
transform -1 0 3070 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1425_
timestamp 1701859473
transform 1 0 2370 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1426_
timestamp 1701859473
transform -1 0 2750 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1427_
timestamp 1701859473
transform 1 0 2710 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1428_
timestamp 1701859473
transform 1 0 3110 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1429_
timestamp 1701859473
transform 1 0 3250 0 1 1830
box -12 -8 32 272
use FILL  FILL_0__1430_
timestamp 1701859473
transform 1 0 3230 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1431_
timestamp 1701859473
transform -1 0 3370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1432_
timestamp 1701859473
transform -1 0 3230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1433_
timestamp 1701859473
transform 1 0 3070 0 -1 2350
box -12 -8 32 272
use FILL  FILL_0__1434_
timestamp 1701859473
transform -1 0 3110 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1435_
timestamp 1701859473
transform 1 0 2930 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1436_
timestamp 1701859473
transform 1 0 2730 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1437_
timestamp 1701859473
transform -1 0 2610 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0__1438_
timestamp 1701859473
transform 1 0 2910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1439_
timestamp 1701859473
transform 1 0 2770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_0__1440_
timestamp 1701859473
transform -1 0 3850 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1441_
timestamp 1701859473
transform 1 0 3450 0 1 1310
box -12 -8 32 272
use FILL  FILL_0__1442_
timestamp 1701859473
transform 1 0 3490 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0__1443_
timestamp 1701859473
transform -1 0 3390 0 1 2350
box -12 -8 32 272
use FILL  FILL_0__1444_
timestamp 1701859473
transform -1 0 2450 0 1 3390
box -12 -8 32 272
use FILL  FILL_0__1445_
timestamp 1701859473
transform -1 0 2610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1446_
timestamp 1701859473
transform -1 0 2850 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1447_
timestamp 1701859473
transform -1 0 2970 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1448_
timestamp 1701859473
transform -1 0 2390 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1449_
timestamp 1701859473
transform -1 0 2750 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1450_
timestamp 1701859473
transform -1 0 1990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1451_
timestamp 1701859473
transform 1 0 1850 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1527_
timestamp 1701859473
transform 1 0 5670 0 1 790
box -12 -8 32 272
use FILL  FILL_0__1528_
timestamp 1701859473
transform -1 0 5690 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1529_
timestamp 1701859473
transform 1 0 5370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0__1530_
timestamp 1701859473
transform 1 0 5110 0 1 2870
box -12 -8 32 272
use FILL  FILL_0__1531_
timestamp 1701859473
transform 1 0 2750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_0__1532_
timestamp 1701859473
transform 1 0 3790 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1533_
timestamp 1701859473
transform 1 0 4050 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1534_
timestamp 1701859473
transform 1 0 4170 0 -1 270
box -12 -8 32 272
use FILL  FILL_0__1535_
timestamp 1701859473
transform 1 0 3930 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert0
timestamp 1701859473
transform -1 0 1470 0 1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert1
timestamp 1701859473
transform 1 0 2130 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert2
timestamp 1701859473
transform 1 0 4770 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert3
timestamp 1701859473
transform 1 0 3650 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert4
timestamp 1701859473
transform 1 0 2130 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert5
timestamp 1701859473
transform 1 0 4130 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert6
timestamp 1701859473
transform -1 0 1350 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert15
timestamp 1701859473
transform -1 0 4730 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert16
timestamp 1701859473
transform -1 0 3510 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert17
timestamp 1701859473
transform -1 0 3950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert18
timestamp 1701859473
transform 1 0 4890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert19
timestamp 1701859473
transform -1 0 1610 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert20
timestamp 1701859473
transform -1 0 4350 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert21
timestamp 1701859473
transform -1 0 1790 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert22
timestamp 1701859473
transform -1 0 4830 0 1 1830
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert23
timestamp 1701859473
transform -1 0 3050 0 -1 790
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert24
timestamp 1701859473
transform 1 0 5030 0 1 270
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert25
timestamp 1701859473
transform -1 0 3010 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert26
timestamp 1701859473
transform 1 0 2990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert27
timestamp 1701859473
transform 1 0 3130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert28
timestamp 1701859473
transform 1 0 2610 0 1 1310
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert29
timestamp 1701859473
transform -1 0 2490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert30
timestamp 1701859473
transform -1 0 4330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert31
timestamp 1701859473
transform -1 0 3470 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert32
timestamp 1701859473
transform 1 0 4590 0 1 4950
box -12 -8 32 272
use FILL  FILL_0_BUFX2_insert33
timestamp 1701859473
transform -1 0 4370 0 1 4430
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 2770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert8
timestamp 1701859473
transform -1 0 1590 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 1730 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert10
timestamp 1701859473
transform -1 0 2330 0 1 2350
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert11
timestamp 1701859473
transform 1 0 4250 0 1 790
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert12
timestamp 1701859473
transform -1 0 3210 0 -1 270
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert13
timestamp 1701859473
transform 1 0 2850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_0_CLKBUF1_insert14
timestamp 1701859473
transform 1 0 4930 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__723_
timestamp 1701859473
transform -1 0 2810 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__724_
timestamp 1701859473
transform -1 0 2610 0 1 790
box -12 -8 32 272
use FILL  FILL_1__725_
timestamp 1701859473
transform -1 0 2690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__726_
timestamp 1701859473
transform 1 0 3330 0 1 270
box -12 -8 32 272
use FILL  FILL_1__727_
timestamp 1701859473
transform 1 0 2890 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__728_
timestamp 1701859473
transform -1 0 3030 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__729_
timestamp 1701859473
transform 1 0 3670 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__730_
timestamp 1701859473
transform 1 0 3570 0 1 270
box -12 -8 32 272
use FILL  FILL_1__731_
timestamp 1701859473
transform -1 0 3490 0 1 270
box -12 -8 32 272
use FILL  FILL_1__732_
timestamp 1701859473
transform -1 0 770 0 1 790
box -12 -8 32 272
use FILL  FILL_1__733_
timestamp 1701859473
transform -1 0 1990 0 1 790
box -12 -8 32 272
use FILL  FILL_1__734_
timestamp 1701859473
transform -1 0 2950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__735_
timestamp 1701859473
transform 1 0 4090 0 1 270
box -12 -8 32 272
use FILL  FILL_1__736_
timestamp 1701859473
transform 1 0 3810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__737_
timestamp 1701859473
transform 1 0 970 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__738_
timestamp 1701859473
transform -1 0 2110 0 1 790
box -12 -8 32 272
use FILL  FILL_1__739_
timestamp 1701859473
transform -1 0 2810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__740_
timestamp 1701859473
transform 1 0 4650 0 1 270
box -12 -8 32 272
use FILL  FILL_1__741_
timestamp 1701859473
transform 1 0 3950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__742_
timestamp 1701859473
transform -1 0 2930 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__743_
timestamp 1701859473
transform 1 0 3070 0 1 270
box -12 -8 32 272
use FILL  FILL_1__744_
timestamp 1701859473
transform -1 0 4450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__745_
timestamp 1701859473
transform 1 0 3670 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__746_
timestamp 1701859473
transform 1 0 2270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__747_
timestamp 1701859473
transform 1 0 3270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__748_
timestamp 1701859473
transform 1 0 3130 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__749_
timestamp 1701859473
transform 1 0 2170 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__750_
timestamp 1701859473
transform -1 0 3250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__751_
timestamp 1701859473
transform 1 0 3370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__752_
timestamp 1701859473
transform 1 0 1650 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__753_
timestamp 1701859473
transform 1 0 3530 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__754_
timestamp 1701859473
transform 1 0 3390 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__755_
timestamp 1701859473
transform -1 0 1430 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__756_
timestamp 1701859473
transform 1 0 2650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__757_
timestamp 1701859473
transform 1 0 2490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__758_
timestamp 1701859473
transform -1 0 2350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__759_
timestamp 1701859473
transform 1 0 2190 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__760_
timestamp 1701859473
transform -1 0 2150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__761_
timestamp 1701859473
transform 1 0 2050 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__762_
timestamp 1701859473
transform -1 0 2150 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__763_
timestamp 1701859473
transform -1 0 2270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__764_
timestamp 1701859473
transform 1 0 2010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__765_
timestamp 1701859473
transform -1 0 2150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__766_
timestamp 1701859473
transform 1 0 3370 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__767_
timestamp 1701859473
transform 1 0 2750 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__768_
timestamp 1701859473
transform -1 0 2890 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__769_
timestamp 1701859473
transform -1 0 4190 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__770_
timestamp 1701859473
transform -1 0 3550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__771_
timestamp 1701859473
transform -1 0 3670 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__772_
timestamp 1701859473
transform -1 0 5410 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__773_
timestamp 1701859473
transform -1 0 4290 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__774_
timestamp 1701859473
transform -1 0 4810 0 1 790
box -12 -8 32 272
use FILL  FILL_1__775_
timestamp 1701859473
transform -1 0 5750 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__776_
timestamp 1701859473
transform 1 0 4910 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__777_
timestamp 1701859473
transform 1 0 5690 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__778_
timestamp 1701859473
transform 1 0 5370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__779_
timestamp 1701859473
transform -1 0 4350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__780_
timestamp 1701859473
transform -1 0 4770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__781_
timestamp 1701859473
transform -1 0 5110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__782_
timestamp 1701859473
transform -1 0 3770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__783_
timestamp 1701859473
transform -1 0 4970 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__784_
timestamp 1701859473
transform 1 0 3830 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__785_
timestamp 1701859473
transform -1 0 3430 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__786_
timestamp 1701859473
transform -1 0 3470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__787_
timestamp 1701859473
transform -1 0 4210 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__788_
timestamp 1701859473
transform -1 0 3550 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__789_
timestamp 1701859473
transform -1 0 3830 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__790_
timestamp 1701859473
transform 1 0 1890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__791_
timestamp 1701859473
transform -1 0 2150 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__792_
timestamp 1701859473
transform 1 0 1990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__793_
timestamp 1701859473
transform 1 0 990 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__794_
timestamp 1701859473
transform 1 0 1610 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__795_
timestamp 1701859473
transform -1 0 1350 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__796_
timestamp 1701859473
transform -1 0 530 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__797_
timestamp 1701859473
transform 1 0 1490 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__798_
timestamp 1701859473
transform 1 0 850 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__799_
timestamp 1701859473
transform 1 0 1510 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__800_
timestamp 1701859473
transform 1 0 2270 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__801_
timestamp 1701859473
transform 1 0 2010 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__802_
timestamp 1701859473
transform -1 0 430 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__803_
timestamp 1701859473
transform -1 0 1230 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__804_
timestamp 1701859473
transform 1 0 670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__805_
timestamp 1701859473
transform -1 0 990 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__806_
timestamp 1701859473
transform 1 0 2250 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__807_
timestamp 1701859473
transform 1 0 1090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__808_
timestamp 1701859473
transform 1 0 990 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__809_
timestamp 1701859473
transform 1 0 1470 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__810_
timestamp 1701859473
transform -1 0 1490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__811_
timestamp 1701859473
transform -1 0 1330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__812_
timestamp 1701859473
transform 1 0 2270 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__813_
timestamp 1701859473
transform 1 0 1650 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__814_
timestamp 1701859473
transform 1 0 3350 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__815_
timestamp 1701859473
transform 1 0 3650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__816_
timestamp 1701859473
transform 1 0 3530 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__817_
timestamp 1701859473
transform 1 0 4450 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__818_
timestamp 1701859473
transform -1 0 4090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__819_
timestamp 1701859473
transform 1 0 3650 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__820_
timestamp 1701859473
transform -1 0 4230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__821_
timestamp 1701859473
transform 1 0 4070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__822_
timestamp 1701859473
transform -1 0 4210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__823_
timestamp 1701859473
transform 1 0 4390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__824_
timestamp 1701859473
transform 1 0 3970 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__825_
timestamp 1701859473
transform -1 0 4110 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__826_
timestamp 1701859473
transform -1 0 4210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__827_
timestamp 1701859473
transform -1 0 3910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__828_
timestamp 1701859473
transform 1 0 4150 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__829_
timestamp 1701859473
transform 1 0 3770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__830_
timestamp 1701859473
transform -1 0 4210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__831_
timestamp 1701859473
transform 1 0 4070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__832_
timestamp 1701859473
transform -1 0 4090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__833_
timestamp 1701859473
transform -1 0 3130 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__834_
timestamp 1701859473
transform 1 0 3370 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__835_
timestamp 1701859473
transform 1 0 3650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__836_
timestamp 1701859473
transform 1 0 3510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__837_
timestamp 1701859473
transform 1 0 3870 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__838_
timestamp 1701859473
transform 1 0 4650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__839_
timestamp 1701859473
transform -1 0 4970 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__840_
timestamp 1701859473
transform 1 0 4510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__841_
timestamp 1701859473
transform 1 0 4790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__842_
timestamp 1701859473
transform -1 0 5110 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__843_
timestamp 1701859473
transform -1 0 4610 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__844_
timestamp 1701859473
transform -1 0 4730 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__845_
timestamp 1701859473
transform -1 0 5710 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__846_
timestamp 1701859473
transform -1 0 3390 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__847_
timestamp 1701859473
transform 1 0 4010 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__848_
timestamp 1701859473
transform 1 0 4330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__849_
timestamp 1701859473
transform 1 0 4510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__850_
timestamp 1701859473
transform -1 0 4250 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__851_
timestamp 1701859473
transform 1 0 4470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__852_
timestamp 1701859473
transform 1 0 4570 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__853_
timestamp 1701859473
transform 1 0 4350 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__854_
timestamp 1701859473
transform 1 0 4270 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__855_
timestamp 1701859473
transform 1 0 4150 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__856_
timestamp 1701859473
transform 1 0 4450 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__857_
timestamp 1701859473
transform 1 0 4590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__858_
timestamp 1701859473
transform -1 0 4610 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__859_
timestamp 1701859473
transform -1 0 4070 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__860_
timestamp 1701859473
transform -1 0 4470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__861_
timestamp 1701859473
transform 1 0 3370 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__862_
timestamp 1701859473
transform 1 0 3610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__863_
timestamp 1701859473
transform -1 0 2390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__864_
timestamp 1701859473
transform -1 0 4650 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__865_
timestamp 1701859473
transform 1 0 3870 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__866_
timestamp 1701859473
transform 1 0 4010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__867_
timestamp 1701859473
transform 1 0 4310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__868_
timestamp 1701859473
transform 1 0 4450 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__869_
timestamp 1701859473
transform 1 0 4850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__870_
timestamp 1701859473
transform 1 0 4730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__871_
timestamp 1701859473
transform 1 0 4290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__872_
timestamp 1701859473
transform 1 0 4730 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__873_
timestamp 1701859473
transform 1 0 5050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__874_
timestamp 1701859473
transform 1 0 5190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__875_
timestamp 1701859473
transform 1 0 5030 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__876_
timestamp 1701859473
transform -1 0 5170 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__877_
timestamp 1701859473
transform -1 0 5470 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__878_
timestamp 1701859473
transform 1 0 5330 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__879_
timestamp 1701859473
transform 1 0 4870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__880_
timestamp 1701859473
transform 1 0 5010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__881_
timestamp 1701859473
transform 1 0 4630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__882_
timestamp 1701859473
transform -1 0 4750 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__883_
timestamp 1701859473
transform 1 0 4410 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__884_
timestamp 1701859473
transform -1 0 4370 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__885_
timestamp 1701859473
transform -1 0 4550 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__886_
timestamp 1701859473
transform 1 0 4210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__887_
timestamp 1701859473
transform -1 0 5070 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__888_
timestamp 1701859473
transform -1 0 4930 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__889_
timestamp 1701859473
transform 1 0 4710 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__890_
timestamp 1701859473
transform 1 0 4770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__891_
timestamp 1701859473
transform -1 0 4650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__892_
timestamp 1701859473
transform 1 0 4890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__893_
timestamp 1701859473
transform 1 0 4710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__894_
timestamp 1701859473
transform 1 0 5050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__895_
timestamp 1701859473
transform 1 0 4770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__896_
timestamp 1701859473
transform 1 0 5090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__897_
timestamp 1701859473
transform 1 0 3330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__898_
timestamp 1701859473
transform 1 0 2750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__899_
timestamp 1701859473
transform 1 0 1770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__900_
timestamp 1701859473
transform -1 0 3290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__901_
timestamp 1701859473
transform 1 0 3210 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__902_
timestamp 1701859473
transform -1 0 3470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__903_
timestamp 1701859473
transform -1 0 5190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__904_
timestamp 1701859473
transform 1 0 4950 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__905_
timestamp 1701859473
transform 1 0 5030 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__906_
timestamp 1701859473
transform 1 0 5450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__907_
timestamp 1701859473
transform -1 0 5250 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__908_
timestamp 1701859473
transform 1 0 5150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__909_
timestamp 1701859473
transform -1 0 5030 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__910_
timestamp 1701859473
transform 1 0 4870 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__911_
timestamp 1701859473
transform -1 0 5390 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__912_
timestamp 1701859473
transform 1 0 5290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__913_
timestamp 1701859473
transform -1 0 5270 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__914_
timestamp 1701859473
transform 1 0 5450 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__915_
timestamp 1701859473
transform 1 0 5590 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__916_
timestamp 1701859473
transform 1 0 5550 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__917_
timestamp 1701859473
transform 1 0 5450 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__918_
timestamp 1701859473
transform -1 0 3610 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__919_
timestamp 1701859473
transform 1 0 4770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__920_
timestamp 1701859473
transform 1 0 5690 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__921_
timestamp 1701859473
transform 1 0 5510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__922_
timestamp 1701859473
transform 1 0 2590 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__923_
timestamp 1701859473
transform -1 0 3070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__924_
timestamp 1701859473
transform -1 0 2910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__925_
timestamp 1701859473
transform -1 0 2510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__926_
timestamp 1701859473
transform 1 0 2950 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__927_
timestamp 1701859473
transform 1 0 2810 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__928_
timestamp 1701859473
transform 1 0 2710 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__929_
timestamp 1701859473
transform -1 0 3110 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__930_
timestamp 1701859473
transform 1 0 3190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__931_
timestamp 1701859473
transform 1 0 3210 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__932_
timestamp 1701859473
transform -1 0 4530 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__933_
timestamp 1701859473
transform 1 0 4890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__934_
timestamp 1701859473
transform 1 0 5210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__935_
timestamp 1701859473
transform -1 0 4470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__936_
timestamp 1701859473
transform 1 0 5290 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__937_
timestamp 1701859473
transform 1 0 5050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__938_
timestamp 1701859473
transform 1 0 5030 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__939_
timestamp 1701859473
transform -1 0 5450 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__940_
timestamp 1701859473
transform 1 0 5730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__941_
timestamp 1701859473
transform -1 0 4510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__942_
timestamp 1701859473
transform -1 0 4650 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__943_
timestamp 1701859473
transform 1 0 4990 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__944_
timestamp 1701859473
transform -1 0 5330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__945_
timestamp 1701859473
transform 1 0 5310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__946_
timestamp 1701859473
transform 1 0 5450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__947_
timestamp 1701859473
transform 1 0 5590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__948_
timestamp 1701859473
transform -1 0 5610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__949_
timestamp 1701859473
transform -1 0 5430 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__950_
timestamp 1701859473
transform 1 0 4630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__951_
timestamp 1701859473
transform -1 0 5090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__952_
timestamp 1701859473
transform -1 0 5470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__953_
timestamp 1701859473
transform 1 0 5130 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__954_
timestamp 1701859473
transform 1 0 5430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__955_
timestamp 1701859473
transform 1 0 5310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__956_
timestamp 1701859473
transform 1 0 5270 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__957_
timestamp 1701859473
transform 1 0 5550 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__958_
timestamp 1701859473
transform -1 0 5610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__959_
timestamp 1701859473
transform 1 0 5590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__960_
timestamp 1701859473
transform 1 0 5290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__961_
timestamp 1701859473
transform -1 0 5630 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__962_
timestamp 1701859473
transform 1 0 5550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__963_
timestamp 1701859473
transform -1 0 5670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__964_
timestamp 1701859473
transform 1 0 5390 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__965_
timestamp 1701859473
transform 1 0 5510 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__966_
timestamp 1701859473
transform 1 0 4670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__967_
timestamp 1701859473
transform -1 0 4550 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__968_
timestamp 1701859473
transform -1 0 4170 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__969_
timestamp 1701859473
transform -1 0 5530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__970_
timestamp 1701859473
transform 1 0 5150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__971_
timestamp 1701859473
transform 1 0 5210 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__972_
timestamp 1701859473
transform -1 0 3170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__973_
timestamp 1701859473
transform 1 0 3390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__974_
timestamp 1701859473
transform 1 0 3830 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__975_
timestamp 1701859473
transform 1 0 4830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__976_
timestamp 1701859473
transform -1 0 4870 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__977_
timestamp 1701859473
transform -1 0 2890 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__978_
timestamp 1701859473
transform -1 0 2590 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__979_
timestamp 1701859473
transform -1 0 2750 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__980_
timestamp 1701859473
transform 1 0 2310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__981_
timestamp 1701859473
transform 1 0 2450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__982_
timestamp 1701859473
transform -1 0 2610 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__983_
timestamp 1701859473
transform 1 0 3010 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__984_
timestamp 1701859473
transform 1 0 2710 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__985_
timestamp 1701859473
transform 1 0 3010 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__986_
timestamp 1701859473
transform 1 0 3110 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__987_
timestamp 1701859473
transform 1 0 3250 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__988_
timestamp 1701859473
transform 1 0 5170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__989_
timestamp 1701859473
transform -1 0 5190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__990_
timestamp 1701859473
transform -1 0 2490 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__991_
timestamp 1701859473
transform -1 0 3630 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__992_
timestamp 1701859473
transform 1 0 3310 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__993_
timestamp 1701859473
transform 1 0 1670 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__994_
timestamp 1701859473
transform -1 0 3490 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__995_
timestamp 1701859473
transform 1 0 3250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__996_
timestamp 1701859473
transform -1 0 3030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__997_
timestamp 1701859473
transform -1 0 2310 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__998_
timestamp 1701859473
transform -1 0 2750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__999_
timestamp 1701859473
transform 1 0 3090 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1000_
timestamp 1701859473
transform 1 0 3110 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1001_
timestamp 1701859473
transform 1 0 4070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1002_
timestamp 1701859473
transform 1 0 4870 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1003_
timestamp 1701859473
transform 1 0 4750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1004_
timestamp 1701859473
transform -1 0 3550 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1005_
timestamp 1701859473
transform 1 0 3390 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1006_
timestamp 1701859473
transform 1 0 4350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1007_
timestamp 1701859473
transform -1 0 4490 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1008_
timestamp 1701859473
transform 1 0 3370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1009_
timestamp 1701859473
transform -1 0 3950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1010_
timestamp 1701859473
transform -1 0 4230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1011_
timestamp 1701859473
transform -1 0 4050 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1012_
timestamp 1701859473
transform 1 0 4050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1013_
timestamp 1701859473
transform -1 0 4950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1014_
timestamp 1701859473
transform 1 0 4570 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1015_
timestamp 1701859473
transform 1 0 4190 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1016_
timestamp 1701859473
transform -1 0 4350 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1017_
timestamp 1701859473
transform -1 0 4210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1018_
timestamp 1701859473
transform -1 0 4090 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1019_
timestamp 1701859473
transform -1 0 3790 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1020_
timestamp 1701859473
transform -1 0 4250 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1021_
timestamp 1701859473
transform -1 0 3550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1022_
timestamp 1701859473
transform -1 0 3770 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1023_
timestamp 1701859473
transform 1 0 3890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1024_
timestamp 1701859473
transform 1 0 3770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1025_
timestamp 1701859473
transform -1 0 3490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1026_
timestamp 1701859473
transform 1 0 5350 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1027_
timestamp 1701859473
transform -1 0 5490 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1028_
timestamp 1701859473
transform 1 0 3670 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1029_
timestamp 1701859473
transform -1 0 3950 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1030_
timestamp 1701859473
transform 1 0 3810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1031_
timestamp 1701859473
transform 1 0 3630 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1032_
timestamp 1701859473
transform 1 0 3790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1033_
timestamp 1701859473
transform -1 0 3930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1034_
timestamp 1701859473
transform -1 0 3750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1035_
timestamp 1701859473
transform -1 0 3750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1036_
timestamp 1701859473
transform -1 0 3610 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1037_
timestamp 1701859473
transform 1 0 3250 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1038_
timestamp 1701859473
transform -1 0 2590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1039_
timestamp 1701859473
transform 1 0 3830 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1040_
timestamp 1701859473
transform -1 0 3910 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1041_
timestamp 1701859473
transform -1 0 2190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1042_
timestamp 1701859473
transform -1 0 1670 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1043_
timestamp 1701859473
transform -1 0 1550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1044_
timestamp 1701859473
transform -1 0 2050 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1045_
timestamp 1701859473
transform -1 0 1910 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1046_
timestamp 1701859473
transform 1 0 1790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1047_
timestamp 1701859473
transform -1 0 2070 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1048_
timestamp 1701859473
transform -1 0 1690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1049_
timestamp 1701859473
transform -1 0 2170 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1050_
timestamp 1701859473
transform 1 0 2030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1051_
timestamp 1701859473
transform -1 0 1930 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1052_
timestamp 1701859473
transform 1 0 1870 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1053_
timestamp 1701859473
transform 1 0 2850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1054_
timestamp 1701859473
transform -1 0 1430 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1055_
timestamp 1701859473
transform 1 0 1310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1056_
timestamp 1701859473
transform 1 0 1270 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1057_
timestamp 1701859473
transform 1 0 1430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1058_
timestamp 1701859473
transform 1 0 1310 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1059_
timestamp 1701859473
transform 1 0 1210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1060_
timestamp 1701859473
transform 1 0 1590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1061_
timestamp 1701859473
transform 1 0 1190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1062_
timestamp 1701859473
transform -1 0 850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1063_
timestamp 1701859473
transform 1 0 930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1064_
timestamp 1701859473
transform 1 0 1730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1065_
timestamp 1701859473
transform -1 0 3170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1066_
timestamp 1701859473
transform 1 0 2590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1067_
timestamp 1701859473
transform 1 0 1070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1068_
timestamp 1701859473
transform -1 0 1750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1069_
timestamp 1701859473
transform -1 0 2450 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1070_
timestamp 1701859473
transform 1 0 1790 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1071_
timestamp 1701859473
transform 1 0 2030 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1072_
timestamp 1701859473
transform 1 0 2190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1073_
timestamp 1701859473
transform 1 0 1990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1074_
timestamp 1701859473
transform 1 0 1590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1075_
timestamp 1701859473
transform 1 0 1890 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1076_
timestamp 1701859473
transform 1 0 2310 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1077_
timestamp 1701859473
transform 1 0 2730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1078_
timestamp 1701859473
transform 1 0 3690 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1079_
timestamp 1701859473
transform 1 0 3730 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1080_
timestamp 1701859473
transform 1 0 2170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1081_
timestamp 1701859473
transform 1 0 2330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1082_
timestamp 1701859473
transform -1 0 2890 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1083_
timestamp 1701859473
transform 1 0 2430 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1084_
timestamp 1701859473
transform 1 0 2590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1085_
timestamp 1701859473
transform 1 0 3010 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1086_
timestamp 1701859473
transform 1 0 2810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1087_
timestamp 1701859473
transform 1 0 2850 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1088_
timestamp 1701859473
transform -1 0 3930 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1089_
timestamp 1701859473
transform 1 0 3630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1090_
timestamp 1701859473
transform 1 0 2670 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1091_
timestamp 1701859473
transform 1 0 2290 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1092_
timestamp 1701859473
transform -1 0 2970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1093_
timestamp 1701859473
transform -1 0 2850 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1094_
timestamp 1701859473
transform 1 0 3770 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1095_
timestamp 1701859473
transform 1 0 4250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1096_
timestamp 1701859473
transform 1 0 4110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1097_
timestamp 1701859473
transform 1 0 1750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1098_
timestamp 1701859473
transform 1 0 3090 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1099_
timestamp 1701859473
transform 1 0 2710 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1100_
timestamp 1701859473
transform -1 0 2590 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1101_
timestamp 1701859473
transform -1 0 2470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1102_
timestamp 1701859473
transform -1 0 2150 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1103_
timestamp 1701859473
transform 1 0 1790 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1104_
timestamp 1701859473
transform -1 0 490 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1105_
timestamp 1701859473
transform -1 0 2090 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1106_
timestamp 1701859473
transform -1 0 1950 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1107_
timestamp 1701859473
transform -1 0 1950 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1108_
timestamp 1701859473
transform -1 0 1430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1109_
timestamp 1701859473
transform -1 0 1510 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1110_
timestamp 1701859473
transform -1 0 1270 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1111_
timestamp 1701859473
transform -1 0 1130 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1112_
timestamp 1701859473
transform -1 0 790 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1113_
timestamp 1701859473
transform -1 0 710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1114_
timestamp 1701859473
transform 1 0 1370 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1115_
timestamp 1701859473
transform -1 0 1130 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1116_
timestamp 1701859473
transform -1 0 1270 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1117_
timestamp 1701859473
transform -1 0 1110 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1118_
timestamp 1701859473
transform -1 0 970 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1119_
timestamp 1701859473
transform -1 0 590 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1120_
timestamp 1701859473
transform -1 0 1150 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1121_
timestamp 1701859473
transform -1 0 1030 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1122_
timestamp 1701859473
transform -1 0 1030 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1123_
timestamp 1701859473
transform -1 0 750 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1124_
timestamp 1701859473
transform -1 0 590 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1125_
timestamp 1701859473
transform 1 0 870 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1126_
timestamp 1701859473
transform -1 0 330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1127_
timestamp 1701859473
transform -1 0 610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1128_
timestamp 1701859473
transform -1 0 330 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1129_
timestamp 1701859473
transform 1 0 1450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1130_
timestamp 1701859473
transform -1 0 1550 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1131_
timestamp 1701859473
transform -1 0 470 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1132_
timestamp 1701859473
transform 1 0 30 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1133_
timestamp 1701859473
transform -1 0 450 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1134_
timestamp 1701859473
transform -1 0 190 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1__1135_
timestamp 1701859473
transform 1 0 170 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1136_
timestamp 1701859473
transform 1 0 170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1137_
timestamp 1701859473
transform -1 0 330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1138_
timestamp 1701859473
transform -1 0 50 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1139_
timestamp 1701859473
transform -1 0 50 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1140_
timestamp 1701859473
transform -1 0 190 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1141_
timestamp 1701859473
transform -1 0 330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1142_
timestamp 1701859473
transform 1 0 30 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1143_
timestamp 1701859473
transform -1 0 50 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1144_
timestamp 1701859473
transform 1 0 170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1145_
timestamp 1701859473
transform 1 0 390 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1146_
timestamp 1701859473
transform -1 0 1350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1147_
timestamp 1701859473
transform 1 0 1350 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1148_
timestamp 1701859473
transform 1 0 170 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1149_
timestamp 1701859473
transform -1 0 290 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1150_
timestamp 1701859473
transform -1 0 970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1151_
timestamp 1701859473
transform 1 0 670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1152_
timestamp 1701859473
transform -1 0 750 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1153_
timestamp 1701859473
transform -1 0 1790 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1154_
timestamp 1701859473
transform 1 0 1510 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1155_
timestamp 1701859473
transform 1 0 1330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1156_
timestamp 1701859473
transform -1 0 1390 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1157_
timestamp 1701859473
transform -1 0 1650 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1158_
timestamp 1701859473
transform -1 0 1250 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1159_
timestamp 1701859473
transform -1 0 1230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1160_
timestamp 1701859473
transform 1 0 1290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1161_
timestamp 1701859473
transform 1 0 1470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1162_
timestamp 1701859473
transform -1 0 1630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1163_
timestamp 1701859473
transform -1 0 1010 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1164_
timestamp 1701859473
transform 1 0 850 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1165_
timestamp 1701859473
transform -1 0 850 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1166_
timestamp 1701859473
transform -1 0 930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1167_
timestamp 1701859473
transform -1 0 790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1168_
timestamp 1701859473
transform 1 0 590 0 1 4950
box -12 -8 32 272
use FILL  FILL_1__1169_
timestamp 1701859473
transform -1 0 710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1170_
timestamp 1701859473
transform -1 0 610 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1171_
timestamp 1701859473
transform 1 0 550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1172_
timestamp 1701859473
transform -1 0 550 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1173_
timestamp 1701859473
transform -1 0 730 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1174_
timestamp 1701859473
transform 1 0 410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1__1175_
timestamp 1701859473
transform -1 0 470 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1176_
timestamp 1701859473
transform -1 0 210 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1177_
timestamp 1701859473
transform 1 0 30 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1178_
timestamp 1701859473
transform -1 0 470 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1179_
timestamp 1701859473
transform -1 0 350 0 1 4430
box -12 -8 32 272
use FILL  FILL_1__1180_
timestamp 1701859473
transform -1 0 330 0 1 3910
box -12 -8 32 272
use FILL  FILL_1__1181_
timestamp 1701859473
transform -1 0 50 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1182_
timestamp 1701859473
transform -1 0 50 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1183_
timestamp 1701859473
transform -1 0 310 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1184_
timestamp 1701859473
transform 1 0 150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1185_
timestamp 1701859473
transform 1 0 30 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1186_
timestamp 1701859473
transform -1 0 290 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1187_
timestamp 1701859473
transform 1 0 310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1188_
timestamp 1701859473
transform 1 0 30 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1189_
timestamp 1701859473
transform -1 0 170 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1190_
timestamp 1701859473
transform 1 0 210 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1191_
timestamp 1701859473
transform 1 0 290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1192_
timestamp 1701859473
transform -1 0 430 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1193_
timestamp 1701859473
transform -1 0 1070 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1194_
timestamp 1701859473
transform -1 0 1250 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1195_
timestamp 1701859473
transform -1 0 890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1__1196_
timestamp 1701859473
transform -1 0 1770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1197_
timestamp 1701859473
transform -1 0 1690 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1198_
timestamp 1701859473
transform -1 0 1570 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1199_
timestamp 1701859473
transform 1 0 1410 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1200_
timestamp 1701859473
transform -1 0 1110 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1201_
timestamp 1701859473
transform 1 0 950 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1202_
timestamp 1701859473
transform 1 0 810 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1203_
timestamp 1701859473
transform 1 0 990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1204_
timestamp 1701859473
transform 1 0 1090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1205_
timestamp 1701859473
transform -1 0 890 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1206_
timestamp 1701859473
transform -1 0 870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1207_
timestamp 1701859473
transform -1 0 730 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1208_
timestamp 1701859473
transform 1 0 570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1209_
timestamp 1701859473
transform -1 0 450 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1210_
timestamp 1701859473
transform 1 0 170 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1211_
timestamp 1701859473
transform 1 0 390 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1212_
timestamp 1701859473
transform 1 0 2950 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1213_
timestamp 1701859473
transform -1 0 3510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1214_
timestamp 1701859473
transform 1 0 510 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1215_
timestamp 1701859473
transform -1 0 670 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1216_
timestamp 1701859473
transform -1 0 170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1217_
timestamp 1701859473
transform -1 0 270 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1218_
timestamp 1701859473
transform -1 0 290 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1219_
timestamp 1701859473
transform 1 0 150 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1220_
timestamp 1701859473
transform 1 0 270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1221_
timestamp 1701859473
transform -1 0 990 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1222_
timestamp 1701859473
transform 1 0 1510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1223_
timestamp 1701859473
transform 1 0 1330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1224_
timestamp 1701859473
transform -1 0 1630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1225_
timestamp 1701859473
transform -1 0 1890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1226_
timestamp 1701859473
transform -1 0 1930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1227_
timestamp 1701859473
transform -1 0 1650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1228_
timestamp 1701859473
transform -1 0 1530 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1229_
timestamp 1701859473
transform 1 0 1110 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1230_
timestamp 1701859473
transform -1 0 690 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1231_
timestamp 1701859473
transform 1 0 30 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1232_
timestamp 1701859473
transform -1 0 150 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1233_
timestamp 1701859473
transform -1 0 50 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1234_
timestamp 1701859473
transform 1 0 30 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1235_
timestamp 1701859473
transform -1 0 50 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1236_
timestamp 1701859473
transform -1 0 50 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1237_
timestamp 1701859473
transform -1 0 190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1238_
timestamp 1701859473
transform -1 0 1210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1239_
timestamp 1701859473
transform 1 0 930 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1240_
timestamp 1701859473
transform -1 0 1090 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1241_
timestamp 1701859473
transform 1 0 430 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1242_
timestamp 1701859473
transform 1 0 790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1243_
timestamp 1701859473
transform 1 0 1290 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1244_
timestamp 1701859473
transform 1 0 1750 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1245_
timestamp 1701859473
transform 1 0 1770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1246_
timestamp 1701859473
transform -1 0 1530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1247_
timestamp 1701859473
transform 1 0 1210 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1248_
timestamp 1701859473
transform -1 0 1090 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1249_
timestamp 1701859473
transform 1 0 670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1250_
timestamp 1701859473
transform -1 0 590 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1251_
timestamp 1701859473
transform 1 0 650 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1252_
timestamp 1701859473
transform 1 0 510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1253_
timestamp 1701859473
transform -1 0 570 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1254_
timestamp 1701859473
transform -1 0 430 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1255_
timestamp 1701859473
transform 1 0 510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1256_
timestamp 1701859473
transform 1 0 750 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1257_
timestamp 1701859473
transform 1 0 790 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1258_
timestamp 1701859473
transform -1 0 950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1259_
timestamp 1701859473
transform -1 0 830 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1260_
timestamp 1701859473
transform 1 0 3410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1261_
timestamp 1701859473
transform -1 0 3410 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1262_
timestamp 1701859473
transform 1 0 3290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1263_
timestamp 1701859473
transform 1 0 3270 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1264_
timestamp 1701859473
transform -1 0 3190 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1265_
timestamp 1701859473
transform 1 0 3290 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1266_
timestamp 1701859473
transform 1 0 4270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1267_
timestamp 1701859473
transform 1 0 4010 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1268_
timestamp 1701859473
transform 1 0 4030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1269_
timestamp 1701859473
transform 1 0 3630 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1270_
timestamp 1701859473
transform 1 0 3510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1271_
timestamp 1701859473
transform -1 0 3770 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1272_
timestamp 1701859473
transform 1 0 3890 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1273_
timestamp 1701859473
transform -1 0 4330 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1274_
timestamp 1701859473
transform 1 0 4270 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1275_
timestamp 1701859473
transform -1 0 4150 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1276_
timestamp 1701859473
transform -1 0 5210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1277_
timestamp 1701859473
transform 1 0 5190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1278_
timestamp 1701859473
transform 1 0 5690 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1279_
timestamp 1701859473
transform 1 0 5670 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1280_
timestamp 1701859473
transform -1 0 4950 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1281_
timestamp 1701859473
transform 1 0 5050 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1282_
timestamp 1701859473
transform -1 0 5730 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1283_
timestamp 1701859473
transform -1 0 5630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1284_
timestamp 1701859473
transform -1 0 5730 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1285_
timestamp 1701859473
transform 1 0 5510 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1286_
timestamp 1701859473
transform 1 0 5330 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1287_
timestamp 1701859473
transform -1 0 5550 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1288_
timestamp 1701859473
transform 1 0 4070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1289_
timestamp 1701859473
transform 1 0 5210 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1290_
timestamp 1701859473
transform 1 0 5330 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1291_
timestamp 1701859473
transform -1 0 5070 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1292_
timestamp 1701859473
transform 1 0 4930 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1293_
timestamp 1701859473
transform -1 0 5670 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1294_
timestamp 1701859473
transform -1 0 5530 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1295_
timestamp 1701859473
transform -1 0 5170 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1296_
timestamp 1701859473
transform 1 0 5030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1297_
timestamp 1701859473
transform 1 0 5250 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1298_
timestamp 1701859473
transform -1 0 5030 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1299_
timestamp 1701859473
transform -1 0 4210 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1300_
timestamp 1701859473
transform 1 0 5170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1301_
timestamp 1701859473
transform 1 0 5370 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1302_
timestamp 1701859473
transform 1 0 5310 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1303_
timestamp 1701859473
transform 1 0 5190 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1304_
timestamp 1701859473
transform -1 0 5210 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1305_
timestamp 1701859473
transform 1 0 5470 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1306_
timestamp 1701859473
transform 1 0 5590 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1307_
timestamp 1701859473
transform -1 0 5150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1308_
timestamp 1701859473
transform 1 0 5230 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1309_
timestamp 1701859473
transform -1 0 5390 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1310_
timestamp 1701859473
transform -1 0 4490 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1311_
timestamp 1701859473
transform -1 0 4890 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1312_
timestamp 1701859473
transform 1 0 4250 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1313_
timestamp 1701859473
transform 1 0 4750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1314_
timestamp 1701859473
transform 1 0 4610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1315_
timestamp 1701859473
transform -1 0 4690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1316_
timestamp 1701859473
transform -1 0 4550 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1317_
timestamp 1701859473
transform 1 0 3930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1318_
timestamp 1701859473
transform 1 0 4370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1319_
timestamp 1701859473
transform -1 0 4510 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1320_
timestamp 1701859473
transform 1 0 4610 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1321_
timestamp 1701859473
transform 1 0 4690 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1322_
timestamp 1701859473
transform 1 0 3970 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1323_
timestamp 1701859473
transform 1 0 4730 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1324_
timestamp 1701859473
transform 1 0 4590 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1325_
timestamp 1701859473
transform 1 0 2170 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1326_
timestamp 1701859473
transform -1 0 4930 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1327_
timestamp 1701859473
transform -1 0 4450 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1328_
timestamp 1701859473
transform 1 0 4550 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1329_
timestamp 1701859473
transform 1 0 4390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1330_
timestamp 1701859473
transform -1 0 4630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1331_
timestamp 1701859473
transform -1 0 4830 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1332_
timestamp 1701859473
transform -1 0 4690 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1333_
timestamp 1701859473
transform 1 0 4550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1334_
timestamp 1701859473
transform -1 0 1650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1335_
timestamp 1701859473
transform -1 0 1790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1336_
timestamp 1701859473
transform 1 0 1610 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1337_
timestamp 1701859473
transform 1 0 1930 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1338_
timestamp 1701859473
transform 1 0 1870 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1339_
timestamp 1701859473
transform -1 0 1850 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1340_
timestamp 1701859473
transform -1 0 1750 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1341_
timestamp 1701859473
transform 1 0 2030 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1342_
timestamp 1701859473
transform -1 0 1610 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1343_
timestamp 1701859473
transform -1 0 1010 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1344_
timestamp 1701859473
transform -1 0 870 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1345_
timestamp 1701859473
transform 1 0 1110 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1346_
timestamp 1701859473
transform -1 0 1230 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1347_
timestamp 1701859473
transform 1 0 1270 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1348_
timestamp 1701859473
transform 1 0 1650 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1349_
timestamp 1701859473
transform -1 0 2450 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1350_
timestamp 1701859473
transform 1 0 2050 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1351_
timestamp 1701859473
transform -1 0 2690 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1352_
timestamp 1701859473
transform 1 0 1510 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1353_
timestamp 1701859473
transform -1 0 1350 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1354_
timestamp 1701859473
transform -1 0 1390 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1355_
timestamp 1701859473
transform -1 0 290 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1356_
timestamp 1701859473
transform -1 0 410 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1357_
timestamp 1701859473
transform 1 0 290 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1358_
timestamp 1701859473
transform 1 0 410 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1359_
timestamp 1701859473
transform 1 0 1870 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1360_
timestamp 1701859473
transform -1 0 1750 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1361_
timestamp 1701859473
transform 1 0 2290 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1362_
timestamp 1701859473
transform -1 0 1250 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1363_
timestamp 1701859473
transform 1 0 1110 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1364_
timestamp 1701859473
transform -1 0 770 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1365_
timestamp 1701859473
transform -1 0 650 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1366_
timestamp 1701859473
transform 1 0 630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1367_
timestamp 1701859473
transform -1 0 670 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1368_
timestamp 1701859473
transform -1 0 950 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1369_
timestamp 1701859473
transform -1 0 1510 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1370_
timestamp 1701859473
transform 1 0 1350 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1371_
timestamp 1701859473
transform 1 0 530 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1372_
timestamp 1701859473
transform -1 0 810 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1373_
timestamp 1701859473
transform -1 0 530 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1374_
timestamp 1701859473
transform 1 0 630 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1375_
timestamp 1701859473
transform -1 0 190 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1376_
timestamp 1701859473
transform 1 0 390 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1377_
timestamp 1701859473
transform -1 0 310 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1378_
timestamp 1701859473
transform -1 0 50 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1379_
timestamp 1701859473
transform 1 0 30 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1380_
timestamp 1701859473
transform 1 0 30 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1381_
timestamp 1701859473
transform 1 0 30 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1382_
timestamp 1701859473
transform 1 0 130 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1383_
timestamp 1701859473
transform 1 0 150 0 -1 790
box -12 -8 32 272
use FILL  FILL_1__1384_
timestamp 1701859473
transform 1 0 130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1385_
timestamp 1701859473
transform -1 0 870 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1386_
timestamp 1701859473
transform -1 0 890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1387_
timestamp 1701859473
transform -1 0 770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1388_
timestamp 1701859473
transform -1 0 550 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1389_
timestamp 1701859473
transform 1 0 290 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1390_
timestamp 1701859473
transform 1 0 450 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1391_
timestamp 1701859473
transform -1 0 610 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1392_
timestamp 1701859473
transform -1 0 410 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1393_
timestamp 1701859473
transform 1 0 390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1394_
timestamp 1701859473
transform -1 0 290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1395_
timestamp 1701859473
transform 1 0 490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1396_
timestamp 1701859473
transform 1 0 870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1397_
timestamp 1701859473
transform -1 0 990 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1398_
timestamp 1701859473
transform -1 0 1250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1399_
timestamp 1701859473
transform -1 0 1090 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1400_
timestamp 1701859473
transform -1 0 1550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1401_
timestamp 1701859473
transform 1 0 1110 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1402_
timestamp 1701859473
transform 1 0 1250 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1403_
timestamp 1701859473
transform 1 0 1390 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1404_
timestamp 1701859473
transform 1 0 1370 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1405_
timestamp 1701859473
transform -1 0 3190 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1406_
timestamp 1701859473
transform 1 0 2450 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1407_
timestamp 1701859473
transform 1 0 2110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1408_
timestamp 1701859473
transform -1 0 2250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1409_
timestamp 1701859473
transform 1 0 3450 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1410_
timestamp 1701859473
transform 1 0 2410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1411_
timestamp 1701859473
transform -1 0 2550 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1412_
timestamp 1701859473
transform -1 0 3570 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1413_
timestamp 1701859473
transform 1 0 2070 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1414_
timestamp 1701859473
transform -1 0 2210 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1415_
timestamp 1701859473
transform -1 0 3730 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1416_
timestamp 1701859473
transform 1 0 2370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1417_
timestamp 1701859473
transform -1 0 2590 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1418_
timestamp 1701859473
transform 1 0 3210 0 1 270
box -12 -8 32 272
use FILL  FILL_1__1419_
timestamp 1701859473
transform 1 0 2130 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1420_
timestamp 1701859473
transform -1 0 2270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1421_
timestamp 1701859473
transform 1 0 2210 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1422_
timestamp 1701859473
transform -1 0 2590 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1423_
timestamp 1701859473
transform -1 0 2730 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1424_
timestamp 1701859473
transform -1 0 3090 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1425_
timestamp 1701859473
transform 1 0 2390 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1426_
timestamp 1701859473
transform -1 0 2770 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1427_
timestamp 1701859473
transform 1 0 2730 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1428_
timestamp 1701859473
transform 1 0 3130 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1429_
timestamp 1701859473
transform 1 0 3270 0 1 1830
box -12 -8 32 272
use FILL  FILL_1__1430_
timestamp 1701859473
transform 1 0 3250 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1431_
timestamp 1701859473
transform -1 0 3390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1432_
timestamp 1701859473
transform -1 0 3250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1433_
timestamp 1701859473
transform 1 0 3090 0 -1 2350
box -12 -8 32 272
use FILL  FILL_1__1434_
timestamp 1701859473
transform -1 0 3130 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1435_
timestamp 1701859473
transform 1 0 2950 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1436_
timestamp 1701859473
transform 1 0 2750 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1437_
timestamp 1701859473
transform -1 0 2630 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1__1438_
timestamp 1701859473
transform 1 0 2930 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1439_
timestamp 1701859473
transform 1 0 2790 0 -1 1310
box -12 -8 32 272
use FILL  FILL_1__1440_
timestamp 1701859473
transform -1 0 3870 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1441_
timestamp 1701859473
transform 1 0 3470 0 1 1310
box -12 -8 32 272
use FILL  FILL_1__1442_
timestamp 1701859473
transform 1 0 3510 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1__1443_
timestamp 1701859473
transform -1 0 3410 0 1 2350
box -12 -8 32 272
use FILL  FILL_1__1444_
timestamp 1701859473
transform -1 0 2470 0 1 3390
box -12 -8 32 272
use FILL  FILL_1__1445_
timestamp 1701859473
transform -1 0 2630 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1446_
timestamp 1701859473
transform -1 0 2870 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1447_
timestamp 1701859473
transform -1 0 2990 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1448_
timestamp 1701859473
transform -1 0 2410 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1449_
timestamp 1701859473
transform -1 0 2770 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1450_
timestamp 1701859473
transform -1 0 2010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1451_
timestamp 1701859473
transform 1 0 1870 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1527_
timestamp 1701859473
transform 1 0 5690 0 1 790
box -12 -8 32 272
use FILL  FILL_1__1528_
timestamp 1701859473
transform -1 0 5710 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1529_
timestamp 1701859473
transform 1 0 5390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1__1530_
timestamp 1701859473
transform 1 0 5130 0 1 2870
box -12 -8 32 272
use FILL  FILL_1__1531_
timestamp 1701859473
transform 1 0 2770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_1__1532_
timestamp 1701859473
transform 1 0 3810 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1533_
timestamp 1701859473
transform 1 0 4070 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1534_
timestamp 1701859473
transform 1 0 4190 0 -1 270
box -12 -8 32 272
use FILL  FILL_1__1535_
timestamp 1701859473
transform 1 0 3950 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert0
timestamp 1701859473
transform -1 0 1490 0 1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert1
timestamp 1701859473
transform 1 0 2150 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert2
timestamp 1701859473
transform 1 0 4790 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert3
timestamp 1701859473
transform 1 0 3670 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert4
timestamp 1701859473
transform 1 0 2150 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert5
timestamp 1701859473
transform 1 0 4150 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert6
timestamp 1701859473
transform -1 0 1370 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert15
timestamp 1701859473
transform -1 0 4750 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert16
timestamp 1701859473
transform -1 0 3530 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert17
timestamp 1701859473
transform -1 0 3970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert18
timestamp 1701859473
transform 1 0 4910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert19
timestamp 1701859473
transform -1 0 1630 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert20
timestamp 1701859473
transform -1 0 4370 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert21
timestamp 1701859473
transform -1 0 1810 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert22
timestamp 1701859473
transform -1 0 4850 0 1 1830
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert23
timestamp 1701859473
transform -1 0 3070 0 -1 790
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert24
timestamp 1701859473
transform 1 0 5050 0 1 270
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert25
timestamp 1701859473
transform -1 0 3030 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert26
timestamp 1701859473
transform 1 0 3010 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert27
timestamp 1701859473
transform 1 0 3150 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert28
timestamp 1701859473
transform 1 0 2630 0 1 1310
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert29
timestamp 1701859473
transform -1 0 2510 0 -1 3390
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert30
timestamp 1701859473
transform -1 0 4350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert31
timestamp 1701859473
transform -1 0 3490 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert32
timestamp 1701859473
transform 1 0 4610 0 1 4950
box -12 -8 32 272
use FILL  FILL_1_BUFX2_insert33
timestamp 1701859473
transform -1 0 4390 0 1 4430
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 2790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert8
timestamp 1701859473
transform -1 0 1610 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 1750 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert10
timestamp 1701859473
transform -1 0 2350 0 1 2350
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert11
timestamp 1701859473
transform 1 0 4270 0 1 790
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert12
timestamp 1701859473
transform -1 0 3230 0 -1 270
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert13
timestamp 1701859473
transform 1 0 2870 0 -1 1830
box -12 -8 32 272
use FILL  FILL_1_CLKBUF1_insert14
timestamp 1701859473
transform 1 0 4950 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__723_
timestamp 1701859473
transform -1 0 2830 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__724_
timestamp 1701859473
transform -1 0 2630 0 1 790
box -12 -8 32 272
use FILL  FILL_2__725_
timestamp 1701859473
transform -1 0 2710 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__726_
timestamp 1701859473
transform 1 0 3350 0 1 270
box -12 -8 32 272
use FILL  FILL_2__727_
timestamp 1701859473
transform 1 0 2910 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__728_
timestamp 1701859473
transform -1 0 3050 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__729_
timestamp 1701859473
transform 1 0 3690 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__730_
timestamp 1701859473
transform 1 0 3590 0 1 270
box -12 -8 32 272
use FILL  FILL_2__731_
timestamp 1701859473
transform -1 0 3510 0 1 270
box -12 -8 32 272
use FILL  FILL_2__732_
timestamp 1701859473
transform -1 0 790 0 1 790
box -12 -8 32 272
use FILL  FILL_2__733_
timestamp 1701859473
transform -1 0 2010 0 1 790
box -12 -8 32 272
use FILL  FILL_2__734_
timestamp 1701859473
transform -1 0 2970 0 1 270
box -12 -8 32 272
use FILL  FILL_2__735_
timestamp 1701859473
transform 1 0 4110 0 1 270
box -12 -8 32 272
use FILL  FILL_2__736_
timestamp 1701859473
transform 1 0 3830 0 1 270
box -12 -8 32 272
use FILL  FILL_2__737_
timestamp 1701859473
transform 1 0 990 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__738_
timestamp 1701859473
transform -1 0 2130 0 1 790
box -12 -8 32 272
use FILL  FILL_2__739_
timestamp 1701859473
transform -1 0 2830 0 1 270
box -12 -8 32 272
use FILL  FILL_2__740_
timestamp 1701859473
transform 1 0 4670 0 1 270
box -12 -8 32 272
use FILL  FILL_2__741_
timestamp 1701859473
transform 1 0 3970 0 1 270
box -12 -8 32 272
use FILL  FILL_2__742_
timestamp 1701859473
transform -1 0 2950 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__743_
timestamp 1701859473
transform 1 0 3090 0 1 270
box -12 -8 32 272
use FILL  FILL_2__744_
timestamp 1701859473
transform -1 0 4470 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__745_
timestamp 1701859473
transform 1 0 3690 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__746_
timestamp 1701859473
transform 1 0 2290 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__747_
timestamp 1701859473
transform 1 0 3290 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__748_
timestamp 1701859473
transform 1 0 3150 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__749_
timestamp 1701859473
transform 1 0 2190 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__750_
timestamp 1701859473
transform -1 0 3270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__751_
timestamp 1701859473
transform 1 0 3390 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__752_
timestamp 1701859473
transform 1 0 1670 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__753_
timestamp 1701859473
transform 1 0 3550 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__754_
timestamp 1701859473
transform 1 0 3410 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__755_
timestamp 1701859473
transform -1 0 1450 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__756_
timestamp 1701859473
transform 1 0 2670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__757_
timestamp 1701859473
transform 1 0 2510 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__758_
timestamp 1701859473
transform -1 0 2370 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__759_
timestamp 1701859473
transform 1 0 2210 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__760_
timestamp 1701859473
transform -1 0 2170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__761_
timestamp 1701859473
transform 1 0 2070 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__762_
timestamp 1701859473
transform -1 0 2170 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__763_
timestamp 1701859473
transform -1 0 2290 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__764_
timestamp 1701859473
transform 1 0 2030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__765_
timestamp 1701859473
transform -1 0 2170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__766_
timestamp 1701859473
transform 1 0 3390 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__767_
timestamp 1701859473
transform 1 0 2770 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__768_
timestamp 1701859473
transform -1 0 2910 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__769_
timestamp 1701859473
transform -1 0 4210 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__770_
timestamp 1701859473
transform -1 0 3570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__771_
timestamp 1701859473
transform -1 0 3690 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__772_
timestamp 1701859473
transform -1 0 5430 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__773_
timestamp 1701859473
transform -1 0 4310 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__774_
timestamp 1701859473
transform -1 0 4830 0 1 790
box -12 -8 32 272
use FILL  FILL_2__775_
timestamp 1701859473
transform -1 0 5770 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__776_
timestamp 1701859473
transform 1 0 4930 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__777_
timestamp 1701859473
transform 1 0 5710 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__778_
timestamp 1701859473
transform 1 0 5390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__779_
timestamp 1701859473
transform -1 0 4370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__780_
timestamp 1701859473
transform -1 0 4790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__781_
timestamp 1701859473
transform -1 0 5130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__782_
timestamp 1701859473
transform -1 0 3790 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__783_
timestamp 1701859473
transform -1 0 4990 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__784_
timestamp 1701859473
transform 1 0 3850 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__785_
timestamp 1701859473
transform -1 0 3450 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__786_
timestamp 1701859473
transform -1 0 3490 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__787_
timestamp 1701859473
transform -1 0 4230 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__788_
timestamp 1701859473
transform -1 0 3570 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__789_
timestamp 1701859473
transform -1 0 3850 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__790_
timestamp 1701859473
transform 1 0 1910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__791_
timestamp 1701859473
transform -1 0 2170 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__792_
timestamp 1701859473
transform 1 0 2010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__793_
timestamp 1701859473
transform 1 0 1010 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__794_
timestamp 1701859473
transform 1 0 1630 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__795_
timestamp 1701859473
transform -1 0 1370 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__796_
timestamp 1701859473
transform -1 0 550 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__797_
timestamp 1701859473
transform 1 0 1510 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__798_
timestamp 1701859473
transform 1 0 870 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__799_
timestamp 1701859473
transform 1 0 1530 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__800_
timestamp 1701859473
transform 1 0 2290 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__801_
timestamp 1701859473
transform 1 0 2030 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__802_
timestamp 1701859473
transform -1 0 450 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__803_
timestamp 1701859473
transform -1 0 1250 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__804_
timestamp 1701859473
transform 1 0 690 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__805_
timestamp 1701859473
transform -1 0 1010 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__806_
timestamp 1701859473
transform 1 0 2270 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__807_
timestamp 1701859473
transform 1 0 1110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__808_
timestamp 1701859473
transform 1 0 1010 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__809_
timestamp 1701859473
transform 1 0 1490 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__810_
timestamp 1701859473
transform -1 0 1510 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__811_
timestamp 1701859473
transform -1 0 1350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__812_
timestamp 1701859473
transform 1 0 2290 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__813_
timestamp 1701859473
transform 1 0 1670 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__814_
timestamp 1701859473
transform 1 0 3370 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__815_
timestamp 1701859473
transform 1 0 3670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__816_
timestamp 1701859473
transform 1 0 3550 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__817_
timestamp 1701859473
transform 1 0 4470 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__818_
timestamp 1701859473
transform -1 0 4110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__819_
timestamp 1701859473
transform 1 0 3670 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__820_
timestamp 1701859473
transform -1 0 4250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__821_
timestamp 1701859473
transform 1 0 4090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__822_
timestamp 1701859473
transform -1 0 4230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__823_
timestamp 1701859473
transform 1 0 4410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__824_
timestamp 1701859473
transform 1 0 3990 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__825_
timestamp 1701859473
transform -1 0 4130 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__826_
timestamp 1701859473
transform -1 0 4230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__827_
timestamp 1701859473
transform -1 0 3930 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__828_
timestamp 1701859473
transform 1 0 4170 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__829_
timestamp 1701859473
transform 1 0 3790 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__830_
timestamp 1701859473
transform -1 0 4230 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__831_
timestamp 1701859473
transform 1 0 4090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__832_
timestamp 1701859473
transform -1 0 4110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__833_
timestamp 1701859473
transform -1 0 3150 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__834_
timestamp 1701859473
transform 1 0 3390 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__835_
timestamp 1701859473
transform 1 0 3670 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__836_
timestamp 1701859473
transform 1 0 3530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__837_
timestamp 1701859473
transform 1 0 3890 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__838_
timestamp 1701859473
transform 1 0 4670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__839_
timestamp 1701859473
transform -1 0 4990 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__840_
timestamp 1701859473
transform 1 0 4530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__841_
timestamp 1701859473
transform 1 0 4810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__842_
timestamp 1701859473
transform -1 0 5130 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__843_
timestamp 1701859473
transform -1 0 4630 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__844_
timestamp 1701859473
transform -1 0 4750 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__845_
timestamp 1701859473
transform -1 0 5730 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__846_
timestamp 1701859473
transform -1 0 3410 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__847_
timestamp 1701859473
transform 1 0 4030 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__848_
timestamp 1701859473
transform 1 0 4350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__849_
timestamp 1701859473
transform 1 0 4530 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__850_
timestamp 1701859473
transform -1 0 4270 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__851_
timestamp 1701859473
transform 1 0 4490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__852_
timestamp 1701859473
transform 1 0 4590 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__853_
timestamp 1701859473
transform 1 0 4370 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__854_
timestamp 1701859473
transform 1 0 4290 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__855_
timestamp 1701859473
transform 1 0 4170 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__856_
timestamp 1701859473
transform 1 0 4470 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__857_
timestamp 1701859473
transform 1 0 4610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__858_
timestamp 1701859473
transform -1 0 4630 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__859_
timestamp 1701859473
transform -1 0 4090 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__860_
timestamp 1701859473
transform -1 0 4490 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__861_
timestamp 1701859473
transform 1 0 3390 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__862_
timestamp 1701859473
transform 1 0 3630 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__863_
timestamp 1701859473
transform -1 0 2410 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__864_
timestamp 1701859473
transform -1 0 4670 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__865_
timestamp 1701859473
transform 1 0 3890 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__866_
timestamp 1701859473
transform 1 0 4030 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__867_
timestamp 1701859473
transform 1 0 4330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__868_
timestamp 1701859473
transform 1 0 4470 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__869_
timestamp 1701859473
transform 1 0 4870 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__870_
timestamp 1701859473
transform 1 0 4750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__871_
timestamp 1701859473
transform 1 0 4310 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__872_
timestamp 1701859473
transform 1 0 4750 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__873_
timestamp 1701859473
transform 1 0 5070 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__874_
timestamp 1701859473
transform 1 0 5210 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__875_
timestamp 1701859473
transform 1 0 5050 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__876_
timestamp 1701859473
transform -1 0 5190 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__877_
timestamp 1701859473
transform -1 0 5490 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__878_
timestamp 1701859473
transform 1 0 5350 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__879_
timestamp 1701859473
transform 1 0 4890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__880_
timestamp 1701859473
transform 1 0 5030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__881_
timestamp 1701859473
transform 1 0 4650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__882_
timestamp 1701859473
transform -1 0 4770 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__883_
timestamp 1701859473
transform 1 0 4430 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__884_
timestamp 1701859473
transform -1 0 4390 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__885_
timestamp 1701859473
transform -1 0 4570 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__886_
timestamp 1701859473
transform 1 0 4230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__887_
timestamp 1701859473
transform -1 0 5090 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__888_
timestamp 1701859473
transform -1 0 4950 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__889_
timestamp 1701859473
transform 1 0 4730 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__890_
timestamp 1701859473
transform 1 0 4790 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__891_
timestamp 1701859473
transform -1 0 4670 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__892_
timestamp 1701859473
transform 1 0 4910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__893_
timestamp 1701859473
transform 1 0 4730 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__894_
timestamp 1701859473
transform 1 0 5070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__895_
timestamp 1701859473
transform 1 0 4790 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__896_
timestamp 1701859473
transform 1 0 5110 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__897_
timestamp 1701859473
transform 1 0 3350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__898_
timestamp 1701859473
transform 1 0 2770 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__899_
timestamp 1701859473
transform 1 0 1790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__900_
timestamp 1701859473
transform -1 0 3310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__901_
timestamp 1701859473
transform 1 0 3230 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__902_
timestamp 1701859473
transform -1 0 3490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__903_
timestamp 1701859473
transform -1 0 5210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__904_
timestamp 1701859473
transform 1 0 4970 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__905_
timestamp 1701859473
transform 1 0 5050 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__906_
timestamp 1701859473
transform 1 0 5470 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__907_
timestamp 1701859473
transform -1 0 5270 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__908_
timestamp 1701859473
transform 1 0 5170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__909_
timestamp 1701859473
transform -1 0 5050 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__910_
timestamp 1701859473
transform 1 0 4890 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__911_
timestamp 1701859473
transform -1 0 5410 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__912_
timestamp 1701859473
transform 1 0 5310 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__913_
timestamp 1701859473
transform -1 0 5290 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__914_
timestamp 1701859473
transform 1 0 5470 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__915_
timestamp 1701859473
transform 1 0 5610 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__916_
timestamp 1701859473
transform 1 0 5570 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__917_
timestamp 1701859473
transform 1 0 5470 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__918_
timestamp 1701859473
transform -1 0 3630 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__919_
timestamp 1701859473
transform 1 0 4790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__920_
timestamp 1701859473
transform 1 0 5710 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__921_
timestamp 1701859473
transform 1 0 5530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__922_
timestamp 1701859473
transform 1 0 2610 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__923_
timestamp 1701859473
transform -1 0 3090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__924_
timestamp 1701859473
transform -1 0 2930 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__925_
timestamp 1701859473
transform -1 0 2530 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__926_
timestamp 1701859473
transform 1 0 2970 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__927_
timestamp 1701859473
transform 1 0 2830 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__928_
timestamp 1701859473
transform 1 0 2730 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__929_
timestamp 1701859473
transform -1 0 3130 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__930_
timestamp 1701859473
transform 1 0 3210 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__931_
timestamp 1701859473
transform 1 0 3230 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__932_
timestamp 1701859473
transform -1 0 4550 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__933_
timestamp 1701859473
transform 1 0 4910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__934_
timestamp 1701859473
transform 1 0 5230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__935_
timestamp 1701859473
transform -1 0 4490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__936_
timestamp 1701859473
transform 1 0 5310 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__937_
timestamp 1701859473
transform 1 0 5070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__938_
timestamp 1701859473
transform 1 0 5050 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__939_
timestamp 1701859473
transform -1 0 5470 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__940_
timestamp 1701859473
transform 1 0 5750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__941_
timestamp 1701859473
transform -1 0 4530 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__942_
timestamp 1701859473
transform -1 0 4670 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__943_
timestamp 1701859473
transform 1 0 5010 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__944_
timestamp 1701859473
transform -1 0 5350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__945_
timestamp 1701859473
transform 1 0 5330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__946_
timestamp 1701859473
transform 1 0 5470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__947_
timestamp 1701859473
transform 1 0 5610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__948_
timestamp 1701859473
transform -1 0 5630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__949_
timestamp 1701859473
transform -1 0 5450 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__950_
timestamp 1701859473
transform 1 0 4650 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__951_
timestamp 1701859473
transform -1 0 5110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__952_
timestamp 1701859473
transform -1 0 5490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__953_
timestamp 1701859473
transform 1 0 5150 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__954_
timestamp 1701859473
transform 1 0 5450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__955_
timestamp 1701859473
transform 1 0 5330 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__956_
timestamp 1701859473
transform 1 0 5290 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__957_
timestamp 1701859473
transform 1 0 5570 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__958_
timestamp 1701859473
transform -1 0 5630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__959_
timestamp 1701859473
transform 1 0 5610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__960_
timestamp 1701859473
transform 1 0 5310 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__961_
timestamp 1701859473
transform -1 0 5650 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__962_
timestamp 1701859473
transform 1 0 5570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__963_
timestamp 1701859473
transform -1 0 5690 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__964_
timestamp 1701859473
transform 1 0 5410 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__965_
timestamp 1701859473
transform 1 0 5530 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__966_
timestamp 1701859473
transform 1 0 4690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__967_
timestamp 1701859473
transform -1 0 4570 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__968_
timestamp 1701859473
transform -1 0 4190 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__969_
timestamp 1701859473
transform -1 0 5550 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__970_
timestamp 1701859473
transform 1 0 5170 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__971_
timestamp 1701859473
transform 1 0 5230 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__972_
timestamp 1701859473
transform -1 0 3190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__973_
timestamp 1701859473
transform 1 0 3410 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__974_
timestamp 1701859473
transform 1 0 3850 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__975_
timestamp 1701859473
transform 1 0 4850 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__976_
timestamp 1701859473
transform -1 0 4890 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__977_
timestamp 1701859473
transform -1 0 2910 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__978_
timestamp 1701859473
transform -1 0 2610 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__979_
timestamp 1701859473
transform -1 0 2770 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__980_
timestamp 1701859473
transform 1 0 2330 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__981_
timestamp 1701859473
transform 1 0 2470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__982_
timestamp 1701859473
transform -1 0 2630 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__983_
timestamp 1701859473
transform 1 0 3030 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__984_
timestamp 1701859473
transform 1 0 2730 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__985_
timestamp 1701859473
transform 1 0 3030 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__986_
timestamp 1701859473
transform 1 0 3130 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__987_
timestamp 1701859473
transform 1 0 3270 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__988_
timestamp 1701859473
transform 1 0 5190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__989_
timestamp 1701859473
transform -1 0 5210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__990_
timestamp 1701859473
transform -1 0 2510 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__991_
timestamp 1701859473
transform -1 0 3650 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__992_
timestamp 1701859473
transform 1 0 3330 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__993_
timestamp 1701859473
transform 1 0 1690 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__994_
timestamp 1701859473
transform -1 0 3510 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__995_
timestamp 1701859473
transform 1 0 3270 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__996_
timestamp 1701859473
transform -1 0 3050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__997_
timestamp 1701859473
transform -1 0 2330 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__998_
timestamp 1701859473
transform -1 0 2770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__999_
timestamp 1701859473
transform 1 0 3110 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1000_
timestamp 1701859473
transform 1 0 3130 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1001_
timestamp 1701859473
transform 1 0 4090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1002_
timestamp 1701859473
transform 1 0 4890 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1003_
timestamp 1701859473
transform 1 0 4770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1004_
timestamp 1701859473
transform -1 0 3570 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1005_
timestamp 1701859473
transform 1 0 3410 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1006_
timestamp 1701859473
transform 1 0 4370 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1007_
timestamp 1701859473
transform -1 0 4510 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1008_
timestamp 1701859473
transform 1 0 3390 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1009_
timestamp 1701859473
transform -1 0 3970 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1010_
timestamp 1701859473
transform -1 0 4250 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1011_
timestamp 1701859473
transform -1 0 4070 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1012_
timestamp 1701859473
transform 1 0 4070 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1013_
timestamp 1701859473
transform -1 0 4970 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1014_
timestamp 1701859473
transform 1 0 4590 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1015_
timestamp 1701859473
transform 1 0 4210 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1016_
timestamp 1701859473
transform -1 0 4370 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1017_
timestamp 1701859473
transform -1 0 4230 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1018_
timestamp 1701859473
transform -1 0 4110 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1019_
timestamp 1701859473
transform -1 0 3810 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1020_
timestamp 1701859473
transform -1 0 4270 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1021_
timestamp 1701859473
transform -1 0 3570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1022_
timestamp 1701859473
transform -1 0 3790 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1023_
timestamp 1701859473
transform 1 0 3910 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1024_
timestamp 1701859473
transform 1 0 3790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1025_
timestamp 1701859473
transform -1 0 3510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1026_
timestamp 1701859473
transform 1 0 5370 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1027_
timestamp 1701859473
transform -1 0 5510 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1028_
timestamp 1701859473
transform 1 0 3690 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1029_
timestamp 1701859473
transform -1 0 3970 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1030_
timestamp 1701859473
transform 1 0 3830 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1031_
timestamp 1701859473
transform 1 0 3650 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1032_
timestamp 1701859473
transform 1 0 3810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1033_
timestamp 1701859473
transform -1 0 3950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1034_
timestamp 1701859473
transform -1 0 3770 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1035_
timestamp 1701859473
transform -1 0 3770 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1036_
timestamp 1701859473
transform -1 0 3630 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1037_
timestamp 1701859473
transform 1 0 3270 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1038_
timestamp 1701859473
transform -1 0 2610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1039_
timestamp 1701859473
transform 1 0 3850 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1040_
timestamp 1701859473
transform -1 0 3930 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1041_
timestamp 1701859473
transform -1 0 2210 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1042_
timestamp 1701859473
transform -1 0 1690 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1043_
timestamp 1701859473
transform -1 0 1570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1044_
timestamp 1701859473
transform -1 0 2070 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1045_
timestamp 1701859473
transform -1 0 1930 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1046_
timestamp 1701859473
transform 1 0 1810 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1047_
timestamp 1701859473
transform -1 0 2090 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1048_
timestamp 1701859473
transform -1 0 1710 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1049_
timestamp 1701859473
transform -1 0 2190 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1050_
timestamp 1701859473
transform 1 0 2050 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1051_
timestamp 1701859473
transform -1 0 1950 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1052_
timestamp 1701859473
transform 1 0 1890 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1053_
timestamp 1701859473
transform 1 0 2870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1054_
timestamp 1701859473
transform -1 0 1450 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1055_
timestamp 1701859473
transform 1 0 1330 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1056_
timestamp 1701859473
transform 1 0 1290 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1057_
timestamp 1701859473
transform 1 0 1450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1058_
timestamp 1701859473
transform 1 0 1330 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1059_
timestamp 1701859473
transform 1 0 1230 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1060_
timestamp 1701859473
transform 1 0 1610 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1061_
timestamp 1701859473
transform 1 0 1210 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1062_
timestamp 1701859473
transform -1 0 870 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1063_
timestamp 1701859473
transform 1 0 950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1064_
timestamp 1701859473
transform 1 0 1750 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1065_
timestamp 1701859473
transform -1 0 3190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1066_
timestamp 1701859473
transform 1 0 2610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1067_
timestamp 1701859473
transform 1 0 1090 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1068_
timestamp 1701859473
transform -1 0 1770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1069_
timestamp 1701859473
transform -1 0 2470 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1070_
timestamp 1701859473
transform 1 0 1810 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1071_
timestamp 1701859473
transform 1 0 2050 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1072_
timestamp 1701859473
transform 1 0 2210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1073_
timestamp 1701859473
transform 1 0 2010 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1074_
timestamp 1701859473
transform 1 0 1610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1075_
timestamp 1701859473
transform 1 0 1910 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1076_
timestamp 1701859473
transform 1 0 2330 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1077_
timestamp 1701859473
transform 1 0 2750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1078_
timestamp 1701859473
transform 1 0 3710 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1079_
timestamp 1701859473
transform 1 0 3750 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1080_
timestamp 1701859473
transform 1 0 2190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1081_
timestamp 1701859473
transform 1 0 2350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1082_
timestamp 1701859473
transform -1 0 2910 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1083_
timestamp 1701859473
transform 1 0 2450 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1084_
timestamp 1701859473
transform 1 0 2610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1085_
timestamp 1701859473
transform 1 0 3030 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1086_
timestamp 1701859473
transform 1 0 2830 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1087_
timestamp 1701859473
transform 1 0 2870 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1088_
timestamp 1701859473
transform -1 0 3950 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1089_
timestamp 1701859473
transform 1 0 3650 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1090_
timestamp 1701859473
transform 1 0 2690 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1091_
timestamp 1701859473
transform 1 0 2310 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1092_
timestamp 1701859473
transform -1 0 2990 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1093_
timestamp 1701859473
transform -1 0 2870 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1094_
timestamp 1701859473
transform 1 0 3790 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1095_
timestamp 1701859473
transform 1 0 4270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1096_
timestamp 1701859473
transform 1 0 4130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1097_
timestamp 1701859473
transform 1 0 1770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1098_
timestamp 1701859473
transform 1 0 3110 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1099_
timestamp 1701859473
transform 1 0 2730 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1100_
timestamp 1701859473
transform -1 0 2610 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1101_
timestamp 1701859473
transform -1 0 2490 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1102_
timestamp 1701859473
transform -1 0 2170 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1103_
timestamp 1701859473
transform 1 0 1810 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1104_
timestamp 1701859473
transform -1 0 510 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1105_
timestamp 1701859473
transform -1 0 2110 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1106_
timestamp 1701859473
transform -1 0 1970 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1107_
timestamp 1701859473
transform -1 0 1970 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1108_
timestamp 1701859473
transform -1 0 1450 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1109_
timestamp 1701859473
transform -1 0 1530 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1110_
timestamp 1701859473
transform -1 0 1290 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1111_
timestamp 1701859473
transform -1 0 1150 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1112_
timestamp 1701859473
transform -1 0 810 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1113_
timestamp 1701859473
transform -1 0 730 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1114_
timestamp 1701859473
transform 1 0 1390 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1115_
timestamp 1701859473
transform -1 0 1150 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1116_
timestamp 1701859473
transform -1 0 1290 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1117_
timestamp 1701859473
transform -1 0 1130 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1118_
timestamp 1701859473
transform -1 0 990 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1119_
timestamp 1701859473
transform -1 0 610 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1120_
timestamp 1701859473
transform -1 0 1170 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1121_
timestamp 1701859473
transform -1 0 1050 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1122_
timestamp 1701859473
transform -1 0 1050 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1123_
timestamp 1701859473
transform -1 0 770 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1124_
timestamp 1701859473
transform -1 0 610 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1125_
timestamp 1701859473
transform 1 0 890 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1126_
timestamp 1701859473
transform -1 0 350 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1127_
timestamp 1701859473
transform -1 0 630 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1128_
timestamp 1701859473
transform -1 0 350 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1129_
timestamp 1701859473
transform 1 0 1470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1130_
timestamp 1701859473
transform -1 0 1570 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1131_
timestamp 1701859473
transform -1 0 490 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1132_
timestamp 1701859473
transform 1 0 50 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1133_
timestamp 1701859473
transform -1 0 470 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1134_
timestamp 1701859473
transform -1 0 210 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2__1135_
timestamp 1701859473
transform 1 0 190 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1136_
timestamp 1701859473
transform 1 0 190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1137_
timestamp 1701859473
transform -1 0 350 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1138_
timestamp 1701859473
transform -1 0 70 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1139_
timestamp 1701859473
transform -1 0 70 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1140_
timestamp 1701859473
transform -1 0 210 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1141_
timestamp 1701859473
transform -1 0 350 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1142_
timestamp 1701859473
transform 1 0 50 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1143_
timestamp 1701859473
transform -1 0 70 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1144_
timestamp 1701859473
transform 1 0 190 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1145_
timestamp 1701859473
transform 1 0 410 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1146_
timestamp 1701859473
transform -1 0 1370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1147_
timestamp 1701859473
transform 1 0 1370 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1148_
timestamp 1701859473
transform 1 0 190 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1149_
timestamp 1701859473
transform -1 0 310 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1150_
timestamp 1701859473
transform -1 0 990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1151_
timestamp 1701859473
transform 1 0 690 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1152_
timestamp 1701859473
transform -1 0 770 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1153_
timestamp 1701859473
transform -1 0 1810 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1154_
timestamp 1701859473
transform 1 0 1530 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1155_
timestamp 1701859473
transform 1 0 1350 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1156_
timestamp 1701859473
transform -1 0 1410 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1157_
timestamp 1701859473
transform -1 0 1670 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1158_
timestamp 1701859473
transform -1 0 1270 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1159_
timestamp 1701859473
transform -1 0 1250 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1160_
timestamp 1701859473
transform 1 0 1310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1161_
timestamp 1701859473
transform 1 0 1490 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1162_
timestamp 1701859473
transform -1 0 1650 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1163_
timestamp 1701859473
transform -1 0 1030 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1164_
timestamp 1701859473
transform 1 0 870 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1165_
timestamp 1701859473
transform -1 0 870 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1166_
timestamp 1701859473
transform -1 0 950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1167_
timestamp 1701859473
transform -1 0 810 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1168_
timestamp 1701859473
transform 1 0 610 0 1 4950
box -12 -8 32 272
use FILL  FILL_2__1169_
timestamp 1701859473
transform -1 0 730 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1170_
timestamp 1701859473
transform -1 0 630 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1171_
timestamp 1701859473
transform 1 0 570 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1172_
timestamp 1701859473
transform -1 0 570 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1173_
timestamp 1701859473
transform -1 0 750 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1174_
timestamp 1701859473
transform 1 0 430 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2__1175_
timestamp 1701859473
transform -1 0 490 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1176_
timestamp 1701859473
transform -1 0 230 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1177_
timestamp 1701859473
transform 1 0 50 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1178_
timestamp 1701859473
transform -1 0 490 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1179_
timestamp 1701859473
transform -1 0 370 0 1 4430
box -12 -8 32 272
use FILL  FILL_2__1180_
timestamp 1701859473
transform -1 0 350 0 1 3910
box -12 -8 32 272
use FILL  FILL_2__1181_
timestamp 1701859473
transform -1 0 70 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1182_
timestamp 1701859473
transform -1 0 70 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1183_
timestamp 1701859473
transform -1 0 330 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1184_
timestamp 1701859473
transform 1 0 170 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1185_
timestamp 1701859473
transform 1 0 50 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1186_
timestamp 1701859473
transform -1 0 310 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1187_
timestamp 1701859473
transform 1 0 330 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1188_
timestamp 1701859473
transform 1 0 50 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1189_
timestamp 1701859473
transform -1 0 190 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1190_
timestamp 1701859473
transform 1 0 230 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1191_
timestamp 1701859473
transform 1 0 310 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1192_
timestamp 1701859473
transform -1 0 450 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1193_
timestamp 1701859473
transform -1 0 1090 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1194_
timestamp 1701859473
transform -1 0 1270 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1195_
timestamp 1701859473
transform -1 0 910 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2__1196_
timestamp 1701859473
transform -1 0 1790 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1197_
timestamp 1701859473
transform -1 0 1710 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1198_
timestamp 1701859473
transform -1 0 1590 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1199_
timestamp 1701859473
transform 1 0 1430 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1200_
timestamp 1701859473
transform -1 0 1130 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1201_
timestamp 1701859473
transform 1 0 970 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1202_
timestamp 1701859473
transform 1 0 830 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1203_
timestamp 1701859473
transform 1 0 1010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1204_
timestamp 1701859473
transform 1 0 1110 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1205_
timestamp 1701859473
transform -1 0 910 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1206_
timestamp 1701859473
transform -1 0 890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1207_
timestamp 1701859473
transform -1 0 750 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1208_
timestamp 1701859473
transform 1 0 590 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1209_
timestamp 1701859473
transform -1 0 470 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1210_
timestamp 1701859473
transform 1 0 190 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1211_
timestamp 1701859473
transform 1 0 410 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1212_
timestamp 1701859473
transform 1 0 2970 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1213_
timestamp 1701859473
transform -1 0 3530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1214_
timestamp 1701859473
transform 1 0 530 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1215_
timestamp 1701859473
transform -1 0 690 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1216_
timestamp 1701859473
transform -1 0 190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1217_
timestamp 1701859473
transform -1 0 290 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1218_
timestamp 1701859473
transform -1 0 310 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1219_
timestamp 1701859473
transform 1 0 170 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1220_
timestamp 1701859473
transform 1 0 290 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1221_
timestamp 1701859473
transform -1 0 1010 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1222_
timestamp 1701859473
transform 1 0 1530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1223_
timestamp 1701859473
transform 1 0 1350 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1224_
timestamp 1701859473
transform -1 0 1650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1225_
timestamp 1701859473
transform -1 0 1910 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1226_
timestamp 1701859473
transform -1 0 1950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1227_
timestamp 1701859473
transform -1 0 1670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1228_
timestamp 1701859473
transform -1 0 1550 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1229_
timestamp 1701859473
transform 1 0 1130 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1230_
timestamp 1701859473
transform -1 0 710 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1231_
timestamp 1701859473
transform 1 0 50 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1232_
timestamp 1701859473
transform -1 0 170 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1233_
timestamp 1701859473
transform -1 0 70 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1234_
timestamp 1701859473
transform 1 0 50 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1235_
timestamp 1701859473
transform -1 0 70 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1236_
timestamp 1701859473
transform -1 0 70 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1237_
timestamp 1701859473
transform -1 0 210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1238_
timestamp 1701859473
transform -1 0 1230 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1239_
timestamp 1701859473
transform 1 0 950 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1240_
timestamp 1701859473
transform -1 0 1110 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1241_
timestamp 1701859473
transform 1 0 450 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1242_
timestamp 1701859473
transform 1 0 810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1243_
timestamp 1701859473
transform 1 0 1310 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1244_
timestamp 1701859473
transform 1 0 1770 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1245_
timestamp 1701859473
transform 1 0 1790 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1246_
timestamp 1701859473
transform -1 0 1550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1247_
timestamp 1701859473
transform 1 0 1230 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1248_
timestamp 1701859473
transform -1 0 1110 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1249_
timestamp 1701859473
transform 1 0 690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1250_
timestamp 1701859473
transform -1 0 610 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1251_
timestamp 1701859473
transform 1 0 670 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1252_
timestamp 1701859473
transform 1 0 530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1253_
timestamp 1701859473
transform -1 0 590 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1254_
timestamp 1701859473
transform -1 0 450 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1255_
timestamp 1701859473
transform 1 0 530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1256_
timestamp 1701859473
transform 1 0 770 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1257_
timestamp 1701859473
transform 1 0 810 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1258_
timestamp 1701859473
transform -1 0 970 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1259_
timestamp 1701859473
transform -1 0 850 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1260_
timestamp 1701859473
transform 1 0 3430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1261_
timestamp 1701859473
transform -1 0 3430 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1262_
timestamp 1701859473
transform 1 0 3310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1263_
timestamp 1701859473
transform 1 0 3290 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1264_
timestamp 1701859473
transform -1 0 3210 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1265_
timestamp 1701859473
transform 1 0 3310 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1266_
timestamp 1701859473
transform 1 0 4290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1267_
timestamp 1701859473
transform 1 0 4030 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1268_
timestamp 1701859473
transform 1 0 4050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1269_
timestamp 1701859473
transform 1 0 3650 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1270_
timestamp 1701859473
transform 1 0 3530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1271_
timestamp 1701859473
transform -1 0 3790 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1272_
timestamp 1701859473
transform 1 0 3910 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1273_
timestamp 1701859473
transform -1 0 4350 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1274_
timestamp 1701859473
transform 1 0 4290 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1275_
timestamp 1701859473
transform -1 0 4170 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1276_
timestamp 1701859473
transform -1 0 5230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1277_
timestamp 1701859473
transform 1 0 5210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1278_
timestamp 1701859473
transform 1 0 5710 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1279_
timestamp 1701859473
transform 1 0 5690 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1280_
timestamp 1701859473
transform -1 0 4970 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1281_
timestamp 1701859473
transform 1 0 5070 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1282_
timestamp 1701859473
transform -1 0 5750 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1283_
timestamp 1701859473
transform -1 0 5650 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1284_
timestamp 1701859473
transform -1 0 5750 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1285_
timestamp 1701859473
transform 1 0 5530 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1286_
timestamp 1701859473
transform 1 0 5350 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1287_
timestamp 1701859473
transform -1 0 5570 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1288_
timestamp 1701859473
transform 1 0 4090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1289_
timestamp 1701859473
transform 1 0 5230 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1290_
timestamp 1701859473
transform 1 0 5350 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1291_
timestamp 1701859473
transform -1 0 5090 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1292_
timestamp 1701859473
transform 1 0 4950 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1293_
timestamp 1701859473
transform -1 0 5690 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1294_
timestamp 1701859473
transform -1 0 5550 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1295_
timestamp 1701859473
transform -1 0 5190 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1296_
timestamp 1701859473
transform 1 0 5050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1297_
timestamp 1701859473
transform 1 0 5270 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1298_
timestamp 1701859473
transform -1 0 5050 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1299_
timestamp 1701859473
transform -1 0 4230 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1300_
timestamp 1701859473
transform 1 0 5190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1301_
timestamp 1701859473
transform 1 0 5390 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1302_
timestamp 1701859473
transform 1 0 5330 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1303_
timestamp 1701859473
transform 1 0 5210 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1304_
timestamp 1701859473
transform -1 0 5230 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1305_
timestamp 1701859473
transform 1 0 5490 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1306_
timestamp 1701859473
transform 1 0 5610 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1307_
timestamp 1701859473
transform -1 0 5170 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1308_
timestamp 1701859473
transform 1 0 5250 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1309_
timestamp 1701859473
transform -1 0 5410 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1310_
timestamp 1701859473
transform -1 0 4510 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1311_
timestamp 1701859473
transform -1 0 4910 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1312_
timestamp 1701859473
transform 1 0 4270 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1313_
timestamp 1701859473
transform 1 0 4770 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1314_
timestamp 1701859473
transform 1 0 4630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1315_
timestamp 1701859473
transform -1 0 4710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1316_
timestamp 1701859473
transform -1 0 4570 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1317_
timestamp 1701859473
transform 1 0 3950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1318_
timestamp 1701859473
transform 1 0 4390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1319_
timestamp 1701859473
transform -1 0 4530 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1320_
timestamp 1701859473
transform 1 0 4630 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1321_
timestamp 1701859473
transform 1 0 4710 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1322_
timestamp 1701859473
transform 1 0 3990 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1323_
timestamp 1701859473
transform 1 0 4750 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1324_
timestamp 1701859473
transform 1 0 4610 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1325_
timestamp 1701859473
transform 1 0 2190 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1326_
timestamp 1701859473
transform -1 0 4950 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1327_
timestamp 1701859473
transform -1 0 4470 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1328_
timestamp 1701859473
transform 1 0 4570 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1329_
timestamp 1701859473
transform 1 0 4410 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1330_
timestamp 1701859473
transform -1 0 4650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1331_
timestamp 1701859473
transform -1 0 4850 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1332_
timestamp 1701859473
transform -1 0 4710 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1333_
timestamp 1701859473
transform 1 0 4570 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1334_
timestamp 1701859473
transform -1 0 1670 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1335_
timestamp 1701859473
transform -1 0 1810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1336_
timestamp 1701859473
transform 1 0 1630 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1337_
timestamp 1701859473
transform 1 0 1950 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1338_
timestamp 1701859473
transform 1 0 1890 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1339_
timestamp 1701859473
transform -1 0 1870 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1340_
timestamp 1701859473
transform -1 0 1770 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1341_
timestamp 1701859473
transform 1 0 2050 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1342_
timestamp 1701859473
transform -1 0 1630 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1343_
timestamp 1701859473
transform -1 0 1030 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1344_
timestamp 1701859473
transform -1 0 890 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1345_
timestamp 1701859473
transform 1 0 1130 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1346_
timestamp 1701859473
transform -1 0 1250 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1347_
timestamp 1701859473
transform 1 0 1290 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1348_
timestamp 1701859473
transform 1 0 1670 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1349_
timestamp 1701859473
transform -1 0 2470 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1350_
timestamp 1701859473
transform 1 0 2070 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1351_
timestamp 1701859473
transform -1 0 2710 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1352_
timestamp 1701859473
transform 1 0 1530 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1353_
timestamp 1701859473
transform -1 0 1370 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1354_
timestamp 1701859473
transform -1 0 1410 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1355_
timestamp 1701859473
transform -1 0 310 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1356_
timestamp 1701859473
transform -1 0 430 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1357_
timestamp 1701859473
transform 1 0 310 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1358_
timestamp 1701859473
transform 1 0 430 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1359_
timestamp 1701859473
transform 1 0 1890 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1360_
timestamp 1701859473
transform -1 0 1770 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1361_
timestamp 1701859473
transform 1 0 2310 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1362_
timestamp 1701859473
transform -1 0 1270 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1363_
timestamp 1701859473
transform 1 0 1130 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1364_
timestamp 1701859473
transform -1 0 790 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1365_
timestamp 1701859473
transform -1 0 670 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1366_
timestamp 1701859473
transform 1 0 650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1367_
timestamp 1701859473
transform -1 0 690 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1368_
timestamp 1701859473
transform -1 0 970 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1369_
timestamp 1701859473
transform -1 0 1530 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1370_
timestamp 1701859473
transform 1 0 1370 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1371_
timestamp 1701859473
transform 1 0 550 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1372_
timestamp 1701859473
transform -1 0 830 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1373_
timestamp 1701859473
transform -1 0 550 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1374_
timestamp 1701859473
transform 1 0 650 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1375_
timestamp 1701859473
transform -1 0 210 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1376_
timestamp 1701859473
transform 1 0 410 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1377_
timestamp 1701859473
transform -1 0 330 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1378_
timestamp 1701859473
transform -1 0 70 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1379_
timestamp 1701859473
transform 1 0 50 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1380_
timestamp 1701859473
transform 1 0 50 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1381_
timestamp 1701859473
transform 1 0 50 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1382_
timestamp 1701859473
transform 1 0 150 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1383_
timestamp 1701859473
transform 1 0 170 0 -1 790
box -12 -8 32 272
use FILL  FILL_2__1384_
timestamp 1701859473
transform 1 0 150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1385_
timestamp 1701859473
transform -1 0 890 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1386_
timestamp 1701859473
transform -1 0 910 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1387_
timestamp 1701859473
transform -1 0 790 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1388_
timestamp 1701859473
transform -1 0 570 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1389_
timestamp 1701859473
transform 1 0 310 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1390_
timestamp 1701859473
transform 1 0 470 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1391_
timestamp 1701859473
transform -1 0 630 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1392_
timestamp 1701859473
transform -1 0 430 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1393_
timestamp 1701859473
transform 1 0 410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1394_
timestamp 1701859473
transform -1 0 310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1395_
timestamp 1701859473
transform 1 0 510 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1396_
timestamp 1701859473
transform 1 0 890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1397_
timestamp 1701859473
transform -1 0 1010 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1398_
timestamp 1701859473
transform -1 0 1270 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1399_
timestamp 1701859473
transform -1 0 1110 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1400_
timestamp 1701859473
transform -1 0 1570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1401_
timestamp 1701859473
transform 1 0 1130 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1402_
timestamp 1701859473
transform 1 0 1270 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1403_
timestamp 1701859473
transform 1 0 1410 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1404_
timestamp 1701859473
transform 1 0 1390 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1405_
timestamp 1701859473
transform -1 0 3210 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1406_
timestamp 1701859473
transform 1 0 2470 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1407_
timestamp 1701859473
transform 1 0 2130 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1408_
timestamp 1701859473
transform -1 0 2270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1409_
timestamp 1701859473
transform 1 0 3470 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1410_
timestamp 1701859473
transform 1 0 2430 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1411_
timestamp 1701859473
transform -1 0 2570 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1412_
timestamp 1701859473
transform -1 0 3590 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1413_
timestamp 1701859473
transform 1 0 2090 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1414_
timestamp 1701859473
transform -1 0 2230 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1415_
timestamp 1701859473
transform -1 0 3750 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1416_
timestamp 1701859473
transform 1 0 2390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1417_
timestamp 1701859473
transform -1 0 2610 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1418_
timestamp 1701859473
transform 1 0 3230 0 1 270
box -12 -8 32 272
use FILL  FILL_2__1419_
timestamp 1701859473
transform 1 0 2150 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1420_
timestamp 1701859473
transform -1 0 2290 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1421_
timestamp 1701859473
transform 1 0 2230 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1422_
timestamp 1701859473
transform -1 0 2610 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1423_
timestamp 1701859473
transform -1 0 2750 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1424_
timestamp 1701859473
transform -1 0 3110 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1425_
timestamp 1701859473
transform 1 0 2410 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1426_
timestamp 1701859473
transform -1 0 2790 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1427_
timestamp 1701859473
transform 1 0 2750 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1428_
timestamp 1701859473
transform 1 0 3150 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1429_
timestamp 1701859473
transform 1 0 3290 0 1 1830
box -12 -8 32 272
use FILL  FILL_2__1430_
timestamp 1701859473
transform 1 0 3270 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1431_
timestamp 1701859473
transform -1 0 3410 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1432_
timestamp 1701859473
transform -1 0 3270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1433_
timestamp 1701859473
transform 1 0 3110 0 -1 2350
box -12 -8 32 272
use FILL  FILL_2__1434_
timestamp 1701859473
transform -1 0 3150 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1435_
timestamp 1701859473
transform 1 0 2970 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1436_
timestamp 1701859473
transform 1 0 2770 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1437_
timestamp 1701859473
transform -1 0 2650 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2__1438_
timestamp 1701859473
transform 1 0 2950 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1439_
timestamp 1701859473
transform 1 0 2810 0 -1 1310
box -12 -8 32 272
use FILL  FILL_2__1440_
timestamp 1701859473
transform -1 0 3890 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1441_
timestamp 1701859473
transform 1 0 3490 0 1 1310
box -12 -8 32 272
use FILL  FILL_2__1442_
timestamp 1701859473
transform 1 0 3530 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2__1443_
timestamp 1701859473
transform -1 0 3430 0 1 2350
box -12 -8 32 272
use FILL  FILL_2__1444_
timestamp 1701859473
transform -1 0 2490 0 1 3390
box -12 -8 32 272
use FILL  FILL_2__1445_
timestamp 1701859473
transform -1 0 2650 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1446_
timestamp 1701859473
transform -1 0 2890 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1447_
timestamp 1701859473
transform -1 0 3010 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1448_
timestamp 1701859473
transform -1 0 2430 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1449_
timestamp 1701859473
transform -1 0 2790 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1450_
timestamp 1701859473
transform -1 0 2030 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1451_
timestamp 1701859473
transform 1 0 1890 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1527_
timestamp 1701859473
transform 1 0 5710 0 1 790
box -12 -8 32 272
use FILL  FILL_2__1528_
timestamp 1701859473
transform -1 0 5730 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1529_
timestamp 1701859473
transform 1 0 5410 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2__1530_
timestamp 1701859473
transform 1 0 5150 0 1 2870
box -12 -8 32 272
use FILL  FILL_2__1531_
timestamp 1701859473
transform 1 0 2790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_2__1532_
timestamp 1701859473
transform 1 0 3830 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1533_
timestamp 1701859473
transform 1 0 4090 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1534_
timestamp 1701859473
transform 1 0 4210 0 -1 270
box -12 -8 32 272
use FILL  FILL_2__1535_
timestamp 1701859473
transform 1 0 3970 0 -1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert0
timestamp 1701859473
transform -1 0 1510 0 1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert1
timestamp 1701859473
transform 1 0 2170 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert2
timestamp 1701859473
transform 1 0 4810 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert3
timestamp 1701859473
transform 1 0 3690 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert4
timestamp 1701859473
transform 1 0 2170 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert5
timestamp 1701859473
transform 1 0 4170 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert6
timestamp 1701859473
transform -1 0 1390 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert15
timestamp 1701859473
transform -1 0 4770 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert16
timestamp 1701859473
transform -1 0 3550 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert17
timestamp 1701859473
transform -1 0 3990 0 -1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert18
timestamp 1701859473
transform 1 0 4930 0 -1 5470
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert19
timestamp 1701859473
transform -1 0 1650 0 1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert20
timestamp 1701859473
transform -1 0 4390 0 -1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert21
timestamp 1701859473
transform -1 0 1830 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert22
timestamp 1701859473
transform -1 0 4870 0 1 1830
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert23
timestamp 1701859473
transform -1 0 3090 0 -1 790
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert24
timestamp 1701859473
transform 1 0 5070 0 1 270
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert25
timestamp 1701859473
transform -1 0 3050 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert26
timestamp 1701859473
transform 1 0 3030 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert27
timestamp 1701859473
transform 1 0 3170 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert28
timestamp 1701859473
transform 1 0 2650 0 1 1310
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert29
timestamp 1701859473
transform -1 0 2530 0 -1 3390
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert30
timestamp 1701859473
transform -1 0 4370 0 -1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert31
timestamp 1701859473
transform -1 0 3510 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert32
timestamp 1701859473
transform 1 0 4630 0 1 4950
box -12 -8 32 272
use FILL  FILL_2_BUFX2_insert33
timestamp 1701859473
transform -1 0 4410 0 1 4430
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert7
timestamp 1701859473
transform -1 0 2810 0 -1 2870
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert8
timestamp 1701859473
transform -1 0 1630 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert9
timestamp 1701859473
transform -1 0 1770 0 -1 270
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert10
timestamp 1701859473
transform -1 0 2370 0 1 2350
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert11
timestamp 1701859473
transform 1 0 4290 0 1 790
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert12
timestamp 1701859473
transform -1 0 3250 0 -1 270
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert13
timestamp 1701859473
transform 1 0 2890 0 -1 1830
box -12 -8 32 272
use FILL  FILL_2_CLKBUF1_insert14
timestamp 1701859473
transform 1 0 4970 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__727_
timestamp 1701859473
transform 1 0 2930 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__735_
timestamp 1701859473
transform 1 0 4130 0 1 270
box -12 -8 32 272
use FILL  FILL_3__742_
timestamp 1701859473
transform -1 0 2970 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__750_
timestamp 1701859473
transform -1 0 3290 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__757_
timestamp 1701859473
transform 1 0 2530 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__765_
timestamp 1701859473
transform -1 0 2190 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__772_
timestamp 1701859473
transform -1 0 5450 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__780_
timestamp 1701859473
transform -1 0 4810 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__788_
timestamp 1701859473
transform -1 0 3590 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__795_
timestamp 1701859473
transform -1 0 1390 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__803_
timestamp 1701859473
transform -1 0 1270 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__810_
timestamp 1701859473
transform -1 0 1530 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__818_
timestamp 1701859473
transform -1 0 4130 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__825_
timestamp 1701859473
transform -1 0 4150 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__833_
timestamp 1701859473
transform -1 0 3170 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__841_
timestamp 1701859473
transform 1 0 4830 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__848_
timestamp 1701859473
transform 1 0 4370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__856_
timestamp 1701859473
transform 1 0 4490 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__863_
timestamp 1701859473
transform -1 0 2430 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__871_
timestamp 1701859473
transform 1 0 4330 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__878_
timestamp 1701859473
transform 1 0 5370 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__886_
timestamp 1701859473
transform 1 0 4250 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__894_
timestamp 1701859473
transform 1 0 5090 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__901_
timestamp 1701859473
transform 1 0 3250 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__909_
timestamp 1701859473
transform -1 0 5070 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__916_
timestamp 1701859473
transform 1 0 5590 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__924_
timestamp 1701859473
transform -1 0 2950 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__931_
timestamp 1701859473
transform 1 0 3250 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__939_
timestamp 1701859473
transform -1 0 5490 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__947_
timestamp 1701859473
transform 1 0 5630 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__954_
timestamp 1701859473
transform 1 0 5470 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__962_
timestamp 1701859473
transform 1 0 5590 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__969_
timestamp 1701859473
transform -1 0 5570 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__977_
timestamp 1701859473
transform -1 0 2930 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__984_
timestamp 1701859473
transform 1 0 2750 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__992_
timestamp 1701859473
transform 1 0 3350 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__999_
timestamp 1701859473
transform 1 0 3130 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1003_
timestamp 1701859473
transform 1 0 4790 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1011_
timestamp 1701859473
transform -1 0 4090 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1018_
timestamp 1701859473
transform -1 0 4130 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1026_
timestamp 1701859473
transform 1 0 5390 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1034_
timestamp 1701859473
transform -1 0 3790 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1041_
timestamp 1701859473
transform -1 0 2230 0 -1 4430
box -12 -8 32 272
use FILL  FILL_3__1049_
timestamp 1701859473
transform -1 0 2210 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1056_
timestamp 1701859473
transform 1 0 1310 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1064_
timestamp 1701859473
transform 1 0 1770 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1071_
timestamp 1701859473
transform 1 0 2070 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1079_
timestamp 1701859473
transform 1 0 3770 0 1 4950
box -12 -8 32 272
use FILL  FILL_3__1087_
timestamp 1701859473
transform 1 0 2890 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1094_
timestamp 1701859473
transform 1 0 3810 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1102_
timestamp 1701859473
transform -1 0 2190 0 -1 4950
box -12 -8 32 272
use FILL  FILL_3__1109_
timestamp 1701859473
transform -1 0 1550 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1117_
timestamp 1701859473
transform -1 0 1150 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1124_
timestamp 1701859473
transform -1 0 630 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1132_
timestamp 1701859473
transform 1 0 70 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3__1140_
timestamp 1701859473
transform -1 0 230 0 1 4430
box -12 -8 32 272
use FILL  FILL_3__1147_
timestamp 1701859473
transform 1 0 1390 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1155_
timestamp 1701859473
transform 1 0 1370 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1162_
timestamp 1701859473
transform -1 0 1670 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1170_
timestamp 1701859473
transform -1 0 650 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1177_
timestamp 1701859473
transform 1 0 70 0 1 3910
box -12 -8 32 272
use FILL  FILL_3__1185_
timestamp 1701859473
transform 1 0 70 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1193_
timestamp 1701859473
transform -1 0 1110 0 -1 3910
box -12 -8 32 272
use FILL  FILL_3__1200_
timestamp 1701859473
transform -1 0 1150 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1208_
timestamp 1701859473
transform 1 0 610 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1215_
timestamp 1701859473
transform -1 0 710 0 1 3390
box -12 -8 32 272
use FILL  FILL_3__1223_
timestamp 1701859473
transform 1 0 1370 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1230_
timestamp 1701859473
transform -1 0 730 0 1 2870
box -12 -8 32 272
use FILL  FILL_3__1238_
timestamp 1701859473
transform -1 0 1250 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1246_
timestamp 1701859473
transform -1 0 1570 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1253_
timestamp 1701859473
transform -1 0 610 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1261_
timestamp 1701859473
transform -1 0 3450 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1268_
timestamp 1701859473
transform 1 0 4070 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1276_
timestamp 1701859473
transform -1 0 5250 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1283_
timestamp 1701859473
transform -1 0 5670 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1291_
timestamp 1701859473
transform -1 0 5110 0 -1 1830
box -12 -8 32 272
use FILL  FILL_3__1299_
timestamp 1701859473
transform -1 0 4250 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1306_
timestamp 1701859473
transform 1 0 5630 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1314_
timestamp 1701859473
transform 1 0 4650 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1321_
timestamp 1701859473
transform 1 0 4730 0 1 1830
box -12 -8 32 272
use FILL  FILL_3__1329_
timestamp 1701859473
transform 1 0 4430 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1336_
timestamp 1701859473
transform 1 0 1650 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1344_
timestamp 1701859473
transform -1 0 910 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1352_
timestamp 1701859473
transform 1 0 1550 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1359_
timestamp 1701859473
transform 1 0 1910 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1367_
timestamp 1701859473
transform -1 0 710 0 -1 790
box -12 -8 32 272
use FILL  FILL_3__1374_
timestamp 1701859473
transform 1 0 670 0 1 270
box -12 -8 32 272
use FILL  FILL_3__1382_
timestamp 1701859473
transform 1 0 170 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1389_
timestamp 1701859473
transform 1 0 330 0 1 790
box -12 -8 32 272
use FILL  FILL_3__1397_
timestamp 1701859473
transform -1 0 1030 0 1 1310
box -12 -8 32 272
use FILL  FILL_3__1404_
timestamp 1701859473
transform 1 0 1410 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1412_
timestamp 1701859473
transform -1 0 3610 0 -1 270
box -12 -8 32 272
use FILL  FILL_3__1420_
timestamp 1701859473
transform -1 0 2310 0 -1 1310
box -12 -8 32 272
use FILL  FILL_3__1427_
timestamp 1701859473
transform 1 0 2770 0 -1 2350
box -12 -8 32 272
use FILL  FILL_3__1435_
timestamp 1701859473
transform 1 0 2990 0 1 2350
box -12 -8 32 272
use FILL  FILL_3__1442_
timestamp 1701859473
transform 1 0 3550 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3__1450_
timestamp 1701859473
transform -1 0 2050 0 -1 3390
box -12 -8 32 272
use FILL  FILL_3__1532_
timestamp 1701859473
transform 1 0 3850 0 -1 270
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert3
timestamp 1701859473
transform 1 0 3710 0 1 2350
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert18
timestamp 1701859473
transform 1 0 4950 0 -1 5470
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert26
timestamp 1701859473
transform 1 0 3050 0 -1 2870
box -12 -8 32 272
use FILL  FILL_3_BUFX2_insert33
timestamp 1701859473
transform -1 0 4430 0 1 4430
box -12 -8 32 272
use FILL  FILL_3_CLKBUF1_insert11
timestamp 1701859473
transform 1 0 4310 0 1 790
box -12 -8 32 272
<< labels >>
flabel metal1 s 5823 2 5883 2 3 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -63 2 -3 2 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 2957 5517 2963 5523 3 FreeSans 16 90 0 0 Cin[4]
port 3 nsew
flabel metal2 s 3037 5517 3043 5523 3 FreeSans 16 90 0 0 Cin[3]
port 4 nsew
flabel metal2 s 4657 5517 4663 5523 3 FreeSans 16 90 0 0 Cin[1]
port 6 nsew
flabel metal2 s 4937 5517 4943 5523 3 FreeSans 16 90 0 0 Cin[0]
port 7 nsew
flabel metal2 s 3757 -23 3763 -17 7 FreeSans 16 270 0 0 Yin[3]
port 18 nsew
flabel metal2 s 3217 -23 3223 -17 7 FreeSans 16 270 0 0 Yin[0]
port 21 nsew
flabel metal3 s -74 3276 -66 3284 7 FreeSans 16 0 0 0 Xin[1]
port 12 nsew
flabel metal3 s -74 3316 -66 3324 7 FreeSans 16 0 0 0 Xin[2]
port 11 nsew
flabel metal3 s -74 3236 -66 3244 7 FreeSans 16 0 0 0 Xin[3]
port 10 nsew
flabel metal3 s -74 3476 -66 3484 7 FreeSans 16 0 0 0 Rdy
port 8 nsew
flabel metal3 s -74 3516 -66 3524 7 FreeSans 16 0 0 0 Xin[0]
port 13 nsew
flabel metal2 s 2597 5517 2603 5523 3 FreeSans 16 90 0 0 Cin[5]
port 2 nsew
flabel metal2 s 3637 5517 3643 5523 3 FreeSans 16 90 0 0 Cin[2]
port 5 nsew
flabel metal2 s 4357 5516 4363 5522 3 FreeSans 16 90 0 0 clk
port 26 nsew
flabel metal3 s 5886 3896 5894 3904 3 FreeSans 16 0 0 0 Xout[3]
port 14 nsew
flabel metal3 s 5886 3176 5894 3184 3 FreeSans 16 0 0 0 Xout[2]
port 15 nsew
flabel metal3 s 5886 3236 5894 3244 3 FreeSans 16 0 0 0 Xout[1]
port 16 nsew
flabel metal3 s 5886 2996 5894 3004 3 FreeSans 16 0 0 0 Xout[0]
port 17 nsew
flabel metal3 s 5886 916 5894 924 3 FreeSans 16 0 0 0 Vld
port 9 nsew
flabel metal2 s 4037 -23 4043 -17 7 FreeSans 16 270 0 0 Yout[3]
port 22 nsew
flabel metal2 s 4157 -23 4163 -17 7 FreeSans 16 270 0 0 Yout[1]
port 24 nsew
flabel metal2 s 4277 -23 4283 -17 7 FreeSans 16 270 0 0 Yout[2]
port 23 nsew
flabel metal2 s 3917 -23 3923 -17 7 FreeSans 16 270 0 0 Yout[0]
port 25 nsew
flabel metal2 s 3657 -23 3663 -17 7 FreeSans 16 270 0 0 Yin[2]
port 19 nsew
flabel metal2 s 3457 -23 3463 -17 7 FreeSans 16 270 0 0 Yin[1]
port 20 nsew
<< properties >>
string FIXED_BBOX -40 -40 5860 5520
<< end >>
