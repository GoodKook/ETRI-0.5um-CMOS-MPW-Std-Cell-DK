* NGSPICE file created from fir_hls.ext - technology: scmos

.subckt OAI21X1 A B C Y vdd gnd
M1000 Y C a_7_14# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1001 a_30_146# A vdd vdd pfet w=12u l=0.6u
+  ad=3.6p pd=12.6u as=25.2p ps=28.2u
M1002 vdd C Y vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=14.4p ps=14.7u
M1003 gnd A a_7_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1004 Y B a_30_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.7u as=3.6p ps=12.6u
M1005 a_7_14# B gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
.ends

.subckt DFFPOSX1 D CLK Q vdd gnd
M1000 vdd Q a_189_206# vdd pfet w=3u l=0.6u
+  ad=10.125p pd=14.7u as=0.9p ps=3.6u
M1001 a_83_186# a_11_14# a_59_14# vdd pfet w=6u l=0.6u
+  ad=3.6p pd=7.2u as=7.2p ps=8.4u
M1002 a_87_10# a_59_14# gnd gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=4.05p ps=5.7u
M1003 gnd CLK a_11_14# gnd nfet w=6u l=0.6u
+  ad=5.85p pd=8.4u as=12.6p ps=16.2u
M1004 gnd a_87_10# a_81_14# gnd nfet w=3u l=0.6u
+  ad=4.05p pd=5.7u as=1.35p ps=3.9u
M1005 a_159_14# a_87_10# gnd gnd nfet w=3u l=0.6u
+  ad=0.9p pd=3.6u as=6.3p ps=10.2u
M1006 a_49_186# D vdd vdd pfet w=6u l=0.6u
+  ad=4.5p pd=7.5u as=11.25p ps=14.4u
M1007 vdd a_87_10# a_83_186# vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=3.6p ps=7.2u
M1008 Q a_167_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=6.975p ps=8.7u
M1009 Q a_167_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=10.125p ps=14.7u
M1010 a_167_14# CLK a_159_14# gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=0.9p ps=3.6u
M1011 a_49_14# D gnd gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=5.85p ps=8.4u
M1012 a_87_10# a_59_14# vdd vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1013 a_59_14# CLK a_49_186# vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=4.5p ps=7.5u
M1014 a_161_186# a_87_10# vdd vdd pfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=12.6p ps=16.2u
M1015 a_189_206# CLK a_167_14# vdd pfet w=3u l=0.6u
+  ad=0.9p pd=3.6u as=6.075p ps=8.4u
M1016 a_59_14# a_11_14# a_49_14# gnd nfet w=3u l=0.6u
+  ad=4.05p pd=5.7u as=1.35p ps=3.9u
M1017 a_187_14# a_11_14# a_167_14# gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=3.6p ps=5.4u
M1018 vdd CLK a_11_14# vdd pfet w=12u l=0.6u
+  ad=11.25p pd=14.4u as=25.2p ps=28.2u
M1019 gnd Q a_187_14# gnd nfet w=3u l=0.6u
+  ad=6.975p pd=8.7u as=1.35p ps=3.9u
M1020 a_167_14# a_11_14# a_161_186# vdd pfet w=6u l=0.6u
+  ad=6.075p pd=8.4u as=1.8p ps=6.6u
M1021 a_81_14# CLK a_59_14# gnd nfet w=3u l=0.6u
+  ad=1.35p pd=3.9u as=4.05p ps=5.7u
.ends

.subckt INVX1 A Y vdd gnd
M1000 Y A gnd gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=6.3p ps=10.2u
M1001 Y A vdd vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=12.6p ps=16.2u
.ends

.subckt NAND2X1 A B Y vdd gnd
M1000 a_27_14# A gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.6p ps=16.2u
M1001 Y B a_27_14# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=2.7p ps=6.9u
M1002 vdd B Y vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1003 Y A vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
.ends

.subckt NOR2X1 A B Y vdd gnd
M1000 a_25_146# A vdd vdd pfet w=12u l=0.6u
+  ad=3.6p pd=12.6u as=25.2p ps=28.2u
M1001 Y A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1002 Y B a_25_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=3.6p ps=12.6u
M1003 gnd B Y gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
.ends

.subckt OR2X2 A B Y vdd gnd
M1000 Y a_7_146# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=6.3p ps=8.4u
M1001 a_25_146# A a_7_146# vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=25.2p ps=28.2u
M1002 a_7_146# A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=6.3p ps=10.2u
M1003 Y a_7_146# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1004 gnd B a_7_146# gnd nfet w=3u l=0.6u
+  ad=6.3p pd=8.4u as=3.6p ps=5.4u
M1005 vdd B a_25_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=5.4p ps=12.9u
.ends

.subckt NAND3X1 A B C Y vdd gnd
M1000 Y C a_34_14# gnd nfet w=9u l=0.6u
+  ad=18.9p pd=22.2u as=2.7p ps=9.6u
M1001 a_26_14# A gnd gnd nfet w=9u l=0.6u
+  ad=2.7p pd=9.6u as=18.9p ps=22.2u
M1002 vdd B Y vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1003 a_34_14# B a_26_14# gnd nfet w=9u l=0.6u
+  ad=2.7p pd=9.6u as=2.7p ps=9.6u
M1004 Y C vdd vdd pfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1005 Y A vdd vdd pfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
.ends

.subckt MUX2X1 A B S Y vdd gnd
M1000 a_75_22# S Y gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=7.2p ps=8.4u
M1001 gnd S a_7_22# gnd nfet w=3u l=0.6u
+  ad=6.3p pd=8.4u as=6.3p ps=10.2u
M1002 Y S a_45_138# vdd pfet w=12u l=0.6u
+  ad=14.49p pd=15.6u as=5.4p ps=12.9u
M1003 gnd A a_75_22# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=2.7p ps=6.9u
M1004 vdd A a_75_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=5.4p ps=12.9u
M1005 a_45_138# B vdd vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=11.7p ps=14.4u
M1006 a_45_22# B gnd gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=6.3p ps=8.4u
M1007 Y a_7_22# a_45_22# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=2.7p ps=6.9u
M1008 a_75_146# a_7_22# Y vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=14.49p ps=15.6u
M1009 vdd S a_7_22# vdd pfet w=6u l=0.6u
+  ad=11.7p pd=14.4u as=12.6p ps=16.2u
.ends

.subckt OAI22X1 A B C D Y vdd gnd
M1000 Y D a_7_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1001 a_25_146# A vdd vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=25.2p ps=28.2u
M1002 a_65_146# D Y vdd pfet w=12u l=0.6u
+  ad=5.4p pd=12.9u as=23.4p ps=15.9u
M1003 gnd A a_7_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1004 a_7_14# C Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1005 a_7_14# B gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1006 Y B a_25_146# vdd pfet w=12u l=0.6u
+  ad=23.4p pd=15.9u as=5.4p ps=12.9u
M1007 vdd C a_65_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=5.4p ps=12.9u
.ends

.subckt AOI21X1 A B C Y vdd gnd
M1000 vdd A a_7_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1001 Y C a_7_146# vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1002 a_28_14# A gnd gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=12.6p ps=16.2u
M1003 Y B a_28_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.7u as=1.8p ps=6.6u
M1004 a_7_146# B vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1005 gnd C Y gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=7.2p ps=8.7u
.ends

.subckt AOI22X1 A B C D Y vdd gnd
M1000 gnd C a_56_14# gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=1.8p ps=6.6u
M1001 vdd A a_7_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1002 Y D a_7_146# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1003 a_28_14# A gnd gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=12.6p ps=16.2u
M1004 Y B a_28_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=1.8p ps=6.6u
M1005 a_7_146# C Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1006 a_7_146# B vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1007 a_56_14# D Y gnd nfet w=6u l=0.6u
+  ad=1.8p pd=6.6u as=7.2p ps=8.4u
.ends

.subckt INVX4 A Y vdd gnd
M1000 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1001 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1002 gnd A Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1003 vdd A Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
.ends

.subckt AND2X2 A B Y vdd gnd
M1000 a_25_14# A a_7_14# gnd nfet w=6u l=0.6u
+  ad=2.7p pd=6.9u as=12.6p ps=16.2u
M1001 gnd B a_25_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=2.7p ps=6.9u
M1002 vdd B a_7_14# vdd pfet w=6u l=0.6u
+  ad=14.4p pd=14.7u as=8.1p ps=8.7u
M1003 Y a_7_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1004 Y a_7_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.7u
M1005 a_7_14# A vdd vdd pfet w=6u l=0.6u
+  ad=8.1p pd=8.7u as=12.6p ps=16.2u
.ends

.subckt INVX2 A Y vdd gnd
M1000 Y A vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=25.2p ps=28.2u
M1001 Y A gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=12.6p ps=16.2u
.ends

.subckt CLKBUF1 A Y vdd gnd
M1000 Y a_105_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1001 a_65_14# a_25_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1002 a_105_14# a_65_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1003 Y a_105_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1004 a_25_14# A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1005 a_65_14# a_25_14# vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1006 a_25_14# A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1007 gnd a_25_14# a_65_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1008 a_105_14# a_65_14# gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1009 gnd a_105_14# Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1010 vdd a_65_14# a_105_14# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1011 vdd a_105_14# Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1012 vdd a_25_14# a_65_14# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1013 gnd A a_25_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1014 vdd A a_25_14# vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1015 gnd a_65_14# a_105_14# gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
.ends

.subckt BUFX2 A Y vdd gnd
M1000 Y a_7_14# vdd vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.7u
M1001 gnd A a_7_14# gnd nfet w=3u l=0.6u
+  ad=7.2p pd=8.7u as=6.3p ps=10.2u
M1002 Y a_7_14# gnd gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.7u
M1003 vdd A a_7_14# vdd pfet w=6u l=0.6u
+  ad=14.4p pd=14.7u as=12.6p ps=16.2u
.ends

.subckt NOR3X1 A B C Y vdd gnd
M1000 gnd B Y gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=3.6p ps=5.4u
M1001 a_7_166# A vdd vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=10.8p ps=11.4u
M1002 a_7_166# B a_65_166# vdd pfet w=9u l=0.6u
+  ad=18.9p pd=22.2u as=10.8p ps=11.4u
M1003 a_65_166# C Y vdd pfet w=9u l=0.6u
+  ad=18.9p pd=22.2u as=10.8p ps=11.4u
M1004 Y C gnd gnd nfet w=3u l=0.6u
+  ad=6.3p pd=10.2u as=3.6p ps=5.4u
M1005 a_65_166# B a_7_166# vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=10.8p ps=11.4u
M1006 vdd A a_7_166# vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=18.9p ps=22.2u
M1007 Y C a_65_166# vdd pfet w=9u l=0.6u
+  ad=10.8p pd=11.4u as=18.9p ps=22.2u
M1008 Y A gnd gnd nfet w=3u l=0.6u
+  ad=3.6p pd=5.4u as=7.2p ps=10.8u
.ends

.subckt INVX8 A Y vdd gnd
M1000 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1001 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=25.2p ps=28.2u
M1002 Y A vdd vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
M1003 Y A gnd gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=12.6p ps=16.2u
M1004 gnd A Y gnd nfet w=6u l=0.6u
+  ad=12.6p pd=16.2u as=7.2p ps=8.4u
M1005 vdd A Y vdd pfet w=12u l=0.6u
+  ad=25.2p pd=28.2u as=14.4p ps=14.4u
M1006 gnd A Y gnd nfet w=6u l=0.6u
+  ad=7.2p pd=8.4u as=7.2p ps=8.4u
M1007 vdd A Y vdd pfet w=12u l=0.6u
+  ad=14.4p pd=14.4u as=14.4p ps=14.4u
.ends

.subckt fir_hls gnd vdd clk ready rst x[7] x[6] x[5] x[4] x[3] x[2] x[1] x[0] y[7]
+ y[6] y[5] y[4] y[3] y[2] y[1] y[0]
X_2037_ _2045_/A _2045_/B _2044_/A _2051_/B vdd gnd OAI21X1
X_2106_ _2106_/A _2106_/B _2106_/C _2169_/A vdd gnd OAI21X1
X_3086_ _3086_/D _3099_/CLK _3086_/Q vdd gnd DFFPOSX1
X_2939_ _3090_/Q _2950_/B vdd gnd INVX1
X_1606_ _1690_/Q _1630_/B _1658_/A vdd gnd NAND2X1
X_2655_ _2665_/A _2655_/B _2656_/C vdd gnd NOR2X1
X_2724_ _3033_/Q _2740_/B _2726_/D vdd gnd NOR2X1
X_1468_ _1468_/A _1692_/Q _1469_/A vdd gnd OR2X2
X_1537_ _1559_/Q _1555_/B _1537_/C _1545_/A vdd gnd NAND3X1
X_2586_ _3062_/Q _3094_/Q _2633_/S _2588_/B vdd gnd MUX2X1
X_3069_ _3069_/D _3101_/CLK _3069_/Q vdd gnd DFFPOSX1
X_2440_ _2440_/D _2535_/CLK _2440_/Q vdd gnd DFFPOSX1
X_2371_ _2386_/A _2371_/B _2385_/A _2375_/C vdd gnd OAI21X1
X_2569_ _3034_/Q _2581_/B _2571_/C vdd gnd NOR2X1
X_2638_ _3075_/Q _3059_/Q _2638_/S _2640_/B vdd gnd MUX2X1
X_2707_ _2957_/S _2707_/B _2890_/A _2860_/A vdd gnd NAND3X1
X_1871_ _2291_/B vdd _1871_/C _2445_/D vdd gnd OAI21X1
X_1940_ _1940_/A _1940_/B _1940_/C _1999_/C vdd gnd NAND3X1
X_2423_ _2423_/A _2424_/C vdd gnd INVX1
X_2285_ _2293_/A _2294_/A _2294_/B _2286_/A vdd gnd OAI21X1
X_2354_ _2364_/A _2363_/A _2355_/A vdd gnd NOR2X1
X_2070_ _2070_/A _2206_/B _2071_/A _2233_/B _2073_/C vdd gnd OAI22X1
X_2972_ _2984_/A _2972_/B _2972_/C _2973_/B vdd gnd OAI21X1
X_1785_ _2442_/Q _2268_/B vdd gnd INVX1
X_1854_ _1916_/A _1861_/C _1860_/C _1988_/A vdd gnd NAND3X1
X_1923_ _1928_/A _1989_/B _1989_/A _1926_/A vdd gnd AOI21X1
X_2406_ _2406_/A _2412_/C _2412_/A vdd gnd NOR2X1
X_2199_ _2375_/B vdd _2199_/C _2199_/D _2451_/D vdd gnd OAI22X1
X_2268_ _2268_/A _2268_/B _2268_/C _2278_/A vdd gnd OAI21X1
X_2337_ _2350_/A _2349_/A _2338_/A vdd gnd NOR2X1
X_1570_ _1570_/D _3061_/CLK _3020_/A vdd gnd DFFPOSX1
X_2053_ _2061_/A _2062_/C _2117_/B vdd gnd NAND2X1
X_2122_ _2122_/A _2146_/C _2156_/A vdd gnd NAND2X1
X_2955_ _2955_/A _2979_/B _2986_/A _2962_/D vdd gnd AOI21X1
X_1768_ vdd _3089_/Q _1769_/C vdd gnd NAND2X1
X_1837_ _1845_/A _1841_/B vdd gnd INVX1
X_1906_ _1906_/A _1974_/C _1932_/A vdd gnd NAND2X1
X_2886_ _3085_/Q _2889_/A vdd gnd INVX1
X_1699_ _1699_/D _3095_/CLK _1699_/Q vdd gnd DFFPOSX1
X_1622_ _1631_/A _2467_/Q _1663_/B vdd gnd NAND2X1
X_2671_ _2783_/A _2985_/D _2985_/A vdd gnd NOR2X1
X_2740_ _3037_/Q _2740_/B _2742_/D vdd gnd NOR2X1
X_1484_ _1484_/A _1484_/B _1484_/C _3110_/A vdd gnd NAND3X1
X_1553_ _1681_/D _1554_/B vdd gnd INVX1
X_2036_ _2040_/C _2069_/C _2040_/B _2045_/B vdd gnd AOI21X1
X_2105_ _2108_/C _2154_/C _2108_/A _2106_/A vdd gnd AOI21X1
X_3085_ _3085_/D _3101_/CLK _3085_/Q vdd gnd DFFPOSX1
X_2938_ _2986_/A _2938_/B _2938_/C _2938_/D _3089_/D vdd gnd AOI22X1
X_2869_ _3032_/Q _2888_/C _2870_/A vdd gnd NAND2X1
X_2723_ _3049_/Q _2726_/A vdd gnd INVX1
X_1536_ vdd _1536_/B _1552_/B vdd gnd NAND2X1
X_1605_ _1657_/B _1657_/A _2318_/A vdd gnd NAND2X1
X_2585_ _3030_/Q _2665_/A _2593_/C vdd gnd NAND2X1
X_2654_ _2885_/A _2879_/B _2988_/A _2654_/D _2655_/B vdd gnd OAI22X1
X_1467_ _1468_/A _1467_/B _1481_/B _1481_/A _3105_/A vdd gnd AOI22X1
X_2019_ _2025_/A _2204_/A _2125_/A _2030_/B vdd gnd OAI21X1
X_3068_ _3068_/D _3101_/CLK _3068_/Q vdd gnd DFFPOSX1
X_2370_ _2370_/A _2384_/B _2385_/A vdd gnd NOR2X1
X_2706_ _2706_/A _2706_/B _2706_/C _2819_/B vdd gnd NAND3X1
X_1519_ _1519_/A x[6] _1520_/C vdd gnd NAND2X1
X_2499_ _2518_/Q _2499_/B _2499_/Y vdd gnd NOR2X1
X_2568_ _3026_/Q _2571_/A vdd gnd INVX1
X_2637_ _3035_/Q _2646_/B vdd gnd INVX1
X_1870_ vdd _1870_/B _1870_/C _1871_/C vdd gnd NAND3X1
X_2353_ _2353_/A _2450_/Q _2364_/A vdd gnd NOR2X1
X_2422_ _2422_/A _2423_/A _2422_/C _2425_/A vdd gnd NAND3X1
X_2284_ _2284_/A _2284_/B _2286_/B vdd gnd NAND2X1
X_1999_ _1999_/A _2066_/A _1999_/C _2050_/A vdd gnd OAI21X1
X_1922_ _1988_/C _1988_/D _1922_/C _1989_/B vdd gnd NAND3X1
X_2971_ _2984_/A _3052_/Q _2972_/C vdd gnd NAND2X1
X_1784_ _2255_/B vdd _1784_/C _2441_/D vdd gnd OAI21X1
X_1853_ _1931_/C _1853_/B _1853_/C _1861_/C vdd gnd OAI21X1
X_2336_ _2336_/A _2449_/Q _2350_/A vdd gnd NOR2X1
X_2405_ _2405_/A _2454_/Q _2406_/A vdd gnd NOR2X1
X_2198_ _2230_/B _2198_/B vdd _2199_/C vdd gnd OAI21X1
X_2267_ _2311_/B _2267_/B _2267_/C _2456_/D vdd gnd OAI21X1
X_2052_ _2052_/A _2107_/B _2052_/C _2061_/A vdd gnd NAND3X1
X_2121_ _2450_/Q _2352_/B vdd gnd INVX1
X_1905_ _1968_/A _1969_/A _1969_/B _1979_/A vdd gnd NAND3X1
X_2954_ _2960_/A _2954_/B _2954_/C _2955_/A vdd gnd OAI21X1
X_2885_ _2885_/A _2889_/B _2885_/C _2885_/D _3084_/D vdd gnd OAI22X1
X_1698_ _1698_/D _2470_/CLK _1698_/Q vdd gnd DFFPOSX1
X_1767_ _2436_/Q _2080_/A vdd gnd INVX1
X_1836_ _2427_/Q _2437_/Q _1845_/A vdd gnd NAND2X1
X_2319_ _2319_/A _2324_/A _2341_/A vdd gnd OR2X2
X_1552_ _1552_/A _1552_/B rst _1561_/D vdd gnd AOI21X1
X_1621_ _1695_/Q _1630_/B _1663_/A vdd gnd NAND2X1
X_2670_ _2708_/B _2988_/B _2991_/B _2712_/B _2704_/B vdd gnd OAI22X1
X_1483_ _1696_/Q _1483_/B _1483_/C _1484_/C vdd gnd NAND3X1
X_2104_ _2104_/A _2104_/B _2104_/C _2108_/C vdd gnd OAI21X1
X_2035_ _2035_/A _2035_/B _2035_/C _2040_/C vdd gnd OAI21X1
X_3084_ _3084_/D _3101_/CLK _3084_/Q vdd gnd DFFPOSX1
X_2937_ _2985_/A _2937_/B _2937_/C _2985_/D _2938_/C vdd gnd AOI22X1
X_2868_ _3080_/Q _2887_/B _2876_/C _2870_/C vdd gnd NAND3X1
X_1819_ _1834_/C _1822_/C _1820_/C vdd gnd NAND2X1
X_2799_ _3065_/Q _2802_/A vdd gnd INVX1
X_2722_ _2722_/A _2742_/B _2722_/C _2722_/D _3048_/D vdd gnd OAI22X1
X_1535_ _1535_/A _1545_/B vdd gnd INVX1
X_1604_ _1604_/A _2461_/Q _1657_/B vdd gnd NAND2X1
X_2584_ _2706_/C _2665_/A vdd gnd INVX4
X_2653_ _3068_/Q _3100_/Q _2661_/S _2654_/D vdd gnd MUX2X1
X_1466_ _1691_/Q _1466_/B _1467_/B vdd gnd NAND2X1
X_3067_ _3067_/D _3099_/CLK _3067_/Q vdd gnd DFFPOSX1
X_2018_ _2431_/Q _2436_/Q _2125_/A vdd gnd AND2X2
X_2636_ _2665_/A _2636_/B _2636_/C _2636_/D _3034_/D vdd gnd AOI22X1
X_2705_ _3046_/Q _2714_/A vdd gnd INVX1
X_1449_ _1693_/Q _1477_/B _1465_/B _1451_/C vdd gnd OAI21X1
X_1518_ _3016_/A _1520_/B vdd gnd INVX1
X_2498_ _2519_/Q _2499_/B vdd gnd INVX1
X_2567_ _2622_/C _2583_/B _2567_/C _2567_/D _3025_/D vdd gnd OAI22X1
X_2283_ _2294_/A _2293_/A _2284_/A vdd gnd NOR2X1
X_2352_ _2352_/A _2352_/B _2363_/A vdd gnd NOR2X1
X_2421_ _2470_/Q _2426_/A _2426_/C vdd gnd NAND2X1
X_1998_ _2011_/C _2066_/A vdd gnd INVX1
X_2619_ _3049_/Q _3041_/Q _2638_/S _2620_/A vdd gnd MUX2X1
X_1852_ _1908_/A _1931_/C vdd gnd INVX1
X_1921_ _1930_/A _1921_/B _1921_/C _1988_/D vdd gnd NAND3X1
X_2970_ _2970_/A _2970_/B _2982_/S _2973_/C vdd gnd MUX2X1
X_1783_ _2427_/Q _2433_/Q vdd _1784_/C vdd gnd NAND3X1
X_2266_ _2456_/Q _2311_/B _2267_/C vdd gnd NAND2X1
X_2335_ _2335_/A _2335_/B _2349_/A vdd gnd NOR2X1
X_2404_ _2405_/A _2454_/Q _2412_/C vdd gnd AND2X2
X_2197_ _2198_/B _2230_/B _2199_/D vdd gnd AND2X2
X_2120_ _2335_/B vdd _2120_/C _2120_/D _2449_/D vdd gnd OAI22X1
X_2051_ _2051_/A _2051_/B _2051_/C _2052_/C vdd gnd NAND3X1
X_1835_ _1861_/A _1860_/C vdd gnd INVX1
X_1904_ _1907_/A _1907_/B _1908_/A _1969_/B vdd gnd OAI21X1
X_2953_ _2960_/A _3075_/Q _2954_/C vdd gnd NAND2X1
X_2884_ _2888_/A _3016_/A _2888_/C _2885_/D vdd gnd AOI21X1
X_1697_ _1697_/D _2469_/CLK _1697_/Q vdd gnd DFFPOSX1
X_1766_ vdd _2025_/A _1766_/C _2435_/D vdd gnd OAI21X1
X_2249_ _2249_/A _2249_/B _2250_/B vdd gnd NOR2X1
X_2318_ _2318_/A _2447_/Q _2324_/A vdd gnd NOR2X1
X_1482_ _1695_/Q _1482_/B _1482_/C _1484_/A vdd gnd OAI21X1
X_1551_ _2533_/B _1551_/B _1552_/A vdd gnd NAND2X1
X_1620_ _1662_/B _1662_/A _2377_/A vdd gnd NAND2X1
X_2103_ _2110_/C _2110_/A _2110_/B _2154_/C vdd gnd NAND3X1
X_3083_ _3083_/D _3099_/CLK _3083_/Q vdd gnd DFFPOSX1
X_2034_ _2068_/A _2068_/B _2068_/C _2069_/C vdd gnd NAND3X1
X_1818_ _1818_/A _1818_/B _1818_/C _1822_/C vdd gnd NAND3X1
X_2936_ _2948_/A _2936_/B _2936_/C _2937_/B vdd gnd OAI21X1
X_2867_ _3000_/A _2887_/B _2888_/A _2870_/B vdd gnd NAND3X1
X_2798_ _2798_/A _2818_/B _2798_/C _2798_/D _3064_/D vdd gnd OAI22X1
X_1749_ _2430_/Q _2179_/A vdd gnd INVX2
X_2652_ _3084_/Q _2885_/A vdd gnd INVX1
X_2721_ _3000_/A _2741_/B _2742_/B _2722_/C vdd gnd OAI21X1
X_1465_ _1474_/A _1465_/B _1465_/C _1481_/B vdd gnd AOI21X1
X_1534_ _1543_/B _1547_/B _1539_/B vdd gnd NAND2X1
X_1603_ _1689_/Q _1630_/B _1657_/A vdd gnd NAND2X1
X_2583_ _2662_/C _2583_/B _2583_/C _2583_/D _3029_/D vdd gnd OAI22X1
X_2017_ _2430_/Q _2437_/Q _2075_/A vdd gnd NAND2X1
X_3066_ _3066_/D _3098_/CLK _3066_/Q vdd gnd DFFPOSX1
X_2919_ _2919_/A _2979_/B _2986_/A _2926_/D vdd gnd AOI21X1
X_2635_ _2665_/A _2635_/B _2636_/C vdd gnd NOR2X1
X_2704_ _2984_/B _2704_/B _2704_/C _2704_/D _3045_/D vdd gnd OAI22X1
X_1448_ _1448_/A _1448_/B _1465_/B vdd gnd AND2X2
X_1517_ _1517_/A _1517_/B _1517_/C _1568_/D vdd gnd OAI21X1
X_2497_ _2511_/B _2512_/B _2497_/Y vdd gnd NOR2X1
X_2566_ _3004_/A _2582_/B _2583_/B _2567_/D vdd gnd OAI21X1
X_3049_ _3049_/D _3098_/CLK _3049_/Q vdd gnd DFFPOSX1
X_2420_ _2420_/A _2420_/B _2420_/C _2469_/D vdd gnd OAI21X1
X_2282_ _2282_/A _2444_/Q _2294_/A vdd gnd NOR2X1
X_2351_ _2353_/A _2352_/A vdd gnd INVX1
X_1997_ _2429_/Q _2438_/Q _2011_/C vdd gnd AND2X2
X_2549_ _2707_/B _2890_/A _2550_/B vdd gnd NAND2X1
X_2618_ _3073_/Q _3057_/Q _2638_/S _2620_/B vdd gnd MUX2X1
X_1851_ _1851_/A _2028_/A _1908_/A vdd gnd NAND2X1
X_1920_ _1980_/A _1980_/C _1930_/B _1988_/C vdd gnd NAND3X1
X_1782_ _2441_/Q _2255_/B vdd gnd INVX1
X_2403_ _2403_/A _2415_/B _2403_/C _2409_/A vdd gnd OAI21X1
X_2196_ _2196_/A _2229_/A _2230_/B vdd gnd NAND2X1
X_2265_ _2265_/A _2268_/C _2267_/B vdd gnd NAND2X1
X_2334_ _2336_/A _2335_/A vdd gnd INVX1
X_2050_ _2050_/A _2107_/A _2050_/C _2107_/B vdd gnd NAND3X1
XCLKBUF1_insert10 clk _3097_/CLK vdd gnd CLKBUF1
X_2952_ _3059_/Q _2954_/B vdd gnd INVX1
X_1765_ vdd _3088_/Q _1766_/C vdd gnd NAND2X1
X_1834_ _1834_/A _1876_/A _1834_/C _1859_/A vdd gnd OAI21X1
X_1903_ _2435_/Q _2430_/Q _1946_/C _1958_/C _1907_/B vdd gnd AOI22X1
X_2883_ _3036_/Q _2887_/B _2885_/C vdd gnd NOR2X1
X_1696_ _1696_/D _2470_/CLK _1696_/Q vdd gnd DFFPOSX1
X_2179_ _2179_/A _2206_/B _2203_/A vdd gnd NOR2X1
X_2248_ _2248_/A _2248_/B vdd _2249_/A vdd gnd OAI21X1
X_2317_ _2339_/A _2319_/A vdd gnd INVX1
X_1481_ _1481_/A _1481_/B _1481_/C _1481_/D _3109_/A vdd gnd AOI22X1
X_1550_ _2481_/Y _1551_/B vdd gnd INVX1
X_2033_ _2033_/A _2066_/C _2040_/B vdd gnd AND2X2
X_2102_ _2102_/A _2102_/B _2154_/A _2106_/B vdd gnd AOI21X1
X_3082_ _3082_/D _3097_/CLK _3082_/Q vdd gnd DFFPOSX1
X_2935_ _2948_/A _3049_/Q _2936_/C vdd gnd NAND2X1
X_1748_ vdd _2071_/A _1748_/C _2429_/D vdd gnd OAI21X1
X_1817_ _2070_/A _2025_/A _1817_/C _1818_/C vdd gnd OAI21X1
X_2866_ _2866_/A _2866_/B _2866_/C _3079_/D vdd gnd NAND3X1
X_2797_ _3000_/A _2817_/B _2818_/B _2798_/C vdd gnd OAI21X1
X_1679_ _1679_/D _3075_/CLK _1679_/Q vdd gnd DFFPOSX1
X_1602_ _1656_/B _1656_/A _2305_/A vdd gnd NAND2X1
X_2582_ _3020_/A _2582_/B _2583_/B _2583_/D vdd gnd OAI21X1
X_2651_ _3028_/Q _2651_/B _2651_/C _2743_/A _2656_/D vdd gnd AOI22X1
X_2720_ _3032_/Q _2740_/B _2722_/D vdd gnd NOR2X1
X_1464_ _1464_/A _1465_/C vdd gnd INVX1
X_1533_ _1537_/C _1535_/A _1533_/C _1547_/B vdd gnd NAND3X1
X_2016_ _2016_/A _2016_/B _2016_/C _2068_/C vdd gnd OAI21X1
X_3065_ _3065_/D _3097_/CLK _3065_/Q vdd gnd DFFPOSX1
X_2918_ _2945_/S _2918_/B _2918_/C _2919_/A vdd gnd OAI21X1
X_2849_ _3016_/A _2853_/B _2853_/C _2850_/A vdd gnd OAI21X1
X_1516_ _1517_/A x[5] _1517_/C vdd gnd NAND2X1
X_2565_ _3033_/Q _2581_/B _2567_/C vdd gnd NOR2X1
X_2634_ _2634_/A _2879_/B _2988_/A _2634_/D _2635_/B vdd gnd OAI22X1
X_2703_ _3020_/A _2703_/B _2704_/B _2704_/D vdd gnd OAI21X1
X_1447_ _1697_/Q _1482_/C _1448_/B vdd gnd NOR2X1
X_2496_ _2507_/B _2512_/B vdd gnd INVX1
X_3048_ _3048_/D _3075_/CLK _3048_/Q vdd gnd DFFPOSX1
X_2281_ _2281_/A _2281_/B _2293_/A vdd gnd NOR2X1
X_2350_ _2350_/A _2389_/B _2364_/B _2357_/A vdd gnd OAI21X1
X_1996_ _1996_/A _1996_/B _1996_/C _2047_/C vdd gnd AOI21X1
X_2548_ _2785_/A _2783_/A _2856_/A vdd gnd NOR2X1
X_2617_ _3033_/Q _2626_/B vdd gnd INVX1
X_2479_ _2511_/C _2509_/B vdd gnd INVX1
X_1781_ vdd _2206_/B _1781_/C _2440_/D vdd gnd OAI21X1
X_1850_ _1856_/B _1876_/C _1853_/C vdd gnd NAND2X1
X_2333_ _2463_/Q _2382_/A _2347_/C vdd gnd NAND2X1
X_2402_ _2412_/B _2403_/C vdd gnd INVX1
X_2195_ _2195_/A _2214_/A _2195_/C _2229_/A vdd gnd NAND3X1
X_2264_ _2264_/A _2264_/B _2264_/C _2265_/A vdd gnd OAI21X1
X_1979_ _1979_/A _1979_/B _1979_/C _1980_/B vdd gnd AOI21X1
X_1902_ _1902_/A _1902_/B _1946_/A _1907_/A vdd gnd AOI21X1
XCLKBUF1_insert11 clk _3087_/CLK vdd gnd CLKBUF1
X_2951_ _3091_/Q _2962_/B vdd gnd INVX1
X_1764_ _2435_/Q _2025_/A vdd gnd INVX2
X_1833_ _2429_/Q _2435_/Q _1876_/A vdd gnd NAND2X1
X_2882_ _2882_/A _2889_/B _2882_/C _2882_/D _3083_/D vdd gnd OAI22X1
X_1695_ _1695_/D _2470_/CLK _1695_/Q vdd gnd DFFPOSX1
X_2316_ _2318_/A _2447_/Q _2339_/A vdd gnd NAND2X1
X_2178_ _2179_/A _2206_/B _2178_/C _2186_/A vdd gnd OAI21X1
X_2247_ _2247_/A _2249_/B vdd gnd INVX1
X_1480_ _1695_/Q _1482_/B _1481_/D vdd gnd NAND2X1
X_2032_ _2041_/C _2041_/B _2069_/A _2045_/A vdd gnd AOI21X1
X_2101_ _2110_/A _2110_/B _2104_/C _2102_/B vdd gnd NAND3X1
X_3081_ _3081_/D _3097_/CLK _3081_/Q vdd gnd DFFPOSX1
X_2934_ _2934_/A _2934_/B _2982_/S _2937_/C vdd gnd MUX2X1
X_2865_ _3031_/Q _2888_/C _2866_/A vdd gnd NAND2X1
X_1678_ _1678_/D _3075_/CLK _1678_/Q vdd gnd DFFPOSX1
X_1747_ vdd _1747_/B _1748_/C vdd gnd NAND2X1
X_1816_ _1816_/A _2071_/A _1839_/A _1818_/B vdd gnd OAI21X1
X_2796_ _3032_/Q _2816_/B _2798_/D vdd gnd NOR2X1
X_1532_ _1559_/Q _1555_/B _1533_/C vdd gnd NOR2X1
X_1601_ _1607_/A _2460_/Q _1656_/B vdd gnd NAND2X1
X_2581_ _3037_/Q _2581_/B _2583_/C vdd gnd NOR2X1
X_2650_ _2650_/A _2650_/B _2667_/B _2651_/C vdd gnd MUX2X1
X_1463_ _1479_/B _1479_/A _1474_/A vdd gnd NAND2X1
X_2015_ _2015_/A _2015_/B _2016_/B vdd gnd AND2X2
X_3064_ _3064_/D _3099_/CLK _3064_/Q vdd gnd DFFPOSX1
X_2917_ _2945_/S _3072_/Q _2918_/C vdd gnd NAND2X1
X_2848_ _3036_/Q _2852_/B _2850_/B vdd gnd NOR2X1
X_2779_ _3037_/Q _2779_/B _2781_/A vdd gnd NOR2X1
X_2702_ _3037_/Q _2702_/B _2704_/C vdd gnd NOR2X1
X_1515_ _3012_/A _1517_/B vdd gnd INVX1
X_2495_ _2495_/A _2511_/C _2511_/B _2743_/A vdd gnd MUX2X1
X_2564_ _3025_/Q _2622_/C vdd gnd INVX1
X_2633_ _3066_/Q _3098_/Q _2633_/S _2634_/D vdd gnd MUX2X1
X_1446_ _1696_/Q _1482_/C vdd gnd INVX1
X_3047_ _3047_/D _3095_/CLK _3047_/Q vdd gnd DFFPOSX1
X_2280_ _2282_/A _2281_/A vdd gnd INVX1
X_1995_ _2049_/C _1996_/C vdd gnd INVX1
X_2616_ _2665_/A _2616_/B _2616_/C _2616_/D _3032_/D vdd gnd AOI22X1
X_2478_ _2524_/Q _2493_/A _2511_/C vdd gnd NAND2X1
X_2547_ _2860_/B _2991_/B _2879_/A _2662_/D _2583_/B vdd gnd OAI22X1
X_1780_ vdd _3093_/Q _1781_/C vdd gnd NAND2X1
X_2332_ _2332_/A _2332_/B _2332_/C _2332_/D _2462_/D vdd gnd AOI22X1
X_2401_ _2468_/Q _2410_/B vdd gnd INVX1
X_2194_ _2194_/A _2194_/B _2195_/C vdd gnd NAND2X1
X_2263_ _2263_/A _2263_/B _2268_/C vdd gnd NAND2X1
X_1978_ _1978_/A _1978_/B _1978_/C _1985_/B vdd gnd OAI21X1
X_1832_ _1832_/A _1864_/A vdd gnd INVX1
X_1901_ _1931_/C _1931_/B _1931_/A _1968_/A vdd gnd NAND3X1
XCLKBUF1_insert12 clk _3101_/CLK vdd gnd CLKBUF1
X_2950_ _2986_/A _2950_/B _2950_/C _2950_/D _3090_/D vdd gnd AOI22X1
X_2881_ _2888_/A _3012_/A _2888_/C _2882_/D vdd gnd AOI21X1
X_1694_ _1694_/D _2470_/CLK _1694_/Q vdd gnd DFFPOSX1
X_1763_ vdd _1816_/A _1763_/C _2434_/D vdd gnd OAI21X1
X_2246_ _2454_/Q _2251_/A vdd gnd INVX1
X_2315_ _2343_/C _2343_/A _2342_/B _2324_/B vdd gnd AOI21X1
X_2177_ _2180_/A _2206_/C _2203_/B _2178_/C vdd gnd OAI21X1
X_2100_ _2124_/A _2100_/B _2100_/C _2110_/B vdd gnd NAND3X1
X_3080_ _3080_/D _3097_/CLK _3080_/Q vdd gnd DFFPOSX1
X_2031_ _2068_/A _2035_/C _2068_/B _2041_/B vdd gnd NAND3X1
X_1815_ _1815_/A _1815_/B _1815_/C _1834_/C vdd gnd NAND3X1
X_2933_ _3081_/Q _3025_/Q _2945_/S _2934_/A vdd gnd MUX2X1
X_2864_ _3079_/Q _2887_/B _2876_/C _2866_/C vdd gnd NAND3X1
X_2795_ _3064_/Q _2798_/A vdd gnd INVX1
X_1677_ _1677_/D _3075_/CLK _1677_/Q vdd gnd DFFPOSX1
X_1746_ _2429_/Q _2071_/A vdd gnd INVX2
X_2229_ _2229_/A _2230_/A _2229_/C _2231_/C vdd gnd OAI21X1
X_1462_ _1691_/Q _1692_/Q _1693_/Q _1479_/B vdd gnd AOI21X1
X_1531_ _1558_/Q _1555_/B vdd gnd INVX1
X_1600_ _1688_/Q _1630_/B _1656_/A vdd gnd NAND2X1
X_2580_ _3029_/Q _2662_/C vdd gnd INVX1
X_3063_ _3063_/D _3095_/CLK _3063_/Q vdd gnd DFFPOSX1
X_2014_ _2435_/Q _2431_/Q _2015_/B vdd gnd NAND2X1
X_2916_ _3056_/Q _2918_/B vdd gnd INVX1
X_2847_ _3076_/Q _2851_/B _2850_/C vdd gnd NAND2X1
X_2778_ _3061_/Q _2779_/B _2778_/C _2781_/C vdd gnd NAND3X1
X_1729_ _1736_/A _1735_/B vdd gnd INVX1
X_2632_ _3082_/Q _2634_/A vdd gnd INVX1
X_2701_ _3045_/Q _2984_/B vdd gnd INVX1
X_1445_ _1695_/Q _1479_/C _1448_/A vdd gnd NOR2X1
X_1514_ _1522_/A _1514_/B _1514_/C _1567_/D vdd gnd OAI21X1
X_2494_ _2508_/C _2495_/A vdd gnd INVX1
X_2563_ _2563_/A _2583_/B _2563_/C _2563_/D _3024_/D vdd gnd OAI22X1
X_3046_ _3046_/D _3075_/CLK _3046_/Q vdd gnd DFFPOSX1
X_1994_ _2062_/A _2056_/B _2054_/B vdd gnd NOR2X1
X_2615_ _2665_/A _2615_/B _2616_/C vdd gnd NOR2X1
X_2477_ _2493_/A _2524_/Q _2511_/A _2507_/B vdd gnd AOI21X1
X_2546_ _2707_/B _2890_/A _2546_/C _2991_/B vdd gnd NAND3X1
X_3029_ _3029_/D _3101_/CLK _3029_/Q vdd gnd DFFPOSX1
X_2400_ _2400_/A _2400_/B _2400_/C _2467_/D vdd gnd OAI21X1
X_2262_ _2264_/B _2264_/A _2263_/B vdd gnd NOR2X1
X_2331_ _2331_/A _2340_/A _2332_/A _2332_/C vdd gnd AOI21X1
X_2193_ _2194_/A _2194_/B _2193_/C _2196_/A vdd gnd NAND3X1
X_1977_ _1996_/B _2049_/C _1996_/A _1978_/B vdd gnd AOI21X1
X_2529_ _2535_/Q _2533_/A vdd gnd INVX1
X_1831_ _2445_/Q _2291_/B vdd gnd INVX1
X_1900_ _1946_/A _1902_/A _1902_/B _1931_/B vdd gnd NAND3X1
X_2880_ _3035_/Q _2887_/B _2882_/C vdd gnd NOR2X1
X_1693_ _1693_/D _2470_/CLK _1693_/Q vdd gnd DFFPOSX1
X_1762_ vdd _3087_/Q _1763_/C vdd gnd NAND2X1
X_2176_ _2204_/A _2176_/B _2248_/A _2203_/B vdd gnd OAI21X1
X_2245_ _2245_/A _2245_/B _2453_/D vdd gnd NAND2X1
X_2314_ _2314_/A _2314_/B _2343_/A vdd gnd AND2X2
X_2030_ _2075_/A _2030_/B _2030_/C _2068_/B vdd gnd NAND3X1
X_2932_ _3065_/Q _3097_/Q _2945_/S _2934_/B vdd gnd MUX2X1
X_1745_ vdd _2070_/A _1745_/C _2428_/D vdd gnd OAI21X1
X_1814_ _2070_/A _2025_/A _1814_/C _1815_/A vdd gnd OAI21X1
X_2863_ _2996_/A _2887_/B _2888_/A _2866_/B vdd gnd NAND3X1
X_2794_ _2794_/A _2818_/B _2794_/C _2794_/D _3063_/D vdd gnd OAI22X1
X_1676_ _1676_/D _3075_/CLK _1676_/Q vdd gnd DFFPOSX1
X_2159_ _2160_/B _2171_/A _2169_/C _2166_/A vdd gnd AOI21X1
X_2228_ _2453_/Q _2382_/A _2245_/A vdd gnd NAND2X1
X_1461_ _1461_/A _1461_/B _1461_/C _1479_/A vdd gnd NAND3X1
X_1530_ _1536_/B _1557_/Q _1535_/A vdd gnd NOR2X1
X_2013_ _2066_/C _2033_/A _2069_/A vdd gnd NAND2X1
X_3062_ _3062_/D _3099_/CLK _3062_/Q vdd gnd DFFPOSX1
X_2915_ _3088_/Q _2926_/B vdd gnd INVX1
X_1728_ _1728_/D _2535_/CLK _1750_/B vdd gnd DFFPOSX1
X_2846_ _2846_/A _2846_/B _2846_/C _3075_/D vdd gnd OAI21X1
X_2777_ _2777_/A _2777_/B _2777_/C _3060_/D vdd gnd OAI21X1
X_1659_ _1659_/A _1659_/B _1665_/C _1691_/D vdd gnd AOI21X1
X_2562_ _3000_/A _2582_/B _2583_/B _2563_/D vdd gnd OAI21X1
X_2631_ _3026_/Q _2651_/B _2631_/C _2743_/A _2636_/D vdd gnd AOI22X1
X_2700_ _2972_/B _2704_/B _2700_/C _2700_/D _3044_/D vdd gnd OAI22X1
X_1444_ _1694_/Q _1479_/C vdd gnd INVX1
X_1513_ _1522_/A x[4] _1514_/C vdd gnd NAND2X1
X_2493_ _2493_/A _2508_/A _2502_/A _2493_/D _2508_/C vdd gnd AOI22X1
X_3045_ _3045_/D _3093_/CLK _3045_/Q vdd gnd DFFPOSX1
X_2829_ _2996_/A _2853_/B _2853_/C _2830_/A vdd gnd OAI21X1
X_1993_ _2117_/A _2117_/C _2056_/B vdd gnd NOR2X1
X_2545_ _2957_/S _2546_/C vdd gnd INVX1
X_2614_ _2614_/A _2879_/B _2988_/A _2614_/D _2615_/B vdd gnd OAI22X1
X_2476_ _2533_/B _2511_/A vdd gnd INVX2
X_3028_ _3028_/D _3101_/CLK _3028_/Q vdd gnd DFFPOSX1
X_2192_ _2195_/A _2214_/A _2193_/C vdd gnd NAND2X1
X_2261_ _2261_/A _2442_/Q _2264_/B vdd gnd NOR2X1
X_2330_ _2339_/B _2330_/B _2340_/A vdd gnd NOR2X1
X_1976_ _1976_/A _1976_/B _1976_/C _1996_/B vdd gnd OAI21X1
X_2528_ _2531_/B _2531_/A _2528_/Y vdd gnd NAND2X1
X_2459_ _2459_/D _2469_/CLK _2459_/Q vdd gnd DFFPOSX1
X_1761_ _2434_/Q _1816_/A vdd gnd INVX1
X_1830_ _2281_/B vdd _1830_/C _1830_/D _2444_/D vdd gnd OAI22X1
X_1692_ _1692_/D _2469_/CLK _1692_/Q vdd gnd DFFPOSX1
X_2313_ _2313_/A _2313_/B _2313_/C _2342_/B vdd gnd OAI21X1
X_2175_ _2431_/Q _2439_/Q _2248_/A vdd gnd NAND2X1
X_2244_ vdd _2244_/B _2251_/C _2245_/B vdd gnd NAND3X1
X_1959_ _2028_/C _2028_/D _2016_/C _2001_/B vdd gnd NAND3X1
X_2931_ _2931_/A _2979_/B _2986_/A _2938_/D vdd gnd AOI21X1
X_1744_ vdd _1756_/B _1745_/C vdd gnd NAND2X1
X_1813_ _1817_/C _1839_/A _1815_/C vdd gnd NAND2X1
X_2862_ _2862_/A _2862_/B _2862_/C _3078_/D vdd gnd NAND3X1
X_2793_ _2996_/A _2817_/B _2818_/B _2794_/C vdd gnd OAI21X1
X_1675_ _1736_/A _1675_/B _1703_/D vdd gnd AND2X2
X_2089_ _2125_/C _2125_/D _2089_/C _2123_/B vdd gnd NAND3X1
X_2158_ _2158_/A _2158_/B _2169_/C vdd gnd NOR2X1
X_2227_ _2227_/A _2227_/B _2452_/D vdd gnd NAND2X1
X_1460_ _1693_/Q _1460_/B _1461_/B vdd gnd NOR2X1
X_2012_ _2012_/A _2012_/B _2012_/C _2033_/A vdd gnd NAND3X1
X_3061_ _3061_/D _3061_/CLK _3061_/Q vdd gnd DFFPOSX1
X_2914_ _2986_/A _2914_/B _2914_/C _2914_/D _3087_/D vdd gnd AOI22X1
X_2845_ _3012_/A _2853_/B _2853_/C _2846_/A vdd gnd OAI21X1
X_1658_ _1658_/A _1658_/B _1658_/C _1690_/D vdd gnd AOI21X1
X_1727_ _1727_/D _3087_/CLK _1747_/B vdd gnd DFFPOSX1
X_2776_ _2780_/A _3016_/A _2780_/C _2777_/B vdd gnd AOI21X1
X_1589_ _1604_/A _2456_/Q _1652_/B vdd gnd NAND2X1
X_1512_ _3008_/A _1514_/B vdd gnd INVX1
X_2492_ _2522_/Q _2493_/D vdd gnd INVX1
X_2561_ _3032_/Q _2581_/B _2563_/C vdd gnd NOR2X1
X_2630_ _2630_/A _2630_/B _2667_/B _2631_/C vdd gnd MUX2X1
X_1443_ _1457_/B _1457_/A _1460_/B _1477_/B vdd gnd AOI21X1
X_3044_ _3044_/D _3093_/CLK _3044_/Q vdd gnd DFFPOSX1
X_2828_ _3031_/Q _2852_/B _2830_/B vdd gnd NOR2X1
X_2759_ _3032_/Q _2779_/B _2761_/A vdd gnd NOR2X1
X_1992_ _1992_/A _2062_/A vdd gnd INVX1
X_2475_ _2493_/A _2508_/A _2517_/D vdd gnd NAND2X1
X_2544_ _2985_/D _2982_/S _2860_/B vdd gnd NAND2X1
X_2613_ _3064_/Q _3096_/Q _2643_/S _2614_/D vdd gnd MUX2X1
X_3027_ _3027_/D _3099_/CLK _3027_/Q vdd gnd DFFPOSX1
X_2191_ _2212_/A _2191_/B _2191_/C _2214_/A vdd gnd NAND3X1
X_2260_ _2268_/A _2268_/B _2264_/A vdd gnd NOR2X1
X_1975_ _2048_/C _2048_/A _2048_/B _2049_/C vdd gnd NAND3X1
X_2458_ _2458_/D _2462_/CLK _2458_/Q vdd gnd DFFPOSX1
X_2527_ _2534_/Q _2530_/A _2531_/A vdd gnd NAND2X1
X_2389_ _2389_/A _2389_/B _2390_/B vdd gnd NOR2X1
X_1691_ _1691_/D _2470_/CLK _1691_/Q vdd gnd DFFPOSX1
X_1760_ vdd _1895_/A _1760_/C _2433_/D vdd gnd OAI21X1
XCLKBUF1_insert0 clk _3098_/CLK vdd gnd CLKBUF1
X_2312_ _2312_/A _2313_/B vdd gnd INVX1
X_2174_ _2432_/Q _2439_/Q _2206_/C vdd gnd NAND2X1
X_2243_ _2243_/A _2243_/B _2251_/C vdd gnd NAND2X1
X_1889_ _2435_/Q _2430_/Q _1946_/A vdd gnd NAND2X1
X_1958_ _1958_/A _1958_/B _1958_/C _1958_/D _1965_/C vdd gnd AOI22X1
X_2930_ _2948_/A _2930_/B _2930_/C _2931_/A vdd gnd OAI21X1
X_2861_ _3030_/Q _2888_/C _2862_/A vdd gnd NAND2X1
X_1674_ vdd rst _1675_/B vdd gnd NOR2X1
X_1743_ _2428_/Q _2070_/A vdd gnd INVX2
X_1812_ _2428_/Q _2435_/Q _1839_/A vdd gnd AND2X2
X_2792_ _3031_/Q _2816_/B _2794_/D vdd gnd NOR2X1
X_2226_ vdd _2226_/B _2226_/C _2227_/B vdd gnd NAND3X1
X_2088_ _2088_/A _2088_/B _2088_/C _2095_/C vdd gnd AOI21X1
X_2157_ _2161_/C _2194_/B _2162_/A _2158_/B vdd gnd AOI21X1
X_3060_ _3060_/D _3101_/CLK _3060_/Q vdd gnd DFFPOSX1
X_2011_ _2070_/A _2233_/B _2011_/C _2012_/C vdd gnd OAI21X1
X_2913_ _2985_/A _2913_/B _2913_/C _2985_/D _2914_/C vdd gnd AOI22X1
X_2844_ _3035_/Q _2852_/B _2846_/B vdd gnd NOR2X1
X_1588_ _1684_/Q _1630_/B _1652_/A vdd gnd NAND2X1
X_1657_ _1657_/A _1657_/B _1658_/C _1689_/D vdd gnd AOI21X1
X_1726_ _1726_/D _2535_/CLK _1756_/B vdd gnd DFFPOSX1
X_2775_ _3036_/Q _2779_/B _2777_/A vdd gnd NOR2X1
X_2209_ _2234_/A _2234_/B _2210_/A vdd gnd NAND2X1
X_1442_ _1690_/Q _1452_/A _1442_/C _1457_/B vdd gnd NAND3X1
X_1511_ _1517_/A _1511_/B _1511_/C _1566_/D vdd gnd OAI21X1
X_2491_ _2491_/A _2505_/A _2491_/C _2511_/C _2743_/B vdd gnd AOI22X1
X_2560_ _3024_/Q _2563_/A vdd gnd INVX1
X_3043_ _3043_/D _3075_/CLK _3043_/Q vdd gnd DFFPOSX1
X_2758_ _3056_/Q _2779_/B _2778_/C _2761_/C vdd gnd NAND3X1
X_2827_ _3071_/Q _2851_/B _2830_/C vdd gnd NAND2X1
X_1709_ _1715_/A _1723_/A vdd gnd INVX1
X_2689_ _3042_/Q _2948_/B vdd gnd INVX1
X_1991_ _1991_/A _1991_/B _1991_/C _2447_/D vdd gnd OAI21X1
X_2612_ _3080_/Q _2614_/A vdd gnd INVX1
X_2474_ _2523_/Q _2508_/A vdd gnd INVX1
X_2543_ _2783_/A _2982_/S vdd gnd INVX4
X_3026_ _3026_/D _3098_/CLK _3026_/Q vdd gnd DFFPOSX1
X_2190_ _2190_/A _2190_/B _2191_/C vdd gnd NAND2X1
X_1974_ _1974_/A _1974_/B _1974_/C _1996_/A vdd gnd OAI21X1
X_2388_ _2388_/A _2388_/B _2389_/A vdd gnd NAND2X1
X_2457_ _2457_/D _2462_/CLK _2457_/Q vdd gnd DFFPOSX1
X_2526_ _2533_/B _2530_/A vdd gnd INVX1
X_3009_ _3009_/A _3021_/B _3009_/C _3009_/D _3098_/D vdd gnd OAI22X1
X_1690_ _1690_/D _2462_/CLK _1690_/Q vdd gnd DFFPOSX1
XCLKBUF1_insert1 clk _3075_/CLK vdd gnd CLKBUF1
X_2242_ _2242_/A _2243_/A vdd gnd INVX1
X_2311_ _2461_/Q _2311_/B _2322_/C vdd gnd NAND2X1
X_2173_ _2173_/A _2180_/A _2185_/A vdd gnd NOR2X1
X_1957_ _1965_/A _1965_/B _2001_/C _1971_/C vdd gnd OAI21X1
X_1888_ _1974_/C _1906_/A _1969_/A vdd gnd AND2X2
X_2509_ _2511_/A _2509_/B _2517_/D _2510_/C vdd gnd OAI21X1
X_1811_ _2434_/Q _2429_/Q _1817_/C vdd gnd AND2X2
X_2860_ _2860_/A _2860_/B _2888_/C vdd gnd NOR2X1
X_2791_ _3063_/Q _2794_/A vdd gnd INVX1
X_1673_ rst _1673_/B _1702_/D vdd gnd NOR2X1
X_1742_ vdd _1800_/A _1742_/C _2427_/D vdd gnd OAI21X1
X_2225_ _2225_/A _2225_/B _2225_/C _2226_/C vdd gnd OAI21X1
X_2087_ _2087_/A _2125_/A _2088_/C vdd gnd AND2X2
X_2156_ _2156_/A _2156_/B _2156_/C _2161_/C vdd gnd NAND3X1
X_2989_ _2989_/A _2989_/B _3019_/B vdd gnd NAND2X1
X_2010_ _2071_/A _2176_/B _2122_/A _2012_/B vdd gnd OAI21X1
X_2912_ _2957_/S _2912_/B _2912_/C _2913_/B vdd gnd OAI21X1
X_1725_ _1725_/D _3087_/CLK _1753_/B vdd gnd DFFPOSX1
X_2843_ _3075_/Q _2851_/B _2846_/C vdd gnd NAND2X1
X_2774_ _3060_/Q _2779_/B _2778_/C _2777_/C vdd gnd NAND3X1
X_1587_ _1651_/B _1651_/A _2252_/A vdd gnd NAND2X1
X_1656_ _1656_/A _1656_/B _1658_/C _1688_/D vdd gnd AOI21X1
X_2139_ _2185_/B _2139_/B _2139_/C _2145_/B vdd gnd OAI21X1
X_2208_ _2234_/B _2234_/A _2235_/A vdd gnd OR2X2
X_1441_ _1688_/Q _1689_/Q _1442_/C vdd gnd AND2X2
X_1510_ _1517_/A x[3] _1511_/C vdd gnd NAND2X1
X_2490_ _2522_/Q _2521_/Q _2530_/Y _2505_/A vdd gnd AOI21X1
X_3042_ _3042_/D _3075_/CLK _3042_/Q vdd gnd DFFPOSX1
X_1708_ _1715_/A _1720_/A _1720_/B _1711_/B vdd gnd OAI21X1
X_2688_ _2936_/B _2704_/B _2688_/C _2688_/D _3041_/D vdd gnd OAI22X1
X_2757_ _2757_/A _2757_/B _2757_/C _3055_/D vdd gnd OAI21X1
X_2826_ _2826_/A _2826_/B _2826_/C _3070_/D vdd gnd OAI21X1
X_1639_ _1639_/A _1639_/B _1676_/D vdd gnd NAND2X1
X_1990_ _2117_/A _2117_/C vdd _1991_/A vdd gnd OAI21X1
X_2542_ _2785_/A _2985_/D vdd gnd INVX4
X_2611_ _3024_/Q _2651_/B _2611_/C _2743_/A _2616_/D vdd gnd AOI22X1
X_2473_ _2530_/Y _2493_/A vdd gnd INVX1
X_3025_ _3025_/D _3097_/CLK _3025_/Q vdd gnd DFFPOSX1
X_2809_ _3012_/A _2817_/B _2818_/B _2810_/C vdd gnd OAI21X1
X_1973_ _1973_/A _1974_/C _1983_/C _1983_/B _1978_/A vdd gnd AOI22X1
X_2525_ _2532_/A _2531_/B vdd gnd INVX1
X_2387_ _2387_/A _2387_/B _2390_/A vdd gnd NAND2X1
X_2456_ _2456_/D _2462_/CLK _2456_/Q vdd gnd DFFPOSX1
X_3008_ _3008_/A _3020_/B _3021_/B _3009_/D vdd gnd OAI21X1
XCLKBUF1_insert2 clk _3099_/CLK vdd gnd CLKBUF1
X_2172_ _2231_/B _2202_/B _2198_/B vdd gnd NOR2X1
X_2241_ _2241_/A _2241_/B _2243_/B vdd gnd NAND2X1
X_2310_ vdd _2310_/B _2310_/C _2460_/D vdd gnd OAI21X1
X_1887_ _1887_/A _1887_/B _1887_/C _1906_/A vdd gnd NAND3X1
X_1956_ _2016_/C _2028_/C _2028_/D _1965_/A vdd gnd AOI21X1
X_2508_ _2508_/A _2508_/B _2508_/C _2510_/B vdd gnd AOI21X1
X_2439_ _2439_/D _2535_/CLK _2439_/Q vdd gnd DFFPOSX1
X_1741_ _1753_/B vdd _1742_/C vdd gnd NAND2X1
X_1810_ _1818_/A _1815_/B vdd gnd INVX1
X_2790_ _2790_/A _2818_/B _2790_/C _2790_/D _3062_/D vdd gnd OAI22X1
X_1672_ rst _1672_/B _1701_/D vdd gnd NOR2X1
X_2155_ _2155_/A _2194_/A _2155_/C _2194_/B vdd gnd NAND3X1
X_2224_ _2230_/A _2225_/C vdd gnd INVX1
X_2086_ _2095_/A _2095_/B _2123_/C _2100_/C vdd gnd OAI21X1
X_1939_ _2070_/A _2176_/B _1974_/B _1940_/A vdd gnd OAI21X1
X_2988_ _2988_/A _2988_/B _2991_/B _2991_/A _3021_/B vdd gnd OAI22X1
X_2911_ _2957_/S _3047_/Q _2912_/C vdd gnd NAND2X1
X_1724_ _1724_/A _1724_/B _1724_/C _1724_/D _1728_/D vdd gnd AOI22X1
X_2842_ _2842_/A _2842_/B _2842_/C _3074_/D vdd gnd OAI21X1
X_2773_ _2773_/A _2773_/B _2773_/C _3059_/D vdd gnd OAI21X1
X_1586_ _2455_/Q _1604_/A _1651_/B vdd gnd NAND2X1
X_1655_ _1655_/A _1655_/B _1666_/C _1687_/D vdd gnd AOI21X1
X_2069_ _2069_/A _2069_/B _2069_/C _2110_/C vdd gnd OAI21X1
X_2138_ _2146_/C _2146_/B _2190_/A _2190_/B vdd gnd NAND3X1
X_2207_ _2248_/A _2248_/B _2207_/C _2234_/B vdd gnd OAI21X1
X_1440_ _1686_/Q _1687_/Q _1452_/A vdd gnd AND2X2
X_3110_ _3110_/A y[7] vdd gnd BUFX2
X_3041_ _3041_/D _3098_/CLK _3041_/Q vdd gnd DFFPOSX1
X_2825_ _2992_/A _2853_/B _2853_/C _2826_/A vdd gnd OAI21X1
X_1638_ _1737_/B _1640_/B _1638_/C _1639_/B vdd gnd NAND3X1
X_1707_ _1719_/B _1720_/B vdd gnd INVX1
X_2687_ _3004_/A _2703_/B _2704_/B _2688_/D vdd gnd OAI21X1
X_2756_ _2780_/A _2996_/A _2780_/C _2757_/B vdd gnd AOI21X1
X_1569_ _1569_/D _3061_/CLK _3016_/A vdd gnd DFFPOSX1
X_2472_ _2507_/A _2516_/D vdd gnd INVX1
X_2541_ _2706_/B _2706_/C _2879_/A vdd gnd NAND2X1
X_2610_ _2610_/A _2610_/B _2667_/B _2611_/C vdd gnd MUX2X1
X_3024_ _3024_/D _3099_/CLK _3024_/Q vdd gnd DFFPOSX1
X_2808_ _3035_/Q _2816_/B _2810_/D vdd gnd NOR2X1
X_2739_ _3053_/Q _2742_/A vdd gnd INVX1
XBUFX2_insert40 _2488_/Y _2638_/S vdd gnd BUFX2
X_1972_ _2048_/A _2048_/B _1976_/C _1983_/C vdd gnd NAND3X1
X_2455_ _2455_/D _2462_/CLK _2455_/Q vdd gnd DFFPOSX1
X_2524_ _2524_/D _2535_/CLK _2524_/Q vdd gnd DFFPOSX1
X_2386_ _2386_/A _2388_/A _2387_/B vdd gnd NAND2X1
X_3007_ _3034_/Q _3019_/B _3009_/C vdd gnd NOR2X1
XCLKBUF1_insert3 clk _2469_/CLK vdd gnd CLKBUF1
X_2171_ _2171_/A _2220_/B _2171_/C _2231_/B vdd gnd OAI21X1
X_2240_ _2241_/A _2242_/A _2241_/B _2244_/B vdd gnd NAND3X1
X_1886_ _1999_/A _1886_/B _1887_/C vdd gnd NAND2X1
X_1955_ _2025_/A _2233_/A _2015_/A _2028_/C vdd gnd OAI21X1
X_2438_ _2438_/D _3087_/CLK _2438_/Q vdd gnd DFFPOSX1
X_2507_ _2507_/A _2507_/B _2507_/C _2522_/D vdd gnd OAI21X1
X_2369_ _2384_/B _2370_/A _2369_/C _2372_/B vdd gnd OAI21X1
X_1671_ _1671_/A _1671_/B _1737_/B _1672_/B vdd gnd OAI21X1
X_1740_ _2427_/Q _1800_/A vdd gnd INVX1
X_2085_ _2089_/C _2125_/D _2125_/C _2095_/A vdd gnd AOI21X1
X_2154_ _2154_/A _2154_/B _2154_/C _2162_/A vdd gnd OAI21X1
X_2223_ _2223_/A _2223_/B _2230_/B _2225_/B vdd gnd AOI21X1
X_2987_ _3094_/Q _2993_/A vdd gnd INVX1
X_1869_ _1869_/A _1869_/B _1870_/C vdd gnd NAND2X1
X_1938_ _2429_/Q _2437_/Q _1974_/B vdd gnd NAND2X1
X_2910_ _2910_/A _2910_/B _2982_/S _2913_/C vdd gnd MUX2X1
X_2841_ _3008_/A _2853_/B _2853_/C _2842_/A vdd gnd OAI21X1
X_1654_ _1654_/A _1654_/B _1658_/C _1686_/D vdd gnd AOI21X1
X_1723_ _1723_/A _1723_/B _1724_/A _1724_/C vdd gnd AOI21X1
X_2772_ _2780_/A _3012_/A _2780_/C _2773_/B vdd gnd AOI21X1
X_1585_ _1683_/Q _1630_/B _1651_/A vdd gnd NAND2X1
X_2206_ _2233_/A _2206_/B _2206_/C _2207_/C vdd gnd OAI21X1
X_2068_ _2068_/A _2068_/B _2068_/C _2069_/B vdd gnd AOI21X1
X_2137_ _2185_/B _2139_/B _2140_/A _2146_/B vdd gnd OAI21X1
X_3040_ _3040_/D _3075_/CLK _3040_/Q vdd gnd DFFPOSX1
X_2824_ _3030_/Q _2852_/B _2826_/B vdd gnd NOR2X1
X_1637_ _1676_/Q _1670_/B _1644_/A _1639_/A vdd gnd NAND3X1
X_1706_ _1723_/B _1720_/A vdd gnd INVX1
X_2686_ _3033_/Q _2702_/B _2688_/C vdd gnd NOR2X1
X_2755_ _3031_/Q _2779_/B _2757_/A vdd gnd NOR2X1
X_1499_ _1557_/Q _2507_/B _2706_/C vdd gnd AND2X2
X_1568_ _1568_/D _3097_/CLK _3012_/A vdd gnd DFFPOSX1
X_2471_ _2522_/Q _2530_/Y _2507_/A vdd gnd NOR2X1
X_2540_ _2602_/B _2667_/B _2668_/C _2662_/D vdd gnd NAND3X1
X_3023_ _3023_/D _3097_/CLK _3023_/Q vdd gnd DFFPOSX1
X_2738_ _2738_/A _2742_/B _2738_/C _2738_/D _3052_/D vdd gnd OAI22X1
X_2807_ _3067_/Q _2810_/A vdd gnd INVX1
X_2669_ _2785_/A _2982_/S _2712_/B vdd gnd NAND2X1
XBUFX2_insert41 _2488_/Y _2643_/S vdd gnd BUFX2
XBUFX2_insert30 _1556_/Q _1536_/B vdd gnd BUFX2
X_1971_ _2002_/A _1971_/B _1971_/C _2048_/B vdd gnd NAND3X1
X_2385_ _2385_/A _2385_/B _2388_/A vdd gnd AND2X2
X_2454_ _2454_/D _2469_/CLK _2454_/Q vdd gnd DFFPOSX1
X_2523_ _2523_/D _2535_/CLK _2523_/Q vdd gnd DFFPOSX1
X_3006_ _3098_/Q _3009_/A vdd gnd INVX1
XCLKBUF1_insert4 clk _3093_/CLK vdd gnd CLKBUF1
X_2170_ _2170_/A _2170_/B _2170_/C _2202_/B vdd gnd AOI21X1
X_1954_ _2028_/A _2087_/A _2016_/C vdd gnd NAND2X1
X_1885_ _2428_/Q _2437_/Q _1999_/A vdd gnd NAND2X1
X_2368_ _2368_/A _2451_/Q _2370_/A vdd gnd NOR2X1
X_2437_ _2437_/D _3087_/CLK _2437_/Q vdd gnd DFFPOSX1
X_2506_ _2508_/B _2506_/B _2507_/B _2507_/C vdd gnd OAI21X1
X_2299_ _2299_/A _2299_/B _2300_/B vdd gnd NAND2X1
X_1670_ _1679_/Q _1670_/B _1670_/C _1671_/A vdd gnd NAND3X1
X_2222_ _2231_/B _2223_/B vdd gnd INVX1
X_2084_ _2125_/A _2125_/B _2089_/C vdd gnd NAND2X1
X_2153_ _2153_/A _2154_/C _2163_/A _2163_/B _2158_/A vdd gnd AOI22X1
X_1937_ _1942_/C _1941_/C _1940_/C vdd gnd NAND2X1
X_2986_ _2986_/A _2986_/B _2986_/C _2986_/D _3093_/D vdd gnd AOI22X1
X_1799_ _1825_/B _1825_/A _1824_/B vdd gnd OR2X2
X_1868_ _1874_/B _1868_/B _1869_/B vdd gnd NOR2X1
X_2840_ _3034_/Q _2852_/B _2842_/B vdd gnd NOR2X1
X_2771_ _3035_/Q _2779_/B _2773_/A vdd gnd NOR2X1
X_1584_ _1604_/A _1630_/B vdd gnd INVX4
X_1653_ _1653_/A _1653_/B _1658_/C _1685_/D vdd gnd AOI21X1
X_1722_ _1750_/B _1724_/B vdd gnd INVX1
X_2205_ _2233_/C _2248_/B vdd gnd INVX1
X_2067_ _2108_/A _2154_/A vdd gnd INVX1
X_2136_ _2136_/A _2136_/B _2139_/B vdd gnd AND2X2
X_2969_ _3084_/Q _3028_/Q _2980_/S _2970_/A vdd gnd MUX2X1
X_1705_ _1753_/B _1724_/A _1712_/A vdd gnd NAND2X1
X_2754_ _3055_/Q _2779_/B _2778_/C _2757_/C vdd gnd NAND3X1
X_2823_ _2853_/B _2852_/B vdd gnd INVX2
X_1567_ _1567_/D _3061_/CLK _3008_/A vdd gnd DFFPOSX1
X_1636_ _1680_/Q _1703_/Q _1736_/A vdd gnd OR2X2
X_2685_ _3041_/Q _2936_/B vdd gnd INVX1
X_1498_ _1557_/Q _2499_/Y _2707_/B vdd gnd AND2X2
X_2119_ vdd _2160_/B _2120_/C vdd gnd NAND2X1
X_3099_ _3099_/D _3099_/CLK _3099_/Q vdd gnd DFFPOSX1
X_2470_ _2470_/D _2470_/CLK _2470_/Q vdd gnd DFFPOSX1
X_3022_ _3022_/D _3098_/CLK _3022_/Q vdd gnd DFFPOSX1
X_2668_ _2706_/B _2706_/C _2668_/C _2988_/B vdd gnd NAND3X1
X_2737_ _3016_/A _2741_/B _2742_/B _2738_/C vdd gnd OAI21X1
X_2806_ _2806_/A _2818_/B _2806_/C _2806_/D _3066_/D vdd gnd OAI22X1
X_1619_ _1619_/A _2466_/Q _1662_/B vdd gnd NAND2X1
X_2599_ _3023_/Q _2651_/B _2599_/C _2743_/A _2606_/D vdd gnd AOI22X1
XBUFX2_insert31 _1556_/Q _1517_/A vdd gnd BUFX2
XBUFX2_insert20 _1734_/Y _1669_/A vdd gnd BUFX2
X_1970_ _2038_/A _2039_/A _2039_/B _2048_/A vdd gnd NAND3X1
X_2522_ _2522_/D _3093_/CLK _2522_/Q vdd gnd DFFPOSX1
X_2384_ _2385_/B _2384_/B _2384_/C _2387_/A vdd gnd AOI21X1
X_2453_ _2453_/D _2470_/CLK _2453_/Q vdd gnd DFFPOSX1
X_3005_ _3005_/A _3021_/B _3005_/C _3005_/D _3097_/D vdd gnd OAI22X1
XCLKBUF1_insert5 clk _2535_/CLK vdd gnd CLKBUF1
X_1884_ _2428_/Q _2437_/Q _1884_/C _1887_/B vdd gnd NAND3X1
X_1953_ _2435_/Q _2432_/Q _2087_/A vdd gnd AND2X2
X_2505_ _2505_/A _2506_/B vdd gnd INVX1
X_2298_ _2314_/A _2343_/C _2299_/A vdd gnd NAND2X1
X_2367_ _2375_/A _2375_/B _2384_/B vdd gnd NOR2X1
X_2436_ _2436_/D _3087_/CLK _2436_/Q vdd gnd DFFPOSX1
X_2152_ _2155_/A _2156_/B _2156_/C _2163_/B vdd gnd NAND3X1
X_2221_ _2221_/A _2221_/B _2232_/A _2223_/A vdd gnd OAI21X1
X_2083_ _2173_/A _2125_/B vdd gnd INVX1
X_1867_ _1874_/A _1869_/A vdd gnd INVX1
X_1936_ _2428_/Q _2438_/Q _1941_/C vdd gnd AND2X2
X_2985_ _2985_/A _2985_/B _2985_/C _2985_/D _2986_/C vdd gnd AOI22X1
X_1798_ _1808_/A _1814_/C _1798_/C _1825_/B vdd gnd OAI21X1
X_2419_ _2424_/A _2424_/B vdd _2420_/B vdd gnd OAI21X1
X_1721_ _1724_/A _1721_/B _1721_/C _1721_/D _1727_/D vdd gnd AOI22X1
X_2770_ _3059_/Q _2779_/B _2778_/C _2773_/C vdd gnd NAND3X1
X_1583_ _1644_/A _1638_/C _1681_/D vdd gnd NOR2X1
X_1652_ _1652_/A _1652_/B _1669_/A _1684_/D vdd gnd AOI21X1
X_2135_ _2136_/B _2136_/A _2185_/B vdd gnd NOR2X1
X_2204_ _2204_/A _2206_/B _2233_/C vdd gnd NOR2X1
X_2066_ _2066_/A _2073_/A _2066_/C _2108_/A vdd gnd OAI21X1
X_1919_ _1988_/B _1988_/A _1922_/C vdd gnd AND2X2
X_2968_ _3068_/Q _3100_/Q _2980_/S _2970_/B vdd gnd MUX2X1
X_2899_ _2956_/S _3046_/Q _2900_/C vdd gnd NAND2X1
X_1704_ _1737_/B _1724_/A vdd gnd INVX2
X_2684_ _2924_/B _2704_/B _2684_/C _2684_/D _3040_/D vdd gnd OAI22X1
X_2753_ _2753_/A _2753_/B _2753_/C _3054_/D vdd gnd OAI21X1
X_2822_ _2822_/A _2860_/A _2853_/B vdd gnd NOR2X1
X_1497_ _1557_/Q _2497_/Y _2706_/B vdd gnd AND2X2
X_1566_ _1566_/D _3097_/CLK _3004_/A vdd gnd DFFPOSX1
X_1635_ _1701_/Q _1673_/B vdd gnd INVX1
X_2049_ _2049_/A _2049_/B _2049_/C _2052_/A vdd gnd OAI21X1
X_2118_ _2221_/A _2221_/B _2118_/C _2160_/B vdd gnd OAI21X1
X_3098_ _3098_/D _3098_/CLK _3098_/Q vdd gnd DFFPOSX1
X_3021_ _3021_/A _3021_/B _3021_/C _3021_/D _3101_/D vdd gnd OAI22X1
X_2805_ _3008_/A _2817_/B _2818_/B _2806_/C vdd gnd OAI21X1
X_1618_ _1694_/Q _1630_/B _1662_/A vdd gnd NAND2X1
X_2667_ _2743_/A _2667_/B _2708_/B vdd gnd NAND2X1
X_2736_ _3036_/Q _2740_/B _2738_/D vdd gnd NOR2X1
X_1549_ rst _1549_/B _1560_/D vdd gnd NOR2X1
X_2598_ _2598_/A _2598_/B _2667_/B _2599_/C vdd gnd MUX2X1
XBUFX2_insert32 _1556_/Q _1519_/A vdd gnd BUFX2
XBUFX2_insert21 _1734_/Y _1666_/C vdd gnd BUFX2
X_2521_ _2521_/D _3093_/CLK _2521_/Q vdd gnd DFFPOSX1
X_2383_ _2467_/Q _2426_/A _2400_/C vdd gnd NAND2X1
X_2452_ _2452_/D _2469_/CLK _2452_/Q vdd gnd DFFPOSX1
X_3004_ _3004_/A _3020_/B _3021_/B _3005_/D vdd gnd OAI21X1
X_2719_ _3048_/Q _2722_/A vdd gnd INVX1
XCLKBUF1_insert6 clk _3095_/CLK vdd gnd CLKBUF1
X_1883_ _1883_/A _1883_/B _1973_/A _1974_/C vdd gnd NAND3X1
X_1952_ _2016_/A _2028_/D vdd gnd INVX1
X_2435_ _2435_/D _3095_/CLK _2435_/Q vdd gnd DFFPOSX1
X_2504_ _2504_/A _2504_/B _2521_/D vdd gnd NAND2X1
X_2297_ _2297_/A _2312_/A _2314_/A vdd gnd NOR2X1
X_2366_ _2368_/A _2375_/A vdd gnd INVX1
X_2082_ _2082_/A _2090_/C _2095_/B vdd gnd NOR2X1
X_2151_ _2190_/B _2151_/B _2151_/C _2156_/B vdd gnd NAND3X1
X_2220_ _2220_/A _2220_/B _2232_/A vdd gnd NOR2X1
X_2984_ _2984_/A _2984_/B _2984_/C _2985_/B vdd gnd OAI21X1
X_1797_ _1895_/A _2071_/A _1834_/A _1798_/C vdd gnd OAI21X1
X_1866_ _1874_/B _1868_/B _1874_/A _1870_/B vdd gnd OAI21X1
X_1935_ _2429_/Q _2437_/Q _1942_/C vdd gnd AND2X2
X_2418_ _2422_/C _2424_/B vdd gnd INVX1
X_2349_ _2349_/A _2364_/B vdd gnd INVX1
X_1651_ _1651_/A _1651_/B _1669_/A _1683_/D vdd gnd AOI21X1
X_1720_ _1720_/A _1720_/B _1721_/D vdd gnd NAND2X1
X_1582_ _1737_/B _1644_/A vdd gnd INVX1
X_2065_ _2107_/B _2107_/A _2106_/C vdd gnd AND2X2
X_2134_ _2139_/C _2140_/B _2140_/C _2190_/A vdd gnd NAND3X1
X_2203_ _2203_/A _2203_/B _2203_/C _2234_/A vdd gnd AOI21X1
X_2967_ _2967_/A _2979_/B _2986_/A _2974_/D vdd gnd AOI21X1
X_1849_ _1856_/B _1856_/C _1876_/C _1916_/A vdd gnd NAND3X1
X_1918_ _1918_/A _1918_/B _1918_/C _1928_/A vdd gnd NAND3X1
X_2898_ _2898_/A _2898_/B _2982_/S _2901_/C vdd gnd MUX2X1
X_2821_ _3070_/Q _2851_/B _2826_/C vdd gnd NAND2X1
X_1634_ _1702_/Q _1668_/B vdd gnd INVX1
X_1703_ _1703_/D _3061_/CLK _1703_/Q vdd gnd DFFPOSX1
X_2683_ _3000_/A _2703_/B _2704_/B _2684_/D vdd gnd OAI21X1
X_2752_ _2780_/A _2992_/A _2780_/C _2753_/B vdd gnd AOI21X1
X_1496_ _1559_/Q _1496_/B _1496_/C _2785_/A vdd gnd OAI21X1
X_1565_ _1565_/D _3061_/CLK _3000_/A vdd gnd DFFPOSX1
X_2048_ _2048_/A _2048_/B _2048_/C _2049_/B vdd gnd AOI21X1
X_2117_ _2117_/A _2117_/B _2117_/C _2221_/B vdd gnd NOR3X1
X_3097_ _3097_/D _3097_/CLK _3097_/Q vdd gnd DFFPOSX1
X_3020_ _3020_/A _3020_/B _3021_/B _3021_/D vdd gnd OAI21X1
X_2804_ _3034_/Q _2816_/B _2806_/D vdd gnd NOR2X1
X_1617_ _1661_/B _1661_/A _2368_/A vdd gnd NAND2X1
X_2597_ _3047_/Q _3039_/Q _2706_/A _2598_/A vdd gnd MUX2X1
X_2666_ _3038_/Q _2900_/B vdd gnd INVX1
X_2735_ _3052_/Q _2738_/A vdd gnd INVX1
X_1479_ _1479_/A _1479_/B _1479_/C _1482_/B vdd gnd AOI21X1
X_1548_ _1559_/Q _1732_/Y _1548_/C _1549_/B vdd gnd NAND3X1
XBUFX2_insert33 _1699_/Q _1607_/A vdd gnd BUFX2
XBUFX2_insert22 _1490_/Y _2984_/A vdd gnd BUFX2
X_2451_ _2451_/D _2469_/CLK _2451_/Q vdd gnd DFFPOSX1
X_2520_ _2520_/D _2535_/CLK _2520_/Q vdd gnd DFFPOSX1
X_2382_ _2382_/A _2382_/B _2382_/C _2382_/D _2466_/D vdd gnd AOI22X1
X_3003_ _3033_/Q _3019_/B _3005_/C vdd gnd NOR2X1
X_2718_ _2718_/A _2742_/B _2718_/C _2718_/D _3047_/D vdd gnd OAI22X1
X_2649_ _3052_/Q _3044_/Q _2661_/S _2650_/A vdd gnd MUX2X1
XCLKBUF1_insert7 clk _3061_/CLK vdd gnd CLKBUF1
X_1882_ _2070_/A _2130_/A _1884_/C _1883_/A vdd gnd OAI21X1
X_1951_ _1960_/C _1960_/B _2016_/A _1965_/B vdd gnd AOI21X1
X_2365_ _2386_/A _2371_/B _2369_/C vdd gnd NOR2X1
X_2434_ _2434_/D _3095_/CLK _2434_/Q vdd gnd DFFPOSX1
X_2503_ _2511_/A _2509_/B _2515_/D _2504_/B vdd gnd OAI21X1
X_2296_ _2312_/A _2297_/A _2296_/C _2299_/B vdd gnd OAI21X1
X_2081_ _2081_/A _2173_/A _2125_/D _2090_/C vdd gnd OAI21X1
X_2150_ _2150_/A _2150_/B _2150_/C _2156_/C vdd gnd OAI21X1
X_1934_ _1943_/A _1940_/B vdd gnd INVX1
X_2983_ _2984_/A _3053_/Q _2984_/C vdd gnd NAND2X1
X_1796_ _2428_/Q _2434_/Q _1834_/A vdd gnd NAND2X1
X_1865_ _1874_/C _1868_/B vdd gnd INVX1
X_2348_ _2464_/Q _2358_/B vdd gnd INVX1
X_2417_ _2422_/A _2424_/A vdd gnd INVX1
X_2279_ _2294_/B _2284_/B vdd gnd INVX1
X_1581_ _1640_/B _1581_/B _1648_/A _1638_/C vdd gnd NAND3X1
X_1650_ _1650_/A _1650_/B _1679_/D vdd gnd NAND2X1
X_2202_ _2231_/B _2202_/B _2202_/C _2218_/C vdd gnd OAI21X1
X_2064_ _2170_/B _2170_/A _2232_/C vdd gnd NAND2X1
X_2133_ _2179_/A _2233_/B _2136_/A _2140_/B vdd gnd OAI21X1
X_1917_ _1980_/A _1921_/B _1921_/C _1918_/C vdd gnd NAND3X1
X_2966_ _2980_/S _2966_/B _2966_/C _2967_/A vdd gnd OAI21X1
X_2897_ _3078_/Q _3022_/Q _2945_/S _2898_/A vdd gnd MUX2X1
X_1779_ _2440_/Q _2206_/B vdd gnd INVX2
X_1848_ _1851_/A _2028_/A _1853_/B _1856_/C vdd gnd AOI21X1
X_2751_ _2822_/A _2991_/B _2780_/C vdd gnd NOR2X1
X_2820_ _2853_/C _2851_/B vdd gnd INVX2
X_1564_ _1564_/D _3101_/CLK _2996_/A vdd gnd DFFPOSX1
X_1633_ _1700_/Q _1667_/B vdd gnd INVX1
X_1702_ _1702_/D _3087_/CLK _1702_/Q vdd gnd DFFPOSX1
X_2682_ _3032_/Q _2702_/B _2684_/C vdd gnd NOR2X1
X_1495_ _1559_/Q _1719_/B _1496_/C vdd gnd NAND2X1
X_2047_ _2047_/A _2047_/B _2047_/C _2062_/C vdd gnd OAI21X1
X_2116_ _2170_/B _2221_/A vdd gnd INVX1
X_3096_ _3096_/D _3099_/CLK _3096_/Q vdd gnd DFFPOSX1
X_2949_ _2985_/A _2949_/B _2949_/C _2985_/D _2950_/C vdd gnd AOI22X1
X_2734_ _2734_/A _2742_/B _2734_/C _2734_/D _3051_/D vdd gnd OAI22X1
X_2803_ _3066_/Q _2806_/A vdd gnd INVX1
X_1547_ _1547_/A _1547_/B rst _1559_/D vdd gnd AOI21X1
X_1616_ _1619_/A _2465_/Q _1661_/B vdd gnd NAND2X1
X_2596_ _3071_/Q _3055_/Q _2706_/A _2598_/B vdd gnd MUX2X1
X_2665_ _2665_/A _2665_/B _2665_/C _2665_/D _3037_/D vdd gnd AOI22X1
X_1478_ _1483_/B _1483_/C _1481_/C vdd gnd NAND2X1
X_3079_ _3079_/D _3099_/CLK _3079_/Q vdd gnd DFFPOSX1
XBUFX2_insert34 _1699_/Q _1619_/A vdd gnd BUFX2
XBUFX2_insert23 _1490_/Y _2948_/A vdd gnd BUFX2
X_2381_ _2381_/A _2381_/B _2382_/A _2382_/D vdd gnd AOI21X1
X_2450_ _2450_/D _2469_/CLK _2450_/Q vdd gnd DFFPOSX1
X_3002_ _3097_/Q _3005_/A vdd gnd INVX1
X_2717_ _2996_/A _2741_/B _2742_/B _2718_/C vdd gnd OAI21X1
X_2579_ _2579_/A _2583_/B _2579_/C _2579_/D _3028_/D vdd gnd OAI22X1
X_2648_ _3076_/Q _3060_/Q _2661_/S _2650_/B vdd gnd MUX2X1
XCLKBUF1_insert8 clk _2462_/CLK vdd gnd CLKBUF1
X_1950_ _2025_/A _2233_/A _1958_/B _1960_/C vdd gnd OAI21X1
X_1881_ _2429_/Q _2436_/Q _1884_/C vdd gnd NAND2X1
X_2502_ _2502_/A _2507_/B _2504_/A vdd gnd NAND2X1
X_2364_ _2364_/A _2364_/B _2364_/C _2386_/A vdd gnd OAI21X1
X_2433_ _2433_/D _3095_/CLK _2433_/Q vdd gnd DFFPOSX1
X_2295_ _2343_/C _2296_/C vdd gnd INVX1
X_2080_ _2080_/A _2204_/A _2131_/A _2125_/D vdd gnd OAI21X1
X_1933_ _2427_/Q _2439_/Q _1943_/A vdd gnd NAND2X1
X_2982_ _2982_/A _2982_/B _2982_/S _2985_/C vdd gnd MUX2X1
X_1795_ _2434_/Q _2429_/Q _1814_/C vdd gnd NAND2X1
X_1864_ _1864_/A _1864_/B _1988_/B _1874_/C vdd gnd NAND3X1
X_2278_ _2278_/A _2278_/B _2278_/C _2294_/B vdd gnd AOI21X1
X_2347_ _2347_/A _2347_/B _2347_/C _2463_/D vdd gnd OAI21X1
X_2416_ _2422_/A _2422_/C _2420_/A vdd gnd NOR2X1
X_1580_ _1677_/Q _1678_/Q _1581_/B vdd gnd NOR2X1
X_2132_ _2136_/A _2136_/B _2140_/C vdd gnd OR2X2
X_2201_ _2230_/B _2202_/C vdd gnd INVX1
X_2063_ _2063_/A _2063_/B _2063_/C _2170_/A vdd gnd NAND3X1
X_1847_ _2433_/Q _2431_/Q _2434_/Q _2430_/Q _1853_/B vdd gnd AOI22X1
X_1916_ _1916_/A _1979_/A _1979_/B _1921_/B vdd gnd NAND3X1
X_2965_ _2980_/S _3076_/Q _2966_/C vdd gnd NAND2X1
X_2896_ _3062_/Q _3094_/Q _2956_/S _2898_/B vdd gnd MUX2X1
X_1778_ vdd _2233_/B _1778_/C _2439_/D vdd gnd OAI21X1
X_1701_ _1701_/D _3087_/CLK _1701_/Q vdd gnd DFFPOSX1
X_2681_ _3040_/Q _2924_/B vdd gnd INVX1
X_2750_ _2819_/A _2988_/B _2780_/A vdd gnd NOR2X1
X_1494_ _2517_/Q _1496_/B vdd gnd INVX1
X_1563_ _1563_/D _3061_/CLK _2992_/A vdd gnd DFFPOSX1
X_1632_ _1666_/B _1666_/A _2423_/A vdd gnd NAND2X1
X_2115_ _2118_/C _2232_/C _2120_/D vdd gnd NOR2X1
X_3095_ _3095_/D _3095_/CLK _3095_/Q vdd gnd DFFPOSX1
X_2046_ _2050_/C _2107_/A _2050_/A _2047_/A vdd gnd AOI21X1
X_2948_ _2948_/A _2948_/B _2948_/C _2949_/B vdd gnd OAI21X1
X_2879_ _2879_/A _2879_/B _2887_/B _2889_/B vdd gnd OAI21X1
X_2664_ _2664_/A _3085_/Q _2665_/A _2665_/D vdd gnd AOI21X1
X_2733_ _3012_/A _2741_/B _2742_/B _2734_/C vdd gnd OAI21X1
X_2802_ _2802_/A _2818_/B _2802_/C _2802_/D _3065_/D vdd gnd OAI22X1
X_1477_ _1693_/Q _1477_/B _1694_/Q _1483_/C vdd gnd OAI21X1
X_1546_ _1546_/A _1548_/C _1547_/A vdd gnd NAND2X1
X_1615_ _1693_/Q _1630_/B _1661_/A vdd gnd NAND2X1
X_2595_ _2662_/D _2651_/B vdd gnd INVX2
X_3078_ _3078_/D _3097_/CLK _3078_/Q vdd gnd DFFPOSX1
X_2029_ _2088_/B _2088_/A _2075_/C _2068_/A vdd gnd NAND3X1
XBUFX2_insert24 _1490_/Y _2980_/S vdd gnd BUFX2
XBUFX2_insert13 _1872_/Y _2358_/A vdd gnd BUFX2
XBUFX2_insert35 _1699_/Q _1631_/A vdd gnd BUFX2
X_2380_ _2381_/A _2381_/B _2382_/C vdd gnd OR2X2
X_3001_ _3001_/A _3021_/B _3001_/C _3001_/D _3096_/D vdd gnd OAI22X1
X_2647_ _3036_/Q _2656_/B vdd gnd INVX1
X_2716_ _3031_/Q _2740_/B _2718_/D vdd gnd NOR2X1
X_1529_ _1537_/C _1529_/B _1529_/C _1543_/B vdd gnd NAND3X1
X_2578_ _3016_/A _2582_/B _2583_/B _2579_/D vdd gnd OAI21X1
XCLKBUF1_insert9 clk _2470_/CLK vdd gnd CLKBUF1
X_1880_ _1886_/B _1880_/B _1973_/A vdd gnd NAND2X1
X_2501_ _2511_/A _2511_/C _2501_/C _2532_/A vdd gnd OAI21X1
X_2294_ _2294_/A _2294_/B _2294_/C _2343_/C vdd gnd OAI21X1
X_2363_ _2363_/A _2364_/C vdd gnd INVX1
X_2432_ _2432_/D _2535_/CLK _2432_/Q vdd gnd DFFPOSX1
X_1863_ _1988_/B _1864_/B _1864_/A _1874_/B vdd gnd AOI21X1
X_1932_ _1932_/A _1932_/B _1968_/A _2048_/C vdd gnd OAI21X1
X_2981_ _3085_/Q _3029_/Q _2984_/A _2982_/A vdd gnd MUX2X1
X_1794_ _2427_/Q _2435_/Q _1825_/A vdd gnd NAND2X1
X_2415_ _2415_/A _2415_/B _2415_/C _2422_/C vdd gnd OAI21X1
X_2277_ _2332_/A _2277_/B _2277_/C _2457_/D vdd gnd OAI21X1
X_2346_ _2360_/A _2389_/B vdd _2347_/A vdd gnd OAI21X1
X_2062_ _2062_/A _2062_/B _2062_/C _2170_/B vdd gnd OAI21X1
X_2131_ _2131_/A _2131_/B _2131_/C _2136_/A vdd gnd OAI21X1
X_2200_ _2452_/Q _2358_/A _2227_/A vdd gnd NAND2X1
X_2964_ _3060_/Q _2966_/B vdd gnd INVX1
X_1777_ vdd _3092_/Q _1778_/C vdd gnd NAND2X1
X_1846_ _2434_/Q _2431_/Q _2028_/A vdd gnd AND2X2
X_1915_ _1979_/C _1915_/B _1921_/C vdd gnd NAND2X1
X_2895_ _2895_/A _2979_/B _2986_/A _2902_/D vdd gnd AOI21X1
X_2329_ _2329_/A _2331_/A vdd gnd INVX1
X_1631_ _1631_/A _2470_/Q _1666_/B vdd gnd NAND2X1
X_1700_ _1700_/D _3087_/CLK _1700_/Q vdd gnd DFFPOSX1
X_2680_ _2912_/B _2704_/B _2680_/C _2680_/D _3039_/D vdd gnd OAI22X1
X_1493_ _1559_/Q _1493_/B _1493_/C _2783_/A vdd gnd OAI21X1
X_1562_ _1562_/D _3093_/CLK _1737_/B vdd gnd DFFPOSX1
X_2045_ _2045_/A _2045_/B _2045_/C _2050_/C vdd gnd OAI21X1
X_2114_ _2220_/A _2118_/C vdd gnd INVX1
X_3094_ _3094_/D _3099_/CLK _3094_/Q vdd gnd DFFPOSX1
X_2947_ _2948_/A _3050_/Q _2948_/C vdd gnd NAND2X1
X_1829_ vdd _1874_/A _1830_/D vdd gnd NAND2X1
X_2878_ _2878_/A _2878_/B _2878_/C _3082_/D vdd gnd NAND3X1
X_2801_ _3004_/A _2817_/B _2818_/B _2802_/C vdd gnd OAI21X1
X_1614_ _1660_/B _1660_/A _2353_/A vdd gnd NAND2X1
X_2594_ _3031_/Q _2606_/B vdd gnd INVX1
X_2663_ _2743_/A _2663_/B _2663_/C _2665_/C vdd gnd AOI21X1
X_2732_ _3035_/Q _2740_/B _2734_/D vdd gnd NOR2X1
X_1476_ _1695_/Q _1483_/B vdd gnd INVX1
X_1545_ _1545_/A _1545_/B _1548_/C vdd gnd NOR2X1
X_2028_ _2028_/A _2087_/A _2028_/C _2028_/D _2035_/C vdd gnd AOI22X1
X_3077_ _3077_/D _3101_/CLK _3077_/Q vdd gnd DFFPOSX1
XBUFX2_insert36 _1699_/Q _1604_/A vdd gnd BUFX2
XBUFX2_insert25 _1490_/Y _2960_/A vdd gnd BUFX2
XBUFX2_insert14 _1872_/Y _2332_/A vdd gnd BUFX2
X_3000_ _3000_/A _3020_/B _3021_/B _3001_/D vdd gnd OAI21X1
X_2577_ _3036_/Q _2581_/B _2579_/C vdd gnd NOR2X1
X_2646_ _2665_/A _2646_/B _2646_/C _2646_/D _3035_/D vdd gnd AOI22X1
X_2715_ _3047_/Q _2718_/A vdd gnd INVX1
X_1459_ _1691_/Q _1459_/B _1461_/A vdd gnd NOR2X1
X_1528_ _1536_/B _1528_/B _1529_/C vdd gnd NOR2X1
X_2431_ _2431_/D _3087_/CLK _2431_/Q vdd gnd DFFPOSX1
X_2500_ _2520_/Q _2501_/C vdd gnd INVX1
X_2293_ _2293_/A _2294_/C vdd gnd INVX1
X_2362_ _2362_/A _2389_/B _2371_/B vdd gnd NOR2X1
X_2629_ _3050_/Q _3042_/Q _2633_/S _2630_/A vdd gnd MUX2X1
X_2980_ _3069_/Q _3101_/Q _2980_/S _2982_/B vdd gnd MUX2X1
X_1793_ _2443_/Q _2270_/B vdd gnd INVX1
X_1862_ _1862_/A _1862_/B _1862_/C _1864_/B vdd gnd NAND3X1
X_1931_ _1931_/A _1931_/B _1931_/C _1932_/B vdd gnd AOI21X1
X_2414_ _2414_/A _2415_/A vdd gnd INVX1
X_2276_ _2457_/Q _2332_/A _2277_/C vdd gnd NAND2X1
X_2345_ _2389_/B _2360_/A _2347_/B vdd gnd AND2X2
X_2061_ _2061_/A _2062_/B vdd gnd INVX1
X_2130_ _2130_/A _2204_/A _2180_/A _2131_/C vdd gnd OAI21X1
X_1914_ _1930_/A _1980_/A vdd gnd INVX1
X_2963_ _3092_/Q _2974_/B vdd gnd INVX1
X_1776_ _2439_/Q _2233_/B vdd gnd INVX2
X_1845_ _1845_/A _1845_/B _1845_/C _1856_/B vdd gnd NAND3X1
X_2894_ _2960_/A _2894_/B _2894_/C _2895_/A vdd gnd OAI21X1
X_2328_ _2330_/B _2339_/B _2329_/A _2332_/D vdd gnd OAI21X1
X_2259_ _2261_/A _2268_/A vdd gnd INVX1
X_1630_ _1698_/Q _1630_/B _1666_/A vdd gnd NAND2X1
X_1492_ _1559_/Q _1723_/B _1493_/C vdd gnd NAND2X1
X_1561_ _1561_/D _2535_/CLK _2533_/B vdd gnd DFFPOSX1
X_2044_ _2044_/A _2044_/B _2044_/C _2107_/A vdd gnd NAND3X1
X_2113_ _2169_/A _2171_/A _2220_/A vdd gnd NAND2X1
X_3093_ _3093_/D _3093_/CLK _3093_/Q vdd gnd DFFPOSX1
X_2946_ _2946_/A _2946_/B _2982_/S _2949_/C vdd gnd MUX2X1
X_2877_ _3034_/Q _2888_/C _2878_/A vdd gnd NAND2X1
X_1759_ vdd _3086_/Q _1760_/C vdd gnd NAND2X1
X_1828_ _1828_/A _1832_/A _1828_/C _1874_/A vdd gnd NAND3X1
X_2731_ _3051_/Q _2734_/A vdd gnd INVX1
X_2800_ _3033_/Q _2816_/B _2802_/D vdd gnd NOR2X1
X_1544_ _1732_/Y _1546_/A vdd gnd INVX1
X_1613_ _1619_/A _2464_/Q _1660_/B vdd gnd NAND2X1
X_2593_ _2665_/A _2593_/B _2593_/C _3030_/D vdd gnd OAI21X1
X_2662_ _2988_/A _2662_/B _2662_/C _2662_/D _2663_/C vdd gnd OAI22X1
X_1475_ _1475_/A _1475_/B _1484_/B _3108_/A vdd gnd NAND3X1
X_2027_ _2035_/A _2035_/B _2068_/C _2041_/C vdd gnd OAI21X1
X_3076_ _3076_/D _3101_/CLK _3076_/Q vdd gnd DFFPOSX1
XBUFX2_insert37 _2488_/Y _2706_/A vdd gnd BUFX2
XBUFX2_insert26 _1490_/Y _2945_/S vdd gnd BUFX2
XBUFX2_insert15 _1872_/Y _2311_/B vdd gnd BUFX2
X_2929_ _2948_/A _3073_/Q _2930_/C vdd gnd NAND2X1
X_2714_ _2714_/A _2742_/B _2714_/C _2714_/D _3046_/D vdd gnd OAI22X1
X_1527_ _1557_/Q _1528_/B vdd gnd INVX1
X_2576_ _3028_/Q _2579_/A vdd gnd INVX1
X_2645_ _2665_/A _2645_/B _2646_/C vdd gnd NOR2X1
X_1458_ _1690_/Q _1459_/B vdd gnd INVX1
X_3059_ _3059_/D _3075_/CLK _3059_/Q vdd gnd DFFPOSX1
X_2361_ _2388_/B _2362_/A vdd gnd INVX1
X_2430_ _2430_/D _2535_/CLK _2430_/Q vdd gnd DFFPOSX1
X_2292_ _2292_/A _2445_/Q _2297_/A vdd gnd NOR2X1
X_2559_ _2559_/A _2583_/B _2559_/C _2559_/D _3023_/D vdd gnd OAI22X1
X_2628_ _3074_/Q _3058_/Q _2638_/S _2630_/B vdd gnd MUX2X1
X_1930_ _1930_/A _1930_/B _1930_/C _1978_/C vdd gnd AOI21X1
X_1792_ _2268_/B vdd _1792_/C _2442_/D vdd gnd OAI21X1
X_1861_ _1861_/A _1916_/A _1861_/C _1862_/B vdd gnd NAND3X1
X_2344_ _2344_/A _2344_/B _2389_/B vdd gnd AND2X2
X_2413_ _2413_/A _2413_/B _2414_/A vdd gnd NOR2X1
X_2275_ _2275_/A _2275_/B _2277_/B vdd gnd NAND2X1
X_2060_ _2449_/Q _2335_/B vdd gnd INVX1
X_1913_ _1930_/A _1980_/C _1930_/B _1918_/B vdd gnd NAND3X1
X_2962_ _2986_/A _2962_/B _2962_/C _2962_/D _3091_/D vdd gnd AOI22X1
X_2893_ _2956_/S _3070_/Q _2894_/C vdd gnd NAND2X1
X_1775_ vdd _2176_/B _1775_/C _2438_/D vdd gnd OAI21X1
X_1844_ _2429_/Q _2435_/Q _1974_/A _1845_/C vdd gnd NAND3X1
X_2258_ _2311_/B _2258_/B _2258_/C _2455_/D vdd gnd OAI21X1
X_2327_ _2327_/A _2448_/Q _2339_/B vdd gnd NOR2X1
X_2189_ _2190_/A _2190_/B _2189_/C _2195_/A vdd gnd NAND3X1
X_1560_ _1560_/D _3061_/CLK _3102_/A vdd gnd DFFPOSX1
X_1491_ _2516_/Q _1493_/B vdd gnd INVX1
X_2112_ _2112_/A _2153_/A _2112_/C _2171_/A vdd gnd NAND3X1
X_2043_ _2051_/C _2051_/B _2051_/A _2047_/B vdd gnd AOI21X1
X_3092_ _3092_/D _3093_/CLK _3092_/Q vdd gnd DFFPOSX1
X_1827_ _1828_/C _1832_/A _1828_/A _1830_/C vdd gnd AOI21X1
X_2945_ _3082_/Q _3026_/Q _2945_/S _2946_/A vdd gnd MUX2X1
X_2876_ _3082_/Q _2887_/B _2876_/C _2878_/C vdd gnd NAND3X1
X_1689_ _1689_/D _2462_/CLK _1689_/Q vdd gnd DFFPOSX1
X_1758_ _2433_/Q _1895_/A vdd gnd INVX1
X_2661_ _3069_/Q _3101_/Q _2661_/S _2662_/B vdd gnd MUX2X1
X_2730_ _2730_/A _2742_/B _2730_/C _2730_/D _3050_/D vdd gnd OAI22X1
X_1474_ _1474_/A _1479_/C _1475_/B vdd gnd OR2X2
X_1543_ _1543_/A _1543_/B _1558_/D vdd gnd NOR2X1
X_1612_ _1692_/Q _1630_/B _1660_/A vdd gnd NAND2X1
X_2592_ _2592_/A _2592_/B _2743_/A _2593_/B vdd gnd MUX2X1
X_3075_ _3075_/D _3075_/CLK _3075_/Q vdd gnd DFFPOSX1
X_2026_ _2075_/C _2088_/B _2088_/A _2035_/A vdd gnd AOI21X1
XBUFX2_insert38 _2488_/Y _2661_/S vdd gnd BUFX2
XBUFX2_insert27 _1490_/Y _2957_/S vdd gnd BUFX2
XBUFX2_insert16 _1872_/Y _2382_/A vdd gnd BUFX2
X_2928_ _3057_/Q _2930_/B vdd gnd INVX1
X_2859_ _3078_/Q _2887_/B _2876_/C _2862_/C vdd gnd NAND3X1
X_2644_ _2882_/A _2879_/B _2988_/A _2644_/D _2645_/B vdd gnd OAI22X1
X_2713_ _2992_/A _2741_/B _2742_/B _2714_/C vdd gnd OAI21X1
X_1457_ _1457_/A _1457_/B _1468_/A vdd gnd NAND2X1
X_1526_ _1558_/Q _1559_/Q _1529_/B vdd gnd NOR2X1
X_2575_ _2575_/A _2583_/B _2575_/C _2575_/D _3027_/D vdd gnd OAI22X1
X_3058_ _3058_/D _3098_/CLK _3058_/Q vdd gnd DFFPOSX1
X_2009_ _2009_/A _2009_/B _2009_/C _2066_/C vdd gnd NAND3X1
X_2291_ _2291_/A _2291_/B _2312_/A vdd gnd NOR2X1
X_2360_ _2360_/A _2360_/B _2388_/B vdd gnd NOR2X1
X_2627_ _3034_/Q _2636_/B vdd gnd INVX1
X_1509_ _3004_/A _1511_/B vdd gnd INVX1
X_2489_ _2508_/B _2491_/A vdd gnd INVX1
X_2558_ _2996_/A _2582_/B _2583_/B _2559_/D vdd gnd OAI21X1
X_1860_ _1860_/A _1979_/C _1860_/C _1862_/C vdd gnd OAI21X1
X_1791_ vdd _1791_/B _1791_/C _1792_/C vdd gnd NAND3X1
X_2274_ _2278_/A _2278_/B _2275_/B vdd gnd OR2X2
X_2343_ _2343_/A _2343_/B _2343_/C _2344_/A vdd gnd NAND3X1
X_2412_ _2412_/A _2412_/B _2412_/C _2415_/C vdd gnd AOI21X1
X_1989_ _1989_/A _1989_/B _1989_/C _2117_/C vdd gnd AOI21X1
X_1843_ _2428_/Q _2436_/Q _1974_/A vdd gnd NAND2X1
X_1912_ _1916_/A _1915_/B _1930_/B vdd gnd NAND2X1
X_2961_ _2985_/A _2961_/B _2961_/C _2985_/D _2962_/C vdd gnd AOI22X1
X_2892_ _3054_/Q _2894_/B vdd gnd INVX1
X_1774_ vdd _3091_/Q _1775_/C vdd gnd NAND2X1
X_2257_ _2455_/Q _2311_/B _2258_/C vdd gnd NAND2X1
X_2326_ _2339_/C _2330_/B vdd gnd INVX1
X_2188_ _2212_/A _2191_/B _2189_/C vdd gnd NAND2X1
X_1490_ _1559_/Q _1490_/B _1490_/C _1490_/Y vdd gnd OAI21X1
X_2042_ _2044_/C _2044_/B _2045_/C _2051_/C vdd gnd NAND3X1
X_2111_ _2154_/B _2111_/B _2154_/A _2112_/C vdd gnd OAI21X1
X_3091_ _3091_/D _3095_/CLK _3091_/Q vdd gnd DFFPOSX1
X_1826_ _1861_/A _1826_/B _1826_/C _1832_/A vdd gnd NAND3X1
X_2944_ _3066_/Q _3098_/Q _2945_/S _2946_/B vdd gnd MUX2X1
X_2875_ _3008_/A _2887_/B _2888_/A _2878_/B vdd gnd NAND3X1
X_1688_ _1688_/D _2462_/CLK _1688_/Q vdd gnd DFFPOSX1
X_1757_ vdd _2204_/A _1757_/C _2432_/D vdd gnd OAI21X1
X_2309_ _2309_/A _2309_/B vdd _2310_/C vdd gnd OAI21X1
X_1611_ _1659_/B _1659_/A _2336_/A vdd gnd NAND2X1
X_2660_ _2660_/A _2660_/B _2667_/B _2663_/B vdd gnd MUX2X1
X_1473_ _1693_/Q _1477_/B _1479_/C _1475_/A vdd gnd OAI21X1
X_1542_ _1557_/Q _2528_/Y _1542_/C _1543_/A vdd gnd NAND3X1
X_2591_ _2591_/A _2591_/B _2743_/B _2592_/A vdd gnd MUX2X1
X_2025_ _2025_/A _2204_/A _2081_/A _2088_/B vdd gnd OAI21X1
X_3074_ _3074_/D _3098_/CLK _3074_/Q vdd gnd DFFPOSX1
X_2927_ _3089_/Q _2938_/B vdd gnd INVX1
X_1809_ _2427_/Q _2436_/Q _1818_/A vdd gnd NAND2X1
XBUFX2_insert39 _2488_/Y _2633_/S vdd gnd BUFX2
XBUFX2_insert28 _1490_/Y _2956_/S vdd gnd BUFX2
XBUFX2_insert17 _1872_/Y _2426_/A vdd gnd BUFX2
X_2858_ _2879_/B _2879_/A _2876_/C vdd gnd OR2X2
X_2789_ _2992_/A _2817_/B _2818_/B _2790_/C vdd gnd OAI21X1
X_2574_ _3012_/A _2582_/B _2583_/B _2575_/D vdd gnd OAI21X1
X_2643_ _3067_/Q _3099_/Q _2643_/S _2644_/D vdd gnd MUX2X1
X_2712_ _2860_/A _2712_/B _2741_/B vdd gnd NOR2X1
X_1456_ _1466_/B _1456_/B _1484_/B _3104_/A vdd gnd OAI21X1
X_1525_ _3102_/A _1537_/C vdd gnd INVX1
X_2008_ _2071_/A _2176_/B _2073_/A _2009_/A vdd gnd OAI21X1
X_3057_ _3057_/D _3098_/CLK _3057_/Q vdd gnd DFFPOSX1
X_2290_ _2292_/A _2291_/A vdd gnd INVX1
X_2557_ _3031_/Q _2581_/B _2559_/C vdd gnd NOR2X1
X_2626_ _2665_/A _2626_/B _2626_/C _2626_/D _3033_/D vdd gnd AOI22X1
X_1439_ _1692_/Q _1460_/B vdd gnd INVX1
X_1508_ _1522_/A _1508_/B _1508_/C _1565_/D vdd gnd OAI21X1
X_2488_ _2491_/C _2511_/C _2515_/D _2488_/Y vdd gnd AOI21X1
X_3109_ _3109_/A y[6] vdd gnd BUFX2
X_1790_ _1800_/A _1816_/A _1808_/A _1791_/B vdd gnd OAI21X1
X_2411_ _2469_/Q _2426_/A _2420_/C vdd gnd NAND2X1
X_2273_ _2278_/B _2278_/A _2275_/A vdd gnd NAND2X1
X_2342_ _2343_/B _2342_/B _2342_/C _2344_/B vdd gnd AOI21X1
X_1988_ _1988_/A _1988_/B _1988_/C _1988_/D _1989_/C vdd gnd AOI22X1
X_2609_ _3048_/Q _3040_/Q _2643_/S _2610_/A vdd gnd MUX2X1
X_2960_ _2960_/A _2960_/B _2960_/C _2961_/B vdd gnd OAI21X1
X_1773_ _2438_/Q _2176_/B vdd gnd INVX2
X_1842_ _2428_/Q _2436_/Q _1876_/A _1845_/B vdd gnd NAND3X1
X_1911_ _1979_/A _1979_/B _1915_/B vdd gnd NAND2X1
X_2891_ _3086_/Q _2902_/B vdd gnd INVX1
X_2187_ _2187_/A _2187_/B _2191_/B vdd gnd NAND2X1
X_2256_ _2256_/A _2264_/C _2258_/B vdd gnd NAND2X1
X_2325_ _2327_/A _2448_/Q _2339_/C vdd gnd NAND2X1
X_2041_ _2069_/A _2041_/B _2041_/C _2044_/B vdd gnd NAND3X1
X_2110_ _2110_/A _2110_/B _2110_/C _2154_/B vdd gnd AOI21X1
X_3090_ _3090_/D _3099_/CLK _3090_/Q vdd gnd DFFPOSX1
X_2943_ _2943_/A _2979_/B _2986_/A _2950_/D vdd gnd AOI21X1
X_1756_ vdd _1756_/B _1757_/C vdd gnd NAND2X1
X_1825_ _1825_/A _1825_/B _1825_/C _1826_/B vdd gnd OAI21X1
X_2874_ _2874_/A _2874_/B _2874_/C _3081_/D vdd gnd NAND3X1
X_1687_ _1687_/D _2470_/CLK _1687_/Q vdd gnd DFFPOSX1
X_2308_ _2308_/A _2314_/B _2309_/B vdd gnd AND2X2
X_2239_ _2250_/A _2239_/B _2242_/A vdd gnd NAND2X1
X_1610_ _1619_/A _2463_/Q _1659_/B vdd gnd NAND2X1
X_2590_ _3070_/Q _3054_/Q _2638_/S _2591_/A vdd gnd MUX2X1
X_1472_ _1474_/A _1472_/B _1481_/B _1481_/A _3107_/A vdd gnd AOI22X1
X_1541_ _1541_/A _1542_/C _1557_/D vdd gnd AND2X2
X_2024_ _2431_/Q _2436_/Q _2081_/A vdd gnd NAND2X1
X_3073_ _3073_/D _3098_/CLK _3073_/Q vdd gnd DFFPOSX1
XBUFX2_insert29 _1556_/Q _1522_/A vdd gnd BUFX2
XBUFX2_insert18 _1734_/Y _1665_/C vdd gnd BUFX2
X_2926_ _2986_/A _2926_/B _2926_/C _2926_/D _3088_/D vdd gnd AOI22X1
X_2857_ _2992_/A _2887_/B _2888_/A _2862_/B vdd gnd NAND3X1
X_1739_ _1739_/D _3093_/CLK _1739_/Q vdd gnd DFFPOSX1
X_1808_ _1808_/A _1814_/C _1825_/C vdd gnd OR2X2
X_2788_ _2860_/A _2991_/A _2817_/B vdd gnd NOR2X1
X_2711_ _3030_/Q _2740_/B _2714_/D vdd gnd NOR2X1
X_1524_ rst _1542_/C vdd gnd INVX1
X_2573_ _3035_/Q _2581_/B _2575_/C vdd gnd NOR2X1
X_2642_ _3083_/Q _2882_/A vdd gnd INVX1
X_1455_ _1690_/Q _1461_/C _1456_/B vdd gnd NOR2X1
X_2007_ _2428_/Q _2439_/Q _2073_/A vdd gnd NAND2X1
X_3056_ _3056_/D _3098_/CLK _3056_/Q vdd gnd DFFPOSX1
X_2909_ _3079_/Q _3023_/Q _2984_/A _2910_/A vdd gnd MUX2X1
X_1507_ _1522_/A x[2] _1508_/C vdd gnd NAND2X1
X_2487_ _2511_/B _2491_/C vdd gnd INVX1
X_2556_ _3023_/Q _2559_/A vdd gnd INVX1
X_2625_ _2664_/A _3081_/Q _2665_/A _2626_/D vdd gnd AOI21X1
X_1438_ _1691_/Q _1457_/A vdd gnd INVX1
X_3108_ _3108_/A y[5] vdd gnd BUFX2
X_3039_ _3039_/D _3095_/CLK _3039_/Q vdd gnd DFFPOSX1
X_2341_ _2341_/A _2341_/B _2343_/B vdd gnd NOR2X1
X_2410_ _2426_/A _2410_/B _2410_/C _2410_/D _2468_/D vdd gnd AOI22X1
X_2272_ _2272_/A _2278_/C _2278_/B vdd gnd NOR2X1
X_1987_ _2063_/A _2063_/C _1991_/B vdd gnd NOR2X1
X_2539_ _2706_/A _2668_/C vdd gnd INVX1
X_2608_ _3072_/Q _3056_/Q _2633_/S _2610_/B vdd gnd MUX2X1
X_1910_ _1979_/C _1979_/A _1979_/B _1980_/C vdd gnd NAND3X1
X_2890_ _2890_/A _2986_/A vdd gnd INVX4
X_1772_ vdd _2130_/A _1772_/C _2437_/D vdd gnd OAI21X1
X_1841_ _1841_/A _1841_/B _1841_/C _1876_/C vdd gnd NAND3X1
X_2324_ _2324_/A _2324_/B _2339_/A _2329_/A vdd gnd OAI21X1
X_2186_ _2186_/A _2186_/B _2187_/A vdd gnd NAND2X1
X_2255_ _2255_/A _2255_/B _2256_/A vdd gnd NAND2X1
X_2040_ _2069_/C _2040_/B _2040_/C _2044_/C vdd gnd NAND3X1
X_2942_ _2948_/A _2942_/B _2942_/C _2943_/A vdd gnd OAI21X1
X_2873_ _3033_/Q _2888_/C _2874_/A vdd gnd NAND2X1
X_1686_ _1686_/D _2462_/CLK _1686_/Q vdd gnd DFFPOSX1
X_1755_ _2432_/Q _2204_/A vdd gnd INVX2
X_1824_ _1825_/C _1824_/B _1824_/C _1828_/C vdd gnd NAND3X1
X_2238_ _2238_/A _2238_/B _2250_/A vdd gnd NAND2X1
X_2307_ _2314_/B _2308_/A _2309_/A vdd gnd NOR2X1
X_2169_ _2169_/A _2171_/A _2169_/C _2170_/C vdd gnd NAND3X1
X_1540_ _2528_/Y _1543_/B _1552_/B _1541_/A vdd gnd OAI21X1
X_1471_ _1693_/Q _1477_/B _1472_/B vdd gnd NAND2X1
X_2023_ _2087_/A _2125_/A _2075_/C vdd gnd NAND2X1
X_3072_ _3072_/D _3098_/CLK _3072_/Q vdd gnd DFFPOSX1
X_1807_ _2444_/Q _2281_/B vdd gnd INVX1
XBUFX2_insert19 _1734_/Y _1658_/C vdd gnd BUFX2
X_2925_ _2985_/A _2925_/B _2925_/C _2985_/D _2926_/C vdd gnd AOI22X1
X_2856_ _2856_/A _2856_/B _2887_/B vdd gnd NAND2X1
X_1669_ _1669_/A _1669_/B _1669_/C _1671_/B vdd gnd OAI21X1
X_1738_ _1738_/D _3093_/CLK _1738_/Q vdd gnd DFFPOSX1
X_2787_ _3030_/Q _2816_/B _2790_/D vdd gnd NOR2X1
X_2710_ _2856_/B _2985_/A _2740_/B vdd gnd NAND2X1
X_1454_ _1457_/B _1466_/B vdd gnd INVX1
X_1523_ _1536_/B _1523_/B _1523_/C _1570_/D vdd gnd OAI21X1
X_2572_ _3027_/Q _2575_/A vdd gnd INVX1
X_2641_ _3027_/Q _2651_/B _2641_/C _2743_/A _2646_/D vdd gnd AOI22X1
X_3055_ _3055_/D _3097_/CLK _3055_/Q vdd gnd DFFPOSX1
X_2006_ _2011_/C _2122_/A _2009_/C vdd gnd NAND2X1
X_2908_ _3063_/Q _3095_/Q _2957_/S _2910_/B vdd gnd MUX2X1
X_2839_ _3074_/Q _2851_/B _2842_/C vdd gnd NAND2X1
X_2624_ _2879_/B _2664_/A vdd gnd INVX1
X_1437_ _1698_/Q _1481_/A vdd gnd INVX1
X_1506_ _3000_/A _1508_/B vdd gnd INVX1
X_2486_ _2509_/B _2511_/B _2518_/D vdd gnd NOR2X1
X_2555_ _2555_/A _2583_/B _2555_/C _2555_/D _3022_/D vdd gnd OAI22X1
X_3107_ _3107_/A y[4] vdd gnd BUFX2
X_3038_ _3038_/D _3075_/CLK _3038_/Q vdd gnd DFFPOSX1
X_2271_ _2271_/A _2443_/Q _2272_/A vdd gnd NOR2X1
X_2340_ _2340_/A _2341_/B vdd gnd INVX1
X_1986_ _2117_/A _2063_/A vdd gnd INVX1
X_2607_ _3032_/Q _2616_/B vdd gnd INVX1
X_2469_ _2469_/D _2469_/CLK _2469_/Q vdd gnd DFFPOSX1
X_2538_ _2743_/B _2667_/B vdd gnd INVX4
X_1840_ _2070_/A _2080_/A _1876_/A _1841_/A vdd gnd OAI21X1
X_1771_ vdd _3090_/Q _1772_/C vdd gnd NAND2X1
X_2254_ _2263_/A _2264_/C vdd gnd INVX1
X_2323_ _2462_/Q _2332_/B vdd gnd INVX1
X_2185_ _2185_/A _2185_/B _2187_/B vdd gnd NOR2X1
X_1969_ _1969_/A _1969_/B _1969_/C _1976_/C vdd gnd AOI21X1
X_1823_ _1861_/A _1826_/C _1824_/C vdd gnd NAND2X1
X_2941_ _2948_/A _3074_/Q _2942_/C vdd gnd NAND2X1
X_2872_ _3081_/Q _2887_/B _2876_/C _2874_/C vdd gnd NAND3X1
X_1685_ _1685_/D _2462_/CLK _1685_/Q vdd gnd DFFPOSX1
X_1754_ vdd _2233_/A _1754_/C _2431_/D vdd gnd OAI21X1
X_2237_ _2238_/B _2238_/A _2239_/B vdd gnd OR2X2
X_2306_ _2313_/A _2306_/B _2314_/B vdd gnd NOR2X1
X_2099_ _2144_/A _2143_/A _2144_/B _2110_/A vdd gnd NAND3X1
X_2168_ _2451_/Q _2375_/B vdd gnd INVX1
X_1470_ _1477_/B _1470_/B _1484_/B _3106_/A vdd gnd OAI21X1
X_3071_ _3071_/D _3097_/CLK _3071_/Q vdd gnd DFFPOSX1
X_2022_ _2075_/A _2088_/A vdd gnd INVX1
X_1806_ _2270_/B vdd _1806_/C _2443_/D vdd gnd OAI21X1
X_2924_ _2960_/A _2924_/B _2924_/C _2925_/B vdd gnd OAI21X1
X_2855_ _2879_/A _2879_/B _2888_/A vdd gnd NOR2X1
X_2786_ _2856_/B _2989_/A _2816_/B vdd gnd NAND2X1
X_1599_ _1655_/B _1655_/A _2292_/A vdd gnd NAND2X1
X_1668_ rst _1668_/B _1700_/D vdd gnd NOR2X1
X_1737_ _1737_/A _1737_/B _1737_/C _1739_/D vdd gnd OAI21X1
X_2640_ _2640_/A _2640_/B _2667_/B _2641_/C vdd gnd MUX2X1
X_1453_ _1461_/C _1453_/B _1484_/B _3103_/A vdd gnd OAI21X1
X_1522_ _1522_/A x[7] _1523_/C vdd gnd NAND2X1
X_2571_ _2571_/A _2583_/B _2571_/C _2571_/D _3026_/D vdd gnd OAI22X1
X_2005_ _2428_/Q _2439_/Q _2122_/A vdd gnd AND2X2
X_3054_ _3054_/D _3075_/CLK _3054_/Q vdd gnd DFFPOSX1
X_2907_ _2907_/A _2979_/B _2986_/A _2914_/D vdd gnd AOI21X1
X_2838_ _2838_/A _2838_/B _2838_/C _3073_/D vdd gnd OAI21X1
X_2769_ _2769_/A _2769_/B _2769_/C _3058_/D vdd gnd OAI21X1
X_2554_ _2992_/A _2582_/B _2583_/B _2555_/D vdd gnd OAI21X1
X_2623_ _2743_/A _2623_/B _2623_/C _2626_/C vdd gnd AOI21X1
X_1436_ _1436_/A _1436_/B _1461_/C vdd gnd NOR2X1
X_1505_ _1517_/A _1505_/B _1505_/C _1564_/D vdd gnd OAI21X1
X_2485_ _2508_/A _2508_/B _2511_/B vdd gnd NAND2X1
X_3106_ _3106_/A y[3] vdd gnd BUFX2
X_3037_ _3037_/D _3061_/CLK _3037_/Q vdd gnd DFFPOSX1
X_2270_ _2270_/A _2270_/B _2278_/C vdd gnd NOR2X1
X_1985_ _1992_/A _1985_/B _2117_/A vdd gnd NAND2X1
X_2537_ _2743_/A _2602_/B vdd gnd INVX1
X_2606_ _2665_/A _2606_/B _2606_/C _2606_/D _3031_/D vdd gnd AOI22X1
X_2399_ _2413_/B _2415_/B vdd _2400_/A vdd gnd OAI21X1
X_2468_ _2468_/D _2470_/CLK _2468_/Q vdd gnd DFFPOSX1
X_1770_ _2437_/Q _2130_/A vdd gnd INVX1
X_2184_ _2185_/A _2185_/B _2184_/C _2212_/A vdd gnd OAI21X1
X_2253_ _2255_/A _2255_/B _2263_/A vdd gnd NOR2X1
X_2322_ _2322_/A _2322_/B _2322_/C _2461_/D vdd gnd OAI21X1
X_1899_ _2433_/Q _2432_/Q _1899_/C _1902_/B vdd gnd NAND3X1
X_1968_ _1968_/A _1969_/C vdd gnd INVX1
X_2940_ _3058_/Q _2942_/B vdd gnd INVX1
X_1753_ vdd _1753_/B _1754_/C vdd gnd NAND2X1
X_1822_ _1851_/A _1834_/C _1822_/C _1861_/A vdd gnd NAND3X1
X_2871_ _3004_/A _2887_/B _2888_/A _2874_/B vdd gnd NAND3X1
X_1684_ _1684_/D _2462_/CLK _1684_/Q vdd gnd DFFPOSX1
X_2167_ _2352_/B vdd _2167_/C _2450_/D vdd gnd OAI21X1
X_2236_ _2247_/A _2236_/B _2238_/B vdd gnd AND2X2
X_2305_ _2305_/A _2446_/Q _2313_/A vdd gnd NOR2X1
X_2098_ _2110_/C _2104_/C vdd gnd INVX1
X_2021_ _2030_/B _2030_/C _2075_/A _2035_/B vdd gnd AOI21X1
X_3070_ _3070_/D _3098_/CLK _3070_/Q vdd gnd DFFPOSX1
X_2923_ _2960_/A _3048_/Q _2924_/C vdd gnd NAND2X1
X_1736_ _1736_/A rst _1737_/C vdd gnd NOR2X1
X_1805_ vdd _1805_/B _1806_/C vdd gnd NAND2X1
X_2854_ _2854_/A _2854_/B _2854_/C _3077_/D vdd gnd OAI21X1
X_2785_ _2785_/A _2982_/S _2989_/A vdd gnd NOR2X1
X_1598_ _1607_/A _2459_/Q _1655_/B vdd gnd NAND2X1
X_1667_ rst _1667_/B _1699_/D vdd gnd NOR2X1
X_2219_ _2229_/A _2225_/A vdd gnd INVX1
X_2570_ _3008_/A _2582_/B _2583_/B _2571_/D vdd gnd OAI21X1
X_1452_ _1452_/A _1688_/Q _1689_/Q _1453_/B vdd gnd AOI21X1
X_1521_ _3020_/A _1523_/B vdd gnd INVX1
X_2004_ _2012_/A _2009_/B vdd gnd INVX1
X_3053_ _3053_/D _3101_/CLK _3053_/Q vdd gnd DFFPOSX1
X_2906_ _2984_/A _2906_/B _2906_/C _2907_/A vdd gnd OAI21X1
X_1719_ _1723_/B _1719_/B _1724_/A _1721_/C vdd gnd AOI21X1
X_2699_ _3016_/A _2703_/B _2704_/B _2700_/D vdd gnd OAI21X1
X_2837_ _3004_/A _2853_/B _2853_/C _2838_/A vdd gnd OAI21X1
X_2768_ _2780_/A _3008_/A _2780_/C _2769_/B vdd gnd AOI21X1
X_1504_ _1519_/A x[1] _1505_/C vdd gnd NAND2X1
X_2553_ _2860_/B _2991_/B _2582_/B vdd gnd NOR2X1
X_2622_ _2988_/A _2622_/B _2622_/C _2662_/D _2623_/C vdd gnd OAI22X1
X_1435_ _1688_/Q _1689_/Q _1436_/B vdd gnd NAND2X1
X_2484_ _2522_/Q _2530_/Y _2521_/Q _2508_/B vdd gnd NOR3X1
X_3105_ _3105_/A y[2] vdd gnd BUFX2
X_3036_ _3036_/D _3101_/CLK _3036_/Q vdd gnd DFFPOSX1
X_1984_ _1984_/A _1984_/B _1984_/C _1992_/A vdd gnd NAND3X1
X_2467_ _2467_/D _2470_/CLK _2467_/Q vdd gnd DFFPOSX1
X_2536_ _3022_/Q _2555_/A vdd gnd INVX1
X_2605_ _2665_/A _2605_/B _2606_/C vdd gnd NOR2X1
X_2398_ _2398_/A _2413_/B vdd gnd INVX1
X_3019_ _3037_/Q _3019_/B _3021_/C vdd gnd NOR2X1
X_2321_ _2341_/A _2324_/B vdd _2322_/A vdd gnd OAI21X1
X_2183_ _2186_/B _2186_/A _2184_/C vdd gnd AND2X2
X_2252_ _2252_/A _2255_/A vdd gnd INVX1
X_1898_ _2434_/Q _2431_/Q _1898_/C _1902_/A vdd gnd NAND3X1
X_1967_ _1976_/A _1976_/B _2048_/C _1983_/B vdd gnd OAI21X1
X_2519_ _2519_/D _3087_/CLK _2519_/Q vdd gnd DFFPOSX1
X_2870_ _2870_/A _2870_/B _2870_/C _3080_/D vdd gnd NAND3X1
X_1683_ _1683_/D _2462_/CLK _1683_/Q vdd gnd DFFPOSX1
X_1752_ _2431_/Q _2233_/A vdd gnd INVX2
X_1821_ _2433_/Q _2430_/Q _1851_/A vdd gnd AND2X2
X_2304_ _2313_/C _2306_/B vdd gnd INVX1
X_2097_ _2104_/A _2104_/B _2110_/C _2102_/A vdd gnd OAI21X1
X_2166_ _2166_/A _2166_/B vdd _2167_/C vdd gnd OAI21X1
X_2235_ _2235_/A _2235_/B _2247_/A vdd gnd OR2X2
X_2999_ _3032_/Q _3019_/B _3001_/C vdd gnd NOR2X1
X_2020_ _2233_/A _2080_/A _2087_/A _2030_/C vdd gnd OAI21X1
X_2922_ _2922_/A _2922_/B _2982_/S _2925_/C vdd gnd MUX2X1
X_2853_ _3020_/A _2853_/B _2853_/C _2854_/A vdd gnd OAI21X1
X_1666_ _1666_/A _1666_/B _1666_/C _1698_/D vdd gnd AOI21X1
X_1735_ _1735_/A _1735_/B rst _1738_/D vdd gnd AOI21X1
X_1804_ _1804_/A _1828_/A _1805_/B vdd gnd NOR2X1
X_2784_ _2819_/B _2988_/A _2860_/A _2991_/A _2818_/B vdd gnd OAI22X1
X_1597_ _1687_/Q _1630_/B _1655_/A vdd gnd NAND2X1
X_2149_ _2156_/A _2155_/A vdd gnd INVX1
X_2218_ _2229_/A _2230_/A _2218_/C _2226_/B vdd gnd NAND3X1
X_1520_ _1536_/B _1520_/B _1520_/C _1569_/D vdd gnd OAI21X1
X_1451_ _1481_/A _1464_/A _1451_/C _1484_/B vdd gnd NAND3X1
X_2003_ _2427_/Q _2440_/Q _2012_/A vdd gnd NAND2X1
X_3052_ _3052_/D _3061_/CLK _3052_/Q vdd gnd DFFPOSX1
X_2905_ _2984_/A _3071_/Q _2906_/C vdd gnd NAND2X1
X_2836_ _3033_/Q _2852_/B _2838_/B vdd gnd NOR2X1
X_1649_ _1678_/Q _1649_/B _1649_/C _1650_/A vdd gnd NAND3X1
X_1718_ _1747_/B _1721_/B vdd gnd INVX1
X_2698_ _3036_/Q _2702_/B _2700_/C vdd gnd NOR2X1
X_2767_ _3034_/Q _2779_/B _2769_/A vdd gnd NOR2X1
X_1503_ _2996_/A _1505_/B vdd gnd INVX1
X_2483_ _2502_/A _2515_/D vdd gnd INVX1
X_2552_ _3030_/Q _2581_/B _2555_/C vdd gnd NOR2X1
X_2621_ _3065_/Q _3097_/Q _2633_/S _2622_/B vdd gnd MUX2X1
X_1434_ _1686_/Q _1687_/Q _1436_/A vdd gnd NAND2X1
X_3104_ _3104_/A y[1] vdd gnd BUFX2
X_3035_ _3035_/D _3099_/CLK _3035_/Q vdd gnd DFFPOSX1
X_2819_ _2819_/A _2819_/B _2860_/A _2822_/A _2853_/C vdd gnd OAI22X1
X_1983_ _2049_/A _1983_/B _1983_/C _1984_/C vdd gnd NAND3X1
X_2604_ _2604_/A _2879_/B _2988_/A _2604_/D _2605_/B vdd gnd OAI22X1
X_2466_ _2466_/D _2470_/CLK _2466_/Q vdd gnd DFFPOSX1
X_2535_ _2535_/D _2535_/CLK _2535_/Q vdd gnd DFFPOSX1
X_2397_ _2398_/A _2397_/B _2400_/B vdd gnd NOR2X1
X_3018_ _3101_/Q _3021_/A vdd gnd INVX1
X_2251_ _2251_/A _2358_/A _2251_/C _2251_/D _2454_/D vdd gnd AOI22X1
X_2320_ _2324_/B _2341_/A _2322_/B vdd gnd AND2X2
X_2182_ _2203_/A _2203_/B _2182_/C _2186_/B vdd gnd NAND3X1
X_1966_ _2039_/B _2038_/A _2039_/A _1976_/B vdd gnd AOI21X1
X_1897_ _2433_/Q _2432_/Q _1898_/C vdd gnd NAND2X1
X_2449_ _2449_/D _2469_/CLK _2449_/Q vdd gnd DFFPOSX1
X_2518_ _2518_/D _3087_/CLK _2518_/Q vdd gnd DFFPOSX1
X_1820_ _1895_/A _2179_/A _1820_/C _1826_/C vdd gnd OAI21X1
X_1682_ _1682_/D _3061_/CLK _1682_/Q vdd gnd DFFPOSX1
X_1751_ vdd _2179_/A _1751_/C _2430_/D vdd gnd OAI21X1
X_2234_ _2234_/A _2234_/B _2235_/B _2236_/B vdd gnd OAI21X1
X_2303_ _2305_/A _2446_/Q _2313_/C vdd gnd NAND2X1
X_2096_ _2144_/B _2143_/A _2144_/A _2104_/B vdd gnd AOI21X1
X_2165_ _2220_/B _2165_/B _2166_/B vdd gnd NOR2X1
X_1949_ _2435_/Q _2431_/Q _2015_/A _1960_/B vdd gnd NAND3X1
X_2998_ _3096_/Q _3001_/A vdd gnd INVX1
X_1803_ _1824_/B _1803_/B _1803_/C _1804_/A vdd gnd AOI21X1
X_2921_ _3080_/Q _3024_/Q _2956_/S _2922_/A vdd gnd MUX2X1
X_2852_ _3037_/Q _2852_/B _2854_/B vdd gnd NOR2X1
X_2783_ _2783_/A _2985_/D _2991_/A vdd gnd NAND2X1
X_1596_ _1654_/B _1654_/A _2282_/A vdd gnd NAND2X1
X_1665_ _1665_/A _1665_/B _1665_/C _1697_/D vdd gnd AOI21X1
X_1734_ _1734_/A _1737_/A _1734_/Y vdd gnd NOR2X1
X_2217_ _2217_/A _2229_/C _2230_/A vdd gnd NAND2X1
X_2079_ _2431_/Q _2437_/Q _2131_/A vdd gnd NAND2X1
X_2148_ _2156_/A _2194_/A _2155_/C _2163_/A vdd gnd NAND3X1
X_1450_ _1696_/Q _1695_/Q _1697_/Q _1464_/A vdd gnd AOI21X1
X_3051_ _3051_/D _3075_/CLK _3051_/Q vdd gnd DFFPOSX1
X_2002_ _2002_/A _2002_/B _2038_/A _2044_/A vdd gnd OAI21X1
X_2904_ _3055_/Q _2906_/B vdd gnd INVX1
X_2835_ _3073_/Q _2851_/B _2838_/C vdd gnd NAND2X1
X_2766_ _3058_/Q _2779_/B _2778_/C _2769_/C vdd gnd NAND3X1
X_1579_ _1670_/B _1679_/Q _1648_/A vdd gnd AND2X2
X_1648_ _1648_/A _1649_/B vdd gnd INVX1
X_1717_ _1717_/A _1717_/B _1717_/C _1726_/D vdd gnd OAI21X1
X_2697_ _3044_/Q _2972_/B vdd gnd INVX1
X_2620_ _2620_/A _2620_/B _2667_/B _2623_/B vdd gnd MUX2X1
X_1502_ _1519_/A _1502_/B _1502_/C _1563_/D vdd gnd OAI21X1
X_2482_ _2530_/Y _2521_/Q _2502_/A vdd gnd NOR2X1
X_2551_ _2856_/A _2989_/B _2581_/B vdd gnd NAND2X1
X_3103_ _3103_/A y[0] vdd gnd BUFX2
X_3034_ _3034_/D _3098_/CLK _3034_/Q vdd gnd DFFPOSX1
X_2749_ _3030_/Q _2779_/B _2753_/A vdd gnd NOR2X1
X_2818_ _2818_/A _2818_/B _2818_/C _2818_/D _3069_/D vdd gnd OAI22X1
X_1982_ _1996_/A _2049_/A vdd gnd INVX1
X_2534_ _2534_/D _3093_/CLK _2534_/Q vdd gnd DFFPOSX1
X_2603_ _3063_/Q _3095_/Q _2706_/A _2604_/D vdd gnd MUX2X1
X_2396_ _2403_/A _2412_/B _2398_/A vdd gnd NOR2X1
X_2465_ _2465_/D _2470_/CLK _2465_/Q vdd gnd DFFPOSX1
X_3017_ _3017_/A _3021_/B _3017_/C _3017_/D _3100_/D vdd gnd OAI22X1
X_2250_ _2250_/A _2250_/B _2251_/D vdd gnd AND2X2
X_2181_ _2203_/C _2182_/C vdd gnd INVX1
X_1965_ _1965_/A _1965_/B _1965_/C _2039_/B vdd gnd OAI21X1
X_1896_ _1958_/D _1958_/C _1946_/C _1931_/A vdd gnd NAND3X1
X_2517_ _2517_/D _2535_/CLK _2517_/Q vdd gnd DFFPOSX1
X_2379_ _2385_/B _2381_/B vdd gnd INVX1
X_2448_ _2448_/D _2469_/CLK _2448_/Q vdd gnd DFFPOSX1
X_1750_ vdd _1750_/B _1751_/C vdd gnd NAND2X1
X_1681_ _1681_/D _3061_/CLK _1682_/D vdd gnd DFFPOSX1
X_2164_ _2171_/C _2164_/B _2220_/B vdd gnd NAND2X1
X_2233_ _2233_/A _2233_/B _2233_/C _2235_/B vdd gnd OAI21X1
X_2302_ _2343_/C _2314_/A _2312_/A _2308_/A vdd gnd AOI21X1
X_2095_ _2095_/A _2095_/B _2095_/C _2144_/B vdd gnd OAI21X1
X_1879_ _2428_/Q _2437_/Q _1880_/B vdd gnd AND2X2
X_1948_ _2434_/Q _2432_/Q _2015_/A vdd gnd NAND2X1
X_2997_ _2997_/A _3021_/B _2997_/C _2997_/D _3095_/D vdd gnd OAI22X1
X_2920_ _3064_/Q _3096_/Q _2956_/S _2922_/B vdd gnd MUX2X1
X_1733_ _1739_/Q _1737_/A vdd gnd INVX1
X_1802_ _1802_/A _1828_/A vdd gnd INVX1
X_2851_ _3077_/Q _2851_/B _2854_/C vdd gnd NAND2X1
X_2782_ _3062_/Q _2790_/A vdd gnd INVX1
X_1595_ _1607_/A _2458_/Q _1654_/B vdd gnd NAND2X1
X_1664_ _1664_/A _1664_/B _1666_/C _1696_/D vdd gnd AOI21X1
X_2147_ _2150_/A _2150_/B _2151_/C _2155_/C vdd gnd OAI21X1
X_2216_ _2216_/A _2216_/B _2229_/C vdd gnd NAND2X1
X_2078_ _2437_/Q _2432_/Q _2173_/A vdd gnd NAND2X1
X_2001_ _2001_/A _2001_/B _2001_/C _2002_/B vdd gnd AOI21X1
X_3050_ _3050_/D _3075_/CLK _3050_/Q vdd gnd DFFPOSX1
X_2903_ _3087_/Q _2914_/B vdd gnd INVX1
X_1716_ _1720_/A _1720_/B _1737_/B _1717_/A vdd gnd OAI21X1
X_2696_ _2960_/B _2704_/B _2696_/C _2696_/D _3043_/D vdd gnd OAI22X1
X_2834_ _2834_/A _2834_/B _2834_/C _3072_/D vdd gnd OAI21X1
X_2765_ _2765_/A _2765_/B _2765_/C _3057_/D vdd gnd OAI21X1
X_1578_ _1676_/Q _1670_/B _1640_/B vdd gnd NAND2X1
X_1647_ _1670_/C _1647_/B _1648_/A _1650_/B vdd gnd OAI21X1
X_2550_ _2957_/S _2550_/B _2989_/B vdd gnd NOR2X1
X_1501_ _1519_/A x[0] _1502_/C vdd gnd NAND2X1
X_2481_ _2481_/A _2481_/Y vdd gnd INVX1
X_3102_ _3102_/A ready vdd gnd BUFX2
X_3033_ _3033_/D _3097_/CLK _3033_/Q vdd gnd DFFPOSX1
X_2679_ _2996_/A _2703_/B _2704_/B _2680_/D vdd gnd OAI21X1
X_2748_ _3054_/Q _2779_/B _2778_/C _2753_/C vdd gnd NAND3X1
X_2817_ _3020_/A _2817_/B _2818_/B _2818_/C vdd gnd OAI21X1
X_1981_ _1996_/A _2049_/C _1996_/B _1984_/B vdd gnd NAND3X1
X_2533_ _2533_/A _2533_/B _2533_/C _2535_/D vdd gnd OAI21X1
X_2602_ _2743_/B _2602_/B _2988_/A vdd gnd NAND2X1
X_2395_ _2395_/A _2453_/Q _2403_/A vdd gnd NOR2X1
X_2464_ _2464_/D _2469_/CLK _2464_/Q vdd gnd DFFPOSX1
X_3016_ _3016_/A _3020_/B _3021_/B _3017_/D vdd gnd OAI21X1
X_2180_ _2180_/A _2206_/C _2203_/C vdd gnd NOR2X1
X_1895_ _1895_/A _2204_/A _1899_/C _1958_/C vdd gnd OAI21X1
X_1964_ _2001_/C _2001_/B _2001_/A _2038_/A vdd gnd NAND3X1
X_2447_ _2447_/D _2469_/CLK _2447_/Q vdd gnd DFFPOSX1
X_2516_ _2516_/D _3093_/CLK _2516_/Q vdd gnd DFFPOSX1
X_2378_ _2378_/A _2384_/C _2385_/B vdd gnd NOR2X1
X_1680_ _1682_/Q _3061_/CLK _1680_/Q vdd gnd DFFPOSX1
X_2301_ _2460_/Q _2310_/B vdd gnd INVX1
X_2163_ _2163_/A _2163_/B _2163_/C _2164_/B vdd gnd NAND3X1
X_2232_ _2232_/A _2232_/B _2232_/C _2241_/B vdd gnd NAND3X1
X_2094_ _2123_/B _2123_/C _2123_/A _2143_/A vdd gnd NAND3X1
X_1878_ _1887_/A _1883_/B vdd gnd INVX1
X_1947_ _2430_/Q _2436_/Q _2016_/A vdd gnd NAND2X1
X_2996_ _2996_/A _3020_/B _3021_/B _2997_/D vdd gnd OAI21X1
X_2850_ _2850_/A _2850_/B _2850_/C _3076_/D vdd gnd OAI21X1
X_1663_ _1663_/A _1663_/B _1666_/C _1695_/D vdd gnd AOI21X1
X_1732_ _1735_/B _1735_/A _1732_/Y vdd gnd NAND2X1
X_1801_ _1803_/C _1803_/B _1824_/B _1802_/A vdd gnd NAND3X1
X_2781_ _2781_/A _2781_/B _2781_/C _3061_/D vdd gnd OAI21X1
X_1594_ _1686_/Q _1630_/B _1654_/A vdd gnd NAND2X1
X_2077_ _2125_/C _2082_/A vdd gnd INVX1
X_2146_ _2190_/A _2146_/B _2146_/C _2150_/B vdd gnd AOI21X1
X_2215_ _2238_/A _2215_/B _2216_/A vdd gnd NOR2X1
X_2979_ _2979_/A _2979_/B _2986_/A _2986_/D vdd gnd AOI21X1
X_2000_ _2050_/A _2051_/A vdd gnd INVX1
X_2902_ _2986_/A _2902_/B _2902_/C _2902_/D _3086_/D vdd gnd AOI22X1
X_2833_ _3000_/A _2853_/B _2853_/C _2834_/A vdd gnd OAI21X1
X_1646_ _1678_/Q _1670_/C vdd gnd INVX1
X_1715_ _1715_/A _1719_/B _1724_/D _1717_/B vdd gnd OAI21X1
X_2695_ _3012_/A _2703_/B _2704_/B _2696_/D vdd gnd OAI21X1
X_2764_ _2780_/A _3004_/A _2780_/C _2765_/B vdd gnd AOI21X1
X_1577_ _1645_/B _1719_/B vdd gnd INVX1
X_2129_ _2431_/Q _2438_/Q _2180_/A vdd gnd NAND2X1
X_1500_ _2992_/A _1502_/B vdd gnd INVX1
X_2480_ _2533_/B _2509_/B _2481_/A vdd gnd NAND2X1
X_3101_ _3101_/D _3101_/CLK _3101_/Q vdd gnd DFFPOSX1
X_3032_ _3032_/D _3099_/CLK _3032_/Q vdd gnd DFFPOSX1
X_2816_ _3037_/Q _2816_/B _2818_/D vdd gnd NOR2X1
X_1629_ _1665_/B _1665_/A _2422_/A vdd gnd NAND2X1
X_2678_ _3031_/Q _2702_/B _2680_/C vdd gnd NOR2X1
X_2747_ _2979_/B _2989_/B _2779_/B vdd gnd NAND2X1
X_1980_ _1980_/A _1980_/B _1980_/C _1984_/A vdd gnd OAI21X1
X_2463_ _2463_/D _2470_/CLK _2463_/Q vdd gnd DFFPOSX1
X_2532_ _2532_/A rst _2533_/C vdd gnd NOR2X1
X_2601_ _2706_/A _2602_/B _2667_/B _2879_/B vdd gnd NAND3X1
X_2394_ _2394_/A _2394_/B _2412_/B vdd gnd NOR2X1
X_3015_ _3036_/Q _3019_/B _3017_/C vdd gnd NOR2X1
X_1894_ _2434_/Q _2431_/Q _1899_/C vdd gnd NAND2X1
X_1963_ _1963_/A _1999_/C _2039_/A vdd gnd AND2X2
X_2446_ _2446_/D _2469_/CLK _2446_/Q vdd gnd DFFPOSX1
X_2515_ _2515_/D _2535_/CLK _2515_/Q vdd gnd DFFPOSX1
X_2377_ _2377_/A _2452_/Q _2378_/A vdd gnd NOR2X1
X_2231_ _2232_/B _2231_/B _2231_/C _2241_/A vdd gnd AOI21X1
X_2300_ _2332_/A _2300_/B _2300_/C _2459_/D vdd gnd OAI21X1
X_2093_ _2124_/A _2144_/A vdd gnd INVX1
X_2162_ _2162_/A _2163_/C vdd gnd INVX1
X_2995_ _3031_/Q _3019_/B _2997_/C vdd gnd NOR2X1
X_1877_ _2427_/Q _2438_/Q _1887_/A vdd gnd NAND2X1
X_1946_ _1946_/A _1946_/B _1946_/C _2001_/C vdd gnd OAI21X1
X_2429_ _2429_/D _3087_/CLK _2429_/Q vdd gnd DFFPOSX1
X_1800_ _1800_/A _2025_/A _1825_/B _1803_/B vdd gnd OAI21X1
X_1662_ _1662_/A _1662_/B _1665_/C _1694_/D vdd gnd AOI21X1
X_1731_ _1738_/Q _1734_/A _1735_/A vdd gnd NAND2X1
X_2780_ _2780_/A _3020_/A _2780_/C _2781_/B vdd gnd AOI21X1
X_1593_ _1653_/B _1653_/A _2271_/A vdd gnd NAND2X1
X_2214_ _2214_/A _2216_/B vdd gnd INVX1
X_2076_ _2179_/A _2176_/B _2125_/C vdd gnd NOR2X1
X_2145_ _2145_/A _2145_/B _2145_/C _2150_/A vdd gnd AOI21X1
X_1929_ _1980_/C _1930_/C vdd gnd INVX1
X_2978_ _2980_/S _2978_/B _2978_/C _2979_/A vdd gnd OAI21X1
X_2763_ _3033_/Q _2779_/B _2765_/A vdd gnd NOR2X1
X_2901_ _2985_/A _2901_/B _2901_/C _2985_/D _2902_/C vdd gnd AOI22X1
X_2832_ _3032_/Q _2852_/B _2834_/B vdd gnd NOR2X1
X_1576_ _1678_/Q _1670_/B _1645_/B vdd gnd NAND2X1
X_1645_ _1678_/Q _1645_/B _1649_/C _1678_/D vdd gnd MUX2X1
X_1714_ _1715_/A _1720_/A _1724_/D vdd gnd NAND2X1
X_2694_ _3035_/Q _2702_/B _2696_/C vdd gnd NOR2X1
X_2059_ _2358_/A _2059_/B _2059_/C _2448_/D vdd gnd OAI21X1
X_2128_ _2432_/Q _2438_/Q _2131_/B vdd gnd NAND2X1
X_3100_ _3100_/D _3101_/CLK _3100_/Q vdd gnd DFFPOSX1
X_3031_ _3031_/D _3097_/CLK _3031_/Q vdd gnd DFFPOSX1
X_2746_ _2822_/A _2979_/B vdd gnd INVX2
X_2815_ _3069_/Q _2818_/A vdd gnd INVX1
X_1559_ _1559_/D _3093_/CLK _1559_/Q vdd gnd DFFPOSX1
X_1628_ _1631_/A _2469_/Q _1665_/B vdd gnd NAND2X1
X_2677_ _3039_/Q _2912_/B vdd gnd INVX1
X_2600_ _3079_/Q _2604_/A vdd gnd INVX1
X_2393_ _2453_/Q _2394_/B vdd gnd INVX1
X_2462_ _2462_/D _2462_/CLK _2462_/Q vdd gnd DFFPOSX1
X_2531_ _2531_/A _2531_/B rst _2534_/D vdd gnd AOI21X1
X_3014_ _3100_/Q _3017_/A vdd gnd INVX1
X_2729_ _3008_/A _2741_/B _2742_/B _2730_/C vdd gnd OAI21X1
X_1962_ _1971_/C _1971_/B _2002_/A _1976_/A vdd gnd AOI21X1
X_1893_ _1958_/A _1958_/B _1946_/C vdd gnd NAND2X1
X_2376_ _2377_/A _2452_/Q _2384_/C vdd gnd AND2X2
X_2445_ _2445_/D _2469_/CLK _2445_/Q vdd gnd DFFPOSX1
X_2514_ _2532_/A _2514_/B _2520_/D vdd gnd AND2X2
X_2230_ _2230_/A _2230_/B _2232_/B vdd gnd NOR2X1
X_2092_ _2100_/C _2100_/B _2124_/A _2104_/A vdd gnd AOI21X1
X_2161_ _2162_/A _2194_/B _2161_/C _2171_/C vdd gnd NAND3X1
X_1945_ _2433_/Q _2432_/Q _2434_/Q _2431_/Q _1946_/B vdd gnd AOI22X1
X_2994_ _3095_/Q _2997_/A vdd gnd INVX1
X_1876_ _1876_/A _1974_/A _1876_/C _1930_/A vdd gnd OAI21X1
X_2359_ _2465_/Q _2382_/A _2373_/C vdd gnd NAND2X1
X_2428_ _2428_/D _2535_/CLK _2428_/Q vdd gnd DFFPOSX1
X_1592_ _1607_/A _2457_/Q _1653_/B vdd gnd NAND2X1
X_1661_ _1661_/A _1661_/B _1665_/C _1693_/D vdd gnd AOI21X1
X_1730_ _1737_/B _1734_/A vdd gnd INVX1
X_2144_ _2144_/A _2144_/B _2144_/C _2151_/C vdd gnd AOI21X1
X_2213_ _2215_/B _2238_/A _2214_/A _2217_/A vdd gnd OAI21X1
X_2075_ _2075_/A _2075_/B _2075_/C _2123_/C vdd gnd OAI21X1
X_1859_ _1859_/A _1862_/A vdd gnd INVX1
X_1928_ _1928_/A _1928_/B _2063_/C vdd gnd NAND2X1
X_2977_ _2980_/S _3077_/Q _2978_/C vdd gnd NAND2X1
X_2900_ _2956_/S _2900_/B _2900_/C _2901_/B vdd gnd OAI21X1
X_1713_ _1756_/B _1724_/A _1717_/C vdd gnd NAND2X1
X_2762_ _3057_/Q _2779_/B _2778_/C _2765_/C vdd gnd NAND3X1
X_2831_ _3072_/Q _2851_/B _2834_/C vdd gnd NAND2X1
X_1575_ _1669_/C _1723_/B vdd gnd INVX1
X_1644_ _1644_/A _1644_/B _1649_/C vdd gnd NOR2X1
X_2693_ _3043_/Q _2960_/B vdd gnd INVX1
X_2127_ _2430_/Q _2439_/Q _2136_/B vdd gnd NAND2X1
X_2058_ _2448_/Q _2358_/A _2059_/C vdd gnd NAND2X1
X_3030_ _3030_/D _3098_/CLK _3030_/Q vdd gnd DFFPOSX1
X_2676_ _2900_/B _2704_/B _2676_/C _2676_/D _3038_/D vdd gnd OAI22X1
X_2745_ _2785_/A _2783_/A _2822_/A vdd gnd NAND2X1
X_2814_ _2814_/A _2818_/B _2814_/C _2814_/D _3068_/D vdd gnd OAI22X1
X_1489_ _1559_/Q _1715_/A _1490_/C vdd gnd NAND2X1
X_1558_ _1558_/D _3093_/CLK _1558_/Q vdd gnd DFFPOSX1
X_1627_ _1697_/Q _1630_/B _1665_/A vdd gnd NAND2X1
X_2530_ _2530_/A _2533_/A _2530_/Y vdd gnd NOR2X1
X_2392_ _2395_/A _2394_/A vdd gnd INVX1
X_2461_ _2461_/D _2462_/CLK _2461_/Q vdd gnd DFFPOSX1
X_3013_ _3013_/A _3021_/B _3013_/C _3013_/D _3099_/D vdd gnd OAI22X1
X_2659_ _3053_/Q _3045_/Q _2661_/S _2660_/A vdd gnd MUX2X1
X_2728_ _3034_/Q _2740_/B _2730_/D vdd gnd NOR2X1
X_1892_ _2434_/Q _2432_/Q _1958_/B vdd gnd AND2X2
X_1961_ _2001_/B _1965_/C _2001_/A _1971_/B vdd gnd NAND3X1
X_2513_ vdd rst _2514_/B vdd gnd NOR2X1
X_2375_ _2375_/A _2375_/B _2375_/C _2381_/A vdd gnd OAI21X1
X_2444_ _2444_/D _3095_/CLK _2444_/Q vdd gnd DFFPOSX1
X_2160_ _2171_/A _2160_/B _2165_/B vdd gnd NAND2X1
X_2091_ _2123_/B _2095_/C _2123_/A _2100_/B vdd gnd NAND3X1
X_1875_ _1988_/A _1988_/B _1918_/A vdd gnd NAND2X1
X_1944_ _1999_/C _1963_/A _2002_/A vdd gnd NAND2X1
X_2993_ _2993_/A _3021_/B _2993_/C _2993_/D _3094_/D vdd gnd OAI22X1
X_2427_ _2427_/D _3087_/CLK _2427_/Q vdd gnd DFFPOSX1
X_2289_ _2459_/Q _2332_/A _2300_/C vdd gnd NAND2X1
X_2358_ _2358_/A _2358_/B _2358_/C _2358_/D _2464_/D vdd gnd AOI22X1
X_1591_ _1685_/Q _1630_/B _1653_/A vdd gnd NAND2X1
X_1660_ _1660_/A _1660_/B _1665_/C _1692_/D vdd gnd AOI21X1
X_2143_ _2143_/A _2144_/C vdd gnd INVX1
X_2212_ _2212_/A _2212_/B _2238_/A vdd gnd NOR2X1
X_2074_ _2087_/A _2125_/A _2075_/B vdd gnd NOR2X1
X_1858_ _1859_/A _1988_/A _1858_/C _1988_/B vdd gnd NAND3X1
X_1927_ _2447_/Q _2358_/A _1991_/C vdd gnd NAND2X1
X_2976_ _3061_/Q _2978_/B vdd gnd INVX1
X_1789_ _1803_/C _1791_/C vdd gnd INVX1
X_2830_ _2830_/A _2830_/B _2830_/C _3071_/D vdd gnd OAI21X1
X_1643_ _1676_/Q _1677_/Q _1670_/B _1644_/B vdd gnd NAND3X1
X_1712_ _1712_/A _1712_/B _1725_/D vdd gnd NAND2X1
X_2692_ _2948_/B _2704_/B _2692_/C _2692_/D _3042_/D vdd gnd OAI22X1
X_2761_ _2761_/A _2761_/B _2761_/C _3056_/D vdd gnd OAI21X1
X_1574_ _1677_/Q _1670_/B _1669_/C vdd gnd NAND2X1
X_2057_ _2057_/A _2057_/B _2059_/B vdd gnd NAND2X1
X_2126_ _2140_/A _2139_/C vdd gnd INVX1
X_2959_ _2960_/A _3051_/Q _2960_/C vdd gnd NAND2X1
X_2813_ _3016_/A _2817_/B _2818_/B _2814_/C vdd gnd OAI21X1
X_1626_ _1664_/B _1664_/A _2405_/A vdd gnd NAND2X1
X_2675_ _2992_/A _2703_/B _2704_/B _2676_/D vdd gnd OAI21X1
X_2744_ _2988_/B _2819_/A _2778_/C vdd gnd OR2X2
X_1488_ _2515_/Q _1490_/B vdd gnd INVX1
X_1557_ _1557_/D _3093_/CLK _1557_/Q vdd gnd DFFPOSX1
X_2109_ _2154_/C _2111_/B vdd gnd INVX1
X_3089_ _3089_/D _3095_/CLK _3089_/Q vdd gnd DFFPOSX1
X_2460_ _2460_/D _2462_/CLK _2460_/Q vdd gnd DFFPOSX1
X_2391_ _2415_/B _2397_/B vdd gnd INVX1
X_3012_ _3012_/A _3020_/B _3021_/B _3013_/D vdd gnd OAI21X1
X_1609_ _1691_/Q _1630_/B _1659_/A vdd gnd NAND2X1
X_2589_ _3046_/Q _3038_/Q _2643_/S _2591_/B vdd gnd MUX2X1
X_2658_ _3077_/Q _3061_/Q _2661_/S _2660_/B vdd gnd MUX2X1
X_2727_ _3050_/Q _2730_/A vdd gnd INVX1
X_1891_ _2433_/Q _2431_/Q _1958_/A vdd gnd AND2X2
X_1960_ _2016_/A _1960_/B _1960_/C _2001_/A vdd gnd NAND3X1
X_2443_ _2443_/D _3095_/CLK _2443_/Q vdd gnd DFFPOSX1
X_2512_ rst _2512_/B _2519_/D vdd gnd NOR2X1
X_2374_ _2466_/Q _2382_/B vdd gnd INVX1
X_2090_ _2179_/A _2176_/B _2090_/C _2123_/A vdd gnd OAI21X1
X_2992_ _2992_/A _3020_/B _3021_/B _2993_/D vdd gnd OAI21X1
X_1874_ _1874_/A _1874_/B _1874_/C _1989_/A vdd gnd OAI21X1
X_1943_ _1943_/A _1943_/B _1943_/C _1963_/A vdd gnd NAND3X1
X_2426_ _2426_/A _2426_/B _2426_/C _2470_/D vdd gnd OAI21X1
X_2288_ _2311_/B _2288_/B _2288_/C _2458_/D vdd gnd OAI21X1
X_2357_ _2357_/A _2360_/B _2358_/A _2358_/D vdd gnd AOI21X1
X_1590_ _1652_/B _1652_/A _2261_/A vdd gnd NAND2X1
X_2073_ _2073_/A _2145_/C _2073_/C _2124_/A vdd gnd OAI21X1
X_2142_ _2150_/C _2190_/B _2151_/B _2194_/A vdd gnd NAND3X1
X_2211_ _2212_/B _2212_/A _2215_/B vdd gnd AND2X2
X_2975_ _3093_/Q _2986_/B vdd gnd INVX1
X_1788_ _1788_/A _1808_/A _1803_/C vdd gnd NOR2X1
X_1857_ _1860_/A _1979_/C _1861_/A _1858_/C vdd gnd OAI21X1
X_1926_ _1926_/A _1926_/B _1926_/C _2446_/D vdd gnd OAI21X1
X_2409_ _2409_/A _2413_/A _2426_/A _2410_/D vdd gnd AOI21X1
X_1642_ _1647_/B _1642_/B _1677_/D vdd gnd AND2X2
X_1711_ _1737_/B _1711_/B _1711_/C _1712_/B vdd gnd NAND3X1
X_2691_ _3008_/A _2703_/B _2704_/B _2692_/D vdd gnd OAI21X1
X_2760_ _2780_/A _3000_/A _2780_/C _2761_/B vdd gnd AOI21X1
X_1573_ _1669_/A _1670_/B vdd gnd INVX2
X_2056_ _2062_/A _2056_/B _2063_/B _2057_/A vdd gnd OAI21X1
X_2125_ _2125_/A _2125_/B _2125_/C _2125_/D _2140_/A vdd gnd AOI22X1
X_1909_ _1932_/A _1909_/B _1909_/C _1979_/B vdd gnd NAND3X1
X_2958_ _2958_/A _2958_/B _2982_/S _2961_/C vdd gnd MUX2X1
X_2889_ _2889_/A _2889_/B _2889_/C _2889_/D _3085_/D vdd gnd OAI22X1
X_2743_ _2743_/A _2743_/B _2819_/A vdd gnd NAND2X1
X_2812_ _3036_/Q _2816_/B _2814_/D vdd gnd NOR2X1
X_1556_ _1556_/D _3061_/CLK _1556_/Q vdd gnd DFFPOSX1
X_1625_ _1631_/A _2468_/Q _1664_/B vdd gnd NAND2X1
X_2674_ _2712_/B _2991_/B _2703_/B vdd gnd NOR2X1
X_1487_ _1559_/Q _1487_/B _1487_/C _2890_/A vdd gnd OAI21X1
X_2039_ _2039_/A _2039_/B _2039_/C _2045_/C vdd gnd AOI21X1
X_2108_ _2108_/A _2154_/C _2108_/C _2153_/A vdd gnd NAND3X1
X_3088_ _3088_/D _3099_/CLK _3088_/Q vdd gnd DFFPOSX1
X_2390_ _2390_/A _2390_/B _2415_/B vdd gnd NOR2X1
X_3011_ _3035_/Q _3019_/B _3013_/C vdd gnd NOR2X1
X_2726_ _2726_/A _2742_/B _2726_/C _2726_/D _3049_/D vdd gnd OAI22X1
X_1539_ _1539_/A _1539_/B _1542_/C _1556_/D vdd gnd OAI21X1
X_1608_ _1658_/B _1658_/A _2327_/A vdd gnd NAND2X1
X_2588_ _2588_/A _2588_/B _2667_/B _2592_/B vdd gnd MUX2X1
X_2657_ _3037_/Q _2665_/B vdd gnd INVX1
X_1890_ _1946_/A _1958_/D vdd gnd INVX1
X_2373_ _2382_/A _2373_/B _2373_/C _2465_/D vdd gnd OAI21X1
X_2442_ _2442_/D _3095_/CLK _2442_/Q vdd gnd DFFPOSX1
X_2511_ _2511_/A _2511_/B _2511_/C _2524_/D vdd gnd OAI21X1
X_2709_ _2860_/A _2856_/B vdd gnd INVX1
X_1942_ _2070_/A _2176_/B _1942_/C _1943_/C vdd gnd OAI21X1
X_2991_ _2991_/A _2991_/B _3020_/B vdd gnd NOR2X1
X_1873_ _2446_/Q _2332_/A _1926_/C vdd gnd NAND2X1
X_2356_ _2357_/A _2360_/B _2358_/C vdd gnd OR2X2
X_2425_ _2425_/A _2425_/B _2426_/B vdd gnd NAND2X1
X_2287_ _2458_/Q _2311_/B _2288_/C vdd gnd NAND2X1
X_2210_ _2210_/A _2235_/A _2212_/B vdd gnd NAND2X1
X_2072_ _2146_/C _2145_/C vdd gnd INVX1
X_2141_ _2145_/C _2145_/B _2145_/A _2151_/B vdd gnd NAND3X1
X_1925_ vdd _1928_/B _1926_/B vdd gnd NAND2X1
X_2974_ _2986_/A _2974_/B _2974_/C _2974_/D _3092_/D vdd gnd AOI22X1
X_1787_ _2433_/Q _2428_/Q _1808_/A vdd gnd NAND2X1
X_1856_ _1876_/C _1856_/B _1856_/C _1860_/A vdd gnd AOI21X1
X_2339_ _2339_/A _2339_/B _2339_/C _2342_/C vdd gnd OAI21X1
X_2408_ _2409_/A _2413_/A _2410_/C vdd gnd OR2X2
X_1572_ _1669_/A _1669_/B _1715_/A vdd gnd NOR2X1
X_1641_ _1677_/Q _1737_/B _1715_/A _1647_/B vdd gnd NAND3X1
X_1710_ _1723_/B _1723_/A _1719_/B _1711_/C vdd gnd OAI21X1
X_2690_ _3034_/Q _2702_/B _2692_/C vdd gnd NOR2X1
X_2124_ _2124_/A _2124_/B _2143_/A _2150_/C vdd gnd OAI21X1
X_2055_ _2117_/B _2063_/B vdd gnd INVX1
X_1839_ _1839_/A _1886_/B _1841_/C vdd gnd NAND2X1
X_1908_ _1908_/A _1931_/B _1931_/A _1909_/B vdd gnd NAND3X1
X_2957_ _3083_/Q _3027_/Q _2957_/S _2958_/A vdd gnd MUX2X1
X_2888_ _2888_/A _3020_/A _2888_/C _2889_/D vdd gnd AOI21X1
X_2742_ _2742_/A _2742_/B _2742_/C _2742_/D _3053_/D vdd gnd OAI22X1
X_2811_ _3068_/Q _2814_/A vdd gnd INVX1
X_1555_ _1555_/A _1555_/B rst _1562_/D vdd gnd AOI21X1
X_1624_ _1696_/Q _1630_/B _1664_/A vdd gnd NAND2X1
X_2673_ _3030_/Q _2702_/B _2676_/C vdd gnd NOR2X1
X_1486_ _1737_/B _1559_/Q _1487_/C vdd gnd NAND2X1
X_2107_ _2107_/A _2107_/B _2112_/A vdd gnd NAND2X1
X_3087_ _3087_/D _3087_/CLK _3087_/Q vdd gnd DFFPOSX1
X_2038_ _2038_/A _2039_/C vdd gnd INVX1
X_3010_ _3099_/Q _3013_/A vdd gnd INVX1
X_2656_ _2665_/A _2656_/B _2656_/C _2656_/D _3036_/D vdd gnd AOI22X1
X_2725_ _3004_/A _2741_/B _2742_/B _2726_/C vdd gnd OAI21X1
X_1469_ _1469_/A _1470_/B vdd gnd INVX1
X_1538_ _1545_/A _1545_/B _1552_/B _1539_/A vdd gnd OAI21X1
X_1607_ _1607_/A _2462_/Q _1658_/B vdd gnd NAND2X1
X_2587_ _3078_/Q _3022_/Q _2633_/S _2588_/A vdd gnd MUX2X1
X_2510_ _2512_/B _2510_/B _2510_/C _2523_/D vdd gnd OAI21X1
X_2372_ _2375_/C _2372_/B _2373_/B vdd gnd NAND2X1
X_2441_ _2441_/D _3095_/CLK _2441_/Q vdd gnd DFFPOSX1
X_2639_ _3051_/Q _3043_/Q _2643_/S _2640_/A vdd gnd MUX2X1
X_2708_ _2819_/B _2708_/B _2712_/B _2860_/A _2742_/B vdd gnd OAI22X1
X_1872_ vdd _1872_/Y vdd gnd INVX8
X_1941_ _2071_/A _2130_/A _1941_/C _1943_/B vdd gnd OAI21X1
X_2990_ _3030_/Q _3019_/B _2993_/C vdd gnd NOR2X1
X_2286_ _2286_/A _2286_/B _2288_/B vdd gnd NAND2X1
X_2355_ _2355_/A _2360_/B vdd gnd INVX1
X_2424_ _2424_/A _2424_/B _2424_/C _2425_/B vdd gnd OAI21X1
X_2140_ _2140_/A _2140_/B _2140_/C _2145_/A vdd gnd NAND3X1
X_2071_ _2071_/A _2206_/B _2146_/C vdd gnd NOR2X1
X_1855_ _1916_/A _1979_/C vdd gnd INVX1
X_1924_ _1928_/A _1989_/B _1989_/A _1928_/B vdd gnd NAND3X1
X_2973_ _2985_/A _2973_/B _2973_/C _2985_/D _2974_/C vdd gnd AOI22X1
X_1786_ _2427_/Q _2434_/Q _1788_/A vdd gnd NAND2X1
X_2269_ _2271_/A _2270_/A vdd gnd INVX1
X_2338_ _2338_/A _2360_/A vdd gnd INVX1
X_2407_ _2412_/A _2413_/A vdd gnd INVX1
X_1571_ _1676_/Q _1669_/B vdd gnd INVX1
X_1640_ _1644_/A _1640_/B _1669_/C _1642_/B vdd gnd OAI21X1
X_2123_ _2123_/A _2123_/B _2123_/C _2124_/B vdd gnd AOI21X1
X_2054_ _2117_/B _2054_/B _2057_/B vdd gnd NAND2X1
X_1838_ _2429_/Q _2436_/Q _1886_/B vdd gnd AND2X2
X_1907_ _1907_/A _1907_/B _1931_/C _1909_/C vdd gnd OAI21X1
X_2956_ _3067_/Q _3099_/Q _2956_/S _2958_/B vdd gnd MUX2X1
X_2887_ _3037_/Q _2887_/B _2889_/C vdd gnd NOR2X1
X_1769_ vdd _2080_/A _1769_/C _2436_/D vdd gnd OAI21X1
X_2672_ _2985_/A _2989_/B _2702_/B vdd gnd NAND2X1
X_2741_ _3020_/A _2741_/B _2742_/B _2742_/C vdd gnd OAI21X1
X_2810_ _2810_/A _2818_/B _2810_/C _2810_/D _3067_/D vdd gnd OAI22X1
X_1485_ _2519_/Q _1557_/Q _1487_/B vdd gnd NAND2X1
X_1554_ _1737_/B _1554_/B _1555_/A vdd gnd NAND2X1
X_1623_ _1663_/B _1663_/A _2395_/A vdd gnd NAND2X1
.ends

