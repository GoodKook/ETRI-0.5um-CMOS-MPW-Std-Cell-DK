/* Verilog module written by vlog2Verilog (qflow) */
/* With bit-blasted vectors */
/* With power connections converted to binary 1, 0 */

module booth_multiplier(
    input clk,
    input [7:0] multIn,
    output [15:0] product,
    input select
);

wire \step3.myadd.fa7.i1  ;
wire \step6.myadd.fa3.cout  ;
wire _588_ ;
wire _168_ ;
wire _800_ ;
wire _60_ ;
wire _397_ ;
wire \step3.myadd.fa2.i1  ;
wire [15:0] _product ;
wire \step3.myadd.fa3.sum  ;
wire \step6.myadd.fa3.i0  ;
wire \step8.myadd.fa1.sum  ;
wire \step1.myadd.x2.i0_bF$buf1  ;
wire \step5.myadd.fa7.i1  ;
wire _703_ ;
wire \step5.myadd.fa2.i1  ;
wire _19_ ;
wire _512_ ;
wire \step8.myadd.fa3.i0  ;
wire \step3.myadd.cin_bF$buf4  ;
wire \step5.myadd.fa5.cout  ;
wire \step3.myadd.fa5.sum  ;
wire _741_ ;
wire _321_ ;
wire \step8.myadd.fa3.sum  ;
wire \step7.myadd.fa7.i1  ;
wire _57_ ;
wire _550_ ;
wire _130_ ;
wire _606_ ;
wire \step5.myadd.cin_bF$buf0  ;
wire \step7.myadd.fa2.i1  ;
wire _835_ ;
wire _415_ ;
wire _95_ ;
wire _644_ ;
wire _224_ ;
wire \step3.myadd.fa7.cout  ;
wire \step3.myadd.fa7.sum  ;
wire _873_ ;
wire _453_ ;
wire \step8.myadd.fa5.sum  ;
wire _509_ ;
wire _682_ ;
wire _262_ ;
wire _738_ ;
wire _318_ ;
wire _491_ ;
wire _547_ ;
wire _127_ ;
wire _776_ ;
wire _356_ ;
wire _585_ ;
wire _165_ ;
wire _394_ ;
wire \step1.myadd.x5.i0  ;
wire \step1.myadd.x1.i0_bF$buf3  ;
wire _679_ ;
wire _259_ ;
wire _488_ ;
wire \step1.myadd.x0.i0  ;
wire _700_ ;
wire _297_ ;
wire _16_ ;
wire \step3.myadd.cin_bF$buf1  ;
wire _54_ ;
wire _603_ ;
wire \step4.myadd.fa6.i1  ;
wire _832_ ;
wire _412_ ;
wire _92_ ;
wire _641_ ;
wire _221_ ;
wire \step4.myadd.fa1.i1  ;
wire _870_ ;
wire _450_ ;
wire _506_ ;
wire \step6.myadd.fa6.i1  ;
wire _735_ ;
wire _315_ ;
wire [7:0] \Q[3]  ;
wire _544_ ;
wire _124_ ;
wire \step1.myadd.x7.i0_bF$buf2  ;
wire \step6.myadd.fa1.i1  ;
wire \step6.myadd.fa1.cout  ;
wire _773_ ;
wire _353_ ;
wire _829_ ;
wire _409_ ;
wire _89_ ;
wire _582_ ;
wire _162_ ;
wire _638_ ;
wire _218_ ;
wire \step8.myadd.fa6.i1  ;
wire _391_ ;
wire _867_ ;
wire _447_ ;
wire \step8.myadd.fa1.i1  ;
wire \step1.myadd.x1.i0_bF$buf0  ;
wire _676_ ;
wire _256_ ;
wire \step4.myadd.fa2.sum  ;
wire \step4.myadd.fa3.cout  ;
wire \step1.myadd.cin_bF$buf2  ;
wire _485_ ;
wire _294_ ;
wire _13_ ;
wire _579_ ;
wire _159_ ;
wire _51_ ;
wire _388_ ;
wire \step4.myadd.fa4.sum  ;
wire _600_ ;
wire _197_ ;
wire \step3.myadd.fa5.cout  ;
wire _7_ ;
wire _503_ ;
wire \step4.myadd.fa6.sum  ;
wire _732_ ;
wire _312_ ;
wire \step8.myadd.fa4.cout  ;
wire _48_ ;
wire \step1.myadd.fa7.cout  ;
wire _541_ ;
wire _121_ ;
wire _770_ ;
wire _350_ ;
wire \step2.myadd.fa4.i0  ;
wire _826_ ;
wire _406_ ;
wire _86_ ;
wire _635_ ;
wire _215_ ;
wire \step4.myadd.fa8.sum  ;
wire _864_ ;
wire _444_ ;
wire \step1.myadd.x0.i0_bF$buf2  ;
wire _673_ ;
wire _253_ ;
wire _729_ ;
wire _309_ ;
wire _482_ ;
wire select ;
wire _538_ ;
wire _118_ ;
wire _291_ ;
wire _10_ ;
wire _767_ ;
wire _347_ ;
wire _576_ ;
wire _156_ ;
wire _385_ ;
wire _194_ ;
wire _899_ ;
wire _479_ ;
wire _288_ ;
wire _4_ ;
wire _500_ ;
wire \step3.myadd.cin  ;
wire _45_ ;
wire \step1.myadd.x6.i0_bF$buf1  ;
wire _823_ ;
wire _403_ ;
wire _83_ ;
wire _632_ ;
wire _212_ ;
wire _861_ ;
wire _441_ ;
wire \step4.myadd.fa1.cout  ;
wire _670_ ;
wire _250_ ;
wire _726_ ;
wire _306_ ;
wire \step5.myadd.fa1.sum  ;
wire _535_ ;
wire _115_ ;
wire _764_ ;
wire _344_ ;
wire _573_ ;
wire _153_ ;
wire \step2.myadd.fa3.cout  ;
wire _629_ ;
wire _209_ ;
wire _382_ ;
wire \step6.myadd.cin_bF$buf2  ;
wire _858_ ;
wire _438_ ;
wire _191_ ;
wire \step3.myadd.fa3.i0  ;
wire \step5.myadd.fa3.sum  ;
wire _667_ ;
wire _247_ ;
wire \step2.myadd.fa7.i1  ;
wire _896_ ;
wire _476_ ;
wire clk_bF$buf0 ;
wire clk_bF$buf1 ;
wire clk_bF$buf2 ;
wire clk_bF$buf3 ;
wire clk_bF$buf4 ;
wire _285_ ;
wire _1_ ;
wire \step2.myadd.fa2.i1  ;
wire \step5.myadd.fa3.i0  ;
wire _42_ ;
wire \step5.myadd.fa5.sum  ;
wire _799_ ;
wire _379_ ;
wire \step1.myadd.x5.i0_bF$buf3  ;
wire _188_ ;
wire _820_ ;
wire _400_ ;
wire _80_ ;
wire \step7.myadd.fa3.i0  ;
wire \step6.myadd.fa4.cout  ;
wire \step5.myadd.fa7.sum  ;
wire _723_ ;
wire _303_ ;
wire _39_ ;
wire _532_ ;
wire _112_ ;
wire \step4.myadd.fa6.cout  ;
wire \step4.myadd.cin_bF$buf3  ;
wire _761_ ;
wire _341_ ;
wire clk ;
wire _817_ ;
wire _77_ ;
wire _570_ ;
wire _150_ ;
wire _626_ ;
wire _206_ ;
wire _855_ ;
wire _435_ ;
wire _664_ ;
wire _244_ ;
wire _893_ ;
wire _473_ ;
wire _529_ ;
wire _109_ ;
wire _282_ ;
wire _758_ ;
wire _338_ ;
wire _567_ ;
wire _147_ ;
wire _796_ ;
wire _376_ ;
wire \step1.myadd.x5.i0_bF$buf0  ;
wire \step8.myadd.fa7.cout  ;
wire _185_ ;
wire \step1.myadd.fa6.i1  ;
wire \step4.myadd.fa7.i0  ;
wire \step1.myadd.fa1.i1  ;
wire _699_ ;
wire _279_ ;
wire _911_ ;
wire \step4.myadd.fa2.i0  ;
wire \step2.myadd.cin_bF$buf4  ;
wire _720_ ;
wire _300_ ;
wire \step3.myadd.fa6.i1  ;
wire _36_ ;
wire \step6.myadd.fa7.i0  ;
wire \step4.myadd.cin_bF$buf0  ;
wire \step3.myadd.fa1.i1  ;
wire _814_ ;
wire _74_ ;
wire \step6.myadd.fa2.i0  ;
wire _623_ ;
wire _203_ ;
wire \step5.myadd.fa6.i1  ;
wire _852_ ;
wire _432_ ;
wire \step8.myadd.fa7.i0  ;
wire _908_ ;
wire _661_ ;
wire _241_ ;
wire \step5.myadd.fa1.i1  ;
wire _717_ ;
wire \step1.myadd.fa4.sum  ;
wire _890_ ;
wire \step8.myadd.fa2.i0  ;
wire _470_ ;
wire \step6.myadd.fa2.sum  ;
wire _526_ ;
wire _106_ ;
wire \step7.myadd.fa6.i1  ;
wire _755_ ;
wire _335_ ;
wire [7:0] \Q[5]  ;
wire _564_ ;
wire _144_ ;
wire \step7.myadd.fa1.i1  ;
wire _793_ ;
wire _373_ ;
wire \step1.myadd.x4.i0_bF$buf2  ;
wire _849_ ;
wire _429_ ;
wire \step1.myadd.fa6.sum  ;
wire _182_ ;
wire \step6.myadd.fa4.sum  ;
wire _658_ ;
wire _238_ ;
wire _887_ ;
wire _467_ ;
wire _696_ ;
wire _276_ ;
wire \step2.myadd.cin_bF$buf1  ;
wire \step1.myadd.fa8.sum  ;
wire \step6.myadd.fa6.sum  ;
wire \step4.myadd.fa4.cout  ;
wire _33_ ;
wire _599_ ;
wire _179_ ;
wire _811_ ;
wire _71_ ;
wire \step1.myadd.x4.i0  ;
wire _620_ ;
wire _200_ ;
wire \step2.myadd.fa6.cout  ;
wire \step6.myadd.fa8.sum  ;
wire _905_ ;
wire \step1.myadd.cin  ;
wire _714_ ;
wire _523_ ;
wire _103_ ;
wire _752_ ;
wire _332_ ;
wire _808_ ;
wire _68_ ;
wire _561_ ;
wire _141_ ;
wire [15:0] product ;
wire \step4.myadd.fa5.i1  ;
wire _617_ ;
wire _790_ ;
wire _370_ ;
wire _846_ ;
wire _426_ ;
wire _655_ ;
wire _235_ ;
wire _884_ ;
wire _464_ ;
wire \step6.myadd.fa5.i1  ;
wire _693_ ;
wire _273_ ;
wire \step6.myadd.fa7.cout  ;
wire _749_ ;
wire _329_ ;
wire _558_ ;
wire _138_ ;
wire _30_ ;
wire _787_ ;
wire _367_ ;
wire \step8.myadd.fa5.i1  ;
wire _596_ ;
wire _176_ ;
wire \step7.myadd.cin_bF$buf4  ;
wire _902_ ;
wire _499_ ;
wire _711_ ;
wire _27_ ;
wire _520_ ;
wire _100_ ;
wire \step7.myadd.fa1.sum  ;
wire _805_ ;
wire _65_ ;
wire _614_ ;
wire \step1.myadd.x3.i0_bF$buf1  ;
wire _843_ ;
wire _423_ ;
wire _652_ ;
wire _232_ ;
wire \step2.myadd.fa5.sum  ;
wire _708_ ;
wire \step7.myadd.fa3.sum  ;
wire _881_ ;
wire _461_ ;
wire \step3.myadd.fa2.cout  ;
wire _517_ ;
wire _690_ ;
wire _270_ ;
wire _746_ ;
wire _326_ ;
wire \step2.myadd.fa3.i0  ;
wire _555_ ;
wire _135_ ;
wire _784_ ;
wire _364_ ;
wire \step2.myadd.fa7.sum  ;
wire \step7.myadd.fa5.sum  ;
wire _593_ ;
wire _173_ ;
wire _649_ ;
wire _229_ ;
wire \step7.myadd.cin_bF$buf1  ;
wire _878_ ;
wire _458_ ;
wire \step2.myadd.fa4.cout  ;
wire _687_ ;
wire _267_ ;
wire _496_ ;
wire \step7.myadd.fa7.sum  ;
wire _24_ ;
wire \step7.myadd.fa3.cout  ;
wire _802_ ;
wire _62_ ;
wire _399_ ;
wire _611_ ;
wire \step1.myadd.x2.i0_bF$buf3  ;
wire _840_ ;
wire _420_ ;
wire _705_ ;
wire [7:0] \Q[0]  ;
wire _514_ ;
wire _743_ ;
wire _323_ ;
wire _59_ ;
wire _552_ ;
wire _132_ ;
wire _608_ ;
wire _781_ ;
wire _361_ ;
wire \step5.myadd.cin_bF$buf2  ;
wire _837_ ;
wire _417_ ;
wire _97_ ;
wire _590_ ;
wire _170_ ;
wire \step4.myadd.fa7.cout  ;
wire _646_ ;
wire _226_ ;
wire _875_ ;
wire _455_ ;
wire _684_ ;
wire _264_ ;
wire _493_ ;
wire _549_ ;
wire _129_ ;
wire _21_ ;
wire _778_ ;
wire _358_ ;
wire \step3.myadd.fa7.i0  ;
wire _587_ ;
wire _167_ ;
wire _396_ ;
wire \step3.myadd.fa2.i0  ;
wire \step2.myadd.fa6.i1  ;
wire \step1.myadd.x2.i0_bF$buf0  ;
wire \step5.myadd.fa7.i0  ;
wire \step2.myadd.fa1.i1  ;
wire _702_ ;
wire _299_ ;
wire \step5.myadd.fa2.i0  ;
wire _18_ ;
wire _511_ ;
wire \step8.myadd.fa2.sum  ;
wire \step3.myadd.cin_bF$buf3  ;
wire _740_ ;
wire _320_ ;
wire \step7.myadd.fa7.i0  ;
wire _56_ ;
wire _605_ ;
wire \step1.myadd.fa2.cout  ;
wire \step7.myadd.fa2.i0  ;
wire _834_ ;
wire _414_ ;
wire _94_ ;
wire \step3.myadd.fa6.sum  ;
wire _643_ ;
wire _223_ ;
wire \step8.myadd.fa4.sum  ;
wire _872_ ;
wire _452_ ;
wire _508_ ;
wire _681_ ;
wire _261_ ;
wire _737_ ;
wire _317_ ;
wire _490_ ;
wire _546_ ;
wire _126_ ;
wire \step3.myadd.fa8.sum  ;
wire _775_ ;
wire _355_ ;
wire \step8.myadd.fa6.sum  ;
wire _584_ ;
wire _164_ ;
wire _393_ ;
wire _869_ ;
wire _449_ ;
wire \step1.myadd.x1.i0_bF$buf2  ;
wire \step5.myadd.fa3.cout  ;
wire _678_ ;
wire _258_ ;
wire \step1.myadd.cin_bF$buf4  ;
wire _487_ ;
wire \step8.myadd.fa8.sum  ;
wire _296_ ;
wire _15_ ;
wire \step3.myadd.cin_bF$buf0  ;
wire _53_ ;
wire _602_ ;
wire \step1.myadd.fa5.i1  ;
wire _199_ ;
wire \step4.myadd.fa6.i0  ;
wire _831_ ;
wire _411_ ;
wire _91_ ;
wire _640_ ;
wire _220_ ;
wire \step4.myadd.fa1.i0  ;
wire _9_ ;
wire _505_ ;
wire \step3.myadd.fa5.i1  ;
wire \step6.myadd.fa6.i0  ;
wire _734_ ;
wire _314_ ;
wire \step2.myadd.fa7.cout  ;
wire _543_ ;
wire _123_ ;
wire \step1.myadd.x7.i0_bF$buf1  ;
wire \step6.myadd.fa1.i0  ;
wire _772_ ;
wire _352_ ;
wire _828_ ;
wire _408_ ;
wire _88_ ;
wire \step5.myadd.fa5.i1  ;
wire _581_ ;
wire _161_ ;
wire _637_ ;
wire _217_ ;
wire \step8.myadd.fa6.i0  ;
wire \step7.myadd.fa6.cout  ;
wire _390_ ;
wire _866_ ;
wire _446_ ;
wire \step8.myadd.fa1.i0  ;
wire _675_ ;
wire _255_ ;
wire \step1.myadd.cin_bF$buf1  ;
wire _484_ ;
wire \step7.myadd.fa5.i1  ;
wire _293_ ;
wire _12_ ;
wire _769_ ;
wire _349_ ;
wire _578_ ;
wire _158_ ;
wire _50_ ;
wire _387_ ;
wire _196_ ;
wire _6_ ;
wire \step4.myadd.fa5.sum  ;
wire _502_ ;
wire _731_ ;
wire _311_ ;
wire _47_ ;
wire _540_ ;
wire _120_ ;
wire \step1.myadd.x6.i0_bF$buf3  ;
wire \step1.myadd.x3.i0  ;
wire _825_ ;
wire _405_ ;
wire _85_ ;
wire \step4.myadd.fa7.sum  ;
wire _634_ ;
wire _214_ ;
wire _863_ ;
wire _443_ ;
wire \step1.myadd.x0.i0_bF$buf1  ;
wire _672_ ;
wire _252_ ;
wire _728_ ;
wire _308_ ;
wire _481_ ;
wire _537_ ;
wire _117_ ;
wire _290_ ;
wire _766_ ;
wire _346_ ;
wire \step4.myadd.fa4.i1  ;
wire \step3.myadd.fa3.cout  ;
wire _575_ ;
wire _155_ ;
wire _384_ ;
wire \step6.myadd.cin_bF$buf4  ;
wire _193_ ;
wire _669_ ;
wire _249_ ;
wire \step8.myadd.fa2.cout  ;
wire \step6.myadd.fa4.i1  ;
wire _898_ ;
wire _478_ ;
wire \step1.myadd.fa5.cout  ;
wire _287_ ;
wire _3_ ;
wire \step8.myadd.fa4.i1  ;
wire _44_ ;
wire \step1.myadd.x6.i0_bF$buf0  ;
wire _822_ ;
wire _402_ ;
wire _82_ ;
wire _631_ ;
wire _211_ ;
wire _860_ ;
wire _440_ ;
wire _725_ ;
wire _305_ ;
wire [7:0] \Q[2]  ;
wire \step5.myadd.fa6.cout  ;
wire _534_ ;
wire _114_ ;
wire _763_ ;
wire _343_ ;
wire _819_ ;
wire _79_ ;
wire _572_ ;
wire _152_ ;
wire _628_ ;
wire _208_ ;
wire _381_ ;
wire \step6.myadd.cin_bF$buf1  ;
wire _857_ ;
wire _437_ ;
wire _190_ ;
wire _666_ ;
wire _246_ ;
wire \step2.myadd.fa7.i0  ;
wire _895_ ;
wire _475_ ;
wire qout_bF$buf0 ;
wire qout_bF$buf1 ;
wire qout_bF$buf2 ;
wire qout_bF$buf3 ;
wire qout_bF$buf4 ;
wire _284_ ;
wire _0_ ;
wire \step2.myadd.fa2.i0  ;
wire _569_ ;
wire _149_ ;
wire _41_ ;
wire _798_ ;
wire _378_ ;
wire \step1.myadd.x5.i0_bF$buf2  ;
wire _187_ ;
wire \step5.myadd.fa6.sum  ;
wire \step1.myadd.fa2.sum  ;
wire \step2.myadd.fa1.cout  ;
wire _722_ ;
wire _302_ ;
wire _38_ ;
wire _531_ ;
wire _111_ ;
wire \step4.myadd.cin_bF$buf2  ;
wire _760_ ;
wire _340_ ;
wire _816_ ;
wire _76_ ;
wire \step5.myadd.fa8.sum  ;
wire _625_ ;
wire _205_ ;
wire _854_ ;
wire _434_ ;
wire _663_ ;
wire _243_ ;
wire \step1.myadd.fa3.cout  ;
wire _719_ ;
wire _892_ ;
wire _472_ ;
wire _528_ ;
wire _108_ ;
wire _281_ ;
wire _757_ ;
wire _337_ ;
wire _566_ ;
wire _146_ ;
wire \step6.myadd.fa2.cout  ;
wire _795_ ;
wire _375_ ;
wire _184_ ;
wire _889_ ;
wire _469_ ;
wire _698_ ;
wire _278_ ;
wire _910_ ;
wire \step2.myadd.cin_bF$buf3  ;
wire \step3.myadd.fa6.i0  ;
wire _35_ ;
wire \step3.myadd.fa1.i0  ;
wire _813_ ;
wire _73_ ;
wire \step2.myadd.fa5.i1  ;
wire _622_ ;
wire _202_ ;
wire \step5.myadd.fa6.i0  ;
wire \step3.myadd.fa6.cout  ;
wire _851_ ;
wire _431_ ;
wire _907_ ;
wire _660_ ;
wire _240_ ;
wire \step5.myadd.fa1.i0  ;
wire _716_ ;
wire _525_ ;
wire _105_ ;
wire \step8.myadd.fa5.cout  ;
wire \step7.myadd.fa6.i0  ;
wire qout ;
wire _754_ ;
wire _334_ ;
wire _563_ ;
wire _143_ ;
wire \step7.myadd.fa1.i0  ;
wire _619_ ;
wire _792_ ;
wire _372_ ;
wire \step1.myadd.x4.i0_bF$buf1  ;
wire _848_ ;
wire _428_ ;
wire _181_ ;
wire _657_ ;
wire _237_ ;
wire _886_ ;
wire _466_ ;
wire _695_ ;
wire _275_ ;
wire \step7.myadd.fa7.cout  ;
wire \step2.myadd.cin_bF$buf0  ;
wire \step2.myadd.fa1.sum  ;
wire _32_ ;
wire _789_ ;
wire _369_ ;
wire _598_ ;
wire _178_ ;
wire _810_ ;
wire _70_ ;
wire \step6.myadd.fa7.sum  ;
wire \step2.myadd.fa3.sum  ;
wire _904_ ;
wire _713_ ;
wire _29_ ;
wire _522_ ;
wire _102_ ;
wire \step6.myadd.cin  ;
wire _751_ ;
wire _331_ ;
wire \step1.myadd.fa4.i1  ;
wire _807_ ;
wire _67_ ;
wire _560_ ;
wire _140_ ;
wire \step4.myadd.fa5.i0  ;
wire _616_ ;
wire \step1.myadd.x3.i0_bF$buf3  ;
wire _845_ ;
wire _425_ ;
wire _654_ ;
wire _234_ ;
wire \step3.myadd.fa4.i1  ;
wire _883_ ;
wire _463_ ;
wire \step4.myadd.fa2.cout  ;
wire \step6.myadd.fa5.i0  ;
wire _519_ ;
wire _692_ ;
wire _272_ ;
wire _748_ ;
wire _328_ ;
wire _557_ ;
wire _137_ ;
wire \step5.myadd.fa4.i1  ;
wire _786_ ;
wire _366_ ;
wire \step8.myadd.fa5.i0  ;
wire _595_ ;
wire _175_ ;
wire \step7.myadd.cin_bF$buf3  ;
wire \step7.myadd.fa4.i1  ;
wire _689_ ;
wire _269_ ;
wire _901_ ;
wire _498_ ;
wire _710_ ;
wire \step8.myadd.fa3.cout  ;
wire _26_ ;
wire \step1.myadd.fa6.cout  ;
wire _804_ ;
wire _64_ ;
wire _613_ ;
wire \step1.myadd.x3.i0_bF$buf0  ;
wire _842_ ;
wire _422_ ;
wire \step6.myadd.fa5.cout  ;
wire _651_ ;
wire _231_ ;
wire _707_ ;
wire _880_ ;
wire _460_ ;
wire _516_ ;
wire \step1.myadd.x7.i0  ;
wire _745_ ;
wire _325_ ;
wire [7:0] \Q[4]  ;
wire _554_ ;
wire _134_ ;
wire \step1.myadd.x2.i0  ;
wire _783_ ;
wire _363_ ;
wire \step5.myadd.cin_bF$buf4  ;
wire _839_ ;
wire _419_ ;
wire _99_ ;
wire _592_ ;
wire _172_ ;
wire _648_ ;
wire _228_ ;
wire \step7.myadd.cin_bF$buf0  ;
wire _877_ ;
wire _457_ ;
wire _686_ ;
wire _266_ ;
wire \step4.myadd.fa8.i1  ;
wire \step7.myadd.fa6.sum  ;
wire _495_ ;
wire \step3.myadd.fa2.sum  ;
wire \step4.myadd.fa3.i1  ;
wire _23_ ;
wire _589_ ;
wire _169_ ;
wire \step6.myadd.fa8.i1  ;
wire _801_ ;
wire _61_ ;
wire _398_ ;
wire _610_ ;
wire \step7.myadd.fa8.sum  ;
wire \step6.myadd.fa3.i1  ;
wire \step1.myadd.x2.i0_bF$buf2  ;
wire \step3.myadd.fa4.sum  ;
wire \step8.myadd.fa8.i1  ;
wire _704_ ;
wire _513_ ;
wire \step8.myadd.fa3.i1  ;
wire _742_ ;
wire _322_ ;
wire _58_ ;
wire _551_ ;
wire _131_ ;
wire _607_ ;
wire \step2.myadd.fa2.cout  ;
wire _780_ ;
wire _360_ ;
wire \step5.myadd.cin_bF$buf1  ;
wire _836_ ;
wire _416_ ;
wire _96_ ;
wire _645_ ;
wire _225_ ;
wire _874_ ;
wire _454_ ;
wire \step7.myadd.fa1.cout  ;
wire _683_ ;
wire _263_ ;
wire _739_ ;
wire _319_ ;
wire _492_ ;
wire _548_ ;
wire _128_ ;
wire _20_ ;
wire _777_ ;
wire _357_ ;
wire _586_ ;
wire _166_ ;
wire _395_ ;
wire \step2.myadd.fa6.i0  ;
wire _489_ ;
wire \step2.myadd.fa1.i0  ;
wire _701_ ;
wire _298_ ;
wire _17_ ;
wire _510_ ;
wire \step3.myadd.cin_bF$buf2  ;
wire \step4.myadd.fa5.cout  ;
wire _55_ ;
wire _604_ ;
wire _833_ ;
wire _413_ ;
wire _93_ ;
wire _642_ ;
wire _222_ ;
wire _871_ ;
wire _451_ ;
wire _507_ ;
wire _680_ ;
wire _260_ ;
wire \step4.myadd.cin  ;
wire _736_ ;
wire _316_ ;
wire select_bF$buf0 ;
wire select_bF$buf1 ;
wire select_bF$buf2 ;
wire select_bF$buf3 ;
wire select_bF$buf4 ;
wire _545_ ;
wire _125_ ;
wire \step1.myadd.x7.i0_bF$buf3  ;
wire _774_ ;
wire _354_ ;
wire \step4.myadd.fa1.sum  ;
wire _583_ ;
wire _163_ ;
wire \step8.myadd.fa6.cout  ;
wire _639_ ;
wire _219_ ;
wire _392_ ;
wire _868_ ;
wire _448_ ;
wire \step1.myadd.x1.i0_bF$buf1  ;
wire _677_ ;
wire _257_ ;
wire \step8.myadd.fa7.sum  ;
wire \step1.myadd.cin_bF$buf3  ;
wire _486_ ;
wire \step4.myadd.fa3.sum  ;
wire _295_ ;
wire _14_ ;
wire _52_ ;
wire _389_ ;
wire _601_ ;
wire _198_ ;
wire _830_ ;
wire _410_ ;
wire _90_ ;
wire _8_ ;
wire _504_ ;
wire \step3.myadd.fa5.i0  ;
wire _733_ ;
wire _313_ ;
wire _49_ ;
wire _542_ ;
wire _122_ ;
wire \step1.myadd.x7.i0_bF$buf0  ;
wire _771_ ;
wire _351_ ;
wire \step2.myadd.fa4.i1  ;
wire \step5.myadd.fa1.cout  ;
wire _827_ ;
wire _407_ ;
wire _87_ ;
wire \step5.myadd.fa5.i0  ;
wire _580_ ;
wire _160_ ;
wire _636_ ;
wire _216_ ;
wire _865_ ;
wire _445_ ;
wire \step1.myadd.x0.i0_bF$buf3  ;
wire _674_ ;
wire _254_ ;
wire \step1.myadd.cin_bF$buf0  ;
wire _483_ ;
wire \step7.myadd.fa5.i0  ;
wire _539_ ;
wire _119_ ;
wire _292_ ;
wire _11_ ;
wire _768_ ;
wire _348_ ;
wire _577_ ;
wire _157_ ;
wire _386_ ;
wire _195_ ;
wire \step2.myadd.fa5.cout  ;
wire _289_ ;
wire _5_ ;
wire _501_ ;
wire _730_ ;
wire _310_ ;
wire \step7.myadd.fa4.cout  ;
wire _46_ ;
wire \step1.myadd.x6.i0_bF$buf2  ;
wire _824_ ;
wire _404_ ;
wire _84_ ;
wire _633_ ;
wire _213_ ;
wire _862_ ;
wire _442_ ;
wire \step1.myadd.x0.i0_bF$buf0  ;
wire _671_ ;
wire _251_ ;
wire \step1.myadd.fa8.i1  ;
wire _727_ ;
wire _307_ ;
wire _480_ ;
wire \step6.myadd.fa6.cout  ;
wire _536_ ;
wire _116_ ;
wire \step1.myadd.fa3.i1  ;
wire \step5.myadd.fa2.sum  ;
wire _765_ ;
wire _345_ ;
wire \step4.myadd.fa4.i0  ;
wire [7:0] \Q[6]  ;
wire _574_ ;
wire _154_ ;
wire \step3.myadd.fa8.i1  ;
wire _383_ ;
wire \step6.myadd.cin_bF$buf3  ;
wire [7:0] multIn ;
wire _859_ ;
wire _439_ ;
wire _192_ ;
wire \step3.myadd.fa3.i1  ;
wire _668_ ;
wire _248_ ;
wire \step6.myadd.fa4.i0  ;
wire \step5.myadd.fa4.sum  ;
wire _897_ ;
wire _477_ ;
wire \step5.myadd.fa8.i1  ;
wire _286_ ;
wire _2_ ;
wire \step5.myadd.fa3.i1  ;
wire \step8.myadd.fa4.i0  ;
wire _43_ ;
wire \step7.myadd.fa8.i1  ;
wire _189_ ;
wire _821_ ;
wire _401_ ;
wire _81_ ;
wire \step7.myadd.fa3.i1  ;
wire _630_ ;
wire _210_ ;
wire \step3.myadd.fa1.cout  ;
wire _724_ ;
wire _304_ ;
wire _533_ ;
wire _113_ ;
wire \step4.myadd.cin_bF$buf4  ;
wire _762_ ;
wire _342_ ;
wire _818_ ;
wire _78_ ;
wire _571_ ;
wire _151_ ;
wire _627_ ;
wire _207_ ;
wire _380_ ;
wire \step6.myadd.cin_bF$buf0  ;
wire _856_ ;
wire _436_ ;
wire _665_ ;
wire _245_ ;
wire \step2.myadd.cin  ;
wire \step1.myadd.x6.i0  ;
wire _894_ ;
wire _474_ ;
wire _283_ ;
wire \step1.myadd.x1.i0  ;
wire _759_ ;
wire _339_ ;
wire \step7.myadd.fa2.cout  ;
wire _568_ ;
wire _148_ ;
wire _40_ ;
wire _797_ ;
wire _377_ ;
wire \step1.myadd.x5.i0_bF$buf1  ;
wire _186_ ;
wire \step4.myadd.fa7.i1  ;
wire \step5.myadd.fa4.cout  ;
wire \step1.myadd.fa1.sum  ;
wire [15:0] _912_ ;
wire \step4.myadd.fa2.i1  ;
wire _721_ ;
wire _301_ ;
wire _37_ ;
wire _530_ ;
wire _110_ ;
wire \step6.myadd.fa7.i1  ;
wire \step4.myadd.cin_bF$buf1  ;
wire _815_ ;
wire \step1.myadd.fa3.sum  ;
wire _75_ ;
wire \step6.myadd.fa2.i1  ;
wire \step6.myadd.fa1.sum  ;
wire _624_ ;
wire _204_ ;
wire _853_ ;
wire _433_ ;
wire \step8.myadd.fa7.i1  ;
wire _909_ ;
wire _662_ ;
wire _242_ ;
wire _718_ ;
wire _891_ ;
wire \step8.myadd.fa2.i1  ;
wire _471_ ;
wire _527_ ;
wire _107_ ;
wire \step1.myadd.fa5.sum  ;
wire _280_ ;
wire \step6.myadd.fa3.sum  ;
wire _756_ ;
wire _336_ ;
wire _565_ ;
wire _145_ ;
wire _794_ ;
wire _374_ ;
wire \step7.myadd.cin  ;
wire \step1.myadd.x4.i0_bF$buf3  ;
wire _183_ ;
wire _659_ ;
wire _239_ ;
wire \step1.myadd.fa7.sum  ;
wire \step6.myadd.fa5.sum  ;
wire _888_ ;
wire _468_ ;
wire _697_ ;
wire _277_ ;
wire \step2.myadd.cin_bF$buf2  ;
wire _34_ ;
wire _812_ ;
wire _72_ ;
wire \step1.myadd.fa1.cout  ;
wire \step2.myadd.fa5.i0  ;
wire _621_ ;
wire _201_ ;
wire _850_ ;
wire _430_ ;
wire _906_ ;
wire _715_ ;
wire [7:0] \Q[1]  ;
wire _524_ ;
wire _104_ ;
wire _753_ ;
wire _333_ ;
wire _809_ ;
wire _69_ ;
wire _562_ ;
wire _142_ ;
wire _618_ ;
wire _791_ ;
wire _371_ ;
wire \step1.myadd.x4.i0_bF$buf0  ;
wire _847_ ;
wire _427_ ;
wire _180_ ;
wire _656_ ;
wire _236_ ;
wire \step5.myadd.fa2.cout  ;
wire _885_ ;
wire _465_ ;
wire _694_ ;
wire _274_ ;
wire _559_ ;
wire _139_ ;
wire _31_ ;
wire _788_ ;
wire _368_ ;
wire \step3.myadd.fa4.cout  ;
wire _597_ ;
wire _177_ ;
wire \step2.myadd.fa2.sum  ;
wire _903_ ;
wire _712_ ;
wire _28_ ;
wire _521_ ;
wire _101_ ;
wire _750_ ;
wire _330_ ;
wire \step2.myadd.fa4.sum  ;
wire _806_ ;
wire \step7.myadd.fa2.sum  ;
wire _66_ ;
wire _615_ ;
wire \step7.myadd.fa5.cout  ;
wire \step1.myadd.x3.i0_bF$buf2  ;
wire _844_ ;
wire _424_ ;
wire _653_ ;
wire _233_ ;
wire \step3.myadd.fa4.i0  ;
wire _709_ ;
wire _882_ ;
wire _462_ ;
wire \step2.myadd.fa6.sum  ;
wire \step7.myadd.fa4.sum  ;
wire _518_ ;
wire \step2.myadd.fa8.i1  ;
wire _691_ ;
wire _271_ ;
wire _747_ ;
wire _327_ ;
wire \step5.myadd.fa7.cout  ;
wire \step2.myadd.fa3.i1  ;
wire _556_ ;
wire _136_ ;
wire \step5.myadd.fa4.i0  ;
wire _785_ ;
wire _365_ ;
wire _594_ ;
wire _174_ ;
wire \step2.myadd.fa8.sum  ;
wire \step7.myadd.cin_bF$buf2  ;
wire _879_ ;
wire _459_ ;
wire \step7.myadd.fa4.i0  ;
wire _688_ ;
wire _268_ ;
wire _900_ ;
wire _497_ ;
wire _25_ ;
wire _803_ ;
wire _63_ ;
wire _612_ ;
wire _841_ ;
wire _421_ ;
wire _650_ ;
wire _230_ ;
wire _706_ ;
wire _515_ ;
wire _744_ ;
wire _324_ ;
wire _553_ ;
wire _133_ ;
wire _609_ ;
wire _782_ ;
wire _362_ ;
wire \step5.myadd.cin_bF$buf3  ;
wire _838_ ;
wire _418_ ;
wire _98_ ;
wire _591_ ;
wire _171_ ;
wire _647_ ;
wire _227_ ;
wire _876_ ;
wire _456_ ;
wire \step8.myadd.fa1.cout  ;
wire \step1.myadd.fa7.i1  ;
wire \step1.myadd.fa4.cout  ;
wire _685_ ;
wire _265_ ;
wire \step3.myadd.fa1.sum  ;
wire \step1.myadd.fa2.i1  ;
wire _494_ ;
wire \step4.myadd.fa3.i0  ;
wire _22_ ;
wire _779_ ;
wire _359_ ;
wire \step5.myadd.cin  ;

BUFX2 BUFX2_insert81 (
    .A(\step5.myadd.cin ),
    .Y(\step5.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert80 (
    .A(\step5.myadd.cin ),
    .Y(\step5.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert79 (
    .A(\step5.myadd.cin ),
    .Y(\step5.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert78 (
    .A(\step5.myadd.cin ),
    .Y(\step5.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert77 (
    .A(\step5.myadd.cin ),
    .Y(\step5.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert76 (
    .A(\step7.myadd.cin ),
    .Y(\step7.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert75 (
    .A(\step7.myadd.cin ),
    .Y(\step7.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert74 (
    .A(\step7.myadd.cin ),
    .Y(\step7.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert73 (
    .A(\step7.myadd.cin ),
    .Y(\step7.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert72 (
    .A(\step7.myadd.cin ),
    .Y(\step7.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert71 (
    .A(\step1.myadd.x1.i0 ),
    .Y(\step1.myadd.x1.i0_bF$buf0 )
);

BUFX2 BUFX2_insert70 (
    .A(\step1.myadd.x1.i0 ),
    .Y(\step1.myadd.x1.i0_bF$buf1 )
);

BUFX2 BUFX2_insert69 (
    .A(\step1.myadd.x1.i0 ),
    .Y(\step1.myadd.x1.i0_bF$buf2 )
);

BUFX2 BUFX2_insert68 (
    .A(\step1.myadd.x1.i0 ),
    .Y(\step1.myadd.x1.i0_bF$buf3 )
);

BUFX2 BUFX2_insert67 (
    .A(\step1.myadd.x6.i0 ),
    .Y(\step1.myadd.x6.i0_bF$buf0 )
);

BUFX2 BUFX2_insert66 (
    .A(\step1.myadd.x6.i0 ),
    .Y(\step1.myadd.x6.i0_bF$buf1 )
);

BUFX2 BUFX2_insert65 (
    .A(\step1.myadd.x6.i0 ),
    .Y(\step1.myadd.x6.i0_bF$buf2 )
);

BUFX2 BUFX2_insert64 (
    .A(\step1.myadd.x6.i0 ),
    .Y(\step1.myadd.x6.i0_bF$buf3 )
);

BUFX2 BUFX2_insert63 (
    .A(\step2.myadd.cin ),
    .Y(\step2.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert62 (
    .A(\step2.myadd.cin ),
    .Y(\step2.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert61 (
    .A(\step2.myadd.cin ),
    .Y(\step2.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert60 (
    .A(\step2.myadd.cin ),
    .Y(\step2.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert59 (
    .A(\step2.myadd.cin ),
    .Y(\step2.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert58 (
    .A(\step4.myadd.cin ),
    .Y(\step4.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert57 (
    .A(\step4.myadd.cin ),
    .Y(\step4.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert56 (
    .A(\step4.myadd.cin ),
    .Y(\step4.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert55 (
    .A(\step4.myadd.cin ),
    .Y(\step4.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert54 (
    .A(\step4.myadd.cin ),
    .Y(\step4.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert53 (
    .A(\step1.myadd.x2.i0 ),
    .Y(\step1.myadd.x2.i0_bF$buf0 )
);

BUFX2 BUFX2_insert52 (
    .A(\step1.myadd.x2.i0 ),
    .Y(\step1.myadd.x2.i0_bF$buf1 )
);

BUFX2 BUFX2_insert51 (
    .A(\step1.myadd.x2.i0 ),
    .Y(\step1.myadd.x2.i0_bF$buf2 )
);

BUFX2 BUFX2_insert50 (
    .A(\step1.myadd.x2.i0 ),
    .Y(\step1.myadd.x2.i0_bF$buf3 )
);

BUFX2 BUFX2_insert49 (
    .A(\step1.myadd.x7.i0 ),
    .Y(\step1.myadd.x7.i0_bF$buf0 )
);

BUFX2 BUFX2_insert48 (
    .A(\step1.myadd.x7.i0 ),
    .Y(\step1.myadd.x7.i0_bF$buf1 )
);

BUFX2 BUFX2_insert47 (
    .A(\step1.myadd.x7.i0 ),
    .Y(\step1.myadd.x7.i0_bF$buf2 )
);

BUFX2 BUFX2_insert46 (
    .A(\step1.myadd.x7.i0 ),
    .Y(\step1.myadd.x7.i0_bF$buf3 )
);

BUFX2 BUFX2_insert45 (
    .A(\step6.myadd.cin ),
    .Y(\step6.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert44 (
    .A(\step6.myadd.cin ),
    .Y(\step6.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert43 (
    .A(\step6.myadd.cin ),
    .Y(\step6.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert42 (
    .A(\step6.myadd.cin ),
    .Y(\step6.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert41 (
    .A(\step6.myadd.cin ),
    .Y(\step6.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert40 (
    .A(qout),
    .Y(qout_bF$buf0)
);

BUFX2 BUFX2_insert39 (
    .A(qout),
    .Y(qout_bF$buf1)
);

BUFX2 BUFX2_insert38 (
    .A(qout),
    .Y(qout_bF$buf2)
);

BUFX2 BUFX2_insert37 (
    .A(qout),
    .Y(qout_bF$buf3)
);

BUFX2 BUFX2_insert36 (
    .A(qout),
    .Y(qout_bF$buf4)
);

BUFX2 BUFX2_insert35 (
    .A(\step1.myadd.x3.i0 ),
    .Y(\step1.myadd.x3.i0_bF$buf0 )
);

BUFX2 BUFX2_insert34 (
    .A(\step1.myadd.x3.i0 ),
    .Y(\step1.myadd.x3.i0_bF$buf1 )
);

BUFX2 BUFX2_insert33 (
    .A(\step1.myadd.x3.i0 ),
    .Y(\step1.myadd.x3.i0_bF$buf2 )
);

BUFX2 BUFX2_insert32 (
    .A(\step1.myadd.x3.i0 ),
    .Y(\step1.myadd.x3.i0_bF$buf3 )
);

BUFX2 BUFX2_insert31 (
    .A(\step1.myadd.cin ),
    .Y(\step1.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert30 (
    .A(\step1.myadd.cin ),
    .Y(\step1.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert29 (
    .A(\step1.myadd.cin ),
    .Y(\step1.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert28 (
    .A(\step1.myadd.cin ),
    .Y(\step1.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert27 (
    .A(\step1.myadd.cin ),
    .Y(\step1.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert26 (
    .A(\step1.myadd.x4.i0 ),
    .Y(\step1.myadd.x4.i0_bF$buf0 )
);

BUFX2 BUFX2_insert25 (
    .A(\step1.myadd.x4.i0 ),
    .Y(\step1.myadd.x4.i0_bF$buf1 )
);

BUFX2 BUFX2_insert24 (
    .A(\step1.myadd.x4.i0 ),
    .Y(\step1.myadd.x4.i0_bF$buf2 )
);

BUFX2 BUFX2_insert23 (
    .A(\step1.myadd.x4.i0 ),
    .Y(\step1.myadd.x4.i0_bF$buf3 )
);

CLKBUF1 CLKBUF1_insert22 (
    .A(clk),
    .Y(clk_bF$buf0)
);

CLKBUF1 CLKBUF1_insert21 (
    .A(clk),
    .Y(clk_bF$buf1)
);

CLKBUF1 CLKBUF1_insert20 (
    .A(clk),
    .Y(clk_bF$buf2)
);

CLKBUF1 CLKBUF1_insert19 (
    .A(clk),
    .Y(clk_bF$buf3)
);

CLKBUF1 CLKBUF1_insert18 (
    .A(clk),
    .Y(clk_bF$buf4)
);

BUFX2 BUFX2_insert17 (
    .A(\step3.myadd.cin ),
    .Y(\step3.myadd.cin_bF$buf0 )
);

BUFX2 BUFX2_insert16 (
    .A(\step3.myadd.cin ),
    .Y(\step3.myadd.cin_bF$buf1 )
);

BUFX2 BUFX2_insert15 (
    .A(\step3.myadd.cin ),
    .Y(\step3.myadd.cin_bF$buf2 )
);

BUFX2 BUFX2_insert14 (
    .A(\step3.myadd.cin ),
    .Y(\step3.myadd.cin_bF$buf3 )
);

BUFX2 BUFX2_insert13 (
    .A(\step3.myadd.cin ),
    .Y(\step3.myadd.cin_bF$buf4 )
);

BUFX2 BUFX2_insert12 (
    .A(select),
    .Y(select_bF$buf0)
);

BUFX2 BUFX2_insert11 (
    .A(select),
    .Y(select_bF$buf1)
);

BUFX2 BUFX2_insert10 (
    .A(select),
    .Y(select_bF$buf2)
);

BUFX2 BUFX2_insert9 (
    .A(select),
    .Y(select_bF$buf3)
);

BUFX2 BUFX2_insert8 (
    .A(select),
    .Y(select_bF$buf4)
);

BUFX2 BUFX2_insert7 (
    .A(\step1.myadd.x0.i0 ),
    .Y(\step1.myadd.x0.i0_bF$buf0 )
);

BUFX2 BUFX2_insert6 (
    .A(\step1.myadd.x0.i0 ),
    .Y(\step1.myadd.x0.i0_bF$buf1 )
);

BUFX2 BUFX2_insert5 (
    .A(\step1.myadd.x0.i0 ),
    .Y(\step1.myadd.x0.i0_bF$buf2 )
);

BUFX2 BUFX2_insert4 (
    .A(\step1.myadd.x0.i0 ),
    .Y(\step1.myadd.x0.i0_bF$buf3 )
);

BUFX2 BUFX2_insert3 (
    .A(\step1.myadd.x5.i0 ),
    .Y(\step1.myadd.x5.i0_bF$buf0 )
);

BUFX2 BUFX2_insert2 (
    .A(\step1.myadd.x5.i0 ),
    .Y(\step1.myadd.x5.i0_bF$buf1 )
);

BUFX2 BUFX2_insert1 (
    .A(\step1.myadd.x5.i0 ),
    .Y(\step1.myadd.x5.i0_bF$buf2 )
);

BUFX2 BUFX2_insert0 (
    .A(\step1.myadd.x5.i0 ),
    .Y(\step1.myadd.x5.i0_bF$buf3 )
);

NAND3X1 _1000_ (
    .A(\step1.myadd.fa3.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_54_)
);

OAI21X1 _1001_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_55_)
);

NAND2X1 _1002_ (
    .A(_55_),
    .B(_54_),
    .Y(\step2.myadd.fa2.i0 )
);

NAND3X1 _1003_ (
    .A(\step1.myadd.fa4.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_56_)
);

OAI21X1 _1004_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_57_)
);

NAND2X1 _1005_ (
    .A(_57_),
    .B(_56_),
    .Y(\step2.myadd.fa3.i0 )
);

NAND3X1 _1006_ (
    .A(\step1.myadd.fa5.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_58_)
);

OAI21X1 _1007_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_59_)
);

NAND2X1 _1008_ (
    .A(_59_),
    .B(_58_),
    .Y(\step2.myadd.fa4.i0 )
);

NAND3X1 _1009_ (
    .A(\step1.myadd.fa6.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_60_)
);

OAI21X1 _1010_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_61_)
);

NAND2X1 _1011_ (
    .A(_61_),
    .B(_60_),
    .Y(\step2.myadd.fa5.i0 )
);

NAND3X1 _1012_ (
    .A(\step1.myadd.fa7.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_62_)
);

OAI21X1 _1013_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_63_)
);

NAND2X1 _1014_ (
    .A(_63_),
    .B(_62_),
    .Y(\step2.myadd.fa6.i0 )
);

NAND3X1 _1015_ (
    .A(\step1.myadd.fa8.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_64_)
);

OAI21X1 _1016_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_65_)
);

NAND2X1 _1017_ (
    .A(_65_),
    .B(_64_),
    .Y(\step2.myadd.fa7.i0 )
);

NAND3X1 _1018_ (
    .A(\step1.myadd.fa1.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_66_)
);

OAI21X1 _1019_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_67_)
);

NAND2X1 _1020_ (
    .A(_67_),
    .B(_66_),
    .Y(\Q[0] [7])
);

AND2X2 _1021_ (
    .A(\step1.myadd.fa1.i1 ),
    .B(\step1.myadd.cin_bF$buf4 ),
    .Y(_71_)
);

NOR2X1 _1022_ (
    .A(\step1.myadd.fa1.i1 ),
    .B(\step1.myadd.cin_bF$buf3 ),
    .Y(_72_)
);

OAI21X1 _1023_ (
    .A(_72_),
    .B(_71_),
    .C(gnd),
    .Y(_73_)
);

INVX1 _1024_ (
    .A(gnd),
    .Y(_74_)
);

NAND2X1 _1025_ (
    .A(\step1.myadd.fa1.i1 ),
    .B(\step1.myadd.cin_bF$buf2 ),
    .Y(_68_)
);

OR2X2 _1026_ (
    .A(\step1.myadd.fa1.i1 ),
    .B(\step1.myadd.cin_bF$buf1 ),
    .Y(_69_)
);

NAND3X1 _1027_ (
    .A(_74_),
    .B(_68_),
    .C(_69_),
    .Y(_70_)
);

NAND2X1 _1028_ (
    .A(_73_),
    .B(_70_),
    .Y(\step1.myadd.fa1.sum )
);

AOI21X1 _1029_ (
    .A(_74_),
    .B(_68_),
    .C(_72_),
    .Y(\step1.myadd.fa1.cout )
);

AND2X2 _1030_ (
    .A(\step1.myadd.fa2.i1 ),
    .B(\step1.myadd.fa1.cout ),
    .Y(_78_)
);

NOR2X1 _1031_ (
    .A(\step1.myadd.fa2.i1 ),
    .B(\step1.myadd.fa1.cout ),
    .Y(_79_)
);

OAI21X1 _1032_ (
    .A(_79_),
    .B(_78_),
    .C(gnd),
    .Y(_80_)
);

INVX1 _1033_ (
    .A(gnd),
    .Y(_81_)
);

NAND2X1 _1034_ (
    .A(\step1.myadd.fa2.i1 ),
    .B(\step1.myadd.fa1.cout ),
    .Y(_75_)
);

OR2X2 _1035_ (
    .A(\step1.myadd.fa2.i1 ),
    .B(\step1.myadd.fa1.cout ),
    .Y(_76_)
);

NAND3X1 _1036_ (
    .A(_81_),
    .B(_75_),
    .C(_76_),
    .Y(_77_)
);

NAND2X1 _1037_ (
    .A(_80_),
    .B(_77_),
    .Y(\step1.myadd.fa2.sum )
);

AOI21X1 _1038_ (
    .A(_81_),
    .B(_75_),
    .C(_79_),
    .Y(\step1.myadd.fa2.cout )
);

AND2X2 _1039_ (
    .A(\step1.myadd.fa3.i1 ),
    .B(\step1.myadd.fa2.cout ),
    .Y(_85_)
);

NOR2X1 _1040_ (
    .A(\step1.myadd.fa3.i1 ),
    .B(\step1.myadd.fa2.cout ),
    .Y(_86_)
);

OAI21X1 _1041_ (
    .A(_86_),
    .B(_85_),
    .C(gnd),
    .Y(_87_)
);

INVX1 _1042_ (
    .A(gnd),
    .Y(_88_)
);

NAND2X1 _1043_ (
    .A(\step1.myadd.fa3.i1 ),
    .B(\step1.myadd.fa2.cout ),
    .Y(_82_)
);

OR2X2 _1044_ (
    .A(\step1.myadd.fa3.i1 ),
    .B(\step1.myadd.fa2.cout ),
    .Y(_83_)
);

NAND3X1 _1045_ (
    .A(_88_),
    .B(_82_),
    .C(_83_),
    .Y(_84_)
);

NAND2X1 _1046_ (
    .A(_87_),
    .B(_84_),
    .Y(\step1.myadd.fa3.sum )
);

AOI21X1 _1047_ (
    .A(_88_),
    .B(_82_),
    .C(_86_),
    .Y(\step1.myadd.fa3.cout )
);

AND2X2 _1048_ (
    .A(\step1.myadd.fa4.i1 ),
    .B(\step1.myadd.fa3.cout ),
    .Y(_92_)
);

NOR2X1 _1049_ (
    .A(\step1.myadd.fa4.i1 ),
    .B(\step1.myadd.fa3.cout ),
    .Y(_93_)
);

OAI21X1 _1050_ (
    .A(_93_),
    .B(_92_),
    .C(gnd),
    .Y(_94_)
);

INVX1 _1051_ (
    .A(gnd),
    .Y(_95_)
);

NAND2X1 _1052_ (
    .A(\step1.myadd.fa4.i1 ),
    .B(\step1.myadd.fa3.cout ),
    .Y(_89_)
);

OR2X2 _1053_ (
    .A(\step1.myadd.fa4.i1 ),
    .B(\step1.myadd.fa3.cout ),
    .Y(_90_)
);

NAND3X1 _1054_ (
    .A(_95_),
    .B(_89_),
    .C(_90_),
    .Y(_91_)
);

NAND2X1 _1055_ (
    .A(_94_),
    .B(_91_),
    .Y(\step1.myadd.fa4.sum )
);

AOI21X1 _1056_ (
    .A(_95_),
    .B(_89_),
    .C(_93_),
    .Y(\step1.myadd.fa4.cout )
);

AND2X2 _1057_ (
    .A(\step1.myadd.fa5.i1 ),
    .B(\step1.myadd.fa4.cout ),
    .Y(_99_)
);

NOR2X1 _1058_ (
    .A(\step1.myadd.fa5.i1 ),
    .B(\step1.myadd.fa4.cout ),
    .Y(_100_)
);

OAI21X1 _1059_ (
    .A(_100_),
    .B(_99_),
    .C(gnd),
    .Y(_101_)
);

INVX1 _1060_ (
    .A(gnd),
    .Y(_102_)
);

NAND2X1 _1061_ (
    .A(\step1.myadd.fa5.i1 ),
    .B(\step1.myadd.fa4.cout ),
    .Y(_96_)
);

OR2X2 _1062_ (
    .A(\step1.myadd.fa5.i1 ),
    .B(\step1.myadd.fa4.cout ),
    .Y(_97_)
);

NAND3X1 _1063_ (
    .A(_102_),
    .B(_96_),
    .C(_97_),
    .Y(_98_)
);

NAND2X1 _1064_ (
    .A(_101_),
    .B(_98_),
    .Y(\step1.myadd.fa5.sum )
);

AOI21X1 _1065_ (
    .A(_102_),
    .B(_96_),
    .C(_100_),
    .Y(\step1.myadd.fa5.cout )
);

AND2X2 _1066_ (
    .A(\step1.myadd.fa6.i1 ),
    .B(\step1.myadd.fa5.cout ),
    .Y(_106_)
);

NOR2X1 _1067_ (
    .A(\step1.myadd.fa6.i1 ),
    .B(\step1.myadd.fa5.cout ),
    .Y(_107_)
);

OAI21X1 _1068_ (
    .A(_107_),
    .B(_106_),
    .C(gnd),
    .Y(_108_)
);

INVX1 _1069_ (
    .A(gnd),
    .Y(_109_)
);

NAND2X1 _1070_ (
    .A(\step1.myadd.fa6.i1 ),
    .B(\step1.myadd.fa5.cout ),
    .Y(_103_)
);

OR2X2 _1071_ (
    .A(\step1.myadd.fa6.i1 ),
    .B(\step1.myadd.fa5.cout ),
    .Y(_104_)
);

NAND3X1 _1072_ (
    .A(_109_),
    .B(_103_),
    .C(_104_),
    .Y(_105_)
);

NAND2X1 _1073_ (
    .A(_108_),
    .B(_105_),
    .Y(\step1.myadd.fa6.sum )
);

AOI21X1 _1074_ (
    .A(_109_),
    .B(_103_),
    .C(_107_),
    .Y(\step1.myadd.fa6.cout )
);

AND2X2 _1075_ (
    .A(\step1.myadd.fa7.i1 ),
    .B(\step1.myadd.fa6.cout ),
    .Y(_113_)
);

NOR2X1 _1076_ (
    .A(\step1.myadd.fa7.i1 ),
    .B(\step1.myadd.fa6.cout ),
    .Y(_114_)
);

OAI21X1 _1077_ (
    .A(_114_),
    .B(_113_),
    .C(gnd),
    .Y(_115_)
);

INVX1 _1078_ (
    .A(gnd),
    .Y(_116_)
);

NAND2X1 _1079_ (
    .A(\step1.myadd.fa7.i1 ),
    .B(\step1.myadd.fa6.cout ),
    .Y(_110_)
);

OR2X2 _1080_ (
    .A(\step1.myadd.fa7.i1 ),
    .B(\step1.myadd.fa6.cout ),
    .Y(_111_)
);

NAND3X1 _1081_ (
    .A(_116_),
    .B(_110_),
    .C(_111_),
    .Y(_112_)
);

NAND2X1 _1082_ (
    .A(_115_),
    .B(_112_),
    .Y(\step1.myadd.fa7.sum )
);

AOI21X1 _1083_ (
    .A(_116_),
    .B(_110_),
    .C(_114_),
    .Y(\step1.myadd.fa7.cout )
);

AND2X2 _1084_ (
    .A(\step1.myadd.fa8.i1 ),
    .B(\step1.myadd.fa7.cout ),
    .Y(_120_)
);

NOR2X1 _1085_ (
    .A(\step1.myadd.fa8.i1 ),
    .B(\step1.myadd.fa7.cout ),
    .Y(_121_)
);

OAI21X1 _1086_ (
    .A(_121_),
    .B(_120_),
    .C(gnd),
    .Y(_122_)
);

INVX1 _1087_ (
    .A(gnd),
    .Y(_123_)
);

NAND2X1 _1088_ (
    .A(\step1.myadd.fa8.i1 ),
    .B(\step1.myadd.fa7.cout ),
    .Y(_117_)
);

OR2X2 _1089_ (
    .A(\step1.myadd.fa8.i1 ),
    .B(\step1.myadd.fa7.cout ),
    .Y(_118_)
);

NAND3X1 _1090_ (
    .A(_123_),
    .B(_117_),
    .C(_118_),
    .Y(_119_)
);

NAND2X1 _1091_ (
    .A(_122_),
    .B(_119_),
    .Y(\step1.myadd.fa8.sum )
);

INVX1 _1092_ (
    .A(\step1.myadd.cin_bF$buf0 ),
    .Y(_124_)
);

NAND2X1 _1093_ (
    .A(\step1.myadd.x0.i0_bF$buf3 ),
    .B(_124_),
    .Y(_125_)
);

INVX1 _1094_ (
    .A(\step1.myadd.x0.i0_bF$buf2 ),
    .Y(_126_)
);

NAND2X1 _1095_ (
    .A(\step1.myadd.cin_bF$buf4 ),
    .B(_126_),
    .Y(_127_)
);

NAND2X1 _1096_ (
    .A(_125_),
    .B(_127_),
    .Y(\step1.myadd.fa1.i1 )
);

INVX1 _1097_ (
    .A(\step1.myadd.cin_bF$buf3 ),
    .Y(_128_)
);

NAND2X1 _1098_ (
    .A(\step1.myadd.x1.i0_bF$buf3 ),
    .B(_128_),
    .Y(_129_)
);

INVX1 _1099_ (
    .A(\step1.myadd.x1.i0_bF$buf2 ),
    .Y(_130_)
);

NAND2X1 _1100_ (
    .A(\step1.myadd.cin_bF$buf2 ),
    .B(_130_),
    .Y(_131_)
);

NAND2X1 _1101_ (
    .A(_129_),
    .B(_131_),
    .Y(\step1.myadd.fa2.i1 )
);

INVX1 _1102_ (
    .A(\step1.myadd.cin_bF$buf1 ),
    .Y(_132_)
);

NAND2X1 _1103_ (
    .A(\step1.myadd.x2.i0_bF$buf3 ),
    .B(_132_),
    .Y(_133_)
);

INVX1 _1104_ (
    .A(\step1.myadd.x2.i0_bF$buf2 ),
    .Y(_134_)
);

NAND2X1 _1105_ (
    .A(\step1.myadd.cin_bF$buf0 ),
    .B(_134_),
    .Y(_135_)
);

NAND2X1 _1106_ (
    .A(_133_),
    .B(_135_),
    .Y(\step1.myadd.fa3.i1 )
);

INVX1 _1107_ (
    .A(\step1.myadd.cin_bF$buf4 ),
    .Y(_136_)
);

NAND2X1 _1108_ (
    .A(\step1.myadd.x3.i0_bF$buf3 ),
    .B(_136_),
    .Y(_137_)
);

INVX1 _1109_ (
    .A(\step1.myadd.x3.i0_bF$buf2 ),
    .Y(_138_)
);

NAND2X1 _1110_ (
    .A(\step1.myadd.cin_bF$buf3 ),
    .B(_138_),
    .Y(_139_)
);

NAND2X1 _1111_ (
    .A(_137_),
    .B(_139_),
    .Y(\step1.myadd.fa4.i1 )
);

INVX1 _1112_ (
    .A(\step1.myadd.cin_bF$buf2 ),
    .Y(_140_)
);

NAND2X1 _1113_ (
    .A(\step1.myadd.x4.i0_bF$buf3 ),
    .B(_140_),
    .Y(_141_)
);

INVX1 _1114_ (
    .A(\step1.myadd.x4.i0_bF$buf2 ),
    .Y(_142_)
);

NAND2X1 _1115_ (
    .A(\step1.myadd.cin_bF$buf1 ),
    .B(_142_),
    .Y(_143_)
);

NAND2X1 _1116_ (
    .A(_141_),
    .B(_143_),
    .Y(\step1.myadd.fa5.i1 )
);

INVX1 _1117_ (
    .A(\step1.myadd.cin_bF$buf0 ),
    .Y(_144_)
);

NAND2X1 _1118_ (
    .A(\step1.myadd.x5.i0_bF$buf3 ),
    .B(_144_),
    .Y(_145_)
);

INVX1 _1119_ (
    .A(\step1.myadd.x5.i0_bF$buf2 ),
    .Y(_146_)
);

NAND2X1 _1120_ (
    .A(\step1.myadd.cin_bF$buf4 ),
    .B(_146_),
    .Y(_147_)
);

NAND2X1 _1121_ (
    .A(_145_),
    .B(_147_),
    .Y(\step1.myadd.fa6.i1 )
);

INVX1 _1122_ (
    .A(\step1.myadd.cin_bF$buf3 ),
    .Y(_148_)
);

NAND2X1 _1123_ (
    .A(\step1.myadd.x6.i0_bF$buf3 ),
    .B(_148_),
    .Y(_149_)
);

INVX1 _1124_ (
    .A(\step1.myadd.x6.i0_bF$buf2 ),
    .Y(_150_)
);

NAND2X1 _1125_ (
    .A(\step1.myadd.cin_bF$buf2 ),
    .B(_150_),
    .Y(_151_)
);

NAND2X1 _1126_ (
    .A(_149_),
    .B(_151_),
    .Y(\step1.myadd.fa7.i1 )
);

INVX1 _1127_ (
    .A(\step1.myadd.cin_bF$buf1 ),
    .Y(_152_)
);

NAND2X1 _1128_ (
    .A(\step1.myadd.x7.i0_bF$buf3 ),
    .B(_152_),
    .Y(_153_)
);

INVX1 _1129_ (
    .A(\step1.myadd.x7.i0_bF$buf2 ),
    .Y(_154_)
);

NAND2X1 _1130_ (
    .A(\step1.myadd.cin_bF$buf0 ),
    .B(_154_),
    .Y(_155_)
);

NAND2X1 _1131_ (
    .A(_153_),
    .B(_155_),
    .Y(\step1.myadd.fa8.i1 )
);

OR2X2 _1132_ (
    .A(\step1.myadd.cin_bF$buf4 ),
    .B(\step2.myadd.cin_bF$buf4 ),
    .Y(_156_)
);

NAND2X1 _1133_ (
    .A(\step1.myadd.cin_bF$buf3 ),
    .B(\step2.myadd.cin_bF$buf3 ),
    .Y(_157_)
);

NAND3X1 _1134_ (
    .A(\step2.myadd.fa2.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_158_)
);

NOR2X1 _1135_ (
    .A(\step1.myadd.cin_bF$buf2 ),
    .B(\step2.myadd.cin_bF$buf2 ),
    .Y(_159_)
);

AND2X2 _1136_ (
    .A(\step1.myadd.cin_bF$buf1 ),
    .B(\step2.myadd.cin_bF$buf1 ),
    .Y(_160_)
);

OAI21X1 _1137_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa2.i0 ),
    .Y(_161_)
);

NAND2X1 _1138_ (
    .A(_161_),
    .B(_158_),
    .Y(\step3.myadd.fa1.i0 )
);

NAND3X1 _1139_ (
    .A(\step2.myadd.fa3.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_162_)
);

OAI21X1 _1140_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa3.i0 ),
    .Y(_163_)
);

NAND2X1 _1141_ (
    .A(_163_),
    .B(_162_),
    .Y(\step3.myadd.fa2.i0 )
);

NAND3X1 _1142_ (
    .A(\step2.myadd.fa4.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_164_)
);

OAI21X1 _1143_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa4.i0 ),
    .Y(_165_)
);

NAND2X1 _1144_ (
    .A(_165_),
    .B(_164_),
    .Y(\step3.myadd.fa3.i0 )
);

NAND3X1 _1145_ (
    .A(\step2.myadd.fa5.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_166_)
);

OAI21X1 _1146_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa5.i0 ),
    .Y(_167_)
);

NAND2X1 _1147_ (
    .A(_167_),
    .B(_166_),
    .Y(\step3.myadd.fa4.i0 )
);

NAND3X1 _1148_ (
    .A(\step2.myadd.fa6.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_168_)
);

OAI21X1 _1149_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa6.i0 ),
    .Y(_169_)
);

NAND2X1 _1150_ (
    .A(_169_),
    .B(_168_),
    .Y(\step3.myadd.fa5.i0 )
);

NAND3X1 _1151_ (
    .A(\step2.myadd.fa7.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_170_)
);

OAI21X1 _1152_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa7.i0 ),
    .Y(_171_)
);

NAND2X1 _1153_ (
    .A(_171_),
    .B(_170_),
    .Y(\step3.myadd.fa6.i0 )
);

NAND3X1 _1154_ (
    .A(\step2.myadd.fa8.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_172_)
);

OAI21X1 _1155_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa7.i0 ),
    .Y(_173_)
);

NAND2X1 _1156_ (
    .A(_173_),
    .B(_172_),
    .Y(\step3.myadd.fa7.i0 )
);

NAND3X1 _1157_ (
    .A(\step2.myadd.fa1.sum ),
    .B(_157_),
    .C(_156_),
    .Y(_174_)
);

OAI21X1 _1158_ (
    .A(_159_),
    .B(_160_),
    .C(\step2.myadd.fa1.i0 ),
    .Y(_175_)
);

NAND2X1 _1159_ (
    .A(_175_),
    .B(_174_),
    .Y(\Q[1] [7])
);

AND2X2 _1160_ (
    .A(\step2.myadd.fa1.i1 ),
    .B(\step2.myadd.cin_bF$buf0 ),
    .Y(_179_)
);

NOR2X1 _1161_ (
    .A(\step2.myadd.fa1.i1 ),
    .B(\step2.myadd.cin_bF$buf4 ),
    .Y(_180_)
);

OAI21X1 _1162_ (
    .A(_180_),
    .B(_179_),
    .C(\step2.myadd.fa1.i0 ),
    .Y(_181_)
);

INVX1 _1163_ (
    .A(\step2.myadd.fa1.i0 ),
    .Y(_182_)
);

NAND2X1 _1164_ (
    .A(\step2.myadd.fa1.i1 ),
    .B(\step2.myadd.cin_bF$buf3 ),
    .Y(_176_)
);

OR2X2 _1165_ (
    .A(\step2.myadd.fa1.i1 ),
    .B(\step2.myadd.cin_bF$buf2 ),
    .Y(_177_)
);

NAND3X1 _1166_ (
    .A(_182_),
    .B(_176_),
    .C(_177_),
    .Y(_178_)
);

NAND2X1 _1167_ (
    .A(_181_),
    .B(_178_),
    .Y(\step2.myadd.fa1.sum )
);

AOI21X1 _1168_ (
    .A(_182_),
    .B(_176_),
    .C(_180_),
    .Y(\step2.myadd.fa1.cout )
);

AND2X2 _1169_ (
    .A(\step2.myadd.fa2.i1 ),
    .B(\step2.myadd.fa1.cout ),
    .Y(_186_)
);

NOR2X1 _1170_ (
    .A(\step2.myadd.fa2.i1 ),
    .B(\step2.myadd.fa1.cout ),
    .Y(_187_)
);

OAI21X1 _1171_ (
    .A(_187_),
    .B(_186_),
    .C(\step2.myadd.fa2.i0 ),
    .Y(_188_)
);

INVX1 _1172_ (
    .A(\step2.myadd.fa2.i0 ),
    .Y(_189_)
);

NAND2X1 _1173_ (
    .A(\step2.myadd.fa2.i1 ),
    .B(\step2.myadd.fa1.cout ),
    .Y(_183_)
);

OR2X2 _1174_ (
    .A(\step2.myadd.fa2.i1 ),
    .B(\step2.myadd.fa1.cout ),
    .Y(_184_)
);

NAND3X1 _1175_ (
    .A(_189_),
    .B(_183_),
    .C(_184_),
    .Y(_185_)
);

NAND2X1 _1176_ (
    .A(_188_),
    .B(_185_),
    .Y(\step2.myadd.fa2.sum )
);

AOI21X1 _1177_ (
    .A(_189_),
    .B(_183_),
    .C(_187_),
    .Y(\step2.myadd.fa2.cout )
);

AND2X2 _1178_ (
    .A(\step2.myadd.fa3.i1 ),
    .B(\step2.myadd.fa2.cout ),
    .Y(_193_)
);

NOR2X1 _1179_ (
    .A(\step2.myadd.fa3.i1 ),
    .B(\step2.myadd.fa2.cout ),
    .Y(_194_)
);

OAI21X1 _1180_ (
    .A(_194_),
    .B(_193_),
    .C(\step2.myadd.fa3.i0 ),
    .Y(_195_)
);

INVX1 _1181_ (
    .A(\step2.myadd.fa3.i0 ),
    .Y(_196_)
);

NAND2X1 _1182_ (
    .A(\step2.myadd.fa3.i1 ),
    .B(\step2.myadd.fa2.cout ),
    .Y(_190_)
);

OR2X2 _1183_ (
    .A(\step2.myadd.fa3.i1 ),
    .B(\step2.myadd.fa2.cout ),
    .Y(_191_)
);

NAND3X1 _1184_ (
    .A(_196_),
    .B(_190_),
    .C(_191_),
    .Y(_192_)
);

NAND2X1 _1185_ (
    .A(_195_),
    .B(_192_),
    .Y(\step2.myadd.fa3.sum )
);

AOI21X1 _1186_ (
    .A(_196_),
    .B(_190_),
    .C(_194_),
    .Y(\step2.myadd.fa3.cout )
);

AND2X2 _1187_ (
    .A(\step2.myadd.fa4.i1 ),
    .B(\step2.myadd.fa3.cout ),
    .Y(_200_)
);

NOR2X1 _1188_ (
    .A(\step2.myadd.fa4.i1 ),
    .B(\step2.myadd.fa3.cout ),
    .Y(_201_)
);

OAI21X1 _1189_ (
    .A(_201_),
    .B(_200_),
    .C(\step2.myadd.fa4.i0 ),
    .Y(_202_)
);

INVX1 _1190_ (
    .A(\step2.myadd.fa4.i0 ),
    .Y(_203_)
);

NAND2X1 _1191_ (
    .A(\step2.myadd.fa4.i1 ),
    .B(\step2.myadd.fa3.cout ),
    .Y(_197_)
);

OR2X2 _1192_ (
    .A(\step2.myadd.fa4.i1 ),
    .B(\step2.myadd.fa3.cout ),
    .Y(_198_)
);

NAND3X1 _1193_ (
    .A(_203_),
    .B(_197_),
    .C(_198_),
    .Y(_199_)
);

NAND2X1 _1194_ (
    .A(_202_),
    .B(_199_),
    .Y(\step2.myadd.fa4.sum )
);

AOI21X1 _1195_ (
    .A(_203_),
    .B(_197_),
    .C(_201_),
    .Y(\step2.myadd.fa4.cout )
);

AND2X2 _1196_ (
    .A(\step2.myadd.fa5.i1 ),
    .B(\step2.myadd.fa4.cout ),
    .Y(_207_)
);

NOR2X1 _1197_ (
    .A(\step2.myadd.fa5.i1 ),
    .B(\step2.myadd.fa4.cout ),
    .Y(_208_)
);

OAI21X1 _1198_ (
    .A(_208_),
    .B(_207_),
    .C(\step2.myadd.fa5.i0 ),
    .Y(_209_)
);

INVX1 _1199_ (
    .A(\step2.myadd.fa5.i0 ),
    .Y(_210_)
);

NAND2X1 _1200_ (
    .A(\step2.myadd.fa5.i1 ),
    .B(\step2.myadd.fa4.cout ),
    .Y(_204_)
);

OR2X2 _1201_ (
    .A(\step2.myadd.fa5.i1 ),
    .B(\step2.myadd.fa4.cout ),
    .Y(_205_)
);

NAND3X1 _1202_ (
    .A(_210_),
    .B(_204_),
    .C(_205_),
    .Y(_206_)
);

NAND2X1 _1203_ (
    .A(_209_),
    .B(_206_),
    .Y(\step2.myadd.fa5.sum )
);

AOI21X1 _1204_ (
    .A(_210_),
    .B(_204_),
    .C(_208_),
    .Y(\step2.myadd.fa5.cout )
);

AND2X2 _1205_ (
    .A(\step2.myadd.fa6.i1 ),
    .B(\step2.myadd.fa5.cout ),
    .Y(_214_)
);

NOR2X1 _1206_ (
    .A(\step2.myadd.fa6.i1 ),
    .B(\step2.myadd.fa5.cout ),
    .Y(_215_)
);

OAI21X1 _1207_ (
    .A(_215_),
    .B(_214_),
    .C(\step2.myadd.fa6.i0 ),
    .Y(_216_)
);

INVX1 _1208_ (
    .A(\step2.myadd.fa6.i0 ),
    .Y(_217_)
);

NAND2X1 _1209_ (
    .A(\step2.myadd.fa6.i1 ),
    .B(\step2.myadd.fa5.cout ),
    .Y(_211_)
);

OR2X2 _1210_ (
    .A(\step2.myadd.fa6.i1 ),
    .B(\step2.myadd.fa5.cout ),
    .Y(_212_)
);

NAND3X1 _1211_ (
    .A(_217_),
    .B(_211_),
    .C(_212_),
    .Y(_213_)
);

NAND2X1 _1212_ (
    .A(_216_),
    .B(_213_),
    .Y(\step2.myadd.fa6.sum )
);

AOI21X1 _1213_ (
    .A(_217_),
    .B(_211_),
    .C(_215_),
    .Y(\step2.myadd.fa6.cout )
);

AND2X2 _1214_ (
    .A(\step2.myadd.fa7.i1 ),
    .B(\step2.myadd.fa6.cout ),
    .Y(_221_)
);

NOR2X1 _1215_ (
    .A(\step2.myadd.fa7.i1 ),
    .B(\step2.myadd.fa6.cout ),
    .Y(_222_)
);

OAI21X1 _1216_ (
    .A(_222_),
    .B(_221_),
    .C(\step2.myadd.fa7.i0 ),
    .Y(_223_)
);

INVX1 _1217_ (
    .A(\step2.myadd.fa7.i0 ),
    .Y(_224_)
);

NAND2X1 _1218_ (
    .A(\step2.myadd.fa7.i1 ),
    .B(\step2.myadd.fa6.cout ),
    .Y(_218_)
);

OR2X2 _1219_ (
    .A(\step2.myadd.fa7.i1 ),
    .B(\step2.myadd.fa6.cout ),
    .Y(_219_)
);

NAND3X1 _1220_ (
    .A(_224_),
    .B(_218_),
    .C(_219_),
    .Y(_220_)
);

NAND2X1 _1221_ (
    .A(_223_),
    .B(_220_),
    .Y(\step2.myadd.fa7.sum )
);

AOI21X1 _1222_ (
    .A(_224_),
    .B(_218_),
    .C(_222_),
    .Y(\step2.myadd.fa7.cout )
);

AND2X2 _1223_ (
    .A(\step2.myadd.fa8.i1 ),
    .B(\step2.myadd.fa7.cout ),
    .Y(_228_)
);

NOR2X1 _1224_ (
    .A(\step2.myadd.fa8.i1 ),
    .B(\step2.myadd.fa7.cout ),
    .Y(_229_)
);

OAI21X1 _1225_ (
    .A(_229_),
    .B(_228_),
    .C(\step2.myadd.fa7.i0 ),
    .Y(_230_)
);

INVX1 _1226_ (
    .A(\step2.myadd.fa7.i0 ),
    .Y(_231_)
);

NAND2X1 _1227_ (
    .A(\step2.myadd.fa8.i1 ),
    .B(\step2.myadd.fa7.cout ),
    .Y(_225_)
);

OR2X2 _1228_ (
    .A(\step2.myadd.fa8.i1 ),
    .B(\step2.myadd.fa7.cout ),
    .Y(_226_)
);

NAND3X1 _1229_ (
    .A(_231_),
    .B(_225_),
    .C(_226_),
    .Y(_227_)
);

NAND2X1 _1230_ (
    .A(_230_),
    .B(_227_),
    .Y(\step2.myadd.fa8.sum )
);

INVX1 _1231_ (
    .A(\step2.myadd.cin_bF$buf1 ),
    .Y(_232_)
);

NAND2X1 _1232_ (
    .A(\step1.myadd.x0.i0_bF$buf1 ),
    .B(_232_),
    .Y(_233_)
);

INVX1 _1233_ (
    .A(\step1.myadd.x0.i0_bF$buf0 ),
    .Y(_234_)
);

NAND2X1 _1234_ (
    .A(\step2.myadd.cin_bF$buf0 ),
    .B(_234_),
    .Y(_235_)
);

NAND2X1 _1235_ (
    .A(_233_),
    .B(_235_),
    .Y(\step2.myadd.fa1.i1 )
);

INVX1 _1236_ (
    .A(\step2.myadd.cin_bF$buf4 ),
    .Y(_236_)
);

NAND2X1 _1237_ (
    .A(\step1.myadd.x1.i0_bF$buf1 ),
    .B(_236_),
    .Y(_237_)
);

INVX1 _1238_ (
    .A(\step1.myadd.x1.i0_bF$buf0 ),
    .Y(_238_)
);

NAND2X1 _1239_ (
    .A(\step2.myadd.cin_bF$buf3 ),
    .B(_238_),
    .Y(_239_)
);

NAND2X1 _1240_ (
    .A(_237_),
    .B(_239_),
    .Y(\step2.myadd.fa2.i1 )
);

INVX1 _1241_ (
    .A(\step2.myadd.cin_bF$buf2 ),
    .Y(_240_)
);

NAND2X1 _1242_ (
    .A(\step1.myadd.x2.i0_bF$buf1 ),
    .B(_240_),
    .Y(_241_)
);

INVX1 _1243_ (
    .A(\step1.myadd.x2.i0_bF$buf0 ),
    .Y(_242_)
);

NAND2X1 _1244_ (
    .A(\step2.myadd.cin_bF$buf1 ),
    .B(_242_),
    .Y(_243_)
);

NAND2X1 _1245_ (
    .A(_241_),
    .B(_243_),
    .Y(\step2.myadd.fa3.i1 )
);

INVX1 _1246_ (
    .A(\step2.myadd.cin_bF$buf0 ),
    .Y(_244_)
);

NAND2X1 _1247_ (
    .A(\step1.myadd.x3.i0_bF$buf1 ),
    .B(_244_),
    .Y(_245_)
);

INVX1 _1248_ (
    .A(\step1.myadd.x3.i0_bF$buf0 ),
    .Y(_246_)
);

NAND2X1 _1249_ (
    .A(\step2.myadd.cin_bF$buf4 ),
    .B(_246_),
    .Y(_247_)
);

NAND2X1 _1250_ (
    .A(_245_),
    .B(_247_),
    .Y(\step2.myadd.fa4.i1 )
);

INVX1 _1251_ (
    .A(\step2.myadd.cin_bF$buf3 ),
    .Y(_248_)
);

NAND2X1 _1252_ (
    .A(\step1.myadd.x4.i0_bF$buf1 ),
    .B(_248_),
    .Y(_249_)
);

INVX1 _1253_ (
    .A(\step1.myadd.x4.i0_bF$buf0 ),
    .Y(_250_)
);

NAND2X1 _1254_ (
    .A(\step2.myadd.cin_bF$buf2 ),
    .B(_250_),
    .Y(_251_)
);

NAND2X1 _1255_ (
    .A(_249_),
    .B(_251_),
    .Y(\step2.myadd.fa5.i1 )
);

INVX1 _1256_ (
    .A(\step2.myadd.cin_bF$buf1 ),
    .Y(_252_)
);

NAND2X1 _1257_ (
    .A(\step1.myadd.x5.i0_bF$buf1 ),
    .B(_252_),
    .Y(_253_)
);

INVX1 _1258_ (
    .A(\step1.myadd.x5.i0_bF$buf0 ),
    .Y(_254_)
);

NAND2X1 _1259_ (
    .A(\step2.myadd.cin_bF$buf0 ),
    .B(_254_),
    .Y(_255_)
);

NAND2X1 _1260_ (
    .A(_253_),
    .B(_255_),
    .Y(\step2.myadd.fa6.i1 )
);

INVX1 _1261_ (
    .A(\step2.myadd.cin_bF$buf4 ),
    .Y(_256_)
);

NAND2X1 _1262_ (
    .A(\step1.myadd.x6.i0_bF$buf1 ),
    .B(_256_),
    .Y(_257_)
);

INVX1 _1263_ (
    .A(\step1.myadd.x6.i0_bF$buf0 ),
    .Y(_258_)
);

NAND2X1 _1264_ (
    .A(\step2.myadd.cin_bF$buf3 ),
    .B(_258_),
    .Y(_259_)
);

NAND2X1 _1265_ (
    .A(_257_),
    .B(_259_),
    .Y(\step2.myadd.fa7.i1 )
);

INVX1 _1266_ (
    .A(\step2.myadd.cin_bF$buf2 ),
    .Y(_260_)
);

NAND2X1 _1267_ (
    .A(\step1.myadd.x7.i0_bF$buf1 ),
    .B(_260_),
    .Y(_261_)
);

INVX1 _1268_ (
    .A(\step1.myadd.x7.i0_bF$buf0 ),
    .Y(_262_)
);

NAND2X1 _1269_ (
    .A(\step2.myadd.cin_bF$buf1 ),
    .B(_262_),
    .Y(_263_)
);

NAND2X1 _1270_ (
    .A(_261_),
    .B(_263_),
    .Y(\step2.myadd.fa8.i1 )
);

OR2X2 _1271_ (
    .A(\step2.myadd.cin_bF$buf0 ),
    .B(\step3.myadd.cin_bF$buf4 ),
    .Y(_264_)
);

NAND2X1 _1272_ (
    .A(\step2.myadd.cin_bF$buf4 ),
    .B(\step3.myadd.cin_bF$buf3 ),
    .Y(_265_)
);

NAND3X1 _1273_ (
    .A(\step3.myadd.fa2.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_266_)
);

NOR2X1 _1274_ (
    .A(\step2.myadd.cin_bF$buf3 ),
    .B(\step3.myadd.cin_bF$buf2 ),
    .Y(_267_)
);

AND2X2 _1275_ (
    .A(\step2.myadd.cin_bF$buf2 ),
    .B(\step3.myadd.cin_bF$buf1 ),
    .Y(_268_)
);

OAI21X1 _1276_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa2.i0 ),
    .Y(_269_)
);

NAND2X1 _1277_ (
    .A(_269_),
    .B(_266_),
    .Y(\step4.myadd.fa1.i0 )
);

NAND3X1 _1278_ (
    .A(\step3.myadd.fa3.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_270_)
);

OAI21X1 _1279_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa3.i0 ),
    .Y(_271_)
);

NAND2X1 _1280_ (
    .A(_271_),
    .B(_270_),
    .Y(\step4.myadd.fa2.i0 )
);

NAND3X1 _1281_ (
    .A(\step3.myadd.fa4.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_272_)
);

OAI21X1 _1282_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa4.i0 ),
    .Y(_273_)
);

NAND2X1 _1283_ (
    .A(_273_),
    .B(_272_),
    .Y(\step4.myadd.fa3.i0 )
);

NAND3X1 _1284_ (
    .A(\step3.myadd.fa5.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_274_)
);

OAI21X1 _1285_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa5.i0 ),
    .Y(_275_)
);

NAND2X1 _1286_ (
    .A(_275_),
    .B(_274_),
    .Y(\step4.myadd.fa4.i0 )
);

NAND3X1 _1287_ (
    .A(\step3.myadd.fa6.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_276_)
);

OAI21X1 _1288_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa6.i0 ),
    .Y(_277_)
);

NAND2X1 _1289_ (
    .A(_277_),
    .B(_276_),
    .Y(\step4.myadd.fa5.i0 )
);

NAND3X1 _1290_ (
    .A(\step3.myadd.fa7.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_278_)
);

OAI21X1 _1291_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa7.i0 ),
    .Y(_279_)
);

NAND2X1 _1292_ (
    .A(_279_),
    .B(_278_),
    .Y(\step4.myadd.fa6.i0 )
);

NAND3X1 _1293_ (
    .A(\step3.myadd.fa8.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_280_)
);

OAI21X1 _1294_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa7.i0 ),
    .Y(_281_)
);

NAND2X1 _1295_ (
    .A(_281_),
    .B(_280_),
    .Y(\step4.myadd.fa7.i0 )
);

NAND3X1 _1296_ (
    .A(\step3.myadd.fa1.sum ),
    .B(_265_),
    .C(_264_),
    .Y(_282_)
);

OAI21X1 _1297_ (
    .A(_267_),
    .B(_268_),
    .C(\step3.myadd.fa1.i0 ),
    .Y(_283_)
);

NAND2X1 _1298_ (
    .A(_283_),
    .B(_282_),
    .Y(\Q[2] [7])
);

AND2X2 _1299_ (
    .A(\step3.myadd.fa1.i1 ),
    .B(\step3.myadd.cin_bF$buf0 ),
    .Y(_287_)
);

NOR2X1 _1300_ (
    .A(\step3.myadd.fa1.i1 ),
    .B(\step3.myadd.cin_bF$buf4 ),
    .Y(_288_)
);

OAI21X1 _1301_ (
    .A(_288_),
    .B(_287_),
    .C(\step3.myadd.fa1.i0 ),
    .Y(_289_)
);

INVX1 _1302_ (
    .A(\step3.myadd.fa1.i0 ),
    .Y(_290_)
);

NAND2X1 _1303_ (
    .A(\step3.myadd.fa1.i1 ),
    .B(\step3.myadd.cin_bF$buf3 ),
    .Y(_284_)
);

OR2X2 _1304_ (
    .A(\step3.myadd.fa1.i1 ),
    .B(\step3.myadd.cin_bF$buf2 ),
    .Y(_285_)
);

NAND3X1 _1305_ (
    .A(_290_),
    .B(_284_),
    .C(_285_),
    .Y(_286_)
);

NAND2X1 _1306_ (
    .A(_289_),
    .B(_286_),
    .Y(\step3.myadd.fa1.sum )
);

AOI21X1 _1307_ (
    .A(_290_),
    .B(_284_),
    .C(_288_),
    .Y(\step3.myadd.fa1.cout )
);

AND2X2 _1308_ (
    .A(\step3.myadd.fa2.i1 ),
    .B(\step3.myadd.fa1.cout ),
    .Y(_294_)
);

NOR2X1 _1309_ (
    .A(\step3.myadd.fa2.i1 ),
    .B(\step3.myadd.fa1.cout ),
    .Y(_295_)
);

OAI21X1 _1310_ (
    .A(_295_),
    .B(_294_),
    .C(\step3.myadd.fa2.i0 ),
    .Y(_296_)
);

INVX1 _1311_ (
    .A(\step3.myadd.fa2.i0 ),
    .Y(_297_)
);

NAND2X1 _1312_ (
    .A(\step3.myadd.fa2.i1 ),
    .B(\step3.myadd.fa1.cout ),
    .Y(_291_)
);

OR2X2 _1313_ (
    .A(\step3.myadd.fa2.i1 ),
    .B(\step3.myadd.fa1.cout ),
    .Y(_292_)
);

NAND3X1 _1314_ (
    .A(_297_),
    .B(_291_),
    .C(_292_),
    .Y(_293_)
);

NAND2X1 _1315_ (
    .A(_296_),
    .B(_293_),
    .Y(\step3.myadd.fa2.sum )
);

AOI21X1 _1316_ (
    .A(_297_),
    .B(_291_),
    .C(_295_),
    .Y(\step3.myadd.fa2.cout )
);

AND2X2 _1317_ (
    .A(\step3.myadd.fa3.i1 ),
    .B(\step3.myadd.fa2.cout ),
    .Y(_301_)
);

NOR2X1 _1318_ (
    .A(\step3.myadd.fa3.i1 ),
    .B(\step3.myadd.fa2.cout ),
    .Y(_302_)
);

OAI21X1 _1319_ (
    .A(_302_),
    .B(_301_),
    .C(\step3.myadd.fa3.i0 ),
    .Y(_303_)
);

INVX1 _1320_ (
    .A(\step3.myadd.fa3.i0 ),
    .Y(_304_)
);

NAND2X1 _1321_ (
    .A(\step3.myadd.fa3.i1 ),
    .B(\step3.myadd.fa2.cout ),
    .Y(_298_)
);

OR2X2 _1322_ (
    .A(\step3.myadd.fa3.i1 ),
    .B(\step3.myadd.fa2.cout ),
    .Y(_299_)
);

NAND3X1 _1323_ (
    .A(_304_),
    .B(_298_),
    .C(_299_),
    .Y(_300_)
);

NAND2X1 _1324_ (
    .A(_303_),
    .B(_300_),
    .Y(\step3.myadd.fa3.sum )
);

AOI21X1 _1325_ (
    .A(_304_),
    .B(_298_),
    .C(_302_),
    .Y(\step3.myadd.fa3.cout )
);

AND2X2 _1326_ (
    .A(\step3.myadd.fa4.i1 ),
    .B(\step3.myadd.fa3.cout ),
    .Y(_308_)
);

NOR2X1 _1327_ (
    .A(\step3.myadd.fa4.i1 ),
    .B(\step3.myadd.fa3.cout ),
    .Y(_309_)
);

OAI21X1 _1328_ (
    .A(_309_),
    .B(_308_),
    .C(\step3.myadd.fa4.i0 ),
    .Y(_310_)
);

INVX1 _1329_ (
    .A(\step3.myadd.fa4.i0 ),
    .Y(_311_)
);

NAND2X1 _1330_ (
    .A(\step3.myadd.fa4.i1 ),
    .B(\step3.myadd.fa3.cout ),
    .Y(_305_)
);

OR2X2 _1331_ (
    .A(\step3.myadd.fa4.i1 ),
    .B(\step3.myadd.fa3.cout ),
    .Y(_306_)
);

NAND3X1 _1332_ (
    .A(_311_),
    .B(_305_),
    .C(_306_),
    .Y(_307_)
);

NAND2X1 _1333_ (
    .A(_310_),
    .B(_307_),
    .Y(\step3.myadd.fa4.sum )
);

AOI21X1 _1334_ (
    .A(_311_),
    .B(_305_),
    .C(_309_),
    .Y(\step3.myadd.fa4.cout )
);

AND2X2 _1335_ (
    .A(\step3.myadd.fa5.i1 ),
    .B(\step3.myadd.fa4.cout ),
    .Y(_315_)
);

NOR2X1 _1336_ (
    .A(\step3.myadd.fa5.i1 ),
    .B(\step3.myadd.fa4.cout ),
    .Y(_316_)
);

OAI21X1 _1337_ (
    .A(_316_),
    .B(_315_),
    .C(\step3.myadd.fa5.i0 ),
    .Y(_317_)
);

INVX1 _1338_ (
    .A(\step3.myadd.fa5.i0 ),
    .Y(_318_)
);

NAND2X1 _1339_ (
    .A(\step3.myadd.fa5.i1 ),
    .B(\step3.myadd.fa4.cout ),
    .Y(_312_)
);

OR2X2 _1340_ (
    .A(\step3.myadd.fa5.i1 ),
    .B(\step3.myadd.fa4.cout ),
    .Y(_313_)
);

NAND3X1 _1341_ (
    .A(_318_),
    .B(_312_),
    .C(_313_),
    .Y(_314_)
);

NAND2X1 _1342_ (
    .A(_317_),
    .B(_314_),
    .Y(\step3.myadd.fa5.sum )
);

AOI21X1 _1343_ (
    .A(_318_),
    .B(_312_),
    .C(_316_),
    .Y(\step3.myadd.fa5.cout )
);

AND2X2 _1344_ (
    .A(\step3.myadd.fa6.i1 ),
    .B(\step3.myadd.fa5.cout ),
    .Y(_322_)
);

NOR2X1 _1345_ (
    .A(\step3.myadd.fa6.i1 ),
    .B(\step3.myadd.fa5.cout ),
    .Y(_323_)
);

OAI21X1 _1346_ (
    .A(_323_),
    .B(_322_),
    .C(\step3.myadd.fa6.i0 ),
    .Y(_324_)
);

INVX1 _1347_ (
    .A(\step3.myadd.fa6.i0 ),
    .Y(_325_)
);

NAND2X1 _1348_ (
    .A(\step3.myadd.fa6.i1 ),
    .B(\step3.myadd.fa5.cout ),
    .Y(_319_)
);

OR2X2 _1349_ (
    .A(\step3.myadd.fa6.i1 ),
    .B(\step3.myadd.fa5.cout ),
    .Y(_320_)
);

NAND3X1 _1350_ (
    .A(_325_),
    .B(_319_),
    .C(_320_),
    .Y(_321_)
);

NAND2X1 _1351_ (
    .A(_324_),
    .B(_321_),
    .Y(\step3.myadd.fa6.sum )
);

AOI21X1 _1352_ (
    .A(_325_),
    .B(_319_),
    .C(_323_),
    .Y(\step3.myadd.fa6.cout )
);

AND2X2 _1353_ (
    .A(\step3.myadd.fa7.i1 ),
    .B(\step3.myadd.fa6.cout ),
    .Y(_329_)
);

NOR2X1 _1354_ (
    .A(\step3.myadd.fa7.i1 ),
    .B(\step3.myadd.fa6.cout ),
    .Y(_330_)
);

OAI21X1 _1355_ (
    .A(_330_),
    .B(_329_),
    .C(\step3.myadd.fa7.i0 ),
    .Y(_331_)
);

INVX1 _1356_ (
    .A(\step3.myadd.fa7.i0 ),
    .Y(_332_)
);

NAND2X1 _1357_ (
    .A(\step3.myadd.fa7.i1 ),
    .B(\step3.myadd.fa6.cout ),
    .Y(_326_)
);

OR2X2 _1358_ (
    .A(\step3.myadd.fa7.i1 ),
    .B(\step3.myadd.fa6.cout ),
    .Y(_327_)
);

NAND3X1 _1359_ (
    .A(_332_),
    .B(_326_),
    .C(_327_),
    .Y(_328_)
);

NAND2X1 _1360_ (
    .A(_331_),
    .B(_328_),
    .Y(\step3.myadd.fa7.sum )
);

AOI21X1 _1361_ (
    .A(_332_),
    .B(_326_),
    .C(_330_),
    .Y(\step3.myadd.fa7.cout )
);

AND2X2 _1362_ (
    .A(\step3.myadd.fa8.i1 ),
    .B(\step3.myadd.fa7.cout ),
    .Y(_336_)
);

NOR2X1 _1363_ (
    .A(\step3.myadd.fa8.i1 ),
    .B(\step3.myadd.fa7.cout ),
    .Y(_337_)
);

OAI21X1 _1364_ (
    .A(_337_),
    .B(_336_),
    .C(\step3.myadd.fa7.i0 ),
    .Y(_338_)
);

INVX1 _1365_ (
    .A(\step3.myadd.fa7.i0 ),
    .Y(_339_)
);

NAND2X1 _1366_ (
    .A(\step3.myadd.fa8.i1 ),
    .B(\step3.myadd.fa7.cout ),
    .Y(_333_)
);

OR2X2 _1367_ (
    .A(\step3.myadd.fa8.i1 ),
    .B(\step3.myadd.fa7.cout ),
    .Y(_334_)
);

NAND3X1 _1368_ (
    .A(_339_),
    .B(_333_),
    .C(_334_),
    .Y(_335_)
);

NAND2X1 _1369_ (
    .A(_338_),
    .B(_335_),
    .Y(\step3.myadd.fa8.sum )
);

INVX1 _1370_ (
    .A(\step3.myadd.cin_bF$buf1 ),
    .Y(_340_)
);

NAND2X1 _1371_ (
    .A(\step1.myadd.x0.i0_bF$buf3 ),
    .B(_340_),
    .Y(_341_)
);

INVX1 _1372_ (
    .A(\step1.myadd.x0.i0_bF$buf2 ),
    .Y(_342_)
);

NAND2X1 _1373_ (
    .A(\step3.myadd.cin_bF$buf0 ),
    .B(_342_),
    .Y(_343_)
);

NAND2X1 _1374_ (
    .A(_341_),
    .B(_343_),
    .Y(\step3.myadd.fa1.i1 )
);

INVX1 _1375_ (
    .A(\step3.myadd.cin_bF$buf4 ),
    .Y(_344_)
);

NAND2X1 _1376_ (
    .A(\step1.myadd.x1.i0_bF$buf3 ),
    .B(_344_),
    .Y(_345_)
);

INVX1 _1377_ (
    .A(\step1.myadd.x1.i0_bF$buf2 ),
    .Y(_346_)
);

NAND2X1 _1378_ (
    .A(\step3.myadd.cin_bF$buf3 ),
    .B(_346_),
    .Y(_347_)
);

NAND2X1 _1379_ (
    .A(_345_),
    .B(_347_),
    .Y(\step3.myadd.fa2.i1 )
);

INVX1 _1380_ (
    .A(\step3.myadd.cin_bF$buf2 ),
    .Y(_348_)
);

NAND2X1 _1381_ (
    .A(\step1.myadd.x2.i0_bF$buf3 ),
    .B(_348_),
    .Y(_349_)
);

INVX1 _1382_ (
    .A(\step1.myadd.x2.i0_bF$buf2 ),
    .Y(_350_)
);

NAND2X1 _1383_ (
    .A(\step3.myadd.cin_bF$buf1 ),
    .B(_350_),
    .Y(_351_)
);

NAND2X1 _1384_ (
    .A(_349_),
    .B(_351_),
    .Y(\step3.myadd.fa3.i1 )
);

INVX1 _1385_ (
    .A(\step3.myadd.cin_bF$buf0 ),
    .Y(_352_)
);

NAND2X1 _1386_ (
    .A(\step1.myadd.x3.i0_bF$buf3 ),
    .B(_352_),
    .Y(_353_)
);

INVX1 _1387_ (
    .A(\step1.myadd.x3.i0_bF$buf2 ),
    .Y(_354_)
);

NAND2X1 _1388_ (
    .A(\step3.myadd.cin_bF$buf4 ),
    .B(_354_),
    .Y(_355_)
);

NAND2X1 _1389_ (
    .A(_353_),
    .B(_355_),
    .Y(\step3.myadd.fa4.i1 )
);

INVX1 _1390_ (
    .A(\step3.myadd.cin_bF$buf3 ),
    .Y(_356_)
);

NAND2X1 _1391_ (
    .A(\step1.myadd.x4.i0_bF$buf3 ),
    .B(_356_),
    .Y(_357_)
);

INVX1 _1392_ (
    .A(\step1.myadd.x4.i0_bF$buf2 ),
    .Y(_358_)
);

NAND2X1 _1393_ (
    .A(\step3.myadd.cin_bF$buf2 ),
    .B(_358_),
    .Y(_359_)
);

NAND2X1 _1394_ (
    .A(_357_),
    .B(_359_),
    .Y(\step3.myadd.fa5.i1 )
);

INVX1 _1395_ (
    .A(\step3.myadd.cin_bF$buf1 ),
    .Y(_360_)
);

NAND2X1 _1396_ (
    .A(\step1.myadd.x5.i0_bF$buf3 ),
    .B(_360_),
    .Y(_361_)
);

INVX1 _1397_ (
    .A(\step1.myadd.x5.i0_bF$buf2 ),
    .Y(_362_)
);

NAND2X1 _1398_ (
    .A(\step3.myadd.cin_bF$buf0 ),
    .B(_362_),
    .Y(_363_)
);

NAND2X1 _1399_ (
    .A(_361_),
    .B(_363_),
    .Y(\step3.myadd.fa6.i1 )
);

INVX1 _1400_ (
    .A(\step3.myadd.cin_bF$buf4 ),
    .Y(_364_)
);

NAND2X1 _1401_ (
    .A(\step1.myadd.x6.i0_bF$buf3 ),
    .B(_364_),
    .Y(_365_)
);

INVX1 _1402_ (
    .A(\step1.myadd.x6.i0_bF$buf2 ),
    .Y(_366_)
);

NAND2X1 _1403_ (
    .A(\step3.myadd.cin_bF$buf3 ),
    .B(_366_),
    .Y(_367_)
);

NAND2X1 _1404_ (
    .A(_365_),
    .B(_367_),
    .Y(\step3.myadd.fa7.i1 )
);

INVX1 _1405_ (
    .A(\step3.myadd.cin_bF$buf2 ),
    .Y(_368_)
);

NAND2X1 _1406_ (
    .A(\step1.myadd.x7.i0_bF$buf3 ),
    .B(_368_),
    .Y(_369_)
);

INVX1 _1407_ (
    .A(\step1.myadd.x7.i0_bF$buf2 ),
    .Y(_370_)
);

NAND2X1 _1408_ (
    .A(\step3.myadd.cin_bF$buf1 ),
    .B(_370_),
    .Y(_371_)
);

NAND2X1 _1409_ (
    .A(_369_),
    .B(_371_),
    .Y(\step3.myadd.fa8.i1 )
);

OR2X2 _1410_ (
    .A(\step3.myadd.cin_bF$buf0 ),
    .B(\step4.myadd.cin_bF$buf4 ),
    .Y(_372_)
);

NAND2X1 _1411_ (
    .A(\step3.myadd.cin_bF$buf4 ),
    .B(\step4.myadd.cin_bF$buf3 ),
    .Y(_373_)
);

NAND3X1 _1412_ (
    .A(\step4.myadd.fa2.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_374_)
);

NOR2X1 _1413_ (
    .A(\step3.myadd.cin_bF$buf3 ),
    .B(\step4.myadd.cin_bF$buf2 ),
    .Y(_375_)
);

AND2X2 _1414_ (
    .A(\step3.myadd.cin_bF$buf2 ),
    .B(\step4.myadd.cin_bF$buf1 ),
    .Y(_376_)
);

OAI21X1 _1415_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa2.i0 ),
    .Y(_377_)
);

NAND2X1 _1416_ (
    .A(_377_),
    .B(_374_),
    .Y(\step5.myadd.fa1.i0 )
);

NAND3X1 _1417_ (
    .A(\step4.myadd.fa3.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_378_)
);

OAI21X1 _1418_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa3.i0 ),
    .Y(_379_)
);

NAND2X1 _1419_ (
    .A(_379_),
    .B(_378_),
    .Y(\step5.myadd.fa2.i0 )
);

NAND3X1 _1420_ (
    .A(\step4.myadd.fa4.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_380_)
);

OAI21X1 _1421_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa4.i0 ),
    .Y(_381_)
);

NAND2X1 _1422_ (
    .A(_381_),
    .B(_380_),
    .Y(\step5.myadd.fa3.i0 )
);

NAND3X1 _1423_ (
    .A(\step4.myadd.fa5.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_382_)
);

OAI21X1 _1424_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa5.i0 ),
    .Y(_383_)
);

NAND2X1 _1425_ (
    .A(_383_),
    .B(_382_),
    .Y(\step5.myadd.fa4.i0 )
);

NAND3X1 _1426_ (
    .A(\step4.myadd.fa6.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_384_)
);

OAI21X1 _1427_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa6.i0 ),
    .Y(_385_)
);

NAND2X1 _1428_ (
    .A(_385_),
    .B(_384_),
    .Y(\step5.myadd.fa5.i0 )
);

NAND3X1 _1429_ (
    .A(\step4.myadd.fa7.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_386_)
);

OAI21X1 _1430_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa7.i0 ),
    .Y(_387_)
);

NAND2X1 _1431_ (
    .A(_387_),
    .B(_386_),
    .Y(\step5.myadd.fa6.i0 )
);

NAND3X1 _1432_ (
    .A(\step4.myadd.fa8.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_388_)
);

OAI21X1 _1433_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa7.i0 ),
    .Y(_389_)
);

NAND2X1 _1434_ (
    .A(_389_),
    .B(_388_),
    .Y(\step5.myadd.fa7.i0 )
);

NAND3X1 _1435_ (
    .A(\step4.myadd.fa1.sum ),
    .B(_373_),
    .C(_372_),
    .Y(_390_)
);

OAI21X1 _1436_ (
    .A(_375_),
    .B(_376_),
    .C(\step4.myadd.fa1.i0 ),
    .Y(_391_)
);

NAND2X1 _1437_ (
    .A(_391_),
    .B(_390_),
    .Y(\Q[3] [7])
);

AND2X2 _1438_ (
    .A(\step4.myadd.fa1.i1 ),
    .B(\step4.myadd.cin_bF$buf0 ),
    .Y(_395_)
);

NOR2X1 _1439_ (
    .A(\step4.myadd.fa1.i1 ),
    .B(\step4.myadd.cin_bF$buf4 ),
    .Y(_396_)
);

OAI21X1 _1440_ (
    .A(_396_),
    .B(_395_),
    .C(\step4.myadd.fa1.i0 ),
    .Y(_397_)
);

INVX1 _1441_ (
    .A(\step4.myadd.fa1.i0 ),
    .Y(_398_)
);

NAND2X1 _1442_ (
    .A(\step4.myadd.fa1.i1 ),
    .B(\step4.myadd.cin_bF$buf3 ),
    .Y(_392_)
);

OR2X2 _1443_ (
    .A(\step4.myadd.fa1.i1 ),
    .B(\step4.myadd.cin_bF$buf2 ),
    .Y(_393_)
);

NAND3X1 _1444_ (
    .A(_398_),
    .B(_392_),
    .C(_393_),
    .Y(_394_)
);

NAND2X1 _1445_ (
    .A(_397_),
    .B(_394_),
    .Y(\step4.myadd.fa1.sum )
);

AOI21X1 _1446_ (
    .A(_398_),
    .B(_392_),
    .C(_396_),
    .Y(\step4.myadd.fa1.cout )
);

AND2X2 _1447_ (
    .A(\step4.myadd.fa2.i1 ),
    .B(\step4.myadd.fa1.cout ),
    .Y(_402_)
);

NOR2X1 _1448_ (
    .A(\step4.myadd.fa2.i1 ),
    .B(\step4.myadd.fa1.cout ),
    .Y(_403_)
);

OAI21X1 _1449_ (
    .A(_403_),
    .B(_402_),
    .C(\step4.myadd.fa2.i0 ),
    .Y(_404_)
);

INVX1 _1450_ (
    .A(\step4.myadd.fa2.i0 ),
    .Y(_405_)
);

NAND2X1 _1451_ (
    .A(\step4.myadd.fa2.i1 ),
    .B(\step4.myadd.fa1.cout ),
    .Y(_399_)
);

OR2X2 _1452_ (
    .A(\step4.myadd.fa2.i1 ),
    .B(\step4.myadd.fa1.cout ),
    .Y(_400_)
);

NAND3X1 _1453_ (
    .A(_405_),
    .B(_399_),
    .C(_400_),
    .Y(_401_)
);

NAND2X1 _1454_ (
    .A(_404_),
    .B(_401_),
    .Y(\step4.myadd.fa2.sum )
);

AOI21X1 _1455_ (
    .A(_405_),
    .B(_399_),
    .C(_403_),
    .Y(\step4.myadd.fa2.cout )
);

AND2X2 _1456_ (
    .A(\step4.myadd.fa3.i1 ),
    .B(\step4.myadd.fa2.cout ),
    .Y(_409_)
);

NOR2X1 _1457_ (
    .A(\step4.myadd.fa3.i1 ),
    .B(\step4.myadd.fa2.cout ),
    .Y(_410_)
);

OAI21X1 _1458_ (
    .A(_410_),
    .B(_409_),
    .C(\step4.myadd.fa3.i0 ),
    .Y(_411_)
);

INVX1 _1459_ (
    .A(\step4.myadd.fa3.i0 ),
    .Y(_412_)
);

NAND2X1 _1460_ (
    .A(\step4.myadd.fa3.i1 ),
    .B(\step4.myadd.fa2.cout ),
    .Y(_406_)
);

OR2X2 _1461_ (
    .A(\step4.myadd.fa3.i1 ),
    .B(\step4.myadd.fa2.cout ),
    .Y(_407_)
);

NAND3X1 _1462_ (
    .A(_412_),
    .B(_406_),
    .C(_407_),
    .Y(_408_)
);

NAND2X1 _1463_ (
    .A(_411_),
    .B(_408_),
    .Y(\step4.myadd.fa3.sum )
);

AOI21X1 _1464_ (
    .A(_412_),
    .B(_406_),
    .C(_410_),
    .Y(\step4.myadd.fa3.cout )
);

AND2X2 _1465_ (
    .A(\step4.myadd.fa4.i1 ),
    .B(\step4.myadd.fa3.cout ),
    .Y(_416_)
);

NOR2X1 _1466_ (
    .A(\step4.myadd.fa4.i1 ),
    .B(\step4.myadd.fa3.cout ),
    .Y(_417_)
);

OAI21X1 _1467_ (
    .A(_417_),
    .B(_416_),
    .C(\step4.myadd.fa4.i0 ),
    .Y(_418_)
);

INVX1 _1468_ (
    .A(\step4.myadd.fa4.i0 ),
    .Y(_419_)
);

NAND2X1 _1469_ (
    .A(\step4.myadd.fa4.i1 ),
    .B(\step4.myadd.fa3.cout ),
    .Y(_413_)
);

OR2X2 _1470_ (
    .A(\step4.myadd.fa4.i1 ),
    .B(\step4.myadd.fa3.cout ),
    .Y(_414_)
);

NAND3X1 _1471_ (
    .A(_419_),
    .B(_413_),
    .C(_414_),
    .Y(_415_)
);

NAND2X1 _1472_ (
    .A(_418_),
    .B(_415_),
    .Y(\step4.myadd.fa4.sum )
);

AOI21X1 _1473_ (
    .A(_419_),
    .B(_413_),
    .C(_417_),
    .Y(\step4.myadd.fa4.cout )
);

AND2X2 _1474_ (
    .A(\step4.myadd.fa5.i1 ),
    .B(\step4.myadd.fa4.cout ),
    .Y(_423_)
);

NOR2X1 _1475_ (
    .A(\step4.myadd.fa5.i1 ),
    .B(\step4.myadd.fa4.cout ),
    .Y(_424_)
);

OAI21X1 _1476_ (
    .A(_424_),
    .B(_423_),
    .C(\step4.myadd.fa5.i0 ),
    .Y(_425_)
);

INVX1 _1477_ (
    .A(\step4.myadd.fa5.i0 ),
    .Y(_426_)
);

NAND2X1 _1478_ (
    .A(\step4.myadd.fa5.i1 ),
    .B(\step4.myadd.fa4.cout ),
    .Y(_420_)
);

OR2X2 _1479_ (
    .A(\step4.myadd.fa5.i1 ),
    .B(\step4.myadd.fa4.cout ),
    .Y(_421_)
);

NAND3X1 _1480_ (
    .A(_426_),
    .B(_420_),
    .C(_421_),
    .Y(_422_)
);

NAND2X1 _1481_ (
    .A(_425_),
    .B(_422_),
    .Y(\step4.myadd.fa5.sum )
);

AOI21X1 _1482_ (
    .A(_426_),
    .B(_420_),
    .C(_424_),
    .Y(\step4.myadd.fa5.cout )
);

AND2X2 _1483_ (
    .A(\step4.myadd.fa6.i1 ),
    .B(\step4.myadd.fa5.cout ),
    .Y(_430_)
);

NOR2X1 _1484_ (
    .A(\step4.myadd.fa6.i1 ),
    .B(\step4.myadd.fa5.cout ),
    .Y(_431_)
);

OAI21X1 _1485_ (
    .A(_431_),
    .B(_430_),
    .C(\step4.myadd.fa6.i0 ),
    .Y(_432_)
);

INVX1 _1486_ (
    .A(\step4.myadd.fa6.i0 ),
    .Y(_433_)
);

NAND2X1 _1487_ (
    .A(\step4.myadd.fa6.i1 ),
    .B(\step4.myadd.fa5.cout ),
    .Y(_427_)
);

OR2X2 _1488_ (
    .A(\step4.myadd.fa6.i1 ),
    .B(\step4.myadd.fa5.cout ),
    .Y(_428_)
);

NAND3X1 _1489_ (
    .A(_433_),
    .B(_427_),
    .C(_428_),
    .Y(_429_)
);

NAND2X1 _1490_ (
    .A(_432_),
    .B(_429_),
    .Y(\step4.myadd.fa6.sum )
);

AOI21X1 _1491_ (
    .A(_433_),
    .B(_427_),
    .C(_431_),
    .Y(\step4.myadd.fa6.cout )
);

AND2X2 _1492_ (
    .A(\step4.myadd.fa7.i1 ),
    .B(\step4.myadd.fa6.cout ),
    .Y(_437_)
);

NOR2X1 _1493_ (
    .A(\step4.myadd.fa7.i1 ),
    .B(\step4.myadd.fa6.cout ),
    .Y(_438_)
);

OAI21X1 _1494_ (
    .A(_438_),
    .B(_437_),
    .C(\step4.myadd.fa7.i0 ),
    .Y(_439_)
);

INVX1 _1495_ (
    .A(\step4.myadd.fa7.i0 ),
    .Y(_440_)
);

NAND2X1 _1496_ (
    .A(\step4.myadd.fa7.i1 ),
    .B(\step4.myadd.fa6.cout ),
    .Y(_434_)
);

OR2X2 _1497_ (
    .A(\step4.myadd.fa7.i1 ),
    .B(\step4.myadd.fa6.cout ),
    .Y(_435_)
);

NAND3X1 _1498_ (
    .A(_440_),
    .B(_434_),
    .C(_435_),
    .Y(_436_)
);

NAND2X1 _1499_ (
    .A(_439_),
    .B(_436_),
    .Y(\step4.myadd.fa7.sum )
);

AOI21X1 _1500_ (
    .A(_440_),
    .B(_434_),
    .C(_438_),
    .Y(\step4.myadd.fa7.cout )
);

AND2X2 _1501_ (
    .A(\step4.myadd.fa8.i1 ),
    .B(\step4.myadd.fa7.cout ),
    .Y(_444_)
);

NOR2X1 _1502_ (
    .A(\step4.myadd.fa8.i1 ),
    .B(\step4.myadd.fa7.cout ),
    .Y(_445_)
);

OAI21X1 _1503_ (
    .A(_445_),
    .B(_444_),
    .C(\step4.myadd.fa7.i0 ),
    .Y(_446_)
);

INVX1 _1504_ (
    .A(\step4.myadd.fa7.i0 ),
    .Y(_447_)
);

NAND2X1 _1505_ (
    .A(\step4.myadd.fa8.i1 ),
    .B(\step4.myadd.fa7.cout ),
    .Y(_441_)
);

OR2X2 _1506_ (
    .A(\step4.myadd.fa8.i1 ),
    .B(\step4.myadd.fa7.cout ),
    .Y(_442_)
);

NAND3X1 _1507_ (
    .A(_447_),
    .B(_441_),
    .C(_442_),
    .Y(_443_)
);

NAND2X1 _1508_ (
    .A(_446_),
    .B(_443_),
    .Y(\step4.myadd.fa8.sum )
);

INVX1 _1509_ (
    .A(\step4.myadd.cin_bF$buf1 ),
    .Y(_448_)
);

NAND2X1 _1510_ (
    .A(\step1.myadd.x0.i0_bF$buf1 ),
    .B(_448_),
    .Y(_449_)
);

INVX1 _1511_ (
    .A(\step1.myadd.x0.i0_bF$buf0 ),
    .Y(_450_)
);

NAND2X1 _1512_ (
    .A(\step4.myadd.cin_bF$buf0 ),
    .B(_450_),
    .Y(_451_)
);

NAND2X1 _1513_ (
    .A(_449_),
    .B(_451_),
    .Y(\step4.myadd.fa1.i1 )
);

INVX1 _1514_ (
    .A(\step4.myadd.cin_bF$buf4 ),
    .Y(_452_)
);

NAND2X1 _1515_ (
    .A(\step1.myadd.x1.i0_bF$buf1 ),
    .B(_452_),
    .Y(_453_)
);

INVX1 _1516_ (
    .A(\step1.myadd.x1.i0_bF$buf0 ),
    .Y(_454_)
);

NAND2X1 _1517_ (
    .A(\step4.myadd.cin_bF$buf3 ),
    .B(_454_),
    .Y(_455_)
);

NAND2X1 _1518_ (
    .A(_453_),
    .B(_455_),
    .Y(\step4.myadd.fa2.i1 )
);

INVX1 _1519_ (
    .A(\step4.myadd.cin_bF$buf2 ),
    .Y(_456_)
);

NAND2X1 _1520_ (
    .A(\step1.myadd.x2.i0_bF$buf1 ),
    .B(_456_),
    .Y(_457_)
);

INVX1 _1521_ (
    .A(\step1.myadd.x2.i0_bF$buf0 ),
    .Y(_458_)
);

NAND2X1 _1522_ (
    .A(\step4.myadd.cin_bF$buf1 ),
    .B(_458_),
    .Y(_459_)
);

NAND2X1 _1523_ (
    .A(_457_),
    .B(_459_),
    .Y(\step4.myadd.fa3.i1 )
);

INVX1 _1524_ (
    .A(\step4.myadd.cin_bF$buf0 ),
    .Y(_460_)
);

NAND2X1 _1525_ (
    .A(\step1.myadd.x3.i0_bF$buf1 ),
    .B(_460_),
    .Y(_461_)
);

INVX1 _1526_ (
    .A(\step1.myadd.x3.i0_bF$buf0 ),
    .Y(_462_)
);

NAND2X1 _1527_ (
    .A(\step4.myadd.cin_bF$buf4 ),
    .B(_462_),
    .Y(_463_)
);

NAND2X1 _1528_ (
    .A(_461_),
    .B(_463_),
    .Y(\step4.myadd.fa4.i1 )
);

INVX1 _1529_ (
    .A(\step4.myadd.cin_bF$buf3 ),
    .Y(_464_)
);

NAND2X1 _1530_ (
    .A(\step1.myadd.x4.i0_bF$buf1 ),
    .B(_464_),
    .Y(_465_)
);

INVX1 _1531_ (
    .A(\step1.myadd.x4.i0_bF$buf0 ),
    .Y(_466_)
);

NAND2X1 _1532_ (
    .A(\step4.myadd.cin_bF$buf2 ),
    .B(_466_),
    .Y(_467_)
);

NAND2X1 _1533_ (
    .A(_465_),
    .B(_467_),
    .Y(\step4.myadd.fa5.i1 )
);

INVX1 _1534_ (
    .A(\step4.myadd.cin_bF$buf1 ),
    .Y(_468_)
);

NAND2X1 _1535_ (
    .A(\step1.myadd.x5.i0_bF$buf1 ),
    .B(_468_),
    .Y(_469_)
);

INVX1 _1536_ (
    .A(\step1.myadd.x5.i0_bF$buf0 ),
    .Y(_470_)
);

NAND2X1 _1537_ (
    .A(\step4.myadd.cin_bF$buf0 ),
    .B(_470_),
    .Y(_471_)
);

NAND2X1 _1538_ (
    .A(_469_),
    .B(_471_),
    .Y(\step4.myadd.fa6.i1 )
);

INVX1 _1539_ (
    .A(\step4.myadd.cin_bF$buf4 ),
    .Y(_472_)
);

NAND2X1 _1540_ (
    .A(\step1.myadd.x6.i0_bF$buf1 ),
    .B(_472_),
    .Y(_473_)
);

INVX1 _1541_ (
    .A(\step1.myadd.x6.i0_bF$buf0 ),
    .Y(_474_)
);

NAND2X1 _1542_ (
    .A(\step4.myadd.cin_bF$buf3 ),
    .B(_474_),
    .Y(_475_)
);

NAND2X1 _1543_ (
    .A(_473_),
    .B(_475_),
    .Y(\step4.myadd.fa7.i1 )
);

INVX1 _1544_ (
    .A(\step4.myadd.cin_bF$buf2 ),
    .Y(_476_)
);

NAND2X1 _1545_ (
    .A(\step1.myadd.x7.i0_bF$buf1 ),
    .B(_476_),
    .Y(_477_)
);

INVX1 _1546_ (
    .A(\step1.myadd.x7.i0_bF$buf0 ),
    .Y(_478_)
);

NAND2X1 _1547_ (
    .A(\step4.myadd.cin_bF$buf1 ),
    .B(_478_),
    .Y(_479_)
);

NAND2X1 _1548_ (
    .A(_477_),
    .B(_479_),
    .Y(\step4.myadd.fa8.i1 )
);

OR2X2 _1549_ (
    .A(\step4.myadd.cin_bF$buf0 ),
    .B(\step5.myadd.cin_bF$buf4 ),
    .Y(_480_)
);

NAND2X1 _1550_ (
    .A(\step4.myadd.cin_bF$buf4 ),
    .B(\step5.myadd.cin_bF$buf3 ),
    .Y(_481_)
);

NAND3X1 _1551_ (
    .A(\step5.myadd.fa2.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_482_)
);

NOR2X1 _1552_ (
    .A(\step4.myadd.cin_bF$buf3 ),
    .B(\step5.myadd.cin_bF$buf2 ),
    .Y(_483_)
);

AND2X2 _1553_ (
    .A(\step4.myadd.cin_bF$buf2 ),
    .B(\step5.myadd.cin_bF$buf1 ),
    .Y(_484_)
);

OAI21X1 _1554_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa2.i0 ),
    .Y(_485_)
);

NAND2X1 _1555_ (
    .A(_485_),
    .B(_482_),
    .Y(\step6.myadd.fa1.i0 )
);

NAND3X1 _1556_ (
    .A(\step5.myadd.fa3.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_486_)
);

OAI21X1 _1557_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa3.i0 ),
    .Y(_487_)
);

NAND2X1 _1558_ (
    .A(_487_),
    .B(_486_),
    .Y(\step6.myadd.fa2.i0 )
);

NAND3X1 _1559_ (
    .A(\step5.myadd.fa4.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_488_)
);

OAI21X1 _1560_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa4.i0 ),
    .Y(_489_)
);

NAND2X1 _1561_ (
    .A(_489_),
    .B(_488_),
    .Y(\step6.myadd.fa3.i0 )
);

NAND3X1 _1562_ (
    .A(\step5.myadd.fa5.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_490_)
);

OAI21X1 _1563_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa5.i0 ),
    .Y(_491_)
);

NAND2X1 _1564_ (
    .A(_491_),
    .B(_490_),
    .Y(\step6.myadd.fa4.i0 )
);

NAND3X1 _1565_ (
    .A(\step5.myadd.fa6.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_492_)
);

OAI21X1 _1566_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa6.i0 ),
    .Y(_493_)
);

NAND2X1 _1567_ (
    .A(_493_),
    .B(_492_),
    .Y(\step6.myadd.fa5.i0 )
);

NAND3X1 _1568_ (
    .A(\step5.myadd.fa7.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_494_)
);

OAI21X1 _1569_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa7.i0 ),
    .Y(_495_)
);

NAND2X1 _1570_ (
    .A(_495_),
    .B(_494_),
    .Y(\step6.myadd.fa6.i0 )
);

NAND3X1 _1571_ (
    .A(\step5.myadd.fa8.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_496_)
);

OAI21X1 _1572_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa7.i0 ),
    .Y(_497_)
);

NAND2X1 _1573_ (
    .A(_497_),
    .B(_496_),
    .Y(\step6.myadd.fa7.i0 )
);

NAND3X1 _1574_ (
    .A(\step5.myadd.fa1.sum ),
    .B(_481_),
    .C(_480_),
    .Y(_498_)
);

OAI21X1 _1575_ (
    .A(_483_),
    .B(_484_),
    .C(\step5.myadd.fa1.i0 ),
    .Y(_499_)
);

NAND2X1 _1576_ (
    .A(_499_),
    .B(_498_),
    .Y(\Q[4] [7])
);

AND2X2 _1577_ (
    .A(\step5.myadd.fa1.i1 ),
    .B(\step5.myadd.cin_bF$buf0 ),
    .Y(_503_)
);

NOR2X1 _1578_ (
    .A(\step5.myadd.fa1.i1 ),
    .B(\step5.myadd.cin_bF$buf4 ),
    .Y(_504_)
);

OAI21X1 _1579_ (
    .A(_504_),
    .B(_503_),
    .C(\step5.myadd.fa1.i0 ),
    .Y(_505_)
);

INVX1 _1580_ (
    .A(\step5.myadd.fa1.i0 ),
    .Y(_506_)
);

NAND2X1 _1581_ (
    .A(\step5.myadd.fa1.i1 ),
    .B(\step5.myadd.cin_bF$buf3 ),
    .Y(_500_)
);

OR2X2 _1582_ (
    .A(\step5.myadd.fa1.i1 ),
    .B(\step5.myadd.cin_bF$buf2 ),
    .Y(_501_)
);

NAND3X1 _1583_ (
    .A(_506_),
    .B(_500_),
    .C(_501_),
    .Y(_502_)
);

NAND2X1 _1584_ (
    .A(_505_),
    .B(_502_),
    .Y(\step5.myadd.fa1.sum )
);

AOI21X1 _1585_ (
    .A(_506_),
    .B(_500_),
    .C(_504_),
    .Y(\step5.myadd.fa1.cout )
);

AND2X2 _1586_ (
    .A(\step5.myadd.fa2.i1 ),
    .B(\step5.myadd.fa1.cout ),
    .Y(_510_)
);

NOR2X1 _1587_ (
    .A(\step5.myadd.fa2.i1 ),
    .B(\step5.myadd.fa1.cout ),
    .Y(_511_)
);

OAI21X1 _1588_ (
    .A(_511_),
    .B(_510_),
    .C(\step5.myadd.fa2.i0 ),
    .Y(_512_)
);

INVX1 _1589_ (
    .A(\step5.myadd.fa2.i0 ),
    .Y(_513_)
);

NAND2X1 _1590_ (
    .A(\step5.myadd.fa2.i1 ),
    .B(\step5.myadd.fa1.cout ),
    .Y(_507_)
);

OR2X2 _1591_ (
    .A(\step5.myadd.fa2.i1 ),
    .B(\step5.myadd.fa1.cout ),
    .Y(_508_)
);

NAND3X1 _1592_ (
    .A(_513_),
    .B(_507_),
    .C(_508_),
    .Y(_509_)
);

NAND2X1 _1593_ (
    .A(_512_),
    .B(_509_),
    .Y(\step5.myadd.fa2.sum )
);

AOI21X1 _1594_ (
    .A(_513_),
    .B(_507_),
    .C(_511_),
    .Y(\step5.myadd.fa2.cout )
);

AND2X2 _1595_ (
    .A(\step5.myadd.fa3.i1 ),
    .B(\step5.myadd.fa2.cout ),
    .Y(_517_)
);

NOR2X1 _1596_ (
    .A(\step5.myadd.fa3.i1 ),
    .B(\step5.myadd.fa2.cout ),
    .Y(_518_)
);

OAI21X1 _1597_ (
    .A(_518_),
    .B(_517_),
    .C(\step5.myadd.fa3.i0 ),
    .Y(_519_)
);

INVX1 _1598_ (
    .A(\step5.myadd.fa3.i0 ),
    .Y(_520_)
);

NAND2X1 _1599_ (
    .A(\step5.myadd.fa3.i1 ),
    .B(\step5.myadd.fa2.cout ),
    .Y(_514_)
);

OR2X2 _1600_ (
    .A(\step5.myadd.fa3.i1 ),
    .B(\step5.myadd.fa2.cout ),
    .Y(_515_)
);

NAND3X1 _1601_ (
    .A(_520_),
    .B(_514_),
    .C(_515_),
    .Y(_516_)
);

NAND2X1 _1602_ (
    .A(_519_),
    .B(_516_),
    .Y(\step5.myadd.fa3.sum )
);

AOI21X1 _1603_ (
    .A(_520_),
    .B(_514_),
    .C(_518_),
    .Y(\step5.myadd.fa3.cout )
);

AND2X2 _1604_ (
    .A(\step5.myadd.fa4.i1 ),
    .B(\step5.myadd.fa3.cout ),
    .Y(_524_)
);

NOR2X1 _1605_ (
    .A(\step5.myadd.fa4.i1 ),
    .B(\step5.myadd.fa3.cout ),
    .Y(_525_)
);

OAI21X1 _1606_ (
    .A(_525_),
    .B(_524_),
    .C(\step5.myadd.fa4.i0 ),
    .Y(_526_)
);

INVX1 _1607_ (
    .A(\step5.myadd.fa4.i0 ),
    .Y(_527_)
);

NAND2X1 _1608_ (
    .A(\step5.myadd.fa4.i1 ),
    .B(\step5.myadd.fa3.cout ),
    .Y(_521_)
);

OR2X2 _1609_ (
    .A(\step5.myadd.fa4.i1 ),
    .B(\step5.myadd.fa3.cout ),
    .Y(_522_)
);

NAND3X1 _1610_ (
    .A(_527_),
    .B(_521_),
    .C(_522_),
    .Y(_523_)
);

NAND2X1 _1611_ (
    .A(_526_),
    .B(_523_),
    .Y(\step5.myadd.fa4.sum )
);

AOI21X1 _1612_ (
    .A(_527_),
    .B(_521_),
    .C(_525_),
    .Y(\step5.myadd.fa4.cout )
);

AND2X2 _1613_ (
    .A(\step5.myadd.fa5.i1 ),
    .B(\step5.myadd.fa4.cout ),
    .Y(_531_)
);

NOR2X1 _1614_ (
    .A(\step5.myadd.fa5.i1 ),
    .B(\step5.myadd.fa4.cout ),
    .Y(_532_)
);

OAI21X1 _1615_ (
    .A(_532_),
    .B(_531_),
    .C(\step5.myadd.fa5.i0 ),
    .Y(_533_)
);

INVX1 _1616_ (
    .A(\step5.myadd.fa5.i0 ),
    .Y(_534_)
);

NAND2X1 _1617_ (
    .A(\step5.myadd.fa5.i1 ),
    .B(\step5.myadd.fa4.cout ),
    .Y(_528_)
);

OR2X2 _1618_ (
    .A(\step5.myadd.fa5.i1 ),
    .B(\step5.myadd.fa4.cout ),
    .Y(_529_)
);

NAND3X1 _1619_ (
    .A(_534_),
    .B(_528_),
    .C(_529_),
    .Y(_530_)
);

NAND2X1 _1620_ (
    .A(_533_),
    .B(_530_),
    .Y(\step5.myadd.fa5.sum )
);

AOI21X1 _1621_ (
    .A(_534_),
    .B(_528_),
    .C(_532_),
    .Y(\step5.myadd.fa5.cout )
);

AND2X2 _1622_ (
    .A(\step5.myadd.fa6.i1 ),
    .B(\step5.myadd.fa5.cout ),
    .Y(_538_)
);

NOR2X1 _1623_ (
    .A(\step5.myadd.fa6.i1 ),
    .B(\step5.myadd.fa5.cout ),
    .Y(_539_)
);

OAI21X1 _1624_ (
    .A(_539_),
    .B(_538_),
    .C(\step5.myadd.fa6.i0 ),
    .Y(_540_)
);

INVX1 _1625_ (
    .A(\step5.myadd.fa6.i0 ),
    .Y(_541_)
);

NAND2X1 _1626_ (
    .A(\step5.myadd.fa6.i1 ),
    .B(\step5.myadd.fa5.cout ),
    .Y(_535_)
);

OR2X2 _1627_ (
    .A(\step5.myadd.fa6.i1 ),
    .B(\step5.myadd.fa5.cout ),
    .Y(_536_)
);

NAND3X1 _1628_ (
    .A(_541_),
    .B(_535_),
    .C(_536_),
    .Y(_537_)
);

NAND2X1 _1629_ (
    .A(_540_),
    .B(_537_),
    .Y(\step5.myadd.fa6.sum )
);

AOI21X1 _1630_ (
    .A(_541_),
    .B(_535_),
    .C(_539_),
    .Y(\step5.myadd.fa6.cout )
);

AND2X2 _1631_ (
    .A(\step5.myadd.fa7.i1 ),
    .B(\step5.myadd.fa6.cout ),
    .Y(_545_)
);

NOR2X1 _1632_ (
    .A(\step5.myadd.fa7.i1 ),
    .B(\step5.myadd.fa6.cout ),
    .Y(_546_)
);

OAI21X1 _1633_ (
    .A(_546_),
    .B(_545_),
    .C(\step5.myadd.fa7.i0 ),
    .Y(_547_)
);

INVX1 _1634_ (
    .A(\step5.myadd.fa7.i0 ),
    .Y(_548_)
);

NAND2X1 _1635_ (
    .A(\step5.myadd.fa7.i1 ),
    .B(\step5.myadd.fa6.cout ),
    .Y(_542_)
);

OR2X2 _1636_ (
    .A(\step5.myadd.fa7.i1 ),
    .B(\step5.myadd.fa6.cout ),
    .Y(_543_)
);

NAND3X1 _1637_ (
    .A(_548_),
    .B(_542_),
    .C(_543_),
    .Y(_544_)
);

NAND2X1 _1638_ (
    .A(_547_),
    .B(_544_),
    .Y(\step5.myadd.fa7.sum )
);

AOI21X1 _1639_ (
    .A(_548_),
    .B(_542_),
    .C(_546_),
    .Y(\step5.myadd.fa7.cout )
);

AND2X2 _1640_ (
    .A(\step5.myadd.fa8.i1 ),
    .B(\step5.myadd.fa7.cout ),
    .Y(_552_)
);

NOR2X1 _1641_ (
    .A(\step5.myadd.fa8.i1 ),
    .B(\step5.myadd.fa7.cout ),
    .Y(_553_)
);

OAI21X1 _1642_ (
    .A(_553_),
    .B(_552_),
    .C(\step5.myadd.fa7.i0 ),
    .Y(_554_)
);

INVX1 _1643_ (
    .A(\step5.myadd.fa7.i0 ),
    .Y(_555_)
);

NAND2X1 _1644_ (
    .A(\step5.myadd.fa8.i1 ),
    .B(\step5.myadd.fa7.cout ),
    .Y(_549_)
);

OR2X2 _1645_ (
    .A(\step5.myadd.fa8.i1 ),
    .B(\step5.myadd.fa7.cout ),
    .Y(_550_)
);

NAND3X1 _1646_ (
    .A(_555_),
    .B(_549_),
    .C(_550_),
    .Y(_551_)
);

NAND2X1 _1647_ (
    .A(_554_),
    .B(_551_),
    .Y(\step5.myadd.fa8.sum )
);

INVX1 _1648_ (
    .A(\step5.myadd.cin_bF$buf1 ),
    .Y(_556_)
);

NAND2X1 _1649_ (
    .A(\step1.myadd.x0.i0_bF$buf3 ),
    .B(_556_),
    .Y(_557_)
);

INVX1 _1650_ (
    .A(\step1.myadd.x0.i0_bF$buf2 ),
    .Y(_558_)
);

NAND2X1 _1651_ (
    .A(\step5.myadd.cin_bF$buf0 ),
    .B(_558_),
    .Y(_559_)
);

NAND2X1 _1652_ (
    .A(_557_),
    .B(_559_),
    .Y(\step5.myadd.fa1.i1 )
);

INVX1 _1653_ (
    .A(\step5.myadd.cin_bF$buf4 ),
    .Y(_560_)
);

NAND2X1 _1654_ (
    .A(\step1.myadd.x1.i0_bF$buf3 ),
    .B(_560_),
    .Y(_561_)
);

INVX1 _1655_ (
    .A(\step1.myadd.x1.i0_bF$buf2 ),
    .Y(_562_)
);

NAND2X1 _1656_ (
    .A(\step5.myadd.cin_bF$buf3 ),
    .B(_562_),
    .Y(_563_)
);

NAND2X1 _1657_ (
    .A(_561_),
    .B(_563_),
    .Y(\step5.myadd.fa2.i1 )
);

INVX1 _1658_ (
    .A(\step5.myadd.cin_bF$buf2 ),
    .Y(_564_)
);

NAND2X1 _1659_ (
    .A(\step1.myadd.x2.i0_bF$buf3 ),
    .B(_564_),
    .Y(_565_)
);

INVX1 _1660_ (
    .A(\step1.myadd.x2.i0_bF$buf2 ),
    .Y(_566_)
);

NAND2X1 _1661_ (
    .A(\step5.myadd.cin_bF$buf1 ),
    .B(_566_),
    .Y(_567_)
);

NAND2X1 _1662_ (
    .A(_565_),
    .B(_567_),
    .Y(\step5.myadd.fa3.i1 )
);

INVX1 _1663_ (
    .A(\step5.myadd.cin_bF$buf0 ),
    .Y(_568_)
);

NAND2X1 _1664_ (
    .A(\step1.myadd.x3.i0_bF$buf3 ),
    .B(_568_),
    .Y(_569_)
);

INVX1 _1665_ (
    .A(\step1.myadd.x3.i0_bF$buf2 ),
    .Y(_570_)
);

NAND2X1 _1666_ (
    .A(\step5.myadd.cin_bF$buf4 ),
    .B(_570_),
    .Y(_571_)
);

NAND2X1 _1667_ (
    .A(_569_),
    .B(_571_),
    .Y(\step5.myadd.fa4.i1 )
);

INVX1 _1668_ (
    .A(\step5.myadd.cin_bF$buf3 ),
    .Y(_572_)
);

NAND2X1 _1669_ (
    .A(\step1.myadd.x4.i0_bF$buf3 ),
    .B(_572_),
    .Y(_573_)
);

INVX1 _1670_ (
    .A(\step1.myadd.x4.i0_bF$buf2 ),
    .Y(_574_)
);

NAND2X1 _1671_ (
    .A(\step5.myadd.cin_bF$buf2 ),
    .B(_574_),
    .Y(_575_)
);

NAND2X1 _1672_ (
    .A(_573_),
    .B(_575_),
    .Y(\step5.myadd.fa5.i1 )
);

INVX1 _1673_ (
    .A(\step5.myadd.cin_bF$buf1 ),
    .Y(_576_)
);

NAND2X1 _1674_ (
    .A(\step1.myadd.x5.i0_bF$buf3 ),
    .B(_576_),
    .Y(_577_)
);

INVX1 _1675_ (
    .A(\step1.myadd.x5.i0_bF$buf2 ),
    .Y(_578_)
);

NAND2X1 _1676_ (
    .A(\step5.myadd.cin_bF$buf0 ),
    .B(_578_),
    .Y(_579_)
);

NAND2X1 _1677_ (
    .A(_577_),
    .B(_579_),
    .Y(\step5.myadd.fa6.i1 )
);

INVX1 _1678_ (
    .A(\step5.myadd.cin_bF$buf4 ),
    .Y(_580_)
);

NAND2X1 _1679_ (
    .A(\step1.myadd.x6.i0_bF$buf3 ),
    .B(_580_),
    .Y(_581_)
);

INVX1 _1680_ (
    .A(\step1.myadd.x6.i0_bF$buf2 ),
    .Y(_582_)
);

NAND2X1 _1681_ (
    .A(\step5.myadd.cin_bF$buf3 ),
    .B(_582_),
    .Y(_583_)
);

NAND2X1 _1682_ (
    .A(_581_),
    .B(_583_),
    .Y(\step5.myadd.fa7.i1 )
);

INVX1 _1683_ (
    .A(\step5.myadd.cin_bF$buf2 ),
    .Y(_584_)
);

NAND2X1 _1684_ (
    .A(\step1.myadd.x7.i0_bF$buf3 ),
    .B(_584_),
    .Y(_585_)
);

INVX1 _1685_ (
    .A(\step1.myadd.x7.i0_bF$buf2 ),
    .Y(_586_)
);

NAND2X1 _1686_ (
    .A(\step5.myadd.cin_bF$buf1 ),
    .B(_586_),
    .Y(_587_)
);

NAND2X1 _1687_ (
    .A(_585_),
    .B(_587_),
    .Y(\step5.myadd.fa8.i1 )
);

OR2X2 _1688_ (
    .A(\step5.myadd.cin_bF$buf0 ),
    .B(\step6.myadd.cin_bF$buf4 ),
    .Y(_588_)
);

NAND2X1 _1689_ (
    .A(\step5.myadd.cin_bF$buf4 ),
    .B(\step6.myadd.cin_bF$buf3 ),
    .Y(_589_)
);

NAND3X1 _1690_ (
    .A(\step6.myadd.fa2.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_590_)
);

NOR2X1 _1691_ (
    .A(\step5.myadd.cin_bF$buf3 ),
    .B(\step6.myadd.cin_bF$buf2 ),
    .Y(_591_)
);

AND2X2 _1692_ (
    .A(\step5.myadd.cin_bF$buf2 ),
    .B(\step6.myadd.cin_bF$buf1 ),
    .Y(_592_)
);

OAI21X1 _1693_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa2.i0 ),
    .Y(_593_)
);

NAND2X1 _1694_ (
    .A(_593_),
    .B(_590_),
    .Y(\step7.myadd.fa1.i0 )
);

NAND3X1 _1695_ (
    .A(\step6.myadd.fa3.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_594_)
);

OAI21X1 _1696_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa3.i0 ),
    .Y(_595_)
);

NAND2X1 _1697_ (
    .A(_595_),
    .B(_594_),
    .Y(\step7.myadd.fa2.i0 )
);

NAND3X1 _1698_ (
    .A(\step6.myadd.fa4.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_596_)
);

OAI21X1 _1699_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa4.i0 ),
    .Y(_597_)
);

NAND2X1 _1700_ (
    .A(_597_),
    .B(_596_),
    .Y(\step7.myadd.fa3.i0 )
);

NAND3X1 _1701_ (
    .A(\step6.myadd.fa5.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_598_)
);

OAI21X1 _1702_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa5.i0 ),
    .Y(_599_)
);

NAND2X1 _1703_ (
    .A(_599_),
    .B(_598_),
    .Y(\step7.myadd.fa4.i0 )
);

NAND3X1 _1704_ (
    .A(\step6.myadd.fa6.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_600_)
);

OAI21X1 _1705_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa6.i0 ),
    .Y(_601_)
);

NAND2X1 _1706_ (
    .A(_601_),
    .B(_600_),
    .Y(\step7.myadd.fa5.i0 )
);

NAND3X1 _1707_ (
    .A(\step6.myadd.fa7.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_602_)
);

OAI21X1 _1708_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa7.i0 ),
    .Y(_603_)
);

NAND2X1 _1709_ (
    .A(_603_),
    .B(_602_),
    .Y(\step7.myadd.fa6.i0 )
);

NAND3X1 _1710_ (
    .A(\step6.myadd.fa8.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_604_)
);

OAI21X1 _1711_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa7.i0 ),
    .Y(_605_)
);

NAND2X1 _1712_ (
    .A(_605_),
    .B(_604_),
    .Y(\step7.myadd.fa7.i0 )
);

NAND3X1 _1713_ (
    .A(\step6.myadd.fa1.sum ),
    .B(_589_),
    .C(_588_),
    .Y(_606_)
);

OAI21X1 _1714_ (
    .A(_591_),
    .B(_592_),
    .C(\step6.myadd.fa1.i0 ),
    .Y(_607_)
);

NAND2X1 _1715_ (
    .A(_607_),
    .B(_606_),
    .Y(\Q[5] [7])
);

AND2X2 _1716_ (
    .A(\step6.myadd.fa1.i1 ),
    .B(\step6.myadd.cin_bF$buf0 ),
    .Y(_611_)
);

NOR2X1 _1717_ (
    .A(\step6.myadd.fa1.i1 ),
    .B(\step6.myadd.cin_bF$buf4 ),
    .Y(_612_)
);

OAI21X1 _1718_ (
    .A(_612_),
    .B(_611_),
    .C(\step6.myadd.fa1.i0 ),
    .Y(_613_)
);

INVX1 _1719_ (
    .A(\step6.myadd.fa1.i0 ),
    .Y(_614_)
);

NAND2X1 _1720_ (
    .A(\step6.myadd.fa1.i1 ),
    .B(\step6.myadd.cin_bF$buf3 ),
    .Y(_608_)
);

OR2X2 _1721_ (
    .A(\step6.myadd.fa1.i1 ),
    .B(\step6.myadd.cin_bF$buf2 ),
    .Y(_609_)
);

NAND3X1 _1722_ (
    .A(_614_),
    .B(_608_),
    .C(_609_),
    .Y(_610_)
);

NAND2X1 _1723_ (
    .A(_613_),
    .B(_610_),
    .Y(\step6.myadd.fa1.sum )
);

AOI21X1 _1724_ (
    .A(_614_),
    .B(_608_),
    .C(_612_),
    .Y(\step6.myadd.fa1.cout )
);

AND2X2 _1725_ (
    .A(\step6.myadd.fa2.i1 ),
    .B(\step6.myadd.fa1.cout ),
    .Y(_618_)
);

NOR2X1 _1726_ (
    .A(\step6.myadd.fa2.i1 ),
    .B(\step6.myadd.fa1.cout ),
    .Y(_619_)
);

OAI21X1 _1727_ (
    .A(_619_),
    .B(_618_),
    .C(\step6.myadd.fa2.i0 ),
    .Y(_620_)
);

INVX1 _1728_ (
    .A(\step6.myadd.fa2.i0 ),
    .Y(_621_)
);

NAND2X1 _1729_ (
    .A(\step6.myadd.fa2.i1 ),
    .B(\step6.myadd.fa1.cout ),
    .Y(_615_)
);

OR2X2 _1730_ (
    .A(\step6.myadd.fa2.i1 ),
    .B(\step6.myadd.fa1.cout ),
    .Y(_616_)
);

NAND3X1 _1731_ (
    .A(_621_),
    .B(_615_),
    .C(_616_),
    .Y(_617_)
);

NAND2X1 _1732_ (
    .A(_620_),
    .B(_617_),
    .Y(\step6.myadd.fa2.sum )
);

AOI21X1 _1733_ (
    .A(_621_),
    .B(_615_),
    .C(_619_),
    .Y(\step6.myadd.fa2.cout )
);

AND2X2 _1734_ (
    .A(\step6.myadd.fa3.i1 ),
    .B(\step6.myadd.fa2.cout ),
    .Y(_625_)
);

NOR2X1 _1735_ (
    .A(\step6.myadd.fa3.i1 ),
    .B(\step6.myadd.fa2.cout ),
    .Y(_626_)
);

OAI21X1 _1736_ (
    .A(_626_),
    .B(_625_),
    .C(\step6.myadd.fa3.i0 ),
    .Y(_627_)
);

INVX1 _1737_ (
    .A(\step6.myadd.fa3.i0 ),
    .Y(_628_)
);

NAND2X1 _1738_ (
    .A(\step6.myadd.fa3.i1 ),
    .B(\step6.myadd.fa2.cout ),
    .Y(_622_)
);

OR2X2 _1739_ (
    .A(\step6.myadd.fa3.i1 ),
    .B(\step6.myadd.fa2.cout ),
    .Y(_623_)
);

NAND3X1 _1740_ (
    .A(_628_),
    .B(_622_),
    .C(_623_),
    .Y(_624_)
);

NAND2X1 _1741_ (
    .A(_627_),
    .B(_624_),
    .Y(\step6.myadd.fa3.sum )
);

AOI21X1 _1742_ (
    .A(_628_),
    .B(_622_),
    .C(_626_),
    .Y(\step6.myadd.fa3.cout )
);

AND2X2 _1743_ (
    .A(\step6.myadd.fa4.i1 ),
    .B(\step6.myadd.fa3.cout ),
    .Y(_632_)
);

NOR2X1 _1744_ (
    .A(\step6.myadd.fa4.i1 ),
    .B(\step6.myadd.fa3.cout ),
    .Y(_633_)
);

OAI21X1 _1745_ (
    .A(_633_),
    .B(_632_),
    .C(\step6.myadd.fa4.i0 ),
    .Y(_634_)
);

INVX1 _1746_ (
    .A(\step6.myadd.fa4.i0 ),
    .Y(_635_)
);

NAND2X1 _1747_ (
    .A(\step6.myadd.fa4.i1 ),
    .B(\step6.myadd.fa3.cout ),
    .Y(_629_)
);

OR2X2 _1748_ (
    .A(\step6.myadd.fa4.i1 ),
    .B(\step6.myadd.fa3.cout ),
    .Y(_630_)
);

NAND3X1 _1749_ (
    .A(_635_),
    .B(_629_),
    .C(_630_),
    .Y(_631_)
);

NAND2X1 _1750_ (
    .A(_634_),
    .B(_631_),
    .Y(\step6.myadd.fa4.sum )
);

AOI21X1 _1751_ (
    .A(_635_),
    .B(_629_),
    .C(_633_),
    .Y(\step6.myadd.fa4.cout )
);

AND2X2 _1752_ (
    .A(\step6.myadd.fa5.i1 ),
    .B(\step6.myadd.fa4.cout ),
    .Y(_639_)
);

NOR2X1 _1753_ (
    .A(\step6.myadd.fa5.i1 ),
    .B(\step6.myadd.fa4.cout ),
    .Y(_640_)
);

OAI21X1 _1754_ (
    .A(_640_),
    .B(_639_),
    .C(\step6.myadd.fa5.i0 ),
    .Y(_641_)
);

INVX1 _1755_ (
    .A(\step6.myadd.fa5.i0 ),
    .Y(_642_)
);

NAND2X1 _1756_ (
    .A(\step6.myadd.fa5.i1 ),
    .B(\step6.myadd.fa4.cout ),
    .Y(_636_)
);

OR2X2 _1757_ (
    .A(\step6.myadd.fa5.i1 ),
    .B(\step6.myadd.fa4.cout ),
    .Y(_637_)
);

NAND3X1 _1758_ (
    .A(_642_),
    .B(_636_),
    .C(_637_),
    .Y(_638_)
);

NAND2X1 _1759_ (
    .A(_641_),
    .B(_638_),
    .Y(\step6.myadd.fa5.sum )
);

AOI21X1 _1760_ (
    .A(_642_),
    .B(_636_),
    .C(_640_),
    .Y(\step6.myadd.fa5.cout )
);

AND2X2 _1761_ (
    .A(\step6.myadd.fa6.i1 ),
    .B(\step6.myadd.fa5.cout ),
    .Y(_646_)
);

NOR2X1 _1762_ (
    .A(\step6.myadd.fa6.i1 ),
    .B(\step6.myadd.fa5.cout ),
    .Y(_647_)
);

OAI21X1 _1763_ (
    .A(_647_),
    .B(_646_),
    .C(\step6.myadd.fa6.i0 ),
    .Y(_648_)
);

INVX1 _1764_ (
    .A(\step6.myadd.fa6.i0 ),
    .Y(_649_)
);

NAND2X1 _1765_ (
    .A(\step6.myadd.fa6.i1 ),
    .B(\step6.myadd.fa5.cout ),
    .Y(_643_)
);

OR2X2 _1766_ (
    .A(\step6.myadd.fa6.i1 ),
    .B(\step6.myadd.fa5.cout ),
    .Y(_644_)
);

NAND3X1 _1767_ (
    .A(_649_),
    .B(_643_),
    .C(_644_),
    .Y(_645_)
);

NAND2X1 _1768_ (
    .A(_648_),
    .B(_645_),
    .Y(\step6.myadd.fa6.sum )
);

AOI21X1 _1769_ (
    .A(_649_),
    .B(_643_),
    .C(_647_),
    .Y(\step6.myadd.fa6.cout )
);

AND2X2 _1770_ (
    .A(\step6.myadd.fa7.i1 ),
    .B(\step6.myadd.fa6.cout ),
    .Y(_653_)
);

NOR2X1 _1771_ (
    .A(\step6.myadd.fa7.i1 ),
    .B(\step6.myadd.fa6.cout ),
    .Y(_654_)
);

OAI21X1 _1772_ (
    .A(_654_),
    .B(_653_),
    .C(\step6.myadd.fa7.i0 ),
    .Y(_655_)
);

INVX1 _1773_ (
    .A(\step6.myadd.fa7.i0 ),
    .Y(_656_)
);

NAND2X1 _1774_ (
    .A(\step6.myadd.fa7.i1 ),
    .B(\step6.myadd.fa6.cout ),
    .Y(_650_)
);

OR2X2 _1775_ (
    .A(\step6.myadd.fa7.i1 ),
    .B(\step6.myadd.fa6.cout ),
    .Y(_651_)
);

NAND3X1 _1776_ (
    .A(_656_),
    .B(_650_),
    .C(_651_),
    .Y(_652_)
);

NAND2X1 _1777_ (
    .A(_655_),
    .B(_652_),
    .Y(\step6.myadd.fa7.sum )
);

AOI21X1 _1778_ (
    .A(_656_),
    .B(_650_),
    .C(_654_),
    .Y(\step6.myadd.fa7.cout )
);

AND2X2 _1779_ (
    .A(\step6.myadd.fa8.i1 ),
    .B(\step6.myadd.fa7.cout ),
    .Y(_660_)
);

NOR2X1 _1780_ (
    .A(\step6.myadd.fa8.i1 ),
    .B(\step6.myadd.fa7.cout ),
    .Y(_661_)
);

OAI21X1 _1781_ (
    .A(_661_),
    .B(_660_),
    .C(\step6.myadd.fa7.i0 ),
    .Y(_662_)
);

INVX1 _1782_ (
    .A(\step6.myadd.fa7.i0 ),
    .Y(_663_)
);

NAND2X1 _1783_ (
    .A(\step6.myadd.fa8.i1 ),
    .B(\step6.myadd.fa7.cout ),
    .Y(_657_)
);

OR2X2 _1784_ (
    .A(\step6.myadd.fa8.i1 ),
    .B(\step6.myadd.fa7.cout ),
    .Y(_658_)
);

NAND3X1 _1785_ (
    .A(_663_),
    .B(_657_),
    .C(_658_),
    .Y(_659_)
);

NAND2X1 _1786_ (
    .A(_662_),
    .B(_659_),
    .Y(\step6.myadd.fa8.sum )
);

INVX1 _1787_ (
    .A(\step6.myadd.cin_bF$buf1 ),
    .Y(_664_)
);

NAND2X1 _1788_ (
    .A(\step1.myadd.x0.i0_bF$buf1 ),
    .B(_664_),
    .Y(_665_)
);

INVX1 _1789_ (
    .A(\step1.myadd.x0.i0_bF$buf0 ),
    .Y(_666_)
);

NAND2X1 _1790_ (
    .A(\step6.myadd.cin_bF$buf0 ),
    .B(_666_),
    .Y(_667_)
);

NAND2X1 _1791_ (
    .A(_665_),
    .B(_667_),
    .Y(\step6.myadd.fa1.i1 )
);

INVX1 _1792_ (
    .A(\step6.myadd.cin_bF$buf4 ),
    .Y(_668_)
);

NAND2X1 _1793_ (
    .A(\step1.myadd.x1.i0_bF$buf1 ),
    .B(_668_),
    .Y(_669_)
);

INVX1 _1794_ (
    .A(\step1.myadd.x1.i0_bF$buf0 ),
    .Y(_670_)
);

NAND2X1 _1795_ (
    .A(\step6.myadd.cin_bF$buf3 ),
    .B(_670_),
    .Y(_671_)
);

NAND2X1 _1796_ (
    .A(_669_),
    .B(_671_),
    .Y(\step6.myadd.fa2.i1 )
);

INVX1 _1797_ (
    .A(\step6.myadd.cin_bF$buf2 ),
    .Y(_672_)
);

NAND2X1 _1798_ (
    .A(\step1.myadd.x2.i0_bF$buf1 ),
    .B(_672_),
    .Y(_673_)
);

INVX1 _1799_ (
    .A(\step1.myadd.x2.i0_bF$buf0 ),
    .Y(_674_)
);

NAND2X1 _1800_ (
    .A(\step6.myadd.cin_bF$buf1 ),
    .B(_674_),
    .Y(_675_)
);

NAND2X1 _1801_ (
    .A(_673_),
    .B(_675_),
    .Y(\step6.myadd.fa3.i1 )
);

INVX1 _1802_ (
    .A(\step6.myadd.cin_bF$buf0 ),
    .Y(_676_)
);

NAND2X1 _1803_ (
    .A(\step1.myadd.x3.i0_bF$buf1 ),
    .B(_676_),
    .Y(_677_)
);

INVX1 _1804_ (
    .A(\step1.myadd.x3.i0_bF$buf0 ),
    .Y(_678_)
);

NAND2X1 _1805_ (
    .A(\step6.myadd.cin_bF$buf4 ),
    .B(_678_),
    .Y(_679_)
);

NAND2X1 _1806_ (
    .A(_677_),
    .B(_679_),
    .Y(\step6.myadd.fa4.i1 )
);

INVX1 _1807_ (
    .A(\step6.myadd.cin_bF$buf3 ),
    .Y(_680_)
);

NAND2X1 _1808_ (
    .A(\step1.myadd.x4.i0_bF$buf1 ),
    .B(_680_),
    .Y(_681_)
);

INVX1 _1809_ (
    .A(\step1.myadd.x4.i0_bF$buf0 ),
    .Y(_682_)
);

NAND2X1 _1810_ (
    .A(\step6.myadd.cin_bF$buf2 ),
    .B(_682_),
    .Y(_683_)
);

NAND2X1 _1811_ (
    .A(_681_),
    .B(_683_),
    .Y(\step6.myadd.fa5.i1 )
);

INVX1 _1812_ (
    .A(\step6.myadd.cin_bF$buf1 ),
    .Y(_684_)
);

NAND2X1 _1813_ (
    .A(\step1.myadd.x5.i0_bF$buf1 ),
    .B(_684_),
    .Y(_685_)
);

INVX1 _1814_ (
    .A(\step1.myadd.x5.i0_bF$buf0 ),
    .Y(_686_)
);

NAND2X1 _1815_ (
    .A(\step6.myadd.cin_bF$buf0 ),
    .B(_686_),
    .Y(_687_)
);

NAND2X1 _1816_ (
    .A(_685_),
    .B(_687_),
    .Y(\step6.myadd.fa6.i1 )
);

INVX1 _1817_ (
    .A(\step6.myadd.cin_bF$buf4 ),
    .Y(_688_)
);

NAND2X1 _1818_ (
    .A(\step1.myadd.x6.i0_bF$buf1 ),
    .B(_688_),
    .Y(_689_)
);

INVX1 _1819_ (
    .A(\step1.myadd.x6.i0_bF$buf0 ),
    .Y(_690_)
);

NAND2X1 _1820_ (
    .A(\step6.myadd.cin_bF$buf3 ),
    .B(_690_),
    .Y(_691_)
);

NAND2X1 _1821_ (
    .A(_689_),
    .B(_691_),
    .Y(\step6.myadd.fa7.i1 )
);

INVX1 _1822_ (
    .A(\step6.myadd.cin_bF$buf2 ),
    .Y(_692_)
);

NAND2X1 _1823_ (
    .A(\step1.myadd.x7.i0_bF$buf1 ),
    .B(_692_),
    .Y(_693_)
);

INVX1 _1824_ (
    .A(\step1.myadd.x7.i0_bF$buf0 ),
    .Y(_694_)
);

NAND2X1 _1825_ (
    .A(\step6.myadd.cin_bF$buf1 ),
    .B(_694_),
    .Y(_695_)
);

NAND2X1 _1826_ (
    .A(_693_),
    .B(_695_),
    .Y(\step6.myadd.fa8.i1 )
);

OR2X2 _1827_ (
    .A(\step6.myadd.cin_bF$buf0 ),
    .B(\step7.myadd.cin_bF$buf4 ),
    .Y(_696_)
);

NAND2X1 _1828_ (
    .A(\step6.myadd.cin_bF$buf4 ),
    .B(\step7.myadd.cin_bF$buf3 ),
    .Y(_697_)
);

NAND3X1 _1829_ (
    .A(\step7.myadd.fa2.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_698_)
);

NOR2X1 _1830_ (
    .A(\step6.myadd.cin_bF$buf3 ),
    .B(\step7.myadd.cin_bF$buf2 ),
    .Y(_699_)
);

AND2X2 _1831_ (
    .A(\step6.myadd.cin_bF$buf2 ),
    .B(\step7.myadd.cin_bF$buf1 ),
    .Y(_700_)
);

OAI21X1 _1832_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa2.i0 ),
    .Y(_701_)
);

NAND2X1 _1833_ (
    .A(_701_),
    .B(_698_),
    .Y(\step8.myadd.fa1.i0 )
);

NAND3X1 _1834_ (
    .A(\step7.myadd.fa3.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_702_)
);

OAI21X1 _1835_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa3.i0 ),
    .Y(_703_)
);

NAND2X1 _1836_ (
    .A(_703_),
    .B(_702_),
    .Y(\step8.myadd.fa2.i0 )
);

NAND3X1 _1837_ (
    .A(\step7.myadd.fa4.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_704_)
);

OAI21X1 _1838_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa4.i0 ),
    .Y(_705_)
);

NAND2X1 _1839_ (
    .A(_705_),
    .B(_704_),
    .Y(\step8.myadd.fa3.i0 )
);

NAND3X1 _1840_ (
    .A(\step7.myadd.fa5.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_706_)
);

OAI21X1 _1841_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa5.i0 ),
    .Y(_707_)
);

NAND2X1 _1842_ (
    .A(_707_),
    .B(_706_),
    .Y(\step8.myadd.fa4.i0 )
);

NAND3X1 _1843_ (
    .A(\step7.myadd.fa6.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_708_)
);

OAI21X1 _1844_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa6.i0 ),
    .Y(_709_)
);

NAND2X1 _1845_ (
    .A(_709_),
    .B(_708_),
    .Y(\step8.myadd.fa5.i0 )
);

NAND3X1 _1846_ (
    .A(\step7.myadd.fa7.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_710_)
);

OAI21X1 _1847_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa7.i0 ),
    .Y(_711_)
);

NAND2X1 _1848_ (
    .A(_711_),
    .B(_710_),
    .Y(\step8.myadd.fa6.i0 )
);

NAND3X1 _1849_ (
    .A(\step7.myadd.fa8.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_712_)
);

OAI21X1 _1850_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa7.i0 ),
    .Y(_713_)
);

NAND2X1 _1851_ (
    .A(_713_),
    .B(_712_),
    .Y(\step8.myadd.fa7.i0 )
);

NAND3X1 _1852_ (
    .A(\step7.myadd.fa1.sum ),
    .B(_697_),
    .C(_696_),
    .Y(_714_)
);

OAI21X1 _1853_ (
    .A(_699_),
    .B(_700_),
    .C(\step7.myadd.fa1.i0 ),
    .Y(_715_)
);

NAND2X1 _1854_ (
    .A(_715_),
    .B(_714_),
    .Y(\Q[6] [7])
);

AND2X2 _1855_ (
    .A(\step7.myadd.fa1.i1 ),
    .B(\step7.myadd.cin_bF$buf0 ),
    .Y(_719_)
);

NOR2X1 _1856_ (
    .A(\step7.myadd.fa1.i1 ),
    .B(\step7.myadd.cin_bF$buf4 ),
    .Y(_720_)
);

OAI21X1 _1857_ (
    .A(_720_),
    .B(_719_),
    .C(\step7.myadd.fa1.i0 ),
    .Y(_721_)
);

INVX1 _1858_ (
    .A(\step7.myadd.fa1.i0 ),
    .Y(_722_)
);

NAND2X1 _1859_ (
    .A(\step7.myadd.fa1.i1 ),
    .B(\step7.myadd.cin_bF$buf3 ),
    .Y(_716_)
);

OR2X2 _1860_ (
    .A(\step7.myadd.fa1.i1 ),
    .B(\step7.myadd.cin_bF$buf2 ),
    .Y(_717_)
);

NAND3X1 _1861_ (
    .A(_722_),
    .B(_716_),
    .C(_717_),
    .Y(_718_)
);

NAND2X1 _1862_ (
    .A(_721_),
    .B(_718_),
    .Y(\step7.myadd.fa1.sum )
);

AOI21X1 _1863_ (
    .A(_722_),
    .B(_716_),
    .C(_720_),
    .Y(\step7.myadd.fa1.cout )
);

AND2X2 _1864_ (
    .A(\step7.myadd.fa2.i1 ),
    .B(\step7.myadd.fa1.cout ),
    .Y(_726_)
);

NOR2X1 _1865_ (
    .A(\step7.myadd.fa2.i1 ),
    .B(\step7.myadd.fa1.cout ),
    .Y(_727_)
);

OAI21X1 _1866_ (
    .A(_727_),
    .B(_726_),
    .C(\step7.myadd.fa2.i0 ),
    .Y(_728_)
);

INVX1 _1867_ (
    .A(\step7.myadd.fa2.i0 ),
    .Y(_729_)
);

NAND2X1 _1868_ (
    .A(\step7.myadd.fa2.i1 ),
    .B(\step7.myadd.fa1.cout ),
    .Y(_723_)
);

OR2X2 _1869_ (
    .A(\step7.myadd.fa2.i1 ),
    .B(\step7.myadd.fa1.cout ),
    .Y(_724_)
);

NAND3X1 _1870_ (
    .A(_729_),
    .B(_723_),
    .C(_724_),
    .Y(_725_)
);

NAND2X1 _1871_ (
    .A(_728_),
    .B(_725_),
    .Y(\step7.myadd.fa2.sum )
);

AOI21X1 _1872_ (
    .A(_729_),
    .B(_723_),
    .C(_727_),
    .Y(\step7.myadd.fa2.cout )
);

AND2X2 _1873_ (
    .A(\step7.myadd.fa3.i1 ),
    .B(\step7.myadd.fa2.cout ),
    .Y(_733_)
);

NOR2X1 _1874_ (
    .A(\step7.myadd.fa3.i1 ),
    .B(\step7.myadd.fa2.cout ),
    .Y(_734_)
);

OAI21X1 _1875_ (
    .A(_734_),
    .B(_733_),
    .C(\step7.myadd.fa3.i0 ),
    .Y(_735_)
);

INVX1 _1876_ (
    .A(\step7.myadd.fa3.i0 ),
    .Y(_736_)
);

NAND2X1 _1877_ (
    .A(\step7.myadd.fa3.i1 ),
    .B(\step7.myadd.fa2.cout ),
    .Y(_730_)
);

OR2X2 _1878_ (
    .A(\step7.myadd.fa3.i1 ),
    .B(\step7.myadd.fa2.cout ),
    .Y(_731_)
);

NAND3X1 _1879_ (
    .A(_736_),
    .B(_730_),
    .C(_731_),
    .Y(_732_)
);

NAND2X1 _1880_ (
    .A(_735_),
    .B(_732_),
    .Y(\step7.myadd.fa3.sum )
);

AOI21X1 _1881_ (
    .A(_736_),
    .B(_730_),
    .C(_734_),
    .Y(\step7.myadd.fa3.cout )
);

AND2X2 _1882_ (
    .A(\step7.myadd.fa4.i1 ),
    .B(\step7.myadd.fa3.cout ),
    .Y(_740_)
);

NOR2X1 _1883_ (
    .A(\step7.myadd.fa4.i1 ),
    .B(\step7.myadd.fa3.cout ),
    .Y(_741_)
);

OAI21X1 _1884_ (
    .A(_741_),
    .B(_740_),
    .C(\step7.myadd.fa4.i0 ),
    .Y(_742_)
);

INVX1 _1885_ (
    .A(\step7.myadd.fa4.i0 ),
    .Y(_743_)
);

NAND2X1 _1886_ (
    .A(\step7.myadd.fa4.i1 ),
    .B(\step7.myadd.fa3.cout ),
    .Y(_737_)
);

OR2X2 _1887_ (
    .A(\step7.myadd.fa4.i1 ),
    .B(\step7.myadd.fa3.cout ),
    .Y(_738_)
);

NAND3X1 _1888_ (
    .A(_743_),
    .B(_737_),
    .C(_738_),
    .Y(_739_)
);

NAND2X1 _1889_ (
    .A(_742_),
    .B(_739_),
    .Y(\step7.myadd.fa4.sum )
);

AOI21X1 _1890_ (
    .A(_743_),
    .B(_737_),
    .C(_741_),
    .Y(\step7.myadd.fa4.cout )
);

AND2X2 _1891_ (
    .A(\step7.myadd.fa5.i1 ),
    .B(\step7.myadd.fa4.cout ),
    .Y(_747_)
);

NOR2X1 _1892_ (
    .A(\step7.myadd.fa5.i1 ),
    .B(\step7.myadd.fa4.cout ),
    .Y(_748_)
);

OAI21X1 _1893_ (
    .A(_748_),
    .B(_747_),
    .C(\step7.myadd.fa5.i0 ),
    .Y(_749_)
);

INVX1 _1894_ (
    .A(\step7.myadd.fa5.i0 ),
    .Y(_750_)
);

NAND2X1 _1895_ (
    .A(\step7.myadd.fa5.i1 ),
    .B(\step7.myadd.fa4.cout ),
    .Y(_744_)
);

OR2X2 _1896_ (
    .A(\step7.myadd.fa5.i1 ),
    .B(\step7.myadd.fa4.cout ),
    .Y(_745_)
);

NAND3X1 _1897_ (
    .A(_750_),
    .B(_744_),
    .C(_745_),
    .Y(_746_)
);

NAND2X1 _1898_ (
    .A(_749_),
    .B(_746_),
    .Y(\step7.myadd.fa5.sum )
);

AOI21X1 _1899_ (
    .A(_750_),
    .B(_744_),
    .C(_748_),
    .Y(\step7.myadd.fa5.cout )
);

AND2X2 _1900_ (
    .A(\step7.myadd.fa6.i1 ),
    .B(\step7.myadd.fa5.cout ),
    .Y(_754_)
);

NOR2X1 _1901_ (
    .A(\step7.myadd.fa6.i1 ),
    .B(\step7.myadd.fa5.cout ),
    .Y(_755_)
);

OAI21X1 _1902_ (
    .A(_755_),
    .B(_754_),
    .C(\step7.myadd.fa6.i0 ),
    .Y(_756_)
);

INVX1 _1903_ (
    .A(\step7.myadd.fa6.i0 ),
    .Y(_757_)
);

NAND2X1 _1904_ (
    .A(\step7.myadd.fa6.i1 ),
    .B(\step7.myadd.fa5.cout ),
    .Y(_751_)
);

OR2X2 _1905_ (
    .A(\step7.myadd.fa6.i1 ),
    .B(\step7.myadd.fa5.cout ),
    .Y(_752_)
);

NAND3X1 _1906_ (
    .A(_757_),
    .B(_751_),
    .C(_752_),
    .Y(_753_)
);

NAND2X1 _1907_ (
    .A(_756_),
    .B(_753_),
    .Y(\step7.myadd.fa6.sum )
);

AOI21X1 _1908_ (
    .A(_757_),
    .B(_751_),
    .C(_755_),
    .Y(\step7.myadd.fa6.cout )
);

AND2X2 _1909_ (
    .A(\step7.myadd.fa7.i1 ),
    .B(\step7.myadd.fa6.cout ),
    .Y(_761_)
);

NOR2X1 _1910_ (
    .A(\step7.myadd.fa7.i1 ),
    .B(\step7.myadd.fa6.cout ),
    .Y(_762_)
);

OAI21X1 _1911_ (
    .A(_762_),
    .B(_761_),
    .C(\step7.myadd.fa7.i0 ),
    .Y(_763_)
);

INVX1 _1912_ (
    .A(\step7.myadd.fa7.i0 ),
    .Y(_764_)
);

NAND2X1 _1913_ (
    .A(\step7.myadd.fa7.i1 ),
    .B(\step7.myadd.fa6.cout ),
    .Y(_758_)
);

OR2X2 _1914_ (
    .A(\step7.myadd.fa7.i1 ),
    .B(\step7.myadd.fa6.cout ),
    .Y(_759_)
);

NAND3X1 _1915_ (
    .A(_764_),
    .B(_758_),
    .C(_759_),
    .Y(_760_)
);

NAND2X1 _1916_ (
    .A(_763_),
    .B(_760_),
    .Y(\step7.myadd.fa7.sum )
);

AOI21X1 _1917_ (
    .A(_764_),
    .B(_758_),
    .C(_762_),
    .Y(\step7.myadd.fa7.cout )
);

AND2X2 _1918_ (
    .A(\step7.myadd.fa8.i1 ),
    .B(\step7.myadd.fa7.cout ),
    .Y(_768_)
);

NOR2X1 _1919_ (
    .A(\step7.myadd.fa8.i1 ),
    .B(\step7.myadd.fa7.cout ),
    .Y(_769_)
);

OAI21X1 _1920_ (
    .A(_769_),
    .B(_768_),
    .C(\step7.myadd.fa7.i0 ),
    .Y(_770_)
);

INVX1 _1921_ (
    .A(\step7.myadd.fa7.i0 ),
    .Y(_771_)
);

NAND2X1 _1922_ (
    .A(\step7.myadd.fa8.i1 ),
    .B(\step7.myadd.fa7.cout ),
    .Y(_765_)
);

OR2X2 _1923_ (
    .A(\step7.myadd.fa8.i1 ),
    .B(\step7.myadd.fa7.cout ),
    .Y(_766_)
);

NAND3X1 _1924_ (
    .A(_771_),
    .B(_765_),
    .C(_766_),
    .Y(_767_)
);

NAND2X1 _1925_ (
    .A(_770_),
    .B(_767_),
    .Y(\step7.myadd.fa8.sum )
);

INVX1 _1926_ (
    .A(\step7.myadd.cin_bF$buf1 ),
    .Y(_772_)
);

NAND2X1 _1927_ (
    .A(\step1.myadd.x0.i0_bF$buf3 ),
    .B(_772_),
    .Y(_773_)
);

INVX1 _1928_ (
    .A(\step1.myadd.x0.i0_bF$buf2 ),
    .Y(_774_)
);

NAND2X1 _1929_ (
    .A(\step7.myadd.cin_bF$buf0 ),
    .B(_774_),
    .Y(_775_)
);

NAND2X1 _1930_ (
    .A(_773_),
    .B(_775_),
    .Y(\step7.myadd.fa1.i1 )
);

INVX1 _1931_ (
    .A(\step7.myadd.cin_bF$buf4 ),
    .Y(_776_)
);

NAND2X1 _1932_ (
    .A(\step1.myadd.x1.i0_bF$buf3 ),
    .B(_776_),
    .Y(_777_)
);

INVX1 _1933_ (
    .A(\step1.myadd.x1.i0_bF$buf2 ),
    .Y(_778_)
);

NAND2X1 _1934_ (
    .A(\step7.myadd.cin_bF$buf3 ),
    .B(_778_),
    .Y(_779_)
);

NAND2X1 _1935_ (
    .A(_777_),
    .B(_779_),
    .Y(\step7.myadd.fa2.i1 )
);

INVX1 _1936_ (
    .A(\step7.myadd.cin_bF$buf2 ),
    .Y(_780_)
);

NAND2X1 _1937_ (
    .A(\step1.myadd.x2.i0_bF$buf3 ),
    .B(_780_),
    .Y(_781_)
);

INVX1 _1938_ (
    .A(\step1.myadd.x2.i0_bF$buf2 ),
    .Y(_782_)
);

NAND2X1 _1939_ (
    .A(\step7.myadd.cin_bF$buf1 ),
    .B(_782_),
    .Y(_783_)
);

NAND2X1 _1940_ (
    .A(_781_),
    .B(_783_),
    .Y(\step7.myadd.fa3.i1 )
);

INVX1 _1941_ (
    .A(\step7.myadd.cin_bF$buf0 ),
    .Y(_784_)
);

NAND2X1 _1942_ (
    .A(\step1.myadd.x3.i0_bF$buf3 ),
    .B(_784_),
    .Y(_785_)
);

INVX1 _1943_ (
    .A(\step1.myadd.x3.i0_bF$buf2 ),
    .Y(_786_)
);

NAND2X1 _1944_ (
    .A(\step7.myadd.cin_bF$buf4 ),
    .B(_786_),
    .Y(_787_)
);

NAND2X1 _1945_ (
    .A(_785_),
    .B(_787_),
    .Y(\step7.myadd.fa4.i1 )
);

INVX1 _1946_ (
    .A(\step7.myadd.cin_bF$buf3 ),
    .Y(_788_)
);

NAND2X1 _1947_ (
    .A(\step1.myadd.x4.i0_bF$buf3 ),
    .B(_788_),
    .Y(_789_)
);

INVX1 _1948_ (
    .A(\step1.myadd.x4.i0_bF$buf2 ),
    .Y(_790_)
);

NAND2X1 _1949_ (
    .A(\step7.myadd.cin_bF$buf2 ),
    .B(_790_),
    .Y(_791_)
);

NAND2X1 _1950_ (
    .A(_789_),
    .B(_791_),
    .Y(\step7.myadd.fa5.i1 )
);

INVX1 _1951_ (
    .A(\step7.myadd.cin_bF$buf1 ),
    .Y(_792_)
);

NAND2X1 _1952_ (
    .A(\step1.myadd.x5.i0_bF$buf3 ),
    .B(_792_),
    .Y(_793_)
);

INVX1 _1953_ (
    .A(\step1.myadd.x5.i0_bF$buf2 ),
    .Y(_794_)
);

NAND2X1 _1954_ (
    .A(\step7.myadd.cin_bF$buf0 ),
    .B(_794_),
    .Y(_795_)
);

NAND2X1 _1955_ (
    .A(_793_),
    .B(_795_),
    .Y(\step7.myadd.fa6.i1 )
);

INVX1 _1956_ (
    .A(\step7.myadd.cin_bF$buf4 ),
    .Y(_796_)
);

NAND2X1 _1957_ (
    .A(\step1.myadd.x6.i0_bF$buf3 ),
    .B(_796_),
    .Y(_797_)
);

INVX1 _1958_ (
    .A(\step1.myadd.x6.i0_bF$buf2 ),
    .Y(_798_)
);

NAND2X1 _1959_ (
    .A(\step7.myadd.cin_bF$buf3 ),
    .B(_798_),
    .Y(_799_)
);

NAND2X1 _1960_ (
    .A(_797_),
    .B(_799_),
    .Y(\step7.myadd.fa7.i1 )
);

INVX1 _1961_ (
    .A(\step7.myadd.cin_bF$buf2 ),
    .Y(_800_)
);

NAND2X1 _1962_ (
    .A(\step1.myadd.x7.i0_bF$buf3 ),
    .B(_800_),
    .Y(_801_)
);

INVX1 _1963_ (
    .A(\step1.myadd.x7.i0_bF$buf2 ),
    .Y(_802_)
);

NAND2X1 _1964_ (
    .A(\step7.myadd.cin_bF$buf1 ),
    .B(_802_),
    .Y(_803_)
);

NAND2X1 _1965_ (
    .A(_801_),
    .B(_803_),
    .Y(\step7.myadd.fa8.i1 )
);

OR2X2 _1966_ (
    .A(\step7.myadd.cin_bF$buf0 ),
    .B(qout_bF$buf4),
    .Y(_804_)
);

NAND2X1 _1967_ (
    .A(\step7.myadd.cin_bF$buf4 ),
    .B(qout_bF$buf3),
    .Y(_805_)
);

NAND3X1 _1968_ (
    .A(\step8.myadd.fa2.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_806_)
);

NOR2X1 _1969_ (
    .A(\step7.myadd.cin_bF$buf3 ),
    .B(qout_bF$buf2),
    .Y(_807_)
);

AND2X2 _1970_ (
    .A(\step7.myadd.cin_bF$buf2 ),
    .B(qout_bF$buf1),
    .Y(_808_)
);

OAI21X1 _1971_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa2.i0 ),
    .Y(_809_)
);

NAND2X1 _1972_ (
    .A(_809_),
    .B(_806_),
    .Y(_product[8])
);

NAND3X1 _1973_ (
    .A(\step8.myadd.fa3.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_810_)
);

OAI21X1 _1974_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa3.i0 ),
    .Y(_811_)
);

NAND2X1 _1975_ (
    .A(_811_),
    .B(_810_),
    .Y(_product[9])
);

NAND3X1 _1976_ (
    .A(\step8.myadd.fa4.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_812_)
);

OAI21X1 _1977_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa4.i0 ),
    .Y(_813_)
);

NAND2X1 _1978_ (
    .A(_813_),
    .B(_812_),
    .Y(_product[10])
);

NAND3X1 _1979_ (
    .A(\step8.myadd.fa5.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_814_)
);

OAI21X1 _1980_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa5.i0 ),
    .Y(_815_)
);

NAND2X1 _1981_ (
    .A(_815_),
    .B(_814_),
    .Y(_product[11])
);

NAND3X1 _1982_ (
    .A(\step8.myadd.fa6.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_816_)
);

OAI21X1 _1983_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa6.i0 ),
    .Y(_817_)
);

NAND2X1 _1984_ (
    .A(_817_),
    .B(_816_),
    .Y(_product[12])
);

NAND3X1 _1985_ (
    .A(\step8.myadd.fa7.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_818_)
);

OAI21X1 _1986_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa7.i0 ),
    .Y(_819_)
);

NAND2X1 _1987_ (
    .A(_819_),
    .B(_818_),
    .Y(_product[13])
);

NAND3X1 _1988_ (
    .A(\step8.myadd.fa8.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_820_)
);

OAI21X1 _1989_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa7.i0 ),
    .Y(_821_)
);

NAND2X1 _1990_ (
    .A(_821_),
    .B(_820_),
    .Y(_product[15])
);

NAND3X1 _1991_ (
    .A(\step8.myadd.fa1.sum ),
    .B(_805_),
    .C(_804_),
    .Y(_822_)
);

OAI21X1 _1992_ (
    .A(_807_),
    .B(_808_),
    .C(\step8.myadd.fa1.i0 ),
    .Y(_823_)
);

NAND2X1 _1993_ (
    .A(_823_),
    .B(_822_),
    .Y(_product[7])
);

AND2X2 _1994_ (
    .A(\step8.myadd.fa1.i1 ),
    .B(qout_bF$buf0),
    .Y(_827_)
);

NOR2X1 _1995_ (
    .A(\step8.myadd.fa1.i1 ),
    .B(qout_bF$buf4),
    .Y(_828_)
);

OAI21X1 _1996_ (
    .A(_828_),
    .B(_827_),
    .C(\step8.myadd.fa1.i0 ),
    .Y(_829_)
);

INVX1 _1997_ (
    .A(\step8.myadd.fa1.i0 ),
    .Y(_830_)
);

NAND2X1 _1998_ (
    .A(\step8.myadd.fa1.i1 ),
    .B(qout_bF$buf3),
    .Y(_824_)
);

OR2X2 _1999_ (
    .A(\step8.myadd.fa1.i1 ),
    .B(qout_bF$buf2),
    .Y(_825_)
);

NAND3X1 _2000_ (
    .A(_830_),
    .B(_824_),
    .C(_825_),
    .Y(_826_)
);

NAND2X1 _2001_ (
    .A(_829_),
    .B(_826_),
    .Y(\step8.myadd.fa1.sum )
);

AOI21X1 _2002_ (
    .A(_830_),
    .B(_824_),
    .C(_828_),
    .Y(\step8.myadd.fa1.cout )
);

AND2X2 _2003_ (
    .A(\step8.myadd.fa2.i1 ),
    .B(\step8.myadd.fa1.cout ),
    .Y(_834_)
);

NOR2X1 _2004_ (
    .A(\step8.myadd.fa2.i1 ),
    .B(\step8.myadd.fa1.cout ),
    .Y(_835_)
);

OAI21X1 _2005_ (
    .A(_835_),
    .B(_834_),
    .C(\step8.myadd.fa2.i0 ),
    .Y(_836_)
);

INVX1 _2006_ (
    .A(\step8.myadd.fa2.i0 ),
    .Y(_837_)
);

NAND2X1 _2007_ (
    .A(\step8.myadd.fa2.i1 ),
    .B(\step8.myadd.fa1.cout ),
    .Y(_831_)
);

OR2X2 _2008_ (
    .A(\step8.myadd.fa2.i1 ),
    .B(\step8.myadd.fa1.cout ),
    .Y(_832_)
);

NAND3X1 _2009_ (
    .A(_837_),
    .B(_831_),
    .C(_832_),
    .Y(_833_)
);

NAND2X1 _2010_ (
    .A(_836_),
    .B(_833_),
    .Y(\step8.myadd.fa2.sum )
);

AOI21X1 _2011_ (
    .A(_837_),
    .B(_831_),
    .C(_835_),
    .Y(\step8.myadd.fa2.cout )
);

AND2X2 _2012_ (
    .A(\step8.myadd.fa3.i1 ),
    .B(\step8.myadd.fa2.cout ),
    .Y(_841_)
);

NOR2X1 _2013_ (
    .A(\step8.myadd.fa3.i1 ),
    .B(\step8.myadd.fa2.cout ),
    .Y(_842_)
);

OAI21X1 _2014_ (
    .A(_842_),
    .B(_841_),
    .C(\step8.myadd.fa3.i0 ),
    .Y(_843_)
);

INVX1 _2015_ (
    .A(\step8.myadd.fa3.i0 ),
    .Y(_844_)
);

NAND2X1 _2016_ (
    .A(\step8.myadd.fa3.i1 ),
    .B(\step8.myadd.fa2.cout ),
    .Y(_838_)
);

OR2X2 _2017_ (
    .A(\step8.myadd.fa3.i1 ),
    .B(\step8.myadd.fa2.cout ),
    .Y(_839_)
);

NAND3X1 _2018_ (
    .A(_844_),
    .B(_838_),
    .C(_839_),
    .Y(_840_)
);

NAND2X1 _2019_ (
    .A(_843_),
    .B(_840_),
    .Y(\step8.myadd.fa3.sum )
);

AOI21X1 _2020_ (
    .A(_844_),
    .B(_838_),
    .C(_842_),
    .Y(\step8.myadd.fa3.cout )
);

AND2X2 _2021_ (
    .A(\step8.myadd.fa4.i1 ),
    .B(\step8.myadd.fa3.cout ),
    .Y(_848_)
);

NOR2X1 _2022_ (
    .A(\step8.myadd.fa4.i1 ),
    .B(\step8.myadd.fa3.cout ),
    .Y(_849_)
);

OAI21X1 _2023_ (
    .A(_849_),
    .B(_848_),
    .C(\step8.myadd.fa4.i0 ),
    .Y(_850_)
);

INVX1 _2024_ (
    .A(\step8.myadd.fa4.i0 ),
    .Y(_851_)
);

NAND2X1 _2025_ (
    .A(\step8.myadd.fa4.i1 ),
    .B(\step8.myadd.fa3.cout ),
    .Y(_845_)
);

OR2X2 _2026_ (
    .A(\step8.myadd.fa4.i1 ),
    .B(\step8.myadd.fa3.cout ),
    .Y(_846_)
);

NAND3X1 _2027_ (
    .A(_851_),
    .B(_845_),
    .C(_846_),
    .Y(_847_)
);

NAND2X1 _2028_ (
    .A(_850_),
    .B(_847_),
    .Y(\step8.myadd.fa4.sum )
);

AOI21X1 _2029_ (
    .A(_851_),
    .B(_845_),
    .C(_849_),
    .Y(\step8.myadd.fa4.cout )
);

AND2X2 _2030_ (
    .A(\step8.myadd.fa5.i1 ),
    .B(\step8.myadd.fa4.cout ),
    .Y(_855_)
);

NOR2X1 _2031_ (
    .A(\step8.myadd.fa5.i1 ),
    .B(\step8.myadd.fa4.cout ),
    .Y(_856_)
);

OAI21X1 _2032_ (
    .A(_856_),
    .B(_855_),
    .C(\step8.myadd.fa5.i0 ),
    .Y(_857_)
);

INVX1 _2033_ (
    .A(\step8.myadd.fa5.i0 ),
    .Y(_858_)
);

NAND2X1 _2034_ (
    .A(\step8.myadd.fa5.i1 ),
    .B(\step8.myadd.fa4.cout ),
    .Y(_852_)
);

OR2X2 _2035_ (
    .A(\step8.myadd.fa5.i1 ),
    .B(\step8.myadd.fa4.cout ),
    .Y(_853_)
);

NAND3X1 _2036_ (
    .A(_858_),
    .B(_852_),
    .C(_853_),
    .Y(_854_)
);

NAND2X1 _2037_ (
    .A(_857_),
    .B(_854_),
    .Y(\step8.myadd.fa5.sum )
);

AOI21X1 _2038_ (
    .A(_858_),
    .B(_852_),
    .C(_856_),
    .Y(\step8.myadd.fa5.cout )
);

AND2X2 _2039_ (
    .A(\step8.myadd.fa6.i1 ),
    .B(\step8.myadd.fa5.cout ),
    .Y(_862_)
);

NOR2X1 _2040_ (
    .A(\step8.myadd.fa6.i1 ),
    .B(\step8.myadd.fa5.cout ),
    .Y(_863_)
);

OAI21X1 _2041_ (
    .A(_863_),
    .B(_862_),
    .C(\step8.myadd.fa6.i0 ),
    .Y(_864_)
);

INVX1 _2042_ (
    .A(\step8.myadd.fa6.i0 ),
    .Y(_865_)
);

NAND2X1 _2043_ (
    .A(\step8.myadd.fa6.i1 ),
    .B(\step8.myadd.fa5.cout ),
    .Y(_859_)
);

OR2X2 _2044_ (
    .A(\step8.myadd.fa6.i1 ),
    .B(\step8.myadd.fa5.cout ),
    .Y(_860_)
);

NAND3X1 _2045_ (
    .A(_865_),
    .B(_859_),
    .C(_860_),
    .Y(_861_)
);

NAND2X1 _2046_ (
    .A(_864_),
    .B(_861_),
    .Y(\step8.myadd.fa6.sum )
);

AOI21X1 _2047_ (
    .A(_865_),
    .B(_859_),
    .C(_863_),
    .Y(\step8.myadd.fa6.cout )
);

AND2X2 _2048_ (
    .A(\step8.myadd.fa7.i1 ),
    .B(\step8.myadd.fa6.cout ),
    .Y(_869_)
);

NOR2X1 _2049_ (
    .A(\step8.myadd.fa7.i1 ),
    .B(\step8.myadd.fa6.cout ),
    .Y(_870_)
);

OAI21X1 _2050_ (
    .A(_870_),
    .B(_869_),
    .C(\step8.myadd.fa7.i0 ),
    .Y(_871_)
);

INVX1 _2051_ (
    .A(\step8.myadd.fa7.i0 ),
    .Y(_872_)
);

NAND2X1 _2052_ (
    .A(\step8.myadd.fa7.i1 ),
    .B(\step8.myadd.fa6.cout ),
    .Y(_866_)
);

OR2X2 _2053_ (
    .A(\step8.myadd.fa7.i1 ),
    .B(\step8.myadd.fa6.cout ),
    .Y(_867_)
);

NAND3X1 _2054_ (
    .A(_872_),
    .B(_866_),
    .C(_867_),
    .Y(_868_)
);

NAND2X1 _2055_ (
    .A(_871_),
    .B(_868_),
    .Y(\step8.myadd.fa7.sum )
);

AOI21X1 _2056_ (
    .A(_872_),
    .B(_866_),
    .C(_870_),
    .Y(\step8.myadd.fa7.cout )
);

AND2X2 _2057_ (
    .A(\step8.myadd.fa8.i1 ),
    .B(\step8.myadd.fa7.cout ),
    .Y(_876_)
);

NOR2X1 _2058_ (
    .A(\step8.myadd.fa8.i1 ),
    .B(\step8.myadd.fa7.cout ),
    .Y(_877_)
);

OAI21X1 _2059_ (
    .A(_877_),
    .B(_876_),
    .C(\step8.myadd.fa7.i0 ),
    .Y(_878_)
);

INVX1 _2060_ (
    .A(\step8.myadd.fa7.i0 ),
    .Y(_879_)
);

NAND2X1 _2061_ (
    .A(\step8.myadd.fa8.i1 ),
    .B(\step8.myadd.fa7.cout ),
    .Y(_873_)
);

OR2X2 _2062_ (
    .A(\step8.myadd.fa8.i1 ),
    .B(\step8.myadd.fa7.cout ),
    .Y(_874_)
);

NAND3X1 _2063_ (
    .A(_879_),
    .B(_873_),
    .C(_874_),
    .Y(_875_)
);

NAND2X1 _2064_ (
    .A(_878_),
    .B(_875_),
    .Y(\step8.myadd.fa8.sum )
);

INVX1 _2065_ (
    .A(qout_bF$buf1),
    .Y(_880_)
);

NAND2X1 _2066_ (
    .A(\step1.myadd.x0.i0_bF$buf1 ),
    .B(_880_),
    .Y(_881_)
);

INVX1 _2067_ (
    .A(\step1.myadd.x0.i0_bF$buf0 ),
    .Y(_882_)
);

NAND2X1 _2068_ (
    .A(qout_bF$buf0),
    .B(_882_),
    .Y(_883_)
);

NAND2X1 _2069_ (
    .A(_881_),
    .B(_883_),
    .Y(\step8.myadd.fa1.i1 )
);

INVX1 _2070_ (
    .A(qout_bF$buf4),
    .Y(_884_)
);

NAND2X1 _2071_ (
    .A(\step1.myadd.x1.i0_bF$buf1 ),
    .B(_884_),
    .Y(_885_)
);

INVX1 _2072_ (
    .A(\step1.myadd.x1.i0_bF$buf0 ),
    .Y(_886_)
);

NAND2X1 _2073_ (
    .A(qout_bF$buf3),
    .B(_886_),
    .Y(_887_)
);

NAND2X1 _2074_ (
    .A(_885_),
    .B(_887_),
    .Y(\step8.myadd.fa2.i1 )
);

INVX1 _2075_ (
    .A(qout_bF$buf2),
    .Y(_888_)
);

NAND2X1 _2076_ (
    .A(\step1.myadd.x2.i0_bF$buf1 ),
    .B(_888_),
    .Y(_889_)
);

INVX1 _2077_ (
    .A(\step1.myadd.x2.i0_bF$buf0 ),
    .Y(_890_)
);

NAND2X1 _2078_ (
    .A(qout_bF$buf1),
    .B(_890_),
    .Y(_891_)
);

NAND2X1 _2079_ (
    .A(_889_),
    .B(_891_),
    .Y(\step8.myadd.fa3.i1 )
);

INVX1 _2080_ (
    .A(qout_bF$buf0),
    .Y(_892_)
);

NAND2X1 _2081_ (
    .A(\step1.myadd.x3.i0_bF$buf1 ),
    .B(_892_),
    .Y(_893_)
);

INVX1 _2082_ (
    .A(\step1.myadd.x3.i0_bF$buf0 ),
    .Y(_894_)
);

NAND2X1 _2083_ (
    .A(qout_bF$buf4),
    .B(_894_),
    .Y(_895_)
);

NAND2X1 _2084_ (
    .A(_893_),
    .B(_895_),
    .Y(\step8.myadd.fa4.i1 )
);

INVX1 _2085_ (
    .A(qout_bF$buf3),
    .Y(_896_)
);

NAND2X1 _2086_ (
    .A(\step1.myadd.x4.i0_bF$buf1 ),
    .B(_896_),
    .Y(_897_)
);

INVX1 _2087_ (
    .A(\step1.myadd.x4.i0_bF$buf0 ),
    .Y(_898_)
);

NAND2X1 _2088_ (
    .A(qout_bF$buf2),
    .B(_898_),
    .Y(_899_)
);

NAND2X1 _2089_ (
    .A(_897_),
    .B(_899_),
    .Y(\step8.myadd.fa5.i1 )
);

INVX1 _2090_ (
    .A(qout_bF$buf1),
    .Y(_900_)
);

NAND2X1 _2091_ (
    .A(\step1.myadd.x5.i0_bF$buf1 ),
    .B(_900_),
    .Y(_901_)
);

INVX1 _2092_ (
    .A(\step1.myadd.x5.i0_bF$buf0 ),
    .Y(_902_)
);

NAND2X1 _2093_ (
    .A(qout_bF$buf0),
    .B(_902_),
    .Y(_903_)
);

NAND2X1 _2094_ (
    .A(_901_),
    .B(_903_),
    .Y(\step8.myadd.fa6.i1 )
);

INVX1 _2095_ (
    .A(qout_bF$buf4),
    .Y(_904_)
);

NAND2X1 _2096_ (
    .A(\step1.myadd.x6.i0_bF$buf1 ),
    .B(_904_),
    .Y(_905_)
);

INVX1 _2097_ (
    .A(\step1.myadd.x6.i0_bF$buf0 ),
    .Y(_906_)
);

NAND2X1 _2098_ (
    .A(qout_bF$buf3),
    .B(_906_),
    .Y(_907_)
);

NAND2X1 _2099_ (
    .A(_905_),
    .B(_907_),
    .Y(\step8.myadd.fa7.i1 )
);

INVX1 _2100_ (
    .A(qout_bF$buf2),
    .Y(_908_)
);

NAND2X1 _2101_ (
    .A(\step1.myadd.x7.i0_bF$buf1 ),
    .B(_908_),
    .Y(_909_)
);

INVX1 _2102_ (
    .A(\step1.myadd.x7.i0_bF$buf0 ),
    .Y(_910_)
);

NAND2X1 _2103_ (
    .A(qout_bF$buf1),
    .B(_910_),
    .Y(_911_)
);

NAND2X1 _2104_ (
    .A(_909_),
    .B(_911_),
    .Y(\step8.myadd.fa8.i1 )
);

BUFX2 _2105_ (
    .A(_912_[0]),
    .Y(product[0])
);

BUFX2 _2106_ (
    .A(_912_[1]),
    .Y(product[1])
);

BUFX2 _2107_ (
    .A(_912_[10]),
    .Y(product[10])
);

BUFX2 _2108_ (
    .A(_912_[11]),
    .Y(product[11])
);

BUFX2 _2109_ (
    .A(_912_[12]),
    .Y(product[12])
);

BUFX2 _2110_ (
    .A(_912_[13]),
    .Y(product[13])
);

BUFX2 _2111_ (
    .A(_912_[14]),
    .Y(product[14])
);

BUFX2 _2112_ (
    .A(_912_[15]),
    .Y(product[15])
);

BUFX2 _2113_ (
    .A(_912_[2]),
    .Y(product[2])
);

BUFX2 _2114_ (
    .A(_912_[3]),
    .Y(product[3])
);

BUFX2 _2115_ (
    .A(_912_[4]),
    .Y(product[4])
);

BUFX2 _2116_ (
    .A(_912_[5]),
    .Y(product[5])
);

BUFX2 _2117_ (
    .A(_912_[6]),
    .Y(product[6])
);

BUFX2 _2118_ (
    .A(_912_[7]),
    .Y(product[7])
);

BUFX2 _2119_ (
    .A(_912_[8]),
    .Y(product[8])
);

BUFX2 _2120_ (
    .A(_912_[9]),
    .Y(product[9])
);

INVX1 _913_ (
    .A(\step1.myadd.cin_bF$buf0 ),
    .Y(_16_)
);

NAND2X1 _914_ (
    .A(multIn[0]),
    .B(select_bF$buf4),
    .Y(_17_)
);

OAI21X1 _915_ (
    .A(select_bF$buf3),
    .B(_16_),
    .C(_17_),
    .Y(_8_)
);

INVX1 _916_ (
    .A(\step2.myadd.cin_bF$buf1 ),
    .Y(_18_)
);

NAND2X1 _917_ (
    .A(select_bF$buf2),
    .B(multIn[1]),
    .Y(_19_)
);

OAI21X1 _918_ (
    .A(select_bF$buf1),
    .B(_18_),
    .C(_19_),
    .Y(_9_)
);

INVX1 _919_ (
    .A(\step3.myadd.cin_bF$buf1 ),
    .Y(_20_)
);

NAND2X1 _920_ (
    .A(select_bF$buf0),
    .B(multIn[2]),
    .Y(_21_)
);

OAI21X1 _921_ (
    .A(select_bF$buf4),
    .B(_20_),
    .C(_21_),
    .Y(_10_)
);

INVX1 _922_ (
    .A(\step4.myadd.cin_bF$buf1 ),
    .Y(_22_)
);

NAND2X1 _923_ (
    .A(select_bF$buf3),
    .B(multIn[3]),
    .Y(_23_)
);

OAI21X1 _924_ (
    .A(select_bF$buf2),
    .B(_22_),
    .C(_23_),
    .Y(_11_)
);

INVX1 _925_ (
    .A(\step5.myadd.cin_bF$buf1 ),
    .Y(_24_)
);

NAND2X1 _926_ (
    .A(select_bF$buf1),
    .B(multIn[4]),
    .Y(_25_)
);

OAI21X1 _927_ (
    .A(select_bF$buf0),
    .B(_24_),
    .C(_25_),
    .Y(_12_)
);

INVX1 _928_ (
    .A(\step6.myadd.cin_bF$buf1 ),
    .Y(_26_)
);

NAND2X1 _929_ (
    .A(select_bF$buf4),
    .B(multIn[5]),
    .Y(_27_)
);

OAI21X1 _930_ (
    .A(select_bF$buf3),
    .B(_26_),
    .C(_27_),
    .Y(_13_)
);

INVX1 _931_ (
    .A(\step7.myadd.cin_bF$buf1 ),
    .Y(_28_)
);

NAND2X1 _932_ (
    .A(select_bF$buf2),
    .B(multIn[6]),
    .Y(_29_)
);

OAI21X1 _933_ (
    .A(select_bF$buf1),
    .B(_28_),
    .C(_29_),
    .Y(_14_)
);

INVX1 _934_ (
    .A(qout_bF$buf0),
    .Y(_30_)
);

NAND2X1 _935_ (
    .A(select_bF$buf0),
    .B(multIn[7]),
    .Y(_31_)
);

OAI21X1 _936_ (
    .A(select_bF$buf4),
    .B(_30_),
    .C(_31_),
    .Y(_15_)
);

INVX1 _937_ (
    .A(multIn[0]),
    .Y(_32_)
);

NAND2X1 _938_ (
    .A(select_bF$buf3),
    .B(\step1.myadd.x0.i0_bF$buf3 ),
    .Y(_33_)
);

OAI21X1 _939_ (
    .A(select_bF$buf2),
    .B(_32_),
    .C(_33_),
    .Y(_0_)
);

INVX1 _940_ (
    .A(multIn[1]),
    .Y(_34_)
);

NAND2X1 _941_ (
    .A(select_bF$buf1),
    .B(\step1.myadd.x1.i0_bF$buf3 ),
    .Y(_35_)
);

OAI21X1 _942_ (
    .A(select_bF$buf0),
    .B(_34_),
    .C(_35_),
    .Y(_1_)
);

INVX1 _943_ (
    .A(multIn[2]),
    .Y(_36_)
);

NAND2X1 _944_ (
    .A(select_bF$buf4),
    .B(\step1.myadd.x2.i0_bF$buf3 ),
    .Y(_37_)
);

OAI21X1 _945_ (
    .A(select_bF$buf3),
    .B(_36_),
    .C(_37_),
    .Y(_2_)
);

INVX1 _946_ (
    .A(multIn[3]),
    .Y(_38_)
);

NAND2X1 _947_ (
    .A(select_bF$buf2),
    .B(\step1.myadd.x3.i0_bF$buf3 ),
    .Y(_39_)
);

OAI21X1 _948_ (
    .A(select_bF$buf1),
    .B(_38_),
    .C(_39_),
    .Y(_3_)
);

INVX1 _949_ (
    .A(multIn[4]),
    .Y(_40_)
);

NAND2X1 _950_ (
    .A(select_bF$buf0),
    .B(\step1.myadd.x4.i0_bF$buf3 ),
    .Y(_41_)
);

OAI21X1 _951_ (
    .A(select_bF$buf4),
    .B(_40_),
    .C(_41_),
    .Y(_4_)
);

INVX1 _952_ (
    .A(multIn[5]),
    .Y(_42_)
);

NAND2X1 _953_ (
    .A(select_bF$buf3),
    .B(\step1.myadd.x5.i0_bF$buf3 ),
    .Y(_43_)
);

OAI21X1 _954_ (
    .A(select_bF$buf2),
    .B(_42_),
    .C(_43_),
    .Y(_5_)
);

INVX1 _955_ (
    .A(multIn[6]),
    .Y(_44_)
);

NAND2X1 _956_ (
    .A(select_bF$buf1),
    .B(\step1.myadd.x6.i0_bF$buf3 ),
    .Y(_45_)
);

OAI21X1 _957_ (
    .A(select_bF$buf0),
    .B(_44_),
    .C(_45_),
    .Y(_6_)
);

INVX1 _958_ (
    .A(multIn[7]),
    .Y(_46_)
);

NAND2X1 _959_ (
    .A(select_bF$buf4),
    .B(\step1.myadd.x7.i0_bF$buf3 ),
    .Y(_47_)
);

OAI21X1 _960_ (
    .A(select_bF$buf3),
    .B(_46_),
    .C(_47_),
    .Y(_7_)
);

DFFPOSX1 _961_ (
    .CLK(clk_bF$buf4),
    .D(_0_),
    .Q(\step1.myadd.x0.i0 )
);

DFFPOSX1 _962_ (
    .CLK(clk_bF$buf3),
    .D(_1_),
    .Q(\step1.myadd.x1.i0 )
);

DFFPOSX1 _963_ (
    .CLK(clk_bF$buf2),
    .D(_2_),
    .Q(\step1.myadd.x2.i0 )
);

DFFPOSX1 _964_ (
    .CLK(clk_bF$buf1),
    .D(_3_),
    .Q(\step1.myadd.x3.i0 )
);

DFFPOSX1 _965_ (
    .CLK(clk_bF$buf0),
    .D(_4_),
    .Q(\step1.myadd.x4.i0 )
);

DFFPOSX1 _966_ (
    .CLK(clk_bF$buf4),
    .D(_5_),
    .Q(\step1.myadd.x5.i0 )
);

DFFPOSX1 _967_ (
    .CLK(clk_bF$buf3),
    .D(_6_),
    .Q(\step1.myadd.x6.i0 )
);

DFFPOSX1 _968_ (
    .CLK(clk_bF$buf2),
    .D(_7_),
    .Q(\step1.myadd.x7.i0 )
);

DFFPOSX1 _969_ (
    .CLK(clk_bF$buf1),
    .D(\Q[0] [7]),
    .Q(_912_[0])
);

DFFPOSX1 _970_ (
    .CLK(clk_bF$buf0),
    .D(\Q[1] [7]),
    .Q(_912_[1])
);

DFFPOSX1 _971_ (
    .CLK(clk_bF$buf4),
    .D(\Q[2] [7]),
    .Q(_912_[2])
);

DFFPOSX1 _972_ (
    .CLK(clk_bF$buf3),
    .D(\Q[3] [7]),
    .Q(_912_[3])
);

DFFPOSX1 _973_ (
    .CLK(clk_bF$buf2),
    .D(\Q[4] [7]),
    .Q(_912_[4])
);

DFFPOSX1 _974_ (
    .CLK(clk_bF$buf1),
    .D(\Q[5] [7]),
    .Q(_912_[5])
);

DFFPOSX1 _975_ (
    .CLK(clk_bF$buf0),
    .D(\Q[6] [7]),
    .Q(_912_[6])
);

DFFPOSX1 _976_ (
    .CLK(clk_bF$buf4),
    .D(_product[7]),
    .Q(_912_[7])
);

DFFPOSX1 _977_ (
    .CLK(clk_bF$buf3),
    .D(_product[8]),
    .Q(_912_[8])
);

DFFPOSX1 _978_ (
    .CLK(clk_bF$buf2),
    .D(_product[9]),
    .Q(_912_[9])
);

DFFPOSX1 _979_ (
    .CLK(clk_bF$buf1),
    .D(_product[10]),
    .Q(_912_[10])
);

DFFPOSX1 _980_ (
    .CLK(clk_bF$buf0),
    .D(_product[11]),
    .Q(_912_[11])
);

DFFPOSX1 _981_ (
    .CLK(clk_bF$buf4),
    .D(_product[12]),
    .Q(_912_[12])
);

DFFPOSX1 _982_ (
    .CLK(clk_bF$buf3),
    .D(_product[13]),
    .Q(_912_[13])
);

DFFPOSX1 _983_ (
    .CLK(clk_bF$buf2),
    .D(_product[15]),
    .Q(_912_[14])
);

DFFPOSX1 _984_ (
    .CLK(clk_bF$buf1),
    .D(_product[15]),
    .Q(_912_[15])
);

DFFPOSX1 _985_ (
    .CLK(clk_bF$buf0),
    .D(_8_),
    .Q(\step1.myadd.cin )
);

DFFPOSX1 _986_ (
    .CLK(clk_bF$buf4),
    .D(_9_),
    .Q(\step2.myadd.cin )
);

DFFPOSX1 _987_ (
    .CLK(clk_bF$buf3),
    .D(_10_),
    .Q(\step3.myadd.cin )
);

DFFPOSX1 _988_ (
    .CLK(clk_bF$buf2),
    .D(_11_),
    .Q(\step4.myadd.cin )
);

DFFPOSX1 _989_ (
    .CLK(clk_bF$buf1),
    .D(_12_),
    .Q(\step5.myadd.cin )
);

DFFPOSX1 _990_ (
    .CLK(clk_bF$buf0),
    .D(_13_),
    .Q(\step6.myadd.cin )
);

DFFPOSX1 _991_ (
    .CLK(clk_bF$buf4),
    .D(_14_),
    .Q(\step7.myadd.cin )
);

DFFPOSX1 _992_ (
    .CLK(clk_bF$buf3),
    .D(_15_),
    .Q(qout)
);

OR2X2 _993_ (
    .A(gnd),
    .B(\step1.myadd.cin_bF$buf4 ),
    .Y(_48_)
);

NAND2X1 _994_ (
    .A(gnd),
    .B(\step1.myadd.cin_bF$buf3 ),
    .Y(_49_)
);

NAND3X1 _995_ (
    .A(\step1.myadd.fa2.sum ),
    .B(_49_),
    .C(_48_),
    .Y(_50_)
);

NOR2X1 _996_ (
    .A(gnd),
    .B(\step1.myadd.cin_bF$buf2 ),
    .Y(_51_)
);

AND2X2 _997_ (
    .A(gnd),
    .B(\step1.myadd.cin_bF$buf1 ),
    .Y(_52_)
);

OAI21X1 _998_ (
    .A(_51_),
    .B(_52_),
    .C(gnd),
    .Y(_53_)
);

NAND2X1 _999_ (
    .A(_53_),
    .B(_50_),
    .Y(\step2.myadd.fa1.i0 )
);

endmodule
