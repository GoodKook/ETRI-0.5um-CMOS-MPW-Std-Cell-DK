* NGSPICE file created from ALU_wrapper.ext - technology: scmos

* Black-box entry subcircuit for FILL abstract view
.subckt FILL gnd vdd
.ends

* Black-box entry subcircuit for NAND2X1 abstract view
.subckt NAND2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX1 abstract view
.subckt INVX1 A Y vdd gnd
.ends

* Black-box entry subcircuit for AOI21X1 abstract view
.subckt AOI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for OAI21X1 abstract view
.subckt OAI21X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for NAND3X1 abstract view
.subckt NAND3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for BUFX2 abstract view
.subckt BUFX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for NOR2X1 abstract view
.subckt NOR2X1 A B Y vdd gnd
.ends

* Black-box entry subcircuit for NOR3X1 abstract view
.subckt NOR3X1 A B C Y vdd gnd
.ends

* Black-box entry subcircuit for AOI22X1 abstract view
.subckt AOI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for INVX2 abstract view
.subckt INVX2 A Y vdd gnd
.ends

* Black-box entry subcircuit for AND2X2 abstract view
.subckt AND2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for OR2X2 abstract view
.subckt OR2X2 A B Y vdd gnd
.ends

* Black-box entry subcircuit for INVX4 abstract view
.subckt INVX4 A Y vdd gnd
.ends

* Black-box entry subcircuit for DFFPOSX1 abstract view
.subckt DFFPOSX1 D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for CLKBUF1 abstract view
.subckt CLKBUF1 A Y vdd gnd
.ends

* Black-box entry subcircuit for OAI22X1 abstract view
.subckt OAI22X1 A B C D Y vdd gnd
.ends

* Black-box entry subcircuit for DFFSR abstract view
.subckt DFFSR R S D CLK Q vdd gnd
.ends

* Black-box entry subcircuit for MUX2X1 abstract view
.subckt MUX2X1 A B S Y vdd gnd
.ends

.subckt ALU_wrapper gnd vdd ABCmd_i[7] ABCmd_i[6] ABCmd_i[5] ABCmd_i[4] ABCmd_i[3]
+ ABCmd_i[2] ABCmd_i[1] ABCmd_i[0] ACC_o[7] ACC_o[6] ACC_o[5] ACC_o[4] ACC_o[3] ACC_o[2]
+ ACC_o[1] ACC_o[0] Done_o LoadA_i LoadB_i LoadCmd_i clk reset
XFILL_0__1759_ gnd vdd FILL
X_1270_ _1288_/B _1288_/A _1374_/A vdd gnd NAND2X1
X_1606_ _1606_/A _1641_/C vdd gnd INVX1
X_1399_ _1399_/A _1416_/A _1470_/B _1407_/A vdd gnd AOI21X1
X_1468_ _1567_/B _1468_/B _1572_/A vdd gnd NAND2X1
X_1537_ _1537_/A _1537_/B _1562_/C vdd gnd NAND2X1
X_981_ _981_/A _984_/B _981_/C _981_/Y vdd gnd OAI21X1
X_1184_ _1184_/A _1343_/A _998_/A _1203_/A vdd gnd OAI21X1
XFILL_0__1527_ gnd vdd FILL
X_1322_ _1564_/A _1574_/A _1323_/A vdd gnd NAND2X1
X_1253_ _1253_/A _1338_/C _1253_/C _1298_/A vdd gnd NAND3X1
X_964_ ABCmd_i[0] _966_/A vdd gnd INVX1
X_1871_ _1874_/B _1874_/A _1871_/C _1872_/C vdd gnd NAND3X1
XFILL_0__1174_ gnd vdd FILL
XBUFX2_insert0 _1668_/Q _974_/A vdd gnd BUFX2
X_1236_ _1236_/A _1236_/B _1236_/C _1238_/C vdd gnd OAI21X1
X_1098_ _991_/A _1621_/B _1101_/B vdd gnd NOR2X1
X_1167_ _1245_/B _1167_/B _1246_/A vdd gnd NAND2X1
X_1305_ _1308_/C _1308_/B _1337_/A _1306_/B vdd gnd AOI21X1
X_947_ _953_/B _947_/B _962_/A _948_/C vdd gnd OAI21X1
X_1785_ _1785_/A _1802_/C _1785_/C _1786_/C vdd gnd AOI21X1
X_1854_ _1869_/B _1874_/A vdd gnd INVX1
X_1219_ _1610_/A _1241_/A _1241_/B _1632_/A vdd gnd NOR3X1
X_1021_ _995_/A _1813_/A _1067_/C _1794_/A _1055_/A vdd gnd AOI22X1
XFILL_0__1775_ gnd vdd FILL
XFILL_0__977_ gnd vdd FILL
XFILL_0__1844_ gnd vdd FILL
X_1004_ _995_/A _1794_/A _994_/A _995_/B _1186_/A vdd gnd AOI22X1
XFILL_0__1011_ gnd vdd FILL
X_1570_ _1626_/A _1604_/A vdd gnd INVX1
X_1699_ ABCmd_i[0] _1843_/A vdd gnd INVX2
X_1768_ _1801_/B _1801_/A _1802_/B vdd gnd AND2X2
X_1837_ _1841_/C _1874_/B vdd gnd INVX1
XFILL_0__1209_ gnd vdd FILL
X_1622_ _1640_/B _1640_/A _1624_/B vdd gnd OR2X2
X_1484_ _1893_/Y _1485_/A vdd gnd INVX1
X_1553_ _1592_/A _1555_/A _1557_/A vdd gnd NAND2X1
XFILL_0__1612_ gnd vdd FILL
X_1536_ _1898_/A _1585_/A vdd gnd INVX1
X_1605_ _1617_/A _1626_/B _1605_/C _1609_/C vdd gnd NAND3X1
X_1467_ _1467_/A _1519_/B _1467_/C _1567_/B vdd gnd NAND3X1
X_1398_ _1398_/A _1416_/C _1470_/B vdd gnd NOR2X1
X_980_ _980_/A _984_/B _981_/C vdd gnd NAND2X1
X_1183_ _995_/A _1184_/A vdd gnd INVX1
X_1321_ _1416_/A _1321_/B _1564_/A vdd gnd NAND2X1
X_1252_ _1255_/B _1255_/A _1253_/C vdd gnd OR2X2
XFILL_0__1457_ gnd vdd FILL
XFILL76350x28950 gnd vdd FILL
X_1519_ _1521_/C _1519_/B _1519_/C _1573_/A vdd gnd NAND3X1
X_963_ reset _963_/Y vdd gnd INVX1
X_1870_ _1876_/A _1872_/B vdd gnd INVX1
X_1235_ _1580_/A _1580_/C _1580_/B _1610_/C vdd gnd NOR3X1
X_1097_ _983_/A _1621_/B vdd gnd INVX4
XBUFX2_insert1 _1668_/Q _1439_/B vdd gnd BUFX2
X_1304_ _1304_/A _1304_/B _1336_/C _1308_/B vdd gnd OAI21X1
X_1166_ _1166_/A _1166_/B _1166_/C _1167_/B vdd gnd NAND3X1
XFILL_0__1860_ gnd vdd FILL
X_946_ LoadCmd_i _962_/A vdd gnd INVX1
X_1784_ ABCmd_i[6] _1785_/C vdd gnd INVX1
X_1853_ _1874_/B _1871_/C _1864_/C vdd gnd NAND2X1
X_1020_ _1067_/C _1794_/A _1057_/A _1055_/C vdd gnd NAND3X1
X_1218_ _1315_/B _1315_/A _1218_/C _1241_/B vdd gnd AOI21X1
X_1149_ _1163_/B _1163_/C _1163_/A _1246_/C vdd gnd NAND3X1
X_929_ _953_/A _941_/A _930_/A vdd gnd NAND2X1
X_1003_ _998_/B _1027_/A _1187_/C vdd gnd OR2X2
X_1698_ ABCmd_i[0] _1845_/A _1845_/D vdd gnd NAND2X1
X_1767_ _1787_/A _1780_/A vdd gnd INVX1
X_1836_ _1836_/A _1836_/B _1836_/C _1875_/A vdd gnd OAI21X1
XFILL_0__1139_ gnd vdd FILL
XFILL76050x25350 gnd vdd FILL
X_1483_ _1897_/A _1535_/A vdd gnd INVX1
X_1621_ _1621_/A _1621_/B _1621_/C _1640_/A vdd gnd OAI21X1
X_1552_ _1552_/A _1552_/B _1552_/C _1592_/A vdd gnd NAND3X1
X_1819_ _1836_/A _1836_/B _1824_/A _1823_/A vdd gnd OAI21X1
X_1535_ _1535_/A _949_/A _1535_/C _1535_/D _1676_/D vdd gnd AOI22X1
X_1604_ _1604_/A _1604_/B _1604_/C _1605_/C vdd gnd NAND3X1
XFILL_0__1542_ gnd vdd FILL
X_1466_ _1466_/A _1466_/B _1466_/C _1467_/C vdd gnd OAI21X1
X_1397_ _1401_/A _1397_/B _1403_/B _1403_/A _1398_/A vdd gnd AOI22X1
X_1182_ _999_/A _1203_/B vdd gnd INVX1
X_1320_ _1642_/C _1642_/A _1643_/A _1574_/A vdd gnd AOI21X1
X_1251_ _1255_/A _1255_/B _1338_/C vdd gnd NAND2X1
XFILL_0__1387_ gnd vdd FILL
X_1518_ _1537_/B _1522_/A _1519_/C vdd gnd NAND2X1
X_1449_ _1449_/A _1449_/B _1456_/B vdd gnd NAND2X1
X_962_ _962_/A _962_/B _962_/C _962_/Y vdd gnd OAI21X1
XFILL_0__1310_ gnd vdd FILL
X_1234_ _1234_/A _1234_/B _1234_/C _1580_/A vdd gnd AOI21X1
X_1096_ _1104_/B _1104_/A _1104_/C _1197_/C vdd gnd NAND3X1
XBUFX2_insert2 _1668_/Q _990_/A vdd gnd BUFX2
X_1303_ _1336_/A _1336_/B _1303_/C _1308_/C vdd gnd NAND3X1
X_1165_ _1165_/A _1165_/B _1245_/A _1245_/B vdd gnd NAND3X1
XFILL_0__992_ gnd vdd FILL
XFILL_0__1790_ gnd vdd FILL
X_945_ _960_/C _952_/C vdd gnd INVX1
X_1783_ _1858_/A _1783_/Y vdd gnd INVX1
XFILL_0__1224_ gnd vdd FILL
X_1852_ _1865_/A _1865_/B _1869_/B _1886_/C vdd gnd OAI21X1
XFILL_0__1155_ gnd vdd FILL
X_1217_ _1316_/B _1580_/B _1217_/C _1610_/A vdd gnd NAND3X1
X_1079_ _995_/B _1343_/A vdd gnd INVX2
X_1148_ _1258_/C _1287_/B _1287_/A _1163_/A vdd gnd OAI21X1
X_928_ _942_/B _942_/C _941_/A vdd gnd NOR2X1
X_1697_ ABCmd_i[1] _1845_/A vdd gnd INVX2
X_1766_ _1785_/A _1766_/Y vdd gnd INVX1
X_1835_ _1841_/C _1871_/C _1861_/B vdd gnd NAND2X1
X_1002_ _1067_/C _1794_/A _1027_/A vdd gnd NAND2X1
XFILL_0__1069_ gnd vdd FILL
XFILL_0__958_ gnd vdd FILL
X_1482_ _949_/A _1482_/B _1482_/C _1675_/D vdd gnd OAI21X1
XFILL_0__1825_ gnd vdd FILL
X_1620_ _1620_/A _1640_/B vdd gnd INVX1
X_1551_ _1593_/A _1552_/A vdd gnd INVX1
X_1749_ ABCmd_i[5] _995_/B _1755_/C vdd gnd NAND2X1
X_1818_ _1818_/A _1818_/B _1875_/B _1824_/A vdd gnd OAI21X1
XFILL76650x150 gnd vdd FILL
XFILL_0__1472_ gnd vdd FILL
X_1534_ _1534_/A _937_/A _949_/A _1535_/D vdd gnd AOI21X1
X_1603_ _1604_/B _1603_/B _1604_/C _1639_/A vdd gnd NAND3X1
X_1396_ _1396_/A _1396_/B _1396_/C _1403_/B vdd gnd NAND3X1
X_1465_ _1465_/A _1465_/B _1465_/C _1466_/B vdd gnd AOI21X1
X_1181_ _998_/A _998_/B _1208_/A vdd gnd NOR2X1
X_1250_ _1250_/A _1250_/B _1250_/C _1255_/B vdd gnd OAI21X1
X_1448_ _1454_/A _1454_/B _1489_/A vdd gnd AND2X2
X_1517_ _1517_/A _1537_/A _1517_/C _1537_/B vdd gnd NAND3X1
X_961_ _961_/A _961_/B _962_/C vdd gnd AND2X2
X_1379_ _1386_/C _1385_/C _1420_/B vdd gnd NAND2X1
X_1095_ _1146_/B _1111_/C _1146_/A _1104_/A vdd gnd OAI21X1
X_1233_ _1478_/B _1529_/A _1529_/B _1580_/C vdd gnd NAND3X1
XFILL_0__1240_ gnd vdd FILL
XBUFX2_insert3 _1668_/Q _1131_/A vdd gnd BUFX2
X_1164_ _1164_/A _1164_/B _1164_/C _1297_/C vdd gnd AOI21X1
X_1302_ _1402_/A _1337_/A vdd gnd INVX1
XFILL_0__1507_ gnd vdd FILL
XFILL_0__1438_ gnd vdd FILL
XFILL76650x57750 gnd vdd FILL
X_944_ _953_/A _949_/A _960_/C vdd gnd NOR2X1
X_1851_ _1881_/B _1880_/A _1869_/C _1869_/B vdd gnd OAI21X1
X_1782_ _1786_/B _1786_/A _1858_/A vdd gnd NAND2X1
X_1216_ _1236_/A _1236_/B _993_/Y _1217_/C vdd gnd OAI21X1
XFILL_0__1085_ gnd vdd FILL
X_1078_ _1083_/C _1084_/C _1082_/C vdd gnd NAND2X1
X_1147_ _1287_/C _1258_/B _1258_/A _1163_/B vdd gnd NAND3X1
XFILL76650x32550 gnd vdd FILL
X_1696_ _1741_/D _1720_/A vdd gnd INVX1
X_1765_ _1787_/B _1765_/B _1785_/A vdd gnd NAND2X1
X_927_ _936_/A _942_/C vdd gnd INVX1
X_1834_ _1834_/A _1834_/B _1869_/A _1841_/C vdd gnd OAI21X1
XFILL_0__1841_ gnd vdd FILL
X_1001_ _1187_/A _1186_/C vdd gnd INVX1
XFILL_0__1755_ gnd vdd FILL
X_1481_ _1481_/A _1481_/B _1481_/C _1481_/D _1482_/B vdd gnd AOI22X1
X_1550_ _1590_/A _1550_/B _1593_/B _1555_/A vdd gnd OAI21X1
X_1748_ _1748_/A _1748_/B _1764_/A _1801_/B vdd gnd OAI21X1
X_1817_ _1881_/A _1818_/B _1818_/A _1875_/B vdd gnd OAI21X1
X_1679_ _1679_/D _1680_/CLK _1900_/A vdd gnd DFFPOSX1
XFILL76350x54150 gnd vdd FILL
X_1533_ _987_/A _1533_/B _1533_/C _1534_/A vdd gnd OAI21X1
X_1602_ _1626_/B _1626_/A _1603_/B vdd gnd NOR2X1
X_1395_ _1466_/A _1466_/C _1395_/C _1403_/A vdd gnd NAND3X1
X_1464_ _1466_/C _1464_/B _1464_/C _1468_/B vdd gnd NAND3X1
X_1180_ _993_/Y _1236_/C vdd gnd INVX1
XFILL_0__1523_ gnd vdd FILL
X_1516_ _1516_/A _1555_/C _1516_/C _1517_/C vdd gnd OAI21X1
X_960_ _960_/A _960_/B _960_/C _961_/B vdd gnd NAND3X1
X_1447_ _1489_/C _1511_/B _1511_/A _1520_/B vdd gnd OAI21X1
X_1378_ _1385_/A _1449_/B _1378_/C _1453_/C vdd gnd NAND3X1
X_1232_ _1232_/A _1232_/B _1232_/C _1529_/A vdd gnd OAI21X1
X_1301_ _1401_/A _1402_/B _1402_/A _1306_/A vdd gnd AOI21X1
XFILL_0__1170_ gnd vdd FILL
XBUFX2_insert4 _1665_/Q _965_/A vdd gnd BUFX2
X_1094_ _1146_/C _1111_/A _1111_/B _1104_/B vdd gnd NAND3X1
X_1163_ _1163_/A _1163_/B _1163_/C _1246_/B vdd gnd AOI21X1
XFILL_0__1368_ gnd vdd FILL
X_943_ LoadB_i _960_/B vdd gnd INVX1
X_1781_ _1787_/A _1781_/B _1787_/B _1786_/B vdd gnd NAND3X1
X_1850_ _1881_/A _1880_/A _1881_/B _1869_/C vdd gnd OAI21X1
X_1215_ _1215_/A _1234_/B _1215_/C _1215_/D _1236_/A vdd gnd AOI22X1
X_1077_ _990_/A _995_/B _1084_/C vdd gnd AND2X2
X_1146_ _1146_/A _1146_/B _1146_/C _1163_/C vdd gnd OAI21X1
XFILL_0__973_ gnd vdd FILL
X_1764_ _1764_/A _1764_/B _1764_/C _1765_/B vdd gnd NAND3X1
XFILL_0__1771_ gnd vdd FILL
X_1902_ _947_/B Done_o vdd gnd BUFX2
XFILL_0__1205_ gnd vdd FILL
X_1833_ _1881_/A _1834_/B _1834_/A _1869_/A vdd gnd OAI21X1
X_1000_ _997_/A _994_/B _1187_/A vdd gnd NAND2X1
X_1695_ ABCmd_i[5] _1716_/B _1741_/D vdd gnd NOR2X1
X_1129_ _1131_/A _1794_/A _1136_/C vdd gnd AND2X2
X_1480_ _1480_/A _952_/C _1481_/B vdd gnd NOR2X1
X_1747_ _1747_/A _1747_/B _1748_/A vdd gnd NOR2X1
X_1816_ _1848_/A _980_/A _1816_/C _1818_/B vdd gnd AOI21X1
X_1678_ _1678_/D _1680_/CLK _1899_/A vdd gnd DFFPOSX1
X_1532_ _1783_/Y _987_/A _1533_/C vdd gnd NAND2X1
XFILL_0__1806_ gnd vdd FILL
X_1601_ _1617_/C _1601_/B _1626_/B vdd gnd NAND2X1
X_1463_ _1519_/B _1467_/A _1464_/C vdd gnd NAND2X1
X_1394_ _1464_/B _1404_/B _1404_/C _1416_/C vdd gnd AOI21X1
XFILL_0__1453_ gnd vdd FILL
X_1377_ _1377_/A _1377_/B _1420_/A vdd gnd AND2X2
X_1515_ _1557_/B _1515_/B _1515_/C _1537_/A vdd gnd NAND3X1
X_1446_ _1489_/B _1511_/B vdd gnd INVX1
X_1093_ _1193_/A _1192_/B _1193_/B _1104_/C vdd gnd OAI21X1
X_1231_ _1231_/A _1232_/B vdd gnd INVX1
XBUFX2_insert5 _1665_/Q _1114_/A vdd gnd BUFX2
X_1300_ _1304_/A _1304_/B _1303_/C _1402_/B vdd gnd OAI21X1
XFILL_0__1298_ gnd vdd FILL
X_1429_ _1429_/A _1429_/B _1487_/B vdd gnd NOR2X1
X_1162_ _1297_/B _1297_/A _1246_/C _1176_/A vdd gnd NAND3X1
X_942_ _953_/A _942_/B _942_/C _949_/B vdd gnd OAI21X1
XFILL75450x54150 gnd vdd FILL
X_1780_ _1780_/A _1802_/B _1789_/B _1786_/A vdd gnd OAI21X1
X_1214_ _1238_/A _1580_/B vdd gnd INVX1
X_1145_ _1164_/B _1164_/A _1164_/C _1297_/A vdd gnd NAND3X1
XFILL76350x39750 gnd vdd FILL
X_1076_ _1267_/C _994_/B _1083_/C vdd gnd AND2X2
XCLKBUF1_insert12 clk _1691_/CLK vdd gnd CLKBUF1
X_1832_ _1848_/A _983_/A _1832_/C _1834_/B vdd gnd AOI21X1
X_1901_ _1901_/A ACC_o[7] vdd gnd BUFX2
X_1694_ _1694_/A _1848_/C ABCmd_i[4] _1716_/B vdd gnd OAI21X1
X_1763_ _1763_/A _1763_/B _1787_/A _1764_/B vdd gnd OAI21X1
XFILL_0__1899_ gnd vdd FILL
X_1128_ _992_/A _995_/B _1152_/B vdd gnd AND2X2
X_1059_ _1813_/A _1548_/A vdd gnd INVX2
XFILL_0__1135_ gnd vdd FILL
XFILL76350x14550 gnd vdd FILL
X_1746_ _1802_/C _1746_/Y vdd gnd INVX1
X_1815_ _1848_/A _980_/A _1848_/C _1816_/C vdd gnd OAI21X1
X_1677_ _1677_/D _1680_/CLK _1898_/A vdd gnd DFFPOSX1
XFILL_0__938_ gnd vdd FILL
XFILL_0__1736_ gnd vdd FILL
X_1531_ _1580_/C _1531_/B _1533_/B vdd gnd NAND2X1
X_1600_ _1600_/A _1600_/B _1600_/C _1617_/C vdd gnd NAND3X1
X_1393_ _1466_/A _1396_/B _1396_/C _1404_/B vdd gnd NAND3X1
X_1462_ _1462_/A _1521_/C _1462_/C _1519_/B vdd gnd NAND3X1
X_1729_ _1759_/A _1729_/B _1729_/C _1747_/A vdd gnd AOI21X1
XFILL76050x36150 gnd vdd FILL
XFILL_0__1383_ gnd vdd FILL
X_1376_ _1453_/B _1420_/C _1453_/A _1465_/A vdd gnd OAI21X1
X_1514_ _1514_/A _1514_/B _1514_/C _1522_/A vdd gnd NAND3X1
X_1445_ _1449_/A _1449_/B _1456_/A _1489_/B vdd gnd NAND3X1
X_1230_ _1530_/A _1478_/B vdd gnd INVX1
XBUFX2_insert6 _1665_/Q _995_/A vdd gnd BUFX2
X_1161_ _1161_/A _1161_/B _1297_/B vdd gnd NAND2X1
X_1092_ _1105_/B _1105_/C _1105_/A _1197_/B vdd gnd NAND3X1
X_941_ _941_/A _949_/A vdd gnd INVX4
X_1428_ _1429_/B _1429_/A _1430_/B vdd gnd AND2X2
X_1359_ _1829_/A _1439_/B _1813_/A _1500_/B _1424_/B vdd gnd AOI22X1
XFILL_0__1220_ gnd vdd FILL
X_1213_ _1234_/B _1234_/C _1234_/A _1238_/A vdd gnd NAND3X1
XFILL_0__1151_ gnd vdd FILL
X_1075_ _1085_/A _1152_/D vdd gnd INVX1
XFILL_0__1418_ gnd vdd FILL
X_1144_ _1287_/A _1287_/C _1258_/B _1164_/B vdd gnd NAND3X1
X_1693_ ABCmd_i[3] _1848_/C vdd gnd INVX4
X_1762_ _1881_/A _1763_/B _1763_/A _1787_/A vdd gnd OAI21X1
X_1831_ _1848_/A _983_/A _1848_/C _1832_/C vdd gnd OAI21X1
XCLKBUF1_insert13 clk _1680_/CLK vdd gnd CLKBUF1
X_1900_ _1900_/A ACC_o[6] vdd gnd BUFX2
XFILL_0__1065_ gnd vdd FILL
X_1127_ _1250_/A _1133_/A vdd gnd INVX1
X_1058_ _1274_/A _1061_/A vdd gnd INVX1
XFILL_0__954_ gnd vdd FILL
XFILL76350x150 gnd vdd FILL
X_1745_ _1745_/A _1764_/C _1802_/C vdd gnd NAND2X1
X_1814_ _1814_/A _1814_/B _1814_/C _1818_/A vdd gnd OAI21X1
XFILL_0__1821_ gnd vdd FILL
X_1676_ _1676_/D _1680_/CLK _1897_/A vdd gnd DFFPOSX1
X_1530_ _1530_/A _1530_/B _1531_/B vdd gnd NAND2X1
X_1392_ _1392_/A _1392_/B _1465_/C _1396_/B vdd gnd OAI21X1
X_1461_ _1461_/A _1461_/B _1461_/C _1462_/C vdd gnd OAI21X1
X_1728_ _1759_/A _1729_/B _1848_/C _1729_/C vdd gnd OAI21X1
X_1659_ _1813_/A _1659_/B _1660_/C vdd gnd NAND2X1
XFILL75450x39750 gnd vdd FILL
X_1513_ _1516_/A _1555_/C _1515_/B _1514_/B vdd gnd OAI21X1
X_1444_ _1449_/A _1449_/B _1456_/A _1489_/C vdd gnd AOI21X1
X_1375_ _1385_/A _1449_/B _1378_/C _1453_/B vdd gnd AOI21X1
XBUFX2_insert7 _1665_/Q _1711_/A vdd gnd BUFX2
XFILL_0__1503_ gnd vdd FILL
X_1091_ _1146_/A _1146_/C _1111_/A _1105_/B vdd gnd NAND3X1
X_1160_ _1166_/A _1165_/B _1245_/A _1161_/A vdd gnd NAND3X1
XFILL_0__1434_ gnd vdd FILL
XFILL75450x14550 gnd vdd FILL
X_1358_ _1363_/C _1364_/C _1424_/C vdd gnd NAND2X1
X_1427_ _1427_/A _1487_/C _1427_/C _1454_/A vdd gnd NAND3X1
X_1289_ _1289_/A _1289_/B _1374_/A _1386_/B vdd gnd AOI21X1
X_940_ LoadA_i _960_/A vdd gnd INVX1
XFILL_0__1081_ gnd vdd FILL
X_1212_ _1212_/A _1212_/B _1212_/C _1234_/A vdd gnd OAI21X1
X_1074_ _980_/A _997_/B _1085_/A vdd gnd NAND2X1
X_1143_ _1143_/A _1143_/B _1287_/A vdd gnd NAND2X1
XFILL_0__1348_ gnd vdd FILL
XFILL_0__1279_ gnd vdd FILL
X_1692_ _970_/A _1694_/A vdd gnd INVX1
X_1761_ _1801_/A _1801_/B _1787_/B vdd gnd NAND2X1
XCLKBUF1_insert14 clk _1682_/CLK vdd gnd CLKBUF1
X_1830_ _1868_/B _1882_/C _1830_/C _1830_/D _1834_/A vdd gnd OAI22X1
X_1126_ _980_/A _994_/B _1250_/A vdd gnd NAND2X1
X_1057_ _1057_/A _1432_/A _1125_/A vdd gnd NAND2X1
XFILL76650x68550 gnd vdd FILL
XFILL_0__1751_ gnd vdd FILL
X_1744_ _1748_/B _1744_/B _1745_/A vdd gnd NAND2X1
X_1675_ _1675_/D _1682_/CLK _1896_/A vdd gnd DFFPOSX1
X_1813_ _1813_/A _1813_/B _1868_/B _1814_/A vdd gnd OAI21X1
XFILL_0__1116_ gnd vdd FILL
X_1109_ _1307_/A _1244_/A vdd gnd INVX1
XFILL76650x43350 gnd vdd FILL
X_1727_ _1727_/A _1727_/B _1727_/C _1747_/B vdd gnd OAI21X1
X_1658_ _978_/A _1664_/B _1658_/C _1685_/D vdd gnd OAI21X1
XFILL_0__1596_ gnd vdd FILL
X_1391_ _1465_/A _1465_/B _1391_/C _1396_/C vdd gnd NAND3X1
X_1460_ _1520_/B _1520_/A _1520_/C _1521_/C vdd gnd NAND3X1
X_1589_ _1589_/A _1621_/C _1640_/C vdd gnd NAND2X1
X_1512_ _1557_/B _1555_/C vdd gnd INVX1
X_1443_ _1450_/B _1450_/A _1456_/A vdd gnd NAND2X1
X_1374_ _1374_/A _1374_/B _1374_/C _1378_/C vdd gnd OAI21X1
XBUFX2_insert8 _934_/Y _1659_/B vdd gnd BUFX2
X_1090_ _1090_/A _1090_/B _1146_/A vdd gnd NAND2X1
X_1357_ _1829_/A _990_/A _1364_/C vdd gnd AND2X2
XFILL_0__1364_ gnd vdd FILL
X_1426_ _1429_/B _1429_/A _1427_/C vdd gnd OR2X2
X_1288_ _1288_/A _1288_/B _1353_/B _1374_/C _1382_/A vdd gnd AOI22X1
X_999_ _999_/A _999_/B _999_/C _999_/Y vdd gnd OAI21X1
X_1211_ _1232_/C _1232_/A _1231_/A _1234_/C vdd gnd OAI21X1
X_1073_ _1088_/B _1088_/A _1088_/C _1111_/C vdd gnd AOI21X1
X_1142_ _1142_/A _1142_/B _1142_/C _1287_/C vdd gnd NAND3X1
X_1409_ _1746_/Y _987_/A _1411_/C vdd gnd NAND2X1
X_1691_ _963_/Y vdd _962_/Y _1691_/CLK _936_/A vdd gnd DFFSR
XCLKBUF1_insert15 clk _1687_/CLK vdd gnd CLKBUF1
X_1760_ _1760_/A _1760_/B _1763_/A _1801_/A vdd gnd MUX2X1
XFILL_0__1201_ gnd vdd FILL
X_1889_ _1891_/A _1891_/B _1890_/C vdd gnd NAND2X1
X_1125_ _1125_/A _1125_/B _1141_/B _1141_/A _1258_/C vdd gnd AOI22X1
X_1056_ _1274_/A _1829_/A _1432_/A vdd gnd AND2X2
X_1743_ _1747_/B _1747_/A _1764_/A _1744_/B vdd gnd OAI21X1
X_1812_ _1845_/A _980_/A _1812_/C _1845_/D _1814_/B vdd gnd AOI22X1
X_1674_ _1674_/D _1688_/CLK _1895_/A vdd gnd DFFPOSX1
XFILL_0__1879_ gnd vdd FILL
XFILL_0__1046_ gnd vdd FILL
X_1039_ _991_/B _1249_/A _1039_/C _1040_/A vdd gnd OAI21X1
X_1108_ _1315_/A _1315_/B _1218_/C _1318_/B vdd gnd NAND3X1
XFILL_0__1802_ gnd vdd FILL
X_1390_ _1396_/A _1466_/A vdd gnd INVX1
X_1657_ _1794_/A _1664_/B _1658_/C vdd gnd NAND2X1
X_1726_ _997_/B _1726_/B _1868_/B _1727_/B vdd gnd OAI21X1
X_1588_ _1590_/A _1590_/D _1621_/C vdd gnd NOR2X1
X_1511_ _1511_/A _1511_/B _1511_/C _1515_/B vdd gnd OAI21X1
X_1442_ _1493_/D _1442_/B _1493_/C _1450_/B vdd gnd OAI21X1
XFILL_0__1716_ gnd vdd FILL
X_1709_ _1709_/A _1709_/B _1740_/A _1741_/A vdd gnd OAI21X1
XFILL_0__1647_ gnd vdd FILL
X_1373_ _1373_/A _1373_/B _1374_/B vdd gnd NOR2X1
XBUFX2_insert9 _934_/Y _1662_/B vdd gnd BUFX2
X_1356_ _1813_/A _1500_/B _1363_/C vdd gnd AND2X2
XFILL_0__1294_ gnd vdd FILL
X_1425_ _1429_/A _1429_/B _1487_/C vdd gnd NAND2X1
X_1287_ _1287_/A _1287_/B _1287_/C _1339_/C vdd gnd OAI21X1
X_998_ _998_/A _998_/B _999_/B vdd gnd AND2X2
X_1210_ _1210_/A _1210_/B _1210_/C _1232_/A vdd gnd AOI21X1
X_1141_ _1141_/A _1141_/B _1141_/C _1258_/B vdd gnd NAND3X1
X_1072_ _1140_/A _1112_/B _1125_/A _1088_/A vdd gnd NAND3X1
X_1408_ _1410_/A _1410_/B _1411_/B vdd gnd AND2X2
XFILL76650x28950 gnd vdd FILL
X_1339_ _1339_/A _1339_/B _1339_/C _1340_/B vdd gnd AOI21X1
X_1690_ _963_/Y vdd _957_/Y _1691_/CLK _953_/A vdd gnd DFFSR
XCLKBUF1_insert16 clk _1688_/CLK vdd gnd CLKBUF1
XFILL_0__1131_ gnd vdd FILL
XFILL_0__1329_ gnd vdd FILL
XFILL_0__1895_ gnd vdd FILL
X_1888_ _1888_/A _1888_/B _1888_/C _1891_/B vdd gnd NAND3X1
X_1055_ _1055_/A _1055_/B _1055_/C _1089_/A vdd gnd OAI21X1
X_1124_ _1271_/A _1277_/B _1277_/C _1141_/A vdd gnd NAND3X1
X_1742_ _1881_/A _1747_/A _1747_/B _1764_/A vdd gnd OAI21X1
X_1673_ _1673_/D _1688_/CLK _988_/A vdd gnd DFFPOSX1
X_1811_ _1813_/A _1813_/B _1812_/C vdd gnd NAND2X1
X_1038_ _994_/B _1249_/A vdd gnd INVX1
X_1107_ _1196_/A _1196_/B _1197_/A _1315_/B vdd gnd OAI21X1
XFILL_0__1732_ gnd vdd FILL
XFILL_0__934_ gnd vdd FILL
X_1656_ _975_/A _1662_/B _1656_/C _1684_/D vdd gnd OAI21X1
X_1725_ ABCmd_i[0] _1725_/B _1726_/B vdd gnd NOR2X1
X_1587_ _1587_/A _1587_/B _1587_/C _1619_/A vdd gnd AOI21X1
XFILL76350x25350 gnd vdd FILL
X_1708_ _997_/B ABCmd_i[5] _1740_/A vdd gnd NAND2X1
XFILL_0__1577_ gnd vdd FILL
X_1372_ _1386_/C _1385_/C _1420_/C vdd gnd NOR2X1
X_1510_ _1515_/C _1557_/B _1516_/C _1514_/C vdd gnd NAND3X1
X_1441_ _1441_/A _1441_/B _1441_/C _1450_/A vdd gnd NAND3X1
X_1639_ _1639_/A _1639_/B _1639_/C _1641_/B vdd gnd AOI21X1
XFILL75750x7350 gnd vdd FILL
XFILL_0__1500_ gnd vdd FILL
X_1424_ _1424_/A _1424_/B _1424_/C _1429_/B vdd gnd OAI21X1
X_1355_ _1424_/A _1368_/A vdd gnd INVX1
X_1286_ _1339_/A _1339_/B _1382_/C _1299_/A vdd gnd NAND3X1
X_997_ _997_/A _997_/B _999_/A vdd gnd NAND2X1
X_1071_ _1112_/A _1140_/C _1140_/B _1088_/B vdd gnd OAI21X1
X_1140_ _1140_/A _1140_/B _1140_/C _1141_/C vdd gnd AOI21X1
XFILL_0__1414_ gnd vdd FILL
X_1407_ _1407_/A _1407_/B _1407_/C _1413_/C vdd gnd OAI21X1
X_1338_ _1338_/A _1338_/B _1338_/C _1396_/A vdd gnd OAI21X1
XFILL76050x150 gnd vdd FILL
X_1269_ _1269_/A _1269_/B _1344_/C _1288_/B vdd gnd NAND3X1
X_1887_ _1887_/A _1888_/B vdd gnd INVX1
X_1054_ _1193_/C _1192_/C _1192_/A _1105_/C vdd gnd AOI21X1
X_1123_ _1277_/A _1271_/C _1271_/B _1141_/B vdd gnd OAI21X1
XFILL_0__1061_ gnd vdd FILL
XFILL_0__1259_ gnd vdd FILL
XFILL_0__950_ gnd vdd FILL
X_1741_ _1741_/A _1741_/B _1741_/C _1741_/D _1748_/B vdd gnd AOI22X1
X_1810_ _1843_/A _980_/A _1813_/B vdd gnd AND2X2
X_1672_ _987_/Y _1688_/CLK _986_/A vdd gnd DFFPOSX1
X_1037_ _993_/A _1152_/A _1040_/C vdd gnd NAND2X1
X_1106_ _1307_/A _1106_/B _1197_/A vdd gnd NAND2X1
XFILL_0__1662_ gnd vdd FILL
X_1655_ _995_/B _1662_/B _1656_/C vdd gnd NAND2X1
X_1724_ _1729_/B _1725_/B vdd gnd INVX1
X_1586_ _1899_/A _1615_/A vdd gnd INVX1
XFILL_0__1027_ gnd vdd FILL
XFILL_0__1593_ gnd vdd FILL
X_1371_ _1449_/B _1385_/A _1386_/C vdd gnd NAND2X1
X_1440_ _1493_/D _1441_/B vdd gnd INVX1
X_1707_ _1868_/B _1739_/B _1709_/B vdd gnd NAND2X1
X_1638_ _1901_/A _1648_/A vdd gnd INVX1
X_1569_ _1627_/A _1627_/B _1626_/A _1576_/B vdd gnd AOI21X1
XFILL_0__1430_ gnd vdd FILL
XFILL76650x3750 gnd vdd FILL
X_1285_ _1374_/C _1353_/B _1353_/A _1339_/B vdd gnd NAND3X1
XFILL76350x7350 gnd vdd FILL
X_1423_ _1499_/A _1621_/B _1429_/A vdd gnd NOR2X1
X_1354_ _1794_/A _980_/A _1424_/A vdd gnd NAND2X1
X_996_ _998_/A _998_/B _999_/C vdd gnd OR2X2
X_1406_ _1564_/B _1406_/B ABCmd_i[7] _1407_/B vdd gnd OAI21X1
X_1070_ _1070_/A _1070_/B _1070_/C _1088_/C vdd gnd AOI21X1
X_1337_ _1337_/A _1337_/B _1401_/A _1404_/C vdd gnd OAI21X1
XFILL_0__1275_ gnd vdd FILL
XFILL_0__1344_ gnd vdd FILL
X_1268_ _1344_/B _1269_/B vdd gnd INVX1
X_1199_ _1244_/A _1244_/B _1307_/C _1201_/B vdd gnd NAND3X1
X_979_ ABCmd_i[5] _981_/A vdd gnd INVX1
X_1053_ _993_/Y _1236_/B _1316_/A _1218_/C vdd gnd OAI21X1
X_1122_ _1142_/C _1142_/B _1142_/A _1287_/B vdd gnd AOI21X1
X_1886_ _1886_/A _1887_/A _1886_/C _1891_/A vdd gnd NAND3X1
XFILL_0__1189_ gnd vdd FILL
X_1740_ _1740_/A _1740_/B _1740_/C _1741_/C vdd gnd NAND3X1
X_1671_ _984_/Y _1687_/CLK _983_/A vdd gnd DFFPOSX1
XFILL_0__1112_ gnd vdd FILL
X_1105_ _1105_/A _1105_/B _1105_/C _1196_/A vdd gnd AOI21X1
X_1869_ _1869_/A _1869_/B _1869_/C _1876_/A vdd gnd OAI21X1
X_1036_ _1131_/A _994_/B _1152_/A vdd gnd AND2X2
X_1654_ _972_/A _956_/C _1654_/C _1683_/D vdd gnd OAI21X1
X_1723_ _1845_/A _1729_/B _1723_/C _1845_/D _1727_/A vdd gnd AOI22X1
X_1585_ _1585_/A _949_/A _1585_/C _1585_/D _1677_/D vdd gnd AOI22X1
X_1019_ _1114_/A _1813_/A _1057_/A vdd gnd AND2X2
XFILL_0__1713_ gnd vdd FILL
X_1370_ _1370_/A _1370_/B _1370_/C _1449_/B vdd gnd NAND3X1
X_1706_ ABCmd_i[0] _1736_/B _1868_/A _1739_/B vdd gnd OAI21X1
X_1637_ _1637_/A _949_/A _1637_/C _1637_/D _1679_/D vdd gnd AOI22X1
X_1568_ _1573_/A _1573_/B _1568_/C _1573_/C _1627_/A vdd gnd AOI22X1
X_1499_ _1499_/A _1590_/D _1539_/B _1509_/C vdd gnd OAI21X1
XFILL76650x54150 gnd vdd FILL
XFILL_0__1360_ gnd vdd FILL
XFILL_0__1627_ gnd vdd FILL
X_1422_ _1487_/A _1427_/A vdd gnd INVX1
X_1353_ _1353_/A _1353_/B _1386_/A _1385_/C vdd gnd AOI21X1
X_1284_ _1352_/A _1352_/B _1353_/B vdd gnd NAND2X1
XFILL_0__1558_ gnd vdd FILL
XBUFX2_insert30 ABCmd_i[2] _1759_/A vdd gnd BUFX2
X_995_ _995_/A _995_/B _998_/B vdd gnd NAND2X1
X_1405_ _1416_/B _1405_/B _1564_/B vdd gnd NAND2X1
X_1198_ _1316_/A _1316_/B _1198_/C _1198_/D _1241_/A vdd gnd AOI22X1
X_1267_ _1813_/A _990_/A _1267_/C _1794_/A _1344_/B vdd gnd AOI22X1
X_1336_ _1336_/A _1336_/B _1336_/C _1337_/B vdd gnd AOI21X1
X_978_ _978_/A _983_/B _978_/C _978_/Y vdd gnd OAI21X1
X_1052_ _1052_/A _1052_/B _1052_/C _1236_/B vdd gnd AOI21X1
X_1121_ _1277_/A _1271_/C _1277_/B _1142_/C vdd gnd OAI21X1
X_1885_ _1885_/A _1885_/B _1887_/A vdd gnd NOR2X1
X_1319_ _1632_/C _1632_/B _1631_/B _1642_/C vdd gnd OAI21X1
X_1670_ _981_/Y _1687_/CLK _980_/A vdd gnd DFFPOSX1
XFILL_0__1875_ gnd vdd FILL
X_1035_ _1044_/A _1040_/B vdd gnd INVX1
X_1104_ _1104_/A _1104_/B _1104_/C _1196_/B vdd gnd AOI21X1
XFILL_0__1042_ gnd vdd FILL
X_1799_ _1799_/A _1799_/B _1808_/A _1805_/A vdd gnd OAI21X1
X_1868_ _1868_/A _1868_/B _1873_/A vdd gnd NOR2X1
X_1653_ _994_/B _956_/C _1654_/C vdd gnd NAND2X1
X_1722_ _997_/B _1729_/B _1843_/A _1723_/C vdd gnd NAND3X1
X_1584_ _1584_/A _937_/A _949_/A _1585_/D vdd gnd AOI21X1
X_1018_ _1187_/A _1186_/A _1187_/C _1048_/C vdd gnd OAI21X1
X_1705_ _989_/A _1868_/A vdd gnd INVX1
X_1636_ _1636_/A _937_/A _949_/A _1637_/D vdd gnd AOI21X1
XFILL_0__1643_ gnd vdd FILL
X_1567_ _1567_/A _1567_/B _1573_/B vdd gnd NAND2X1
X_1498_ _1539_/C _1498_/B _1539_/B vdd gnd NAND2X1
XFILL_0__1290_ gnd vdd FILL
XFILL_0__1488_ gnd vdd FILL
X_1421_ _995_/B _986_/A _1487_/A vdd gnd NAND2X1
X_1283_ _1373_/A _1373_/B _1374_/C vdd gnd NAND2X1
X_1352_ _1352_/A _1352_/B _1386_/A vdd gnd NOR2X1
XBUFX2_insert31 ABCmd_i[2] _1849_/A vdd gnd BUFX2
XBUFX2_insert20 _953_/Y _987_/B vdd gnd BUFX2
X_1619_ _1619_/A _1619_/B _1619_/C _1620_/A vdd gnd OAI21X1
X_994_ _994_/A _994_/B _998_/A vdd gnd NAND2X1
X_1335_ _1335_/A _960_/C _1606_/A _1407_/C vdd gnd OAI21X1
X_1197_ _1197_/A _1197_/B _1197_/C _1198_/D vdd gnd NAND3X1
X_1404_ _1464_/B _1404_/B _1404_/C _1416_/B vdd gnd NAND3X1
X_1266_ _1266_/A _1266_/B _1344_/C vdd gnd NAND2X1
X_977_ _977_/A _983_/B _978_/C vdd gnd NAND2X1
XFILL_0__1891_ gnd vdd FILL
XFILL_0__1325_ gnd vdd FILL
X_1884_ _1884_/A _1884_/B _1885_/B vdd gnd NOR2X1
X_1051_ _1052_/B _1052_/A _1052_/C _1316_/A vdd gnd NAND3X1
X_1318_ _1318_/A _1318_/B _1318_/C _1632_/B vdd gnd AOI21X1
X_1120_ _1120_/A _1120_/B _1271_/C vdd gnd NOR2X1
X_1249_ _1249_/A _1621_/B _1255_/A vdd gnd NOR2X1
XFILL75750x54150 gnd vdd FILL
X_1034_ _989_/A _980_/A _1044_/A vdd gnd NAND2X1
X_1103_ _1197_/B _1197_/C _1196_/C _1315_/A vdd gnd NAND3X1
X_1798_ _1881_/A _1799_/B _1799_/A _1808_/A vdd gnd OAI21X1
XFILL_0__930_ gnd vdd FILL
X_1867_ _1867_/A _1867_/B ABCmd_i[6] _1878_/B vdd gnd OAI21X1
XFILL76650x39750 gnd vdd FILL
X_1721_ ABCmd_i[5] _994_/B _1727_/C vdd gnd NAND2X1
X_1652_ _969_/A _1659_/B _1652_/C _1682_/D vdd gnd OAI21X1
X_1017_ _1212_/C _1212_/B _1215_/A _1052_/C vdd gnd OAI21X1
X_1583_ _987_/A _1583_/B _1583_/C _1584_/A vdd gnd OAI21X1
XFILL76050x10950 gnd vdd FILL
XFILL76650x14550 gnd vdd FILL
XFILL_0_BUFX2_insert0 gnd vdd FILL
X_1704_ _1711_/A _1736_/B vdd gnd INVX1
XFILL_0__1007_ gnd vdd FILL
X_1635_ _987_/A _1635_/B _1635_/C _1636_/A vdd gnd OAI21X1
X_1566_ _1566_/A _1568_/C _1566_/C _1627_/B vdd gnd NAND3X1
XFILL_0__1573_ gnd vdd FILL
X_1497_ _986_/A _1590_/D vdd gnd INVX2
X_1420_ _1420_/A _1420_/B _1420_/C _1461_/C vdd gnd AOI21X1
X_1351_ _1377_/B _1377_/A _1453_/A vdd gnd NAND2X1
X_1282_ _1288_/A _1288_/B _1353_/A vdd gnd AND2X2
X_1618_ _1629_/A _1639_/B vdd gnd INVX1
X_1549_ _1552_/B _1552_/C _1593_/B vdd gnd NAND2X1
XBUFX2_insert10 _934_/Y _956_/C vdd gnd BUFX2
XBUFX2_insert32 ABCmd_i[2] _1848_/A vdd gnd BUFX2
XFILL_0__1410_ gnd vdd FILL
XFILL76350x36150 gnd vdd FILL
X_993_ _993_/A _993_/B _993_/Y vdd gnd NAND2X1
XBUFX2_insert21 _1669_/Q _992_/A vdd gnd BUFX2
XFILL_0__1341_ gnd vdd FILL
X_1334_ _953_/A _949_/A ABCmd_i[7] _1606_/A vdd gnd OAI21X1
XFILL_0__1608_ gnd vdd FILL
X_1196_ _1196_/A _1196_/B _1196_/C _1198_/C vdd gnd OAI21X1
X_1403_ _1403_/A _1403_/B _1403_/C _1405_/B vdd gnd NAND3X1
X_1265_ _1344_/A _1269_/A vdd gnd INVX1
X_976_ ABCmd_i[4] _978_/A vdd gnd INVX1
X_1883_ _1883_/A _1883_/B _1884_/B vdd gnd NAND2X1
XFILL_0__1186_ gnd vdd FILL
X_1050_ _1192_/A _1192_/B _1193_/A _1052_/A vdd gnd OAI21X1
XFILL_0__1255_ gnd vdd FILL
X_1317_ _1318_/B _1318_/C _1318_/A _1631_/B vdd gnd NAND3X1
X_1179_ _1643_/A _1642_/B vdd gnd INVX1
X_1248_ _1338_/A _1253_/A vdd gnd INVX1
X_959_ _959_/A _959_/B _959_/C _959_/D _961_/A vdd gnd AOI22X1
X_1102_ _1106_/B _1307_/A _1196_/C vdd gnd AND2X2
X_1797_ _1849_/A _977_/A _1797_/C _1799_/B vdd gnd AOI21X1
XFILL_0_BUFX2_insert31 gnd vdd FILL
X_1866_ _1888_/A _1888_/C _1878_/A vdd gnd NAND2X1
X_1033_ _1047_/B _1047_/A _1047_/C _1193_/C vdd gnd NAND3X1
X_1720_ _1720_/A _1720_/B _1720_/C _1733_/B vdd gnd OAI21X1
X_1651_ _997_/B _1659_/B _1652_/C vdd gnd NAND2X1
X_1016_ _1016_/A _1016_/B _999_/Y _1212_/B vdd gnd AOI21X1
X_1582_ _1859_/B _987_/A _1583_/C vdd gnd NAND2X1
XFILL_0__1856_ gnd vdd FILL
XFILL_0__989_ gnd vdd FILL
XFILL_0__1023_ gnd vdd FILL
X_1849_ _1849_/A _986_/A _1849_/C _1880_/A vdd gnd AOI21X1
X_1703_ ABCmd_i[5] _1868_/B vdd gnd INVX2
X_1634_ _1867_/B _987_/A _1635_/C vdd gnd NAND2X1
X_1565_ _1572_/B _1572_/A _1568_/C vdd gnd NOR2X1
X_1496_ _1496_/A _1539_/C _1498_/B _1509_/B vdd gnd NAND3X1
X_1350_ _1418_/B _1350_/B _1418_/A _1377_/B vdd gnd OAI21X1
X_1281_ _1289_/B _1374_/A _1289_/A _1339_/A vdd gnd NAND3X1
X_1479_ ABCmd_i[7] _1766_/Y _1480_/A vdd gnd NOR2X1
XFILL_0__1624_ gnd vdd FILL
X_1617_ _1617_/A _1626_/B _1617_/C _1629_/A vdd gnd OAI21X1
X_1548_ _1548_/A _1590_/D _1548_/C _1587_/C _1552_/B vdd gnd OAI22X1
XBUFX2_insert11 _934_/Y _1664_/B vdd gnd BUFX2
XBUFX2_insert22 _1669_/Q _977_/A vdd gnd BUFX2
X_992_ _992_/A _997_/B _993_/A vdd gnd AND2X2
XFILL75750x39750 gnd vdd FILL
X_1333_ _1879_/C _1335_/A vdd gnd INVX1
X_1195_ _1236_/C _1237_/B _1316_/A _1316_/B vdd gnd NAND3X1
XFILL_0__1538_ gnd vdd FILL
XFILL_0__1469_ gnd vdd FILL
X_1402_ _1402_/A _1402_/B _1402_/C _1403_/C vdd gnd AOI21X1
XFILL_0__1271_ gnd vdd FILL
X_1264_ _1344_/A _1264_/B _1264_/C _1288_/A vdd gnd NAND3X1
X_975_ _975_/A _984_/B _975_/C _975_/Y vdd gnd OAI21X1
X_1882_ _1883_/B _1883_/A _1882_/C _1885_/A vdd gnd AOI21X1
XFILL75750x14550 gnd vdd FILL
X_1316_ _1316_/A _1316_/B _1316_/C _1318_/A vdd gnd NAND3X1
X_1178_ _1313_/C _1313_/B _1318_/B _1643_/A vdd gnd AOI21X1
X_1247_ _986_/A _997_/B _1338_/A vdd gnd NAND2X1
X_958_ _972_/B _959_/A vdd gnd INVX1
X_1796_ _1849_/A _977_/A _1848_/C _1797_/C vdd gnd OAI21X1
XFILL_0__1872_ gnd vdd FILL
X_1865_ _1865_/A _1865_/B _1874_/A _1888_/C vdd gnd OAI21X1
X_1032_ _1070_/A _1055_/B _1055_/C _1047_/B vdd gnd NAND3X1
X_1101_ _1101_/A _1101_/B _1106_/B vdd gnd OR2X2
XFILL_0__1306_ gnd vdd FILL
X_1650_ _966_/A _1659_/B _1650_/C _1681_/D vdd gnd OAI21X1
XFILL_0__1786_ gnd vdd FILL
X_1015_ _1039_/C _1232_/C _1189_/B _1212_/C vdd gnd OAI21X1
X_1581_ _1581_/A _1581_/B _1583_/B vdd gnd NAND2X1
XFILL75450x36150 gnd vdd FILL
X_1779_ _1781_/B _1789_/B vdd gnd INVX1
X_1848_ _1848_/A _986_/A _1848_/C _1849_/C vdd gnd OAI21X1
XFILL76350x64950 gnd vdd FILL
X_1702_ _1711_/A _1702_/B _1845_/D _1702_/D _1709_/A vdd gnd AOI22X1
X_1633_ _1633_/A _1633_/B _1635_/B vdd gnd NAND2X1
X_1564_ _1564_/A _1564_/B _1566_/C vdd gnd NOR2X1
X_1495_ _1495_/A _1495_/B _1498_/B vdd gnd OR2X2
X_1616_ _1900_/A _1637_/A vdd gnd INVX1
X_1547_ _1621_/B _1547_/B _1587_/C vdd gnd NOR2X1
X_1280_ _1352_/A _1373_/B _1289_/B vdd gnd NAND2X1
XFILL_0__1554_ gnd vdd FILL
X_1478_ _1478_/A _1478_/B ABCmd_i[7] _1481_/A vdd gnd OAI21X1
X_991_ _991_/A _991_/B _993_/B vdd gnd NOR2X1
XBUFX2_insert23 _1669_/Q _1500_/B vdd gnd BUFX2
X_1332_ _1895_/A _1413_/A vdd gnd INVX1
X_1194_ _1215_/D _1215_/C _1194_/C _1237_/B vdd gnd NAND3X1
X_1401_ _1401_/A _1402_/C vdd gnd INVX1
X_1263_ _1364_/B _1499_/A _1266_/B _1264_/C vdd gnd OAI21X1
XFILL_0__1399_ gnd vdd FILL
X_974_ _974_/A _984_/B _975_/C vdd gnd NAND2X1
X_1881_ _1881_/A _1881_/B _1883_/B vdd gnd NAND2X1
X_1315_ _1315_/A _1315_/B _1316_/C vdd gnd NAND2X1
X_1246_ _1246_/A _1246_/B _1246_/C _1336_/C vdd gnd OAI21X1
X_1177_ _1307_/A _1244_/B _1307_/C _1313_/B vdd gnd NAND3X1
X_957_ _957_/A _957_/B _957_/Y vdd gnd OR2X2
X_1795_ _1795_/A _1795_/B _1795_/C _1799_/A vdd gnd OAI21X1
X_1864_ _1869_/A _1869_/B _1864_/C _1888_/A vdd gnd NAND3X1
XFILL_0__1236_ gnd vdd FILL
X_1031_ _1055_/A _1070_/C _1070_/B _1047_/A vdd gnd OAI21X1
X_1100_ _1101_/B _1101_/A _1307_/A vdd gnd NAND2X1
XFILL_0_BUFX2_insert11 gnd vdd FILL
X_1229_ _1477_/C _1477_/B _1477_/A _1530_/A vdd gnd NAND3X1
X_1580_ _1580_/A _1580_/B _1580_/C _1581_/A vdd gnd OAI21X1
X_1778_ _1778_/A _1778_/B _1788_/A _1781_/B vdd gnd OAI21X1
X_1847_ _1847_/A _1847_/B _1847_/C _1881_/B vdd gnd OAI21X1
X_1014_ _991_/A _1364_/B _1099_/A _1189_/B vdd gnd OAI21X1
XFILL_0_BUFX2_insert3 gnd vdd FILL
X_1701_ _989_/A ABCmd_i[1] _1702_/B vdd gnd NAND2X1
XFILL_0__1837_ gnd vdd FILL
X_1632_ _1632_/A _1632_/B _1632_/C _1633_/B vdd gnd OAI21X1
X_1563_ _1617_/A _1563_/B _1626_/A vdd gnd NAND2X1
X_1494_ _1495_/B _1495_/A _1539_/C vdd gnd NAND2X1
XFILL_0__1484_ gnd vdd FILL
X_1477_ _1477_/A _1477_/B _1477_/C _1478_/A vdd gnd AOI21X1
X_1615_ _1615_/A _949_/A _1615_/C _1615_/D _1678_/D vdd gnd AOI22X1
XBUFX2_insert24 _1669_/Q _1267_/C vdd gnd BUFX2
X_1546_ _1587_/B _1587_/A _1552_/C vdd gnd NAND2X1
X_990_ _990_/A _991_/B vdd gnd INVX2
X_1331_ _988_/Y _941_/A _1331_/C _1673_/D vdd gnd OAI21X1
X_1400_ _1564_/A _1574_/A _1416_/A _1406_/B vdd gnd OAI21X1
X_1529_ _1529_/A _1529_/B _1530_/B vdd gnd NAND2X1
X_1193_ _1193_/A _1193_/B _1193_/C _1215_/D vdd gnd NAND3X1
X_1262_ _1813_/A _1439_/B _1266_/B vdd gnd AND2X2
X_973_ ABCmd_i[3] _975_/A vdd gnd INVX1
X_1880_ _1880_/A _1883_/A vdd gnd INVX1
X_1314_ _1610_/A _1318_/C vdd gnd INVX1
XFILL_0__1321_ gnd vdd FILL
XFILL_0__1519_ gnd vdd FILL
X_1245_ _1245_/A _1245_/B _1402_/A vdd gnd NAND2X1
X_1176_ _1176_/A _1176_/B _1176_/C _1307_/C vdd gnd NAND3X1
X_956_ _959_/B _972_/B _956_/C _959_/D _957_/B vdd gnd OAI22X1
X_1863_ _1863_/A _1863_/B _1863_/Y vdd gnd AND2X2
X_1030_ _1186_/C _1187_/B _1186_/B _1047_/C vdd gnd AOI21X1
XFILL_0__1166_ gnd vdd FILL
X_1794_ _1794_/A _1794_/B _1868_/B _1795_/A vdd gnd OAI21X1
X_1228_ _1228_/A _1228_/B _1228_/C _1477_/B vdd gnd OAI21X1
XFILL_0_BUFX2_insert23 gnd vdd FILL
X_1159_ _1621_/B _1159_/B _1159_/C _1165_/B vdd gnd OAI21X1
X_939_ _959_/C _939_/B LoadB_i _950_/B vdd gnd OAI21X1
X_1777_ _1881_/A _1778_/B _1778_/A _1788_/A vdd gnd OAI21X1
X_1846_ _1884_/A _1846_/B _1868_/B _1847_/A vdd gnd OAI21X1
X_1013_ _1131_/A _997_/B _1099_/A vdd gnd NAND2X1
X_1700_ _1711_/A _1843_/A _1702_/D vdd gnd NAND2X1
XFILL_0__1767_ gnd vdd FILL
XFILL_0__969_ gnd vdd FILL
XFILL_0__1003_ gnd vdd FILL
X_1631_ _1631_/A _1631_/B _1631_/C _1633_/A vdd gnd NAND3X1
X_1562_ _1562_/A _1598_/B _1562_/C _1617_/A vdd gnd NAND3X1
X_1493_ _1493_/A _1505_/C _1493_/C _1493_/D _1495_/A vdd gnd OAI22X1
X_1829_ _1829_/A _1829_/B _1868_/B _1830_/C vdd gnd OAI21X1
XBUFX2_insert25 _1666_/Q _1729_/B vdd gnd BUFX2
X_1476_ _1476_/A _960_/C _1481_/D vdd gnd NOR2X1
X_1614_ _1614_/A _1614_/B _949_/A _1615_/D vdd gnd AOI21X1
X_1545_ _983_/A _1545_/B _1548_/C _1587_/A vdd gnd AOI21X1
XFILL76650x25350 gnd vdd FILL
X_1330_ _941_/A _1330_/B _1331_/C vdd gnd NAND2X1
X_1192_ _1192_/A _1192_/B _1192_/C _1215_/C vdd gnd OAI21X1
XFILL_0__1604_ gnd vdd FILL
X_1261_ _1548_/A _991_/B _1266_/A _1264_/B vdd gnd OAI21X1
X_972_ _972_/A _972_/B _972_/C _972_/Y vdd gnd OAI21X1
X_1528_ _1528_/A _1528_/B _1528_/C _1535_/C vdd gnd OAI21X1
X_1459_ _1521_/A _1459_/B _1459_/C _1467_/A vdd gnd NAND3X1
XFILL_0__1182_ gnd vdd FILL
X_1313_ _1318_/B _1313_/B _1313_/C _1642_/A vdd gnd NAND3X1
XFILL_0__1251_ gnd vdd FILL
X_1244_ _1244_/A _1244_/B _1244_/C _1306_/C vdd gnd AOI21X1
X_1175_ _1175_/A _1175_/B _1175_/C _1244_/B vdd gnd NAND3X1
XFILL_0__1449_ gnd vdd FILL
X_955_ LoadB_i _962_/A _959_/D vdd gnd NOR2X1
X_1793_ _1845_/A _977_/A _1793_/C _1845_/D _1795_/B vdd gnd AOI22X1
X_1227_ _1410_/A _1410_/B _1477_/C vdd gnd NOR2X1
X_1862_ _1879_/B _1879_/C _1863_/A vdd gnd NOR2X1
XFILL_0__1096_ gnd vdd FILL
X_1158_ _1158_/A _1158_/B _1245_/A vdd gnd NAND2X1
X_1089_ _1089_/A _1125_/B _1089_/C _1146_/C vdd gnd NAND3X1
XFILL_0__985_ gnd vdd FILL
X_938_ LoadCmd_i _962_/B _939_/B vdd gnd NOR2X1
X_1776_ _1849_/A _974_/A _1776_/C _1778_/B vdd gnd AOI21X1
X_1845_ _1845_/A _986_/A _1845_/C _1845_/D _1847_/B vdd gnd AOI22X1
XFILL_0__1852_ gnd vdd FILL
XFILL_0__1217_ gnd vdd FILL
X_1012_ _1267_/C _1364_/B vdd gnd INVX2
X_1630_ _1641_/C _1630_/B _1630_/C _1637_/C vdd gnd NAND3X1
X_1561_ _1561_/A _1561_/B _1563_/B vdd gnd NAND2X1
X_1492_ _1548_/A _1621_/B _1495_/B vdd gnd NOR2X1
XFILL_0__1697_ gnd vdd FILL
X_1759_ _1759_/A _1848_/C _1760_/B _1760_/A vdd gnd OAI21X1
X_1828_ _1845_/A _983_/A _1828_/C _1845_/D _1830_/D vdd gnd AOI22X1
XFILL_0__1620_ gnd vdd FILL
X_1613_ _987_/A _1613_/B _953_/A _1614_/B vdd gnd AOI21X1
X_1475_ ABCmd_i[7] _1863_/Y _1476_/A vdd gnd NOR2X1
X_1544_ _1589_/A _1545_/B _1548_/C vdd gnd NOR2X1
XBUFX2_insert26 _1666_/Q _1067_/C vdd gnd BUFX2
XFILL_0__1534_ gnd vdd FILL
X_1191_ _1202_/A _1202_/B _1212_/A _1194_/C vdd gnd AOI21X1
X_1260_ _1267_/C _1794_/A _1266_/A vdd gnd AND2X2
XFILL_0__1465_ gnd vdd FILL
X_1527_ _1527_/A _1527_/B ABCmd_i[7] _1528_/B vdd gnd OAI21X1
X_1389_ _1396_/A _1466_/C _1395_/C _1464_/B vdd gnd NAND3X1
X_1458_ _1461_/A _1461_/B _1520_/C _1459_/B vdd gnd OAI21X1
X_971_ _997_/A _972_/B _972_/C vdd gnd NAND2X1
X_1243_ _1643_/B _1643_/C _1642_/B _1566_/A vdd gnd OAI21X1
X_1312_ _1470_/A _1566_/A _1399_/A vdd gnd NAND2X1
XFILL_0__1379_ gnd vdd FILL
X_1174_ _1244_/C _1307_/B _1244_/A _1313_/C vdd gnd OAI21X1
X_954_ LoadA_i _962_/A _959_/B vdd gnd NOR2X1
X_1792_ _1794_/A _1794_/B _1793_/C vdd gnd NAND2X1
X_1226_ _989_/A _994_/A _1410_/B vdd gnd NAND2X1
X_1861_ _1861_/A _1861_/B _1861_/C _1879_/B vdd gnd NAND3X1
X_1157_ _1165_/A _1166_/B _1166_/C _1161_/B vdd gnd NAND3X1
XFILL_0__1302_ gnd vdd FILL
X_1088_ _1088_/A _1088_/B _1088_/C _1111_/A vdd gnd NAND3X1
X_937_ _937_/A _953_/B _947_/B _962_/B vdd gnd AOI21X1
XFILL_0__1782_ gnd vdd FILL
X_1011_ _992_/A _997_/B _1039_/C vdd gnd NAND2X1
X_1775_ _1849_/A _974_/A _1848_/C _1776_/C vdd gnd OAI21X1
X_1844_ _1884_/A _1846_/B _1845_/C vdd gnd NAND2X1
X_1209_ _1210_/C _1210_/B _1210_/A _1231_/A vdd gnd NAND3X1
XFILL_0__1147_ gnd vdd FILL
X_1560_ _1562_/A _1598_/B _1561_/A vdd gnd NAND2X1
X_1758_ _1763_/B _1760_/B vdd gnd INVX1
X_1689_ vdd _963_/Y _950_/Y _1691_/CLK _942_/B vdd gnd DFFSR
X_1827_ _1829_/A _1829_/B _1828_/C vdd gnd NAND2X1
X_1491_ _1539_/A _1496_/A vdd gnd INVX1
XFILL_0__1748_ gnd vdd FILL
XFILL_0__1817_ gnd vdd FILL
X_1612_ _1867_/A _1613_/B vdd gnd INVX1
X_1474_ _1524_/C _1474_/B ABCmd_i[7] _1481_/C vdd gnd OAI21X1
X_1543_ _1621_/A _1621_/B _1589_/A vdd gnd NOR2X1
XFILL_0__1550_ gnd vdd FILL
XBUFX2_insert27 _1666_/Q _1274_/A vdd gnd BUFX2
X_1190_ _1190_/A _1190_/B _1190_/C _1202_/B vdd gnd NAND3X1
XFILL_0__1395_ gnd vdd FILL
X_1526_ _1572_/B _1527_/A vdd gnd INVX1
X_1388_ _1392_/B _1392_/A _1391_/C _1395_/C vdd gnd OAI21X1
X_1457_ _1457_/A _1457_/B _1511_/A _1461_/B vdd gnd AOI21X1
X_970_ _970_/A _972_/A vdd gnd INVX1
XFILL76350x50550 gnd vdd FILL
X_1242_ _1631_/C _1631_/A _1632_/A _1643_/C vdd gnd AOI21X1
X_1311_ _1321_/B _1416_/A _1470_/A vdd gnd AND2X2
X_1173_ _1175_/B _1175_/A _1175_/C _1244_/C vdd gnd AOI21X1
X_953_ _953_/A _953_/B _953_/Y vdd gnd NAND2X1
X_1509_ _1509_/A _1509_/B _1509_/C _1557_/B vdd gnd NAND3X1
X_1791_ _1843_/A _977_/A _1794_/B vdd gnd AND2X2
XFILL_0__1232_ gnd vdd FILL
X_1860_ _1867_/A _1861_/C vdd gnd INVX1
X_1225_ _1225_/A _1225_/B _1477_/A vdd gnd NAND2X1
X_1087_ _1146_/B _1111_/C _1111_/B _1105_/A vdd gnd OAI21X1
X_1156_ _1158_/A _1159_/C _1166_/B vdd gnd NAND2X1
X_936_ _936_/A _936_/B _953_/B vdd gnd NOR2X1
X_1010_ _993_/B _1232_/C vdd gnd INVX1
X_1774_ _1774_/A _1774_/B _1774_/C _1778_/A vdd gnd OAI21X1
X_1843_ _1843_/A _986_/A _1846_/B vdd gnd AND2X2
X_1208_ _1208_/A _999_/B _999_/A _1210_/B vdd gnd OAI21X1
XFILL_0__1077_ gnd vdd FILL
X_1139_ _1258_/C _1287_/B _1258_/A _1164_/A vdd gnd OAI21X1
XFILL_0_BUFX2_insert7 gnd vdd FILL
X_1826_ _1843_/A _983_/A _1829_/B vdd gnd AND2X2
XFILL_0__1833_ gnd vdd FILL
X_1490_ _1794_/A _986_/A _1539_/A vdd gnd NAND2X1
X_1757_ _1759_/A _997_/A _1757_/C _1763_/B vdd gnd AOI21X1
X_1688_ _1688_/D _1688_/CLK _1884_/A vdd gnd DFFPOSX1
XFILL_0__1480_ gnd vdd FILL
X_1611_ _1611_/A _1631_/C ABCmd_i[7] _1614_/A vdd gnd OAI21X1
X_1473_ _1525_/B _1525_/A _1474_/B vdd gnd NOR2X1
X_1542_ _1548_/A _1590_/D _1587_/B vdd gnd NOR2X1
XBUFX2_insert28 _1666_/Q _994_/A vdd gnd BUFX2
XBUFX2_insert17 _953_/Y _984_/B vdd gnd BUFX2
X_1809_ ABCmd_i[5] _1829_/A _1814_/C vdd gnd NAND2X1
X_1525_ _1525_/A _1525_/B _1525_/C _1527_/B vdd gnd AOI21X1
X_1387_ _1387_/A _1387_/B _1453_/A _1392_/A vdd gnd AOI21X1
X_1456_ _1456_/A _1456_/B _1457_/B vdd gnd NAND2X1
X_1241_ _1241_/A _1241_/B _1610_/A _1631_/A vdd gnd OAI21X1
X_1172_ _1246_/A _1297_/A _1246_/C _1175_/A vdd gnd NAND3X1
XFILL_0__1515_ gnd vdd FILL
X_1310_ _1310_/A _1397_/B _1310_/C _1416_/A vdd gnd NAND3X1
X_1439_ _1884_/A _1439_/B _1829_/A _1500_/B _1493_/D vdd gnd AOI22X1
X_1508_ _1516_/A _1515_/C vdd gnd INVX1
X_952_ _952_/A _962_/B _952_/C _957_/A vdd gnd OAI21X1
X_1790_ ABCmd_i[5] _1813_/A _1795_/C vdd gnd NAND2X1
XFILL_0__1162_ gnd vdd FILL
X_1224_ _1228_/A _1228_/B _1225_/B vdd gnd NOR2X1
X_1086_ _1090_/B _1090_/A _1111_/B vdd gnd AND2X2
XFILL_0_BUFX2_insert27 gnd vdd FILL
X_1155_ _1621_/B _1159_/B _1158_/A vdd gnd NOR2X1
X_935_ _956_/C _959_/C vdd gnd INVX1
X_1842_ ABCmd_i[5] ABCmd_i[4] _1847_/C vdd gnd NAND2X1
X_1773_ _995_/B _1773_/B _1868_/B _1774_/A vdd gnd OAI21X1
X_1207_ _998_/A _1410_/A _1228_/C _1228_/A _1210_/C vdd gnd OAI22X1
X_1138_ _1143_/B _1143_/A _1258_/A vdd gnd AND2X2
X_1069_ _1089_/C _1125_/B _1089_/A _1146_/B vdd gnd AOI21X1
XFILL_0__1763_ gnd vdd FILL
XFILL_0__965_ gnd vdd FILL
X_1756_ _1759_/A _997_/A _1848_/C _1757_/C vdd gnd OAI21X1
X_1687_ _1687_/D _1687_/CLK _1829_/A vdd gnd DFFPOSX1
X_1825_ _1884_/A _1882_/C vdd gnd INVX1
X_1610_ _1610_/A _1610_/B _1610_/C _1611_/A vdd gnd AOI21X1
XBUFX2_insert29 ABCmd_i[2] _970_/A vdd gnd BUFX2
X_1739_ _1868_/B _1739_/B _1739_/C _1740_/C vdd gnd NAND3X1
XBUFX2_insert18 _953_/Y _983_/B vdd gnd BUFX2
X_1808_ _1808_/A _1836_/A vdd gnd INVX1
X_1472_ _1572_/A _1525_/B vdd gnd INVX1
X_1541_ _1884_/A _1590_/A vdd gnd INVX1
XFILL76350x10950 gnd vdd FILL
XFILL_0__1531_ gnd vdd FILL
X_1524_ _1525_/C _1572_/B _1524_/C _1528_/A vdd gnd NOR3X1
XFILL_0__1600_ gnd vdd FILL
X_1455_ _1456_/B _1456_/A _1457_/A vdd gnd OR2X2
X_1386_ _1386_/A _1386_/B _1386_/C _1387_/B vdd gnd OAI21X1
X_1240_ _1632_/C _1631_/C vdd gnd INVX1
X_1171_ _1246_/B _1297_/C _1297_/B _1175_/B vdd gnd OAI21X1
XFILL_0__1445_ gnd vdd FILL
X_1507_ _1509_/C _1509_/B _1509_/A _1516_/A vdd gnd AOI21X1
X_1438_ _1442_/B _1441_/C vdd gnd INVX1
X_1369_ _1369_/A _1432_/A _1370_/A vdd gnd NOR2X1
X_951_ LoadA_i LoadB_i _962_/A _952_/A vdd gnd OAI21X1
XFILL76650x36150 gnd vdd FILL
XFILL_0__1092_ gnd vdd FILL
X_1223_ _998_/A _1410_/A _1228_/B vdd gnd NOR2X1
X_1085_ _1085_/A _1085_/B _1085_/C _1090_/B vdd gnd NAND3X1
X_1154_ _1621_/B _1159_/B _1158_/B _1166_/C vdd gnd OAI21X1
XFILL_0__981_ gnd vdd FILL
X_1772_ _1845_/A _974_/A _1772_/C _1845_/D _1774_/B vdd gnd AOI22X1
X_934_ _936_/B _934_/B _934_/Y vdd gnd NAND2X1
X_1841_ _1875_/A _1875_/B _1841_/C _1865_/B vdd gnd AOI21X1
XFILL_0__1213_ gnd vdd FILL
X_1206_ _965_/A _994_/B _994_/A _997_/B _1228_/A vdd gnd AOI22X1
X_1137_ _1250_/A _1137_/B _1137_/C _1143_/B vdd gnd NAND3X1
X_1068_ _1112_/A _1140_/C _1112_/B _1089_/C vdd gnd OAI21X1
XFILL_0__1693_ gnd vdd FILL
X_1755_ _1755_/A _1755_/B _1755_/C _1763_/A vdd gnd OAI21X1
X_1686_ _1686_/D _1687_/CLK _1813_/A vdd gnd DFFPOSX1
X_1824_ _1824_/A _1824_/B _1875_/B _1871_/C vdd gnd OAI21X1
XFILL_0__1127_ gnd vdd FILL
XFILL_0__1058_ gnd vdd FILL
XBUFX2_insert19 _953_/Y _972_/B vdd gnd BUFX2
X_1807_ _1836_/B _1807_/B _1859_/B vdd gnd NOR2X1
X_1471_ _1574_/A _1574_/B _1471_/C _1525_/A vdd gnd OAI21X1
X_1540_ _1559_/A _1599_/A vdd gnd INVX1
X_1738_ _1738_/A _1738_/B _1739_/C vdd gnd NAND2X1
X_1669_ _978_/Y _1680_/CLK _1669_/Q vdd gnd DFFPOSX1
X_1523_ _1567_/A _1573_/A _1572_/B vdd gnd NAND2X1
XFILL_0__1461_ gnd vdd FILL
X_1454_ _1454_/A _1454_/B _1511_/C _1489_/B _1461_/A vdd gnd AOI22X1
XFILL_0__1728_ gnd vdd FILL
X_1385_ _1385_/A _1449_/B _1385_/C _1387_/A vdd gnd NAND3X1
X_1170_ _1197_/B _1196_/C _1196_/A _1175_/C vdd gnd AOI21X1
X_1299_ _1299_/A _1299_/B _1340_/A _1304_/B vdd gnd AOI21X1
XFILL_0__1375_ gnd vdd FILL
X_1368_ _1368_/A _1368_/B _1424_/C _1370_/B vdd gnd NAND3X1
X_1506_ _1547_/B _1506_/B _1509_/A vdd gnd AND2X2
X_1437_ _1493_/A _1505_/C _1442_/B vdd gnd NOR2X1
X_950_ _950_/A _950_/B _950_/Y vdd gnd NAND2X1
X_1222_ _1228_/C _1225_/A vdd gnd INVX1
X_1084_ _1364_/B _1249_/A _1084_/C _1085_/C vdd gnd OAI21X1
X_1153_ _1159_/C _1158_/B vdd gnd INVX1
X_1771_ _995_/B _1773_/B _1772_/C vdd gnd NAND2X1
X_933_ _936_/A _937_/A _934_/B vdd gnd NOR2X1
X_1840_ _1869_/A _1865_/A vdd gnd INVX1
XFILL_0__1143_ gnd vdd FILL
X_1205_ _989_/A _997_/A _1228_/C vdd gnd NAND2X1
X_1067_ _1114_/A _1829_/A _1067_/C _1813_/A _1112_/A vdd gnd AOI22X1
X_1136_ _1364_/B _1343_/A _1136_/C _1137_/C vdd gnd OAI21X1
X_1754_ _994_/B _1754_/B _1868_/B _1755_/A vdd gnd OAI21X1
X_1685_ _1685_/D _1688_/CLK _1794_/A vdd gnd DFFPOSX1
X_1823_ _1823_/A _1823_/B _1867_/A vdd gnd NAND2X1
X_1119_ _1274_/A _1884_/A _1120_/B vdd gnd NAND2X1
XFILL_0__946_ gnd vdd FILL
XFILL_0__1744_ gnd vdd FILL
XFILL_0__1813_ gnd vdd FILL
XFILL75750x36150 gnd vdd FILL
X_1470_ _1470_/A _1470_/B _1574_/B vdd gnd NAND2X1
X_1668_ _975_/Y _1687_/CLK _1668_/Q vdd gnd DFFPOSX1
X_1737_ _1868_/A _1845_/A _965_/A _1738_/A vdd gnd OAI21X1
X_1806_ _1820_/B _1820_/A _1807_/B vdd gnd NOR2X1
X_1599_ _1599_/A _1599_/B _1599_/C _1600_/C vdd gnd OAI21X1
XFILL76650x64950 gnd vdd FILL
XFILL_0__1391_ gnd vdd FILL
XFILL_0__1658_ gnd vdd FILL
XFILL_0__1589_ gnd vdd FILL
X_1384_ _1420_/B _1453_/C _1420_/A _1392_/B vdd gnd AOI21X1
X_1453_ _1453_/A _1453_/B _1453_/C _1520_/C vdd gnd OAI21X1
X_1522_ _1522_/A _1537_/B _1522_/C _1567_/A vdd gnd NAND3X1
X_1505_ _1621_/A _1550_/B _1505_/C _1506_/B vdd gnd OAI21X1
X_1436_ _1884_/A _1500_/B _1505_/C vdd gnd NAND2X1
X_1367_ _1424_/A _1367_/B _1367_/C _1370_/C vdd gnd NAND3X1
X_1298_ _1298_/A _1298_/B _1340_/C _1383_/B _1304_/A vdd gnd AOI22X1
XFILL_0_BUFX2_insert19 gnd vdd FILL
X_1221_ _993_/B _1231_/A _1221_/C _1529_/B vdd gnd NAND3X1
X_1152_ _1152_/A _1152_/B _1152_/C _1152_/D _1159_/C vdd gnd AOI22X1
X_1083_ _991_/B _1343_/A _1083_/C _1085_/B vdd gnd OAI21X1
X_1419_ _1462_/A _1521_/A vdd gnd INVX1
XFILL_0__1426_ gnd vdd FILL
XFILL76350x61350 gnd vdd FILL
X_1770_ _1843_/A _974_/A _1773_/B vdd gnd AND2X2
X_932_ _953_/A _937_/A vdd gnd INVX2
X_1204_ _965_/A _997_/B _1410_/A vdd gnd NAND2X1
X_1899_ _1899_/A ACC_o[5] vdd gnd BUFX2
X_1066_ _1066_/A _1279_/A _1140_/C vdd gnd NOR2X1
XFILL_0__1073_ gnd vdd FILL
X_1135_ _991_/B _1499_/A _1152_/B _1137_/B vdd gnd OAI21X1
X_1684_ _1684_/D _1691_/CLK _995_/B vdd gnd DFFPOSX1
X_1753_ _1845_/A _997_/A _1753_/C _1845_/D _1755_/B vdd gnd AOI22X1
X_1822_ _1836_/C _1824_/B _1823_/B vdd gnd NAND2X1
X_1049_ _1099_/C _1049_/B _1193_/A vdd gnd NAND2X1
X_1118_ _1271_/A _1271_/B _1277_/C _1142_/B vdd gnd NAND3X1
X_1736_ ABCmd_i[1] _1736_/B ABCmd_i[0] _1738_/B vdd gnd MUX2X1
X_1667_ _972_/Y _1682_/CLK _997_/A vdd gnd DFFPOSX1
X_1805_ _1805_/A _1820_/B vdd gnd INVX1
XFILL_0__1108_ gnd vdd FILL
X_1598_ _1599_/C _1598_/B _1598_/C _1601_/B vdd gnd NAND3X1
X_1383_ _1383_/A _1383_/B _1383_/C _1391_/C vdd gnd AOI21X1
X_1452_ _1520_/B _1520_/A _1461_/C _1459_/C vdd gnd NAND3X1
X_1521_ _1521_/A _1521_/B _1521_/C _1522_/C vdd gnd OAI21X1
X_1719_ _1734_/A _1741_/A _1720_/B vdd gnd NOR2X1
XFILL_0__1511_ gnd vdd FILL
X_1504_ _980_/A _1550_/B vdd gnd INVX1
XFILL_0__1709_ gnd vdd FILL
X_1297_ _1297_/A _1297_/B _1297_/C _1303_/C vdd gnd AOI21X1
X_1366_ _1432_/A _1369_/A _1366_/C _1366_/D _1385_/A vdd gnd OAI22X1
X_1435_ _1829_/A _1439_/B _1493_/A vdd gnd NAND2X1
X_1220_ _1232_/A _1221_/C vdd gnd INVX1
X_1151_ _1166_/A _1165_/A vdd gnd INVX1
X_1082_ _1152_/C _1152_/D _1082_/C _1090_/A vdd gnd NAND3X1
XFILL_0__1356_ gnd vdd FILL
X_1418_ _1418_/A _1418_/B _1418_/C _1462_/A vdd gnd OAI21X1
X_1349_ _1349_/A _1349_/B _1418_/B vdd gnd NOR2X1
X_931_ _942_/B _936_/B vdd gnd INVX1
X_1203_ _1203_/A _1203_/B _999_/C _1210_/A vdd gnd NAND3X1
X_1065_ _1067_/C _1829_/A _1279_/A vdd gnd NAND2X1
X_1134_ _1794_/A _1499_/A vdd gnd INVX1
XFILL_0__961_ gnd vdd FILL
X_1898_ _1898_/A ACC_o[4] vdd gnd BUFX2
X_1752_ _994_/B _1754_/B _1753_/C vdd gnd NAND2X1
X_1683_ _1683_/D _1691_/CLK _994_/B vdd gnd DFFPOSX1
X_1821_ _1824_/A _1836_/C vdd gnd INVX1
XFILL_0__1124_ gnd vdd FILL
X_1048_ _1048_/A _1048_/B _1048_/C _1192_/B vdd gnd AOI21X1
X_1117_ _1277_/B _1271_/B vdd gnd INVX1
X_1735_ _970_/A _1848_/C _1740_/B _1741_/B vdd gnd OAI21X1
X_1804_ _1858_/A _1804_/B _1804_/C _1820_/A vdd gnd OAI21X1
X_1666_ _969_/Y _1682_/CLK _1666_/Q vdd gnd DFFPOSX1
XFILL_0__1038_ gnd vdd FILL
X_1597_ _1600_/A _1600_/B _1598_/C vdd gnd NAND2X1
XFILL_0__927_ gnd vdd FILL
X_1382_ _1382_/A _1386_/B _1382_/C _1383_/C vdd gnd NOR3X1
X_1520_ _1520_/A _1520_/B _1520_/C _1521_/B vdd gnd AOI21X1
X_1451_ _1511_/C _1489_/B _1489_/A _1520_/A vdd gnd NAND3X1
X_1649_ _989_/A _1659_/B _1650_/C vdd gnd NAND2X1
X_1718_ _1718_/A _1857_/A vdd gnd INVX1
XFILL_0__1372_ gnd vdd FILL
XFILL_0__1441_ gnd vdd FILL
XFILL_0__1639_ gnd vdd FILL
X_1503_ _1545_/B _1547_/B vdd gnd INVX1
X_1296_ _1336_/A _1336_/B _1336_/C _1401_/A vdd gnd NAND3X1
X_1434_ _1493_/C _1441_/A vdd gnd INVX1
X_1365_ _1367_/B _1367_/C _1424_/A _1366_/D vdd gnd AOI21X1
X_1150_ _989_/A _986_/A _1166_/A vdd gnd NAND2X1
X_1417_ _1573_/C _1471_/C vdd gnd INVX1
X_1081_ _991_/B _1343_/A _1099_/B _1152_/C vdd gnd OAI21X1
XFILL_0__1286_ gnd vdd FILL
X_930_ _930_/A _947_/B vdd gnd INVX1
XFILL75450x7350 gnd vdd FILL
X_1348_ _1349_/B _1349_/A _1350_/B vdd gnd AND2X2
X_1279_ _1279_/A _1369_/A _1279_/C _1352_/A vdd gnd OAI21X1
X_1202_ _1202_/A _1202_/B _1215_/A _1234_/B vdd gnd NAND3X1
X_1133_ _1133_/A _1133_/B _1250_/C _1143_/A vdd gnd NAND3X1
X_1064_ _1140_/A _1140_/B _1125_/A _1125_/B vdd gnd NAND3X1
X_1897_ _1897_/A ACC_o[3] vdd gnd BUFX2
X_1820_ _1820_/A _1820_/B _1836_/A _1824_/B vdd gnd AOI21X1
X_1751_ ABCmd_i[0] _1751_/B _1754_/B vdd gnd NOR2X1
X_1682_ _1682_/D _1682_/CLK _997_/B vdd gnd DFFPOSX1
XFILL_0__1887_ gnd vdd FILL
XFILL_0__1054_ gnd vdd FILL
X_1047_ _1047_/A _1047_/B _1047_/C _1192_/A vdd gnd AOI21X1
X_1116_ _997_/A _1813_/A _1277_/B vdd gnd NAND2X1
X_1734_ _1734_/A _1740_/B vdd gnd INVX1
X_1665_ _966_/Y _1682_/CLK _1665_/Q vdd gnd DFFPOSX1
XFILL_0__1810_ gnd vdd FILL
X_1803_ ABCmd_i[6] _1857_/B _1804_/B vdd gnd NAND2X1
X_1596_ _1619_/B _1619_/A _1600_/B vdd gnd OR2X2
XFILL_0__1724_ gnd vdd FILL
X_1381_ _1465_/B _1465_/A _1465_/C _1466_/C vdd gnd NAND3X1
X_1450_ _1450_/A _1450_/B _1456_/B _1511_/C vdd gnd NAND3X1
XFILL_0__1655_ gnd vdd FILL
X_1717_ _1717_/A _1717_/B _1718_/A vdd gnd NAND2X1
X_1579_ _1610_/C _1581_/B vdd gnd INVX1
X_1648_ _1648_/A _949_/A _1648_/C _1648_/D _1680_/D vdd gnd AOI22X1
XFILL_0__1569_ gnd vdd FILL
X_1364_ _1548_/A _1364_/B _1364_/C _1367_/C vdd gnd OAI21X1
X_1502_ _1502_/A _1593_/A _1545_/B vdd gnd NOR2X1
X_1295_ _1383_/B _1340_/C _1383_/A _1336_/B vdd gnd NAND3X1
X_1433_ _1813_/A _980_/A _1493_/C vdd gnd NAND2X1
X_1080_ _992_/A _994_/B _1099_/B vdd gnd NAND2X1
X_1347_ _1347_/A _1418_/C _1347_/C _1377_/A vdd gnd NAND3X1
X_1278_ _1278_/A _1279_/C vdd gnd INVX1
X_1416_ _1416_/A _1416_/B _1416_/C _1573_/C vdd gnd AOI21X1
X_1201_ _1201_/A _1201_/B _1241_/A _1643_/B vdd gnd AOI21X1
X_1896_ _1896_/A ACC_o[2] vdd gnd BUFX2
X_989_ _989_/A _991_/A vdd gnd INVX1
XFILL_0__1406_ gnd vdd FILL
X_1063_ _1112_/B _1140_/B vdd gnd INVX1
X_1132_ _1250_/B _1133_/B vdd gnd INVX1
XFILL76350x3750 gnd vdd FILL
XFILL_0__1337_ gnd vdd FILL
XFILL76050x7350 gnd vdd FILL
X_1681_ _1681_/D _1691_/CLK _989_/A vdd gnd DFFPOSX1
X_1750_ _997_/A _1751_/B vdd gnd INVX1
X_1046_ _1193_/B _1193_/C _1192_/C _1052_/B vdd gnd NAND3X1
X_1115_ _1277_/A _1271_/A vdd gnd INVX1
XFILL_0__942_ gnd vdd FILL
X_1879_ ABCmd_i[6] _1879_/B _1879_/C _1890_/B vdd gnd NAND3X1
XFILL_0__1740_ gnd vdd FILL
X_1733_ _1733_/A _1733_/B _1764_/C vdd gnd NAND2X1
X_1802_ _1802_/A _1802_/B _1802_/C _1857_/B vdd gnd OAI21X1
X_1664_ _987_/A _1664_/B _1664_/C _1688_/D vdd gnd OAI21X1
X_1029_ _1048_/B _1048_/A _1048_/C _1193_/B vdd gnd NAND3X1
X_1595_ _1619_/A _1619_/B _1600_/A vdd gnd NAND2X1
X_1380_ _1453_/C _1420_/B _1420_/A _1465_/B vdd gnd NAND3X1
X_1716_ ABCmd_i[5] _1716_/B _1716_/C _1717_/A vdd gnd OAI21X1
XFILL_0__1585_ gnd vdd FILL
X_1647_ _1647_/A _937_/A _949_/A _1648_/D vdd gnd AOI21X1
X_1578_ _952_/C _1578_/B _1578_/C _1585_/C vdd gnd NAND3X1
XFILL_0__1019_ gnd vdd FILL
X_1363_ _1621_/A _991_/B _1363_/C _1367_/B vdd gnd OAI21X1
X_1501_ _1884_/A _980_/A _1593_/A vdd gnd NAND2X1
X_1294_ _1382_/A _1386_/B _1382_/C _1383_/B vdd gnd OAI21X1
X_1432_ _1432_/A _1432_/B _1449_/A vdd gnd NAND2X1
XFILL76050x28950 gnd vdd FILL
XFILL_0__1422_ gnd vdd FILL
X_1415_ _1470_/A _1470_/B _1566_/A _1469_/A vdd gnd NAND3X1
X_1346_ _1349_/B _1349_/A _1347_/C vdd gnd OR2X2
X_1277_ _1277_/A _1277_/B _1277_/C _1373_/B vdd gnd OAI21X1
XFILL76650x50550 gnd vdd FILL
X_988_ _988_/A _988_/Y vdd gnd INVX1
X_1895_ _1895_/A ACC_o[1] vdd gnd BUFX2
X_1131_ _1131_/A _1794_/A _992_/A _995_/B _1250_/B vdd gnd AOI22X1
XFILL_0__1267_ gnd vdd FILL
X_1062_ _997_/A _1794_/A _1112_/B vdd gnd NAND2X1
X_1200_ _1244_/C _1307_/B _1307_/A _1201_/A vdd gnd OAI21X1
X_1329_ _1329_/A _1329_/B _1329_/C _1330_/B vdd gnd OAI21X1
X_1680_ _1680_/D _1680_/CLK _1901_/A vdd gnd DFFPOSX1
X_1114_ _1114_/A _1884_/A _1274_/A _1829_/A _1277_/A vdd gnd AOI22X1
X_1878_ _1878_/A _1878_/B _1890_/A _1892_/A vdd gnd OAI21X1
X_1045_ _1049_/B _1099_/C _1192_/C vdd gnd AND2X2
X_1732_ _1732_/A _1732_/B _1747_/B _1733_/A vdd gnd MUX2X1
X_1801_ _1801_/A _1801_/B _1802_/A vdd gnd NOR2X1
X_1663_ _1884_/A _1664_/B _1664_/C vdd gnd NAND2X1
XFILL_0__1868_ gnd vdd FILL
X_1028_ _1055_/A _1070_/C _1055_/B _1048_/A vdd gnd OAI21X1
X_1594_ _1594_/A _1619_/C _1619_/B vdd gnd NAND2X1
XFILL_0__1104_ gnd vdd FILL
X_1715_ _1716_/C _1720_/A _1717_/B vdd gnd OR2X2
X_1646_ _987_/A _1646_/B _1646_/C _1647_/A vdd gnd OAI21X1
X_1577_ ABCmd_i[7] _1892_/A _1578_/B vdd gnd OR2X2
X_1362_ _1829_/A _1621_/A vdd gnd INVX2
X_1500_ _1829_/A _1500_/B _1502_/A vdd gnd NAND2X1
X_1293_ _1339_/A _1339_/B _1339_/C _1340_/C vdd gnd NAND3X1
X_1431_ _1454_/B _1454_/A _1511_/A vdd gnd NAND2X1
XFILL_0__1705_ gnd vdd FILL
X_1629_ _1629_/A _1629_/B _1629_/C _1630_/C vdd gnd OAI21X1
X_1414_ _942_/B _942_/C _1896_/A _1482_/C vdd gnd OAI21X1
X_1345_ _1349_/A _1349_/B _1418_/C vdd gnd NAND2X1
X_1276_ _1373_/A _1352_/B _1289_/A vdd gnd NAND2X1
XFILL_0__1352_ gnd vdd FILL
X_1894_ _988_/A ACC_o[0] vdd gnd BUFX2
X_987_ _987_/A _987_/B _987_/C _987_/Y vdd gnd OAI21X1
XFILL_0__1197_ gnd vdd FILL
X_1130_ _1152_/B _1136_/C _1250_/C vdd gnd NAND2X1
X_1061_ _1061_/A _1548_/A _1120_/A _1140_/A vdd gnd OAI21X1
X_1328_ _1857_/A ABCmd_i[7] _960_/C _1329_/B vdd gnd OAI21X1
X_1259_ _980_/A _995_/B _1344_/A vdd gnd NAND2X1
XFILL_0__1120_ gnd vdd FILL
X_1877_ _1877_/A _1877_/B _1890_/A vdd gnd AND2X2
X_1044_ _1044_/A _1044_/B _1044_/C _1049_/B vdd gnd NAND3X1
X_1113_ _1114_/A _1884_/A _1432_/A _1277_/C vdd gnd NAND3X1
X_1731_ _1759_/A _1848_/C _1732_/B _1732_/A vdd gnd OAI21X1
X_1662_ _984_/A _1662_/B _1662_/C _1687_/D vdd gnd OAI21X1
XFILL_0__1798_ gnd vdd FILL
X_1800_ _1800_/A _1804_/C _1805_/A _1836_/B vdd gnd AOI21X1
XFILL_0__1034_ gnd vdd FILL
X_1027_ _1027_/A _1066_/A _1070_/C vdd gnd NOR2X1
X_1593_ _1593_/A _1593_/B _1593_/C _1594_/A vdd gnd OAI21X1
X_1714_ _1741_/A _1734_/A _1720_/C _1716_/C vdd gnd OAI21X1
X_1645_ _1879_/C _987_/A _1646_/C vdd gnd NAND2X1
X_1576_ _1576_/A _1576_/B ABCmd_i[7] _1578_/C vdd gnd OAI21X1
XFILL76650x7350 gnd vdd FILL
X_1430_ _1487_/B _1430_/B _1487_/A _1454_/B vdd gnd OAI21X1
XFILL_0__1635_ gnd vdd FILL
X_1628_ _1639_/C _1629_/C vdd gnd INVX1
X_1292_ _1298_/A _1298_/B _1383_/A vdd gnd AND2X2
X_1361_ _1424_/C _1368_/B _1368_/A _1366_/C vdd gnd AOI21X1
X_1559_ _1559_/A _1599_/C _1559_/C _1598_/B vdd gnd NAND3X1
XFILL76650x10950 gnd vdd FILL
X_1413_ _1413_/A _949_/A _1413_/C _1413_/D _1674_/D vdd gnd AOI22X1
XFILL_0__1282_ gnd vdd FILL
X_1275_ _1432_/B _1432_/A _1278_/A _1373_/A vdd gnd AOI21X1
X_1344_ _1344_/A _1344_/B _1344_/C _1349_/B vdd gnd OAI21X1
XFILL76350x57750 gnd vdd FILL
X_986_ _986_/A _987_/B _987_/C vdd gnd NAND2X1
XFILL_0__1403_ gnd vdd FILL
X_1060_ _1114_/A _1829_/A _1120_/A vdd gnd NAND2X1
X_1327_ _965_/A _989_/A _987_/A _1329_/A vdd gnd AOI21X1
X_1893_ _1893_/A _1893_/B _1893_/Y vdd gnd NAND2X1
X_1189_ _993_/Y _1189_/B _1202_/A vdd gnd AND2X2
XFILL75750x150 gnd vdd FILL
X_1258_ _1258_/A _1258_/B _1258_/C _1382_/C vdd gnd AOI21X1
XFILL_0__1050_ gnd vdd FILL
X_969_ _969_/A _987_/B _969_/C _969_/Y vdd gnd OAI21X1
XFILL_0__1883_ gnd vdd FILL
X_1876_ _1876_/A _1876_/B _1876_/C _1877_/A vdd gnd OAI21X1
XFILL_0__1317_ gnd vdd FILL
X_1043_ _1364_/B _1159_/B _1152_/A _1044_/C vdd gnd OAI21X1
XFILL_0__1248_ gnd vdd FILL
X_1112_ _1112_/A _1112_/B _1125_/A _1142_/A vdd gnd OAI21X1
X_1730_ _1747_/A _1732_/B vdd gnd INVX1
X_1661_ _1829_/A _1662_/B _1662_/C vdd gnd NAND2X1
X_1592_ _1592_/A _1593_/C _1619_/C vdd gnd OR2X2
X_1859_ _1859_/A _1859_/B _1863_/B vdd gnd NOR2X1
X_1026_ _995_/A _1813_/A _1066_/A vdd gnd NAND2X1
XFILL_0__1720_ gnd vdd FILL
XFILL_0__1651_ gnd vdd FILL
XFILL76050x54150 gnd vdd FILL
X_1713_ _1881_/A _1734_/A _1741_/A _1720_/C vdd gnd OAI21X1
X_1009_ _1016_/B _999_/Y _1016_/A _1215_/A vdd gnd NAND3X1
X_1575_ _1604_/C _1604_/B _1604_/A _1576_/A vdd gnd AOI21X1
X_1644_ _1644_/A _1644_/B _1646_/B vdd gnd NAND2X1
XFILL_0__1565_ gnd vdd FILL
X_1291_ _1340_/A _1299_/B _1299_/A _1336_/A vdd gnd NAND3X1
XFILL_0__1496_ gnd vdd FILL
X_1360_ _1424_/B _1368_/B vdd gnd INVX1
X_1627_ _1627_/A _1627_/B _1627_/C _1629_/B vdd gnd AOI21X1
X_1489_ _1489_/A _1489_/B _1489_/C _1516_/C vdd gnd AOI21X1
X_1558_ _1599_/B _1559_/C vdd gnd INVX1
XFILL_0_CLKBUF1_insert15 gnd vdd FILL
X_1412_ _1412_/A _937_/A _949_/A _1413_/D vdd gnd AOI21X1
X_1343_ _1343_/A _1621_/B _1349_/A vdd gnd NOR2X1
X_1274_ _1274_/A _1884_/A _997_/A _1829_/A _1278_/A vdd gnd AOI22X1
X_985_ ABCmd_i[7] _987_/A vdd gnd INVX4
X_1326_ _987_/A _1326_/B _1326_/C _1329_/C vdd gnd OAI21X1
X_1188_ _1190_/C _1190_/A _1190_/B _1212_/A vdd gnd AOI21X1
XFILL_0__1333_ gnd vdd FILL
X_1892_ _1892_/A _1892_/B _1893_/B vdd gnd NAND2X1
X_1257_ _1298_/B _1298_/A _1340_/A vdd gnd NAND2X1
X_968_ _994_/A _987_/B _969_/C vdd gnd NAND2X1
X_1875_ _1875_/A _1875_/B _1875_/C _1876_/B vdd gnd AOI21X1
X_1111_ _1111_/A _1111_/B _1111_/C _1164_/C vdd gnd AOI21X1
X_1042_ _997_/B _1159_/B vdd gnd INVX1
XFILL_0__1178_ gnd vdd FILL
X_1309_ _1402_/A _1402_/B _1401_/A _1397_/B vdd gnd NAND3X1
X_1660_ _981_/A _1662_/B _1660_/C _1686_/D vdd gnd OAI21X1
X_1591_ _1591_/A _1640_/C _1593_/C vdd gnd NAND2X1
XFILL75750x10950 gnd vdd FILL
X_1789_ _1789_/A _1789_/B _1789_/C _1804_/C vdd gnd AOI21X1
X_1858_ _1858_/A _1858_/B _1859_/A vdd gnd NAND2X1
X_1025_ _1070_/A _1070_/B _1055_/C _1048_/B vdd gnd NAND3X1
X_1712_ _970_/A _1848_/C _1881_/A vdd gnd NOR2X1
XFILL_0__1779_ gnd vdd FILL
XFILL_0__1848_ gnd vdd FILL
XFILL_0__1015_ gnd vdd FILL
XFILL_0__1581_ gnd vdd FILL
X_1643_ _1643_/A _1643_/B _1643_/C _1644_/A vdd gnd OAI21X1
X_1574_ _1574_/A _1574_/B _1574_/C _1604_/C vdd gnd OAI21X1
X_1008_ _1186_/A _1186_/B _1187_/A _1016_/B vdd gnd OAI21X1
X_1290_ _1382_/A _1386_/B _1339_/C _1299_/B vdd gnd OAI21X1
X_1626_ _1626_/A _1626_/B _1627_/C vdd gnd OR2X2
X_1488_ _1517_/A _1514_/A vdd gnd INVX1
X_1557_ _1557_/A _1557_/B _1599_/C vdd gnd OR2X2
X_1411_ _1411_/A _1411_/B _1411_/C _1412_/A vdd gnd OAI21X1
XFILL_0__1616_ gnd vdd FILL
X_1609_ _1639_/A _1609_/B _1609_/C _1615_/C vdd gnd NAND3X1
X_1342_ _1418_/A _1347_/A vdd gnd INVX1
X_1273_ _1369_/A _1432_/B vdd gnd INVX1
X_984_ _984_/A _984_/B _984_/C _984_/Y vdd gnd OAI21X1
X_1325_ _1325_/A _960_/C _1326_/C vdd gnd NOR2X1
X_1891_ _1891_/A _1891_/B _1892_/B vdd gnd AND2X2
X_1256_ _1338_/B _1256_/B _1338_/A _1298_/B vdd gnd OAI21X1
XFILL_0__1263_ gnd vdd FILL
XFILL76050x39750 gnd vdd FILL
X_1187_ _1187_/A _1187_/B _1187_/C _1190_/C vdd gnd NAND3X1
X_967_ ABCmd_i[1] _969_/A vdd gnd INVX1
X_1041_ _991_/B _1249_/A _993_/A _1044_/B vdd gnd OAI21X1
X_1110_ _1197_/A _1196_/B _1197_/C _1176_/C vdd gnd OAI21X1
X_1874_ _1874_/A _1874_/B _1875_/C vdd gnd NAND2X1
X_1239_ _1610_/A _1610_/B _1610_/C _1632_/C vdd gnd NAND3X1
X_1308_ _1337_/A _1308_/B _1308_/C _1310_/A vdd gnd NAND3X1
XFILL76650x61350 gnd vdd FILL
XFILL_0__1100_ gnd vdd FILL
XFILL76050x14550 gnd vdd FILL
X_1788_ _1788_/A _1789_/C vdd gnd INVX1
X_1857_ _1857_/A _1857_/B _1858_/B vdd gnd NOR2X1
XFILL_0__1864_ gnd vdd FILL
X_1024_ _1055_/B _1070_/B vdd gnd INVX1
X_1590_ _1590_/A _1621_/B _1621_/A _1590_/D _1591_/A vdd gnd OAI22X1
X_1711_ _1711_/A _970_/A _1711_/C _1734_/A vdd gnd AOI21X1
X_1642_ _1642_/A _1642_/B _1642_/C _1644_/B vdd gnd NAND3X1
X_1573_ _1573_/A _1573_/B _1573_/C _1574_/C vdd gnd AOI21X1
X_1007_ _998_/B _1027_/A _1186_/B vdd gnd NOR2X1
XFILL_0__1701_ gnd vdd FILL
X_1625_ _1639_/C _1639_/B _1639_/A _1630_/B vdd gnd NAND3X1
X_1487_ _1487_/A _1487_/B _1487_/C _1517_/A vdd gnd OAI21X1
X_1556_ _1599_/B _1556_/B _1599_/A _1562_/A vdd gnd OAI21X1
X_1410_ _1410_/A _1410_/B ABCmd_i[7] _1411_/A vdd gnd OAI21X1
XFILL_0__1546_ gnd vdd FILL
X_1341_ _994_/B _986_/A _1418_/A vdd gnd NAND2X1
X_1272_ _1884_/A _997_/A _1369_/A vdd gnd NAND2X1
X_1608_ _1608_/A _1641_/C _1609_/B vdd gnd AND2X2
X_1539_ _1539_/A _1539_/B _1539_/C _1559_/A vdd gnd OAI21X1
X_983_ _983_/A _983_/B _984_/C vdd gnd NAND2X1
X_1890_ _1890_/A _1890_/B _1890_/C _1893_/A vdd gnd NAND3X1
XFILL_0__1193_ gnd vdd FILL
X_1324_ ABCmd_i[7] _1820_/A _1325_/A vdd gnd NOR2X1
X_1186_ _1186_/A _1186_/B _1186_/C _1190_/A vdd gnd OAI21X1
X_1255_ _1255_/A _1255_/B _1338_/B vdd gnd NOR2X1
X_966_ _966_/A _983_/B _966_/C _966_/Y vdd gnd OAI21X1
X_1040_ _1040_/A _1040_/B _1040_/C _1099_/C vdd gnd NAND3X1
X_1873_ _1873_/A _1876_/C vdd gnd INVX1
X_1238_ _1238_/A _1238_/B _1238_/C _1610_/B vdd gnd NAND3X1
X_1307_ _1307_/A _1307_/B _1307_/C _1310_/C vdd gnd OAI21X1
X_1169_ _1176_/B _1176_/A _1176_/C _1307_/B vdd gnd AOI21X1
X_949_ _949_/A _949_/B _949_/C _960_/A _950_/A vdd gnd AOI22X1
XFILL_0__1794_ gnd vdd FILL
XFILL_0__996_ gnd vdd FILL
XFILL_0__1228_ gnd vdd FILL
XFILL_0__1030_ gnd vdd FILL
X_1023_ _997_/A _995_/B _1055_/B vdd gnd NAND2X1
X_1787_ _1787_/A _1787_/B _1789_/A vdd gnd NAND2X1
X_1856_ _1886_/A _1886_/C _1879_/C vdd gnd NAND2X1
X_1710_ _1711_/A _970_/A _1848_/C _1711_/C vdd gnd OAI21X1
X_1641_ _1641_/A _1641_/B _1641_/C _1648_/C vdd gnd OAI21X1
X_1572_ _1572_/A _1572_/B _1572_/C _1604_/B vdd gnd OAI21X1
X_1839_ _1861_/A _1861_/B _1867_/B vdd gnd NAND2X1
X_1006_ _1187_/B _1186_/C _1187_/C _1016_/A vdd gnd NAND3X1
XFILL_0__1829_ gnd vdd FILL
X_1624_ _1624_/A _1624_/B _1639_/C vdd gnd NAND2X1
XFILL_0__1631_ gnd vdd FILL
X_1486_ _1567_/B _1525_/C vdd gnd INVX1
XFILL_0__1562_ gnd vdd FILL
X_1555_ _1555_/A _1592_/A _1555_/C _1599_/B vdd gnd AOI21X1
XFILL_0__1476_ gnd vdd FILL
X_1340_ _1340_/A _1340_/B _1340_/C _1465_/C vdd gnd OAI21X1
X_1271_ _1271_/A _1271_/B _1271_/C _1352_/B vdd gnd AOI21X1
X_1607_ _1626_/B _1617_/A _1608_/A vdd gnd OR2X2
X_1538_ _1562_/C _1561_/B vdd gnd INVX1
X_1469_ _1469_/A _1471_/C _1572_/A _1524_/C vdd gnd AOI21X1
XFILL75450x150 gnd vdd FILL
X_982_ ABCmd_i[6] _984_/A vdd gnd INVX1
X_1185_ _1203_/B _1203_/A _1208_/A _1190_/B vdd gnd AOI21X1
X_1323_ _1323_/A _1399_/A _1326_/B vdd gnd AND2X2
X_1254_ _1255_/B _1255_/A _1256_/B vdd gnd AND2X2
X_965_ _965_/A _983_/B _966_/C vdd gnd NAND2X1
X_1872_ _1873_/A _1872_/B _1872_/C _1877_/B vdd gnd NAND3X1
XFILL_0__1313_ gnd vdd FILL
X_1306_ _1306_/A _1306_/B _1306_/C _1321_/B vdd gnd OAI21X1
XFILL_0__1244_ gnd vdd FILL
X_1237_ _993_/Y _1237_/B _1316_/A _1238_/B vdd gnd NAND3X1
X_1099_ _1099_/A _1099_/B _1099_/C _1101_/A vdd gnd OAI21X1
X_1168_ _1246_/B _1297_/C _1246_/A _1176_/B vdd gnd OAI21X1
X_948_ _960_/B _952_/C _948_/C _949_/C vdd gnd OAI21X1
X_1022_ _1055_/A _1070_/A vdd gnd INVX1
X_1786_ _1786_/A _1786_/B _1786_/C _1800_/A vdd gnd NAND3X1
X_1855_ _1869_/A _1874_/A _1864_/C _1886_/A vdd gnd NAND3X1
XFILL_0__1158_ gnd vdd FILL
XFILL_0__1089_ gnd vdd FILL
XFILL76350x43350 gnd vdd FILL
X_1838_ _1875_/B _1874_/B _1875_/A _1861_/A vdd gnd NAND3X1
X_1005_ _1186_/A _1187_/B vdd gnd INVX1
X_1640_ _1640_/A _1640_/B _1640_/C _1641_/A vdd gnd OAI21X1
X_1571_ _1573_/A _1573_/B _1572_/C vdd gnd NAND2X1
X_1769_ ABCmd_i[5] _1794_/A _1774_/C vdd gnd NAND2X1
X_1485_ _1485_/A _960_/C _1606_/A _1528_/C vdd gnd OAI21X1
X_1623_ _1640_/A _1640_/B _1624_/A vdd gnd NAND2X1
X_1554_ _1557_/B _1557_/A _1556_/B vdd gnd NOR2X1
XFILL_0__1492_ gnd vdd FILL
.ends

