magic
tech scmos
magscale 1 3
timestamp 1569140870
<< checkpaint >>
rect -50 -50 300 300
<< ndiffusion >>
rect 75 75 175 175
<< metal1 >>
rect 75 75 175 175
use ntap_CDNS_7230122529123  ntap_CDNS_7230122529123_0
timestamp 1569140870
transform 1 0 72 0 1 72
box 4 4 102 102
use ptap_ring_ndiode_CDNS_7230122529121  ptap_ring_ndiode_CDNS_7230122529121_0
timestamp 1569140870
transform 1 0 0 0 1 0
box 10 10 240 240
<< end >>
